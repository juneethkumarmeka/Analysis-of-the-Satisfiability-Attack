module basic_2500_25000_3000_8_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nand U0 (N_0,In_1627,In_1691);
or U1 (N_1,In_1349,In_613);
nand U2 (N_2,In_703,In_318);
nand U3 (N_3,In_1625,In_1571);
and U4 (N_4,In_347,In_1637);
xor U5 (N_5,In_1404,In_548);
and U6 (N_6,In_1649,In_1333);
xnor U7 (N_7,In_711,In_1476);
nand U8 (N_8,In_2377,In_596);
nor U9 (N_9,In_1165,In_1825);
and U10 (N_10,In_1918,In_1018);
nor U11 (N_11,In_453,In_499);
xor U12 (N_12,In_212,In_198);
nand U13 (N_13,In_1535,In_1143);
nand U14 (N_14,In_2018,In_1945);
xor U15 (N_15,In_1700,In_1051);
nor U16 (N_16,In_154,In_666);
nor U17 (N_17,In_1460,In_1414);
xnor U18 (N_18,In_693,In_936);
nor U19 (N_19,In_1240,In_676);
and U20 (N_20,In_399,In_2277);
or U21 (N_21,In_1829,In_259);
nand U22 (N_22,In_2192,In_2310);
nand U23 (N_23,In_2327,In_1620);
or U24 (N_24,In_1305,In_36);
or U25 (N_25,In_1807,In_1693);
and U26 (N_26,In_969,In_721);
nand U27 (N_27,In_858,In_956);
and U28 (N_28,In_1530,In_1034);
and U29 (N_29,In_2118,In_1548);
nand U30 (N_30,In_716,In_2467);
nor U31 (N_31,In_719,In_639);
and U32 (N_32,In_1148,In_106);
nor U33 (N_33,In_602,In_1408);
nand U34 (N_34,In_350,In_994);
nand U35 (N_35,In_127,In_2158);
nand U36 (N_36,In_2132,In_678);
or U37 (N_37,In_1208,In_637);
nor U38 (N_38,In_2110,In_576);
xnor U39 (N_39,In_995,In_2037);
or U40 (N_40,In_2226,In_1689);
nor U41 (N_41,In_2446,In_873);
nand U42 (N_42,In_1737,In_1216);
xor U43 (N_43,In_1366,In_765);
nand U44 (N_44,In_770,In_2249);
and U45 (N_45,In_1618,In_18);
nand U46 (N_46,In_1009,In_1000);
and U47 (N_47,In_293,In_1576);
nand U48 (N_48,In_798,In_1298);
nand U49 (N_49,In_124,In_1919);
xor U50 (N_50,In_308,In_1699);
and U51 (N_51,In_57,In_433);
and U52 (N_52,In_482,In_1037);
or U53 (N_53,In_2430,In_2116);
nand U54 (N_54,In_1959,In_1776);
nand U55 (N_55,In_1407,In_1008);
and U56 (N_56,In_1002,In_253);
nor U57 (N_57,In_1753,In_1083);
nor U58 (N_58,In_589,In_1426);
and U59 (N_59,In_2129,In_249);
or U60 (N_60,In_432,In_2356);
or U61 (N_61,In_2415,In_1715);
and U62 (N_62,In_2330,In_1277);
or U63 (N_63,In_1154,In_1482);
xnor U64 (N_64,In_986,In_420);
or U65 (N_65,In_2094,In_2397);
nor U66 (N_66,In_1123,In_606);
and U67 (N_67,In_1757,In_583);
nand U68 (N_68,In_1995,In_413);
and U69 (N_69,In_486,In_918);
or U70 (N_70,In_774,In_2391);
nand U71 (N_71,In_704,In_2191);
or U72 (N_72,In_1915,In_2027);
or U73 (N_73,In_44,In_954);
or U74 (N_74,In_1067,In_1924);
xor U75 (N_75,In_1734,In_1522);
xnor U76 (N_76,In_1076,In_1219);
nand U77 (N_77,In_1336,In_2239);
nor U78 (N_78,In_1974,In_1690);
and U79 (N_79,In_2342,In_2151);
or U80 (N_80,In_56,In_1955);
and U81 (N_81,In_1505,In_310);
xor U82 (N_82,In_2026,In_1434);
or U83 (N_83,In_980,In_2312);
and U84 (N_84,In_1373,In_1702);
nand U85 (N_85,In_642,In_1279);
nor U86 (N_86,In_1678,In_1072);
nor U87 (N_87,In_1615,In_1095);
or U88 (N_88,In_11,In_832);
or U89 (N_89,In_1790,In_117);
nor U90 (N_90,In_2228,In_1852);
and U91 (N_91,In_2296,In_377);
and U92 (N_92,In_1934,In_845);
xor U93 (N_93,In_2081,In_1064);
nor U94 (N_94,In_248,In_552);
nand U95 (N_95,In_1580,In_315);
and U96 (N_96,In_547,In_1958);
nor U97 (N_97,In_1747,In_138);
nand U98 (N_98,In_1015,In_343);
and U99 (N_99,In_788,In_2180);
nor U100 (N_100,In_1348,In_1192);
and U101 (N_101,In_1012,In_992);
or U102 (N_102,In_1106,In_1759);
nand U103 (N_103,In_1888,In_940);
and U104 (N_104,In_2302,In_368);
nand U105 (N_105,In_1722,In_1116);
xor U106 (N_106,In_444,In_254);
nand U107 (N_107,In_62,In_644);
nor U108 (N_108,In_1473,In_1338);
xnor U109 (N_109,In_2058,In_1384);
nor U110 (N_110,In_1268,In_1446);
or U111 (N_111,In_963,In_2346);
or U112 (N_112,In_632,In_1783);
and U113 (N_113,In_1409,In_2044);
and U114 (N_114,In_387,In_495);
or U115 (N_115,In_1329,In_2285);
or U116 (N_116,In_1654,In_730);
xnor U117 (N_117,In_278,In_148);
nor U118 (N_118,In_722,In_1978);
and U119 (N_119,In_1812,In_2365);
xnor U120 (N_120,In_1883,In_706);
and U121 (N_121,In_1103,In_1029);
and U122 (N_122,In_191,In_1272);
and U123 (N_123,In_2208,In_917);
nor U124 (N_124,In_1508,In_1956);
nor U125 (N_125,In_1014,In_939);
nand U126 (N_126,In_1511,In_2381);
nor U127 (N_127,In_814,In_2144);
nor U128 (N_128,In_2413,In_2259);
and U129 (N_129,In_1245,In_1592);
or U130 (N_130,In_1808,In_1249);
nor U131 (N_131,In_574,In_338);
and U132 (N_132,In_1781,In_727);
or U133 (N_133,In_623,In_2219);
or U134 (N_134,In_1805,In_1677);
xor U135 (N_135,In_285,In_900);
nand U136 (N_136,In_1447,In_800);
nor U137 (N_137,In_2344,In_115);
or U138 (N_138,In_2085,In_1971);
or U139 (N_139,In_1417,In_1480);
and U140 (N_140,In_1102,In_67);
nor U141 (N_141,In_1612,In_94);
and U142 (N_142,In_861,In_1112);
or U143 (N_143,In_2177,In_593);
and U144 (N_144,In_1452,In_192);
nand U145 (N_145,In_1821,In_833);
nand U146 (N_146,In_2078,In_2126);
or U147 (N_147,In_1844,In_2362);
and U148 (N_148,In_1491,In_1894);
or U149 (N_149,In_610,In_111);
or U150 (N_150,In_846,In_1193);
and U151 (N_151,In_1146,In_745);
nor U152 (N_152,In_648,In_1179);
or U153 (N_153,In_512,In_829);
and U154 (N_154,In_649,In_1742);
nand U155 (N_155,In_1319,In_65);
xor U156 (N_156,In_523,In_738);
nor U157 (N_157,In_640,In_1731);
nand U158 (N_158,In_749,In_1098);
nor U159 (N_159,In_2231,In_2486);
nor U160 (N_160,In_81,In_764);
xor U161 (N_161,In_408,In_2420);
xor U162 (N_162,In_634,In_1975);
nand U163 (N_163,In_1496,In_233);
nand U164 (N_164,In_342,In_234);
and U165 (N_165,In_965,In_540);
and U166 (N_166,In_1949,In_1282);
and U167 (N_167,In_4,In_2087);
and U168 (N_168,In_712,In_1785);
xnor U169 (N_169,In_1954,In_2477);
nand U170 (N_170,In_1428,In_805);
nor U171 (N_171,In_2246,In_2015);
or U172 (N_172,In_454,In_2222);
xor U173 (N_173,In_431,In_2393);
xor U174 (N_174,In_511,In_654);
and U175 (N_175,In_2384,In_1914);
and U176 (N_176,In_51,In_1190);
nand U177 (N_177,In_2097,In_1773);
nand U178 (N_178,In_2074,In_333);
or U179 (N_179,In_529,In_867);
and U180 (N_180,In_2120,In_2066);
xnor U181 (N_181,In_1784,In_1077);
xnor U182 (N_182,In_1787,In_16);
and U183 (N_183,In_1565,In_79);
xnor U184 (N_184,In_675,In_1679);
or U185 (N_185,In_1387,In_2388);
or U186 (N_186,In_1831,In_1944);
nand U187 (N_187,In_1564,In_513);
or U188 (N_188,In_945,In_313);
and U189 (N_189,In_1743,In_2375);
xor U190 (N_190,In_840,In_549);
or U191 (N_191,In_1751,In_1262);
xnor U192 (N_192,In_919,In_2326);
nor U193 (N_193,In_502,In_503);
and U194 (N_194,In_1292,In_2103);
or U195 (N_195,In_159,In_2334);
and U196 (N_196,In_2202,In_1232);
nand U197 (N_197,In_2360,In_1218);
or U198 (N_198,In_113,In_2261);
and U199 (N_199,In_1343,In_1642);
nand U200 (N_200,In_95,In_1019);
nand U201 (N_201,In_443,In_2347);
nand U202 (N_202,In_2034,In_265);
xor U203 (N_203,In_2279,In_448);
nand U204 (N_204,In_35,In_1799);
and U205 (N_205,In_163,In_277);
xor U206 (N_206,In_59,In_1855);
and U207 (N_207,In_756,In_1539);
nor U208 (N_208,In_1090,In_2445);
nor U209 (N_209,In_354,In_695);
nor U210 (N_210,In_471,In_2145);
xnor U211 (N_211,In_799,In_2499);
xnor U212 (N_212,In_1750,In_1011);
nor U213 (N_213,In_1641,In_2492);
xor U214 (N_214,In_859,In_686);
nor U215 (N_215,In_677,In_1161);
xnor U216 (N_216,In_2468,In_517);
and U217 (N_217,In_819,In_1741);
nor U218 (N_218,In_1286,In_1477);
and U219 (N_219,In_1285,In_605);
xnor U220 (N_220,In_620,In_83);
and U221 (N_221,In_1345,In_20);
nor U222 (N_222,In_2050,In_1151);
nor U223 (N_223,In_1624,In_2456);
and U224 (N_224,In_720,In_532);
nand U225 (N_225,In_1220,In_755);
xor U226 (N_226,In_2159,In_1598);
nand U227 (N_227,In_524,In_1501);
xnor U228 (N_228,In_1206,In_2021);
nor U229 (N_229,In_1858,In_2271);
nand U230 (N_230,In_1411,In_2088);
and U231 (N_231,In_1467,In_1695);
or U232 (N_232,In_1092,In_2176);
xor U233 (N_233,In_2369,In_638);
and U234 (N_234,In_2282,In_1801);
nor U235 (N_235,In_1705,In_331);
and U236 (N_236,In_1712,In_1614);
or U237 (N_237,In_926,In_2476);
nand U238 (N_238,In_668,In_1004);
xor U239 (N_239,In_1435,In_417);
xnor U240 (N_240,In_1466,In_1109);
nor U241 (N_241,In_88,In_1068);
or U242 (N_242,In_1517,In_2153);
xnor U243 (N_243,In_1257,In_207);
or U244 (N_244,In_1039,In_1010);
or U245 (N_245,In_824,In_2341);
nor U246 (N_246,In_1122,In_1114);
and U247 (N_247,In_209,In_674);
nand U248 (N_248,In_1431,In_694);
nor U249 (N_249,In_1557,In_683);
nand U250 (N_250,In_1374,In_1323);
xnor U251 (N_251,In_1880,In_932);
and U252 (N_252,In_2287,In_337);
xnor U253 (N_253,In_1965,In_2214);
xor U254 (N_254,In_2041,In_2216);
nor U255 (N_255,In_2458,In_978);
and U256 (N_256,In_551,In_2395);
nor U257 (N_257,In_1720,In_1896);
and U258 (N_258,In_1320,In_2028);
nor U259 (N_259,In_1385,In_2442);
or U260 (N_260,In_1890,In_2303);
nand U261 (N_261,In_1342,In_758);
or U262 (N_262,In_2367,In_72);
and U263 (N_263,In_1033,In_617);
and U264 (N_264,In_380,In_1516);
xnor U265 (N_265,In_815,In_223);
nand U266 (N_266,In_2183,In_1041);
xor U267 (N_267,In_1487,In_311);
nor U268 (N_268,In_14,In_1779);
and U269 (N_269,In_484,In_2127);
xor U270 (N_270,In_863,In_741);
xor U271 (N_271,In_1465,In_550);
and U272 (N_272,In_1261,In_587);
or U273 (N_273,In_1500,In_460);
nor U274 (N_274,In_1656,In_142);
nand U275 (N_275,In_518,In_2412);
xnor U276 (N_276,In_1623,In_2432);
nand U277 (N_277,In_1160,In_2464);
nand U278 (N_278,In_1449,In_2429);
nand U279 (N_279,In_625,In_1199);
or U280 (N_280,In_1271,In_1777);
or U281 (N_281,In_401,In_615);
xor U282 (N_282,In_1952,In_276);
and U283 (N_283,In_1827,In_915);
xnor U284 (N_284,In_904,In_1900);
and U285 (N_285,In_1723,In_2055);
xnor U286 (N_286,In_787,In_1352);
nor U287 (N_287,In_288,In_1479);
xnor U288 (N_288,In_1363,In_944);
or U289 (N_289,In_870,In_2290);
nor U290 (N_290,In_1652,In_2165);
nand U291 (N_291,In_627,In_769);
nand U292 (N_292,In_174,In_1128);
nor U293 (N_293,In_466,In_1802);
nor U294 (N_294,In_1075,In_469);
or U295 (N_295,In_957,In_1927);
xor U296 (N_296,In_137,In_437);
and U297 (N_297,In_2233,In_1484);
and U298 (N_298,In_2431,In_1904);
xor U299 (N_299,In_1846,In_323);
and U300 (N_300,In_435,In_129);
nand U301 (N_301,In_1241,In_1817);
xnor U302 (N_302,In_221,In_101);
xnor U303 (N_303,In_1707,In_1430);
nand U304 (N_304,In_2286,In_145);
and U305 (N_305,In_2318,In_427);
and U306 (N_306,In_171,In_1059);
nor U307 (N_307,In_2406,In_705);
nor U308 (N_308,In_2010,In_2134);
xor U309 (N_309,In_2163,In_737);
nor U310 (N_310,In_412,In_2421);
nand U311 (N_311,In_1023,In_1244);
nor U312 (N_312,In_852,In_450);
or U313 (N_313,In_2090,In_1383);
and U314 (N_314,In_1943,In_2247);
and U315 (N_315,In_1767,In_1658);
nor U316 (N_316,In_2004,In_1645);
or U317 (N_317,In_2073,In_1322);
nand U318 (N_318,In_2150,In_419);
nand U319 (N_319,In_2109,In_2280);
nand U320 (N_320,In_384,In_242);
or U321 (N_321,In_421,In_1818);
xnor U322 (N_322,In_813,In_1729);
and U323 (N_323,In_2045,In_383);
nor U324 (N_324,In_2426,In_2253);
and U325 (N_325,In_700,In_2308);
or U326 (N_326,In_1830,In_1930);
and U327 (N_327,In_1605,In_530);
and U328 (N_328,In_984,In_2465);
xnor U329 (N_329,In_1183,In_2368);
nor U330 (N_330,In_892,In_1486);
or U331 (N_331,In_268,In_1925);
nand U332 (N_332,In_210,In_560);
nand U333 (N_333,In_988,In_2380);
nor U334 (N_334,In_1736,In_2416);
nand U335 (N_335,In_2077,In_960);
xnor U336 (N_336,In_1696,In_1203);
or U337 (N_337,In_2352,In_881);
nand U338 (N_338,In_921,In_1101);
xor U339 (N_339,In_2471,In_275);
nor U340 (N_340,In_2053,In_2457);
or U341 (N_341,In_1356,In_330);
or U342 (N_342,In_568,In_736);
nand U343 (N_343,In_842,In_5);
nand U344 (N_344,In_89,In_1892);
nor U345 (N_345,In_1003,In_2289);
and U346 (N_346,In_1823,In_2351);
nor U347 (N_347,In_753,In_2440);
nand U348 (N_348,In_327,In_1406);
xnor U349 (N_349,In_1278,In_848);
nand U350 (N_350,In_894,In_2104);
nor U351 (N_351,In_60,In_261);
and U352 (N_352,In_1124,In_836);
or U353 (N_353,In_2425,In_319);
nand U354 (N_354,In_239,In_785);
xor U355 (N_355,In_1171,In_2376);
nand U356 (N_356,In_1226,In_537);
and U357 (N_357,In_1439,In_1440);
and U358 (N_358,In_2455,In_1795);
xor U359 (N_359,In_152,In_2059);
xor U360 (N_360,In_526,In_373);
or U361 (N_361,In_1224,In_476);
nor U362 (N_362,In_1659,In_1086);
and U363 (N_363,In_1512,In_1158);
nand U364 (N_364,In_656,In_1275);
nand U365 (N_365,In_743,In_717);
xnor U366 (N_366,In_1584,In_1375);
xnor U367 (N_367,In_463,In_2130);
or U368 (N_368,In_2181,In_1231);
or U369 (N_369,In_1339,In_1593);
nand U370 (N_370,In_2122,In_1026);
and U371 (N_371,In_821,In_49);
or U372 (N_372,In_1770,In_780);
or U373 (N_373,In_2011,In_382);
or U374 (N_374,In_2459,In_1221);
or U375 (N_375,In_1875,In_2101);
nand U376 (N_376,In_750,In_2254);
nand U377 (N_377,In_993,In_82);
nand U378 (N_378,In_2046,In_2453);
nor U379 (N_379,In_803,In_2491);
nor U380 (N_380,In_226,In_1215);
nand U381 (N_381,In_1071,In_2343);
and U382 (N_382,In_2402,In_595);
or U383 (N_383,In_2349,In_312);
nand U384 (N_384,In_979,In_173);
nand U385 (N_385,In_1429,In_2294);
nand U386 (N_386,In_914,In_1503);
nand U387 (N_387,In_1942,In_1537);
and U388 (N_388,In_747,In_1263);
nand U389 (N_389,In_2371,In_1188);
or U390 (N_390,In_2305,In_1456);
nor U391 (N_391,In_205,In_1881);
nor U392 (N_392,In_1481,In_2284);
nor U393 (N_393,In_621,In_2418);
xor U394 (N_394,In_559,In_733);
and U395 (N_395,In_2333,In_1066);
or U396 (N_396,In_657,In_1873);
and U397 (N_397,In_2098,In_726);
and U398 (N_398,In_2329,In_2481);
or U399 (N_399,In_1433,In_1813);
and U400 (N_400,In_2175,In_1816);
xnor U401 (N_401,In_818,In_1842);
nor U402 (N_402,In_1893,In_394);
xor U403 (N_403,In_628,In_179);
xor U404 (N_404,In_473,In_2039);
nor U405 (N_405,In_2063,In_1572);
and U406 (N_406,In_1299,In_884);
and U407 (N_407,In_497,In_1520);
nor U408 (N_408,In_297,In_1786);
xnor U409 (N_409,In_2485,In_161);
xnor U410 (N_410,In_378,In_2032);
nand U411 (N_411,In_515,In_238);
and U412 (N_412,In_2203,In_2339);
or U413 (N_413,In_168,In_1254);
nor U414 (N_414,In_1669,In_1317);
and U415 (N_415,In_2324,In_599);
nand U416 (N_416,In_1990,In_70);
or U417 (N_417,In_977,In_663);
nor U418 (N_418,In_1464,In_1718);
nor U419 (N_419,In_42,In_876);
nor U420 (N_420,In_1591,In_17);
or U421 (N_421,In_1362,In_1588);
or U422 (N_422,In_2187,In_1388);
nor U423 (N_423,In_1402,In_1399);
xnor U424 (N_424,In_797,In_1248);
and U425 (N_425,In_2307,In_2366);
xor U426 (N_426,In_2115,In_352);
and U427 (N_427,In_1028,In_1681);
xnor U428 (N_428,In_533,In_566);
nor U429 (N_429,In_1526,In_355);
or U430 (N_430,In_2317,In_902);
xnor U431 (N_431,In_1964,In_1040);
nor U432 (N_432,In_197,In_1176);
nand U433 (N_433,In_329,In_1867);
xnor U434 (N_434,In_1814,In_2178);
xor U435 (N_435,In_1252,In_506);
nor U436 (N_436,In_215,In_2060);
nand U437 (N_437,In_1771,In_735);
nor U438 (N_438,In_1657,In_77);
and U439 (N_439,In_664,In_1330);
and U440 (N_440,In_1191,In_230);
and U441 (N_441,In_1749,In_1653);
nor U442 (N_442,In_91,In_316);
nand U443 (N_443,In_2267,In_1613);
and U444 (N_444,In_1543,In_869);
xnor U445 (N_445,In_1532,In_1967);
and U446 (N_446,In_32,In_1913);
nand U447 (N_447,In_366,In_1984);
or U448 (N_448,In_2245,In_591);
xnor U449 (N_449,In_1885,In_1989);
nand U450 (N_450,In_651,In_2436);
nor U451 (N_451,In_2298,In_1586);
or U452 (N_452,In_584,In_231);
nor U453 (N_453,In_725,In_150);
and U454 (N_454,In_157,In_1212);
and U455 (N_455,In_2099,In_472);
or U456 (N_456,In_1251,In_440);
or U457 (N_457,In_2469,In_607);
nand U458 (N_458,In_302,In_1201);
or U459 (N_459,In_570,In_775);
nand U460 (N_460,In_1765,In_2378);
xnor U461 (N_461,In_1643,In_2198);
nor U462 (N_462,In_1302,In_2174);
xnor U463 (N_463,In_913,In_768);
xor U464 (N_464,In_164,In_284);
xor U465 (N_465,In_1761,In_1910);
and U466 (N_466,In_303,In_1562);
and U467 (N_467,In_1514,In_1169);
and U468 (N_468,In_2067,In_214);
xor U469 (N_469,In_1863,In_1044);
nor U470 (N_470,In_983,In_1583);
xnor U471 (N_471,In_348,In_562);
or U472 (N_472,In_1550,In_425);
and U473 (N_473,In_2209,In_521);
xnor U474 (N_474,In_685,In_1992);
xor U475 (N_475,In_1048,In_2064);
and U476 (N_476,In_219,In_897);
nand U477 (N_477,In_2408,In_100);
nand U478 (N_478,In_761,In_2407);
nand U479 (N_479,In_1754,In_860);
or U480 (N_480,In_1928,In_1933);
nand U481 (N_481,In_23,In_353);
nor U482 (N_482,In_1337,In_184);
xor U483 (N_483,In_554,In_1675);
nand U484 (N_484,In_2114,In_1360);
nor U485 (N_485,In_825,In_976);
and U486 (N_486,In_1144,In_455);
and U487 (N_487,In_135,In_1309);
nor U488 (N_488,In_478,In_692);
or U489 (N_489,In_2119,In_1833);
xnor U490 (N_490,In_2042,In_1209);
or U491 (N_491,In_1136,In_1256);
and U492 (N_492,In_1444,In_786);
or U493 (N_493,In_2139,In_227);
or U494 (N_494,In_388,In_1382);
or U495 (N_495,In_1401,In_1554);
xor U496 (N_496,In_1493,In_905);
nor U497 (N_497,In_1567,In_2162);
nor U498 (N_498,In_1458,In_2225);
nand U499 (N_499,In_2197,In_376);
or U500 (N_500,In_2359,In_2229);
xnor U501 (N_501,In_359,In_1214);
nor U502 (N_502,In_1606,In_1443);
or U503 (N_503,In_2196,In_2314);
xor U504 (N_504,In_2156,In_2323);
nor U505 (N_505,In_696,In_565);
xor U506 (N_506,In_1521,In_1912);
or U507 (N_507,In_305,In_477);
xor U508 (N_508,In_2185,In_853);
xor U509 (N_509,In_1926,In_781);
and U510 (N_510,In_1175,In_114);
nand U511 (N_511,In_175,In_1621);
nor U512 (N_512,In_2264,In_1324);
or U513 (N_513,In_1422,In_2061);
nor U514 (N_514,In_1436,In_563);
xnor U515 (N_515,In_760,In_2437);
xor U516 (N_516,In_1764,In_2211);
nand U517 (N_517,In_1,In_1834);
nand U518 (N_518,In_1899,In_224);
nor U519 (N_519,In_2451,In_2172);
and U520 (N_520,In_908,In_1869);
nor U521 (N_521,In_1983,In_1365);
and U522 (N_522,In_2112,In_1709);
nand U523 (N_523,In_1703,In_740);
xor U524 (N_524,In_1735,In_1545);
xor U525 (N_525,In_2300,In_1727);
and U526 (N_526,In_30,In_1579);
nor U527 (N_527,In_1381,In_496);
and U528 (N_528,In_494,In_1310);
nor U529 (N_529,In_1970,In_652);
and U530 (N_530,In_2005,In_631);
or U531 (N_531,In_713,In_1782);
or U532 (N_532,In_2404,In_1358);
nand U533 (N_533,In_392,In_1105);
nand U534 (N_534,In_2137,In_1811);
or U535 (N_535,In_2155,In_300);
xnor U536 (N_536,In_837,In_162);
and U537 (N_537,In_489,In_199);
or U538 (N_538,In_1993,In_1636);
or U539 (N_539,In_779,In_1631);
nand U540 (N_540,In_1534,In_2292);
nor U541 (N_541,In_186,In_1202);
nor U542 (N_542,In_2257,In_103);
and U543 (N_543,In_1376,In_2309);
and U544 (N_544,In_409,In_1181);
or U545 (N_545,In_1140,In_682);
or U546 (N_546,In_1716,In_2013);
nor U547 (N_547,In_1239,In_282);
or U548 (N_548,In_865,In_601);
and U549 (N_549,In_415,In_949);
and U550 (N_550,In_734,In_1062);
nand U551 (N_551,In_834,In_1270);
nor U552 (N_552,In_754,In_2017);
nor U553 (N_553,In_1344,In_1167);
nand U554 (N_554,In_158,In_260);
and U555 (N_555,In_292,In_1663);
nand U556 (N_556,In_126,In_1932);
or U557 (N_557,In_2111,In_2398);
or U558 (N_558,In_1629,In_912);
or U559 (N_559,In_927,In_2070);
nor U560 (N_560,In_133,In_1025);
nand U561 (N_561,In_2385,In_189);
nor U562 (N_562,In_609,In_1483);
and U563 (N_563,In_1774,In_1237);
and U564 (N_564,In_262,In_180);
xnor U565 (N_565,In_404,In_2474);
nand U566 (N_566,In_470,In_220);
nor U567 (N_567,In_1921,In_2452);
nor U568 (N_568,In_1052,In_929);
nor U569 (N_569,In_1826,In_479);
or U570 (N_570,In_2071,In_1845);
and U571 (N_571,In_2207,In_2396);
nand U572 (N_572,In_1851,In_2128);
nand U573 (N_573,In_46,In_531);
and U574 (N_574,In_1180,In_322);
and U575 (N_575,In_1648,In_2301);
nand U576 (N_576,In_449,In_1198);
nand U577 (N_577,In_2399,In_1638);
nor U578 (N_578,In_828,In_48);
nor U579 (N_579,In_1457,In_294);
and U580 (N_580,In_1523,In_2361);
xor U581 (N_581,In_603,In_2401);
xor U582 (N_582,In_2454,In_1939);
nand U583 (N_583,In_2234,In_92);
and U584 (N_584,In_538,In_2251);
xor U585 (N_585,In_1472,In_177);
xnor U586 (N_586,In_616,In_1471);
xor U587 (N_587,In_2164,In_1536);
nor U588 (N_588,In_938,In_742);
or U589 (N_589,In_1108,In_235);
nand U590 (N_590,In_794,In_714);
and U591 (N_591,In_951,In_370);
and U592 (N_592,In_2188,In_1544);
nand U593 (N_593,In_1755,In_429);
nand U594 (N_594,In_1178,In_975);
and U595 (N_595,In_1985,In_78);
xor U596 (N_596,In_1130,In_21);
xor U597 (N_597,In_190,In_255);
nor U598 (N_598,In_931,In_608);
and U599 (N_599,In_0,In_2173);
and U600 (N_600,In_363,In_2353);
xor U601 (N_601,In_964,In_1389);
nor U602 (N_602,In_2470,In_2093);
xor U603 (N_603,In_1698,In_1552);
nor U604 (N_604,In_105,In_86);
and U605 (N_605,In_349,In_1016);
nor U606 (N_606,In_1726,In_240);
nand U607 (N_607,In_1288,In_1459);
nor U608 (N_608,In_2478,In_1570);
nand U609 (N_609,In_1877,In_2379);
nand U610 (N_610,In_320,In_1832);
and U611 (N_611,In_1671,In_1980);
nor U612 (N_612,In_2210,In_1916);
nor U613 (N_613,In_365,In_2147);
or U614 (N_614,In_519,In_1223);
nor U615 (N_615,In_462,In_1468);
nor U616 (N_616,In_2328,In_522);
and U617 (N_617,In_534,In_345);
or U618 (N_618,In_1021,In_1253);
or U619 (N_619,In_558,In_630);
xor U620 (N_620,In_1451,In_1207);
or U621 (N_621,In_1788,In_123);
nor U622 (N_622,In_116,In_1312);
and U623 (N_623,In_1478,In_2258);
and U624 (N_624,In_1131,In_1730);
and U625 (N_625,In_271,In_1184);
nand U626 (N_626,In_1866,In_1555);
xor U627 (N_627,In_400,In_1266);
nand U628 (N_628,In_2386,In_514);
and U629 (N_629,In_999,In_281);
and U630 (N_630,In_1088,In_636);
nand U631 (N_631,In_360,In_2062);
nand U632 (N_632,In_1841,In_458);
nand U633 (N_633,In_1152,In_1581);
or U634 (N_634,In_2102,In_1332);
nor U635 (N_635,In_1664,In_2206);
nand U636 (N_636,In_811,In_2200);
nor U637 (N_637,In_2480,In_1822);
xnor U638 (N_638,In_1917,In_2218);
and U639 (N_639,In_1168,In_2113);
xnor U640 (N_640,In_959,In_1334);
nand U641 (N_641,In_2283,In_941);
xnor U642 (N_642,In_1427,In_996);
and U643 (N_643,In_291,In_868);
and U644 (N_644,In_134,In_822);
nand U645 (N_645,In_1574,In_2171);
and U646 (N_646,In_1093,In_325);
nand U647 (N_647,In_2269,In_1864);
nand U648 (N_648,In_9,In_2472);
or U649 (N_649,In_626,In_1903);
and U650 (N_650,In_28,In_2387);
or U651 (N_651,In_237,In_1073);
and U652 (N_652,In_1423,In_2023);
or U653 (N_653,In_1284,In_367);
nor U654 (N_654,In_724,In_650);
nand U655 (N_655,In_2291,In_1596);
and U656 (N_656,In_139,In_1839);
or U657 (N_657,In_2293,In_681);
xor U658 (N_658,In_1878,In_2428);
or U659 (N_659,In_1665,In_1556);
nand U660 (N_660,In_2484,In_2444);
and U661 (N_661,In_410,In_879);
nand U662 (N_662,In_1475,In_689);
and U663 (N_663,In_985,In_1020);
xor U664 (N_664,In_1089,In_1999);
or U665 (N_665,In_2466,In_1617);
nor U666 (N_666,In_1533,In_1603);
nand U667 (N_667,In_2410,In_87);
nand U668 (N_668,In_806,In_2003);
nand U669 (N_669,In_452,In_441);
and U670 (N_670,In_1540,In_1670);
or U671 (N_671,In_418,In_1968);
xnor U672 (N_672,In_545,In_2096);
xor U673 (N_673,In_1791,In_1835);
or U674 (N_674,In_385,In_2179);
and U675 (N_675,In_1361,In_998);
and U676 (N_676,In_864,In_2166);
nor U677 (N_677,In_1630,In_202);
nor U678 (N_678,In_1474,In_459);
or U679 (N_679,In_1289,In_2138);
nand U680 (N_680,In_2095,In_588);
xor U681 (N_681,In_166,In_709);
nand U682 (N_682,In_567,In_1518);
or U683 (N_683,In_2160,In_1963);
nor U684 (N_684,In_2092,In_1229);
and U685 (N_685,In_2498,In_1997);
or U686 (N_686,In_326,In_2443);
xnor U687 (N_687,In_1056,In_1394);
and U688 (N_688,In_1159,In_97);
and U689 (N_689,In_1174,In_6);
nand U690 (N_690,In_1081,In_1941);
nand U691 (N_691,In_109,In_746);
xor U692 (N_692,In_1094,In_796);
and U693 (N_693,In_600,In_375);
or U694 (N_694,In_2135,In_1135);
xnor U695 (N_695,In_1082,In_1300);
nor U696 (N_696,In_793,In_835);
and U697 (N_697,In_1355,In_128);
xor U698 (N_698,In_306,In_66);
xnor U699 (N_699,In_699,In_193);
xor U700 (N_700,In_1515,In_855);
xnor U701 (N_701,In_1682,In_176);
and U702 (N_702,In_490,In_1354);
xnor U703 (N_703,In_1017,In_1469);
nor U704 (N_704,In_2068,In_592);
and U705 (N_705,In_389,In_2048);
nand U706 (N_706,In_1668,In_906);
nand U707 (N_707,In_263,In_1838);
and U708 (N_708,In_1870,In_1155);
or U709 (N_709,In_922,In_317);
or U710 (N_710,In_475,In_53);
nor U711 (N_711,In_911,In_874);
xnor U712 (N_712,In_895,In_2148);
nor U713 (N_713,In_1397,In_1994);
and U714 (N_714,In_1549,In_544);
nand U715 (N_715,In_296,In_1290);
nor U716 (N_716,In_357,In_1230);
nor U717 (N_717,In_1837,In_1121);
xnor U718 (N_718,In_1326,In_165);
and U719 (N_719,In_1147,In_1987);
nand U720 (N_720,In_2392,In_1644);
or U721 (N_721,In_1577,In_195);
or U722 (N_722,In_228,In_2422);
nor U723 (N_723,In_1861,In_1398);
and U724 (N_724,In_928,In_1872);
xnor U725 (N_725,In_1347,In_402);
or U726 (N_726,In_468,In_456);
nand U727 (N_727,In_1820,In_661);
nor U728 (N_728,In_270,In_2167);
and U729 (N_729,In_2370,In_2019);
nor U730 (N_730,In_2275,In_447);
xor U731 (N_731,In_1156,In_54);
xor U732 (N_732,In_1553,In_1711);
nor U733 (N_733,In_1796,In_2332);
nand U734 (N_734,In_1857,In_1929);
xnor U735 (N_735,In_390,In_1738);
nor U736 (N_736,In_31,In_2409);
nor U737 (N_737,In_393,In_888);
xnor U738 (N_738,In_1951,In_1499);
nor U739 (N_739,In_791,In_997);
or U740 (N_740,In_182,In_1905);
xnor U741 (N_741,In_1824,In_1946);
nor U742 (N_742,In_1291,In_1884);
nand U743 (N_743,In_1868,In_1400);
or U744 (N_744,In_374,In_1306);
xnor U745 (N_745,In_334,In_1055);
nor U746 (N_746,In_1045,In_776);
and U747 (N_747,In_1316,In_187);
xor U748 (N_748,In_898,In_2320);
or U749 (N_749,In_1227,In_2363);
xor U750 (N_750,In_1424,In_85);
nor U751 (N_751,In_789,In_411);
nor U752 (N_752,In_1119,In_2319);
or U753 (N_753,In_1217,In_856);
xor U754 (N_754,In_527,In_2036);
or U755 (N_755,In_2414,In_577);
nand U756 (N_756,In_188,In_1335);
or U757 (N_757,In_2051,In_1504);
nor U758 (N_758,In_1461,In_204);
nor U759 (N_759,In_422,In_1745);
and U760 (N_760,In_827,In_1611);
nand U761 (N_761,In_1281,In_658);
and U762 (N_762,In_1107,In_2265);
nor U763 (N_763,In_141,In_546);
nor U764 (N_764,In_1351,In_119);
or U765 (N_765,In_1986,In_525);
and U766 (N_766,In_76,In_1962);
nand U767 (N_767,In_336,In_1038);
xor U768 (N_768,In_1099,In_885);
xnor U769 (N_769,In_762,In_1173);
nand U770 (N_770,In_633,In_492);
and U771 (N_771,In_10,In_2439);
xor U772 (N_772,In_1007,In_1819);
or U773 (N_773,In_1455,In_2383);
and U774 (N_774,In_485,In_968);
xor U775 (N_775,In_1639,In_1717);
or U776 (N_776,In_136,In_206);
nor U777 (N_777,In_1024,In_1196);
nand U778 (N_778,In_147,In_2189);
or U779 (N_779,In_22,In_1981);
nor U780 (N_780,In_2002,In_1247);
or U781 (N_781,In_1937,In_2461);
or U782 (N_782,In_1710,In_1953);
nor U783 (N_783,In_792,In_1810);
nand U784 (N_784,In_1142,In_1666);
or U785 (N_785,In_539,In_1157);
or U786 (N_786,In_272,In_1874);
xor U787 (N_787,In_1922,In_1441);
nand U788 (N_788,In_2136,In_1804);
xor U789 (N_789,In_1728,In_1882);
nor U790 (N_790,In_680,In_19);
nor U791 (N_791,In_820,In_71);
or U792 (N_792,In_594,In_1590);
or U793 (N_793,In_1719,In_771);
nand U794 (N_794,In_847,In_1573);
or U795 (N_795,In_324,In_2108);
nor U796 (N_796,In_2124,In_2056);
or U797 (N_797,In_2295,In_2012);
nor U798 (N_798,In_1887,In_2255);
or U799 (N_799,In_2357,In_1442);
nor U800 (N_800,In_2400,In_1166);
nor U801 (N_801,In_1134,In_1233);
xnor U802 (N_802,In_1672,In_896);
xnor U803 (N_803,In_2086,In_2043);
nor U804 (N_804,In_1463,In_991);
nor U805 (N_805,In_536,In_1437);
nand U806 (N_806,In_208,In_1704);
nor U807 (N_807,In_1138,In_1769);
nor U808 (N_808,In_1961,In_1380);
xor U809 (N_809,In_1485,In_33);
nor U810 (N_810,In_1100,In_1558);
xnor U811 (N_811,In_2217,In_1996);
nor U812 (N_812,In_575,In_1027);
nand U813 (N_813,In_1507,In_93);
nand U814 (N_814,In_972,In_406);
nor U815 (N_815,In_1575,In_1561);
nor U816 (N_816,In_614,In_2125);
nor U817 (N_817,In_2205,In_217);
xnor U818 (N_818,In_807,In_1714);
nand U819 (N_819,In_1488,In_2157);
xnor U820 (N_820,In_598,In_120);
and U821 (N_821,In_314,In_1043);
nor U822 (N_822,In_505,In_710);
or U823 (N_823,In_37,In_1849);
and U824 (N_824,In_1889,In_573);
nor U825 (N_825,In_843,In_1364);
xor U826 (N_826,In_773,In_118);
xnor U827 (N_827,In_1162,In_1448);
nor U828 (N_828,In_1204,In_391);
xnor U829 (N_829,In_2495,In_183);
or U830 (N_830,In_2288,In_950);
or U831 (N_831,In_1379,In_467);
and U832 (N_832,In_1748,In_509);
nand U833 (N_833,In_407,In_1070);
nand U834 (N_834,In_857,In_1848);
and U835 (N_835,In_772,In_201);
or U836 (N_836,In_1906,In_140);
nor U837 (N_837,In_586,In_2014);
or U838 (N_838,In_2049,In_1662);
nor U839 (N_839,In_952,In_943);
and U840 (N_840,In_2154,In_1110);
nand U841 (N_841,In_500,In_1368);
or U842 (N_842,In_358,In_55);
xnor U843 (N_843,In_2201,In_2411);
or U844 (N_844,In_2140,In_1104);
nand U845 (N_845,In_619,In_1308);
and U846 (N_846,In_543,In_1862);
or U847 (N_847,In_2268,In_751);
xnor U848 (N_848,In_2035,In_1065);
and U849 (N_849,In_2262,In_1314);
xor U850 (N_850,In_823,In_1594);
and U851 (N_851,In_569,In_1210);
nor U852 (N_852,In_252,In_1497);
nand U853 (N_853,In_582,In_1137);
and U854 (N_854,In_2297,In_701);
and U855 (N_855,In_886,In_1547);
xnor U856 (N_856,In_1972,In_1315);
and U857 (N_857,In_1265,In_782);
and U858 (N_858,In_830,In_2213);
nor U859 (N_859,In_298,In_1050);
xor U860 (N_860,In_2348,In_1129);
and U861 (N_861,In_2345,In_1634);
nand U862 (N_862,In_2260,In_1260);
and U863 (N_863,In_264,In_1234);
nand U864 (N_864,In_1806,In_1908);
xor U865 (N_865,In_2030,In_809);
or U866 (N_866,In_102,In_1153);
xnor U867 (N_867,In_2270,In_424);
nor U868 (N_868,In_436,In_344);
xor U869 (N_869,In_535,In_1694);
and U870 (N_870,In_1622,In_2244);
nor U871 (N_871,In_446,In_1139);
or U872 (N_872,In_763,In_889);
nand U873 (N_873,In_1600,In_1006);
and U874 (N_874,In_2355,In_2024);
nand U875 (N_875,In_810,In_501);
xnor U876 (N_876,In_1988,In_2054);
nand U877 (N_877,In_2389,In_2186);
xnor U878 (N_878,In_1935,In_2435);
and U879 (N_879,In_2463,In_850);
and U880 (N_880,In_715,In_731);
or U881 (N_881,In_2084,In_2076);
and U882 (N_882,In_1898,In_1280);
or U883 (N_883,In_930,In_26);
or U884 (N_884,In_1325,In_241);
nor U885 (N_885,In_1133,In_2281);
nand U886 (N_886,In_108,In_1421);
or U887 (N_887,In_660,In_2450);
nor U888 (N_888,In_2315,In_52);
nand U889 (N_889,In_1969,In_1931);
or U890 (N_890,In_104,In_1792);
nor U891 (N_891,In_2335,In_966);
nand U892 (N_892,In_2141,In_653);
xor U893 (N_893,In_346,In_1651);
nor U894 (N_894,In_266,In_572);
nand U895 (N_895,In_624,In_491);
and U896 (N_896,In_2082,In_2350);
xnor U897 (N_897,In_372,In_1200);
nor U898 (N_898,In_341,In_178);
or U899 (N_899,In_1087,In_1840);
or U900 (N_900,In_2161,In_1489);
and U901 (N_901,In_1120,In_1413);
xor U902 (N_902,In_1947,In_1966);
xor U903 (N_903,In_1766,In_1390);
nor U904 (N_904,In_1327,In_2117);
nand U905 (N_905,In_1392,In_1836);
or U906 (N_906,In_2131,In_1746);
nand U907 (N_907,In_1982,In_461);
nor U908 (N_908,In_2497,In_1495);
or U909 (N_909,In_1405,In_1684);
xor U910 (N_910,In_34,In_1163);
or U911 (N_911,In_1371,In_1490);
or U912 (N_912,In_507,In_804);
nor U913 (N_913,In_110,In_7);
or U914 (N_914,In_1307,In_15);
and U915 (N_915,In_1793,In_1506);
or U916 (N_916,In_2146,In_672);
nand U917 (N_917,In_1789,In_1420);
and U918 (N_918,In_1074,In_256);
nor U919 (N_919,In_541,In_1991);
and U920 (N_920,In_1803,In_643);
or U921 (N_921,In_1030,In_1843);
nand U922 (N_922,In_1053,In_1891);
and U923 (N_923,In_1304,In_2007);
nor U924 (N_924,In_2221,In_47);
and U925 (N_925,In_590,In_1902);
xor U926 (N_926,In_1650,In_1940);
nand U927 (N_927,In_222,In_2419);
nand U928 (N_928,In_2405,In_2106);
nand U929 (N_929,In_581,In_1559);
nor U930 (N_930,In_185,In_1740);
xnor U931 (N_931,In_1189,In_1242);
nor U932 (N_932,In_1524,In_688);
and U933 (N_933,In_38,In_1186);
or U934 (N_934,In_1775,In_2475);
and U935 (N_935,In_817,In_1412);
xor U936 (N_936,In_1492,In_1607);
xnor U937 (N_937,In_2069,In_2133);
xnor U938 (N_938,In_1205,In_131);
xnor U939 (N_939,In_2215,In_381);
nor U940 (N_940,In_2299,In_901);
or U941 (N_941,In_579,In_795);
xnor U942 (N_942,In_2204,In_618);
or U943 (N_943,In_1047,In_2075);
or U944 (N_944,In_2448,In_556);
xor U945 (N_945,In_887,In_816);
and U946 (N_946,In_1509,In_1920);
or U947 (N_947,In_2252,In_2169);
and U948 (N_948,In_1674,In_1113);
or U949 (N_949,In_597,In_1372);
xnor U950 (N_950,In_784,In_2338);
xnor U951 (N_951,In_2276,In_428);
xnor U952 (N_952,In_481,In_1566);
nor U953 (N_953,In_2487,In_580);
nor U954 (N_954,In_2242,In_647);
or U955 (N_955,In_1378,In_151);
and U956 (N_956,In_971,In_1568);
or U957 (N_957,In_854,In_2273);
nand U958 (N_958,In_1510,In_2337);
nand U959 (N_959,In_982,In_872);
and U960 (N_960,In_2313,In_1115);
nand U961 (N_961,In_283,In_1111);
and U962 (N_962,In_1321,In_61);
and U963 (N_963,In_2194,In_416);
and U964 (N_964,In_1069,In_457);
and U965 (N_965,In_578,In_2009);
nor U966 (N_966,In_172,In_783);
xor U967 (N_967,In_1850,In_236);
and U968 (N_968,In_1697,In_1415);
or U969 (N_969,In_1293,In_1798);
xnor U970 (N_970,In_1117,In_112);
xor U971 (N_971,In_920,In_1462);
nand U972 (N_972,In_1494,In_925);
xnor U973 (N_973,In_1527,In_662);
and U974 (N_974,In_2072,In_39);
and U975 (N_975,In_1528,In_280);
or U976 (N_976,In_1454,In_2168);
nor U977 (N_977,In_493,In_1118);
or U978 (N_978,In_1778,In_2274);
nand U979 (N_979,In_812,In_923);
nand U980 (N_980,In_274,In_2100);
and U981 (N_981,In_1255,In_1246);
nand U982 (N_982,In_1708,In_1901);
xnor U983 (N_983,In_1125,In_1259);
nand U984 (N_984,In_916,In_671);
nand U985 (N_985,In_2190,In_2438);
nor U986 (N_986,In_1313,In_2031);
or U987 (N_987,In_2022,In_430);
nand U988 (N_988,In_2394,In_1706);
nor U989 (N_989,In_1762,In_1541);
nand U990 (N_990,In_130,In_1688);
nor U991 (N_991,In_438,In_1060);
nor U992 (N_992,In_1768,In_1815);
and U993 (N_993,In_1854,In_1236);
nand U994 (N_994,In_670,In_2306);
or U995 (N_995,In_1560,In_122);
nor U996 (N_996,In_132,In_1228);
nand U997 (N_997,In_2372,In_1311);
xnor U998 (N_998,In_1097,In_1936);
and U999 (N_999,In_1973,In_759);
nor U1000 (N_1000,In_2184,In_2083);
or U1001 (N_1001,In_723,In_395);
nand U1002 (N_1002,In_1177,In_1367);
or U1003 (N_1003,In_2025,In_328);
xor U1004 (N_1004,In_2236,In_1350);
and U1005 (N_1005,In_1713,In_989);
nand U1006 (N_1006,In_646,In_748);
or U1007 (N_1007,In_153,In_910);
or U1008 (N_1008,In_1318,In_1979);
nand U1009 (N_1009,In_1425,In_1610);
and U1010 (N_1010,In_1150,In_160);
xor U1011 (N_1011,In_155,In_2489);
nand U1012 (N_1012,In_143,In_2494);
and U1013 (N_1013,In_1187,In_321);
nand U1014 (N_1014,In_1410,In_1998);
and U1015 (N_1015,In_1907,In_1063);
or U1016 (N_1016,In_2220,In_2182);
and U1017 (N_1017,In_414,In_2142);
and U1018 (N_1018,In_1628,In_246);
nor U1019 (N_1019,In_2033,In_877);
xnor U1020 (N_1020,In_2322,In_1626);
or U1021 (N_1021,In_144,In_1724);
nor U1022 (N_1022,In_146,In_2040);
nor U1023 (N_1023,In_622,In_831);
xor U1024 (N_1024,In_181,In_946);
nor U1025 (N_1025,In_1609,In_1084);
nand U1026 (N_1026,In_213,In_1859);
nand U1027 (N_1027,In_1346,In_2462);
and U1028 (N_1028,In_69,In_510);
or U1029 (N_1029,In_1701,In_1127);
nor U1030 (N_1030,In_1078,In_1800);
nor U1031 (N_1031,In_2170,In_200);
xor U1032 (N_1032,In_1772,In_273);
nand U1033 (N_1033,In_1599,In_1911);
xor U1034 (N_1034,In_244,In_2235);
xor U1035 (N_1035,In_555,In_1976);
and U1036 (N_1036,In_2364,In_398);
xnor U1037 (N_1037,In_1195,In_2250);
and U1038 (N_1038,In_2052,In_1847);
nor U1039 (N_1039,In_2240,In_553);
nand U1040 (N_1040,In_2316,In_64);
nor U1041 (N_1041,In_170,In_851);
and U1042 (N_1042,In_1341,In_2029);
xnor U1043 (N_1043,In_396,In_893);
and U1044 (N_1044,In_684,In_891);
and U1045 (N_1045,In_1871,In_766);
nor U1046 (N_1046,In_295,In_1225);
or U1047 (N_1047,In_1733,In_1238);
nor U1048 (N_1048,In_844,In_1054);
or U1049 (N_1049,In_1616,In_1295);
nor U1050 (N_1050,In_1529,In_2382);
or U1051 (N_1051,In_1977,In_970);
or U1052 (N_1052,In_948,In_1418);
and U1053 (N_1053,In_883,In_1164);
or U1054 (N_1054,In_838,In_947);
nor U1055 (N_1055,In_1357,In_1331);
or U1056 (N_1056,In_45,In_962);
nor U1057 (N_1057,In_1276,In_1646);
nor U1058 (N_1058,In_464,In_2121);
or U1059 (N_1059,In_974,In_1660);
xnor U1060 (N_1060,In_702,In_1923);
nand U1061 (N_1061,In_335,In_1595);
nor U1062 (N_1062,In_1692,In_903);
nand U1063 (N_1063,In_955,In_245);
xnor U1064 (N_1064,In_981,In_1036);
nand U1065 (N_1065,In_1760,In_74);
nand U1066 (N_1066,In_1001,In_2460);
or U1067 (N_1067,In_301,In_2449);
nor U1068 (N_1068,In_299,In_909);
nor U1069 (N_1069,In_1264,In_707);
xnor U1070 (N_1070,In_2331,In_1445);
nand U1071 (N_1071,In_371,In_1909);
nand U1072 (N_1072,In_194,In_665);
and U1073 (N_1073,In_1683,In_1601);
or U1074 (N_1074,In_1563,In_1126);
nor U1075 (N_1075,In_1589,In_1531);
nor U1076 (N_1076,In_1582,In_286);
nor U1077 (N_1077,In_445,In_1369);
xnor U1078 (N_1078,In_1853,In_487);
nor U1079 (N_1079,In_2149,In_1604);
nor U1080 (N_1080,In_1393,In_1676);
or U1081 (N_1081,In_1865,In_287);
xor U1082 (N_1082,In_2001,In_1667);
and U1083 (N_1083,In_3,In_2325);
nor U1084 (N_1084,In_937,In_73);
nand U1085 (N_1085,In_604,In_2152);
or U1086 (N_1086,In_516,In_2473);
and U1087 (N_1087,In_967,In_564);
or U1088 (N_1088,In_504,In_2482);
or U1089 (N_1089,In_29,In_2340);
and U1090 (N_1090,In_1303,In_1551);
or U1091 (N_1091,In_1273,In_1432);
nor U1092 (N_1092,In_465,In_340);
and U1093 (N_1093,In_1132,In_2311);
nand U1094 (N_1094,In_612,In_1633);
nand U1095 (N_1095,In_1856,In_1647);
nor U1096 (N_1096,In_1395,In_1403);
nor U1097 (N_1097,In_987,In_718);
or U1098 (N_1098,In_12,In_1035);
and U1099 (N_1099,In_2123,In_2232);
nand U1100 (N_1100,In_426,In_728);
xnor U1101 (N_1101,In_2256,In_1950);
nor U1102 (N_1102,In_2424,In_2272);
nand U1103 (N_1103,In_1057,In_1608);
nand U1104 (N_1104,In_403,In_1957);
nor U1105 (N_1105,In_2091,In_1453);
or U1106 (N_1106,In_880,In_2403);
nand U1107 (N_1107,In_1752,In_1585);
and U1108 (N_1108,In_40,In_247);
xnor U1109 (N_1109,In_790,In_2263);
and U1110 (N_1110,In_752,In_1895);
nor U1111 (N_1111,In_953,In_935);
or U1112 (N_1112,In_1519,In_1438);
nor U1113 (N_1113,In_229,In_571);
nor U1114 (N_1114,In_1661,In_1739);
xor U1115 (N_1115,In_1243,In_480);
xor U1116 (N_1116,In_1269,In_2373);
or U1117 (N_1117,In_1049,In_1274);
and U1118 (N_1118,In_871,In_364);
and U1119 (N_1119,In_2266,In_1525);
nand U1120 (N_1120,In_1149,In_203);
or U1121 (N_1121,In_225,In_361);
nand U1122 (N_1122,In_739,In_862);
or U1123 (N_1123,In_80,In_2065);
xnor U1124 (N_1124,In_1296,In_2199);
nor U1125 (N_1125,In_2496,In_934);
and U1126 (N_1126,In_1013,In_2105);
xnor U1127 (N_1127,In_258,In_2358);
or U1128 (N_1128,In_890,In_1640);
nor U1129 (N_1129,In_121,In_1450);
and U1130 (N_1130,In_801,In_942);
nand U1131 (N_1131,In_2423,In_1340);
nand U1132 (N_1132,In_1756,In_1960);
or U1133 (N_1133,In_405,In_243);
xor U1134 (N_1134,In_1597,In_2079);
nand U1135 (N_1135,In_2490,In_2374);
and U1136 (N_1136,In_2441,In_933);
xnor U1137 (N_1137,In_826,In_757);
xnor U1138 (N_1138,In_1419,In_1938);
and U1139 (N_1139,In_1619,In_1079);
or U1140 (N_1140,In_8,In_1328);
and U1141 (N_1141,In_2488,In_958);
nor U1142 (N_1142,In_907,In_1022);
xnor U1143 (N_1143,In_1294,In_1058);
nor U1144 (N_1144,In_1546,In_483);
nand U1145 (N_1145,In_304,In_508);
or U1146 (N_1146,In_1513,In_1032);
and U1147 (N_1147,In_339,In_961);
or U1148 (N_1148,In_13,In_307);
xor U1149 (N_1149,In_269,In_99);
nand U1150 (N_1150,In_27,In_655);
or U1151 (N_1151,In_211,In_1725);
and U1152 (N_1152,In_2417,In_488);
or U1153 (N_1153,In_1297,In_2427);
nand U1154 (N_1154,In_2,In_673);
or U1155 (N_1155,In_667,In_778);
nand U1156 (N_1156,In_58,In_2223);
xor U1157 (N_1157,In_520,In_1353);
and U1158 (N_1158,In_423,In_1185);
xnor U1159 (N_1159,In_1758,In_1182);
nor U1160 (N_1160,In_2107,In_50);
nor U1161 (N_1161,In_882,In_1170);
nand U1162 (N_1162,In_1879,In_41);
nand U1163 (N_1163,In_1258,In_2493);
or U1164 (N_1164,In_1377,In_90);
or U1165 (N_1165,In_1396,In_1213);
nand U1166 (N_1166,In_2243,In_849);
nor U1167 (N_1167,In_899,In_802);
and U1168 (N_1168,In_2483,In_1096);
xnor U1169 (N_1169,In_2212,In_439);
xnor U1170 (N_1170,In_1732,In_1578);
and U1171 (N_1171,In_267,In_232);
nor U1172 (N_1172,In_2321,In_1287);
nor U1173 (N_1173,In_1172,In_1721);
nand U1174 (N_1174,In_1194,In_2089);
nor U1175 (N_1175,In_2304,In_369);
nand U1176 (N_1176,In_1538,In_645);
or U1177 (N_1177,In_878,In_1794);
or U1178 (N_1178,In_635,In_1046);
nand U1179 (N_1179,In_1632,In_611);
or U1180 (N_1180,In_2434,In_250);
and U1181 (N_1181,In_351,In_196);
and U1182 (N_1182,In_279,In_63);
xnor U1183 (N_1183,In_2006,In_1359);
and U1184 (N_1184,In_1860,In_218);
and U1185 (N_1185,In_2278,In_474);
and U1186 (N_1186,In_2230,In_1301);
nand U1187 (N_1187,In_149,In_1542);
nor U1188 (N_1188,In_669,In_1267);
and U1189 (N_1189,In_68,In_216);
nor U1190 (N_1190,In_96,In_1416);
nor U1191 (N_1191,In_451,In_1886);
and U1192 (N_1192,In_1080,In_585);
nor U1193 (N_1193,In_767,In_25);
nor U1194 (N_1194,In_1635,In_1780);
xnor U1195 (N_1195,In_542,In_1005);
nor U1196 (N_1196,In_1602,In_1250);
xor U1197 (N_1197,In_498,In_2237);
nand U1198 (N_1198,In_698,In_2193);
or U1199 (N_1199,In_2008,In_2227);
and U1200 (N_1200,In_442,In_309);
nor U1201 (N_1201,In_332,In_1687);
xnor U1202 (N_1202,In_2354,In_1680);
and U1203 (N_1203,In_1948,In_659);
nor U1204 (N_1204,In_561,In_2020);
nor U1205 (N_1205,In_732,In_1897);
or U1206 (N_1206,In_2195,In_1470);
or U1207 (N_1207,In_2143,In_1763);
nor U1208 (N_1208,In_1222,In_1211);
and U1209 (N_1209,In_2248,In_156);
nand U1210 (N_1210,In_729,In_1141);
nor U1211 (N_1211,In_98,In_744);
and U1212 (N_1212,In_1685,In_434);
nor U1213 (N_1213,In_251,In_866);
or U1214 (N_1214,In_777,In_1655);
or U1215 (N_1215,In_2038,In_839);
nor U1216 (N_1216,In_691,In_75);
or U1217 (N_1217,In_990,In_1587);
xor U1218 (N_1218,In_2241,In_1061);
or U1219 (N_1219,In_125,In_362);
and U1220 (N_1220,In_973,In_289);
nand U1221 (N_1221,In_557,In_697);
xnor U1222 (N_1222,In_290,In_1091);
xnor U1223 (N_1223,In_2080,In_356);
nor U1224 (N_1224,In_1809,In_1145);
nor U1225 (N_1225,In_379,In_1876);
and U1226 (N_1226,In_2447,In_2336);
and U1227 (N_1227,In_2390,In_1283);
nor U1228 (N_1228,In_1197,In_2000);
and U1229 (N_1229,In_708,In_24);
and U1230 (N_1230,In_1031,In_1797);
nand U1231 (N_1231,In_1502,In_808);
xnor U1232 (N_1232,In_2224,In_2047);
or U1233 (N_1233,In_2433,In_690);
and U1234 (N_1234,In_2016,In_257);
and U1235 (N_1235,In_629,In_2479);
xnor U1236 (N_1236,In_167,In_1744);
nor U1237 (N_1237,In_1673,In_169);
and U1238 (N_1238,In_841,In_687);
nand U1239 (N_1239,In_1085,In_1391);
or U1240 (N_1240,In_1498,In_1042);
xor U1241 (N_1241,In_107,In_1686);
and U1242 (N_1242,In_641,In_84);
and U1243 (N_1243,In_1386,In_875);
or U1244 (N_1244,In_43,In_1828);
or U1245 (N_1245,In_397,In_1370);
nor U1246 (N_1246,In_386,In_679);
and U1247 (N_1247,In_2238,In_1569);
and U1248 (N_1248,In_528,In_1235);
or U1249 (N_1249,In_924,In_2057);
xor U1250 (N_1250,In_1791,In_1331);
or U1251 (N_1251,In_828,In_664);
or U1252 (N_1252,In_770,In_268);
and U1253 (N_1253,In_965,In_410);
or U1254 (N_1254,In_1060,In_1771);
or U1255 (N_1255,In_1492,In_2131);
nor U1256 (N_1256,In_451,In_1137);
or U1257 (N_1257,In_1709,In_2269);
xnor U1258 (N_1258,In_1450,In_164);
nand U1259 (N_1259,In_1285,In_384);
and U1260 (N_1260,In_435,In_2204);
and U1261 (N_1261,In_1444,In_1218);
xnor U1262 (N_1262,In_510,In_405);
xnor U1263 (N_1263,In_645,In_59);
or U1264 (N_1264,In_40,In_346);
nand U1265 (N_1265,In_911,In_98);
nor U1266 (N_1266,In_1495,In_2169);
nor U1267 (N_1267,In_1011,In_2453);
or U1268 (N_1268,In_1426,In_747);
xnor U1269 (N_1269,In_966,In_151);
xnor U1270 (N_1270,In_2156,In_2345);
and U1271 (N_1271,In_57,In_775);
nor U1272 (N_1272,In_1047,In_1736);
nand U1273 (N_1273,In_364,In_1561);
nand U1274 (N_1274,In_352,In_138);
nor U1275 (N_1275,In_2208,In_2268);
xnor U1276 (N_1276,In_1085,In_2070);
nor U1277 (N_1277,In_1750,In_618);
xnor U1278 (N_1278,In_266,In_652);
or U1279 (N_1279,In_2299,In_298);
nand U1280 (N_1280,In_122,In_2116);
and U1281 (N_1281,In_374,In_1506);
xor U1282 (N_1282,In_1631,In_437);
or U1283 (N_1283,In_2166,In_1378);
nand U1284 (N_1284,In_1374,In_1400);
xnor U1285 (N_1285,In_45,In_711);
xnor U1286 (N_1286,In_1120,In_2283);
nor U1287 (N_1287,In_1761,In_1877);
or U1288 (N_1288,In_167,In_1867);
or U1289 (N_1289,In_1976,In_1798);
nor U1290 (N_1290,In_754,In_367);
nand U1291 (N_1291,In_2347,In_1318);
or U1292 (N_1292,In_137,In_464);
xor U1293 (N_1293,In_898,In_342);
or U1294 (N_1294,In_276,In_608);
and U1295 (N_1295,In_1329,In_95);
and U1296 (N_1296,In_1812,In_355);
xor U1297 (N_1297,In_2483,In_2036);
or U1298 (N_1298,In_2195,In_2062);
and U1299 (N_1299,In_685,In_190);
and U1300 (N_1300,In_1609,In_2249);
xnor U1301 (N_1301,In_1208,In_574);
or U1302 (N_1302,In_2007,In_2120);
nand U1303 (N_1303,In_1731,In_1968);
nor U1304 (N_1304,In_2186,In_1542);
and U1305 (N_1305,In_2283,In_1610);
and U1306 (N_1306,In_2013,In_568);
or U1307 (N_1307,In_253,In_1969);
and U1308 (N_1308,In_2219,In_2426);
xor U1309 (N_1309,In_1057,In_1940);
or U1310 (N_1310,In_974,In_699);
nor U1311 (N_1311,In_2252,In_2019);
or U1312 (N_1312,In_931,In_663);
and U1313 (N_1313,In_1253,In_1753);
and U1314 (N_1314,In_1193,In_1030);
or U1315 (N_1315,In_766,In_1453);
or U1316 (N_1316,In_619,In_1652);
and U1317 (N_1317,In_118,In_865);
nand U1318 (N_1318,In_414,In_623);
or U1319 (N_1319,In_2154,In_2062);
nor U1320 (N_1320,In_2213,In_1530);
nand U1321 (N_1321,In_2327,In_26);
or U1322 (N_1322,In_185,In_476);
nand U1323 (N_1323,In_1838,In_273);
nand U1324 (N_1324,In_493,In_1026);
nand U1325 (N_1325,In_1186,In_967);
xnor U1326 (N_1326,In_1333,In_1607);
nand U1327 (N_1327,In_380,In_2316);
nand U1328 (N_1328,In_820,In_1087);
xor U1329 (N_1329,In_1224,In_99);
nor U1330 (N_1330,In_2018,In_135);
or U1331 (N_1331,In_1686,In_1795);
and U1332 (N_1332,In_328,In_300);
nor U1333 (N_1333,In_2052,In_1662);
nand U1334 (N_1334,In_1646,In_1);
xnor U1335 (N_1335,In_805,In_2331);
and U1336 (N_1336,In_777,In_2061);
nor U1337 (N_1337,In_1566,In_506);
or U1338 (N_1338,In_2171,In_2004);
and U1339 (N_1339,In_984,In_1729);
nor U1340 (N_1340,In_1299,In_1037);
xnor U1341 (N_1341,In_517,In_1740);
nor U1342 (N_1342,In_2006,In_295);
or U1343 (N_1343,In_2238,In_2229);
nand U1344 (N_1344,In_1840,In_339);
and U1345 (N_1345,In_2384,In_881);
nand U1346 (N_1346,In_2111,In_342);
nand U1347 (N_1347,In_1756,In_1181);
xor U1348 (N_1348,In_2153,In_1317);
or U1349 (N_1349,In_672,In_1423);
or U1350 (N_1350,In_2062,In_2412);
or U1351 (N_1351,In_1725,In_1246);
xor U1352 (N_1352,In_7,In_1798);
and U1353 (N_1353,In_1372,In_2268);
and U1354 (N_1354,In_1570,In_663);
nor U1355 (N_1355,In_1678,In_2110);
and U1356 (N_1356,In_2075,In_565);
xnor U1357 (N_1357,In_2187,In_1545);
nor U1358 (N_1358,In_1590,In_714);
nand U1359 (N_1359,In_66,In_1411);
nand U1360 (N_1360,In_2445,In_1390);
or U1361 (N_1361,In_774,In_1790);
nor U1362 (N_1362,In_729,In_1363);
or U1363 (N_1363,In_712,In_872);
and U1364 (N_1364,In_2059,In_784);
or U1365 (N_1365,In_13,In_1981);
nor U1366 (N_1366,In_736,In_1985);
xnor U1367 (N_1367,In_761,In_1578);
xnor U1368 (N_1368,In_2426,In_1912);
and U1369 (N_1369,In_1166,In_603);
nor U1370 (N_1370,In_1809,In_1349);
xnor U1371 (N_1371,In_1850,In_643);
nor U1372 (N_1372,In_1342,In_1185);
nor U1373 (N_1373,In_544,In_752);
nor U1374 (N_1374,In_319,In_748);
nor U1375 (N_1375,In_347,In_2194);
xor U1376 (N_1376,In_1467,In_412);
xnor U1377 (N_1377,In_453,In_2366);
or U1378 (N_1378,In_2421,In_2133);
nor U1379 (N_1379,In_2382,In_2112);
and U1380 (N_1380,In_1864,In_2094);
nand U1381 (N_1381,In_225,In_1911);
xnor U1382 (N_1382,In_2199,In_455);
nand U1383 (N_1383,In_822,In_2026);
nor U1384 (N_1384,In_780,In_291);
nor U1385 (N_1385,In_1701,In_2335);
xor U1386 (N_1386,In_1532,In_2196);
and U1387 (N_1387,In_411,In_2198);
nand U1388 (N_1388,In_441,In_1561);
nand U1389 (N_1389,In_306,In_2118);
nand U1390 (N_1390,In_734,In_848);
and U1391 (N_1391,In_613,In_272);
xnor U1392 (N_1392,In_2002,In_1687);
nand U1393 (N_1393,In_1968,In_1280);
and U1394 (N_1394,In_1248,In_640);
or U1395 (N_1395,In_1779,In_2188);
xnor U1396 (N_1396,In_1644,In_810);
nor U1397 (N_1397,In_767,In_2017);
or U1398 (N_1398,In_1693,In_1834);
nand U1399 (N_1399,In_2038,In_2154);
and U1400 (N_1400,In_1393,In_1891);
nand U1401 (N_1401,In_794,In_1452);
and U1402 (N_1402,In_685,In_1239);
or U1403 (N_1403,In_2450,In_2114);
or U1404 (N_1404,In_1150,In_2027);
xor U1405 (N_1405,In_72,In_1450);
nor U1406 (N_1406,In_1814,In_2468);
nor U1407 (N_1407,In_996,In_2278);
xor U1408 (N_1408,In_2264,In_341);
nand U1409 (N_1409,In_1441,In_357);
or U1410 (N_1410,In_191,In_1673);
xnor U1411 (N_1411,In_1400,In_77);
nor U1412 (N_1412,In_1297,In_1031);
nand U1413 (N_1413,In_2466,In_2499);
nand U1414 (N_1414,In_1168,In_2301);
or U1415 (N_1415,In_17,In_1549);
nor U1416 (N_1416,In_788,In_2299);
nor U1417 (N_1417,In_488,In_1631);
nand U1418 (N_1418,In_1382,In_422);
or U1419 (N_1419,In_1712,In_1852);
nor U1420 (N_1420,In_1664,In_353);
or U1421 (N_1421,In_725,In_921);
or U1422 (N_1422,In_1745,In_2387);
or U1423 (N_1423,In_510,In_945);
or U1424 (N_1424,In_189,In_2093);
and U1425 (N_1425,In_1580,In_502);
or U1426 (N_1426,In_1401,In_2407);
xnor U1427 (N_1427,In_268,In_1247);
and U1428 (N_1428,In_1441,In_777);
nor U1429 (N_1429,In_1257,In_1215);
and U1430 (N_1430,In_752,In_1423);
nor U1431 (N_1431,In_2078,In_376);
and U1432 (N_1432,In_1272,In_1336);
and U1433 (N_1433,In_1395,In_1032);
or U1434 (N_1434,In_898,In_704);
nand U1435 (N_1435,In_1007,In_1460);
xor U1436 (N_1436,In_2041,In_2212);
and U1437 (N_1437,In_2079,In_1661);
nand U1438 (N_1438,In_708,In_1713);
xnor U1439 (N_1439,In_410,In_256);
nand U1440 (N_1440,In_1510,In_1917);
nand U1441 (N_1441,In_629,In_2079);
nand U1442 (N_1442,In_2227,In_1415);
nor U1443 (N_1443,In_1673,In_1632);
xnor U1444 (N_1444,In_719,In_2280);
nand U1445 (N_1445,In_1803,In_2286);
or U1446 (N_1446,In_682,In_826);
xnor U1447 (N_1447,In_142,In_1897);
xor U1448 (N_1448,In_2339,In_381);
nor U1449 (N_1449,In_1938,In_1213);
nor U1450 (N_1450,In_733,In_1383);
or U1451 (N_1451,In_1169,In_1690);
nand U1452 (N_1452,In_98,In_7);
and U1453 (N_1453,In_2455,In_1118);
xnor U1454 (N_1454,In_1931,In_4);
and U1455 (N_1455,In_1790,In_548);
xor U1456 (N_1456,In_674,In_1487);
nand U1457 (N_1457,In_1811,In_1736);
nor U1458 (N_1458,In_984,In_2121);
nor U1459 (N_1459,In_294,In_767);
or U1460 (N_1460,In_1127,In_588);
nor U1461 (N_1461,In_1216,In_346);
and U1462 (N_1462,In_748,In_1076);
nor U1463 (N_1463,In_1553,In_2405);
or U1464 (N_1464,In_1283,In_1164);
nor U1465 (N_1465,In_307,In_1639);
or U1466 (N_1466,In_1194,In_947);
and U1467 (N_1467,In_1570,In_1614);
nor U1468 (N_1468,In_1563,In_1164);
xor U1469 (N_1469,In_659,In_1077);
and U1470 (N_1470,In_1764,In_477);
nand U1471 (N_1471,In_1991,In_2399);
nor U1472 (N_1472,In_701,In_488);
nand U1473 (N_1473,In_1353,In_1634);
or U1474 (N_1474,In_1409,In_1082);
and U1475 (N_1475,In_1502,In_2480);
and U1476 (N_1476,In_1139,In_1966);
and U1477 (N_1477,In_82,In_1329);
nand U1478 (N_1478,In_1824,In_1811);
or U1479 (N_1479,In_996,In_152);
nor U1480 (N_1480,In_1073,In_963);
and U1481 (N_1481,In_33,In_2121);
nor U1482 (N_1482,In_267,In_756);
and U1483 (N_1483,In_352,In_188);
nor U1484 (N_1484,In_710,In_677);
or U1485 (N_1485,In_1289,In_2198);
and U1486 (N_1486,In_639,In_207);
nand U1487 (N_1487,In_1948,In_306);
xnor U1488 (N_1488,In_877,In_274);
xor U1489 (N_1489,In_673,In_598);
or U1490 (N_1490,In_1641,In_1262);
xor U1491 (N_1491,In_1811,In_1002);
or U1492 (N_1492,In_2142,In_2054);
nor U1493 (N_1493,In_1645,In_365);
nor U1494 (N_1494,In_1132,In_49);
or U1495 (N_1495,In_1359,In_724);
or U1496 (N_1496,In_335,In_2019);
nor U1497 (N_1497,In_807,In_2359);
nand U1498 (N_1498,In_1291,In_1814);
xnor U1499 (N_1499,In_1205,In_1156);
xnor U1500 (N_1500,In_1085,In_654);
xor U1501 (N_1501,In_2174,In_650);
and U1502 (N_1502,In_1159,In_1354);
nor U1503 (N_1503,In_2063,In_1905);
or U1504 (N_1504,In_2286,In_1410);
nor U1505 (N_1505,In_1700,In_163);
or U1506 (N_1506,In_2132,In_2303);
nand U1507 (N_1507,In_2487,In_1326);
and U1508 (N_1508,In_518,In_333);
or U1509 (N_1509,In_1291,In_2129);
or U1510 (N_1510,In_1484,In_1011);
xor U1511 (N_1511,In_1655,In_844);
xor U1512 (N_1512,In_1586,In_1114);
and U1513 (N_1513,In_2176,In_705);
nand U1514 (N_1514,In_161,In_1501);
nor U1515 (N_1515,In_1759,In_1772);
nor U1516 (N_1516,In_2488,In_570);
xnor U1517 (N_1517,In_2182,In_1173);
nor U1518 (N_1518,In_1030,In_2034);
and U1519 (N_1519,In_605,In_452);
and U1520 (N_1520,In_1088,In_1115);
nand U1521 (N_1521,In_1577,In_1025);
and U1522 (N_1522,In_2307,In_319);
or U1523 (N_1523,In_1140,In_1769);
xnor U1524 (N_1524,In_284,In_315);
nand U1525 (N_1525,In_1554,In_172);
and U1526 (N_1526,In_810,In_2028);
or U1527 (N_1527,In_1472,In_1974);
and U1528 (N_1528,In_1093,In_363);
and U1529 (N_1529,In_1605,In_2059);
xnor U1530 (N_1530,In_84,In_2221);
or U1531 (N_1531,In_1730,In_2148);
nand U1532 (N_1532,In_580,In_2493);
nor U1533 (N_1533,In_1344,In_1555);
or U1534 (N_1534,In_1868,In_769);
xor U1535 (N_1535,In_207,In_2497);
and U1536 (N_1536,In_35,In_76);
xnor U1537 (N_1537,In_1679,In_1638);
xnor U1538 (N_1538,In_1818,In_2474);
nor U1539 (N_1539,In_729,In_2323);
and U1540 (N_1540,In_1970,In_904);
nand U1541 (N_1541,In_453,In_2023);
or U1542 (N_1542,In_1202,In_1918);
nand U1543 (N_1543,In_993,In_1859);
nor U1544 (N_1544,In_1960,In_874);
nand U1545 (N_1545,In_438,In_264);
or U1546 (N_1546,In_1546,In_209);
xnor U1547 (N_1547,In_1813,In_1167);
xor U1548 (N_1548,In_371,In_626);
nand U1549 (N_1549,In_211,In_1899);
nor U1550 (N_1550,In_314,In_1850);
nor U1551 (N_1551,In_810,In_1021);
nor U1552 (N_1552,In_10,In_1281);
and U1553 (N_1553,In_316,In_1706);
nand U1554 (N_1554,In_582,In_96);
nor U1555 (N_1555,In_892,In_1157);
xor U1556 (N_1556,In_2235,In_1792);
xnor U1557 (N_1557,In_193,In_799);
nand U1558 (N_1558,In_1337,In_212);
nand U1559 (N_1559,In_992,In_1533);
or U1560 (N_1560,In_1390,In_414);
nor U1561 (N_1561,In_1121,In_536);
and U1562 (N_1562,In_2187,In_543);
and U1563 (N_1563,In_2207,In_2183);
nor U1564 (N_1564,In_1998,In_1743);
or U1565 (N_1565,In_1669,In_39);
and U1566 (N_1566,In_926,In_587);
or U1567 (N_1567,In_453,In_1837);
and U1568 (N_1568,In_433,In_859);
and U1569 (N_1569,In_2074,In_2368);
nor U1570 (N_1570,In_609,In_1167);
nor U1571 (N_1571,In_991,In_2466);
xor U1572 (N_1572,In_1858,In_179);
nand U1573 (N_1573,In_1028,In_1523);
and U1574 (N_1574,In_1550,In_2183);
and U1575 (N_1575,In_2076,In_1210);
nand U1576 (N_1576,In_25,In_699);
nand U1577 (N_1577,In_636,In_987);
nand U1578 (N_1578,In_1874,In_2297);
nor U1579 (N_1579,In_901,In_2363);
and U1580 (N_1580,In_38,In_146);
xnor U1581 (N_1581,In_1838,In_154);
xor U1582 (N_1582,In_1631,In_1149);
nand U1583 (N_1583,In_1037,In_2416);
xor U1584 (N_1584,In_1911,In_2319);
and U1585 (N_1585,In_1362,In_244);
and U1586 (N_1586,In_2390,In_1486);
xnor U1587 (N_1587,In_1849,In_170);
nor U1588 (N_1588,In_1412,In_56);
xnor U1589 (N_1589,In_265,In_1673);
and U1590 (N_1590,In_1589,In_86);
nand U1591 (N_1591,In_648,In_514);
or U1592 (N_1592,In_156,In_423);
and U1593 (N_1593,In_1091,In_1842);
or U1594 (N_1594,In_1520,In_859);
nand U1595 (N_1595,In_450,In_22);
nor U1596 (N_1596,In_1779,In_355);
xor U1597 (N_1597,In_1478,In_1026);
or U1598 (N_1598,In_1746,In_2048);
nor U1599 (N_1599,In_1599,In_1194);
xor U1600 (N_1600,In_971,In_200);
nor U1601 (N_1601,In_772,In_1373);
nor U1602 (N_1602,In_68,In_2015);
xor U1603 (N_1603,In_1094,In_2200);
nand U1604 (N_1604,In_122,In_789);
and U1605 (N_1605,In_282,In_1682);
nand U1606 (N_1606,In_1485,In_37);
nand U1607 (N_1607,In_2375,In_338);
nor U1608 (N_1608,In_2419,In_2345);
or U1609 (N_1609,In_1650,In_1205);
nand U1610 (N_1610,In_725,In_1811);
nor U1611 (N_1611,In_1170,In_332);
and U1612 (N_1612,In_2412,In_1143);
xor U1613 (N_1613,In_1929,In_1075);
and U1614 (N_1614,In_618,In_920);
and U1615 (N_1615,In_641,In_1136);
and U1616 (N_1616,In_1973,In_2033);
nor U1617 (N_1617,In_657,In_989);
xnor U1618 (N_1618,In_153,In_1882);
nand U1619 (N_1619,In_386,In_1169);
and U1620 (N_1620,In_1131,In_365);
xnor U1621 (N_1621,In_1158,In_1287);
nand U1622 (N_1622,In_1778,In_776);
or U1623 (N_1623,In_1226,In_456);
or U1624 (N_1624,In_102,In_1126);
nor U1625 (N_1625,In_618,In_2473);
xnor U1626 (N_1626,In_784,In_745);
nand U1627 (N_1627,In_1997,In_1968);
nand U1628 (N_1628,In_68,In_2);
nand U1629 (N_1629,In_2419,In_2233);
or U1630 (N_1630,In_1103,In_1022);
or U1631 (N_1631,In_304,In_1555);
or U1632 (N_1632,In_2417,In_199);
nor U1633 (N_1633,In_1314,In_1425);
or U1634 (N_1634,In_1927,In_1537);
and U1635 (N_1635,In_535,In_2434);
or U1636 (N_1636,In_459,In_2061);
and U1637 (N_1637,In_1732,In_1788);
nor U1638 (N_1638,In_65,In_1242);
nor U1639 (N_1639,In_448,In_1583);
or U1640 (N_1640,In_794,In_1891);
xor U1641 (N_1641,In_866,In_845);
nor U1642 (N_1642,In_2096,In_547);
xor U1643 (N_1643,In_270,In_2144);
nor U1644 (N_1644,In_1500,In_1948);
or U1645 (N_1645,In_1580,In_19);
xor U1646 (N_1646,In_2067,In_1449);
or U1647 (N_1647,In_822,In_2393);
and U1648 (N_1648,In_1992,In_666);
xor U1649 (N_1649,In_390,In_73);
or U1650 (N_1650,In_171,In_2306);
nand U1651 (N_1651,In_990,In_137);
xnor U1652 (N_1652,In_697,In_232);
nor U1653 (N_1653,In_1516,In_103);
and U1654 (N_1654,In_775,In_594);
xnor U1655 (N_1655,In_1425,In_2056);
and U1656 (N_1656,In_1754,In_508);
and U1657 (N_1657,In_2088,In_1349);
or U1658 (N_1658,In_2130,In_2350);
xnor U1659 (N_1659,In_1785,In_1889);
xor U1660 (N_1660,In_1227,In_1476);
and U1661 (N_1661,In_8,In_709);
or U1662 (N_1662,In_1517,In_2151);
and U1663 (N_1663,In_1112,In_1092);
or U1664 (N_1664,In_467,In_770);
and U1665 (N_1665,In_1157,In_516);
nand U1666 (N_1666,In_2358,In_2223);
xnor U1667 (N_1667,In_1758,In_1765);
nand U1668 (N_1668,In_1030,In_1242);
nand U1669 (N_1669,In_190,In_379);
nor U1670 (N_1670,In_2098,In_293);
and U1671 (N_1671,In_1485,In_1742);
nand U1672 (N_1672,In_2302,In_1391);
nor U1673 (N_1673,In_73,In_876);
nor U1674 (N_1674,In_1551,In_930);
nor U1675 (N_1675,In_1684,In_1312);
and U1676 (N_1676,In_1106,In_1842);
xor U1677 (N_1677,In_1188,In_2353);
nand U1678 (N_1678,In_652,In_653);
or U1679 (N_1679,In_1487,In_522);
and U1680 (N_1680,In_1051,In_1448);
and U1681 (N_1681,In_1601,In_114);
and U1682 (N_1682,In_1665,In_180);
or U1683 (N_1683,In_1234,In_702);
xor U1684 (N_1684,In_2344,In_2337);
and U1685 (N_1685,In_2206,In_1867);
and U1686 (N_1686,In_723,In_1517);
xor U1687 (N_1687,In_150,In_495);
nand U1688 (N_1688,In_1247,In_1958);
and U1689 (N_1689,In_2483,In_128);
nand U1690 (N_1690,In_1814,In_1303);
or U1691 (N_1691,In_254,In_468);
xnor U1692 (N_1692,In_1853,In_2228);
nand U1693 (N_1693,In_608,In_661);
and U1694 (N_1694,In_2493,In_2469);
or U1695 (N_1695,In_2081,In_2482);
xnor U1696 (N_1696,In_2204,In_978);
nand U1697 (N_1697,In_2179,In_931);
nand U1698 (N_1698,In_1627,In_2495);
xnor U1699 (N_1699,In_10,In_1539);
nor U1700 (N_1700,In_706,In_788);
nor U1701 (N_1701,In_1274,In_2161);
and U1702 (N_1702,In_132,In_295);
and U1703 (N_1703,In_1302,In_207);
xnor U1704 (N_1704,In_1234,In_1122);
nand U1705 (N_1705,In_1884,In_245);
nor U1706 (N_1706,In_1783,In_1931);
nor U1707 (N_1707,In_2470,In_672);
nor U1708 (N_1708,In_887,In_2210);
xnor U1709 (N_1709,In_1468,In_2310);
nand U1710 (N_1710,In_928,In_599);
nand U1711 (N_1711,In_828,In_35);
xor U1712 (N_1712,In_2045,In_13);
xor U1713 (N_1713,In_2277,In_1885);
or U1714 (N_1714,In_474,In_1664);
xor U1715 (N_1715,In_33,In_841);
or U1716 (N_1716,In_1983,In_2361);
nand U1717 (N_1717,In_2333,In_1008);
xor U1718 (N_1718,In_2489,In_1404);
and U1719 (N_1719,In_1971,In_315);
or U1720 (N_1720,In_2029,In_2186);
or U1721 (N_1721,In_1510,In_1914);
and U1722 (N_1722,In_2132,In_1552);
or U1723 (N_1723,In_2322,In_449);
nand U1724 (N_1724,In_1998,In_2422);
or U1725 (N_1725,In_976,In_2000);
and U1726 (N_1726,In_1841,In_2153);
nor U1727 (N_1727,In_233,In_694);
nor U1728 (N_1728,In_1984,In_1747);
and U1729 (N_1729,In_1313,In_2160);
nor U1730 (N_1730,In_817,In_2237);
or U1731 (N_1731,In_2079,In_1720);
nand U1732 (N_1732,In_1164,In_2059);
nor U1733 (N_1733,In_2294,In_965);
or U1734 (N_1734,In_321,In_2053);
nand U1735 (N_1735,In_2240,In_790);
nor U1736 (N_1736,In_509,In_2222);
nor U1737 (N_1737,In_339,In_1913);
and U1738 (N_1738,In_1341,In_2499);
nor U1739 (N_1739,In_1562,In_797);
xor U1740 (N_1740,In_246,In_1880);
nor U1741 (N_1741,In_960,In_1112);
and U1742 (N_1742,In_2377,In_1640);
nand U1743 (N_1743,In_330,In_1224);
nor U1744 (N_1744,In_2189,In_2285);
nor U1745 (N_1745,In_68,In_495);
nor U1746 (N_1746,In_1850,In_882);
and U1747 (N_1747,In_728,In_1210);
or U1748 (N_1748,In_1220,In_2343);
or U1749 (N_1749,In_2421,In_1574);
or U1750 (N_1750,In_934,In_2376);
and U1751 (N_1751,In_908,In_4);
nand U1752 (N_1752,In_1141,In_1496);
and U1753 (N_1753,In_1203,In_666);
or U1754 (N_1754,In_2426,In_2007);
nand U1755 (N_1755,In_2097,In_63);
and U1756 (N_1756,In_616,In_888);
nor U1757 (N_1757,In_2318,In_739);
nand U1758 (N_1758,In_250,In_1445);
and U1759 (N_1759,In_538,In_844);
xor U1760 (N_1760,In_1339,In_1220);
xor U1761 (N_1761,In_931,In_1241);
nand U1762 (N_1762,In_1625,In_315);
and U1763 (N_1763,In_2222,In_2044);
nand U1764 (N_1764,In_361,In_936);
xnor U1765 (N_1765,In_1459,In_1342);
nand U1766 (N_1766,In_341,In_1620);
nor U1767 (N_1767,In_1240,In_471);
nor U1768 (N_1768,In_2359,In_1528);
and U1769 (N_1769,In_49,In_281);
or U1770 (N_1770,In_1700,In_195);
and U1771 (N_1771,In_1414,In_360);
or U1772 (N_1772,In_1487,In_957);
nor U1773 (N_1773,In_264,In_1049);
and U1774 (N_1774,In_2310,In_1635);
nor U1775 (N_1775,In_2325,In_110);
nand U1776 (N_1776,In_2413,In_29);
nor U1777 (N_1777,In_271,In_586);
nor U1778 (N_1778,In_1764,In_2129);
and U1779 (N_1779,In_2095,In_460);
xnor U1780 (N_1780,In_1281,In_220);
xor U1781 (N_1781,In_719,In_2068);
or U1782 (N_1782,In_2088,In_1368);
nand U1783 (N_1783,In_618,In_328);
or U1784 (N_1784,In_2480,In_2070);
nand U1785 (N_1785,In_349,In_1798);
nor U1786 (N_1786,In_637,In_173);
or U1787 (N_1787,In_917,In_1944);
nor U1788 (N_1788,In_1463,In_2486);
xnor U1789 (N_1789,In_52,In_910);
and U1790 (N_1790,In_2156,In_1363);
and U1791 (N_1791,In_1827,In_164);
and U1792 (N_1792,In_545,In_167);
or U1793 (N_1793,In_1626,In_2477);
and U1794 (N_1794,In_2179,In_2487);
nor U1795 (N_1795,In_2374,In_765);
or U1796 (N_1796,In_1803,In_1242);
and U1797 (N_1797,In_2379,In_1759);
nand U1798 (N_1798,In_534,In_832);
nor U1799 (N_1799,In_654,In_1892);
xnor U1800 (N_1800,In_189,In_2195);
nand U1801 (N_1801,In_455,In_1487);
xnor U1802 (N_1802,In_2141,In_1869);
and U1803 (N_1803,In_2410,In_806);
nor U1804 (N_1804,In_1472,In_491);
nand U1805 (N_1805,In_1376,In_896);
nand U1806 (N_1806,In_1122,In_875);
or U1807 (N_1807,In_1384,In_1204);
xor U1808 (N_1808,In_1869,In_1210);
nor U1809 (N_1809,In_1286,In_152);
or U1810 (N_1810,In_1977,In_1014);
nand U1811 (N_1811,In_665,In_1834);
and U1812 (N_1812,In_2119,In_954);
nor U1813 (N_1813,In_1921,In_118);
nor U1814 (N_1814,In_2203,In_2322);
and U1815 (N_1815,In_925,In_311);
or U1816 (N_1816,In_844,In_1270);
or U1817 (N_1817,In_343,In_68);
nor U1818 (N_1818,In_529,In_789);
nor U1819 (N_1819,In_1971,In_2455);
nor U1820 (N_1820,In_1038,In_319);
nor U1821 (N_1821,In_1552,In_572);
nand U1822 (N_1822,In_1093,In_697);
or U1823 (N_1823,In_705,In_1226);
nand U1824 (N_1824,In_458,In_896);
nor U1825 (N_1825,In_519,In_254);
or U1826 (N_1826,In_1969,In_1435);
xor U1827 (N_1827,In_1389,In_1289);
nor U1828 (N_1828,In_1264,In_68);
xnor U1829 (N_1829,In_463,In_1276);
and U1830 (N_1830,In_182,In_1333);
and U1831 (N_1831,In_57,In_2083);
and U1832 (N_1832,In_1113,In_672);
nor U1833 (N_1833,In_1438,In_2220);
xnor U1834 (N_1834,In_1177,In_82);
and U1835 (N_1835,In_2107,In_930);
or U1836 (N_1836,In_47,In_1827);
nand U1837 (N_1837,In_1000,In_1274);
and U1838 (N_1838,In_1742,In_1484);
and U1839 (N_1839,In_2370,In_163);
nor U1840 (N_1840,In_1900,In_2460);
or U1841 (N_1841,In_804,In_628);
and U1842 (N_1842,In_545,In_2144);
and U1843 (N_1843,In_1788,In_1866);
nor U1844 (N_1844,In_83,In_1102);
and U1845 (N_1845,In_1443,In_2271);
nor U1846 (N_1846,In_623,In_624);
nand U1847 (N_1847,In_394,In_897);
nand U1848 (N_1848,In_538,In_218);
and U1849 (N_1849,In_2240,In_303);
xnor U1850 (N_1850,In_1953,In_2456);
or U1851 (N_1851,In_481,In_75);
and U1852 (N_1852,In_213,In_2025);
or U1853 (N_1853,In_705,In_2078);
and U1854 (N_1854,In_1495,In_2232);
or U1855 (N_1855,In_1850,In_851);
nand U1856 (N_1856,In_2368,In_42);
nand U1857 (N_1857,In_80,In_1506);
xor U1858 (N_1858,In_2385,In_1566);
and U1859 (N_1859,In_2046,In_303);
nor U1860 (N_1860,In_46,In_393);
or U1861 (N_1861,In_824,In_594);
nor U1862 (N_1862,In_1017,In_1998);
or U1863 (N_1863,In_1150,In_2023);
nor U1864 (N_1864,In_1933,In_2105);
nor U1865 (N_1865,In_37,In_1382);
xor U1866 (N_1866,In_812,In_720);
nor U1867 (N_1867,In_1095,In_415);
and U1868 (N_1868,In_1265,In_934);
and U1869 (N_1869,In_1893,In_2463);
nor U1870 (N_1870,In_2136,In_2285);
nor U1871 (N_1871,In_1686,In_802);
nand U1872 (N_1872,In_2233,In_1102);
nand U1873 (N_1873,In_2373,In_2091);
nor U1874 (N_1874,In_2423,In_71);
xor U1875 (N_1875,In_1415,In_1181);
or U1876 (N_1876,In_1160,In_1198);
nand U1877 (N_1877,In_912,In_59);
and U1878 (N_1878,In_1260,In_1380);
xor U1879 (N_1879,In_1748,In_2459);
and U1880 (N_1880,In_2179,In_819);
or U1881 (N_1881,In_2037,In_804);
nor U1882 (N_1882,In_2042,In_2080);
xor U1883 (N_1883,In_2293,In_962);
nor U1884 (N_1884,In_2416,In_2448);
nor U1885 (N_1885,In_1182,In_1656);
nand U1886 (N_1886,In_1099,In_690);
nand U1887 (N_1887,In_1826,In_229);
nor U1888 (N_1888,In_111,In_2092);
and U1889 (N_1889,In_552,In_64);
xor U1890 (N_1890,In_917,In_87);
nor U1891 (N_1891,In_1873,In_1137);
nor U1892 (N_1892,In_1235,In_1044);
xnor U1893 (N_1893,In_2370,In_2086);
nand U1894 (N_1894,In_110,In_919);
nand U1895 (N_1895,In_1482,In_1739);
xor U1896 (N_1896,In_1818,In_2079);
xnor U1897 (N_1897,In_1528,In_1875);
and U1898 (N_1898,In_805,In_1707);
nor U1899 (N_1899,In_1485,In_462);
and U1900 (N_1900,In_164,In_793);
or U1901 (N_1901,In_1419,In_285);
xor U1902 (N_1902,In_1595,In_427);
or U1903 (N_1903,In_1236,In_992);
nand U1904 (N_1904,In_1177,In_1443);
nor U1905 (N_1905,In_279,In_1206);
nor U1906 (N_1906,In_2193,In_1228);
or U1907 (N_1907,In_590,In_230);
or U1908 (N_1908,In_1927,In_22);
and U1909 (N_1909,In_1121,In_2150);
and U1910 (N_1910,In_2386,In_1666);
nand U1911 (N_1911,In_868,In_356);
or U1912 (N_1912,In_2201,In_1985);
or U1913 (N_1913,In_123,In_368);
and U1914 (N_1914,In_499,In_1841);
xor U1915 (N_1915,In_2414,In_1080);
or U1916 (N_1916,In_1629,In_6);
or U1917 (N_1917,In_2231,In_1624);
xor U1918 (N_1918,In_2147,In_1449);
and U1919 (N_1919,In_730,In_842);
nor U1920 (N_1920,In_789,In_104);
and U1921 (N_1921,In_1789,In_1783);
or U1922 (N_1922,In_873,In_734);
nand U1923 (N_1923,In_549,In_1062);
or U1924 (N_1924,In_2249,In_273);
nand U1925 (N_1925,In_2425,In_364);
nor U1926 (N_1926,In_1166,In_1812);
and U1927 (N_1927,In_752,In_415);
nand U1928 (N_1928,In_1948,In_1394);
or U1929 (N_1929,In_1740,In_2137);
xor U1930 (N_1930,In_1986,In_1693);
nand U1931 (N_1931,In_2497,In_391);
nand U1932 (N_1932,In_1838,In_212);
nor U1933 (N_1933,In_2459,In_784);
nor U1934 (N_1934,In_2215,In_2283);
or U1935 (N_1935,In_942,In_1335);
xnor U1936 (N_1936,In_1817,In_115);
nand U1937 (N_1937,In_911,In_698);
or U1938 (N_1938,In_991,In_1319);
nor U1939 (N_1939,In_1490,In_1681);
and U1940 (N_1940,In_490,In_866);
and U1941 (N_1941,In_1326,In_123);
nor U1942 (N_1942,In_2280,In_1119);
or U1943 (N_1943,In_268,In_508);
and U1944 (N_1944,In_204,In_1987);
or U1945 (N_1945,In_173,In_1678);
xnor U1946 (N_1946,In_867,In_249);
or U1947 (N_1947,In_1393,In_2187);
xnor U1948 (N_1948,In_1552,In_653);
nand U1949 (N_1949,In_1235,In_2021);
and U1950 (N_1950,In_1277,In_2249);
xor U1951 (N_1951,In_815,In_1612);
or U1952 (N_1952,In_395,In_1689);
nand U1953 (N_1953,In_1735,In_248);
xnor U1954 (N_1954,In_2464,In_1089);
xnor U1955 (N_1955,In_2227,In_1476);
nor U1956 (N_1956,In_1837,In_1229);
xor U1957 (N_1957,In_684,In_171);
or U1958 (N_1958,In_108,In_154);
xnor U1959 (N_1959,In_1595,In_2083);
nor U1960 (N_1960,In_1187,In_1981);
or U1961 (N_1961,In_2074,In_2357);
nor U1962 (N_1962,In_1745,In_46);
xnor U1963 (N_1963,In_1976,In_1991);
or U1964 (N_1964,In_1490,In_40);
nand U1965 (N_1965,In_1673,In_1532);
xor U1966 (N_1966,In_265,In_1648);
and U1967 (N_1967,In_968,In_2372);
and U1968 (N_1968,In_183,In_697);
nand U1969 (N_1969,In_2393,In_2023);
and U1970 (N_1970,In_426,In_1178);
nor U1971 (N_1971,In_571,In_48);
nor U1972 (N_1972,In_2339,In_2105);
and U1973 (N_1973,In_1370,In_1947);
nor U1974 (N_1974,In_246,In_389);
or U1975 (N_1975,In_1127,In_609);
and U1976 (N_1976,In_2393,In_2333);
and U1977 (N_1977,In_1397,In_492);
nand U1978 (N_1978,In_1796,In_1222);
nand U1979 (N_1979,In_2219,In_411);
or U1980 (N_1980,In_300,In_1766);
or U1981 (N_1981,In_1176,In_1518);
nor U1982 (N_1982,In_2441,In_1298);
nor U1983 (N_1983,In_1951,In_182);
nand U1984 (N_1984,In_880,In_1923);
nor U1985 (N_1985,In_1821,In_792);
nand U1986 (N_1986,In_2005,In_1995);
nand U1987 (N_1987,In_1755,In_758);
and U1988 (N_1988,In_1714,In_1238);
nand U1989 (N_1989,In_39,In_319);
or U1990 (N_1990,In_689,In_842);
xnor U1991 (N_1991,In_1011,In_1869);
nor U1992 (N_1992,In_111,In_1383);
or U1993 (N_1993,In_784,In_1240);
or U1994 (N_1994,In_1748,In_541);
nor U1995 (N_1995,In_2265,In_1577);
and U1996 (N_1996,In_1499,In_1307);
xnor U1997 (N_1997,In_2266,In_2033);
nand U1998 (N_1998,In_593,In_113);
nor U1999 (N_1999,In_45,In_1489);
and U2000 (N_2000,In_282,In_1705);
and U2001 (N_2001,In_1608,In_2263);
xor U2002 (N_2002,In_1621,In_18);
nor U2003 (N_2003,In_2097,In_661);
xor U2004 (N_2004,In_2353,In_205);
nand U2005 (N_2005,In_1958,In_1594);
nand U2006 (N_2006,In_84,In_1690);
xnor U2007 (N_2007,In_2271,In_194);
nor U2008 (N_2008,In_394,In_514);
xor U2009 (N_2009,In_439,In_1434);
xor U2010 (N_2010,In_312,In_842);
nor U2011 (N_2011,In_630,In_1034);
nor U2012 (N_2012,In_1115,In_764);
and U2013 (N_2013,In_298,In_1640);
xor U2014 (N_2014,In_1479,In_513);
and U2015 (N_2015,In_945,In_1015);
nand U2016 (N_2016,In_355,In_275);
nor U2017 (N_2017,In_1018,In_679);
nand U2018 (N_2018,In_2204,In_893);
or U2019 (N_2019,In_90,In_1177);
nor U2020 (N_2020,In_715,In_1931);
nand U2021 (N_2021,In_1876,In_894);
and U2022 (N_2022,In_506,In_1440);
xnor U2023 (N_2023,In_34,In_768);
nand U2024 (N_2024,In_1969,In_2064);
and U2025 (N_2025,In_526,In_1837);
xor U2026 (N_2026,In_2353,In_341);
or U2027 (N_2027,In_917,In_841);
or U2028 (N_2028,In_1230,In_1595);
and U2029 (N_2029,In_2146,In_601);
nor U2030 (N_2030,In_1635,In_113);
xor U2031 (N_2031,In_534,In_774);
nor U2032 (N_2032,In_1324,In_1411);
nand U2033 (N_2033,In_561,In_337);
nand U2034 (N_2034,In_1029,In_260);
nor U2035 (N_2035,In_2068,In_285);
nand U2036 (N_2036,In_266,In_1169);
xor U2037 (N_2037,In_732,In_1251);
nand U2038 (N_2038,In_1049,In_986);
and U2039 (N_2039,In_336,In_903);
or U2040 (N_2040,In_2192,In_707);
nor U2041 (N_2041,In_1340,In_2139);
nor U2042 (N_2042,In_2473,In_431);
nor U2043 (N_2043,In_2182,In_2227);
nor U2044 (N_2044,In_886,In_455);
nor U2045 (N_2045,In_1314,In_482);
or U2046 (N_2046,In_844,In_943);
xnor U2047 (N_2047,In_1200,In_1934);
xnor U2048 (N_2048,In_566,In_857);
or U2049 (N_2049,In_904,In_1729);
or U2050 (N_2050,In_2134,In_147);
and U2051 (N_2051,In_85,In_1683);
xor U2052 (N_2052,In_534,In_2478);
nand U2053 (N_2053,In_269,In_1627);
nor U2054 (N_2054,In_867,In_598);
nor U2055 (N_2055,In_1753,In_422);
nor U2056 (N_2056,In_347,In_782);
and U2057 (N_2057,In_1815,In_1853);
or U2058 (N_2058,In_307,In_2185);
and U2059 (N_2059,In_1507,In_2182);
nand U2060 (N_2060,In_860,In_2412);
or U2061 (N_2061,In_2218,In_28);
nor U2062 (N_2062,In_201,In_72);
nand U2063 (N_2063,In_2324,In_1445);
nor U2064 (N_2064,In_941,In_2332);
or U2065 (N_2065,In_828,In_406);
or U2066 (N_2066,In_2418,In_1581);
and U2067 (N_2067,In_570,In_78);
nand U2068 (N_2068,In_2069,In_803);
nor U2069 (N_2069,In_1489,In_2209);
nand U2070 (N_2070,In_2198,In_2363);
xor U2071 (N_2071,In_291,In_85);
xnor U2072 (N_2072,In_2163,In_890);
or U2073 (N_2073,In_2231,In_1132);
xnor U2074 (N_2074,In_1183,In_1171);
or U2075 (N_2075,In_1631,In_1178);
and U2076 (N_2076,In_239,In_308);
nand U2077 (N_2077,In_630,In_406);
nor U2078 (N_2078,In_368,In_2280);
or U2079 (N_2079,In_916,In_1310);
nor U2080 (N_2080,In_1974,In_1216);
nor U2081 (N_2081,In_49,In_25);
nand U2082 (N_2082,In_686,In_20);
nand U2083 (N_2083,In_1583,In_1457);
nand U2084 (N_2084,In_1320,In_405);
nand U2085 (N_2085,In_2396,In_4);
and U2086 (N_2086,In_316,In_1631);
nor U2087 (N_2087,In_344,In_1792);
nor U2088 (N_2088,In_1806,In_994);
and U2089 (N_2089,In_1750,In_1959);
or U2090 (N_2090,In_2278,In_1617);
nor U2091 (N_2091,In_2080,In_756);
or U2092 (N_2092,In_162,In_1298);
or U2093 (N_2093,In_2192,In_1812);
and U2094 (N_2094,In_1469,In_2012);
xnor U2095 (N_2095,In_542,In_981);
xnor U2096 (N_2096,In_1311,In_2495);
xor U2097 (N_2097,In_509,In_1746);
and U2098 (N_2098,In_477,In_128);
nor U2099 (N_2099,In_789,In_1310);
nor U2100 (N_2100,In_77,In_2089);
nand U2101 (N_2101,In_170,In_1016);
nand U2102 (N_2102,In_1626,In_905);
or U2103 (N_2103,In_1083,In_640);
or U2104 (N_2104,In_1365,In_1539);
and U2105 (N_2105,In_326,In_2252);
or U2106 (N_2106,In_721,In_1112);
and U2107 (N_2107,In_271,In_1985);
nor U2108 (N_2108,In_1148,In_1915);
and U2109 (N_2109,In_577,In_165);
or U2110 (N_2110,In_195,In_651);
nand U2111 (N_2111,In_2211,In_1041);
nand U2112 (N_2112,In_1262,In_2368);
and U2113 (N_2113,In_1858,In_1331);
or U2114 (N_2114,In_908,In_2476);
and U2115 (N_2115,In_2499,In_385);
and U2116 (N_2116,In_1884,In_2125);
nand U2117 (N_2117,In_253,In_1829);
nand U2118 (N_2118,In_132,In_140);
and U2119 (N_2119,In_1901,In_998);
xnor U2120 (N_2120,In_107,In_48);
or U2121 (N_2121,In_2421,In_1469);
xor U2122 (N_2122,In_2287,In_1553);
xor U2123 (N_2123,In_532,In_1550);
xor U2124 (N_2124,In_759,In_1471);
or U2125 (N_2125,In_313,In_886);
nand U2126 (N_2126,In_1699,In_616);
xor U2127 (N_2127,In_451,In_1682);
nor U2128 (N_2128,In_830,In_144);
nor U2129 (N_2129,In_137,In_1681);
xor U2130 (N_2130,In_1038,In_1051);
nor U2131 (N_2131,In_959,In_1802);
and U2132 (N_2132,In_1058,In_424);
nor U2133 (N_2133,In_1541,In_2034);
or U2134 (N_2134,In_1985,In_1879);
or U2135 (N_2135,In_1186,In_1840);
and U2136 (N_2136,In_1719,In_381);
and U2137 (N_2137,In_1965,In_903);
nor U2138 (N_2138,In_227,In_1420);
or U2139 (N_2139,In_625,In_420);
nor U2140 (N_2140,In_883,In_1445);
nand U2141 (N_2141,In_2162,In_905);
and U2142 (N_2142,In_2314,In_1773);
nand U2143 (N_2143,In_230,In_2267);
nand U2144 (N_2144,In_180,In_593);
or U2145 (N_2145,In_1335,In_2180);
nand U2146 (N_2146,In_1095,In_728);
xor U2147 (N_2147,In_673,In_671);
and U2148 (N_2148,In_329,In_389);
xor U2149 (N_2149,In_1050,In_746);
or U2150 (N_2150,In_618,In_1598);
nand U2151 (N_2151,In_2407,In_370);
nand U2152 (N_2152,In_332,In_995);
nand U2153 (N_2153,In_2077,In_2367);
nor U2154 (N_2154,In_1470,In_1048);
xnor U2155 (N_2155,In_2448,In_68);
nor U2156 (N_2156,In_80,In_528);
nand U2157 (N_2157,In_1041,In_2205);
nor U2158 (N_2158,In_78,In_2179);
and U2159 (N_2159,In_72,In_1014);
nand U2160 (N_2160,In_2072,In_1718);
nand U2161 (N_2161,In_1486,In_1201);
nor U2162 (N_2162,In_1574,In_1414);
nor U2163 (N_2163,In_1169,In_1505);
or U2164 (N_2164,In_1413,In_2313);
xnor U2165 (N_2165,In_2082,In_1777);
nor U2166 (N_2166,In_199,In_1660);
xor U2167 (N_2167,In_2110,In_2317);
xnor U2168 (N_2168,In_1640,In_1660);
xor U2169 (N_2169,In_1890,In_1267);
and U2170 (N_2170,In_1383,In_1028);
nand U2171 (N_2171,In_2085,In_262);
nand U2172 (N_2172,In_1042,In_1862);
or U2173 (N_2173,In_500,In_382);
nand U2174 (N_2174,In_14,In_123);
nor U2175 (N_2175,In_81,In_1815);
xor U2176 (N_2176,In_2374,In_1516);
or U2177 (N_2177,In_2246,In_1674);
and U2178 (N_2178,In_1442,In_2497);
nor U2179 (N_2179,In_1133,In_2111);
and U2180 (N_2180,In_1043,In_2307);
xnor U2181 (N_2181,In_1575,In_1571);
nor U2182 (N_2182,In_1779,In_43);
nand U2183 (N_2183,In_1455,In_140);
nor U2184 (N_2184,In_57,In_2471);
and U2185 (N_2185,In_2048,In_1831);
or U2186 (N_2186,In_1945,In_922);
xnor U2187 (N_2187,In_567,In_135);
or U2188 (N_2188,In_492,In_2385);
nor U2189 (N_2189,In_2005,In_124);
nand U2190 (N_2190,In_639,In_558);
nor U2191 (N_2191,In_724,In_1968);
or U2192 (N_2192,In_1726,In_249);
xnor U2193 (N_2193,In_1759,In_1852);
nand U2194 (N_2194,In_2363,In_1263);
xor U2195 (N_2195,In_2005,In_220);
xor U2196 (N_2196,In_2141,In_505);
xnor U2197 (N_2197,In_1951,In_2090);
nor U2198 (N_2198,In_1860,In_709);
or U2199 (N_2199,In_1591,In_1364);
xor U2200 (N_2200,In_2492,In_355);
xnor U2201 (N_2201,In_993,In_267);
and U2202 (N_2202,In_1698,In_4);
xor U2203 (N_2203,In_291,In_2348);
or U2204 (N_2204,In_2158,In_499);
nor U2205 (N_2205,In_1984,In_1412);
and U2206 (N_2206,In_403,In_716);
nand U2207 (N_2207,In_396,In_2323);
xor U2208 (N_2208,In_237,In_2443);
and U2209 (N_2209,In_2257,In_900);
or U2210 (N_2210,In_174,In_855);
and U2211 (N_2211,In_1321,In_646);
nand U2212 (N_2212,In_250,In_73);
nor U2213 (N_2213,In_262,In_1665);
xor U2214 (N_2214,In_1966,In_408);
xor U2215 (N_2215,In_839,In_1486);
xnor U2216 (N_2216,In_1728,In_1082);
nor U2217 (N_2217,In_70,In_2477);
nand U2218 (N_2218,In_1072,In_462);
nand U2219 (N_2219,In_1243,In_1424);
nand U2220 (N_2220,In_452,In_958);
or U2221 (N_2221,In_59,In_1751);
nor U2222 (N_2222,In_2291,In_1370);
and U2223 (N_2223,In_483,In_1091);
xor U2224 (N_2224,In_1649,In_1811);
or U2225 (N_2225,In_1426,In_1303);
nor U2226 (N_2226,In_2218,In_1136);
nand U2227 (N_2227,In_1787,In_1080);
nor U2228 (N_2228,In_1309,In_1064);
and U2229 (N_2229,In_2075,In_2185);
xnor U2230 (N_2230,In_278,In_1136);
xnor U2231 (N_2231,In_1482,In_1214);
and U2232 (N_2232,In_526,In_1466);
and U2233 (N_2233,In_2161,In_1334);
nor U2234 (N_2234,In_1653,In_1564);
xnor U2235 (N_2235,In_390,In_1229);
and U2236 (N_2236,In_143,In_1298);
or U2237 (N_2237,In_621,In_945);
nand U2238 (N_2238,In_1033,In_923);
and U2239 (N_2239,In_1289,In_97);
nor U2240 (N_2240,In_1896,In_565);
nor U2241 (N_2241,In_453,In_367);
or U2242 (N_2242,In_1106,In_2010);
and U2243 (N_2243,In_2100,In_411);
or U2244 (N_2244,In_1832,In_1912);
nand U2245 (N_2245,In_1067,In_940);
xnor U2246 (N_2246,In_182,In_1605);
nand U2247 (N_2247,In_2454,In_1081);
nor U2248 (N_2248,In_1395,In_1553);
xnor U2249 (N_2249,In_1182,In_539);
and U2250 (N_2250,In_288,In_1053);
and U2251 (N_2251,In_1614,In_2198);
xnor U2252 (N_2252,In_457,In_1979);
or U2253 (N_2253,In_183,In_1922);
and U2254 (N_2254,In_173,In_990);
or U2255 (N_2255,In_442,In_644);
and U2256 (N_2256,In_1435,In_861);
nor U2257 (N_2257,In_885,In_1273);
or U2258 (N_2258,In_1368,In_225);
nor U2259 (N_2259,In_1686,In_1023);
and U2260 (N_2260,In_410,In_1893);
xor U2261 (N_2261,In_1711,In_2111);
or U2262 (N_2262,In_1110,In_1446);
nand U2263 (N_2263,In_724,In_733);
and U2264 (N_2264,In_810,In_2487);
and U2265 (N_2265,In_411,In_2351);
nor U2266 (N_2266,In_2350,In_1917);
xor U2267 (N_2267,In_864,In_897);
nor U2268 (N_2268,In_1607,In_2183);
nor U2269 (N_2269,In_1101,In_763);
nand U2270 (N_2270,In_452,In_2266);
nand U2271 (N_2271,In_1191,In_1102);
nand U2272 (N_2272,In_1878,In_2482);
or U2273 (N_2273,In_294,In_1192);
xor U2274 (N_2274,In_2154,In_1530);
xnor U2275 (N_2275,In_2105,In_292);
and U2276 (N_2276,In_340,In_1579);
nand U2277 (N_2277,In_748,In_858);
nor U2278 (N_2278,In_2167,In_613);
nand U2279 (N_2279,In_63,In_488);
nor U2280 (N_2280,In_1,In_2426);
or U2281 (N_2281,In_1881,In_1434);
and U2282 (N_2282,In_2334,In_1347);
nor U2283 (N_2283,In_661,In_923);
and U2284 (N_2284,In_905,In_509);
and U2285 (N_2285,In_1249,In_149);
and U2286 (N_2286,In_855,In_1688);
and U2287 (N_2287,In_1537,In_1364);
nor U2288 (N_2288,In_1292,In_1031);
or U2289 (N_2289,In_891,In_2486);
and U2290 (N_2290,In_1223,In_2030);
xnor U2291 (N_2291,In_1986,In_1665);
or U2292 (N_2292,In_274,In_745);
nor U2293 (N_2293,In_576,In_1875);
nor U2294 (N_2294,In_1254,In_1869);
or U2295 (N_2295,In_230,In_2235);
nor U2296 (N_2296,In_1699,In_1027);
nor U2297 (N_2297,In_1211,In_482);
and U2298 (N_2298,In_195,In_989);
nor U2299 (N_2299,In_512,In_1360);
or U2300 (N_2300,In_1143,In_417);
and U2301 (N_2301,In_1620,In_1680);
or U2302 (N_2302,In_2257,In_1115);
and U2303 (N_2303,In_254,In_343);
nor U2304 (N_2304,In_1342,In_2327);
or U2305 (N_2305,In_2191,In_658);
and U2306 (N_2306,In_53,In_834);
and U2307 (N_2307,In_879,In_2241);
nand U2308 (N_2308,In_1531,In_268);
nand U2309 (N_2309,In_290,In_2041);
nor U2310 (N_2310,In_1126,In_879);
xnor U2311 (N_2311,In_796,In_1350);
nand U2312 (N_2312,In_2335,In_716);
nand U2313 (N_2313,In_2148,In_1945);
nor U2314 (N_2314,In_558,In_2133);
and U2315 (N_2315,In_2083,In_1350);
nand U2316 (N_2316,In_470,In_1815);
nor U2317 (N_2317,In_325,In_2289);
nand U2318 (N_2318,In_467,In_1536);
and U2319 (N_2319,In_458,In_2326);
or U2320 (N_2320,In_411,In_151);
and U2321 (N_2321,In_1120,In_275);
nor U2322 (N_2322,In_390,In_1663);
xor U2323 (N_2323,In_311,In_878);
xnor U2324 (N_2324,In_1430,In_546);
xnor U2325 (N_2325,In_1460,In_251);
nand U2326 (N_2326,In_1671,In_223);
nor U2327 (N_2327,In_259,In_11);
nand U2328 (N_2328,In_1459,In_1700);
or U2329 (N_2329,In_1624,In_165);
xor U2330 (N_2330,In_1135,In_878);
or U2331 (N_2331,In_220,In_1698);
or U2332 (N_2332,In_1731,In_2160);
nor U2333 (N_2333,In_1338,In_891);
or U2334 (N_2334,In_64,In_1945);
nand U2335 (N_2335,In_1902,In_740);
and U2336 (N_2336,In_1605,In_1299);
and U2337 (N_2337,In_391,In_1636);
nor U2338 (N_2338,In_1093,In_5);
nor U2339 (N_2339,In_2308,In_351);
nor U2340 (N_2340,In_1079,In_2437);
xnor U2341 (N_2341,In_450,In_1687);
or U2342 (N_2342,In_630,In_695);
or U2343 (N_2343,In_1740,In_1736);
xnor U2344 (N_2344,In_1971,In_926);
nand U2345 (N_2345,In_118,In_1214);
or U2346 (N_2346,In_124,In_2036);
nor U2347 (N_2347,In_1756,In_872);
nand U2348 (N_2348,In_2076,In_1133);
and U2349 (N_2349,In_1788,In_98);
xor U2350 (N_2350,In_1956,In_65);
nand U2351 (N_2351,In_2125,In_2485);
nor U2352 (N_2352,In_329,In_182);
or U2353 (N_2353,In_1818,In_1930);
or U2354 (N_2354,In_519,In_857);
nand U2355 (N_2355,In_633,In_566);
or U2356 (N_2356,In_1877,In_1726);
nand U2357 (N_2357,In_1560,In_1180);
or U2358 (N_2358,In_1156,In_115);
nor U2359 (N_2359,In_419,In_1386);
or U2360 (N_2360,In_711,In_977);
and U2361 (N_2361,In_1402,In_887);
and U2362 (N_2362,In_2419,In_2457);
nor U2363 (N_2363,In_845,In_2024);
and U2364 (N_2364,In_2199,In_1023);
xor U2365 (N_2365,In_1936,In_1315);
xor U2366 (N_2366,In_1234,In_2245);
nor U2367 (N_2367,In_909,In_1515);
or U2368 (N_2368,In_995,In_1120);
xor U2369 (N_2369,In_2280,In_1554);
nor U2370 (N_2370,In_2303,In_2299);
and U2371 (N_2371,In_1092,In_1203);
nor U2372 (N_2372,In_2179,In_1423);
nand U2373 (N_2373,In_2474,In_1210);
and U2374 (N_2374,In_2095,In_1385);
nand U2375 (N_2375,In_1122,In_87);
nand U2376 (N_2376,In_2178,In_2210);
nor U2377 (N_2377,In_709,In_2460);
nor U2378 (N_2378,In_2216,In_1067);
or U2379 (N_2379,In_894,In_1507);
and U2380 (N_2380,In_2066,In_706);
nor U2381 (N_2381,In_1204,In_136);
and U2382 (N_2382,In_146,In_1019);
nor U2383 (N_2383,In_816,In_460);
or U2384 (N_2384,In_2481,In_542);
nand U2385 (N_2385,In_1483,In_265);
nand U2386 (N_2386,In_983,In_811);
nor U2387 (N_2387,In_1811,In_2010);
or U2388 (N_2388,In_1295,In_38);
nand U2389 (N_2389,In_2258,In_645);
or U2390 (N_2390,In_1614,In_1949);
xor U2391 (N_2391,In_1586,In_1422);
or U2392 (N_2392,In_1555,In_1744);
nor U2393 (N_2393,In_1590,In_288);
or U2394 (N_2394,In_593,In_205);
nand U2395 (N_2395,In_1659,In_1988);
xnor U2396 (N_2396,In_748,In_341);
nor U2397 (N_2397,In_386,In_1938);
xnor U2398 (N_2398,In_1687,In_2400);
xor U2399 (N_2399,In_1996,In_158);
or U2400 (N_2400,In_424,In_1424);
nand U2401 (N_2401,In_1960,In_1962);
or U2402 (N_2402,In_1385,In_922);
xor U2403 (N_2403,In_830,In_1111);
or U2404 (N_2404,In_2388,In_2455);
xnor U2405 (N_2405,In_1448,In_2195);
xnor U2406 (N_2406,In_1106,In_2148);
or U2407 (N_2407,In_1828,In_1625);
nand U2408 (N_2408,In_443,In_654);
nand U2409 (N_2409,In_2050,In_941);
and U2410 (N_2410,In_2236,In_942);
nor U2411 (N_2411,In_29,In_2183);
nor U2412 (N_2412,In_2067,In_1504);
and U2413 (N_2413,In_1759,In_794);
xnor U2414 (N_2414,In_223,In_2052);
nor U2415 (N_2415,In_1561,In_743);
nand U2416 (N_2416,In_2455,In_572);
and U2417 (N_2417,In_2434,In_460);
or U2418 (N_2418,In_1065,In_19);
or U2419 (N_2419,In_144,In_798);
or U2420 (N_2420,In_560,In_2147);
nand U2421 (N_2421,In_6,In_427);
nor U2422 (N_2422,In_256,In_459);
xor U2423 (N_2423,In_1110,In_339);
nor U2424 (N_2424,In_687,In_1593);
nand U2425 (N_2425,In_1040,In_1070);
xor U2426 (N_2426,In_416,In_1110);
and U2427 (N_2427,In_785,In_2331);
nor U2428 (N_2428,In_829,In_1300);
xnor U2429 (N_2429,In_2488,In_2332);
nand U2430 (N_2430,In_457,In_2186);
or U2431 (N_2431,In_992,In_1105);
or U2432 (N_2432,In_2266,In_2220);
or U2433 (N_2433,In_1625,In_1427);
nand U2434 (N_2434,In_2307,In_1831);
nand U2435 (N_2435,In_2328,In_628);
or U2436 (N_2436,In_1624,In_1639);
nand U2437 (N_2437,In_711,In_1103);
nand U2438 (N_2438,In_23,In_1943);
nor U2439 (N_2439,In_748,In_1972);
and U2440 (N_2440,In_2222,In_2042);
xnor U2441 (N_2441,In_1480,In_380);
nand U2442 (N_2442,In_1381,In_669);
nand U2443 (N_2443,In_308,In_1173);
xor U2444 (N_2444,In_2149,In_1374);
nor U2445 (N_2445,In_1340,In_111);
nand U2446 (N_2446,In_1433,In_1523);
and U2447 (N_2447,In_2103,In_162);
xnor U2448 (N_2448,In_143,In_267);
nor U2449 (N_2449,In_547,In_1363);
and U2450 (N_2450,In_744,In_1918);
or U2451 (N_2451,In_520,In_726);
nor U2452 (N_2452,In_1042,In_1230);
or U2453 (N_2453,In_410,In_1122);
nand U2454 (N_2454,In_629,In_1525);
xor U2455 (N_2455,In_738,In_1591);
nand U2456 (N_2456,In_1238,In_911);
and U2457 (N_2457,In_830,In_531);
nand U2458 (N_2458,In_2381,In_1905);
nor U2459 (N_2459,In_792,In_585);
or U2460 (N_2460,In_494,In_101);
nand U2461 (N_2461,In_2464,In_1525);
nor U2462 (N_2462,In_346,In_181);
nor U2463 (N_2463,In_1788,In_453);
and U2464 (N_2464,In_1238,In_2006);
or U2465 (N_2465,In_1414,In_290);
nand U2466 (N_2466,In_1600,In_1203);
nand U2467 (N_2467,In_220,In_1893);
xor U2468 (N_2468,In_361,In_588);
or U2469 (N_2469,In_2004,In_817);
nor U2470 (N_2470,In_34,In_1701);
or U2471 (N_2471,In_1367,In_1530);
nand U2472 (N_2472,In_1147,In_302);
or U2473 (N_2473,In_1872,In_1531);
nand U2474 (N_2474,In_1405,In_241);
xor U2475 (N_2475,In_669,In_189);
xnor U2476 (N_2476,In_2326,In_2441);
or U2477 (N_2477,In_943,In_2169);
and U2478 (N_2478,In_2390,In_2181);
nor U2479 (N_2479,In_1991,In_675);
or U2480 (N_2480,In_1375,In_813);
nor U2481 (N_2481,In_169,In_2437);
nor U2482 (N_2482,In_850,In_2067);
and U2483 (N_2483,In_352,In_1113);
nor U2484 (N_2484,In_650,In_1803);
nor U2485 (N_2485,In_346,In_2051);
or U2486 (N_2486,In_1842,In_1691);
or U2487 (N_2487,In_1357,In_1355);
nor U2488 (N_2488,In_681,In_1954);
and U2489 (N_2489,In_19,In_1048);
and U2490 (N_2490,In_2071,In_1514);
xor U2491 (N_2491,In_2241,In_2441);
nor U2492 (N_2492,In_1882,In_2426);
nand U2493 (N_2493,In_1803,In_1358);
or U2494 (N_2494,In_1386,In_1100);
and U2495 (N_2495,In_2028,In_589);
nor U2496 (N_2496,In_720,In_2116);
nand U2497 (N_2497,In_269,In_1609);
xor U2498 (N_2498,In_811,In_1696);
nor U2499 (N_2499,In_935,In_1441);
or U2500 (N_2500,In_56,In_1576);
nand U2501 (N_2501,In_1549,In_1907);
xor U2502 (N_2502,In_149,In_2378);
or U2503 (N_2503,In_2354,In_872);
and U2504 (N_2504,In_391,In_1989);
and U2505 (N_2505,In_2338,In_1679);
nor U2506 (N_2506,In_1838,In_845);
nand U2507 (N_2507,In_517,In_1417);
nor U2508 (N_2508,In_154,In_510);
or U2509 (N_2509,In_1356,In_1347);
and U2510 (N_2510,In_1048,In_1287);
nor U2511 (N_2511,In_227,In_1298);
or U2512 (N_2512,In_1557,In_52);
and U2513 (N_2513,In_1169,In_1435);
xor U2514 (N_2514,In_2205,In_1968);
and U2515 (N_2515,In_1594,In_1100);
nor U2516 (N_2516,In_1434,In_1774);
or U2517 (N_2517,In_2203,In_2038);
and U2518 (N_2518,In_1483,In_1903);
nand U2519 (N_2519,In_1673,In_635);
nor U2520 (N_2520,In_489,In_768);
and U2521 (N_2521,In_1444,In_1614);
and U2522 (N_2522,In_2220,In_2278);
xnor U2523 (N_2523,In_2315,In_1428);
xnor U2524 (N_2524,In_978,In_1015);
nand U2525 (N_2525,In_44,In_2440);
xor U2526 (N_2526,In_736,In_1566);
xor U2527 (N_2527,In_281,In_2497);
nand U2528 (N_2528,In_709,In_361);
nor U2529 (N_2529,In_2234,In_530);
and U2530 (N_2530,In_1163,In_623);
xnor U2531 (N_2531,In_1415,In_1040);
nand U2532 (N_2532,In_1174,In_569);
xor U2533 (N_2533,In_379,In_2023);
nand U2534 (N_2534,In_543,In_970);
nor U2535 (N_2535,In_2245,In_1376);
or U2536 (N_2536,In_2290,In_1522);
nand U2537 (N_2537,In_715,In_2402);
nand U2538 (N_2538,In_702,In_1497);
or U2539 (N_2539,In_1405,In_2424);
and U2540 (N_2540,In_597,In_351);
and U2541 (N_2541,In_2024,In_2460);
nand U2542 (N_2542,In_75,In_2235);
or U2543 (N_2543,In_372,In_979);
or U2544 (N_2544,In_764,In_93);
nand U2545 (N_2545,In_353,In_2454);
nand U2546 (N_2546,In_1047,In_1786);
nor U2547 (N_2547,In_1831,In_193);
xor U2548 (N_2548,In_73,In_184);
nand U2549 (N_2549,In_2384,In_1948);
or U2550 (N_2550,In_1276,In_1819);
nor U2551 (N_2551,In_383,In_790);
nor U2552 (N_2552,In_1421,In_816);
xor U2553 (N_2553,In_883,In_1909);
nand U2554 (N_2554,In_2437,In_1608);
nand U2555 (N_2555,In_518,In_1355);
nand U2556 (N_2556,In_700,In_1648);
xnor U2557 (N_2557,In_1835,In_2488);
or U2558 (N_2558,In_1679,In_1341);
nor U2559 (N_2559,In_2306,In_1394);
xnor U2560 (N_2560,In_770,In_697);
or U2561 (N_2561,In_1002,In_2126);
and U2562 (N_2562,In_2060,In_344);
nor U2563 (N_2563,In_33,In_685);
nand U2564 (N_2564,In_1484,In_698);
xnor U2565 (N_2565,In_321,In_2298);
xor U2566 (N_2566,In_678,In_2447);
xor U2567 (N_2567,In_760,In_819);
or U2568 (N_2568,In_1976,In_2070);
nand U2569 (N_2569,In_414,In_1745);
or U2570 (N_2570,In_2013,In_233);
and U2571 (N_2571,In_1013,In_1108);
and U2572 (N_2572,In_1318,In_113);
nand U2573 (N_2573,In_1992,In_627);
and U2574 (N_2574,In_1119,In_416);
xnor U2575 (N_2575,In_183,In_332);
or U2576 (N_2576,In_1806,In_2396);
and U2577 (N_2577,In_1556,In_424);
xor U2578 (N_2578,In_1512,In_914);
nand U2579 (N_2579,In_36,In_679);
nor U2580 (N_2580,In_185,In_1971);
nand U2581 (N_2581,In_853,In_605);
nor U2582 (N_2582,In_1916,In_689);
and U2583 (N_2583,In_1640,In_1212);
nand U2584 (N_2584,In_1691,In_1713);
nor U2585 (N_2585,In_1200,In_860);
xor U2586 (N_2586,In_1709,In_2412);
and U2587 (N_2587,In_2171,In_633);
nor U2588 (N_2588,In_2342,In_400);
nor U2589 (N_2589,In_1287,In_554);
and U2590 (N_2590,In_1825,In_598);
xor U2591 (N_2591,In_2203,In_1818);
or U2592 (N_2592,In_628,In_1201);
and U2593 (N_2593,In_206,In_866);
and U2594 (N_2594,In_1404,In_1317);
xnor U2595 (N_2595,In_165,In_624);
and U2596 (N_2596,In_422,In_1906);
or U2597 (N_2597,In_295,In_1772);
nor U2598 (N_2598,In_1682,In_836);
xor U2599 (N_2599,In_1335,In_133);
nand U2600 (N_2600,In_548,In_2009);
nand U2601 (N_2601,In_1913,In_1641);
xnor U2602 (N_2602,In_480,In_1368);
nand U2603 (N_2603,In_2035,In_2149);
or U2604 (N_2604,In_1926,In_231);
or U2605 (N_2605,In_275,In_770);
and U2606 (N_2606,In_209,In_1676);
nor U2607 (N_2607,In_439,In_1740);
xnor U2608 (N_2608,In_207,In_952);
xnor U2609 (N_2609,In_1130,In_271);
nand U2610 (N_2610,In_1055,In_1723);
or U2611 (N_2611,In_592,In_2167);
nor U2612 (N_2612,In_2055,In_701);
xnor U2613 (N_2613,In_2338,In_2462);
xor U2614 (N_2614,In_20,In_125);
and U2615 (N_2615,In_229,In_1);
or U2616 (N_2616,In_1048,In_2225);
and U2617 (N_2617,In_1336,In_2081);
xor U2618 (N_2618,In_51,In_498);
nand U2619 (N_2619,In_1464,In_1664);
nand U2620 (N_2620,In_853,In_1131);
xor U2621 (N_2621,In_784,In_128);
and U2622 (N_2622,In_308,In_950);
nand U2623 (N_2623,In_2223,In_350);
xnor U2624 (N_2624,In_1447,In_652);
and U2625 (N_2625,In_152,In_384);
nand U2626 (N_2626,In_1590,In_844);
xor U2627 (N_2627,In_1402,In_51);
nand U2628 (N_2628,In_2070,In_406);
nor U2629 (N_2629,In_754,In_1641);
xnor U2630 (N_2630,In_1587,In_494);
xor U2631 (N_2631,In_1905,In_443);
and U2632 (N_2632,In_621,In_799);
and U2633 (N_2633,In_1163,In_2356);
or U2634 (N_2634,In_2148,In_2472);
and U2635 (N_2635,In_547,In_74);
or U2636 (N_2636,In_1337,In_1335);
and U2637 (N_2637,In_1620,In_1290);
xor U2638 (N_2638,In_508,In_1966);
nand U2639 (N_2639,In_2094,In_1517);
nor U2640 (N_2640,In_299,In_417);
nor U2641 (N_2641,In_2004,In_730);
xnor U2642 (N_2642,In_446,In_1547);
xnor U2643 (N_2643,In_333,In_708);
or U2644 (N_2644,In_2026,In_1912);
or U2645 (N_2645,In_1631,In_595);
nand U2646 (N_2646,In_1751,In_2162);
nor U2647 (N_2647,In_1978,In_390);
nand U2648 (N_2648,In_1988,In_1854);
nand U2649 (N_2649,In_1960,In_3);
and U2650 (N_2650,In_964,In_166);
or U2651 (N_2651,In_1560,In_1193);
xor U2652 (N_2652,In_619,In_1623);
or U2653 (N_2653,In_609,In_689);
or U2654 (N_2654,In_1661,In_475);
and U2655 (N_2655,In_831,In_1588);
and U2656 (N_2656,In_1360,In_1100);
nor U2657 (N_2657,In_1492,In_651);
or U2658 (N_2658,In_2402,In_1645);
and U2659 (N_2659,In_1952,In_2099);
and U2660 (N_2660,In_1055,In_744);
nand U2661 (N_2661,In_1495,In_1415);
nor U2662 (N_2662,In_492,In_135);
nor U2663 (N_2663,In_2210,In_2017);
xnor U2664 (N_2664,In_945,In_1453);
nand U2665 (N_2665,In_356,In_1311);
nor U2666 (N_2666,In_55,In_757);
nor U2667 (N_2667,In_1031,In_933);
or U2668 (N_2668,In_1515,In_716);
or U2669 (N_2669,In_1574,In_1965);
xnor U2670 (N_2670,In_469,In_1113);
nand U2671 (N_2671,In_2056,In_521);
xnor U2672 (N_2672,In_1250,In_120);
or U2673 (N_2673,In_2094,In_39);
or U2674 (N_2674,In_1065,In_1279);
nand U2675 (N_2675,In_2136,In_197);
nand U2676 (N_2676,In_277,In_2162);
xor U2677 (N_2677,In_1845,In_213);
nand U2678 (N_2678,In_2418,In_1935);
nand U2679 (N_2679,In_1244,In_487);
nor U2680 (N_2680,In_2134,In_1647);
nand U2681 (N_2681,In_1150,In_1691);
nand U2682 (N_2682,In_2065,In_2355);
nand U2683 (N_2683,In_2361,In_891);
nor U2684 (N_2684,In_226,In_51);
xor U2685 (N_2685,In_453,In_1042);
nor U2686 (N_2686,In_913,In_71);
nor U2687 (N_2687,In_691,In_1674);
nor U2688 (N_2688,In_1487,In_617);
nand U2689 (N_2689,In_2296,In_782);
nor U2690 (N_2690,In_1854,In_233);
and U2691 (N_2691,In_586,In_876);
nor U2692 (N_2692,In_467,In_1181);
nand U2693 (N_2693,In_2424,In_2328);
xor U2694 (N_2694,In_506,In_591);
nand U2695 (N_2695,In_1182,In_553);
nor U2696 (N_2696,In_262,In_896);
nand U2697 (N_2697,In_940,In_1930);
xor U2698 (N_2698,In_387,In_2441);
and U2699 (N_2699,In_1749,In_1914);
xor U2700 (N_2700,In_70,In_727);
or U2701 (N_2701,In_394,In_1162);
xor U2702 (N_2702,In_1553,In_611);
nand U2703 (N_2703,In_338,In_1746);
nor U2704 (N_2704,In_1537,In_1886);
nor U2705 (N_2705,In_387,In_1030);
or U2706 (N_2706,In_213,In_993);
and U2707 (N_2707,In_685,In_1993);
or U2708 (N_2708,In_912,In_196);
or U2709 (N_2709,In_1114,In_2023);
or U2710 (N_2710,In_1943,In_1889);
nand U2711 (N_2711,In_341,In_1494);
and U2712 (N_2712,In_2316,In_1360);
xnor U2713 (N_2713,In_1903,In_472);
and U2714 (N_2714,In_2235,In_2271);
nand U2715 (N_2715,In_1523,In_2181);
nor U2716 (N_2716,In_641,In_2252);
nor U2717 (N_2717,In_1794,In_2229);
or U2718 (N_2718,In_695,In_2324);
xnor U2719 (N_2719,In_2304,In_1603);
nand U2720 (N_2720,In_2197,In_199);
nor U2721 (N_2721,In_1754,In_2075);
xor U2722 (N_2722,In_2221,In_2328);
nor U2723 (N_2723,In_93,In_2287);
nand U2724 (N_2724,In_1882,In_1006);
or U2725 (N_2725,In_555,In_881);
or U2726 (N_2726,In_2268,In_90);
nor U2727 (N_2727,In_527,In_1820);
and U2728 (N_2728,In_221,In_1702);
nand U2729 (N_2729,In_780,In_1903);
xor U2730 (N_2730,In_1404,In_876);
xor U2731 (N_2731,In_2290,In_1500);
and U2732 (N_2732,In_1826,In_1559);
xnor U2733 (N_2733,In_1454,In_578);
or U2734 (N_2734,In_2055,In_559);
nand U2735 (N_2735,In_763,In_939);
nor U2736 (N_2736,In_6,In_2200);
nand U2737 (N_2737,In_2463,In_2314);
or U2738 (N_2738,In_1721,In_2067);
xnor U2739 (N_2739,In_1623,In_1573);
xor U2740 (N_2740,In_1743,In_850);
or U2741 (N_2741,In_1939,In_225);
nand U2742 (N_2742,In_57,In_1167);
nand U2743 (N_2743,In_1152,In_260);
nor U2744 (N_2744,In_2340,In_2054);
nor U2745 (N_2745,In_487,In_2429);
nor U2746 (N_2746,In_2234,In_1832);
or U2747 (N_2747,In_1412,In_149);
or U2748 (N_2748,In_2257,In_1149);
nand U2749 (N_2749,In_1218,In_1507);
xor U2750 (N_2750,In_2469,In_483);
and U2751 (N_2751,In_288,In_154);
or U2752 (N_2752,In_859,In_2307);
or U2753 (N_2753,In_1711,In_510);
nand U2754 (N_2754,In_398,In_983);
and U2755 (N_2755,In_1758,In_1571);
nor U2756 (N_2756,In_1543,In_979);
xnor U2757 (N_2757,In_1184,In_1796);
or U2758 (N_2758,In_1730,In_930);
nor U2759 (N_2759,In_728,In_2053);
xor U2760 (N_2760,In_2135,In_216);
and U2761 (N_2761,In_1173,In_1954);
or U2762 (N_2762,In_903,In_85);
or U2763 (N_2763,In_1581,In_952);
xnor U2764 (N_2764,In_1454,In_1316);
nand U2765 (N_2765,In_2009,In_1480);
nand U2766 (N_2766,In_1003,In_816);
or U2767 (N_2767,In_763,In_952);
xor U2768 (N_2768,In_1538,In_443);
nor U2769 (N_2769,In_522,In_2261);
and U2770 (N_2770,In_984,In_2340);
nand U2771 (N_2771,In_1455,In_1672);
and U2772 (N_2772,In_1465,In_1308);
nand U2773 (N_2773,In_2214,In_4);
nand U2774 (N_2774,In_2257,In_654);
or U2775 (N_2775,In_919,In_78);
nor U2776 (N_2776,In_777,In_302);
or U2777 (N_2777,In_1176,In_1074);
nand U2778 (N_2778,In_892,In_1642);
nor U2779 (N_2779,In_120,In_741);
and U2780 (N_2780,In_1757,In_1374);
or U2781 (N_2781,In_2001,In_1252);
and U2782 (N_2782,In_1196,In_1722);
nand U2783 (N_2783,In_1799,In_2217);
xnor U2784 (N_2784,In_970,In_1408);
xnor U2785 (N_2785,In_447,In_95);
or U2786 (N_2786,In_328,In_2032);
nor U2787 (N_2787,In_2368,In_2274);
nor U2788 (N_2788,In_2007,In_777);
xnor U2789 (N_2789,In_2374,In_2314);
or U2790 (N_2790,In_231,In_1895);
nor U2791 (N_2791,In_1785,In_2272);
nor U2792 (N_2792,In_293,In_1398);
or U2793 (N_2793,In_954,In_97);
nand U2794 (N_2794,In_331,In_2283);
nor U2795 (N_2795,In_1012,In_887);
nor U2796 (N_2796,In_448,In_540);
or U2797 (N_2797,In_2420,In_1517);
nand U2798 (N_2798,In_240,In_1868);
or U2799 (N_2799,In_2471,In_424);
nor U2800 (N_2800,In_1316,In_2340);
xnor U2801 (N_2801,In_752,In_1518);
or U2802 (N_2802,In_550,In_711);
xor U2803 (N_2803,In_2331,In_2167);
nor U2804 (N_2804,In_158,In_585);
or U2805 (N_2805,In_776,In_1452);
nand U2806 (N_2806,In_1851,In_1256);
or U2807 (N_2807,In_1800,In_389);
and U2808 (N_2808,In_1056,In_2384);
nand U2809 (N_2809,In_237,In_458);
xor U2810 (N_2810,In_734,In_1111);
and U2811 (N_2811,In_1114,In_2381);
nand U2812 (N_2812,In_727,In_2421);
nor U2813 (N_2813,In_1800,In_2031);
nand U2814 (N_2814,In_446,In_544);
or U2815 (N_2815,In_744,In_980);
and U2816 (N_2816,In_1913,In_1826);
nand U2817 (N_2817,In_12,In_1896);
and U2818 (N_2818,In_848,In_1120);
and U2819 (N_2819,In_1789,In_983);
xor U2820 (N_2820,In_588,In_586);
and U2821 (N_2821,In_1805,In_64);
or U2822 (N_2822,In_2268,In_2315);
nor U2823 (N_2823,In_1475,In_394);
nand U2824 (N_2824,In_480,In_1403);
and U2825 (N_2825,In_2313,In_1087);
nand U2826 (N_2826,In_2192,In_256);
or U2827 (N_2827,In_1849,In_1712);
xnor U2828 (N_2828,In_1181,In_1429);
or U2829 (N_2829,In_910,In_1020);
and U2830 (N_2830,In_177,In_1432);
or U2831 (N_2831,In_1812,In_921);
xnor U2832 (N_2832,In_573,In_137);
and U2833 (N_2833,In_1580,In_492);
xor U2834 (N_2834,In_635,In_1307);
nand U2835 (N_2835,In_853,In_2053);
or U2836 (N_2836,In_219,In_2188);
nand U2837 (N_2837,In_2393,In_2238);
or U2838 (N_2838,In_616,In_1911);
xor U2839 (N_2839,In_560,In_2384);
nand U2840 (N_2840,In_1318,In_2058);
xnor U2841 (N_2841,In_1874,In_1487);
nand U2842 (N_2842,In_1007,In_1154);
xnor U2843 (N_2843,In_2474,In_1448);
nor U2844 (N_2844,In_2261,In_1029);
xnor U2845 (N_2845,In_1272,In_950);
nand U2846 (N_2846,In_1105,In_386);
and U2847 (N_2847,In_196,In_186);
and U2848 (N_2848,In_792,In_2005);
nand U2849 (N_2849,In_180,In_41);
and U2850 (N_2850,In_2089,In_1577);
nor U2851 (N_2851,In_1150,In_1303);
or U2852 (N_2852,In_2454,In_771);
nor U2853 (N_2853,In_2030,In_904);
nand U2854 (N_2854,In_579,In_668);
and U2855 (N_2855,In_1960,In_152);
xor U2856 (N_2856,In_1259,In_1492);
nor U2857 (N_2857,In_1765,In_2240);
and U2858 (N_2858,In_1130,In_234);
nand U2859 (N_2859,In_1148,In_1354);
xnor U2860 (N_2860,In_996,In_2306);
or U2861 (N_2861,In_901,In_2229);
or U2862 (N_2862,In_29,In_1046);
and U2863 (N_2863,In_2321,In_1433);
xor U2864 (N_2864,In_24,In_1758);
or U2865 (N_2865,In_712,In_170);
or U2866 (N_2866,In_797,In_859);
and U2867 (N_2867,In_1241,In_1590);
xor U2868 (N_2868,In_1016,In_621);
xor U2869 (N_2869,In_1656,In_1763);
or U2870 (N_2870,In_302,In_1593);
nand U2871 (N_2871,In_1419,In_515);
xor U2872 (N_2872,In_1644,In_249);
or U2873 (N_2873,In_697,In_410);
or U2874 (N_2874,In_968,In_2208);
or U2875 (N_2875,In_1533,In_1124);
nor U2876 (N_2876,In_2123,In_1270);
nand U2877 (N_2877,In_2349,In_1212);
nand U2878 (N_2878,In_2131,In_1224);
or U2879 (N_2879,In_1972,In_842);
or U2880 (N_2880,In_769,In_635);
nor U2881 (N_2881,In_2119,In_1550);
xnor U2882 (N_2882,In_2319,In_2224);
xnor U2883 (N_2883,In_40,In_2465);
xor U2884 (N_2884,In_1099,In_698);
nor U2885 (N_2885,In_2229,In_1478);
nand U2886 (N_2886,In_1748,In_1484);
or U2887 (N_2887,In_2366,In_2332);
nor U2888 (N_2888,In_15,In_2011);
nor U2889 (N_2889,In_613,In_1371);
or U2890 (N_2890,In_2381,In_2035);
nand U2891 (N_2891,In_1244,In_1820);
xnor U2892 (N_2892,In_1661,In_1181);
nand U2893 (N_2893,In_1432,In_1282);
xor U2894 (N_2894,In_2471,In_1533);
nand U2895 (N_2895,In_580,In_2190);
nand U2896 (N_2896,In_1413,In_1138);
nand U2897 (N_2897,In_1977,In_1480);
nor U2898 (N_2898,In_1476,In_921);
nand U2899 (N_2899,In_1051,In_2150);
or U2900 (N_2900,In_1273,In_1805);
and U2901 (N_2901,In_979,In_341);
xor U2902 (N_2902,In_47,In_1252);
xor U2903 (N_2903,In_813,In_80);
and U2904 (N_2904,In_1948,In_942);
xnor U2905 (N_2905,In_1465,In_2271);
nor U2906 (N_2906,In_447,In_1378);
or U2907 (N_2907,In_964,In_441);
or U2908 (N_2908,In_2038,In_882);
nor U2909 (N_2909,In_1023,In_2377);
nor U2910 (N_2910,In_436,In_1725);
and U2911 (N_2911,In_1886,In_514);
or U2912 (N_2912,In_1461,In_2304);
nand U2913 (N_2913,In_863,In_2459);
nor U2914 (N_2914,In_1509,In_1155);
nor U2915 (N_2915,In_1234,In_1677);
or U2916 (N_2916,In_1531,In_2287);
xnor U2917 (N_2917,In_2296,In_727);
or U2918 (N_2918,In_1500,In_1203);
xor U2919 (N_2919,In_1912,In_1316);
xnor U2920 (N_2920,In_644,In_739);
nor U2921 (N_2921,In_2197,In_1649);
or U2922 (N_2922,In_779,In_381);
and U2923 (N_2923,In_579,In_2362);
and U2924 (N_2924,In_1641,In_2020);
xor U2925 (N_2925,In_1431,In_501);
nor U2926 (N_2926,In_2315,In_2149);
and U2927 (N_2927,In_369,In_309);
xor U2928 (N_2928,In_2222,In_57);
xnor U2929 (N_2929,In_1956,In_272);
nor U2930 (N_2930,In_1634,In_1318);
nand U2931 (N_2931,In_457,In_785);
nand U2932 (N_2932,In_1884,In_30);
and U2933 (N_2933,In_1596,In_922);
and U2934 (N_2934,In_1654,In_2425);
and U2935 (N_2935,In_2005,In_1639);
and U2936 (N_2936,In_772,In_1206);
xor U2937 (N_2937,In_634,In_1505);
or U2938 (N_2938,In_400,In_1272);
xnor U2939 (N_2939,In_1926,In_1260);
nor U2940 (N_2940,In_864,In_432);
nand U2941 (N_2941,In_1647,In_1017);
nand U2942 (N_2942,In_614,In_1890);
xor U2943 (N_2943,In_1470,In_578);
and U2944 (N_2944,In_893,In_1975);
and U2945 (N_2945,In_269,In_1515);
and U2946 (N_2946,In_1492,In_76);
or U2947 (N_2947,In_1362,In_1101);
xor U2948 (N_2948,In_2033,In_2238);
or U2949 (N_2949,In_781,In_242);
xnor U2950 (N_2950,In_2447,In_86);
and U2951 (N_2951,In_1071,In_267);
xor U2952 (N_2952,In_366,In_243);
nor U2953 (N_2953,In_1699,In_1809);
xor U2954 (N_2954,In_2400,In_1679);
nand U2955 (N_2955,In_932,In_196);
nor U2956 (N_2956,In_1889,In_1347);
or U2957 (N_2957,In_989,In_707);
xnor U2958 (N_2958,In_1495,In_87);
nor U2959 (N_2959,In_1885,In_1705);
nor U2960 (N_2960,In_1661,In_535);
nand U2961 (N_2961,In_1677,In_2406);
or U2962 (N_2962,In_1745,In_958);
xnor U2963 (N_2963,In_2251,In_287);
nor U2964 (N_2964,In_1035,In_2492);
and U2965 (N_2965,In_1094,In_592);
nor U2966 (N_2966,In_2120,In_146);
nand U2967 (N_2967,In_205,In_650);
or U2968 (N_2968,In_2111,In_926);
or U2969 (N_2969,In_1328,In_1351);
xnor U2970 (N_2970,In_1638,In_549);
nand U2971 (N_2971,In_1815,In_2117);
nand U2972 (N_2972,In_339,In_61);
and U2973 (N_2973,In_1680,In_1065);
nor U2974 (N_2974,In_2135,In_743);
xor U2975 (N_2975,In_830,In_1422);
xnor U2976 (N_2976,In_2273,In_1062);
nor U2977 (N_2977,In_45,In_1568);
or U2978 (N_2978,In_2492,In_123);
or U2979 (N_2979,In_54,In_1388);
or U2980 (N_2980,In_1061,In_480);
and U2981 (N_2981,In_1742,In_956);
or U2982 (N_2982,In_60,In_883);
and U2983 (N_2983,In_2090,In_916);
nand U2984 (N_2984,In_2034,In_1226);
nand U2985 (N_2985,In_2158,In_794);
or U2986 (N_2986,In_551,In_2443);
and U2987 (N_2987,In_2385,In_742);
or U2988 (N_2988,In_2110,In_2375);
nor U2989 (N_2989,In_2430,In_1959);
and U2990 (N_2990,In_1689,In_2064);
nand U2991 (N_2991,In_1142,In_1844);
nor U2992 (N_2992,In_1402,In_1030);
and U2993 (N_2993,In_170,In_61);
or U2994 (N_2994,In_1440,In_999);
xnor U2995 (N_2995,In_2060,In_565);
xor U2996 (N_2996,In_357,In_1438);
and U2997 (N_2997,In_2260,In_1071);
xnor U2998 (N_2998,In_1512,In_2449);
nor U2999 (N_2999,In_299,In_185);
and U3000 (N_3000,In_389,In_2303);
or U3001 (N_3001,In_1288,In_16);
or U3002 (N_3002,In_292,In_256);
and U3003 (N_3003,In_436,In_2423);
xnor U3004 (N_3004,In_431,In_2464);
or U3005 (N_3005,In_1367,In_1479);
nor U3006 (N_3006,In_2237,In_2366);
nand U3007 (N_3007,In_300,In_706);
nand U3008 (N_3008,In_659,In_2488);
nor U3009 (N_3009,In_1432,In_619);
nor U3010 (N_3010,In_833,In_1186);
xor U3011 (N_3011,In_249,In_386);
nor U3012 (N_3012,In_1896,In_2161);
or U3013 (N_3013,In_1370,In_926);
xnor U3014 (N_3014,In_383,In_18);
nor U3015 (N_3015,In_645,In_760);
nand U3016 (N_3016,In_1597,In_2083);
xor U3017 (N_3017,In_2496,In_1562);
xnor U3018 (N_3018,In_1885,In_2127);
and U3019 (N_3019,In_1888,In_308);
and U3020 (N_3020,In_1498,In_50);
and U3021 (N_3021,In_1199,In_497);
nand U3022 (N_3022,In_1086,In_237);
xnor U3023 (N_3023,In_2448,In_1826);
nand U3024 (N_3024,In_908,In_1718);
or U3025 (N_3025,In_1651,In_459);
and U3026 (N_3026,In_1637,In_764);
nand U3027 (N_3027,In_2,In_628);
or U3028 (N_3028,In_264,In_623);
and U3029 (N_3029,In_866,In_1773);
and U3030 (N_3030,In_62,In_781);
nor U3031 (N_3031,In_1032,In_1700);
xnor U3032 (N_3032,In_1831,In_971);
nor U3033 (N_3033,In_1163,In_2327);
and U3034 (N_3034,In_1619,In_1228);
and U3035 (N_3035,In_1901,In_2066);
nand U3036 (N_3036,In_460,In_2106);
nor U3037 (N_3037,In_2155,In_868);
or U3038 (N_3038,In_909,In_934);
nor U3039 (N_3039,In_378,In_1100);
or U3040 (N_3040,In_644,In_1890);
nand U3041 (N_3041,In_940,In_2344);
nand U3042 (N_3042,In_1372,In_1729);
and U3043 (N_3043,In_695,In_2141);
xnor U3044 (N_3044,In_1798,In_1940);
nand U3045 (N_3045,In_147,In_1033);
or U3046 (N_3046,In_923,In_734);
nand U3047 (N_3047,In_671,In_2439);
nor U3048 (N_3048,In_131,In_2421);
xnor U3049 (N_3049,In_726,In_2482);
or U3050 (N_3050,In_1419,In_2214);
nor U3051 (N_3051,In_1544,In_814);
nor U3052 (N_3052,In_136,In_990);
and U3053 (N_3053,In_576,In_2135);
nor U3054 (N_3054,In_386,In_1348);
or U3055 (N_3055,In_262,In_1271);
or U3056 (N_3056,In_1393,In_1601);
nor U3057 (N_3057,In_162,In_2114);
or U3058 (N_3058,In_829,In_1212);
nand U3059 (N_3059,In_2024,In_1207);
or U3060 (N_3060,In_994,In_1532);
xnor U3061 (N_3061,In_194,In_591);
xnor U3062 (N_3062,In_2028,In_1071);
xor U3063 (N_3063,In_1969,In_1260);
or U3064 (N_3064,In_896,In_2495);
nand U3065 (N_3065,In_2151,In_2160);
nor U3066 (N_3066,In_2081,In_731);
xor U3067 (N_3067,In_838,In_2368);
and U3068 (N_3068,In_1779,In_746);
nand U3069 (N_3069,In_2004,In_2022);
nor U3070 (N_3070,In_817,In_713);
nor U3071 (N_3071,In_524,In_530);
and U3072 (N_3072,In_975,In_917);
nand U3073 (N_3073,In_2047,In_502);
or U3074 (N_3074,In_530,In_822);
and U3075 (N_3075,In_1829,In_1332);
and U3076 (N_3076,In_688,In_2321);
nand U3077 (N_3077,In_621,In_2208);
or U3078 (N_3078,In_1886,In_1733);
or U3079 (N_3079,In_963,In_1112);
nand U3080 (N_3080,In_1688,In_519);
or U3081 (N_3081,In_1860,In_1564);
or U3082 (N_3082,In_1677,In_1133);
or U3083 (N_3083,In_1500,In_115);
or U3084 (N_3084,In_1849,In_324);
nor U3085 (N_3085,In_183,In_2091);
xor U3086 (N_3086,In_1041,In_2013);
nor U3087 (N_3087,In_2050,In_1378);
nand U3088 (N_3088,In_1416,In_6);
xnor U3089 (N_3089,In_1895,In_2162);
nand U3090 (N_3090,In_229,In_973);
and U3091 (N_3091,In_402,In_1164);
and U3092 (N_3092,In_1985,In_53);
or U3093 (N_3093,In_1263,In_1140);
xor U3094 (N_3094,In_1115,In_207);
nand U3095 (N_3095,In_411,In_1077);
xnor U3096 (N_3096,In_32,In_1744);
or U3097 (N_3097,In_626,In_90);
and U3098 (N_3098,In_123,In_162);
nand U3099 (N_3099,In_653,In_2424);
and U3100 (N_3100,In_1290,In_633);
nor U3101 (N_3101,In_1356,In_1563);
and U3102 (N_3102,In_1107,In_2330);
or U3103 (N_3103,In_703,In_722);
or U3104 (N_3104,In_1790,In_1641);
xnor U3105 (N_3105,In_2157,In_1740);
xor U3106 (N_3106,In_727,In_1138);
xor U3107 (N_3107,In_1994,In_2421);
xnor U3108 (N_3108,In_2036,In_1628);
nor U3109 (N_3109,In_1498,In_174);
and U3110 (N_3110,In_1927,In_1375);
nor U3111 (N_3111,In_2449,In_691);
nand U3112 (N_3112,In_1950,In_2179);
nor U3113 (N_3113,In_1723,In_1896);
nor U3114 (N_3114,In_584,In_943);
nand U3115 (N_3115,In_1417,In_1431);
or U3116 (N_3116,In_540,In_2097);
xor U3117 (N_3117,In_1858,In_2388);
nand U3118 (N_3118,In_806,In_1313);
nor U3119 (N_3119,In_766,In_1807);
xor U3120 (N_3120,In_1806,In_2424);
and U3121 (N_3121,In_2226,In_1180);
xnor U3122 (N_3122,In_242,In_1295);
xnor U3123 (N_3123,In_2340,In_5);
and U3124 (N_3124,In_1649,In_385);
or U3125 (N_3125,N_2283,N_2666);
and U3126 (N_3126,N_1275,N_1669);
or U3127 (N_3127,N_2346,N_286);
nand U3128 (N_3128,N_2811,N_1362);
nor U3129 (N_3129,N_2113,N_1714);
xnor U3130 (N_3130,N_2493,N_192);
xor U3131 (N_3131,N_721,N_1179);
xnor U3132 (N_3132,N_2287,N_167);
nand U3133 (N_3133,N_512,N_1839);
nand U3134 (N_3134,N_20,N_688);
and U3135 (N_3135,N_1074,N_1671);
nand U3136 (N_3136,N_733,N_2567);
and U3137 (N_3137,N_2463,N_862);
xor U3138 (N_3138,N_366,N_827);
or U3139 (N_3139,N_703,N_2832);
xnor U3140 (N_3140,N_1633,N_121);
or U3141 (N_3141,N_2830,N_2216);
xor U3142 (N_3142,N_3015,N_1116);
nand U3143 (N_3143,N_147,N_2397);
nand U3144 (N_3144,N_763,N_2232);
nor U3145 (N_3145,N_842,N_2071);
or U3146 (N_3146,N_1568,N_2664);
nand U3147 (N_3147,N_527,N_1399);
nand U3148 (N_3148,N_406,N_2987);
and U3149 (N_3149,N_2098,N_1016);
or U3150 (N_3150,N_1637,N_1348);
and U3151 (N_3151,N_71,N_1073);
nor U3152 (N_3152,N_964,N_1648);
and U3153 (N_3153,N_2030,N_3011);
nand U3154 (N_3154,N_2360,N_2227);
or U3155 (N_3155,N_4,N_2824);
or U3156 (N_3156,N_1639,N_1578);
or U3157 (N_3157,N_1543,N_2236);
or U3158 (N_3158,N_1619,N_706);
nand U3159 (N_3159,N_2288,N_2056);
nand U3160 (N_3160,N_2398,N_2197);
and U3161 (N_3161,N_1207,N_2210);
xor U3162 (N_3162,N_1065,N_3097);
nor U3163 (N_3163,N_2436,N_1511);
or U3164 (N_3164,N_2701,N_1412);
nor U3165 (N_3165,N_2069,N_2779);
and U3166 (N_3166,N_438,N_2912);
nor U3167 (N_3167,N_3021,N_3085);
nor U3168 (N_3168,N_2704,N_2728);
nor U3169 (N_3169,N_321,N_1503);
nor U3170 (N_3170,N_1397,N_689);
nand U3171 (N_3171,N_1475,N_793);
nand U3172 (N_3172,N_1172,N_1313);
nor U3173 (N_3173,N_160,N_1898);
and U3174 (N_3174,N_3067,N_93);
xnor U3175 (N_3175,N_1486,N_2184);
or U3176 (N_3176,N_3107,N_2383);
nor U3177 (N_3177,N_2776,N_1783);
and U3178 (N_3178,N_193,N_2538);
and U3179 (N_3179,N_1319,N_87);
and U3180 (N_3180,N_1444,N_77);
or U3181 (N_3181,N_2928,N_2042);
nand U3182 (N_3182,N_1332,N_2315);
xor U3183 (N_3183,N_2583,N_2437);
or U3184 (N_3184,N_1934,N_1258);
and U3185 (N_3185,N_2768,N_630);
or U3186 (N_3186,N_351,N_2057);
nand U3187 (N_3187,N_2087,N_2316);
nor U3188 (N_3188,N_2485,N_1973);
and U3189 (N_3189,N_3003,N_2376);
nand U3190 (N_3190,N_1952,N_694);
or U3191 (N_3191,N_2963,N_1247);
nand U3192 (N_3192,N_938,N_549);
nor U3193 (N_3193,N_681,N_1910);
nor U3194 (N_3194,N_2469,N_38);
or U3195 (N_3195,N_801,N_1560);
and U3196 (N_3196,N_385,N_1478);
and U3197 (N_3197,N_2791,N_2708);
nor U3198 (N_3198,N_2818,N_26);
xor U3199 (N_3199,N_1244,N_104);
nor U3200 (N_3200,N_568,N_2931);
nand U3201 (N_3201,N_687,N_80);
nand U3202 (N_3202,N_2771,N_854);
and U3203 (N_3203,N_381,N_1050);
and U3204 (N_3204,N_1420,N_2082);
and U3205 (N_3205,N_62,N_2500);
xnor U3206 (N_3206,N_2626,N_3084);
xor U3207 (N_3207,N_948,N_914);
xnor U3208 (N_3208,N_1526,N_51);
xor U3209 (N_3209,N_922,N_1308);
and U3210 (N_3210,N_1328,N_1810);
nor U3211 (N_3211,N_2909,N_2792);
xor U3212 (N_3212,N_504,N_560);
nand U3213 (N_3213,N_2599,N_1510);
nand U3214 (N_3214,N_184,N_2003);
nand U3215 (N_3215,N_1438,N_3010);
nand U3216 (N_3216,N_3047,N_430);
nor U3217 (N_3217,N_1583,N_954);
or U3218 (N_3218,N_2377,N_777);
or U3219 (N_3219,N_389,N_2093);
nor U3220 (N_3220,N_672,N_2486);
or U3221 (N_3221,N_136,N_979);
or U3222 (N_3222,N_875,N_205);
or U3223 (N_3223,N_408,N_2359);
and U3224 (N_3224,N_1216,N_2411);
xor U3225 (N_3225,N_1201,N_985);
nor U3226 (N_3226,N_8,N_1142);
nor U3227 (N_3227,N_1445,N_2100);
and U3228 (N_3228,N_2644,N_2009);
nor U3229 (N_3229,N_1271,N_856);
or U3230 (N_3230,N_370,N_25);
nor U3231 (N_3231,N_2781,N_2074);
or U3232 (N_3232,N_828,N_781);
or U3233 (N_3233,N_2324,N_316);
xor U3234 (N_3234,N_1889,N_3022);
and U3235 (N_3235,N_989,N_1311);
nand U3236 (N_3236,N_2535,N_3034);
xor U3237 (N_3237,N_2340,N_186);
and U3238 (N_3238,N_2494,N_1873);
xor U3239 (N_3239,N_131,N_1352);
nor U3240 (N_3240,N_1989,N_181);
and U3241 (N_3241,N_1390,N_2660);
and U3242 (N_3242,N_287,N_332);
nor U3243 (N_3243,N_1573,N_520);
or U3244 (N_3244,N_2410,N_259);
and U3245 (N_3245,N_343,N_1758);
or U3246 (N_3246,N_1559,N_900);
or U3247 (N_3247,N_678,N_2630);
and U3248 (N_3248,N_276,N_1139);
nand U3249 (N_3249,N_731,N_753);
or U3250 (N_3250,N_1092,N_2778);
xnor U3251 (N_3251,N_1620,N_2145);
nand U3252 (N_3252,N_2477,N_2204);
xnor U3253 (N_3253,N_227,N_2264);
nand U3254 (N_3254,N_570,N_1488);
and U3255 (N_3255,N_1832,N_2503);
xnor U3256 (N_3256,N_418,N_2610);
and U3257 (N_3257,N_3076,N_1256);
xor U3258 (N_3258,N_3091,N_2980);
nor U3259 (N_3259,N_249,N_2180);
nand U3260 (N_3260,N_1598,N_1572);
or U3261 (N_3261,N_398,N_2070);
nor U3262 (N_3262,N_1751,N_3102);
nand U3263 (N_3263,N_1931,N_2426);
or U3264 (N_3264,N_274,N_1415);
nand U3265 (N_3265,N_546,N_596);
or U3266 (N_3266,N_890,N_1705);
and U3267 (N_3267,N_2171,N_10);
nor U3268 (N_3268,N_3096,N_2347);
or U3269 (N_3269,N_340,N_2140);
xor U3270 (N_3270,N_617,N_2829);
or U3271 (N_3271,N_2616,N_1351);
and U3272 (N_3272,N_283,N_2044);
nand U3273 (N_3273,N_1457,N_830);
nand U3274 (N_3274,N_2531,N_1377);
nor U3275 (N_3275,N_544,N_1630);
xnor U3276 (N_3276,N_2689,N_1966);
nor U3277 (N_3277,N_2373,N_1701);
or U3278 (N_3278,N_727,N_870);
nor U3279 (N_3279,N_1281,N_1782);
nand U3280 (N_3280,N_909,N_1997);
nor U3281 (N_3281,N_1237,N_2352);
or U3282 (N_3282,N_2192,N_867);
nand U3283 (N_3283,N_2220,N_1760);
or U3284 (N_3284,N_1697,N_2577);
and U3285 (N_3285,N_2101,N_991);
nand U3286 (N_3286,N_2586,N_707);
or U3287 (N_3287,N_2266,N_2391);
nor U3288 (N_3288,N_2941,N_978);
nor U3289 (N_3289,N_743,N_2008);
and U3290 (N_3290,N_409,N_3012);
or U3291 (N_3291,N_2260,N_1833);
nor U3292 (N_3292,N_3090,N_2984);
nor U3293 (N_3293,N_2631,N_1191);
nor U3294 (N_3294,N_3002,N_869);
or U3295 (N_3295,N_1431,N_1106);
xor U3296 (N_3296,N_224,N_2520);
xor U3297 (N_3297,N_3033,N_602);
nor U3298 (N_3298,N_493,N_159);
xnor U3299 (N_3299,N_3078,N_2050);
or U3300 (N_3300,N_2143,N_1450);
nor U3301 (N_3301,N_2951,N_3109);
and U3302 (N_3302,N_3074,N_2303);
xnor U3303 (N_3303,N_1978,N_122);
nand U3304 (N_3304,N_1436,N_1233);
nand U3305 (N_3305,N_756,N_605);
or U3306 (N_3306,N_814,N_1880);
nor U3307 (N_3307,N_3122,N_1871);
and U3308 (N_3308,N_105,N_986);
nand U3309 (N_3309,N_1921,N_1946);
xnor U3310 (N_3310,N_2942,N_1707);
nand U3311 (N_3311,N_2453,N_2096);
or U3312 (N_3312,N_637,N_1658);
and U3313 (N_3313,N_2461,N_2713);
or U3314 (N_3314,N_950,N_2843);
nand U3315 (N_3315,N_156,N_3001);
xnor U3316 (N_3316,N_174,N_3110);
nand U3317 (N_3317,N_2130,N_1563);
and U3318 (N_3318,N_2823,N_2851);
nor U3319 (N_3319,N_2627,N_658);
and U3320 (N_3320,N_2684,N_1939);
and U3321 (N_3321,N_2466,N_2000);
and U3322 (N_3322,N_2696,N_2226);
or U3323 (N_3323,N_894,N_1688);
and U3324 (N_3324,N_3028,N_2891);
xnor U3325 (N_3325,N_2517,N_2409);
xnor U3326 (N_3326,N_916,N_2723);
nor U3327 (N_3327,N_117,N_3104);
and U3328 (N_3328,N_1158,N_2923);
nor U3329 (N_3329,N_754,N_2425);
xnor U3330 (N_3330,N_2556,N_171);
xor U3331 (N_3331,N_214,N_1122);
nand U3332 (N_3332,N_1301,N_507);
nor U3333 (N_3333,N_2849,N_1534);
or U3334 (N_3334,N_2010,N_2046);
nand U3335 (N_3335,N_3040,N_1015);
nor U3336 (N_3336,N_1059,N_2196);
nand U3337 (N_3337,N_2319,N_168);
or U3338 (N_3338,N_1204,N_2566);
or U3339 (N_3339,N_1235,N_593);
and U3340 (N_3340,N_3008,N_755);
nand U3341 (N_3341,N_1603,N_1675);
nor U3342 (N_3342,N_1339,N_1212);
xor U3343 (N_3343,N_2183,N_857);
nand U3344 (N_3344,N_1435,N_317);
and U3345 (N_3345,N_639,N_2747);
and U3346 (N_3346,N_2919,N_2972);
nor U3347 (N_3347,N_1899,N_2798);
and U3348 (N_3348,N_1144,N_1005);
xnor U3349 (N_3349,N_1003,N_2362);
nor U3350 (N_3350,N_1780,N_268);
and U3351 (N_3351,N_550,N_1029);
xor U3352 (N_3352,N_597,N_2430);
or U3353 (N_3353,N_1721,N_107);
xor U3354 (N_3354,N_1298,N_846);
xnor U3355 (N_3355,N_50,N_2602);
nand U3356 (N_3356,N_2393,N_1395);
and U3357 (N_3357,N_1115,N_2270);
or U3358 (N_3358,N_1335,N_1490);
or U3359 (N_3359,N_2814,N_348);
and U3360 (N_3360,N_2205,N_1803);
or U3361 (N_3361,N_988,N_803);
xor U3362 (N_3362,N_2203,N_1944);
xnor U3363 (N_3363,N_2557,N_2403);
nor U3364 (N_3364,N_2526,N_2793);
nand U3365 (N_3365,N_671,N_661);
and U3366 (N_3366,N_838,N_2725);
and U3367 (N_3367,N_1464,N_809);
xor U3368 (N_3368,N_936,N_543);
nand U3369 (N_3369,N_3006,N_494);
xor U3370 (N_3370,N_565,N_1553);
nand U3371 (N_3371,N_812,N_1433);
xor U3372 (N_3372,N_864,N_280);
and U3373 (N_3373,N_2257,N_1755);
nor U3374 (N_3374,N_1804,N_85);
nand U3375 (N_3375,N_2129,N_464);
or U3376 (N_3376,N_2871,N_1355);
nand U3377 (N_3377,N_217,N_1268);
xnor U3378 (N_3378,N_3086,N_319);
and U3379 (N_3379,N_1866,N_164);
nor U3380 (N_3380,N_613,N_2939);
or U3381 (N_3381,N_514,N_1641);
and U3382 (N_3382,N_1717,N_1481);
nand U3383 (N_3383,N_2935,N_715);
or U3384 (N_3384,N_903,N_2570);
nor U3385 (N_3385,N_1571,N_2253);
or U3386 (N_3386,N_1911,N_212);
nand U3387 (N_3387,N_2005,N_1402);
nor U3388 (N_3388,N_2677,N_2958);
xor U3389 (N_3389,N_2518,N_1590);
nand U3390 (N_3390,N_307,N_3114);
or U3391 (N_3391,N_1231,N_1292);
nor U3392 (N_3392,N_804,N_1032);
and U3393 (N_3393,N_54,N_2353);
and U3394 (N_3394,N_1887,N_1725);
xnor U3395 (N_3395,N_2142,N_879);
nor U3396 (N_3396,N_1213,N_2608);
or U3397 (N_3397,N_2863,N_253);
nor U3398 (N_3398,N_2846,N_1632);
nand U3399 (N_3399,N_2640,N_1859);
and U3400 (N_3400,N_187,N_1738);
and U3401 (N_3401,N_1733,N_1229);
and U3402 (N_3402,N_1089,N_2614);
nand U3403 (N_3403,N_3088,N_505);
nor U3404 (N_3404,N_373,N_1564);
nand U3405 (N_3405,N_1561,N_1223);
xor U3406 (N_3406,N_2431,N_897);
nor U3407 (N_3407,N_1737,N_2777);
nand U3408 (N_3408,N_1709,N_225);
nor U3409 (N_3409,N_1774,N_2451);
nand U3410 (N_3410,N_347,N_1631);
nand U3411 (N_3411,N_2548,N_1263);
and U3412 (N_3412,N_545,N_200);
nand U3413 (N_3413,N_2222,N_334);
or U3414 (N_3414,N_825,N_518);
or U3415 (N_3415,N_1358,N_1702);
xnor U3416 (N_3416,N_2527,N_2473);
nand U3417 (N_3417,N_1775,N_482);
or U3418 (N_3418,N_810,N_2209);
xor U3419 (N_3419,N_270,N_2712);
or U3420 (N_3420,N_1090,N_2529);
nor U3421 (N_3421,N_502,N_1055);
nor U3422 (N_3422,N_152,N_2173);
xnor U3423 (N_3423,N_2982,N_2867);
and U3424 (N_3424,N_1326,N_2737);
or U3425 (N_3425,N_263,N_1638);
or U3426 (N_3426,N_623,N_439);
and U3427 (N_3427,N_1754,N_1398);
nand U3428 (N_3428,N_431,N_1967);
or U3429 (N_3429,N_1980,N_650);
nor U3430 (N_3430,N_2158,N_1801);
or U3431 (N_3431,N_1267,N_260);
nor U3432 (N_3432,N_1024,N_760);
nand U3433 (N_3433,N_3036,N_1596);
and U3434 (N_3434,N_2131,N_2174);
nand U3435 (N_3435,N_2041,N_1240);
nand U3436 (N_3436,N_3106,N_1891);
or U3437 (N_3437,N_1888,N_1894);
nor U3438 (N_3438,N_2094,N_2642);
xor U3439 (N_3439,N_1706,N_76);
xor U3440 (N_3440,N_1035,N_81);
or U3441 (N_3441,N_1805,N_330);
and U3442 (N_3442,N_2903,N_443);
nor U3443 (N_3443,N_1236,N_1072);
and U3444 (N_3444,N_169,N_742);
or U3445 (N_3445,N_1276,N_1466);
or U3446 (N_3446,N_1941,N_665);
xor U3447 (N_3447,N_2746,N_957);
nor U3448 (N_3448,N_920,N_1574);
xor U3449 (N_3449,N_2399,N_886);
xnor U3450 (N_3450,N_3058,N_2679);
xor U3451 (N_3451,N_1716,N_877);
or U3452 (N_3452,N_1672,N_2820);
nor U3453 (N_3453,N_2047,N_2123);
or U3454 (N_3454,N_1196,N_2955);
nand U3455 (N_3455,N_3068,N_693);
xnor U3456 (N_3456,N_874,N_344);
nand U3457 (N_3457,N_974,N_1011);
and U3458 (N_3458,N_2167,N_816);
and U3459 (N_3459,N_2657,N_1948);
or U3460 (N_3460,N_2974,N_1699);
nand U3461 (N_3461,N_1876,N_2134);
or U3462 (N_3462,N_525,N_1926);
nor U3463 (N_3463,N_2394,N_2124);
nor U3464 (N_3464,N_2943,N_2036);
or U3465 (N_3465,N_2692,N_2975);
or U3466 (N_3466,N_2693,N_1130);
or U3467 (N_3467,N_2541,N_972);
xnor U3468 (N_3468,N_3079,N_2992);
nand U3469 (N_3469,N_1777,N_2565);
xor U3470 (N_3470,N_752,N_341);
and U3471 (N_3471,N_2784,N_1977);
nand U3472 (N_3472,N_1455,N_2540);
or U3473 (N_3473,N_1593,N_2351);
and U3474 (N_3474,N_364,N_194);
nor U3475 (N_3475,N_849,N_2248);
or U3476 (N_3476,N_60,N_151);
and U3477 (N_3477,N_1101,N_281);
nand U3478 (N_3478,N_822,N_626);
nor U3479 (N_3479,N_2545,N_1291);
nand U3480 (N_3480,N_1517,N_1499);
nor U3481 (N_3481,N_2193,N_2294);
and U3482 (N_3482,N_2081,N_2363);
xor U3483 (N_3483,N_1537,N_2827);
or U3484 (N_3484,N_2555,N_509);
nand U3485 (N_3485,N_454,N_1834);
and U3486 (N_3486,N_2967,N_496);
and U3487 (N_3487,N_2886,N_1047);
or U3488 (N_3488,N_3089,N_2029);
or U3489 (N_3489,N_817,N_2813);
nand U3490 (N_3490,N_1163,N_1576);
or U3491 (N_3491,N_1219,N_573);
nor U3492 (N_3492,N_1245,N_918);
nor U3493 (N_3493,N_1660,N_2787);
nand U3494 (N_3494,N_587,N_2097);
and U3495 (N_3495,N_1947,N_946);
or U3496 (N_3496,N_436,N_163);
and U3497 (N_3497,N_2854,N_1286);
or U3498 (N_3498,N_65,N_1359);
nor U3499 (N_3499,N_2900,N_1719);
or U3500 (N_3500,N_1950,N_984);
nor U3501 (N_3501,N_1821,N_649);
xor U3502 (N_3502,N_23,N_1868);
and U3503 (N_3503,N_161,N_999);
and U3504 (N_3504,N_1062,N_1806);
nand U3505 (N_3505,N_851,N_1329);
or U3506 (N_3506,N_487,N_295);
or U3507 (N_3507,N_2960,N_2905);
and U3508 (N_3508,N_480,N_52);
nand U3509 (N_3509,N_1396,N_1018);
xnor U3510 (N_3510,N_2976,N_1831);
and U3511 (N_3511,N_1369,N_3101);
nand U3512 (N_3512,N_3044,N_2803);
and U3513 (N_3513,N_2705,N_254);
or U3514 (N_3514,N_1604,N_981);
nor U3515 (N_3515,N_2,N_1673);
xor U3516 (N_3516,N_177,N_2001);
and U3517 (N_3517,N_483,N_1850);
nor U3518 (N_3518,N_711,N_1260);
xnor U3519 (N_3519,N_1976,N_844);
or U3520 (N_3520,N_1188,N_273);
and U3521 (N_3521,N_241,N_638);
nand U3522 (N_3522,N_1651,N_1079);
xor U3523 (N_3523,N_2831,N_1808);
and U3524 (N_3524,N_2511,N_435);
nor U3525 (N_3525,N_998,N_1470);
xor U3526 (N_3526,N_2293,N_1279);
nor U3527 (N_3527,N_2277,N_2388);
nor U3528 (N_3528,N_2132,N_2265);
and U3529 (N_3529,N_1509,N_2498);
nand U3530 (N_3530,N_2501,N_1487);
and U3531 (N_3531,N_2629,N_138);
nand U3532 (N_3532,N_2625,N_1676);
nand U3533 (N_3533,N_1974,N_2439);
and U3534 (N_3534,N_896,N_2429);
and U3535 (N_3535,N_1538,N_1273);
nand U3536 (N_3536,N_614,N_2215);
and U3537 (N_3537,N_2990,N_1371);
or U3538 (N_3538,N_667,N_2613);
nor U3539 (N_3539,N_262,N_2638);
nor U3540 (N_3540,N_718,N_675);
and U3541 (N_3541,N_1012,N_19);
nand U3542 (N_3542,N_537,N_495);
nor U3543 (N_3543,N_377,N_2414);
or U3544 (N_3544,N_1798,N_577);
xor U3545 (N_3545,N_2957,N_2729);
xor U3546 (N_3546,N_2547,N_668);
nand U3547 (N_3547,N_1192,N_240);
xor U3548 (N_3548,N_2994,N_2048);
and U3549 (N_3549,N_2135,N_3071);
xnor U3550 (N_3550,N_243,N_2482);
nor U3551 (N_3551,N_172,N_2594);
nand U3552 (N_3552,N_1811,N_2387);
nor U3553 (N_3553,N_2648,N_2218);
or U3554 (N_3554,N_692,N_2187);
nand U3555 (N_3555,N_1463,N_2874);
or U3556 (N_3556,N_1284,N_2952);
nor U3557 (N_3557,N_2106,N_2032);
nand U3558 (N_3558,N_726,N_404);
xnor U3559 (N_3559,N_2420,N_769);
nand U3560 (N_3560,N_350,N_572);
xnor U3561 (N_3561,N_2489,N_1141);
or U3562 (N_3562,N_314,N_445);
nor U3563 (N_3563,N_2111,N_1556);
nor U3564 (N_3564,N_1346,N_446);
nor U3565 (N_3565,N_2786,N_934);
and U3566 (N_3566,N_2744,N_532);
nand U3567 (N_3567,N_1713,N_2736);
nand U3568 (N_3568,N_79,N_137);
and U3569 (N_3569,N_229,N_589);
or U3570 (N_3570,N_1041,N_1209);
or U3571 (N_3571,N_403,N_2006);
xor U3572 (N_3572,N_651,N_2754);
or U3573 (N_3573,N_2060,N_2881);
nor U3574 (N_3574,N_1925,N_500);
or U3575 (N_3575,N_2457,N_1796);
or U3576 (N_3576,N_795,N_746);
nor U3577 (N_3577,N_624,N_2372);
nor U3578 (N_3578,N_3105,N_218);
nand U3579 (N_3579,N_2929,N_2890);
xor U3580 (N_3580,N_1127,N_1456);
nand U3581 (N_3581,N_1070,N_557);
and U3582 (N_3582,N_2685,N_1150);
or U3583 (N_3583,N_1935,N_3094);
xor U3584 (N_3584,N_1968,N_852);
nand U3585 (N_3585,N_2973,N_963);
nor U3586 (N_3586,N_1442,N_1228);
xor U3587 (N_3587,N_819,N_547);
or U3588 (N_3588,N_1290,N_656);
or U3589 (N_3589,N_2983,N_2138);
and U3590 (N_3590,N_386,N_1856);
xor U3591 (N_3591,N_2932,N_2231);
and U3592 (N_3592,N_18,N_2572);
and U3593 (N_3593,N_2505,N_2936);
xnor U3594 (N_3594,N_292,N_949);
nor U3595 (N_3595,N_1984,N_2937);
xnor U3596 (N_3596,N_2026,N_2213);
and U3597 (N_3597,N_3123,N_1994);
and U3598 (N_3598,N_583,N_1093);
nand U3599 (N_3599,N_2024,N_53);
nand U3600 (N_3600,N_5,N_329);
or U3601 (N_3601,N_2152,N_3017);
and U3602 (N_3602,N_1120,N_3075);
nand U3603 (N_3603,N_1535,N_1274);
and U3604 (N_3604,N_1121,N_2714);
nand U3605 (N_3605,N_673,N_889);
nand U3606 (N_3606,N_1333,N_2949);
or U3607 (N_3607,N_1447,N_808);
nor U3608 (N_3608,N_2358,N_2571);
nor U3609 (N_3609,N_1813,N_1541);
or U3610 (N_3610,N_1265,N_100);
and U3611 (N_3611,N_2875,N_2504);
xor U3612 (N_3612,N_1527,N_1722);
nor U3613 (N_3613,N_1756,N_1847);
and U3614 (N_3614,N_664,N_170);
and U3615 (N_3615,N_798,N_1861);
xnor U3616 (N_3616,N_1105,N_2079);
xor U3617 (N_3617,N_539,N_1140);
nor U3618 (N_3618,N_2267,N_33);
nand U3619 (N_3619,N_772,N_997);
xnor U3620 (N_3620,N_1913,N_298);
nor U3621 (N_3621,N_1642,N_43);
and U3622 (N_3622,N_2752,N_695);
nand U3623 (N_3623,N_1595,N_2945);
xnor U3624 (N_3624,N_1242,N_1908);
xor U3625 (N_3625,N_1965,N_2918);
xnor U3626 (N_3626,N_388,N_2336);
and U3627 (N_3627,N_1682,N_1173);
xor U3628 (N_3628,N_935,N_1909);
nor U3629 (N_3629,N_908,N_2534);
and U3630 (N_3630,N_2745,N_2406);
xnor U3631 (N_3631,N_3045,N_1460);
or U3632 (N_3632,N_2624,N_396);
nand U3633 (N_3633,N_375,N_2427);
nor U3634 (N_3634,N_1567,N_1109);
xor U3635 (N_3635,N_1277,N_326);
nor U3636 (N_3636,N_222,N_9);
or U3637 (N_3637,N_1698,N_1076);
or U3638 (N_3638,N_148,N_2715);
and U3639 (N_3639,N_2062,N_476);
and U3640 (N_3640,N_1496,N_1695);
and U3641 (N_3641,N_1958,N_1215);
and U3642 (N_3642,N_1477,N_2665);
or U3643 (N_3643,N_2603,N_2561);
or U3644 (N_3644,N_2760,N_2102);
or U3645 (N_3645,N_663,N_1498);
nand U3646 (N_3646,N_625,N_2646);
or U3647 (N_3647,N_2782,N_2458);
nor U3648 (N_3648,N_1042,N_1224);
or U3649 (N_3649,N_2576,N_3098);
nand U3650 (N_3650,N_2883,N_2168);
xnor U3651 (N_3651,N_2718,N_1791);
or U3652 (N_3652,N_427,N_548);
nand U3653 (N_3653,N_2528,N_2698);
nor U3654 (N_3654,N_1610,N_2780);
xor U3655 (N_3655,N_3054,N_1221);
and U3656 (N_3656,N_248,N_2761);
nor U3657 (N_3657,N_1975,N_21);
or U3658 (N_3658,N_2332,N_685);
or U3659 (N_3659,N_2611,N_322);
and U3660 (N_3660,N_2585,N_729);
or U3661 (N_3661,N_1452,N_1837);
or U3662 (N_3662,N_1581,N_2924);
or U3663 (N_3663,N_2165,N_2107);
or U3664 (N_3664,N_961,N_739);
and U3665 (N_3665,N_2964,N_670);
or U3666 (N_3666,N_1685,N_925);
xor U3667 (N_3667,N_716,N_1829);
or U3668 (N_3668,N_578,N_1184);
nand U3669 (N_3669,N_1776,N_1300);
nor U3670 (N_3670,N_2066,N_858);
xnor U3671 (N_3671,N_264,N_2136);
nor U3672 (N_3672,N_1828,N_1732);
or U3673 (N_3673,N_1649,N_2930);
nor U3674 (N_3674,N_1374,N_2968);
nor U3675 (N_3675,N_2112,N_2118);
nand U3676 (N_3676,N_1960,N_2166);
nor U3677 (N_3677,N_2769,N_284);
and U3678 (N_3678,N_1315,N_919);
and U3679 (N_3679,N_648,N_1491);
and U3680 (N_3680,N_643,N_556);
or U3681 (N_3681,N_473,N_271);
or U3682 (N_3682,N_1647,N_2396);
nand U3683 (N_3683,N_2464,N_95);
and U3684 (N_3684,N_2099,N_2822);
or U3685 (N_3685,N_2126,N_128);
or U3686 (N_3686,N_2177,N_799);
xnor U3687 (N_3687,N_839,N_677);
and U3688 (N_3688,N_1425,N_3103);
xnor U3689 (N_3689,N_1683,N_2054);
nand U3690 (N_3690,N_1835,N_1205);
xor U3691 (N_3691,N_2933,N_1111);
xnor U3692 (N_3692,N_1746,N_616);
nand U3693 (N_3693,N_309,N_2395);
nor U3694 (N_3694,N_2889,N_1174);
or U3695 (N_3695,N_3093,N_1680);
nand U3696 (N_3696,N_258,N_866);
or U3697 (N_3697,N_92,N_554);
or U3698 (N_3698,N_365,N_3020);
nor U3699 (N_3699,N_2741,N_165);
xnor U3700 (N_3700,N_982,N_1885);
nand U3701 (N_3701,N_1124,N_2038);
or U3702 (N_3702,N_1112,N_3112);
or U3703 (N_3703,N_1670,N_444);
nor U3704 (N_3704,N_2908,N_182);
nor U3705 (N_3705,N_2022,N_3059);
nor U3706 (N_3706,N_829,N_1148);
or U3707 (N_3707,N_2225,N_118);
nand U3708 (N_3708,N_876,N_2125);
xnor U3709 (N_3709,N_868,N_2826);
nand U3710 (N_3710,N_1336,N_1366);
or U3711 (N_3711,N_2276,N_202);
nand U3712 (N_3712,N_94,N_2299);
nand U3713 (N_3713,N_3087,N_3080);
nor U3714 (N_3714,N_789,N_2766);
nor U3715 (N_3715,N_2053,N_1650);
nor U3716 (N_3716,N_2224,N_407);
and U3717 (N_3717,N_2250,N_2151);
and U3718 (N_3718,N_1364,N_2775);
nand U3719 (N_3719,N_530,N_2615);
nand U3720 (N_3720,N_618,N_367);
or U3721 (N_3721,N_1513,N_645);
or U3722 (N_3722,N_1986,N_1605);
xor U3723 (N_3723,N_2510,N_1378);
and U3724 (N_3724,N_74,N_336);
or U3725 (N_3725,N_536,N_1167);
nor U3726 (N_3726,N_551,N_3081);
and U3727 (N_3727,N_1061,N_1820);
nand U3728 (N_3728,N_2072,N_747);
and U3729 (N_3729,N_2885,N_1118);
nor U3730 (N_3730,N_2211,N_1694);
or U3731 (N_3731,N_1762,N_1817);
nor U3732 (N_3732,N_153,N_2483);
or U3733 (N_3733,N_2650,N_3055);
nand U3734 (N_3734,N_2734,N_2163);
nor U3735 (N_3735,N_1489,N_1867);
nor U3736 (N_3736,N_1519,N_740);
xnor U3737 (N_3737,N_2433,N_2590);
or U3738 (N_3738,N_1819,N_2921);
nand U3739 (N_3739,N_2088,N_40);
nor U3740 (N_3740,N_3121,N_1031);
nor U3741 (N_3741,N_1907,N_179);
or U3742 (N_3742,N_1334,N_1533);
or U3743 (N_3743,N_2806,N_22);
nor U3744 (N_3744,N_1004,N_2658);
and U3745 (N_3745,N_1906,N_1068);
nor U3746 (N_3746,N_2195,N_1446);
or U3747 (N_3747,N_1690,N_2687);
and U3748 (N_3748,N_11,N_102);
and U3749 (N_3749,N_951,N_228);
xor U3750 (N_3750,N_2953,N_1394);
nor U3751 (N_3751,N_2068,N_3046);
nor U3752 (N_3752,N_859,N_125);
nand U3753 (N_3753,N_973,N_178);
nor U3754 (N_3754,N_2179,N_1849);
nor U3755 (N_3755,N_993,N_368);
xor U3756 (N_3756,N_1045,N_682);
or U3757 (N_3757,N_2750,N_969);
or U3758 (N_3758,N_1953,N_2837);
nand U3759 (N_3759,N_208,N_2285);
nor U3760 (N_3760,N_1959,N_2799);
nand U3761 (N_3761,N_2756,N_2200);
or U3762 (N_3762,N_511,N_2855);
xnor U3763 (N_3763,N_1350,N_2893);
nand U3764 (N_3764,N_2311,N_1440);
nor U3765 (N_3765,N_2966,N_1858);
and U3766 (N_3766,N_1063,N_1646);
or U3767 (N_3767,N_1383,N_751);
or U3768 (N_3768,N_2977,N_1904);
xnor U3769 (N_3769,N_1057,N_929);
nor U3770 (N_3770,N_244,N_579);
xnor U3771 (N_3771,N_2350,N_2021);
nor U3772 (N_3772,N_256,N_1022);
nand U3773 (N_3773,N_109,N_1927);
nor U3774 (N_3774,N_1154,N_451);
nor U3775 (N_3775,N_1961,N_741);
and U3776 (N_3776,N_598,N_2917);
nor U3777 (N_3777,N_1998,N_2812);
xnor U3778 (N_3778,N_1919,N_272);
and U3779 (N_3779,N_2019,N_1627);
and U3780 (N_3780,N_1465,N_3060);
and U3781 (N_3781,N_485,N_1294);
nand U3782 (N_3782,N_2765,N_108);
nor U3783 (N_3783,N_1303,N_528);
nor U3784 (N_3784,N_1614,N_246);
nand U3785 (N_3785,N_2310,N_2895);
or U3786 (N_3786,N_3099,N_1153);
nor U3787 (N_3787,N_2341,N_124);
or U3788 (N_3788,N_2845,N_2127);
nand U3789 (N_3789,N_1807,N_303);
or U3790 (N_3790,N_1500,N_1544);
nor U3791 (N_3791,N_745,N_1266);
nand U3792 (N_3792,N_2051,N_173);
and U3793 (N_3793,N_1608,N_1686);
or U3794 (N_3794,N_2002,N_379);
nand U3795 (N_3795,N_765,N_2465);
nor U3796 (N_3796,N_1429,N_355);
or U3797 (N_3797,N_2580,N_2105);
xor U3798 (N_3798,N_1097,N_2927);
and U3799 (N_3799,N_2554,N_2011);
and U3800 (N_3800,N_2156,N_1038);
nor U3801 (N_3801,N_150,N_2274);
nor U3802 (N_3802,N_697,N_405);
xor U3803 (N_3803,N_1391,N_1853);
nand U3804 (N_3804,N_17,N_1417);
nand U3805 (N_3805,N_603,N_157);
nor U3806 (N_3806,N_70,N_1789);
xnor U3807 (N_3807,N_1626,N_1107);
or U3808 (N_3808,N_2839,N_2542);
nor U3809 (N_3809,N_2591,N_1193);
xor U3810 (N_3810,N_628,N_1748);
and U3811 (N_3811,N_1532,N_2742);
xor U3812 (N_3812,N_197,N_2753);
and U3813 (N_3813,N_449,N_1165);
and U3814 (N_3814,N_424,N_977);
nor U3815 (N_3815,N_860,N_1640);
nor U3816 (N_3816,N_275,N_1652);
xnor U3817 (N_3817,N_204,N_2246);
nand U3818 (N_3818,N_2998,N_615);
xnor U3819 (N_3819,N_2017,N_2674);
nor U3820 (N_3820,N_470,N_2012);
and U3821 (N_3821,N_1851,N_2934);
nor U3822 (N_3822,N_1720,N_2219);
and U3823 (N_3823,N_1177,N_2263);
or U3824 (N_3824,N_126,N_251);
or U3825 (N_3825,N_2407,N_155);
nand U3826 (N_3826,N_2441,N_300);
nand U3827 (N_3827,N_1028,N_609);
or U3828 (N_3828,N_1225,N_1250);
xnor U3829 (N_3829,N_720,N_2244);
and U3830 (N_3830,N_2380,N_2726);
nor U3831 (N_3831,N_1129,N_2848);
nor U3832 (N_3832,N_882,N_2522);
xor U3833 (N_3833,N_2673,N_1667);
xnor U3834 (N_3834,N_928,N_231);
xor U3835 (N_3835,N_383,N_2161);
nand U3836 (N_3836,N_1386,N_1232);
nor U3837 (N_3837,N_2331,N_1629);
or U3838 (N_3838,N_722,N_2361);
and U3839 (N_3839,N_106,N_101);
nor U3840 (N_3840,N_1200,N_135);
xor U3841 (N_3841,N_764,N_1666);
or U3842 (N_3842,N_1723,N_2835);
and U3843 (N_3843,N_2035,N_2816);
or U3844 (N_3844,N_1060,N_58);
nand U3845 (N_3845,N_2743,N_2027);
nand U3846 (N_3846,N_2334,N_1185);
nand U3847 (N_3847,N_2065,N_782);
or U3848 (N_3848,N_824,N_2198);
nand U3849 (N_3849,N_399,N_1795);
or U3850 (N_3850,N_2188,N_59);
and U3851 (N_3851,N_813,N_3018);
nand U3852 (N_3852,N_2413,N_1971);
xor U3853 (N_3853,N_704,N_2575);
xor U3854 (N_3854,N_2379,N_1307);
nor U3855 (N_3855,N_1996,N_907);
and U3856 (N_3856,N_91,N_2878);
nand U3857 (N_3857,N_2058,N_306);
nand U3858 (N_3858,N_555,N_1384);
nand U3859 (N_3859,N_190,N_2600);
or U3860 (N_3860,N_1186,N_2016);
and U3861 (N_3861,N_506,N_995);
nand U3862 (N_3862,N_635,N_1159);
nor U3863 (N_3863,N_2122,N_437);
nand U3864 (N_3864,N_788,N_1423);
and U3865 (N_3865,N_1548,N_1710);
and U3866 (N_3866,N_2993,N_2349);
nand U3867 (N_3867,N_2080,N_372);
or U3868 (N_3868,N_2110,N_1084);
or U3869 (N_3869,N_279,N_2004);
xor U3870 (N_3870,N_1146,N_1788);
xor U3871 (N_3871,N_1882,N_662);
or U3872 (N_3872,N_2335,N_47);
or U3873 (N_3873,N_1078,N_2488);
and U3874 (N_3874,N_2617,N_2833);
nand U3875 (N_3875,N_1001,N_1017);
or U3876 (N_3876,N_818,N_2748);
or U3877 (N_3877,N_1530,N_1987);
or U3878 (N_3878,N_2530,N_2445);
nor U3879 (N_3879,N_447,N_581);
or U3880 (N_3880,N_748,N_2295);
nand U3881 (N_3881,N_2898,N_655);
nand U3882 (N_3882,N_2185,N_209);
nor U3883 (N_3883,N_1718,N_1825);
xor U3884 (N_3884,N_422,N_1317);
and U3885 (N_3885,N_1202,N_2690);
xnor U3886 (N_3886,N_2468,N_636);
and U3887 (N_3887,N_534,N_792);
and U3888 (N_3888,N_911,N_776);
and U3889 (N_3889,N_1347,N_1584);
xor U3890 (N_3890,N_2320,N_481);
and U3891 (N_3891,N_1227,N_1432);
xor U3892 (N_3892,N_696,N_850);
and U3893 (N_3893,N_166,N_1338);
or U3894 (N_3894,N_620,N_1113);
or U3895 (N_3895,N_1249,N_1905);
or U3896 (N_3896,N_2719,N_2172);
nand U3897 (N_3897,N_3007,N_831);
nand U3898 (N_3898,N_3030,N_1006);
nor U3899 (N_3899,N_1524,N_1692);
nor U3900 (N_3900,N_3056,N_1178);
nand U3901 (N_3901,N_836,N_1766);
nor U3902 (N_3902,N_66,N_3038);
xnor U3903 (N_3903,N_807,N_2852);
or U3904 (N_3904,N_2419,N_943);
xnor U3905 (N_3905,N_1768,N_2015);
nand U3906 (N_3906,N_2278,N_955);
or U3907 (N_3907,N_1039,N_714);
and U3908 (N_3908,N_2774,N_1761);
nor U3909 (N_3909,N_2366,N_299);
and U3910 (N_3910,N_2706,N_2537);
or U3911 (N_3911,N_1474,N_771);
nand U3912 (N_3912,N_1387,N_1504);
nand U3913 (N_3913,N_1551,N_2181);
and U3914 (N_3914,N_1239,N_1816);
nand U3915 (N_3915,N_342,N_1623);
nand U3916 (N_3916,N_576,N_2460);
nor U3917 (N_3917,N_2670,N_1119);
and U3918 (N_3918,N_175,N_2233);
or U3919 (N_3919,N_1133,N_2049);
or U3920 (N_3920,N_2256,N_2717);
nand U3921 (N_3921,N_2507,N_1408);
and U3922 (N_3922,N_1659,N_1983);
nand U3923 (N_3923,N_352,N_2880);
or U3924 (N_3924,N_201,N_1739);
or U3925 (N_3925,N_183,N_2868);
nor U3926 (N_3926,N_2539,N_2367);
and U3927 (N_3927,N_1995,N_2269);
or U3928 (N_3928,N_448,N_2730);
and U3929 (N_3929,N_2817,N_2447);
xnor U3930 (N_3930,N_811,N_232);
xnor U3931 (N_3931,N_84,N_2479);
or U3932 (N_3932,N_1539,N_2667);
nor U3933 (N_3933,N_881,N_735);
or U3934 (N_3934,N_2508,N_3113);
nand U3935 (N_3935,N_442,N_1327);
or U3936 (N_3936,N_1181,N_676);
nand U3937 (N_3937,N_2609,N_2302);
and U3938 (N_3938,N_2996,N_2651);
nor U3939 (N_3939,N_417,N_1248);
xnor U3940 (N_3940,N_1752,N_1392);
nor U3941 (N_3941,N_2523,N_2328);
xnor U3942 (N_3942,N_2206,N_1135);
and U3943 (N_3943,N_460,N_600);
xnor U3944 (N_3944,N_3070,N_2858);
and U3945 (N_3945,N_1067,N_1197);
xnor U3946 (N_3946,N_1495,N_1254);
or U3947 (N_3947,N_387,N_611);
xor U3948 (N_3948,N_1288,N_1745);
nand U3949 (N_3949,N_2502,N_2758);
or U3950 (N_3950,N_1013,N_2757);
nor U3951 (N_3951,N_2601,N_1166);
and U3952 (N_3952,N_325,N_72);
nand U3953 (N_3953,N_2095,N_1514);
and U3954 (N_3954,N_732,N_2033);
and U3955 (N_3955,N_749,N_1075);
nor U3956 (N_3956,N_15,N_2703);
and U3957 (N_3957,N_2438,N_1508);
or U3958 (N_3958,N_1822,N_28);
and U3959 (N_3959,N_1878,N_1380);
xnor U3960 (N_3960,N_288,N_2378);
or U3961 (N_3961,N_2045,N_2077);
nor U3962 (N_3962,N_3026,N_2401);
xor U3963 (N_3963,N_297,N_1840);
and U3964 (N_3964,N_338,N_191);
or U3965 (N_3965,N_610,N_1940);
nand U3966 (N_3966,N_2308,N_2533);
nor U3967 (N_3967,N_2271,N_2739);
and U3968 (N_3968,N_2740,N_785);
xor U3969 (N_3969,N_2620,N_1747);
nor U3970 (N_3970,N_56,N_2133);
nor U3971 (N_3971,N_1597,N_2327);
nor U3972 (N_3972,N_2532,N_1662);
xor U3973 (N_3973,N_926,N_679);
or U3974 (N_3974,N_1349,N_2089);
xor U3975 (N_3975,N_2861,N_2598);
or U3976 (N_3976,N_2842,N_933);
nand U3977 (N_3977,N_767,N_3108);
nand U3978 (N_3978,N_552,N_1424);
xnor U3979 (N_3979,N_942,N_1388);
or U3980 (N_3980,N_2979,N_133);
and U3981 (N_3981,N_561,N_1606);
nand U3982 (N_3982,N_1886,N_2978);
or U3983 (N_3983,N_472,N_63);
or U3984 (N_3984,N_1963,N_2911);
xor U3985 (N_3985,N_2345,N_2551);
and U3986 (N_3986,N_2767,N_1373);
xnor U3987 (N_3987,N_1515,N_761);
nand U3988 (N_3988,N_2536,N_1657);
or U3989 (N_3989,N_3064,N_1160);
or U3990 (N_3990,N_699,N_1845);
and U3991 (N_3991,N_3073,N_2178);
nand U3992 (N_3992,N_2386,N_2800);
nor U3993 (N_3993,N_185,N_2596);
xnor U3994 (N_3994,N_2724,N_835);
nor U3995 (N_3995,N_1404,N_730);
and U3996 (N_3996,N_2954,N_1624);
nor U3997 (N_3997,N_805,N_2470);
and U3998 (N_3998,N_2194,N_2141);
nor U3999 (N_3999,N_2971,N_2495);
or U4000 (N_4000,N_1957,N_2034);
or U4001 (N_4001,N_2595,N_3116);
or U4002 (N_4002,N_474,N_1800);
nand U4003 (N_4003,N_2422,N_1473);
or U4004 (N_4004,N_2487,N_2584);
and U4005 (N_4005,N_2697,N_2564);
nor U4006 (N_4006,N_1484,N_2462);
or U4007 (N_4007,N_215,N_2888);
or U4008 (N_4008,N_1033,N_1428);
and U4009 (N_4009,N_116,N_2691);
and U4010 (N_4010,N_524,N_1703);
nor U4011 (N_4011,N_1763,N_30);
or U4012 (N_4012,N_3077,N_112);
and U4013 (N_4013,N_783,N_1654);
or U4014 (N_4014,N_2859,N_2434);
xnor U4015 (N_4015,N_1087,N_146);
nand U4016 (N_4016,N_2031,N_206);
and U4017 (N_4017,N_3025,N_55);
nor U4018 (N_4018,N_1485,N_210);
nor U4019 (N_4019,N_2497,N_2659);
nor U4020 (N_4020,N_1622,N_2338);
or U4021 (N_4021,N_2318,N_1982);
and U4022 (N_4022,N_567,N_1501);
nor U4023 (N_4023,N_36,N_1570);
nor U4024 (N_4024,N_1790,N_2446);
or U4025 (N_4025,N_3119,N_1152);
nor U4026 (N_4026,N_608,N_1051);
nor U4027 (N_4027,N_823,N_1869);
or U4028 (N_4028,N_2249,N_1356);
xor U4029 (N_4029,N_1125,N_1009);
and U4030 (N_4030,N_2139,N_586);
or U4031 (N_4031,N_1314,N_478);
xor U4032 (N_4032,N_73,N_356);
nand U4033 (N_4033,N_1030,N_574);
nand U4034 (N_4034,N_646,N_1027);
xor U4035 (N_4035,N_1049,N_1036);
xor U4036 (N_4036,N_235,N_2450);
nor U4037 (N_4037,N_708,N_815);
or U4038 (N_4038,N_1881,N_1981);
or U4039 (N_4039,N_2251,N_1080);
nand U4040 (N_4040,N_2645,N_1838);
or U4041 (N_4041,N_230,N_2240);
nor U4042 (N_4042,N_794,N_1687);
nand U4043 (N_4043,N_362,N_2546);
or U4044 (N_4044,N_1764,N_674);
nand U4045 (N_4045,N_725,N_1618);
nand U4046 (N_4046,N_96,N_2573);
or U4047 (N_4047,N_2343,N_2108);
nand U4048 (N_4048,N_2467,N_2735);
nand U4049 (N_4049,N_1194,N_2669);
or U4050 (N_4050,N_1674,N_369);
xnor U4051 (N_4051,N_349,N_1183);
nor U4052 (N_4052,N_775,N_320);
or U4053 (N_4053,N_2239,N_311);
nor U4054 (N_4054,N_980,N_1600);
xor U4055 (N_4055,N_2797,N_1528);
nor U4056 (N_4056,N_2506,N_1222);
nor U4057 (N_4057,N_923,N_2675);
or U4058 (N_4058,N_2559,N_1874);
xnor U4059 (N_4059,N_1297,N_2568);
and U4060 (N_4060,N_335,N_2922);
nor U4061 (N_4061,N_921,N_2115);
nor U4062 (N_4062,N_629,N_686);
or U4063 (N_4063,N_2553,N_469);
and U4064 (N_4064,N_1661,N_2484);
nor U4065 (N_4065,N_1750,N_901);
xnor U4066 (N_4066,N_491,N_1785);
nand U4067 (N_4067,N_479,N_114);
nor U4068 (N_4068,N_1520,N_1321);
or U4069 (N_4069,N_2290,N_2090);
or U4070 (N_4070,N_1712,N_1407);
and U4071 (N_4071,N_1025,N_2699);
or U4072 (N_4072,N_1331,N_2879);
nor U4073 (N_4073,N_1612,N_346);
xor U4074 (N_4074,N_2633,N_2720);
or U4075 (N_4075,N_1979,N_1744);
nand U4076 (N_4076,N_2969,N_457);
nor U4077 (N_4077,N_2809,N_2157);
nor U4078 (N_4078,N_660,N_1769);
or U4079 (N_4079,N_2821,N_2763);
nand U4080 (N_4080,N_2063,N_69);
xor U4081 (N_4081,N_1014,N_1757);
and U4082 (N_4082,N_2007,N_1787);
and U4083 (N_4083,N_1287,N_1360);
nand U4084 (N_4084,N_2214,N_353);
or U4085 (N_4085,N_1134,N_425);
nor U4086 (N_4086,N_1582,N_1208);
nor U4087 (N_4087,N_134,N_604);
nor U4088 (N_4088,N_1525,N_1023);
xnor U4089 (N_4089,N_3066,N_1110);
and U4090 (N_4090,N_308,N_891);
and U4091 (N_4091,N_1427,N_1220);
nor U4092 (N_4092,N_1189,N_400);
and U4093 (N_4093,N_959,N_2412);
nor U4094 (N_4094,N_0,N_2150);
or U4095 (N_4095,N_207,N_1943);
nor U4096 (N_4096,N_841,N_2710);
and U4097 (N_4097,N_768,N_3005);
or U4098 (N_4098,N_3023,N_2904);
xor U4099 (N_4099,N_1594,N_1198);
and U4100 (N_4100,N_289,N_1865);
nand U4101 (N_4101,N_2623,N_2296);
and U4102 (N_4102,N_1592,N_1422);
or U4103 (N_4103,N_1430,N_1345);
nand U4104 (N_4104,N_2374,N_766);
and U4105 (N_4105,N_1877,N_595);
and U4106 (N_4106,N_2176,N_1729);
nand U4107 (N_4107,N_2424,N_315);
and U4108 (N_4108,N_2578,N_1988);
or U4109 (N_4109,N_750,N_1354);
xnor U4110 (N_4110,N_1382,N_2435);
or U4111 (N_4111,N_1043,N_2170);
or U4112 (N_4112,N_1552,N_2281);
nor U4113 (N_4113,N_2558,N_1765);
or U4114 (N_4114,N_1132,N_2783);
xor U4115 (N_4115,N_1007,N_1554);
nand U4116 (N_4116,N_1330,N_2490);
and U4117 (N_4117,N_2882,N_67);
nand U4118 (N_4118,N_2521,N_845);
and U4119 (N_4119,N_774,N_2947);
or U4120 (N_4120,N_123,N_3092);
and U4121 (N_4121,N_1305,N_269);
nor U4122 (N_4122,N_2120,N_498);
nand U4123 (N_4123,N_2731,N_1773);
nor U4124 (N_4124,N_2091,N_571);
or U4125 (N_4125,N_992,N_1353);
nand U4126 (N_4126,N_428,N_873);
nand U4127 (N_4127,N_2920,N_1414);
nor U4128 (N_4128,N_1128,N_1679);
nor U4129 (N_4129,N_391,N_1863);
nand U4130 (N_4130,N_910,N_2654);
and U4131 (N_4131,N_1162,N_780);
and U4132 (N_4132,N_2589,N_1214);
xnor U4133 (N_4133,N_2959,N_2579);
nand U4134 (N_4134,N_88,N_3111);
nor U4135 (N_4135,N_1879,N_1368);
nand U4136 (N_4136,N_35,N_333);
and U4137 (N_4137,N_3042,N_1058);
nor U4138 (N_4138,N_2864,N_1409);
xor U4139 (N_4139,N_2313,N_467);
nand U4140 (N_4140,N_1884,N_2459);
or U4141 (N_4141,N_410,N_2329);
and U4142 (N_4142,N_2865,N_2906);
nor U4143 (N_4143,N_2086,N_2997);
xor U4144 (N_4144,N_501,N_1964);
nand U4145 (N_4145,N_144,N_990);
and U4146 (N_4146,N_3053,N_1052);
nand U4147 (N_4147,N_529,N_3024);
and U4148 (N_4148,N_2228,N_1969);
xnor U4149 (N_4149,N_905,N_32);
xnor U4150 (N_4150,N_558,N_1890);
nor U4151 (N_4151,N_2668,N_1734);
and U4152 (N_4152,N_1401,N_158);
or U4153 (N_4153,N_132,N_2711);
xor U4154 (N_4154,N_3095,N_1824);
nand U4155 (N_4155,N_2040,N_1230);
nor U4156 (N_4156,N_1634,N_290);
nand U4157 (N_4157,N_429,N_1441);
nand U4158 (N_4158,N_3013,N_1443);
nand U4159 (N_4159,N_698,N_759);
nand U4160 (N_4160,N_945,N_736);
xnor U4161 (N_4161,N_503,N_2732);
nor U4162 (N_4162,N_832,N_39);
xor U4163 (N_4163,N_266,N_770);
nand U4164 (N_4164,N_2064,N_2709);
nand U4165 (N_4165,N_441,N_354);
and U4166 (N_4166,N_458,N_2805);
xor U4167 (N_4167,N_1678,N_1999);
nor U4168 (N_4168,N_2915,N_2452);
nor U4169 (N_4169,N_162,N_962);
nand U4170 (N_4170,N_522,N_1468);
nand U4171 (N_4171,N_2662,N_2672);
xnor U4172 (N_4172,N_956,N_1531);
nor U4173 (N_4173,N_1385,N_2344);
nand U4174 (N_4174,N_394,N_2275);
or U4175 (N_4175,N_2075,N_2902);
nor U4176 (N_4176,N_3049,N_7);
nand U4177 (N_4177,N_1962,N_1367);
nand U4178 (N_4178,N_3009,N_872);
nor U4179 (N_4179,N_2686,N_1730);
nor U4180 (N_4180,N_1545,N_2819);
nand U4181 (N_4181,N_2901,N_723);
xor U4182 (N_4182,N_705,N_1895);
nor U4183 (N_4183,N_1846,N_2873);
nand U4184 (N_4184,N_3120,N_531);
xnor U4185 (N_4185,N_2162,N_1403);
and U4186 (N_4186,N_778,N_944);
nor U4187 (N_4187,N_1451,N_401);
xor U4188 (N_4188,N_1434,N_2948);
nand U4189 (N_4189,N_1299,N_1772);
or U4190 (N_4190,N_2014,N_960);
and U4191 (N_4191,N_1915,N_2280);
and U4192 (N_4192,N_2292,N_1523);
and U4193 (N_4193,N_2291,N_213);
nand U4194 (N_4194,N_1026,N_3048);
nor U4195 (N_4195,N_376,N_1095);
xnor U4196 (N_4196,N_2513,N_2392);
and U4197 (N_4197,N_145,N_3062);
nor U4198 (N_4198,N_1020,N_1749);
or U4199 (N_4199,N_1040,N_1342);
nand U4200 (N_4200,N_3031,N_1082);
nand U4201 (N_4201,N_913,N_861);
or U4202 (N_4202,N_1771,N_2417);
nand U4203 (N_4203,N_790,N_1818);
nand U4204 (N_4204,N_2581,N_2678);
and U4205 (N_4205,N_1546,N_2230);
xnor U4206 (N_4206,N_220,N_2258);
and U4207 (N_4207,N_2104,N_1094);
and U4208 (N_4208,N_1289,N_1529);
xor U4209 (N_4209,N_1691,N_1376);
and U4210 (N_4210,N_2628,N_2671);
and U4211 (N_4211,N_2789,N_363);
or U4212 (N_4212,N_2877,N_806);
nand U4213 (N_4213,N_2259,N_255);
nor U4214 (N_4214,N_46,N_641);
or U4215 (N_4215,N_382,N_1814);
or U4216 (N_4216,N_294,N_2405);
and U4217 (N_4217,N_2389,N_1100);
nand U4218 (N_4218,N_2635,N_797);
nor U4219 (N_4219,N_1615,N_2128);
and U4220 (N_4220,N_1728,N_2330);
nor U4221 (N_4221,N_1278,N_2241);
or U4222 (N_4222,N_1096,N_607);
and U4223 (N_4223,N_3083,N_758);
nor U4224 (N_4224,N_2847,N_1064);
xnor U4225 (N_4225,N_1857,N_415);
xnor U4226 (N_4226,N_78,N_1137);
xnor U4227 (N_4227,N_466,N_784);
and U4228 (N_4228,N_1826,N_2619);
xor U4229 (N_4229,N_2284,N_1086);
and U4230 (N_4230,N_541,N_2802);
xor U4231 (N_4231,N_2085,N_2872);
or U4232 (N_4232,N_2606,N_2159);
or U4233 (N_4233,N_968,N_601);
xor U4234 (N_4234,N_2492,N_1589);
xnor U4235 (N_4235,N_820,N_75);
nor U4236 (N_4236,N_455,N_517);
or U4237 (N_4237,N_1665,N_1453);
and U4238 (N_4238,N_930,N_1037);
nand U4239 (N_4239,N_2995,N_939);
nor U4240 (N_4240,N_345,N_690);
and U4241 (N_4241,N_1643,N_1411);
or U4242 (N_4242,N_1741,N_304);
or U4243 (N_4243,N_1617,N_2301);
nor U4244 (N_4244,N_1852,N_1203);
nand U4245 (N_4245,N_2416,N_318);
and U4246 (N_4246,N_1211,N_2999);
or U4247 (N_4247,N_1601,N_2309);
nor U4248 (N_4248,N_1171,N_2268);
nand U4249 (N_4249,N_724,N_1970);
and U4250 (N_4250,N_257,N_2073);
nand U4251 (N_4251,N_265,N_2037);
xor U4252 (N_4252,N_141,N_1285);
xor U4253 (N_4253,N_2762,N_234);
or U4254 (N_4254,N_843,N_757);
nand U4255 (N_4255,N_1187,N_585);
xor U4256 (N_4256,N_2384,N_1972);
nor U4257 (N_4257,N_1416,N_1325);
nor U4258 (N_4258,N_2423,N_433);
xnor U4259 (N_4259,N_2907,N_2755);
and U4260 (N_4260,N_965,N_2509);
nand U4261 (N_4261,N_1149,N_2146);
xor U4262 (N_4262,N_2807,N_564);
xnor U4263 (N_4263,N_1677,N_1797);
or U4264 (N_4264,N_143,N_119);
nand U4265 (N_4265,N_1199,N_475);
nor U4266 (N_4266,N_1557,N_633);
or U4267 (N_4267,N_1238,N_302);
or U4268 (N_4268,N_2876,N_99);
or U4269 (N_4269,N_1770,N_2884);
or U4270 (N_4270,N_489,N_1131);
xor U4271 (N_4271,N_1341,N_1602);
xor U4272 (N_4272,N_883,N_2323);
nand U4273 (N_4273,N_2892,N_2682);
nand U4274 (N_4274,N_463,N_2234);
xor U4275 (N_4275,N_3072,N_154);
nand U4276 (N_4276,N_657,N_1827);
xor U4277 (N_4277,N_233,N_700);
nand U4278 (N_4278,N_2229,N_459);
and U4279 (N_4279,N_2634,N_1778);
or U4280 (N_4280,N_2639,N_1462);
nand U4281 (N_4281,N_1081,N_14);
nand U4282 (N_4282,N_486,N_2255);
xor U4283 (N_4283,N_996,N_2788);
xor U4284 (N_4284,N_1169,N_1123);
nand U4285 (N_4285,N_1613,N_2857);
or U4286 (N_4286,N_2305,N_2560);
or U4287 (N_4287,N_90,N_277);
or U4288 (N_4288,N_1426,N_1864);
or U4289 (N_4289,N_2149,N_2279);
nor U4290 (N_4290,N_2607,N_1916);
xnor U4291 (N_4291,N_1413,N_719);
nor U4292 (N_4292,N_1098,N_713);
nand U4293 (N_4293,N_397,N_1010);
nand U4294 (N_4294,N_1180,N_669);
nand U4295 (N_4295,N_250,N_1454);
and U4296 (N_4296,N_2655,N_411);
nand U4297 (N_4297,N_3004,N_1071);
or U4298 (N_4298,N_293,N_360);
nand U4299 (N_4299,N_2137,N_2897);
xnor U4300 (N_4300,N_237,N_640);
nand U4301 (N_4301,N_2084,N_1034);
nor U4302 (N_4302,N_987,N_236);
or U4303 (N_4303,N_453,N_1823);
nor U4304 (N_4304,N_1316,N_1389);
or U4305 (N_4305,N_684,N_1920);
and U4306 (N_4306,N_419,N_1255);
nor U4307 (N_4307,N_895,N_1439);
or U4308 (N_4308,N_2790,N_1664);
nand U4309 (N_4309,N_2622,N_2365);
xnor U4310 (N_4310,N_2860,N_888);
nand U4311 (N_4311,N_2364,N_709);
nand U4312 (N_4312,N_2306,N_1951);
nand U4313 (N_4313,N_2562,N_3027);
or U4314 (N_4314,N_1418,N_223);
nor U4315 (N_4315,N_2444,N_2235);
and U4316 (N_4316,N_1054,N_261);
nand U4317 (N_4317,N_1860,N_1400);
nand U4318 (N_4318,N_983,N_2148);
and U4319 (N_4319,N_2550,N_738);
nor U4320 (N_4320,N_2563,N_1753);
nand U4321 (N_4321,N_2749,N_2632);
nor U4322 (N_4322,N_855,N_2801);
and U4323 (N_4323,N_2965,N_1304);
or U4324 (N_4324,N_1103,N_2039);
xor U4325 (N_4325,N_3124,N_426);
xnor U4326 (N_4326,N_2569,N_654);
or U4327 (N_4327,N_3063,N_450);
nor U4328 (N_4328,N_1252,N_2593);
or U4329 (N_4329,N_1312,N_1653);
xnor U4330 (N_4330,N_1217,N_1902);
and U4331 (N_4331,N_737,N_2810);
nor U4332 (N_4332,N_421,N_1136);
or U4333 (N_4333,N_452,N_1437);
and U4334 (N_4334,N_2989,N_717);
and U4335 (N_4335,N_2160,N_402);
or U4336 (N_4336,N_622,N_2496);
and U4337 (N_4337,N_899,N_2443);
nand U4338 (N_4338,N_1168,N_521);
nor U4339 (N_4339,N_2649,N_932);
or U4340 (N_4340,N_374,N_802);
xnor U4341 (N_4341,N_1901,N_1251);
and U4342 (N_4342,N_2544,N_2342);
nand U4343 (N_4343,N_1502,N_1611);
nor U4344 (N_4344,N_3032,N_282);
xor U4345 (N_4345,N_540,N_2896);
xnor U4346 (N_4346,N_1340,N_2604);
or U4347 (N_4347,N_328,N_2841);
nand U4348 (N_4348,N_647,N_413);
nor U4349 (N_4349,N_2169,N_57);
nand U4350 (N_4350,N_1956,N_1270);
nand U4351 (N_4351,N_2289,N_1549);
nor U4352 (N_4352,N_533,N_2061);
nor U4353 (N_4353,N_2472,N_878);
xnor U4354 (N_4354,N_2317,N_1767);
xnor U4355 (N_4355,N_198,N_1104);
xnor U4356 (N_4356,N_1588,N_2175);
nor U4357 (N_4357,N_44,N_2223);
and U4358 (N_4358,N_2455,N_416);
xor U4359 (N_4359,N_1715,N_2300);
nor U4360 (N_4360,N_2371,N_1458);
xor U4361 (N_4361,N_461,N_1985);
xnor U4362 (N_4362,N_2986,N_2261);
or U4363 (N_4363,N_2653,N_941);
nand U4364 (N_4364,N_2944,N_1932);
nand U4365 (N_4365,N_710,N_2956);
xnor U4366 (N_4366,N_2314,N_666);
and U4367 (N_4367,N_3118,N_331);
and U4368 (N_4368,N_2368,N_2076);
nor U4369 (N_4369,N_471,N_1226);
and U4370 (N_4370,N_966,N_327);
xor U4371 (N_4371,N_1793,N_2390);
xnor U4372 (N_4372,N_1812,N_1585);
nand U4373 (N_4373,N_591,N_510);
or U4374 (N_4374,N_2023,N_542);
xnor U4375 (N_4375,N_1000,N_2681);
xor U4376 (N_4376,N_1518,N_1938);
nand U4377 (N_4377,N_1704,N_2844);
or U4378 (N_4378,N_1506,N_139);
and U4379 (N_4379,N_1176,N_1261);
xnor U4380 (N_4380,N_3117,N_833);
nand U4381 (N_4381,N_2190,N_1143);
and U4382 (N_4382,N_884,N_115);
and U4383 (N_4383,N_323,N_2910);
and U4384 (N_4384,N_1393,N_762);
or U4385 (N_4385,N_61,N_1306);
and U4386 (N_4386,N_1262,N_2273);
and U4387 (N_4387,N_975,N_2913);
xnor U4388 (N_4388,N_902,N_390);
nor U4389 (N_4389,N_83,N_2764);
nand U4390 (N_4390,N_1740,N_683);
and U4391 (N_4391,N_1912,N_2092);
or U4392 (N_4392,N_940,N_242);
nand U4393 (N_4393,N_834,N_2815);
xnor U4394 (N_4394,N_1540,N_41);
xor U4395 (N_4395,N_563,N_2421);
or U4396 (N_4396,N_2676,N_606);
xnor U4397 (N_4397,N_2199,N_2612);
xor U4398 (N_4398,N_120,N_1565);
and U4399 (N_4399,N_1875,N_1577);
nand U4400 (N_4400,N_2840,N_3041);
xor U4401 (N_4401,N_1164,N_2597);
nand U4402 (N_4402,N_1145,N_142);
nor U4403 (N_4403,N_1253,N_2970);
nand U4404 (N_4404,N_278,N_6);
xnor U4405 (N_4405,N_1609,N_1522);
nor U4406 (N_4406,N_2894,N_2870);
and U4407 (N_4407,N_3115,N_1645);
nor U4408 (N_4408,N_384,N_1655);
xor U4409 (N_4409,N_519,N_1365);
or U4410 (N_4410,N_2245,N_848);
or U4411 (N_4411,N_590,N_1069);
or U4412 (N_4412,N_291,N_2304);
and U4413 (N_4413,N_488,N_2552);
xnor U4414 (N_4414,N_86,N_619);
or U4415 (N_4415,N_339,N_1218);
nor U4416 (N_4416,N_1580,N_2962);
nand U4417 (N_4417,N_2333,N_1046);
nor U4418 (N_4418,N_826,N_245);
xor U4419 (N_4419,N_2018,N_1296);
xor U4420 (N_4420,N_1155,N_2938);
or U4421 (N_4421,N_1663,N_1467);
or U4422 (N_4422,N_734,N_1917);
and U4423 (N_4423,N_1318,N_2449);
nor U4424 (N_4424,N_2722,N_702);
and U4425 (N_4425,N_2028,N_1234);
or U4426 (N_4426,N_1493,N_296);
nand U4427 (N_4427,N_779,N_2661);
nor U4428 (N_4428,N_621,N_2297);
nand U4429 (N_4429,N_1836,N_2772);
or U4430 (N_4430,N_27,N_2116);
or U4431 (N_4431,N_1844,N_680);
nor U4432 (N_4432,N_1830,N_1743);
nor U4433 (N_4433,N_2621,N_1512);
nor U4434 (N_4434,N_432,N_2083);
xor U4435 (N_4435,N_1170,N_553);
and U4436 (N_4436,N_2147,N_1019);
nor U4437 (N_4437,N_312,N_1621);
nor U4438 (N_4438,N_2432,N_2476);
xnor U4439 (N_4439,N_1302,N_2153);
nand U4440 (N_4440,N_712,N_1903);
or U4441 (N_4441,N_1700,N_2588);
xnor U4442 (N_4442,N_1269,N_1862);
xnor U4443 (N_4443,N_247,N_140);
nor U4444 (N_4444,N_3057,N_2926);
or U4445 (N_4445,N_2950,N_1282);
or U4446 (N_4446,N_180,N_2785);
nand U4447 (N_4447,N_2400,N_559);
and U4448 (N_4448,N_359,N_2925);
nand U4449 (N_4449,N_1794,N_958);
and U4450 (N_4450,N_2914,N_1521);
and U4451 (N_4451,N_2759,N_1536);
xor U4452 (N_4452,N_1883,N_267);
and U4453 (N_4453,N_1542,N_1117);
xnor U4454 (N_4454,N_2512,N_931);
or U4455 (N_4455,N_976,N_2262);
nand U4456 (N_4456,N_1922,N_1379);
nand U4457 (N_4457,N_2549,N_1628);
nor U4458 (N_4458,N_238,N_2491);
or U4459 (N_4459,N_847,N_2751);
nand U4460 (N_4460,N_627,N_642);
or U4461 (N_4461,N_310,N_2688);
and U4462 (N_4462,N_2415,N_221);
nand U4463 (N_4463,N_2582,N_1668);
nor U4464 (N_4464,N_1942,N_837);
nand U4465 (N_4465,N_917,N_915);
nand U4466 (N_4466,N_2155,N_3);
nor U4467 (N_4467,N_1587,N_1147);
xor U4468 (N_4468,N_1558,N_821);
nand U4469 (N_4469,N_1406,N_2282);
or U4470 (N_4470,N_1257,N_2985);
xnor U4471 (N_4471,N_2796,N_1656);
and U4472 (N_4472,N_592,N_2637);
xor U4473 (N_4473,N_2866,N_49);
nor U4474 (N_4474,N_337,N_1);
nand U4475 (N_4475,N_1053,N_490);
nor U4476 (N_4476,N_2525,N_195);
or U4477 (N_4477,N_1693,N_1480);
and U4478 (N_4478,N_2804,N_45);
xor U4479 (N_4479,N_2707,N_1083);
or U4480 (N_4480,N_2440,N_301);
nor U4481 (N_4481,N_1479,N_1896);
xor U4482 (N_4482,N_110,N_1492);
xnor U4483 (N_4483,N_1138,N_644);
nand U4484 (N_4484,N_1102,N_1295);
nand U4485 (N_4485,N_523,N_653);
or U4486 (N_4486,N_652,N_971);
xor U4487 (N_4487,N_1410,N_2418);
xnor U4488 (N_4488,N_1724,N_2357);
or U4489 (N_4489,N_2663,N_111);
nor U4490 (N_4490,N_1175,N_199);
and U4491 (N_4491,N_2647,N_2052);
xor U4492 (N_4492,N_1344,N_588);
or U4493 (N_4493,N_3037,N_1923);
nor U4494 (N_4494,N_324,N_1742);
or U4495 (N_4495,N_149,N_1099);
xnor U4496 (N_4496,N_1370,N_2254);
xnor U4497 (N_4497,N_2773,N_2733);
and U4498 (N_4498,N_1727,N_1708);
and U4499 (N_4499,N_2481,N_1924);
nor U4500 (N_4500,N_1243,N_127);
nor U4501 (N_4501,N_82,N_393);
or U4502 (N_4502,N_632,N_1293);
nor U4503 (N_4503,N_1085,N_1802);
nor U4504 (N_4504,N_513,N_3061);
or U4505 (N_4505,N_1992,N_1799);
or U4506 (N_4506,N_29,N_2025);
xor U4507 (N_4507,N_1320,N_97);
or U4508 (N_4508,N_2702,N_1644);
nor U4509 (N_4509,N_2946,N_937);
and U4510 (N_4510,N_994,N_1021);
and U4511 (N_4511,N_1469,N_2402);
nor U4512 (N_4512,N_2850,N_2716);
nor U4513 (N_4513,N_580,N_582);
nand U4514 (N_4514,N_967,N_1579);
or U4515 (N_4515,N_1990,N_492);
xor U4516 (N_4516,N_1870,N_2862);
and U4517 (N_4517,N_1736,N_3052);
xnor U4518 (N_4518,N_1337,N_1264);
xor U4519 (N_4519,N_2519,N_1108);
xor U4520 (N_4520,N_358,N_594);
and U4521 (N_4521,N_129,N_2899);
nor U4522 (N_4522,N_2574,N_2991);
nor U4523 (N_4523,N_1616,N_2238);
and U4524 (N_4524,N_2916,N_1246);
and U4525 (N_4525,N_3014,N_226);
nor U4526 (N_4526,N_634,N_1048);
and U4527 (N_4527,N_3039,N_2321);
nand U4528 (N_4528,N_2212,N_515);
nor U4529 (N_4529,N_1343,N_357);
and U4530 (N_4530,N_2020,N_1562);
or U4531 (N_4531,N_1841,N_1625);
xnor U4532 (N_4532,N_1936,N_285);
and U4533 (N_4533,N_1945,N_440);
nor U4534 (N_4534,N_1363,N_2337);
or U4535 (N_4535,N_2656,N_2770);
and U4536 (N_4536,N_786,N_42);
xor U4537 (N_4537,N_1516,N_691);
nor U4538 (N_4538,N_2961,N_1497);
xnor U4539 (N_4539,N_2694,N_569);
or U4540 (N_4540,N_871,N_2117);
or U4541 (N_4541,N_1792,N_1696);
and U4542 (N_4542,N_2307,N_1735);
or U4543 (N_4543,N_176,N_1843);
nand U4544 (N_4544,N_12,N_1854);
or U4545 (N_4545,N_535,N_2059);
xor U4546 (N_4546,N_2191,N_2700);
xor U4547 (N_4547,N_2201,N_3000);
or U4548 (N_4548,N_1091,N_2605);
nor U4549 (N_4549,N_2242,N_1151);
and U4550 (N_4550,N_1586,N_2326);
nor U4551 (N_4551,N_1933,N_216);
xor U4552 (N_4552,N_3043,N_371);
xnor U4553 (N_4553,N_631,N_787);
or U4554 (N_4554,N_1607,N_2499);
or U4555 (N_4555,N_103,N_1993);
nand U4556 (N_4556,N_2182,N_456);
xor U4557 (N_4557,N_1900,N_1779);
xor U4558 (N_4558,N_791,N_203);
xor U4559 (N_4559,N_1635,N_2186);
xnor U4560 (N_4560,N_1459,N_2587);
or U4561 (N_4561,N_1681,N_1283);
xor U4562 (N_4562,N_1077,N_2836);
or U4563 (N_4563,N_1114,N_1784);
or U4564 (N_4564,N_1088,N_2738);
xnor U4565 (N_4565,N_1711,N_1190);
nor U4566 (N_4566,N_2808,N_2454);
nor U4567 (N_4567,N_130,N_612);
nor U4568 (N_4568,N_1930,N_953);
and U4569 (N_4569,N_1381,N_599);
nand U4570 (N_4570,N_484,N_2370);
nor U4571 (N_4571,N_380,N_434);
xnor U4572 (N_4572,N_1892,N_392);
nor U4573 (N_4573,N_952,N_64);
or U4574 (N_4574,N_2794,N_2825);
nand U4575 (N_4575,N_2067,N_2869);
xnor U4576 (N_4576,N_305,N_1461);
and U4577 (N_4577,N_13,N_744);
nand U4578 (N_4578,N_2382,N_1955);
nand U4579 (N_4579,N_1507,N_3082);
nor U4580 (N_4580,N_2543,N_2339);
xnor U4581 (N_4581,N_2078,N_2515);
xnor U4582 (N_4582,N_887,N_3019);
or U4583 (N_4583,N_1781,N_1448);
and U4584 (N_4584,N_893,N_796);
xnor U4585 (N_4585,N_538,N_2322);
nor U4586 (N_4586,N_2636,N_189);
xnor U4587 (N_4587,N_414,N_2055);
nor U4588 (N_4588,N_2189,N_840);
nand U4589 (N_4589,N_2408,N_98);
and U4590 (N_4590,N_924,N_2325);
nor U4591 (N_4591,N_2114,N_2478);
xor U4592 (N_4592,N_1815,N_2592);
xor U4593 (N_4593,N_912,N_2043);
xor U4594 (N_4594,N_1126,N_1272);
nand U4595 (N_4595,N_465,N_1575);
and U4596 (N_4596,N_2683,N_2516);
and U4597 (N_4597,N_2252,N_2514);
nand U4598 (N_4598,N_1419,N_526);
and U4599 (N_4599,N_2164,N_927);
nor U4600 (N_4600,N_1476,N_1421);
xor U4601 (N_4601,N_2103,N_1483);
and U4602 (N_4602,N_1472,N_2355);
xnor U4603 (N_4603,N_1449,N_2795);
and U4604 (N_4604,N_2834,N_1591);
nand U4605 (N_4605,N_1555,N_1324);
xnor U4606 (N_4606,N_1002,N_2298);
or U4607 (N_4607,N_1195,N_1929);
nor U4608 (N_4608,N_2988,N_1786);
nor U4609 (N_4609,N_378,N_659);
nor U4610 (N_4610,N_2217,N_773);
nand U4611 (N_4611,N_2641,N_499);
and U4612 (N_4612,N_1161,N_1569);
nand U4613 (N_4613,N_37,N_566);
nand U4614 (N_4614,N_508,N_2442);
or U4615 (N_4615,N_1842,N_1918);
xnor U4616 (N_4616,N_1731,N_1182);
xnor U4617 (N_4617,N_2154,N_395);
nor U4618 (N_4618,N_2348,N_3035);
xnor U4619 (N_4619,N_728,N_1210);
xor U4620 (N_4620,N_2109,N_1008);
nand U4621 (N_4621,N_1949,N_1482);
nor U4622 (N_4622,N_2119,N_1928);
nand U4623 (N_4623,N_2652,N_1991);
nor U4624 (N_4624,N_701,N_885);
nor U4625 (N_4625,N_1056,N_1689);
nor U4626 (N_4626,N_853,N_16);
nor U4627 (N_4627,N_1375,N_892);
and U4628 (N_4628,N_31,N_211);
and U4629 (N_4629,N_2208,N_2471);
nand U4630 (N_4630,N_1372,N_3069);
and U4631 (N_4631,N_898,N_2828);
and U4632 (N_4632,N_947,N_1405);
nor U4633 (N_4633,N_24,N_1809);
nor U4634 (N_4634,N_412,N_1759);
nor U4635 (N_4635,N_2456,N_1361);
and U4636 (N_4636,N_2448,N_863);
or U4637 (N_4637,N_2981,N_89);
nor U4638 (N_4638,N_1937,N_1156);
and U4639 (N_4639,N_3065,N_3051);
nand U4640 (N_4640,N_1309,N_462);
xnor U4641 (N_4641,N_2838,N_2247);
nor U4642 (N_4642,N_2237,N_1322);
xor U4643 (N_4643,N_188,N_906);
or U4644 (N_4644,N_34,N_1280);
or U4645 (N_4645,N_1855,N_1505);
nand U4646 (N_4646,N_1259,N_3016);
and U4647 (N_4647,N_423,N_1726);
nor U4648 (N_4648,N_1914,N_1494);
nor U4649 (N_4649,N_2312,N_196);
nand U4650 (N_4650,N_2480,N_313);
xnor U4651 (N_4651,N_2695,N_800);
and U4652 (N_4652,N_562,N_239);
and U4653 (N_4653,N_1471,N_2680);
or U4654 (N_4654,N_1066,N_2369);
nor U4655 (N_4655,N_113,N_516);
nand U4656 (N_4656,N_477,N_2221);
or U4657 (N_4657,N_1897,N_2721);
nor U4658 (N_4658,N_3029,N_865);
nor U4659 (N_4659,N_1241,N_2121);
xor U4660 (N_4660,N_1566,N_2207);
nand U4661 (N_4661,N_68,N_2272);
xor U4662 (N_4662,N_2375,N_970);
or U4663 (N_4663,N_2887,N_361);
nor U4664 (N_4664,N_2856,N_1872);
or U4665 (N_4665,N_2404,N_1157);
nor U4666 (N_4666,N_584,N_1684);
or U4667 (N_4667,N_2475,N_2727);
xor U4668 (N_4668,N_48,N_3100);
and U4669 (N_4669,N_2618,N_2202);
and U4670 (N_4670,N_420,N_2524);
nand U4671 (N_4671,N_2643,N_468);
or U4672 (N_4672,N_2013,N_2286);
or U4673 (N_4673,N_1547,N_1954);
nor U4674 (N_4674,N_2381,N_252);
nand U4675 (N_4675,N_497,N_880);
xor U4676 (N_4676,N_2385,N_575);
nand U4677 (N_4677,N_2354,N_1599);
nand U4678 (N_4678,N_2144,N_1636);
nor U4679 (N_4679,N_1848,N_1310);
nand U4680 (N_4680,N_1357,N_1893);
xor U4681 (N_4681,N_2356,N_2474);
nor U4682 (N_4682,N_2428,N_219);
nor U4683 (N_4683,N_2243,N_1323);
nor U4684 (N_4684,N_2853,N_1206);
xor U4685 (N_4685,N_2940,N_904);
xnor U4686 (N_4686,N_1550,N_3050);
nor U4687 (N_4687,N_1044,N_892);
nand U4688 (N_4688,N_3052,N_2766);
xnor U4689 (N_4689,N_1424,N_1992);
nor U4690 (N_4690,N_93,N_2325);
nand U4691 (N_4691,N_1704,N_2066);
nand U4692 (N_4692,N_150,N_1939);
or U4693 (N_4693,N_2142,N_3045);
xnor U4694 (N_4694,N_983,N_1783);
nor U4695 (N_4695,N_1298,N_2212);
or U4696 (N_4696,N_1283,N_795);
and U4697 (N_4697,N_623,N_823);
nand U4698 (N_4698,N_1939,N_2172);
and U4699 (N_4699,N_2286,N_485);
or U4700 (N_4700,N_1792,N_3080);
and U4701 (N_4701,N_2141,N_630);
nand U4702 (N_4702,N_387,N_2441);
nand U4703 (N_4703,N_2399,N_286);
or U4704 (N_4704,N_3035,N_1868);
and U4705 (N_4705,N_1638,N_523);
nor U4706 (N_4706,N_2208,N_1403);
or U4707 (N_4707,N_2648,N_1735);
xor U4708 (N_4708,N_2924,N_2582);
nand U4709 (N_4709,N_1863,N_2421);
xnor U4710 (N_4710,N_3075,N_2814);
nor U4711 (N_4711,N_2445,N_990);
xnor U4712 (N_4712,N_2231,N_3107);
nor U4713 (N_4713,N_856,N_3048);
nand U4714 (N_4714,N_1386,N_598);
xnor U4715 (N_4715,N_1227,N_907);
nand U4716 (N_4716,N_196,N_2204);
or U4717 (N_4717,N_731,N_1007);
and U4718 (N_4718,N_959,N_1744);
xnor U4719 (N_4719,N_299,N_914);
nand U4720 (N_4720,N_308,N_1837);
nor U4721 (N_4721,N_1463,N_1715);
or U4722 (N_4722,N_351,N_950);
nand U4723 (N_4723,N_2059,N_1934);
nor U4724 (N_4724,N_2011,N_442);
nand U4725 (N_4725,N_1845,N_2904);
nand U4726 (N_4726,N_3020,N_252);
or U4727 (N_4727,N_108,N_2303);
nor U4728 (N_4728,N_3052,N_2922);
nor U4729 (N_4729,N_1685,N_1666);
nor U4730 (N_4730,N_2703,N_2909);
and U4731 (N_4731,N_491,N_2861);
xor U4732 (N_4732,N_2830,N_1473);
or U4733 (N_4733,N_2800,N_687);
xor U4734 (N_4734,N_490,N_1819);
nand U4735 (N_4735,N_2328,N_1060);
and U4736 (N_4736,N_491,N_611);
or U4737 (N_4737,N_2464,N_287);
nor U4738 (N_4738,N_597,N_1017);
nand U4739 (N_4739,N_2016,N_1470);
and U4740 (N_4740,N_800,N_2056);
and U4741 (N_4741,N_1040,N_2364);
nor U4742 (N_4742,N_2497,N_3104);
nand U4743 (N_4743,N_598,N_235);
nand U4744 (N_4744,N_1104,N_902);
xnor U4745 (N_4745,N_2452,N_231);
and U4746 (N_4746,N_2274,N_846);
nand U4747 (N_4747,N_1016,N_2065);
nor U4748 (N_4748,N_368,N_1695);
and U4749 (N_4749,N_184,N_1669);
and U4750 (N_4750,N_2030,N_2549);
or U4751 (N_4751,N_1528,N_1051);
or U4752 (N_4752,N_1485,N_1790);
and U4753 (N_4753,N_1647,N_379);
xnor U4754 (N_4754,N_2866,N_208);
nor U4755 (N_4755,N_1461,N_1437);
nor U4756 (N_4756,N_1436,N_1933);
or U4757 (N_4757,N_368,N_2815);
nor U4758 (N_4758,N_1187,N_2741);
nor U4759 (N_4759,N_106,N_404);
nand U4760 (N_4760,N_2095,N_2324);
nand U4761 (N_4761,N_2931,N_2161);
xor U4762 (N_4762,N_2795,N_860);
or U4763 (N_4763,N_2727,N_689);
xor U4764 (N_4764,N_2856,N_2354);
and U4765 (N_4765,N_3093,N_2077);
and U4766 (N_4766,N_37,N_1853);
and U4767 (N_4767,N_2712,N_1635);
xnor U4768 (N_4768,N_933,N_318);
and U4769 (N_4769,N_887,N_674);
xnor U4770 (N_4770,N_2339,N_1248);
or U4771 (N_4771,N_1269,N_2128);
nand U4772 (N_4772,N_2681,N_490);
nor U4773 (N_4773,N_639,N_475);
and U4774 (N_4774,N_2868,N_2541);
xnor U4775 (N_4775,N_2713,N_1261);
nor U4776 (N_4776,N_905,N_3016);
and U4777 (N_4777,N_2090,N_2404);
and U4778 (N_4778,N_1596,N_1621);
xnor U4779 (N_4779,N_892,N_2929);
or U4780 (N_4780,N_344,N_2601);
or U4781 (N_4781,N_706,N_1986);
nor U4782 (N_4782,N_926,N_1492);
or U4783 (N_4783,N_2199,N_601);
or U4784 (N_4784,N_315,N_545);
or U4785 (N_4785,N_1228,N_2524);
nand U4786 (N_4786,N_2709,N_2082);
nand U4787 (N_4787,N_2531,N_2625);
nor U4788 (N_4788,N_880,N_946);
nand U4789 (N_4789,N_1967,N_964);
and U4790 (N_4790,N_2073,N_1138);
nand U4791 (N_4791,N_1935,N_132);
and U4792 (N_4792,N_2166,N_2724);
and U4793 (N_4793,N_1726,N_426);
xnor U4794 (N_4794,N_2133,N_2901);
or U4795 (N_4795,N_1977,N_1693);
nand U4796 (N_4796,N_129,N_658);
nand U4797 (N_4797,N_1035,N_541);
and U4798 (N_4798,N_2090,N_378);
xnor U4799 (N_4799,N_1583,N_931);
and U4800 (N_4800,N_2736,N_2696);
nor U4801 (N_4801,N_1592,N_2375);
nor U4802 (N_4802,N_526,N_417);
and U4803 (N_4803,N_89,N_824);
nand U4804 (N_4804,N_180,N_2456);
or U4805 (N_4805,N_2085,N_901);
nand U4806 (N_4806,N_2816,N_2829);
or U4807 (N_4807,N_814,N_2421);
and U4808 (N_4808,N_2754,N_1962);
xor U4809 (N_4809,N_265,N_966);
nand U4810 (N_4810,N_2636,N_1841);
xnor U4811 (N_4811,N_2639,N_1875);
xnor U4812 (N_4812,N_504,N_1204);
nand U4813 (N_4813,N_2847,N_1811);
nor U4814 (N_4814,N_2451,N_2368);
nor U4815 (N_4815,N_2273,N_516);
and U4816 (N_4816,N_2452,N_2776);
nor U4817 (N_4817,N_2286,N_1269);
nor U4818 (N_4818,N_2571,N_2542);
or U4819 (N_4819,N_122,N_505);
nand U4820 (N_4820,N_2857,N_1582);
xnor U4821 (N_4821,N_2306,N_1218);
and U4822 (N_4822,N_2477,N_1649);
xnor U4823 (N_4823,N_1673,N_2648);
nand U4824 (N_4824,N_2781,N_136);
and U4825 (N_4825,N_1780,N_819);
and U4826 (N_4826,N_2342,N_3023);
nand U4827 (N_4827,N_724,N_1578);
and U4828 (N_4828,N_2882,N_1562);
nand U4829 (N_4829,N_368,N_1925);
nor U4830 (N_4830,N_2665,N_2162);
xor U4831 (N_4831,N_1211,N_2262);
xor U4832 (N_4832,N_1182,N_1415);
and U4833 (N_4833,N_338,N_1417);
nor U4834 (N_4834,N_1142,N_1328);
xor U4835 (N_4835,N_2190,N_1534);
nor U4836 (N_4836,N_3111,N_717);
and U4837 (N_4837,N_1063,N_113);
nor U4838 (N_4838,N_1690,N_138);
nand U4839 (N_4839,N_2539,N_2689);
xor U4840 (N_4840,N_1068,N_3117);
nand U4841 (N_4841,N_2287,N_421);
xor U4842 (N_4842,N_231,N_404);
or U4843 (N_4843,N_3078,N_941);
xor U4844 (N_4844,N_192,N_2382);
and U4845 (N_4845,N_1255,N_207);
nand U4846 (N_4846,N_2611,N_2306);
xnor U4847 (N_4847,N_627,N_428);
nand U4848 (N_4848,N_2197,N_1402);
xnor U4849 (N_4849,N_1414,N_639);
or U4850 (N_4850,N_2202,N_343);
nor U4851 (N_4851,N_1705,N_1435);
and U4852 (N_4852,N_41,N_2140);
xor U4853 (N_4853,N_1536,N_2225);
nor U4854 (N_4854,N_440,N_2860);
nor U4855 (N_4855,N_413,N_2854);
and U4856 (N_4856,N_1709,N_902);
nand U4857 (N_4857,N_2418,N_360);
or U4858 (N_4858,N_2283,N_2368);
nand U4859 (N_4859,N_2495,N_762);
nor U4860 (N_4860,N_785,N_1063);
nand U4861 (N_4861,N_2252,N_3100);
xnor U4862 (N_4862,N_2974,N_3123);
xor U4863 (N_4863,N_2038,N_385);
nor U4864 (N_4864,N_2035,N_2371);
xnor U4865 (N_4865,N_2375,N_1860);
or U4866 (N_4866,N_1813,N_3081);
and U4867 (N_4867,N_7,N_359);
nor U4868 (N_4868,N_590,N_845);
xor U4869 (N_4869,N_994,N_2199);
xnor U4870 (N_4870,N_1567,N_409);
nand U4871 (N_4871,N_451,N_2634);
nor U4872 (N_4872,N_2550,N_1405);
or U4873 (N_4873,N_2788,N_104);
nand U4874 (N_4874,N_15,N_747);
nor U4875 (N_4875,N_2628,N_923);
xor U4876 (N_4876,N_2965,N_870);
or U4877 (N_4877,N_1641,N_184);
or U4878 (N_4878,N_2422,N_1089);
nand U4879 (N_4879,N_945,N_2821);
nor U4880 (N_4880,N_1956,N_261);
xnor U4881 (N_4881,N_3091,N_1601);
xnor U4882 (N_4882,N_2957,N_2184);
and U4883 (N_4883,N_1359,N_1334);
nand U4884 (N_4884,N_2307,N_2551);
nor U4885 (N_4885,N_2314,N_1995);
nor U4886 (N_4886,N_511,N_1689);
xor U4887 (N_4887,N_1426,N_1497);
nor U4888 (N_4888,N_689,N_2793);
xor U4889 (N_4889,N_2670,N_3044);
xor U4890 (N_4890,N_2855,N_1573);
nor U4891 (N_4891,N_1994,N_3001);
xor U4892 (N_4892,N_564,N_1114);
and U4893 (N_4893,N_2964,N_1417);
nand U4894 (N_4894,N_1701,N_24);
or U4895 (N_4895,N_1653,N_406);
and U4896 (N_4896,N_2817,N_756);
xor U4897 (N_4897,N_2103,N_468);
and U4898 (N_4898,N_2024,N_1421);
or U4899 (N_4899,N_1371,N_935);
or U4900 (N_4900,N_2472,N_619);
nor U4901 (N_4901,N_5,N_1326);
nand U4902 (N_4902,N_2214,N_612);
nand U4903 (N_4903,N_2913,N_1526);
xnor U4904 (N_4904,N_2643,N_88);
nand U4905 (N_4905,N_1647,N_1035);
xor U4906 (N_4906,N_3012,N_87);
nor U4907 (N_4907,N_2388,N_1340);
nor U4908 (N_4908,N_338,N_638);
and U4909 (N_4909,N_2777,N_2404);
and U4910 (N_4910,N_296,N_2570);
nand U4911 (N_4911,N_962,N_810);
or U4912 (N_4912,N_2308,N_1725);
and U4913 (N_4913,N_391,N_2823);
and U4914 (N_4914,N_2234,N_3093);
nand U4915 (N_4915,N_1859,N_2832);
nand U4916 (N_4916,N_1107,N_2411);
and U4917 (N_4917,N_489,N_567);
and U4918 (N_4918,N_1795,N_2967);
or U4919 (N_4919,N_1705,N_2876);
and U4920 (N_4920,N_2597,N_925);
xor U4921 (N_4921,N_695,N_678);
nor U4922 (N_4922,N_2603,N_2046);
xnor U4923 (N_4923,N_2199,N_753);
xor U4924 (N_4924,N_884,N_268);
and U4925 (N_4925,N_180,N_301);
or U4926 (N_4926,N_1943,N_1128);
and U4927 (N_4927,N_2265,N_2811);
nand U4928 (N_4928,N_3013,N_208);
nand U4929 (N_4929,N_1385,N_1271);
xnor U4930 (N_4930,N_2794,N_1901);
nor U4931 (N_4931,N_450,N_2203);
xor U4932 (N_4932,N_216,N_2034);
nand U4933 (N_4933,N_1405,N_2709);
or U4934 (N_4934,N_2112,N_250);
or U4935 (N_4935,N_1170,N_2466);
nand U4936 (N_4936,N_2590,N_2227);
or U4937 (N_4937,N_2206,N_710);
or U4938 (N_4938,N_2924,N_868);
nand U4939 (N_4939,N_1753,N_2784);
and U4940 (N_4940,N_2557,N_1455);
xnor U4941 (N_4941,N_1103,N_713);
or U4942 (N_4942,N_2819,N_1265);
nand U4943 (N_4943,N_596,N_1678);
nor U4944 (N_4944,N_1960,N_2378);
nand U4945 (N_4945,N_1667,N_216);
xor U4946 (N_4946,N_628,N_1515);
xnor U4947 (N_4947,N_1835,N_2230);
or U4948 (N_4948,N_2870,N_857);
nor U4949 (N_4949,N_2394,N_2821);
or U4950 (N_4950,N_1930,N_2212);
nand U4951 (N_4951,N_1087,N_1311);
and U4952 (N_4952,N_376,N_593);
nor U4953 (N_4953,N_1585,N_222);
nor U4954 (N_4954,N_1643,N_2045);
or U4955 (N_4955,N_1786,N_2599);
and U4956 (N_4956,N_797,N_1038);
nor U4957 (N_4957,N_1571,N_1882);
xor U4958 (N_4958,N_2146,N_1193);
xor U4959 (N_4959,N_808,N_2851);
nor U4960 (N_4960,N_1723,N_886);
or U4961 (N_4961,N_1950,N_2432);
and U4962 (N_4962,N_2592,N_741);
nor U4963 (N_4963,N_2012,N_1900);
nand U4964 (N_4964,N_1124,N_1072);
or U4965 (N_4965,N_2547,N_433);
nand U4966 (N_4966,N_2853,N_2663);
and U4967 (N_4967,N_1119,N_2091);
and U4968 (N_4968,N_2277,N_1940);
nor U4969 (N_4969,N_1256,N_3052);
nand U4970 (N_4970,N_2640,N_22);
nand U4971 (N_4971,N_1505,N_1122);
nor U4972 (N_4972,N_1892,N_2536);
nor U4973 (N_4973,N_2577,N_1193);
or U4974 (N_4974,N_2410,N_2170);
xor U4975 (N_4975,N_2267,N_1488);
and U4976 (N_4976,N_979,N_543);
and U4977 (N_4977,N_1989,N_1311);
and U4978 (N_4978,N_142,N_145);
and U4979 (N_4979,N_2641,N_2465);
xor U4980 (N_4980,N_160,N_1810);
nor U4981 (N_4981,N_2046,N_1713);
or U4982 (N_4982,N_2794,N_933);
nand U4983 (N_4983,N_1472,N_2918);
nor U4984 (N_4984,N_2974,N_2605);
and U4985 (N_4985,N_647,N_88);
or U4986 (N_4986,N_902,N_1947);
xnor U4987 (N_4987,N_2161,N_586);
and U4988 (N_4988,N_1590,N_587);
or U4989 (N_4989,N_2788,N_1692);
and U4990 (N_4990,N_655,N_799);
or U4991 (N_4991,N_2464,N_1561);
xor U4992 (N_4992,N_1162,N_2100);
and U4993 (N_4993,N_887,N_2503);
and U4994 (N_4994,N_914,N_976);
nand U4995 (N_4995,N_65,N_160);
and U4996 (N_4996,N_2845,N_3094);
and U4997 (N_4997,N_647,N_1883);
xnor U4998 (N_4998,N_976,N_2471);
and U4999 (N_4999,N_2788,N_279);
nand U5000 (N_5000,N_2791,N_2493);
or U5001 (N_5001,N_1249,N_2295);
nor U5002 (N_5002,N_2029,N_1178);
nor U5003 (N_5003,N_2226,N_353);
nor U5004 (N_5004,N_2314,N_2834);
xnor U5005 (N_5005,N_149,N_2657);
nand U5006 (N_5006,N_3112,N_1820);
nand U5007 (N_5007,N_1917,N_498);
xor U5008 (N_5008,N_2474,N_1833);
nor U5009 (N_5009,N_895,N_2556);
or U5010 (N_5010,N_228,N_2196);
or U5011 (N_5011,N_2323,N_2776);
and U5012 (N_5012,N_2531,N_1090);
and U5013 (N_5013,N_447,N_2378);
nor U5014 (N_5014,N_2574,N_2914);
xnor U5015 (N_5015,N_1585,N_1014);
nand U5016 (N_5016,N_1652,N_948);
and U5017 (N_5017,N_3037,N_366);
nand U5018 (N_5018,N_2934,N_894);
and U5019 (N_5019,N_930,N_395);
xnor U5020 (N_5020,N_2572,N_1017);
nor U5021 (N_5021,N_1138,N_6);
or U5022 (N_5022,N_1006,N_2772);
and U5023 (N_5023,N_1370,N_2943);
and U5024 (N_5024,N_2463,N_23);
nor U5025 (N_5025,N_1079,N_2109);
and U5026 (N_5026,N_956,N_430);
nand U5027 (N_5027,N_1443,N_1693);
xor U5028 (N_5028,N_2746,N_625);
nor U5029 (N_5029,N_270,N_1800);
and U5030 (N_5030,N_2077,N_1558);
nor U5031 (N_5031,N_841,N_2627);
or U5032 (N_5032,N_1687,N_2839);
nor U5033 (N_5033,N_3007,N_2936);
or U5034 (N_5034,N_1274,N_396);
xor U5035 (N_5035,N_879,N_801);
or U5036 (N_5036,N_2487,N_2071);
and U5037 (N_5037,N_259,N_1792);
or U5038 (N_5038,N_527,N_2826);
and U5039 (N_5039,N_137,N_698);
nand U5040 (N_5040,N_68,N_2676);
nor U5041 (N_5041,N_1181,N_1036);
or U5042 (N_5042,N_1165,N_2004);
nand U5043 (N_5043,N_1776,N_2837);
nor U5044 (N_5044,N_2215,N_1324);
or U5045 (N_5045,N_348,N_1188);
nand U5046 (N_5046,N_202,N_638);
xor U5047 (N_5047,N_645,N_1211);
and U5048 (N_5048,N_1594,N_959);
nand U5049 (N_5049,N_1461,N_1910);
xnor U5050 (N_5050,N_1551,N_1915);
nor U5051 (N_5051,N_652,N_1780);
and U5052 (N_5052,N_2728,N_278);
or U5053 (N_5053,N_2257,N_182);
xor U5054 (N_5054,N_1713,N_460);
xor U5055 (N_5055,N_2515,N_911);
xnor U5056 (N_5056,N_1983,N_73);
and U5057 (N_5057,N_1125,N_2941);
nor U5058 (N_5058,N_1014,N_2032);
or U5059 (N_5059,N_1438,N_20);
xor U5060 (N_5060,N_1638,N_1621);
or U5061 (N_5061,N_2347,N_793);
nand U5062 (N_5062,N_2941,N_1208);
and U5063 (N_5063,N_1868,N_1899);
xor U5064 (N_5064,N_1597,N_2256);
and U5065 (N_5065,N_222,N_1328);
nor U5066 (N_5066,N_3088,N_225);
or U5067 (N_5067,N_2006,N_2827);
nor U5068 (N_5068,N_1999,N_1584);
and U5069 (N_5069,N_1529,N_2160);
xnor U5070 (N_5070,N_1906,N_1627);
nand U5071 (N_5071,N_203,N_3098);
and U5072 (N_5072,N_1641,N_2393);
nand U5073 (N_5073,N_1626,N_2764);
nand U5074 (N_5074,N_3049,N_1033);
nand U5075 (N_5075,N_663,N_2279);
and U5076 (N_5076,N_2218,N_888);
xor U5077 (N_5077,N_1231,N_2078);
or U5078 (N_5078,N_1528,N_91);
and U5079 (N_5079,N_2439,N_1287);
and U5080 (N_5080,N_2945,N_576);
or U5081 (N_5081,N_2817,N_2586);
nor U5082 (N_5082,N_2693,N_2718);
xnor U5083 (N_5083,N_872,N_1614);
xnor U5084 (N_5084,N_1383,N_743);
and U5085 (N_5085,N_153,N_1026);
or U5086 (N_5086,N_2874,N_521);
and U5087 (N_5087,N_2548,N_3009);
and U5088 (N_5088,N_653,N_2920);
nand U5089 (N_5089,N_923,N_1610);
or U5090 (N_5090,N_2202,N_761);
and U5091 (N_5091,N_1748,N_2009);
nand U5092 (N_5092,N_389,N_1044);
or U5093 (N_5093,N_1251,N_1766);
and U5094 (N_5094,N_945,N_1791);
nor U5095 (N_5095,N_1877,N_2421);
nand U5096 (N_5096,N_1382,N_2068);
or U5097 (N_5097,N_1030,N_1241);
and U5098 (N_5098,N_1823,N_1068);
or U5099 (N_5099,N_2937,N_2808);
nand U5100 (N_5100,N_2766,N_2335);
nand U5101 (N_5101,N_1727,N_1844);
and U5102 (N_5102,N_1307,N_1122);
nor U5103 (N_5103,N_2396,N_2816);
nand U5104 (N_5104,N_1074,N_162);
nand U5105 (N_5105,N_614,N_2523);
nor U5106 (N_5106,N_1160,N_1021);
nor U5107 (N_5107,N_2348,N_956);
nand U5108 (N_5108,N_926,N_1778);
nor U5109 (N_5109,N_2044,N_1336);
nand U5110 (N_5110,N_2762,N_2746);
nand U5111 (N_5111,N_249,N_2780);
xnor U5112 (N_5112,N_298,N_2327);
xor U5113 (N_5113,N_496,N_1928);
and U5114 (N_5114,N_578,N_2992);
nand U5115 (N_5115,N_1549,N_1330);
and U5116 (N_5116,N_2379,N_549);
and U5117 (N_5117,N_1019,N_1189);
nor U5118 (N_5118,N_2683,N_2666);
and U5119 (N_5119,N_2569,N_238);
and U5120 (N_5120,N_134,N_934);
xnor U5121 (N_5121,N_1436,N_30);
nor U5122 (N_5122,N_1545,N_1844);
or U5123 (N_5123,N_596,N_1562);
nor U5124 (N_5124,N_2945,N_1818);
and U5125 (N_5125,N_733,N_1188);
and U5126 (N_5126,N_3105,N_2432);
nand U5127 (N_5127,N_3113,N_31);
nand U5128 (N_5128,N_1577,N_1498);
xor U5129 (N_5129,N_2420,N_3115);
xnor U5130 (N_5130,N_2430,N_1413);
or U5131 (N_5131,N_1829,N_1257);
xor U5132 (N_5132,N_2182,N_1471);
xnor U5133 (N_5133,N_1543,N_57);
xnor U5134 (N_5134,N_1661,N_1899);
xor U5135 (N_5135,N_3060,N_2554);
xnor U5136 (N_5136,N_1194,N_1398);
nor U5137 (N_5137,N_1436,N_2824);
nand U5138 (N_5138,N_1720,N_1915);
nand U5139 (N_5139,N_2550,N_3052);
xnor U5140 (N_5140,N_186,N_555);
nand U5141 (N_5141,N_696,N_1164);
or U5142 (N_5142,N_2490,N_1029);
xnor U5143 (N_5143,N_2738,N_2051);
xor U5144 (N_5144,N_1105,N_1418);
and U5145 (N_5145,N_1940,N_493);
nand U5146 (N_5146,N_2342,N_1784);
nand U5147 (N_5147,N_814,N_1241);
and U5148 (N_5148,N_1942,N_474);
xnor U5149 (N_5149,N_2068,N_209);
xor U5150 (N_5150,N_2767,N_2015);
and U5151 (N_5151,N_2356,N_739);
or U5152 (N_5152,N_25,N_1436);
and U5153 (N_5153,N_95,N_2985);
or U5154 (N_5154,N_897,N_2244);
nor U5155 (N_5155,N_1566,N_2550);
nand U5156 (N_5156,N_1929,N_910);
or U5157 (N_5157,N_2319,N_269);
nor U5158 (N_5158,N_3025,N_2637);
nor U5159 (N_5159,N_841,N_2424);
nand U5160 (N_5160,N_861,N_2720);
xnor U5161 (N_5161,N_2605,N_900);
nand U5162 (N_5162,N_1252,N_51);
and U5163 (N_5163,N_898,N_3081);
xor U5164 (N_5164,N_1799,N_1708);
xnor U5165 (N_5165,N_2945,N_368);
or U5166 (N_5166,N_888,N_2082);
and U5167 (N_5167,N_1654,N_2283);
nand U5168 (N_5168,N_916,N_598);
nor U5169 (N_5169,N_2015,N_222);
or U5170 (N_5170,N_257,N_215);
nor U5171 (N_5171,N_1073,N_264);
nor U5172 (N_5172,N_2505,N_1183);
and U5173 (N_5173,N_498,N_581);
nand U5174 (N_5174,N_2071,N_2705);
and U5175 (N_5175,N_611,N_2371);
or U5176 (N_5176,N_37,N_3096);
xnor U5177 (N_5177,N_186,N_2935);
xor U5178 (N_5178,N_2641,N_1514);
nor U5179 (N_5179,N_2332,N_2232);
or U5180 (N_5180,N_2485,N_502);
or U5181 (N_5181,N_2005,N_2995);
xor U5182 (N_5182,N_1063,N_1410);
or U5183 (N_5183,N_1808,N_1141);
and U5184 (N_5184,N_1069,N_2634);
nand U5185 (N_5185,N_1007,N_1464);
nor U5186 (N_5186,N_3073,N_2440);
nor U5187 (N_5187,N_2126,N_2777);
or U5188 (N_5188,N_1736,N_2232);
xor U5189 (N_5189,N_1498,N_1461);
nor U5190 (N_5190,N_2640,N_1705);
or U5191 (N_5191,N_2366,N_1370);
or U5192 (N_5192,N_1460,N_834);
xor U5193 (N_5193,N_998,N_1972);
and U5194 (N_5194,N_2696,N_1435);
xor U5195 (N_5195,N_583,N_2503);
xor U5196 (N_5196,N_3007,N_953);
xnor U5197 (N_5197,N_366,N_683);
nor U5198 (N_5198,N_2499,N_427);
or U5199 (N_5199,N_429,N_2127);
or U5200 (N_5200,N_728,N_2369);
nand U5201 (N_5201,N_3051,N_2807);
xnor U5202 (N_5202,N_420,N_711);
nand U5203 (N_5203,N_2971,N_2802);
nor U5204 (N_5204,N_1866,N_591);
nor U5205 (N_5205,N_1333,N_765);
or U5206 (N_5206,N_2969,N_2598);
xor U5207 (N_5207,N_81,N_2638);
or U5208 (N_5208,N_1659,N_2615);
xor U5209 (N_5209,N_323,N_1887);
and U5210 (N_5210,N_1457,N_1489);
or U5211 (N_5211,N_2465,N_2768);
or U5212 (N_5212,N_648,N_1018);
and U5213 (N_5213,N_1643,N_293);
nor U5214 (N_5214,N_661,N_2561);
nor U5215 (N_5215,N_458,N_336);
nor U5216 (N_5216,N_597,N_1413);
or U5217 (N_5217,N_2212,N_1184);
nand U5218 (N_5218,N_847,N_2707);
xnor U5219 (N_5219,N_501,N_1601);
and U5220 (N_5220,N_1935,N_2219);
nor U5221 (N_5221,N_2015,N_3082);
and U5222 (N_5222,N_2432,N_3033);
nor U5223 (N_5223,N_298,N_2025);
or U5224 (N_5224,N_592,N_1228);
nor U5225 (N_5225,N_2227,N_2718);
and U5226 (N_5226,N_777,N_1295);
nor U5227 (N_5227,N_2723,N_2214);
nor U5228 (N_5228,N_348,N_1350);
xnor U5229 (N_5229,N_1703,N_1546);
nor U5230 (N_5230,N_1433,N_365);
and U5231 (N_5231,N_2401,N_2649);
xor U5232 (N_5232,N_3033,N_2535);
nor U5233 (N_5233,N_1732,N_880);
or U5234 (N_5234,N_1956,N_26);
xnor U5235 (N_5235,N_2092,N_2611);
nor U5236 (N_5236,N_1115,N_2994);
nand U5237 (N_5237,N_626,N_662);
nand U5238 (N_5238,N_13,N_2622);
nand U5239 (N_5239,N_1232,N_1118);
xnor U5240 (N_5240,N_1749,N_906);
or U5241 (N_5241,N_2849,N_637);
nor U5242 (N_5242,N_145,N_1505);
or U5243 (N_5243,N_2990,N_564);
nor U5244 (N_5244,N_1577,N_2053);
and U5245 (N_5245,N_2981,N_1549);
or U5246 (N_5246,N_2395,N_2786);
and U5247 (N_5247,N_922,N_1393);
nand U5248 (N_5248,N_1981,N_1948);
nand U5249 (N_5249,N_84,N_1081);
nor U5250 (N_5250,N_2442,N_3118);
nand U5251 (N_5251,N_776,N_2086);
nand U5252 (N_5252,N_2864,N_841);
xor U5253 (N_5253,N_3070,N_1635);
nand U5254 (N_5254,N_2173,N_2961);
nand U5255 (N_5255,N_2914,N_2189);
nor U5256 (N_5256,N_2592,N_1013);
nand U5257 (N_5257,N_1011,N_66);
nand U5258 (N_5258,N_1622,N_2893);
and U5259 (N_5259,N_462,N_2987);
and U5260 (N_5260,N_242,N_812);
nand U5261 (N_5261,N_1876,N_1998);
and U5262 (N_5262,N_2977,N_871);
xnor U5263 (N_5263,N_1152,N_2254);
or U5264 (N_5264,N_431,N_2202);
or U5265 (N_5265,N_12,N_1206);
nor U5266 (N_5266,N_2087,N_393);
or U5267 (N_5267,N_1649,N_946);
xor U5268 (N_5268,N_1726,N_2517);
xor U5269 (N_5269,N_1890,N_2370);
nor U5270 (N_5270,N_1700,N_1136);
xnor U5271 (N_5271,N_221,N_1702);
nor U5272 (N_5272,N_1164,N_1840);
or U5273 (N_5273,N_1699,N_988);
nor U5274 (N_5274,N_566,N_764);
xnor U5275 (N_5275,N_555,N_2286);
and U5276 (N_5276,N_1260,N_2568);
xnor U5277 (N_5277,N_100,N_835);
and U5278 (N_5278,N_270,N_2334);
nand U5279 (N_5279,N_1898,N_1435);
xnor U5280 (N_5280,N_1579,N_1862);
nor U5281 (N_5281,N_1952,N_1003);
nor U5282 (N_5282,N_1975,N_2187);
nand U5283 (N_5283,N_2472,N_472);
or U5284 (N_5284,N_532,N_2178);
or U5285 (N_5285,N_413,N_474);
nand U5286 (N_5286,N_580,N_2486);
nand U5287 (N_5287,N_2175,N_2438);
nor U5288 (N_5288,N_62,N_268);
xnor U5289 (N_5289,N_2305,N_385);
nand U5290 (N_5290,N_3124,N_158);
and U5291 (N_5291,N_2784,N_2725);
xor U5292 (N_5292,N_1071,N_213);
and U5293 (N_5293,N_2642,N_537);
or U5294 (N_5294,N_2790,N_3108);
or U5295 (N_5295,N_2952,N_730);
and U5296 (N_5296,N_1284,N_714);
nand U5297 (N_5297,N_1748,N_2997);
and U5298 (N_5298,N_2784,N_3101);
and U5299 (N_5299,N_200,N_1795);
nand U5300 (N_5300,N_493,N_1198);
nor U5301 (N_5301,N_2454,N_2624);
nand U5302 (N_5302,N_2939,N_1232);
xor U5303 (N_5303,N_189,N_3080);
nand U5304 (N_5304,N_1552,N_724);
or U5305 (N_5305,N_1559,N_1913);
and U5306 (N_5306,N_876,N_2698);
xor U5307 (N_5307,N_1494,N_1007);
xnor U5308 (N_5308,N_1607,N_878);
nor U5309 (N_5309,N_2105,N_670);
nor U5310 (N_5310,N_133,N_2498);
xnor U5311 (N_5311,N_2696,N_1268);
xor U5312 (N_5312,N_1159,N_1068);
and U5313 (N_5313,N_1614,N_1708);
xnor U5314 (N_5314,N_240,N_935);
nand U5315 (N_5315,N_1380,N_2780);
nor U5316 (N_5316,N_134,N_2100);
or U5317 (N_5317,N_59,N_1683);
or U5318 (N_5318,N_1850,N_2789);
nor U5319 (N_5319,N_915,N_612);
nand U5320 (N_5320,N_2521,N_1760);
xor U5321 (N_5321,N_869,N_1794);
or U5322 (N_5322,N_1799,N_1131);
nand U5323 (N_5323,N_1619,N_1852);
or U5324 (N_5324,N_2662,N_2408);
nand U5325 (N_5325,N_1163,N_1160);
nor U5326 (N_5326,N_2478,N_2210);
xnor U5327 (N_5327,N_2193,N_1443);
nor U5328 (N_5328,N_920,N_1402);
nor U5329 (N_5329,N_951,N_773);
and U5330 (N_5330,N_2031,N_360);
nor U5331 (N_5331,N_838,N_1362);
and U5332 (N_5332,N_2058,N_1255);
and U5333 (N_5333,N_1543,N_3090);
or U5334 (N_5334,N_2491,N_2892);
xor U5335 (N_5335,N_15,N_2559);
xnor U5336 (N_5336,N_2116,N_2296);
and U5337 (N_5337,N_2929,N_2948);
xor U5338 (N_5338,N_2821,N_2777);
nand U5339 (N_5339,N_2842,N_1987);
nor U5340 (N_5340,N_291,N_1618);
nand U5341 (N_5341,N_1255,N_573);
nor U5342 (N_5342,N_445,N_1035);
nor U5343 (N_5343,N_378,N_1916);
and U5344 (N_5344,N_2133,N_409);
or U5345 (N_5345,N_2742,N_1224);
and U5346 (N_5346,N_287,N_2400);
xnor U5347 (N_5347,N_1842,N_145);
and U5348 (N_5348,N_2032,N_1582);
xor U5349 (N_5349,N_316,N_788);
and U5350 (N_5350,N_981,N_1157);
and U5351 (N_5351,N_2887,N_45);
nor U5352 (N_5352,N_1063,N_1974);
nand U5353 (N_5353,N_2049,N_325);
nand U5354 (N_5354,N_1643,N_1090);
nand U5355 (N_5355,N_1367,N_756);
xor U5356 (N_5356,N_2853,N_2596);
and U5357 (N_5357,N_311,N_3027);
nand U5358 (N_5358,N_1408,N_3044);
or U5359 (N_5359,N_1683,N_1005);
nor U5360 (N_5360,N_1839,N_1761);
nor U5361 (N_5361,N_1493,N_1628);
or U5362 (N_5362,N_1880,N_580);
or U5363 (N_5363,N_1322,N_1776);
nand U5364 (N_5364,N_2124,N_902);
nor U5365 (N_5365,N_1936,N_1651);
xnor U5366 (N_5366,N_937,N_332);
or U5367 (N_5367,N_1335,N_1935);
nand U5368 (N_5368,N_922,N_3124);
or U5369 (N_5369,N_3018,N_1483);
nor U5370 (N_5370,N_1580,N_161);
nor U5371 (N_5371,N_2719,N_104);
or U5372 (N_5372,N_639,N_2578);
or U5373 (N_5373,N_3007,N_1245);
or U5374 (N_5374,N_1578,N_731);
and U5375 (N_5375,N_2861,N_2929);
nand U5376 (N_5376,N_2701,N_2319);
xnor U5377 (N_5377,N_2571,N_2488);
nor U5378 (N_5378,N_793,N_1539);
or U5379 (N_5379,N_2234,N_960);
or U5380 (N_5380,N_105,N_1217);
xnor U5381 (N_5381,N_824,N_1092);
or U5382 (N_5382,N_943,N_2517);
xor U5383 (N_5383,N_2830,N_2392);
xnor U5384 (N_5384,N_2210,N_1505);
or U5385 (N_5385,N_1616,N_2319);
or U5386 (N_5386,N_807,N_1911);
xor U5387 (N_5387,N_1887,N_844);
or U5388 (N_5388,N_3014,N_209);
nand U5389 (N_5389,N_544,N_1827);
nand U5390 (N_5390,N_551,N_2140);
and U5391 (N_5391,N_140,N_1170);
nor U5392 (N_5392,N_2885,N_2526);
or U5393 (N_5393,N_2519,N_2429);
xnor U5394 (N_5394,N_2589,N_1133);
and U5395 (N_5395,N_2582,N_1667);
or U5396 (N_5396,N_334,N_2077);
and U5397 (N_5397,N_3061,N_1653);
nor U5398 (N_5398,N_618,N_2998);
and U5399 (N_5399,N_1123,N_781);
or U5400 (N_5400,N_134,N_2643);
nor U5401 (N_5401,N_607,N_1063);
nand U5402 (N_5402,N_1398,N_607);
nand U5403 (N_5403,N_2118,N_1004);
and U5404 (N_5404,N_2822,N_716);
nand U5405 (N_5405,N_1763,N_2998);
or U5406 (N_5406,N_2946,N_2871);
xor U5407 (N_5407,N_408,N_1370);
xor U5408 (N_5408,N_1023,N_1241);
nand U5409 (N_5409,N_648,N_1697);
nor U5410 (N_5410,N_2101,N_2410);
or U5411 (N_5411,N_1114,N_1049);
or U5412 (N_5412,N_1739,N_1201);
or U5413 (N_5413,N_1940,N_2183);
or U5414 (N_5414,N_682,N_389);
nor U5415 (N_5415,N_2828,N_329);
xnor U5416 (N_5416,N_2125,N_2141);
nand U5417 (N_5417,N_907,N_2652);
or U5418 (N_5418,N_84,N_893);
nand U5419 (N_5419,N_1866,N_518);
nand U5420 (N_5420,N_2651,N_1587);
nand U5421 (N_5421,N_1537,N_1845);
nand U5422 (N_5422,N_1249,N_759);
or U5423 (N_5423,N_298,N_2093);
xor U5424 (N_5424,N_2351,N_2962);
and U5425 (N_5425,N_2232,N_835);
and U5426 (N_5426,N_3121,N_306);
nand U5427 (N_5427,N_1992,N_814);
nor U5428 (N_5428,N_49,N_2045);
and U5429 (N_5429,N_2925,N_2322);
or U5430 (N_5430,N_2532,N_2681);
and U5431 (N_5431,N_3083,N_2901);
or U5432 (N_5432,N_2349,N_68);
nor U5433 (N_5433,N_2607,N_419);
nor U5434 (N_5434,N_158,N_2503);
and U5435 (N_5435,N_3113,N_2741);
nor U5436 (N_5436,N_2721,N_2193);
or U5437 (N_5437,N_2149,N_378);
xor U5438 (N_5438,N_2594,N_2287);
nand U5439 (N_5439,N_360,N_2648);
nor U5440 (N_5440,N_711,N_1803);
xor U5441 (N_5441,N_1779,N_537);
xor U5442 (N_5442,N_2351,N_853);
or U5443 (N_5443,N_3011,N_1844);
nor U5444 (N_5444,N_1397,N_257);
nor U5445 (N_5445,N_2823,N_2210);
nand U5446 (N_5446,N_1285,N_647);
nor U5447 (N_5447,N_234,N_1575);
nor U5448 (N_5448,N_1695,N_1843);
nor U5449 (N_5449,N_3023,N_2014);
or U5450 (N_5450,N_1471,N_693);
xor U5451 (N_5451,N_2200,N_587);
xnor U5452 (N_5452,N_1746,N_638);
and U5453 (N_5453,N_603,N_1817);
nand U5454 (N_5454,N_2754,N_547);
or U5455 (N_5455,N_1474,N_1693);
or U5456 (N_5456,N_1340,N_1928);
xor U5457 (N_5457,N_2488,N_2896);
xnor U5458 (N_5458,N_32,N_1673);
and U5459 (N_5459,N_472,N_2737);
and U5460 (N_5460,N_3029,N_175);
xnor U5461 (N_5461,N_62,N_2746);
and U5462 (N_5462,N_2870,N_1777);
nor U5463 (N_5463,N_2035,N_2950);
nand U5464 (N_5464,N_3036,N_464);
xor U5465 (N_5465,N_2853,N_2966);
xnor U5466 (N_5466,N_2973,N_2529);
xor U5467 (N_5467,N_1921,N_785);
nor U5468 (N_5468,N_40,N_2575);
xor U5469 (N_5469,N_2097,N_2106);
xor U5470 (N_5470,N_1157,N_1432);
nor U5471 (N_5471,N_374,N_1309);
xor U5472 (N_5472,N_111,N_1957);
and U5473 (N_5473,N_2697,N_405);
xnor U5474 (N_5474,N_1743,N_559);
nand U5475 (N_5475,N_393,N_1348);
xor U5476 (N_5476,N_1987,N_1066);
and U5477 (N_5477,N_2788,N_3068);
xor U5478 (N_5478,N_365,N_2862);
and U5479 (N_5479,N_1871,N_1924);
or U5480 (N_5480,N_132,N_2150);
xor U5481 (N_5481,N_270,N_1000);
nand U5482 (N_5482,N_2620,N_2411);
nor U5483 (N_5483,N_1377,N_622);
or U5484 (N_5484,N_3019,N_2578);
xor U5485 (N_5485,N_2714,N_517);
nand U5486 (N_5486,N_2598,N_704);
or U5487 (N_5487,N_2168,N_1007);
and U5488 (N_5488,N_791,N_1349);
nor U5489 (N_5489,N_980,N_408);
xor U5490 (N_5490,N_760,N_2947);
and U5491 (N_5491,N_2419,N_1948);
and U5492 (N_5492,N_1475,N_1518);
nor U5493 (N_5493,N_2603,N_2251);
nand U5494 (N_5494,N_659,N_1611);
and U5495 (N_5495,N_2064,N_1832);
nand U5496 (N_5496,N_2642,N_1033);
nor U5497 (N_5497,N_780,N_71);
nor U5498 (N_5498,N_925,N_3030);
and U5499 (N_5499,N_691,N_3071);
and U5500 (N_5500,N_2488,N_2861);
xnor U5501 (N_5501,N_2017,N_2590);
or U5502 (N_5502,N_1951,N_2252);
nand U5503 (N_5503,N_259,N_2184);
nand U5504 (N_5504,N_590,N_1188);
and U5505 (N_5505,N_1513,N_1969);
nand U5506 (N_5506,N_2447,N_315);
or U5507 (N_5507,N_304,N_2832);
nor U5508 (N_5508,N_2226,N_1601);
nor U5509 (N_5509,N_1798,N_2384);
xor U5510 (N_5510,N_2691,N_141);
nor U5511 (N_5511,N_1214,N_2779);
or U5512 (N_5512,N_1761,N_2926);
nand U5513 (N_5513,N_3053,N_1460);
or U5514 (N_5514,N_461,N_1284);
xor U5515 (N_5515,N_2025,N_697);
nand U5516 (N_5516,N_319,N_1534);
and U5517 (N_5517,N_158,N_361);
or U5518 (N_5518,N_519,N_2276);
nor U5519 (N_5519,N_2891,N_2436);
or U5520 (N_5520,N_5,N_252);
nor U5521 (N_5521,N_1238,N_1277);
xor U5522 (N_5522,N_586,N_235);
and U5523 (N_5523,N_311,N_3083);
nand U5524 (N_5524,N_506,N_1996);
xnor U5525 (N_5525,N_2559,N_1904);
xnor U5526 (N_5526,N_2412,N_1184);
nand U5527 (N_5527,N_741,N_2850);
nor U5528 (N_5528,N_89,N_2839);
or U5529 (N_5529,N_1717,N_1759);
nand U5530 (N_5530,N_1807,N_1986);
xnor U5531 (N_5531,N_2063,N_1143);
or U5532 (N_5532,N_2311,N_167);
and U5533 (N_5533,N_2510,N_654);
nor U5534 (N_5534,N_2688,N_1810);
or U5535 (N_5535,N_1680,N_1258);
nor U5536 (N_5536,N_1945,N_3006);
nor U5537 (N_5537,N_1926,N_2092);
and U5538 (N_5538,N_83,N_2407);
nand U5539 (N_5539,N_1805,N_1405);
and U5540 (N_5540,N_106,N_2333);
nand U5541 (N_5541,N_2791,N_1444);
and U5542 (N_5542,N_2671,N_2858);
nor U5543 (N_5543,N_159,N_701);
or U5544 (N_5544,N_788,N_1085);
nand U5545 (N_5545,N_1228,N_457);
nand U5546 (N_5546,N_1807,N_661);
and U5547 (N_5547,N_1753,N_2474);
xnor U5548 (N_5548,N_2160,N_2365);
or U5549 (N_5549,N_2669,N_2395);
xor U5550 (N_5550,N_825,N_823);
xor U5551 (N_5551,N_222,N_1754);
xor U5552 (N_5552,N_1314,N_1744);
or U5553 (N_5553,N_1374,N_1364);
xnor U5554 (N_5554,N_1883,N_1526);
nand U5555 (N_5555,N_2560,N_900);
or U5556 (N_5556,N_994,N_3121);
or U5557 (N_5557,N_2248,N_2659);
or U5558 (N_5558,N_895,N_1731);
nand U5559 (N_5559,N_129,N_2698);
xnor U5560 (N_5560,N_2890,N_2790);
nor U5561 (N_5561,N_2631,N_1328);
nor U5562 (N_5562,N_1135,N_628);
nand U5563 (N_5563,N_2455,N_823);
nor U5564 (N_5564,N_2440,N_2408);
nand U5565 (N_5565,N_718,N_2251);
nor U5566 (N_5566,N_1202,N_3057);
nor U5567 (N_5567,N_1817,N_2983);
and U5568 (N_5568,N_3034,N_873);
and U5569 (N_5569,N_2068,N_1847);
nand U5570 (N_5570,N_769,N_1751);
or U5571 (N_5571,N_1186,N_43);
or U5572 (N_5572,N_1244,N_493);
nand U5573 (N_5573,N_2330,N_2465);
nor U5574 (N_5574,N_1986,N_876);
nor U5575 (N_5575,N_228,N_2617);
and U5576 (N_5576,N_1218,N_2914);
xor U5577 (N_5577,N_1459,N_547);
nor U5578 (N_5578,N_3086,N_1210);
nor U5579 (N_5579,N_4,N_337);
xor U5580 (N_5580,N_424,N_1027);
nor U5581 (N_5581,N_222,N_2077);
xnor U5582 (N_5582,N_1571,N_2088);
nand U5583 (N_5583,N_2982,N_2250);
and U5584 (N_5584,N_3087,N_2994);
or U5585 (N_5585,N_2069,N_1210);
or U5586 (N_5586,N_2956,N_2250);
xor U5587 (N_5587,N_1128,N_1974);
or U5588 (N_5588,N_962,N_1710);
and U5589 (N_5589,N_1237,N_3016);
nor U5590 (N_5590,N_1885,N_2057);
nor U5591 (N_5591,N_3047,N_2466);
and U5592 (N_5592,N_2682,N_207);
nor U5593 (N_5593,N_1027,N_1071);
xnor U5594 (N_5594,N_1037,N_2679);
and U5595 (N_5595,N_3095,N_518);
or U5596 (N_5596,N_1427,N_574);
or U5597 (N_5597,N_338,N_193);
and U5598 (N_5598,N_2679,N_185);
nor U5599 (N_5599,N_686,N_1896);
nor U5600 (N_5600,N_584,N_2238);
or U5601 (N_5601,N_1564,N_295);
or U5602 (N_5602,N_1536,N_2063);
xor U5603 (N_5603,N_172,N_153);
xor U5604 (N_5604,N_483,N_2835);
and U5605 (N_5605,N_3123,N_2109);
xnor U5606 (N_5606,N_415,N_1645);
xnor U5607 (N_5607,N_3066,N_1395);
nor U5608 (N_5608,N_1015,N_1198);
nor U5609 (N_5609,N_2969,N_1132);
nor U5610 (N_5610,N_460,N_2933);
and U5611 (N_5611,N_2121,N_1633);
xnor U5612 (N_5612,N_373,N_3118);
nand U5613 (N_5613,N_1384,N_2299);
nand U5614 (N_5614,N_1136,N_2304);
nor U5615 (N_5615,N_2190,N_2713);
nand U5616 (N_5616,N_1932,N_2150);
and U5617 (N_5617,N_32,N_1816);
xor U5618 (N_5618,N_1337,N_2642);
and U5619 (N_5619,N_1947,N_1957);
nand U5620 (N_5620,N_2134,N_1772);
and U5621 (N_5621,N_2083,N_2114);
xor U5622 (N_5622,N_1074,N_223);
nand U5623 (N_5623,N_2401,N_2371);
or U5624 (N_5624,N_2365,N_673);
xor U5625 (N_5625,N_1361,N_2346);
nor U5626 (N_5626,N_1624,N_828);
and U5627 (N_5627,N_1168,N_296);
nor U5628 (N_5628,N_1083,N_627);
nand U5629 (N_5629,N_1570,N_159);
xnor U5630 (N_5630,N_417,N_1849);
nand U5631 (N_5631,N_602,N_495);
nand U5632 (N_5632,N_1755,N_2859);
nor U5633 (N_5633,N_1220,N_2134);
xor U5634 (N_5634,N_1098,N_1806);
nor U5635 (N_5635,N_958,N_1834);
and U5636 (N_5636,N_727,N_281);
and U5637 (N_5637,N_731,N_1232);
nand U5638 (N_5638,N_2322,N_2192);
and U5639 (N_5639,N_1409,N_1185);
or U5640 (N_5640,N_1234,N_1148);
or U5641 (N_5641,N_2645,N_959);
nand U5642 (N_5642,N_3046,N_2569);
or U5643 (N_5643,N_1012,N_1950);
and U5644 (N_5644,N_1240,N_1187);
xor U5645 (N_5645,N_1212,N_2871);
nand U5646 (N_5646,N_1097,N_1160);
nor U5647 (N_5647,N_1343,N_2548);
xnor U5648 (N_5648,N_191,N_1475);
or U5649 (N_5649,N_215,N_1867);
nor U5650 (N_5650,N_200,N_1678);
or U5651 (N_5651,N_2912,N_2187);
or U5652 (N_5652,N_2315,N_728);
and U5653 (N_5653,N_2085,N_513);
xnor U5654 (N_5654,N_3100,N_692);
xnor U5655 (N_5655,N_584,N_1916);
xor U5656 (N_5656,N_2394,N_781);
or U5657 (N_5657,N_2992,N_2359);
or U5658 (N_5658,N_2916,N_929);
xnor U5659 (N_5659,N_1505,N_2331);
or U5660 (N_5660,N_963,N_729);
nor U5661 (N_5661,N_477,N_1845);
nand U5662 (N_5662,N_2765,N_1550);
nand U5663 (N_5663,N_2257,N_3088);
nand U5664 (N_5664,N_678,N_473);
nand U5665 (N_5665,N_317,N_991);
or U5666 (N_5666,N_2995,N_1797);
or U5667 (N_5667,N_1773,N_1315);
and U5668 (N_5668,N_1291,N_2780);
or U5669 (N_5669,N_3099,N_2707);
nand U5670 (N_5670,N_2981,N_2849);
or U5671 (N_5671,N_1855,N_2000);
nand U5672 (N_5672,N_23,N_394);
nand U5673 (N_5673,N_2604,N_2003);
nand U5674 (N_5674,N_372,N_1343);
and U5675 (N_5675,N_1572,N_305);
xor U5676 (N_5676,N_1163,N_2573);
and U5677 (N_5677,N_876,N_3066);
nor U5678 (N_5678,N_1943,N_1122);
xnor U5679 (N_5679,N_2712,N_2217);
nand U5680 (N_5680,N_1720,N_671);
xnor U5681 (N_5681,N_2372,N_2871);
and U5682 (N_5682,N_1872,N_2477);
xnor U5683 (N_5683,N_128,N_309);
nand U5684 (N_5684,N_2694,N_1013);
and U5685 (N_5685,N_1729,N_2517);
nand U5686 (N_5686,N_1351,N_564);
and U5687 (N_5687,N_1635,N_644);
nor U5688 (N_5688,N_1099,N_2099);
xor U5689 (N_5689,N_824,N_849);
nand U5690 (N_5690,N_2997,N_1582);
nand U5691 (N_5691,N_183,N_1756);
or U5692 (N_5692,N_60,N_517);
and U5693 (N_5693,N_2325,N_550);
nor U5694 (N_5694,N_2505,N_1102);
and U5695 (N_5695,N_2734,N_1507);
and U5696 (N_5696,N_3040,N_2944);
nor U5697 (N_5697,N_2282,N_2490);
or U5698 (N_5698,N_703,N_1256);
xnor U5699 (N_5699,N_1555,N_894);
xnor U5700 (N_5700,N_1719,N_2587);
or U5701 (N_5701,N_2606,N_2776);
or U5702 (N_5702,N_3036,N_2603);
or U5703 (N_5703,N_874,N_761);
and U5704 (N_5704,N_2241,N_406);
and U5705 (N_5705,N_2330,N_2828);
xnor U5706 (N_5706,N_3091,N_2260);
xnor U5707 (N_5707,N_1166,N_3112);
and U5708 (N_5708,N_895,N_1635);
and U5709 (N_5709,N_2199,N_2017);
and U5710 (N_5710,N_3103,N_1772);
or U5711 (N_5711,N_780,N_1739);
xnor U5712 (N_5712,N_509,N_30);
xor U5713 (N_5713,N_2051,N_2242);
nand U5714 (N_5714,N_816,N_1358);
or U5715 (N_5715,N_2779,N_1670);
xor U5716 (N_5716,N_2713,N_2863);
nand U5717 (N_5717,N_958,N_1445);
xnor U5718 (N_5718,N_807,N_2678);
or U5719 (N_5719,N_679,N_539);
nor U5720 (N_5720,N_2900,N_2728);
nand U5721 (N_5721,N_565,N_1613);
and U5722 (N_5722,N_1965,N_251);
or U5723 (N_5723,N_2997,N_2643);
or U5724 (N_5724,N_890,N_1170);
nor U5725 (N_5725,N_2040,N_617);
nor U5726 (N_5726,N_1981,N_1310);
or U5727 (N_5727,N_2432,N_985);
nand U5728 (N_5728,N_3103,N_2128);
nor U5729 (N_5729,N_2229,N_688);
nand U5730 (N_5730,N_2742,N_1675);
or U5731 (N_5731,N_427,N_2261);
nor U5732 (N_5732,N_2183,N_2044);
or U5733 (N_5733,N_2248,N_202);
or U5734 (N_5734,N_235,N_1359);
nor U5735 (N_5735,N_1329,N_2837);
nor U5736 (N_5736,N_214,N_968);
nand U5737 (N_5737,N_1201,N_933);
nand U5738 (N_5738,N_2269,N_336);
xor U5739 (N_5739,N_2813,N_2822);
nor U5740 (N_5740,N_1637,N_2867);
xnor U5741 (N_5741,N_810,N_1991);
nor U5742 (N_5742,N_2862,N_1569);
nor U5743 (N_5743,N_2035,N_3062);
nor U5744 (N_5744,N_1180,N_2252);
or U5745 (N_5745,N_2523,N_2194);
and U5746 (N_5746,N_2244,N_110);
nor U5747 (N_5747,N_1253,N_1428);
nand U5748 (N_5748,N_1496,N_1996);
and U5749 (N_5749,N_2351,N_188);
nand U5750 (N_5750,N_2619,N_3031);
xnor U5751 (N_5751,N_1792,N_2318);
xor U5752 (N_5752,N_69,N_3011);
or U5753 (N_5753,N_1822,N_475);
xnor U5754 (N_5754,N_658,N_2667);
and U5755 (N_5755,N_1232,N_1684);
xnor U5756 (N_5756,N_923,N_600);
xnor U5757 (N_5757,N_1401,N_851);
xor U5758 (N_5758,N_1059,N_1659);
nand U5759 (N_5759,N_2057,N_961);
and U5760 (N_5760,N_913,N_1557);
or U5761 (N_5761,N_135,N_357);
or U5762 (N_5762,N_2067,N_2533);
and U5763 (N_5763,N_1370,N_872);
xnor U5764 (N_5764,N_2943,N_533);
nand U5765 (N_5765,N_15,N_2711);
nand U5766 (N_5766,N_930,N_1970);
and U5767 (N_5767,N_1236,N_319);
and U5768 (N_5768,N_2624,N_1060);
nor U5769 (N_5769,N_1101,N_1102);
xor U5770 (N_5770,N_215,N_2722);
xor U5771 (N_5771,N_2021,N_2316);
or U5772 (N_5772,N_228,N_1681);
nand U5773 (N_5773,N_2425,N_1178);
nor U5774 (N_5774,N_1148,N_1308);
nand U5775 (N_5775,N_494,N_1115);
and U5776 (N_5776,N_3043,N_1333);
or U5777 (N_5777,N_421,N_509);
and U5778 (N_5778,N_2389,N_1010);
nor U5779 (N_5779,N_1979,N_2881);
nor U5780 (N_5780,N_1567,N_360);
or U5781 (N_5781,N_2262,N_3083);
and U5782 (N_5782,N_1892,N_1703);
or U5783 (N_5783,N_3077,N_1389);
nor U5784 (N_5784,N_1491,N_1435);
nor U5785 (N_5785,N_1623,N_1634);
nor U5786 (N_5786,N_1751,N_2402);
xor U5787 (N_5787,N_332,N_818);
xnor U5788 (N_5788,N_2486,N_851);
nand U5789 (N_5789,N_253,N_1246);
xnor U5790 (N_5790,N_1994,N_1819);
nand U5791 (N_5791,N_2595,N_929);
xnor U5792 (N_5792,N_415,N_579);
nor U5793 (N_5793,N_981,N_1452);
or U5794 (N_5794,N_2935,N_1713);
nand U5795 (N_5795,N_256,N_121);
nand U5796 (N_5796,N_2656,N_967);
or U5797 (N_5797,N_1806,N_1708);
and U5798 (N_5798,N_1052,N_1817);
or U5799 (N_5799,N_2528,N_405);
and U5800 (N_5800,N_2212,N_902);
or U5801 (N_5801,N_2803,N_945);
nor U5802 (N_5802,N_370,N_1443);
xor U5803 (N_5803,N_2047,N_585);
and U5804 (N_5804,N_1820,N_1734);
nand U5805 (N_5805,N_312,N_260);
or U5806 (N_5806,N_1107,N_2124);
nand U5807 (N_5807,N_1463,N_2089);
or U5808 (N_5808,N_357,N_665);
and U5809 (N_5809,N_1401,N_811);
nand U5810 (N_5810,N_2880,N_2688);
xor U5811 (N_5811,N_2441,N_549);
nand U5812 (N_5812,N_1431,N_2609);
xor U5813 (N_5813,N_562,N_1067);
nor U5814 (N_5814,N_1800,N_2596);
xor U5815 (N_5815,N_73,N_656);
nand U5816 (N_5816,N_2669,N_1900);
nor U5817 (N_5817,N_1605,N_321);
xnor U5818 (N_5818,N_1114,N_3048);
or U5819 (N_5819,N_793,N_1137);
nand U5820 (N_5820,N_973,N_1639);
xor U5821 (N_5821,N_977,N_409);
and U5822 (N_5822,N_1600,N_1781);
nand U5823 (N_5823,N_1518,N_2457);
xor U5824 (N_5824,N_810,N_1835);
nand U5825 (N_5825,N_1467,N_339);
and U5826 (N_5826,N_2926,N_502);
xor U5827 (N_5827,N_2202,N_2900);
nand U5828 (N_5828,N_2614,N_2391);
or U5829 (N_5829,N_140,N_1162);
and U5830 (N_5830,N_173,N_1309);
nand U5831 (N_5831,N_582,N_1092);
or U5832 (N_5832,N_794,N_2233);
xor U5833 (N_5833,N_2275,N_66);
nor U5834 (N_5834,N_1786,N_2208);
nor U5835 (N_5835,N_1371,N_2390);
nor U5836 (N_5836,N_1753,N_2389);
nand U5837 (N_5837,N_346,N_1076);
xnor U5838 (N_5838,N_1445,N_829);
xnor U5839 (N_5839,N_2452,N_1554);
nor U5840 (N_5840,N_2083,N_75);
or U5841 (N_5841,N_2070,N_154);
nor U5842 (N_5842,N_1158,N_1122);
or U5843 (N_5843,N_2436,N_2175);
or U5844 (N_5844,N_807,N_2841);
xnor U5845 (N_5845,N_97,N_2952);
nand U5846 (N_5846,N_2217,N_2658);
and U5847 (N_5847,N_1573,N_495);
xnor U5848 (N_5848,N_2679,N_2498);
nor U5849 (N_5849,N_956,N_682);
xor U5850 (N_5850,N_1627,N_2846);
xor U5851 (N_5851,N_2346,N_2541);
nand U5852 (N_5852,N_259,N_306);
nor U5853 (N_5853,N_1924,N_15);
xnor U5854 (N_5854,N_1610,N_2109);
nand U5855 (N_5855,N_1970,N_1481);
xor U5856 (N_5856,N_1867,N_2250);
nor U5857 (N_5857,N_2857,N_2804);
nand U5858 (N_5858,N_2426,N_111);
nor U5859 (N_5859,N_1308,N_1641);
nor U5860 (N_5860,N_3023,N_215);
and U5861 (N_5861,N_1160,N_1036);
xor U5862 (N_5862,N_1157,N_2109);
xnor U5863 (N_5863,N_1317,N_1497);
or U5864 (N_5864,N_295,N_186);
and U5865 (N_5865,N_393,N_62);
xnor U5866 (N_5866,N_1708,N_2366);
or U5867 (N_5867,N_1956,N_1296);
nor U5868 (N_5868,N_256,N_289);
nor U5869 (N_5869,N_2367,N_1960);
xnor U5870 (N_5870,N_855,N_1748);
xnor U5871 (N_5871,N_149,N_1280);
nand U5872 (N_5872,N_758,N_2459);
and U5873 (N_5873,N_1361,N_2922);
or U5874 (N_5874,N_241,N_3034);
xor U5875 (N_5875,N_2136,N_797);
and U5876 (N_5876,N_1946,N_713);
nor U5877 (N_5877,N_1191,N_930);
xnor U5878 (N_5878,N_370,N_2785);
nor U5879 (N_5879,N_48,N_1374);
xor U5880 (N_5880,N_2269,N_1358);
or U5881 (N_5881,N_2660,N_1008);
xnor U5882 (N_5882,N_510,N_1755);
nor U5883 (N_5883,N_1865,N_1845);
nor U5884 (N_5884,N_121,N_2778);
and U5885 (N_5885,N_1112,N_2647);
and U5886 (N_5886,N_2021,N_2599);
or U5887 (N_5887,N_99,N_289);
nand U5888 (N_5888,N_2894,N_221);
nand U5889 (N_5889,N_2639,N_2370);
or U5890 (N_5890,N_2894,N_396);
and U5891 (N_5891,N_2039,N_1133);
and U5892 (N_5892,N_2389,N_465);
xnor U5893 (N_5893,N_431,N_2853);
nand U5894 (N_5894,N_2647,N_667);
or U5895 (N_5895,N_1802,N_2921);
xor U5896 (N_5896,N_29,N_2706);
xor U5897 (N_5897,N_1889,N_352);
or U5898 (N_5898,N_483,N_547);
or U5899 (N_5899,N_2363,N_36);
nor U5900 (N_5900,N_2647,N_2922);
nand U5901 (N_5901,N_1009,N_589);
xor U5902 (N_5902,N_867,N_252);
xnor U5903 (N_5903,N_910,N_1747);
nor U5904 (N_5904,N_1537,N_1848);
nand U5905 (N_5905,N_2660,N_2990);
or U5906 (N_5906,N_2534,N_537);
nand U5907 (N_5907,N_2283,N_1506);
xor U5908 (N_5908,N_664,N_2873);
or U5909 (N_5909,N_1617,N_1910);
xor U5910 (N_5910,N_1036,N_1066);
xnor U5911 (N_5911,N_2197,N_462);
or U5912 (N_5912,N_1362,N_955);
nand U5913 (N_5913,N_2121,N_2030);
and U5914 (N_5914,N_2370,N_1584);
or U5915 (N_5915,N_2919,N_2135);
nand U5916 (N_5916,N_2514,N_1693);
and U5917 (N_5917,N_1956,N_827);
nor U5918 (N_5918,N_442,N_108);
and U5919 (N_5919,N_883,N_2041);
or U5920 (N_5920,N_220,N_2436);
and U5921 (N_5921,N_660,N_1185);
or U5922 (N_5922,N_1319,N_2428);
nor U5923 (N_5923,N_2164,N_1155);
and U5924 (N_5924,N_1366,N_324);
nand U5925 (N_5925,N_2114,N_2238);
nand U5926 (N_5926,N_1212,N_2253);
or U5927 (N_5927,N_2138,N_2842);
nor U5928 (N_5928,N_1321,N_1631);
nor U5929 (N_5929,N_131,N_1200);
or U5930 (N_5930,N_2186,N_2708);
nor U5931 (N_5931,N_194,N_1738);
nand U5932 (N_5932,N_1362,N_1807);
nand U5933 (N_5933,N_172,N_1858);
xor U5934 (N_5934,N_3081,N_1128);
or U5935 (N_5935,N_1950,N_2818);
and U5936 (N_5936,N_2133,N_2009);
nand U5937 (N_5937,N_1106,N_1761);
or U5938 (N_5938,N_3123,N_679);
xnor U5939 (N_5939,N_2833,N_2100);
or U5940 (N_5940,N_1124,N_2621);
and U5941 (N_5941,N_1188,N_31);
nor U5942 (N_5942,N_2522,N_413);
nor U5943 (N_5943,N_1216,N_1047);
xor U5944 (N_5944,N_2816,N_2767);
xnor U5945 (N_5945,N_2114,N_913);
or U5946 (N_5946,N_849,N_1007);
nor U5947 (N_5947,N_1062,N_707);
xnor U5948 (N_5948,N_1570,N_2416);
xor U5949 (N_5949,N_626,N_1043);
nand U5950 (N_5950,N_626,N_428);
or U5951 (N_5951,N_1739,N_2519);
xnor U5952 (N_5952,N_2305,N_23);
and U5953 (N_5953,N_2170,N_43);
and U5954 (N_5954,N_444,N_2509);
or U5955 (N_5955,N_3045,N_2647);
and U5956 (N_5956,N_775,N_2820);
nand U5957 (N_5957,N_1015,N_2286);
or U5958 (N_5958,N_2804,N_2720);
nand U5959 (N_5959,N_1861,N_1965);
nor U5960 (N_5960,N_2455,N_142);
xnor U5961 (N_5961,N_970,N_1307);
nand U5962 (N_5962,N_1726,N_3023);
xnor U5963 (N_5963,N_1375,N_1440);
xor U5964 (N_5964,N_880,N_141);
and U5965 (N_5965,N_2825,N_1396);
nor U5966 (N_5966,N_955,N_2609);
nor U5967 (N_5967,N_2123,N_1659);
xnor U5968 (N_5968,N_142,N_286);
xor U5969 (N_5969,N_1935,N_2266);
xnor U5970 (N_5970,N_869,N_2709);
nor U5971 (N_5971,N_2731,N_1674);
and U5972 (N_5972,N_2851,N_1099);
and U5973 (N_5973,N_181,N_342);
xnor U5974 (N_5974,N_2917,N_601);
or U5975 (N_5975,N_2500,N_385);
nand U5976 (N_5976,N_2268,N_1229);
and U5977 (N_5977,N_3115,N_520);
or U5978 (N_5978,N_72,N_2435);
xnor U5979 (N_5979,N_2491,N_831);
nand U5980 (N_5980,N_1981,N_2291);
nand U5981 (N_5981,N_1296,N_1228);
xnor U5982 (N_5982,N_1422,N_1191);
and U5983 (N_5983,N_3098,N_1648);
xor U5984 (N_5984,N_538,N_1740);
nand U5985 (N_5985,N_102,N_1396);
or U5986 (N_5986,N_2161,N_75);
or U5987 (N_5987,N_850,N_2948);
nand U5988 (N_5988,N_1619,N_131);
and U5989 (N_5989,N_2427,N_2997);
and U5990 (N_5990,N_1657,N_611);
or U5991 (N_5991,N_1990,N_1415);
nand U5992 (N_5992,N_1237,N_1336);
nor U5993 (N_5993,N_1264,N_1698);
or U5994 (N_5994,N_1523,N_759);
and U5995 (N_5995,N_2433,N_3079);
xor U5996 (N_5996,N_1813,N_1817);
nand U5997 (N_5997,N_1244,N_1003);
or U5998 (N_5998,N_2805,N_2051);
nor U5999 (N_5999,N_1045,N_1912);
xnor U6000 (N_6000,N_192,N_3106);
and U6001 (N_6001,N_2304,N_1429);
nand U6002 (N_6002,N_1292,N_1589);
or U6003 (N_6003,N_866,N_684);
or U6004 (N_6004,N_1272,N_1092);
or U6005 (N_6005,N_1558,N_2197);
or U6006 (N_6006,N_1780,N_1698);
or U6007 (N_6007,N_895,N_3092);
xnor U6008 (N_6008,N_2573,N_1152);
nor U6009 (N_6009,N_3115,N_1819);
nor U6010 (N_6010,N_755,N_747);
nand U6011 (N_6011,N_671,N_1716);
nor U6012 (N_6012,N_1956,N_2934);
or U6013 (N_6013,N_723,N_2161);
nand U6014 (N_6014,N_2321,N_2920);
or U6015 (N_6015,N_305,N_30);
or U6016 (N_6016,N_2493,N_1398);
and U6017 (N_6017,N_2705,N_1336);
xnor U6018 (N_6018,N_2133,N_1495);
nand U6019 (N_6019,N_399,N_1719);
nor U6020 (N_6020,N_356,N_698);
nor U6021 (N_6021,N_198,N_2934);
or U6022 (N_6022,N_723,N_2599);
or U6023 (N_6023,N_1250,N_2342);
xor U6024 (N_6024,N_2160,N_2244);
xor U6025 (N_6025,N_1475,N_2573);
xor U6026 (N_6026,N_2348,N_2234);
or U6027 (N_6027,N_901,N_724);
nor U6028 (N_6028,N_704,N_3038);
nand U6029 (N_6029,N_241,N_443);
xor U6030 (N_6030,N_3116,N_1551);
or U6031 (N_6031,N_2180,N_672);
xnor U6032 (N_6032,N_385,N_1312);
and U6033 (N_6033,N_665,N_1485);
nor U6034 (N_6034,N_593,N_2648);
nand U6035 (N_6035,N_886,N_1420);
nor U6036 (N_6036,N_1259,N_2132);
xnor U6037 (N_6037,N_2671,N_576);
nand U6038 (N_6038,N_331,N_2035);
nor U6039 (N_6039,N_925,N_1659);
or U6040 (N_6040,N_2889,N_104);
and U6041 (N_6041,N_2951,N_807);
and U6042 (N_6042,N_3025,N_3094);
or U6043 (N_6043,N_1900,N_2310);
and U6044 (N_6044,N_2042,N_2734);
nor U6045 (N_6045,N_2349,N_2775);
nor U6046 (N_6046,N_599,N_1984);
nand U6047 (N_6047,N_1094,N_2505);
nand U6048 (N_6048,N_1620,N_136);
nor U6049 (N_6049,N_2075,N_1259);
or U6050 (N_6050,N_2319,N_2556);
xnor U6051 (N_6051,N_1906,N_2275);
xnor U6052 (N_6052,N_328,N_1824);
and U6053 (N_6053,N_2281,N_692);
xnor U6054 (N_6054,N_2748,N_1050);
xnor U6055 (N_6055,N_2239,N_1477);
nor U6056 (N_6056,N_1813,N_129);
and U6057 (N_6057,N_1355,N_854);
nand U6058 (N_6058,N_132,N_329);
nor U6059 (N_6059,N_1980,N_34);
or U6060 (N_6060,N_2762,N_3098);
nand U6061 (N_6061,N_2112,N_3015);
xnor U6062 (N_6062,N_1852,N_694);
xnor U6063 (N_6063,N_1242,N_1337);
nand U6064 (N_6064,N_1002,N_3012);
and U6065 (N_6065,N_296,N_2103);
and U6066 (N_6066,N_909,N_2917);
xnor U6067 (N_6067,N_3068,N_1554);
nor U6068 (N_6068,N_304,N_336);
nand U6069 (N_6069,N_1196,N_2018);
or U6070 (N_6070,N_2090,N_2513);
and U6071 (N_6071,N_1942,N_2571);
and U6072 (N_6072,N_2844,N_1568);
xnor U6073 (N_6073,N_1162,N_2517);
or U6074 (N_6074,N_2829,N_940);
nor U6075 (N_6075,N_2290,N_877);
nand U6076 (N_6076,N_2860,N_2021);
nor U6077 (N_6077,N_1762,N_2713);
nor U6078 (N_6078,N_1031,N_400);
xor U6079 (N_6079,N_2996,N_1055);
nor U6080 (N_6080,N_2424,N_2552);
or U6081 (N_6081,N_31,N_666);
nor U6082 (N_6082,N_1186,N_370);
xnor U6083 (N_6083,N_410,N_2808);
nand U6084 (N_6084,N_2870,N_245);
and U6085 (N_6085,N_210,N_2799);
xor U6086 (N_6086,N_1941,N_985);
nand U6087 (N_6087,N_100,N_246);
nor U6088 (N_6088,N_1241,N_644);
xor U6089 (N_6089,N_2278,N_2097);
and U6090 (N_6090,N_856,N_1759);
nand U6091 (N_6091,N_1312,N_925);
and U6092 (N_6092,N_1616,N_2614);
or U6093 (N_6093,N_578,N_2290);
nand U6094 (N_6094,N_1682,N_1729);
nor U6095 (N_6095,N_1036,N_350);
and U6096 (N_6096,N_3030,N_2790);
and U6097 (N_6097,N_2304,N_1307);
nor U6098 (N_6098,N_2951,N_707);
nor U6099 (N_6099,N_1268,N_1494);
or U6100 (N_6100,N_1145,N_1391);
xor U6101 (N_6101,N_1111,N_1946);
xor U6102 (N_6102,N_2953,N_783);
xor U6103 (N_6103,N_2936,N_2686);
xnor U6104 (N_6104,N_1305,N_1757);
or U6105 (N_6105,N_2759,N_2998);
nor U6106 (N_6106,N_758,N_217);
nand U6107 (N_6107,N_507,N_2848);
nand U6108 (N_6108,N_2148,N_1493);
or U6109 (N_6109,N_1363,N_3074);
nor U6110 (N_6110,N_2007,N_2541);
or U6111 (N_6111,N_2427,N_2794);
nand U6112 (N_6112,N_2406,N_1945);
and U6113 (N_6113,N_2203,N_72);
and U6114 (N_6114,N_2569,N_656);
xor U6115 (N_6115,N_364,N_1203);
nor U6116 (N_6116,N_237,N_2157);
or U6117 (N_6117,N_50,N_2269);
xnor U6118 (N_6118,N_1832,N_1219);
and U6119 (N_6119,N_2236,N_1814);
or U6120 (N_6120,N_616,N_42);
nor U6121 (N_6121,N_1374,N_2014);
nand U6122 (N_6122,N_1158,N_2860);
or U6123 (N_6123,N_1553,N_1588);
nand U6124 (N_6124,N_361,N_2621);
xor U6125 (N_6125,N_2644,N_2426);
or U6126 (N_6126,N_1609,N_726);
or U6127 (N_6127,N_1311,N_3112);
xor U6128 (N_6128,N_837,N_985);
nor U6129 (N_6129,N_1707,N_1031);
or U6130 (N_6130,N_1607,N_868);
nand U6131 (N_6131,N_974,N_3111);
and U6132 (N_6132,N_2932,N_1115);
or U6133 (N_6133,N_131,N_2819);
and U6134 (N_6134,N_1354,N_1066);
nor U6135 (N_6135,N_2879,N_1133);
nor U6136 (N_6136,N_2681,N_2386);
nand U6137 (N_6137,N_3082,N_2386);
nor U6138 (N_6138,N_887,N_1001);
or U6139 (N_6139,N_2110,N_682);
nor U6140 (N_6140,N_761,N_3045);
and U6141 (N_6141,N_2204,N_2038);
or U6142 (N_6142,N_460,N_1140);
xor U6143 (N_6143,N_1450,N_3101);
and U6144 (N_6144,N_2238,N_927);
xor U6145 (N_6145,N_368,N_317);
or U6146 (N_6146,N_2674,N_2813);
or U6147 (N_6147,N_721,N_1468);
xor U6148 (N_6148,N_1856,N_1696);
nor U6149 (N_6149,N_366,N_2515);
and U6150 (N_6150,N_1016,N_338);
and U6151 (N_6151,N_1445,N_1664);
nand U6152 (N_6152,N_6,N_917);
and U6153 (N_6153,N_2973,N_126);
nor U6154 (N_6154,N_1068,N_1789);
xor U6155 (N_6155,N_1177,N_28);
nand U6156 (N_6156,N_2015,N_2994);
and U6157 (N_6157,N_746,N_1302);
nand U6158 (N_6158,N_1875,N_1440);
or U6159 (N_6159,N_319,N_1921);
xnor U6160 (N_6160,N_2246,N_2560);
or U6161 (N_6161,N_1766,N_2639);
xnor U6162 (N_6162,N_2608,N_166);
xnor U6163 (N_6163,N_303,N_2806);
or U6164 (N_6164,N_2567,N_738);
nor U6165 (N_6165,N_3039,N_791);
and U6166 (N_6166,N_936,N_480);
and U6167 (N_6167,N_1336,N_2317);
or U6168 (N_6168,N_3053,N_3095);
or U6169 (N_6169,N_2814,N_2221);
or U6170 (N_6170,N_2292,N_2819);
nor U6171 (N_6171,N_2583,N_2);
xor U6172 (N_6172,N_746,N_1790);
nor U6173 (N_6173,N_1766,N_966);
nand U6174 (N_6174,N_1723,N_367);
xnor U6175 (N_6175,N_2328,N_1406);
or U6176 (N_6176,N_1937,N_2198);
nor U6177 (N_6177,N_1342,N_2166);
nor U6178 (N_6178,N_1165,N_668);
nand U6179 (N_6179,N_809,N_2534);
nor U6180 (N_6180,N_1182,N_1246);
nand U6181 (N_6181,N_2852,N_1319);
nand U6182 (N_6182,N_2880,N_2386);
nand U6183 (N_6183,N_2095,N_1471);
or U6184 (N_6184,N_2170,N_3117);
xnor U6185 (N_6185,N_1677,N_964);
nor U6186 (N_6186,N_3101,N_566);
nor U6187 (N_6187,N_1501,N_2170);
nand U6188 (N_6188,N_1381,N_933);
nor U6189 (N_6189,N_1180,N_1866);
xor U6190 (N_6190,N_2825,N_734);
and U6191 (N_6191,N_1249,N_2622);
and U6192 (N_6192,N_1251,N_1310);
nand U6193 (N_6193,N_2113,N_2438);
nand U6194 (N_6194,N_1455,N_2469);
or U6195 (N_6195,N_2666,N_1858);
nand U6196 (N_6196,N_2248,N_475);
nand U6197 (N_6197,N_660,N_2786);
nor U6198 (N_6198,N_973,N_448);
and U6199 (N_6199,N_1327,N_3046);
xor U6200 (N_6200,N_1057,N_1994);
or U6201 (N_6201,N_1276,N_229);
xor U6202 (N_6202,N_274,N_3039);
xor U6203 (N_6203,N_2260,N_2980);
and U6204 (N_6204,N_820,N_541);
and U6205 (N_6205,N_106,N_136);
nand U6206 (N_6206,N_2638,N_182);
or U6207 (N_6207,N_1622,N_2958);
nor U6208 (N_6208,N_245,N_347);
nand U6209 (N_6209,N_2200,N_656);
and U6210 (N_6210,N_1555,N_2405);
xnor U6211 (N_6211,N_1650,N_1384);
and U6212 (N_6212,N_1489,N_2880);
or U6213 (N_6213,N_545,N_1158);
or U6214 (N_6214,N_223,N_2217);
xor U6215 (N_6215,N_2102,N_2569);
nand U6216 (N_6216,N_1744,N_2607);
xor U6217 (N_6217,N_999,N_630);
nor U6218 (N_6218,N_3068,N_302);
xnor U6219 (N_6219,N_1307,N_3120);
nor U6220 (N_6220,N_1294,N_2756);
or U6221 (N_6221,N_2475,N_261);
and U6222 (N_6222,N_1474,N_2528);
or U6223 (N_6223,N_1177,N_2106);
nand U6224 (N_6224,N_2306,N_518);
or U6225 (N_6225,N_2422,N_2791);
or U6226 (N_6226,N_1853,N_53);
xnor U6227 (N_6227,N_2518,N_1404);
nor U6228 (N_6228,N_265,N_1276);
nand U6229 (N_6229,N_754,N_1185);
nand U6230 (N_6230,N_1870,N_2216);
xor U6231 (N_6231,N_780,N_1460);
or U6232 (N_6232,N_2071,N_2109);
nand U6233 (N_6233,N_862,N_2326);
xnor U6234 (N_6234,N_269,N_2292);
nor U6235 (N_6235,N_1233,N_2691);
xor U6236 (N_6236,N_46,N_867);
or U6237 (N_6237,N_2401,N_356);
nor U6238 (N_6238,N_2377,N_2317);
nor U6239 (N_6239,N_1558,N_547);
nand U6240 (N_6240,N_2187,N_340);
nor U6241 (N_6241,N_128,N_1376);
nand U6242 (N_6242,N_1780,N_1069);
xor U6243 (N_6243,N_1924,N_2150);
xnor U6244 (N_6244,N_839,N_673);
and U6245 (N_6245,N_1043,N_269);
nor U6246 (N_6246,N_73,N_1727);
or U6247 (N_6247,N_978,N_1335);
xor U6248 (N_6248,N_173,N_129);
and U6249 (N_6249,N_335,N_1405);
or U6250 (N_6250,N_5339,N_5286);
xor U6251 (N_6251,N_3980,N_5549);
nand U6252 (N_6252,N_5178,N_5236);
nor U6253 (N_6253,N_4991,N_5095);
or U6254 (N_6254,N_3924,N_3140);
and U6255 (N_6255,N_4738,N_3446);
nand U6256 (N_6256,N_5189,N_5381);
nand U6257 (N_6257,N_6055,N_5393);
xor U6258 (N_6258,N_5616,N_5647);
nor U6259 (N_6259,N_5235,N_5800);
xnor U6260 (N_6260,N_5551,N_3670);
nand U6261 (N_6261,N_3815,N_3428);
and U6262 (N_6262,N_5994,N_3400);
or U6263 (N_6263,N_4503,N_3675);
xnor U6264 (N_6264,N_5972,N_4277);
xor U6265 (N_6265,N_3659,N_3649);
nor U6266 (N_6266,N_4719,N_5300);
nor U6267 (N_6267,N_4588,N_3759);
nor U6268 (N_6268,N_5051,N_5259);
xor U6269 (N_6269,N_4021,N_4649);
nor U6270 (N_6270,N_3286,N_3385);
nor U6271 (N_6271,N_4710,N_3389);
nand U6272 (N_6272,N_4753,N_3483);
nor U6273 (N_6273,N_3343,N_4650);
xnor U6274 (N_6274,N_3854,N_4733);
and U6275 (N_6275,N_3193,N_5359);
nand U6276 (N_6276,N_4884,N_4903);
nand U6277 (N_6277,N_6037,N_3474);
and U6278 (N_6278,N_4613,N_5498);
xor U6279 (N_6279,N_4105,N_4458);
xor U6280 (N_6280,N_4469,N_5078);
and U6281 (N_6281,N_3831,N_3674);
nand U6282 (N_6282,N_4915,N_4846);
nand U6283 (N_6283,N_5639,N_4533);
nand U6284 (N_6284,N_6153,N_3168);
nand U6285 (N_6285,N_3973,N_3608);
nand U6286 (N_6286,N_5501,N_3653);
xnor U6287 (N_6287,N_5684,N_3233);
or U6288 (N_6288,N_5042,N_3956);
or U6289 (N_6289,N_5443,N_4525);
nor U6290 (N_6290,N_4102,N_3497);
and U6291 (N_6291,N_4468,N_5998);
and U6292 (N_6292,N_4055,N_4434);
or U6293 (N_6293,N_5249,N_4078);
nor U6294 (N_6294,N_6061,N_5055);
nor U6295 (N_6295,N_4000,N_3868);
xor U6296 (N_6296,N_4068,N_4638);
nor U6297 (N_6297,N_4621,N_4653);
nor U6298 (N_6298,N_3901,N_5390);
nor U6299 (N_6299,N_6160,N_3421);
or U6300 (N_6300,N_4729,N_5480);
or U6301 (N_6301,N_3988,N_3452);
and U6302 (N_6302,N_4803,N_3787);
or U6303 (N_6303,N_3412,N_4894);
nor U6304 (N_6304,N_3906,N_6092);
nor U6305 (N_6305,N_3426,N_4788);
nand U6306 (N_6306,N_5168,N_5840);
nor U6307 (N_6307,N_4866,N_4930);
nand U6308 (N_6308,N_5242,N_4839);
or U6309 (N_6309,N_4791,N_4700);
nor U6310 (N_6310,N_3641,N_3833);
or U6311 (N_6311,N_5538,N_4426);
and U6312 (N_6312,N_3645,N_4331);
or U6313 (N_6313,N_4361,N_3779);
nand U6314 (N_6314,N_4197,N_4233);
and U6315 (N_6315,N_4770,N_4948);
xor U6316 (N_6316,N_5196,N_5985);
nand U6317 (N_6317,N_4848,N_5212);
and U6318 (N_6318,N_3609,N_5417);
nand U6319 (N_6319,N_3972,N_4965);
nor U6320 (N_6320,N_6012,N_3276);
or U6321 (N_6321,N_4179,N_4306);
nor U6322 (N_6322,N_3558,N_5150);
xnor U6323 (N_6323,N_6050,N_4294);
nor U6324 (N_6324,N_3741,N_6210);
nand U6325 (N_6325,N_3699,N_4040);
nand U6326 (N_6326,N_4027,N_4919);
nand U6327 (N_6327,N_5920,N_3561);
or U6328 (N_6328,N_5522,N_5869);
xnor U6329 (N_6329,N_5823,N_5354);
nand U6330 (N_6330,N_5026,N_3437);
or U6331 (N_6331,N_5872,N_5370);
nor U6332 (N_6332,N_5743,N_5490);
or U6333 (N_6333,N_3777,N_3520);
nor U6334 (N_6334,N_3161,N_3163);
or U6335 (N_6335,N_4366,N_3993);
and U6336 (N_6336,N_5137,N_4432);
and U6337 (N_6337,N_6045,N_3642);
or U6338 (N_6338,N_5697,N_3771);
nor U6339 (N_6339,N_4928,N_3480);
nand U6340 (N_6340,N_3733,N_4881);
nand U6341 (N_6341,N_3475,N_4013);
and U6342 (N_6342,N_3295,N_3309);
and U6343 (N_6343,N_3834,N_3877);
xnor U6344 (N_6344,N_3555,N_4995);
and U6345 (N_6345,N_3795,N_4499);
and U6346 (N_6346,N_5730,N_4768);
or U6347 (N_6347,N_4993,N_4139);
nor U6348 (N_6348,N_5158,N_4180);
nand U6349 (N_6349,N_6211,N_4832);
nand U6350 (N_6350,N_5890,N_5266);
or U6351 (N_6351,N_5919,N_5086);
xnor U6352 (N_6352,N_4560,N_4545);
nand U6353 (N_6353,N_5624,N_6146);
or U6354 (N_6354,N_5626,N_4085);
and U6355 (N_6355,N_5588,N_3842);
and U6356 (N_6356,N_5757,N_4612);
and U6357 (N_6357,N_3300,N_3467);
or U6358 (N_6358,N_5247,N_4913);
nor U6359 (N_6359,N_5815,N_5599);
and U6360 (N_6360,N_5958,N_4527);
nor U6361 (N_6361,N_3616,N_5532);
nor U6362 (N_6362,N_3442,N_6095);
nor U6363 (N_6363,N_3856,N_5533);
or U6364 (N_6364,N_4904,N_3563);
nand U6365 (N_6365,N_5713,N_4441);
or U6366 (N_6366,N_3619,N_5008);
and U6367 (N_6367,N_5967,N_3324);
or U6368 (N_6368,N_3361,N_5272);
and U6369 (N_6369,N_5251,N_4604);
nor U6370 (N_6370,N_6207,N_4216);
xor U6371 (N_6371,N_4611,N_3549);
xnor U6372 (N_6372,N_4654,N_6178);
and U6373 (N_6373,N_5939,N_5604);
nand U6374 (N_6374,N_3496,N_6234);
nor U6375 (N_6375,N_3661,N_5736);
nand U6376 (N_6376,N_4367,N_3349);
xnor U6377 (N_6377,N_3604,N_3692);
and U6378 (N_6378,N_3534,N_3603);
and U6379 (N_6379,N_5722,N_5237);
or U6380 (N_6380,N_5067,N_3967);
nor U6381 (N_6381,N_5877,N_4393);
and U6382 (N_6382,N_4888,N_5864);
xor U6383 (N_6383,N_3600,N_4648);
or U6384 (N_6384,N_6036,N_6057);
nand U6385 (N_6385,N_5573,N_5441);
nor U6386 (N_6386,N_4822,N_4845);
or U6387 (N_6387,N_4130,N_4844);
and U6388 (N_6388,N_5152,N_4629);
xor U6389 (N_6389,N_4228,N_5682);
xnor U6390 (N_6390,N_4978,N_5561);
or U6391 (N_6391,N_3635,N_5453);
xnor U6392 (N_6392,N_5197,N_4573);
and U6393 (N_6393,N_5819,N_5625);
and U6394 (N_6394,N_3648,N_4644);
and U6395 (N_6395,N_5646,N_5644);
xor U6396 (N_6396,N_4676,N_4515);
nor U6397 (N_6397,N_5628,N_4299);
nand U6398 (N_6398,N_6104,N_4395);
and U6399 (N_6399,N_4012,N_6106);
or U6400 (N_6400,N_6137,N_6103);
and U6401 (N_6401,N_6059,N_3362);
nand U6402 (N_6402,N_4608,N_4637);
nor U6403 (N_6403,N_4798,N_4632);
or U6404 (N_6404,N_4797,N_4261);
and U6405 (N_6405,N_4988,N_5411);
or U6406 (N_6406,N_5737,N_3895);
nand U6407 (N_6407,N_3263,N_4544);
nor U6408 (N_6408,N_3241,N_5494);
nor U6409 (N_6409,N_4581,N_3680);
nand U6410 (N_6410,N_4529,N_4742);
and U6411 (N_6411,N_3229,N_3138);
nor U6412 (N_6412,N_5516,N_5089);
or U6413 (N_6413,N_4015,N_3929);
or U6414 (N_6414,N_3387,N_4308);
nor U6415 (N_6415,N_6019,N_3850);
nand U6416 (N_6416,N_4119,N_5712);
nand U6417 (N_6417,N_3162,N_3843);
and U6418 (N_6418,N_6079,N_4833);
nor U6419 (N_6419,N_5185,N_3872);
nand U6420 (N_6420,N_4429,N_5933);
xnor U6421 (N_6421,N_3957,N_5668);
nor U6422 (N_6422,N_4643,N_6082);
xnor U6423 (N_6423,N_4156,N_5653);
nor U6424 (N_6424,N_3274,N_4257);
or U6425 (N_6425,N_4996,N_5975);
or U6426 (N_6426,N_5087,N_6001);
or U6427 (N_6427,N_4475,N_3369);
and U6428 (N_6428,N_4062,N_4728);
nor U6429 (N_6429,N_4661,N_5692);
nand U6430 (N_6430,N_5085,N_5955);
nor U6431 (N_6431,N_6201,N_5327);
nand U6432 (N_6432,N_5333,N_6063);
or U6433 (N_6433,N_3197,N_6217);
nor U6434 (N_6434,N_5775,N_5611);
nor U6435 (N_6435,N_5426,N_3152);
and U6436 (N_6436,N_5881,N_5316);
and U6437 (N_6437,N_6085,N_5288);
nor U6438 (N_6438,N_3338,N_5544);
nor U6439 (N_6439,N_3789,N_5418);
nor U6440 (N_6440,N_3390,N_3577);
and U6441 (N_6441,N_4967,N_4399);
nor U6442 (N_6442,N_6196,N_5733);
nand U6443 (N_6443,N_5155,N_5543);
xnor U6444 (N_6444,N_5768,N_5485);
xnor U6445 (N_6445,N_5121,N_3847);
nor U6446 (N_6446,N_4989,N_4309);
nor U6447 (N_6447,N_3944,N_3271);
nand U6448 (N_6448,N_3125,N_4779);
xnor U6449 (N_6449,N_3678,N_4633);
or U6450 (N_6450,N_3298,N_5341);
nand U6451 (N_6451,N_3432,N_3943);
or U6452 (N_6452,N_4704,N_5622);
nor U6453 (N_6453,N_3727,N_5927);
or U6454 (N_6454,N_3738,N_4708);
nand U6455 (N_6455,N_3990,N_5818);
nand U6456 (N_6456,N_4543,N_3468);
nand U6457 (N_6457,N_3874,N_3593);
and U6458 (N_6458,N_4950,N_5889);
nor U6459 (N_6459,N_3702,N_4445);
or U6460 (N_6460,N_3694,N_3585);
xnor U6461 (N_6461,N_5946,N_5780);
or U6462 (N_6462,N_3855,N_5157);
nor U6463 (N_6463,N_4064,N_3935);
xnor U6464 (N_6464,N_5493,N_4173);
and U6465 (N_6465,N_5725,N_5854);
and U6466 (N_6466,N_5245,N_4072);
nand U6467 (N_6467,N_4730,N_4590);
xnor U6468 (N_6468,N_5965,N_6134);
or U6469 (N_6469,N_4196,N_4325);
or U6470 (N_6470,N_6167,N_5399);
and U6471 (N_6471,N_4087,N_3624);
xor U6472 (N_6472,N_5641,N_4524);
and U6473 (N_6473,N_5904,N_5499);
xor U6474 (N_6474,N_3752,N_6020);
or U6475 (N_6475,N_5314,N_4722);
nor U6476 (N_6476,N_4615,N_3920);
and U6477 (N_6477,N_3154,N_3453);
xnor U6478 (N_6478,N_5224,N_5753);
nand U6479 (N_6479,N_5790,N_3742);
nor U6480 (N_6480,N_3544,N_5307);
or U6481 (N_6481,N_3537,N_5378);
nor U6482 (N_6482,N_6048,N_4528);
nor U6483 (N_6483,N_3755,N_3199);
nand U6484 (N_6484,N_6145,N_5739);
and U6485 (N_6485,N_4418,N_4307);
nand U6486 (N_6486,N_6028,N_5861);
nand U6487 (N_6487,N_4271,N_3866);
or U6488 (N_6488,N_6084,N_3605);
xnor U6489 (N_6489,N_5253,N_3296);
xor U6490 (N_6490,N_5460,N_3490);
or U6491 (N_6491,N_5326,N_3451);
nand U6492 (N_6492,N_5813,N_4935);
or U6493 (N_6493,N_5062,N_3717);
nand U6494 (N_6494,N_5782,N_5868);
nand U6495 (N_6495,N_4767,N_3402);
nor U6496 (N_6496,N_4416,N_4954);
or U6497 (N_6497,N_4014,N_6204);
nor U6498 (N_6498,N_4360,N_4103);
nand U6499 (N_6499,N_3858,N_4242);
or U6500 (N_6500,N_6081,N_3769);
and U6501 (N_6501,N_4582,N_3739);
xnor U6502 (N_6502,N_3501,N_3912);
xnor U6503 (N_6503,N_4564,N_5814);
nor U6504 (N_6504,N_6011,N_4371);
nand U6505 (N_6505,N_4138,N_3591);
and U6506 (N_6506,N_4131,N_6141);
and U6507 (N_6507,N_4902,N_5252);
nand U6508 (N_6508,N_5824,N_4016);
nand U6509 (N_6509,N_4781,N_5620);
and U6510 (N_6510,N_4603,N_5321);
and U6511 (N_6511,N_3970,N_3379);
and U6512 (N_6512,N_3457,N_5837);
xnor U6513 (N_6513,N_6129,N_5787);
xor U6514 (N_6514,N_4635,N_5896);
nand U6515 (N_6515,N_4069,N_4404);
and U6516 (N_6516,N_3705,N_5074);
nor U6517 (N_6517,N_5570,N_6174);
xor U6518 (N_6518,N_5360,N_4813);
nand U6519 (N_6519,N_5512,N_4720);
nand U6520 (N_6520,N_3218,N_5357);
nand U6521 (N_6521,N_3838,N_5268);
nor U6522 (N_6522,N_3191,N_3841);
nand U6523 (N_6523,N_4448,N_4470);
xor U6524 (N_6524,N_5820,N_5015);
and U6525 (N_6525,N_4319,N_4454);
and U6526 (N_6526,N_5822,N_5984);
or U6527 (N_6527,N_3620,N_5020);
xnor U6528 (N_6528,N_4758,N_5079);
and U6529 (N_6529,N_6071,N_3355);
xnor U6530 (N_6530,N_4091,N_4741);
nor U6531 (N_6531,N_4933,N_4034);
nor U6532 (N_6532,N_5634,N_3332);
or U6533 (N_6533,N_6169,N_5884);
nand U6534 (N_6534,N_5546,N_3169);
xnor U6535 (N_6535,N_5263,N_5349);
and U6536 (N_6536,N_5190,N_6040);
and U6537 (N_6537,N_4706,N_5658);
or U6538 (N_6538,N_4314,N_3293);
or U6539 (N_6539,N_3356,N_4721);
and U6540 (N_6540,N_5076,N_5829);
and U6541 (N_6541,N_5232,N_5275);
and U6542 (N_6542,N_4958,N_4641);
and U6543 (N_6543,N_5291,N_5104);
nand U6544 (N_6544,N_4421,N_4726);
xor U6545 (N_6545,N_5465,N_5594);
nand U6546 (N_6546,N_5982,N_3198);
nand U6547 (N_6547,N_5080,N_3433);
or U6548 (N_6548,N_3150,N_3597);
or U6549 (N_6549,N_4122,N_4843);
or U6550 (N_6550,N_6166,N_6030);
xnor U6551 (N_6551,N_5540,N_4780);
nor U6552 (N_6552,N_3305,N_4011);
or U6553 (N_6553,N_4032,N_5656);
nand U6554 (N_6554,N_5161,N_4268);
and U6555 (N_6555,N_3275,N_3628);
or U6556 (N_6556,N_5997,N_6076);
xnor U6557 (N_6557,N_4807,N_3547);
xnor U6558 (N_6558,N_5090,N_6144);
or U6559 (N_6559,N_4323,N_4514);
nand U6560 (N_6560,N_4795,N_5781);
xor U6561 (N_6561,N_6111,N_4941);
nand U6562 (N_6562,N_3599,N_4553);
xor U6563 (N_6563,N_6124,N_4990);
nand U6564 (N_6564,N_4235,N_3627);
xnor U6565 (N_6565,N_5070,N_5388);
nand U6566 (N_6566,N_5001,N_4177);
and U6567 (N_6567,N_3588,N_4279);
xnor U6568 (N_6568,N_4402,N_5223);
and U6569 (N_6569,N_5748,N_5772);
nor U6570 (N_6570,N_3553,N_4743);
or U6571 (N_6571,N_3947,N_4141);
nor U6572 (N_6572,N_5483,N_4058);
and U6573 (N_6573,N_5298,N_4760);
or U6574 (N_6574,N_3350,N_3489);
nand U6575 (N_6575,N_5747,N_3646);
and U6576 (N_6576,N_3745,N_5174);
and U6577 (N_6577,N_6164,N_3840);
nand U6578 (N_6578,N_3346,N_5821);
or U6579 (N_6579,N_5694,N_4566);
nor U6580 (N_6580,N_3846,N_3859);
nand U6581 (N_6581,N_6015,N_5574);
and U6582 (N_6582,N_4424,N_5510);
xnor U6583 (N_6583,N_5749,N_3601);
xor U6584 (N_6584,N_3592,N_3499);
and U6585 (N_6585,N_4818,N_6155);
or U6586 (N_6586,N_5099,N_3244);
and U6587 (N_6587,N_5332,N_4980);
nor U6588 (N_6588,N_3887,N_4053);
nor U6589 (N_6589,N_6097,N_3285);
nand U6590 (N_6590,N_4183,N_5862);
and U6591 (N_6591,N_5595,N_5687);
and U6592 (N_6592,N_3910,N_3148);
and U6593 (N_6593,N_5505,N_3710);
nand U6594 (N_6594,N_3340,N_3449);
xor U6595 (N_6595,N_6127,N_5598);
nor U6596 (N_6596,N_5906,N_3417);
nor U6597 (N_6597,N_6123,N_4232);
nand U6598 (N_6598,N_3987,N_6147);
xnor U6599 (N_6599,N_3961,N_3318);
and U6600 (N_6600,N_4971,N_5053);
nor U6601 (N_6601,N_4898,N_5226);
or U6602 (N_6602,N_5392,N_3266);
or U6603 (N_6603,N_5587,N_4801);
nand U6604 (N_6604,N_3292,N_6130);
and U6605 (N_6605,N_3896,N_4814);
and U6606 (N_6606,N_5165,N_4479);
nand U6607 (N_6607,N_4678,N_3477);
nand U6608 (N_6608,N_5631,N_3481);
or U6609 (N_6609,N_5180,N_6185);
xor U6610 (N_6610,N_4519,N_5885);
nor U6611 (N_6611,N_5206,N_5382);
and U6612 (N_6612,N_4230,N_4773);
and U6613 (N_6613,N_6175,N_5844);
nand U6614 (N_6614,N_3236,N_4892);
nand U6615 (N_6615,N_5179,N_6107);
xor U6616 (N_6616,N_5239,N_4570);
and U6617 (N_6617,N_4596,N_4302);
or U6618 (N_6618,N_4276,N_5852);
nand U6619 (N_6619,N_5627,N_6068);
xor U6620 (N_6620,N_4185,N_3398);
or U6621 (N_6621,N_3936,N_3950);
or U6622 (N_6622,N_6220,N_3135);
nor U6623 (N_6623,N_3882,N_3806);
nand U6624 (N_6624,N_4410,N_3239);
nand U6625 (N_6625,N_4060,N_6026);
nand U6626 (N_6626,N_4217,N_5222);
nor U6627 (N_6627,N_3676,N_5164);
or U6628 (N_6628,N_4838,N_5683);
xnor U6629 (N_6629,N_5066,N_5841);
xor U6630 (N_6630,N_5106,N_5233);
or U6631 (N_6631,N_4628,N_3278);
xnor U6632 (N_6632,N_4447,N_6139);
and U6633 (N_6633,N_4220,N_4374);
or U6634 (N_6634,N_3429,N_3227);
and U6635 (N_6635,N_3223,N_5913);
xor U6636 (N_6636,N_3413,N_3982);
xor U6637 (N_6637,N_5308,N_4029);
or U6638 (N_6638,N_3458,N_3826);
and U6639 (N_6639,N_3261,N_4994);
and U6640 (N_6640,N_5706,N_5582);
or U6641 (N_6641,N_4534,N_5111);
xnor U6642 (N_6642,N_5715,N_6034);
nor U6643 (N_6643,N_4229,N_3319);
or U6644 (N_6644,N_5836,N_3788);
and U6645 (N_6645,N_3818,N_5437);
nand U6646 (N_6646,N_3574,N_3482);
and U6647 (N_6647,N_4384,N_4984);
and U6648 (N_6648,N_3767,N_3723);
xor U6649 (N_6649,N_4358,N_3918);
xor U6650 (N_6650,N_5006,N_4736);
or U6651 (N_6651,N_3322,N_3884);
and U6652 (N_6652,N_5888,N_3992);
and U6653 (N_6653,N_4681,N_5947);
and U6654 (N_6654,N_5924,N_3210);
or U6655 (N_6655,N_4858,N_4121);
and U6656 (N_6656,N_5575,N_4574);
xor U6657 (N_6657,N_3253,N_3167);
nor U6658 (N_6658,N_4254,N_3822);
and U6659 (N_6659,N_5279,N_4695);
and U6660 (N_6660,N_5870,N_3875);
nor U6661 (N_6661,N_4398,N_5000);
nor U6662 (N_6662,N_5711,N_4090);
nor U6663 (N_6663,N_6236,N_4218);
or U6664 (N_6664,N_5839,N_4518);
nor U6665 (N_6665,N_3893,N_3165);
or U6666 (N_6666,N_6237,N_3258);
nand U6667 (N_6667,N_4703,N_5909);
or U6668 (N_6668,N_3704,N_4214);
xor U6669 (N_6669,N_4457,N_4381);
and U6670 (N_6670,N_4076,N_3283);
nor U6671 (N_6671,N_4042,N_6086);
nand U6672 (N_6672,N_5192,N_4655);
nor U6673 (N_6673,N_3391,N_4101);
xor U6674 (N_6674,N_4098,N_5312);
or U6675 (N_6675,N_3317,N_4097);
and U6676 (N_6676,N_3958,N_4847);
nand U6677 (N_6677,N_3321,N_4289);
nor U6678 (N_6678,N_3246,N_5583);
or U6679 (N_6679,N_5094,N_3845);
nand U6680 (N_6680,N_4198,N_4243);
xor U6681 (N_6681,N_5696,N_5718);
nand U6682 (N_6682,N_3539,N_3303);
or U6683 (N_6683,N_5433,N_5458);
and U6684 (N_6684,N_4920,N_3825);
xnor U6685 (N_6685,N_4487,N_4940);
nand U6686 (N_6686,N_4617,N_3685);
nand U6687 (N_6687,N_4199,N_5132);
or U6688 (N_6688,N_4472,N_3540);
nand U6689 (N_6689,N_4043,N_3757);
nand U6690 (N_6690,N_5709,N_5428);
or U6691 (N_6691,N_4662,N_4956);
xor U6692 (N_6692,N_4107,N_5073);
nor U6693 (N_6693,N_4482,N_5645);
or U6694 (N_6694,N_5457,N_4620);
nand U6695 (N_6695,N_4473,N_3171);
and U6696 (N_6696,N_3633,N_5531);
or U6697 (N_6697,N_3312,N_5491);
or U6698 (N_6698,N_4070,N_5567);
nor U6699 (N_6699,N_3508,N_4431);
nand U6700 (N_6700,N_5408,N_3572);
nand U6701 (N_6701,N_4598,N_5126);
and U6702 (N_6702,N_3126,N_5119);
and U6703 (N_6703,N_5557,N_4373);
nand U6704 (N_6704,N_5274,N_5334);
nor U6705 (N_6705,N_5803,N_3695);
nor U6706 (N_6706,N_3701,N_6023);
and U6707 (N_6707,N_3509,N_5315);
and U6708 (N_6708,N_5169,N_3470);
nor U6709 (N_6709,N_3775,N_4422);
nand U6710 (N_6710,N_5619,N_4129);
and U6711 (N_6711,N_3147,N_6024);
nor U6712 (N_6712,N_4250,N_5717);
or U6713 (N_6713,N_3780,N_5419);
nor U6714 (N_6714,N_4835,N_4976);
or U6715 (N_6715,N_3743,N_3792);
or U6716 (N_6716,N_5936,N_5935);
and U6717 (N_6717,N_4089,N_4831);
and U6718 (N_6718,N_4718,N_6161);
nand U6719 (N_6719,N_3339,N_3976);
and U6720 (N_6720,N_4449,N_5667);
nand U6721 (N_6721,N_5415,N_4411);
nand U6722 (N_6722,N_5723,N_3344);
nor U6723 (N_6723,N_5296,N_4075);
and U6724 (N_6724,N_3625,N_6245);
nor U6725 (N_6725,N_6003,N_4462);
nor U6726 (N_6726,N_4341,N_4536);
or U6727 (N_6727,N_3697,N_3673);
or U6728 (N_6728,N_4133,N_5665);
nor U6729 (N_6729,N_5934,N_3479);
nor U6730 (N_6730,N_5088,N_5211);
and U6731 (N_6731,N_5338,N_4267);
xnor U6732 (N_6732,N_6002,N_3360);
and U6733 (N_6733,N_3358,N_3892);
nand U6734 (N_6734,N_5110,N_5795);
nand U6735 (N_6735,N_3201,N_5843);
or U6736 (N_6736,N_5203,N_4631);
or U6737 (N_6737,N_4096,N_4348);
nand U6738 (N_6738,N_5130,N_4137);
nand U6739 (N_6739,N_3443,N_4328);
xor U6740 (N_6740,N_3216,N_4663);
xor U6741 (N_6741,N_4819,N_5082);
nor U6742 (N_6742,N_5993,N_6078);
or U6743 (N_6743,N_3240,N_5578);
xnor U6744 (N_6744,N_5964,N_5773);
nand U6745 (N_6745,N_3889,N_6053);
nand U6746 (N_6746,N_4158,N_4310);
nor U6747 (N_6747,N_5097,N_3411);
nand U6748 (N_6748,N_5014,N_3662);
nand U6749 (N_6749,N_3923,N_3153);
or U6750 (N_6750,N_4375,N_5123);
nand U6751 (N_6751,N_4538,N_4282);
xor U6752 (N_6752,N_5720,N_5591);
and U6753 (N_6753,N_5833,N_3985);
nand U6754 (N_6754,N_4713,N_4178);
nand U6755 (N_6755,N_4986,N_3431);
xor U6756 (N_6756,N_4312,N_5755);
or U6757 (N_6757,N_5636,N_3994);
nand U6758 (N_6758,N_4561,N_5365);
or U6759 (N_6759,N_3602,N_5637);
nand U6760 (N_6760,N_4711,N_3914);
nand U6761 (N_6761,N_5019,N_5470);
and U6762 (N_6762,N_5960,N_4002);
nand U6763 (N_6763,N_3804,N_5735);
or U6764 (N_6764,N_3925,N_4446);
or U6765 (N_6765,N_4587,N_4999);
nor U6766 (N_6766,N_3528,N_3819);
and U6767 (N_6767,N_4322,N_3459);
nor U6768 (N_6768,N_3415,N_5534);
and U6769 (N_6769,N_5004,N_5260);
and U6770 (N_6770,N_6008,N_3181);
xor U6771 (N_6771,N_5462,N_5873);
nand U6772 (N_6772,N_4531,N_4512);
or U6773 (N_6773,N_4377,N_3280);
and U6774 (N_6774,N_6177,N_4626);
nand U6775 (N_6775,N_5902,N_4925);
and U6776 (N_6776,N_5876,N_5900);
nor U6777 (N_6777,N_4117,N_3200);
nand U6778 (N_6778,N_4646,N_3464);
or U6779 (N_6779,N_3460,N_5537);
and U6780 (N_6780,N_5506,N_4305);
xor U6781 (N_6781,N_5700,N_4132);
xor U6782 (N_6782,N_3188,N_6136);
and U6783 (N_6783,N_5250,N_4281);
or U6784 (N_6784,N_3381,N_5439);
or U6785 (N_6785,N_5035,N_5704);
nand U6786 (N_6786,N_5745,N_3933);
and U6787 (N_6787,N_3991,N_3272);
or U6788 (N_6788,N_3485,N_4318);
nand U6789 (N_6789,N_5234,N_3983);
nand U6790 (N_6790,N_4864,N_6073);
nand U6791 (N_6791,N_3128,N_4315);
xnor U6792 (N_6792,N_5827,N_6215);
xnor U6793 (N_6793,N_3851,N_3986);
xor U6794 (N_6794,N_3488,N_5865);
and U6795 (N_6795,N_4048,N_3237);
or U6796 (N_6796,N_4247,N_4923);
nor U6797 (N_6797,N_4660,N_3587);
xnor U6798 (N_6798,N_3419,N_5227);
nor U6799 (N_6799,N_5895,N_5352);
or U6800 (N_6800,N_5596,N_4747);
and U6801 (N_6801,N_3878,N_4606);
or U6802 (N_6802,N_5949,N_5487);
or U6803 (N_6803,N_3471,N_3960);
nor U6804 (N_6804,N_3213,N_6089);
nor U6805 (N_6805,N_4916,N_5423);
and U6806 (N_6806,N_6044,N_4192);
and U6807 (N_6807,N_4998,N_5013);
nor U6808 (N_6808,N_5740,N_3813);
nor U6809 (N_6809,N_4272,N_5530);
or U6810 (N_6810,N_5010,N_4840);
nand U6811 (N_6811,N_6041,N_5509);
and U6812 (N_6812,N_5792,N_4987);
xnor U6813 (N_6813,N_3824,N_3665);
xnor U6814 (N_6814,N_3331,N_4672);
nand U6815 (N_6815,N_5134,N_5003);
nand U6816 (N_6816,N_3159,N_4008);
nand U6817 (N_6817,N_4657,N_3857);
and U6818 (N_6818,N_3219,N_5287);
xor U6819 (N_6819,N_3905,N_4280);
or U6820 (N_6820,N_3731,N_3919);
xnor U6821 (N_6821,N_3796,N_3626);
nor U6822 (N_6822,N_5771,N_3690);
xnor U6823 (N_6823,N_4221,N_5576);
nand U6824 (N_6824,N_4204,N_4423);
nor U6825 (N_6825,N_5701,N_5802);
or U6826 (N_6826,N_3450,N_3518);
nand U6827 (N_6827,N_3915,N_6142);
and U6828 (N_6828,N_3926,N_4551);
nor U6829 (N_6829,N_4213,N_5779);
or U6830 (N_6830,N_3902,N_3713);
nand U6831 (N_6831,N_4815,N_5167);
nor U6832 (N_6832,N_3316,N_3684);
and U6833 (N_6833,N_4752,N_3352);
and U6834 (N_6834,N_4580,N_5801);
or U6835 (N_6835,N_5175,N_4751);
nor U6836 (N_6836,N_4018,N_5068);
nor U6837 (N_6837,N_4406,N_6062);
xnor U6838 (N_6838,N_4882,N_6066);
xnor U6839 (N_6839,N_4968,N_3578);
nand U6840 (N_6840,N_5216,N_3820);
and U6841 (N_6841,N_6243,N_5559);
and U6842 (N_6842,N_3364,N_3311);
nor U6843 (N_6843,N_6056,N_5244);
nand U6844 (N_6844,N_5615,N_3869);
xor U6845 (N_6845,N_4051,N_4383);
xnor U6846 (N_6846,N_5071,N_5660);
and U6847 (N_6847,N_5220,N_5447);
and U6848 (N_6848,N_4554,N_5793);
nor U6849 (N_6849,N_3310,N_5666);
xor U6850 (N_6850,N_5347,N_5271);
nand U6851 (N_6851,N_5845,N_3885);
xnor U6852 (N_6852,N_5690,N_4949);
xnor U6853 (N_6853,N_3234,N_4802);
or U6854 (N_6854,N_3394,N_5048);
xnor U6855 (N_6855,N_6227,N_4771);
xnor U6856 (N_6856,N_3337,N_3308);
or U6857 (N_6857,N_3870,N_4876);
xnor U6858 (N_6858,N_3786,N_3979);
or U6859 (N_6859,N_5776,N_5649);
or U6860 (N_6860,N_6183,N_3844);
xor U6861 (N_6861,N_5897,N_5593);
nand U6862 (N_6862,N_5109,N_5995);
and U6863 (N_6863,N_3535,N_5767);
nor U6864 (N_6864,N_4350,N_5689);
xor U6865 (N_6865,N_4749,N_3584);
nand U6866 (N_6866,N_3158,N_4300);
xor U6867 (N_6867,N_4931,N_3761);
nor U6868 (N_6868,N_6115,N_3890);
nand U6869 (N_6869,N_6189,N_5856);
or U6870 (N_6870,N_4828,N_4498);
xor U6871 (N_6871,N_4205,N_6051);
and U6872 (N_6872,N_5804,N_3329);
nand U6873 (N_6873,N_5096,N_4568);
and U6874 (N_6874,N_5932,N_3289);
nor U6875 (N_6875,N_4522,N_5602);
xor U6876 (N_6876,N_4493,N_4094);
nand U6877 (N_6877,N_3839,N_6031);
xnor U6878 (N_6878,N_3636,N_4073);
nand U6879 (N_6879,N_3177,N_4263);
nand U6880 (N_6880,N_3865,N_4372);
or U6881 (N_6881,N_5041,N_3969);
nand U6882 (N_6882,N_3533,N_5784);
nand U6883 (N_6883,N_5218,N_3629);
and U6884 (N_6884,N_3380,N_4557);
nand U6885 (N_6885,N_3862,N_3984);
nand U6886 (N_6886,N_5072,N_5049);
nand U6887 (N_6887,N_3209,N_4960);
or U6888 (N_6888,N_5077,N_6170);
nor U6889 (N_6889,N_3512,N_5681);
xnor U6890 (N_6890,N_5560,N_5763);
xor U6891 (N_6891,N_5698,N_4900);
nor U6892 (N_6892,N_3781,N_5944);
nor U6893 (N_6893,N_3744,N_6232);
and U6894 (N_6894,N_4966,N_5038);
nor U6895 (N_6895,N_4036,N_5970);
nand U6896 (N_6896,N_3758,N_5515);
xor U6897 (N_6897,N_5948,N_5961);
nor U6898 (N_6898,N_4356,N_5999);
nor U6899 (N_6899,N_5507,N_3610);
or U6900 (N_6900,N_6156,N_4298);
nor U6901 (N_6901,N_4144,N_3800);
nand U6902 (N_6902,N_5808,N_3934);
xor U6903 (N_6903,N_5971,N_5210);
nand U6904 (N_6904,N_4264,N_6248);
or U6905 (N_6905,N_4513,N_5761);
nand U6906 (N_6906,N_3320,N_3273);
xnor U6907 (N_6907,N_3754,N_6180);
nand U6908 (N_6908,N_4118,N_4744);
and U6909 (N_6909,N_4093,N_5240);
nand U6910 (N_6910,N_5422,N_5794);
nand U6911 (N_6911,N_5313,N_3288);
and U6912 (N_6912,N_5350,N_3618);
or U6913 (N_6913,N_3746,N_6173);
xnor U6914 (N_6914,N_5117,N_3637);
nand U6915 (N_6915,N_4202,N_3484);
nand U6916 (N_6916,N_5355,N_5609);
nor U6917 (N_6917,N_4380,N_5131);
and U6918 (N_6918,N_5759,N_4579);
nor U6919 (N_6919,N_4509,N_6007);
and U6920 (N_6920,N_3998,N_4269);
or U6921 (N_6921,N_3807,N_4645);
nor U6922 (N_6922,N_5926,N_3397);
nand U6923 (N_6923,N_4125,N_3538);
or U6924 (N_6924,N_3196,N_5874);
or U6925 (N_6925,N_3232,N_6018);
xnor U6926 (N_6926,N_3166,N_4160);
nand U6927 (N_6927,N_5269,N_3517);
nand U6928 (N_6928,N_3712,N_4020);
nand U6929 (N_6929,N_3916,N_4420);
nor U6930 (N_6930,N_3864,N_5254);
nor U6931 (N_6931,N_5477,N_4973);
or U6932 (N_6932,N_3439,N_5769);
nand U6933 (N_6933,N_4151,N_4208);
nand U6934 (N_6934,N_3170,N_5817);
nor U6935 (N_6935,N_4346,N_5809);
and U6936 (N_6936,N_3526,N_4083);
xor U6937 (N_6937,N_3607,N_4853);
and U6938 (N_6938,N_3736,N_4452);
or U6939 (N_6939,N_4616,N_5517);
nor U6940 (N_6940,N_5978,N_5405);
xnor U6941 (N_6941,N_3975,N_4918);
and U6942 (N_6942,N_3725,N_4686);
and U6943 (N_6943,N_3357,N_3632);
xor U6944 (N_6944,N_5299,N_3613);
nor U6945 (N_6945,N_5416,N_3784);
nand U6946 (N_6946,N_5114,N_4901);
xnor U6947 (N_6947,N_3478,N_5832);
xor U6948 (N_6948,N_4150,N_4401);
or U6949 (N_6949,N_3595,N_5762);
xnor U6950 (N_6950,N_5219,N_4555);
or U6951 (N_6951,N_4754,N_3359);
and U6952 (N_6952,N_4389,N_4688);
nand U6953 (N_6953,N_3830,N_4863);
xnor U6954 (N_6954,N_4591,N_4505);
nor U6955 (N_6955,N_3282,N_5601);
xor U6956 (N_6956,N_4149,N_3566);
nor U6957 (N_6957,N_4031,N_6027);
and U6958 (N_6958,N_4258,N_5063);
nand U6959 (N_6959,N_3968,N_3911);
xor U6960 (N_6960,N_3622,N_6101);
or U6961 (N_6961,N_3336,N_5075);
nand U6962 (N_6962,N_4274,N_5040);
and U6963 (N_6963,N_4508,N_5918);
and U6964 (N_6964,N_4099,N_4057);
nand U6965 (N_6965,N_5451,N_3404);
xor U6966 (N_6966,N_4549,N_5688);
and U6967 (N_6967,N_4761,N_5142);
nor U6968 (N_6968,N_5193,N_5005);
nor U6969 (N_6969,N_4886,N_5811);
or U6970 (N_6970,N_4163,N_5430);
xor U6971 (N_6971,N_5280,N_5486);
and U6972 (N_6972,N_5482,N_5729);
xnor U6973 (N_6973,N_3334,N_3267);
xnor U6974 (N_6974,N_3374,N_3903);
and U6975 (N_6975,N_3644,N_6072);
nor U6976 (N_6976,N_3559,N_5526);
or U6977 (N_6977,N_3879,N_4811);
nand U6978 (N_6978,N_5788,N_3959);
xnor U6979 (N_6979,N_4127,N_5225);
xnor U6980 (N_6980,N_5432,N_3821);
and U6981 (N_6981,N_4735,N_6098);
nor U6982 (N_6982,N_4927,N_6143);
or U6983 (N_6983,N_6179,N_4727);
and U6984 (N_6984,N_6091,N_3269);
xor U6985 (N_6985,N_3214,N_3502);
or U6986 (N_6986,N_4100,N_4540);
nand U6987 (N_6987,N_4619,N_3594);
or U6988 (N_6988,N_4005,N_3527);
nand U6989 (N_6989,N_4981,N_6029);
or U6990 (N_6990,N_3491,N_4456);
nor U6991 (N_6991,N_5642,N_4772);
nand U6992 (N_6992,N_5317,N_6090);
or U6993 (N_6993,N_4285,N_5514);
nor U6994 (N_6994,N_4186,N_6119);
or U6995 (N_6995,N_4656,N_5708);
xnor U6996 (N_6996,N_4044,N_4465);
or U6997 (N_6997,N_5579,N_6224);
or U6998 (N_6998,N_4190,N_6096);
or U6999 (N_6999,N_5553,N_4288);
nand U7000 (N_7000,N_5584,N_4669);
xnor U7001 (N_7001,N_3711,N_6241);
nand U7002 (N_7002,N_3207,N_3230);
nor U7003 (N_7003,N_3650,N_4891);
nand U7004 (N_7004,N_6083,N_5112);
and U7005 (N_7005,N_4796,N_3963);
and U7006 (N_7006,N_6032,N_4262);
xnor U7007 (N_7007,N_3463,N_5484);
nand U7008 (N_7008,N_4658,N_5524);
nand U7009 (N_7009,N_5977,N_5659);
and U7010 (N_7010,N_5860,N_5894);
xor U7011 (N_7011,N_4504,N_4732);
nand U7012 (N_7012,N_4219,N_3951);
nor U7013 (N_7013,N_4397,N_3794);
or U7014 (N_7014,N_3899,N_4764);
xnor U7015 (N_7015,N_5992,N_4834);
xor U7016 (N_7016,N_4246,N_4701);
xnor U7017 (N_7017,N_5304,N_5282);
nor U7018 (N_7018,N_3799,N_6077);
or U7019 (N_7019,N_3651,N_6016);
xor U7020 (N_7020,N_5492,N_4689);
xor U7021 (N_7021,N_4548,N_4270);
nor U7022 (N_7022,N_3598,N_3515);
and U7023 (N_7023,N_4942,N_4856);
nor U7024 (N_7024,N_5466,N_5398);
nor U7025 (N_7025,N_5425,N_4575);
nand U7026 (N_7026,N_4789,N_4985);
nor U7027 (N_7027,N_5034,N_5166);
or U7028 (N_7028,N_3764,N_4387);
xnor U7029 (N_7029,N_6000,N_3791);
nand U7030 (N_7030,N_3424,N_3371);
nor U7031 (N_7031,N_4953,N_4460);
nor U7032 (N_7032,N_4041,N_3259);
or U7033 (N_7033,N_4652,N_6049);
nor U7034 (N_7034,N_5396,N_4455);
nand U7035 (N_7035,N_5140,N_4790);
xor U7036 (N_7036,N_4614,N_4970);
nand U7037 (N_7037,N_3953,N_5045);
xor U7038 (N_7038,N_6163,N_5760);
nand U7039 (N_7039,N_5963,N_5734);
or U7040 (N_7040,N_5607,N_5107);
and U7041 (N_7041,N_3715,N_4273);
nand U7042 (N_7042,N_5675,N_3252);
or U7043 (N_7043,N_3291,N_4225);
xnor U7044 (N_7044,N_4775,N_4388);
xnor U7045 (N_7045,N_4917,N_3436);
or U7046 (N_7046,N_5475,N_4176);
and U7047 (N_7047,N_4240,N_5379);
nor U7048 (N_7048,N_4909,N_5618);
xor U7049 (N_7049,N_5640,N_6233);
nor U7050 (N_7050,N_4241,N_4433);
and U7051 (N_7051,N_6087,N_4413);
xnor U7052 (N_7052,N_3255,N_4687);
xor U7053 (N_7053,N_5581,N_3615);
nand U7054 (N_7054,N_4291,N_3183);
nor U7055 (N_7055,N_5144,N_6131);
xor U7056 (N_7056,N_5309,N_4408);
xor U7057 (N_7057,N_3456,N_4463);
or U7058 (N_7058,N_5127,N_3341);
or U7059 (N_7059,N_3681,N_5262);
or U7060 (N_7060,N_5928,N_4396);
nand U7061 (N_7061,N_5556,N_4164);
nor U7062 (N_7062,N_3287,N_5842);
xnor U7063 (N_7063,N_3511,N_5785);
xnor U7064 (N_7064,N_5941,N_4222);
nand U7065 (N_7065,N_5141,N_5907);
nor U7066 (N_7066,N_3194,N_5329);
and U7067 (N_7067,N_4576,N_4207);
xnor U7068 (N_7068,N_3965,N_6060);
nor U7069 (N_7069,N_3643,N_3455);
nor U7070 (N_7070,N_4464,N_3823);
and U7071 (N_7071,N_4114,N_3297);
nand U7072 (N_7072,N_3137,N_5143);
xnor U7073 (N_7073,N_5903,N_5566);
or U7074 (N_7074,N_6132,N_3465);
nor U7075 (N_7075,N_6110,N_4516);
or U7076 (N_7076,N_4128,N_4143);
or U7077 (N_7077,N_6221,N_5261);
or U7078 (N_7078,N_3220,N_4379);
nand U7079 (N_7079,N_4175,N_5727);
xor U7080 (N_7080,N_5548,N_5783);
nor U7081 (N_7081,N_4024,N_4625);
and U7082 (N_7082,N_4592,N_4947);
nor U7083 (N_7083,N_4354,N_4782);
and U7084 (N_7084,N_4067,N_5265);
nor U7085 (N_7085,N_5145,N_3557);
nor U7086 (N_7086,N_4019,N_3330);
xor U7087 (N_7087,N_3671,N_4339);
or U7088 (N_7088,N_4148,N_5562);
nand U7089 (N_7089,N_4244,N_4238);
xor U7090 (N_7090,N_4890,N_4668);
nor U7091 (N_7091,N_3243,N_4237);
xor U7092 (N_7092,N_5791,N_5092);
xnor U7093 (N_7093,N_3139,N_4001);
and U7094 (N_7094,N_4808,N_3848);
nor U7095 (N_7095,N_3427,N_5917);
and U7096 (N_7096,N_5100,N_3546);
or U7097 (N_7097,N_4889,N_5680);
and U7098 (N_7098,N_3590,N_3703);
or U7099 (N_7099,N_5061,N_5409);
and U7100 (N_7100,N_5027,N_4777);
nand U7101 (N_7101,N_5159,N_4203);
nand U7102 (N_7102,N_5886,N_5545);
nor U7103 (N_7103,N_5495,N_6122);
and U7104 (N_7104,N_4106,N_5449);
and U7105 (N_7105,N_3611,N_4785);
or U7106 (N_7106,N_4113,N_3268);
xnor U7107 (N_7107,N_4206,N_3376);
and U7108 (N_7108,N_4737,N_3149);
xor U7109 (N_7109,N_3623,N_4142);
and U7110 (N_7110,N_6010,N_5916);
or U7111 (N_7111,N_3793,N_4709);
xnor U7112 (N_7112,N_5950,N_4082);
nor U7113 (N_7113,N_3173,N_5413);
nand U7114 (N_7114,N_3212,N_3897);
nand U7115 (N_7115,N_3500,N_5479);
and U7116 (N_7116,N_4523,N_4326);
xor U7117 (N_7117,N_3634,N_5032);
and U7118 (N_7118,N_3146,N_5796);
nand U7119 (N_7119,N_5098,N_5362);
nor U7120 (N_7120,N_3401,N_3801);
and U7121 (N_7121,N_6202,N_4870);
nand U7122 (N_7122,N_5281,N_4414);
or U7123 (N_7123,N_3913,N_5930);
or U7124 (N_7124,N_4820,N_5328);
nor U7125 (N_7125,N_5922,N_4520);
or U7126 (N_7126,N_6100,N_5770);
xor U7127 (N_7127,N_5209,N_4723);
nand U7128 (N_7128,N_6194,N_4914);
or U7129 (N_7129,N_5243,N_6158);
xor U7130 (N_7130,N_4227,N_6209);
or U7131 (N_7131,N_5853,N_5580);
and U7132 (N_7132,N_6014,N_3964);
xnor U7133 (N_7133,N_4333,N_4517);
nand U7134 (N_7134,N_6190,N_5292);
and U7135 (N_7135,N_3722,N_3222);
xnor U7136 (N_7136,N_4526,N_3989);
nand U7137 (N_7137,N_4731,N_4922);
and U7138 (N_7138,N_3672,N_5199);
nand U7139 (N_7139,N_3867,N_5478);
xnor U7140 (N_7140,N_4481,N_4936);
and U7141 (N_7141,N_4295,N_3304);
xor U7142 (N_7142,N_3127,N_5957);
xor U7143 (N_7143,N_6064,N_6117);
nor U7144 (N_7144,N_5702,N_3469);
or U7145 (N_7145,N_3410,N_4030);
nand U7146 (N_7146,N_3407,N_4364);
xor U7147 (N_7147,N_4108,N_4926);
or U7148 (N_7148,N_4546,N_5305);
nand U7149 (N_7149,N_6033,N_4869);
xnor U7150 (N_7150,N_4699,N_5311);
nand U7151 (N_7151,N_5346,N_3714);
or U7152 (N_7152,N_4442,N_4368);
xor U7153 (N_7153,N_3270,N_4172);
or U7154 (N_7154,N_5407,N_6198);
and U7155 (N_7155,N_4039,N_4154);
xor U7156 (N_7156,N_5875,N_5828);
nor U7157 (N_7157,N_3492,N_4542);
and U7158 (N_7158,N_3564,N_4830);
or U7159 (N_7159,N_3730,N_6070);
nor U7160 (N_7160,N_4647,N_6065);
or U7161 (N_7161,N_5979,N_5914);
nand U7162 (N_7162,N_6004,N_5987);
xor U7163 (N_7163,N_5878,N_5489);
or U7164 (N_7164,N_4541,N_4471);
or U7165 (N_7165,N_5966,N_4092);
nand U7166 (N_7166,N_5459,N_5774);
and U7167 (N_7167,N_3955,N_4571);
xnor U7168 (N_7168,N_5529,N_4038);
xnor U7169 (N_7169,N_4490,N_4969);
nor U7170 (N_7170,N_3688,N_6239);
or U7171 (N_7171,N_4249,N_4826);
and U7172 (N_7172,N_4417,N_4146);
or U7173 (N_7173,N_3718,N_4849);
xnor U7174 (N_7174,N_5318,N_4715);
or U7175 (N_7175,N_4209,N_6240);
nand U7176 (N_7176,N_3802,N_4712);
nor U7177 (N_7177,N_5855,N_4799);
xor U7178 (N_7178,N_4618,N_3414);
or U7179 (N_7179,N_3748,N_3721);
xnor U7180 (N_7180,N_4724,N_5427);
or U7181 (N_7181,N_5125,N_4682);
and U7182 (N_7182,N_4607,N_5614);
nand U7183 (N_7183,N_5617,N_5367);
and U7184 (N_7184,N_4924,N_5481);
or U7185 (N_7185,N_3829,N_3724);
nand U7186 (N_7186,N_4806,N_4056);
xnor U7187 (N_7187,N_3871,N_4734);
xnor U7188 (N_7188,N_3894,N_4182);
nand U7189 (N_7189,N_5741,N_5691);
nor U7190 (N_7190,N_3386,N_5023);
and U7191 (N_7191,N_3174,N_4521);
nand U7192 (N_7192,N_4774,N_4316);
nand U7193 (N_7193,N_3803,N_4787);
xnor U7194 (N_7194,N_3811,N_4677);
nand U7195 (N_7195,N_5044,N_5871);
xor U7196 (N_7196,N_4705,N_5882);
or U7197 (N_7197,N_3617,N_5940);
or U7198 (N_7198,N_4665,N_4337);
nand U7199 (N_7199,N_5805,N_4115);
xor U7200 (N_7200,N_3768,N_5989);
and U7201 (N_7201,N_5600,N_4211);
nor U7202 (N_7202,N_5497,N_3997);
nand U7203 (N_7203,N_5612,N_4266);
nand U7204 (N_7204,N_4725,N_3348);
and U7205 (N_7205,N_5520,N_4977);
nand U7206 (N_7206,N_5945,N_5385);
and U7207 (N_7207,N_4292,N_4327);
or U7208 (N_7208,N_5508,N_4004);
or U7209 (N_7209,N_4155,N_4698);
or U7210 (N_7210,N_5377,N_5629);
nor U7211 (N_7211,N_5424,N_3828);
xor U7212 (N_7212,N_6118,N_5335);
xor U7213 (N_7213,N_3448,N_4899);
nor U7214 (N_7214,N_6052,N_3996);
xor U7215 (N_7215,N_4278,N_4578);
nand U7216 (N_7216,N_4303,N_5571);
nor U7217 (N_7217,N_4992,N_5632);
xor U7218 (N_7218,N_6105,N_4461);
xnor U7219 (N_7219,N_4673,N_3257);
xor U7220 (N_7220,N_4439,N_5651);
nor U7221 (N_7221,N_5135,N_3814);
and U7222 (N_7222,N_5172,N_3494);
nand U7223 (N_7223,N_4052,N_5905);
xor U7224 (N_7224,N_4405,N_3542);
nor U7225 (N_7225,N_5440,N_5858);
nor U7226 (N_7226,N_4483,N_5968);
or U7227 (N_7227,N_3580,N_3917);
nand U7228 (N_7228,N_6009,N_5990);
and U7229 (N_7229,N_4167,N_5257);
xnor U7230 (N_7230,N_3805,N_4939);
nor U7231 (N_7231,N_5988,N_5671);
nor U7232 (N_7232,N_5009,N_6075);
or U7233 (N_7233,N_4577,N_6203);
nand U7234 (N_7234,N_6116,N_5438);
nor U7235 (N_7235,N_3406,N_4809);
nand U7236 (N_7236,N_4756,N_3370);
and U7237 (N_7237,N_4344,N_5420);
nand U7238 (N_7238,N_6222,N_4357);
or U7239 (N_7239,N_3383,N_5542);
xnor U7240 (N_7240,N_6181,N_3187);
and U7241 (N_7241,N_5431,N_3582);
nand U7242 (N_7242,N_6188,N_3543);
xor U7243 (N_7243,N_3773,N_3256);
xnor U7244 (N_7244,N_5319,N_6128);
or U7245 (N_7245,N_3422,N_4634);
xor U7246 (N_7246,N_5214,N_4017);
nor U7247 (N_7247,N_3189,N_5695);
nor U7248 (N_7248,N_5170,N_3353);
nor U7249 (N_7249,N_4290,N_4955);
xnor U7250 (N_7250,N_6126,N_5290);
or U7251 (N_7251,N_4874,N_3836);
or U7252 (N_7252,N_5397,N_3217);
nand U7253 (N_7253,N_5434,N_3909);
or U7254 (N_7254,N_5059,N_3368);
and U7255 (N_7255,N_3776,N_3284);
nand U7256 (N_7256,N_5181,N_3962);
nor U7257 (N_7257,N_4412,N_4755);
xnor U7258 (N_7258,N_4390,N_4565);
or U7259 (N_7259,N_4793,N_3363);
and U7260 (N_7260,N_4400,N_3208);
or U7261 (N_7261,N_5807,N_3709);
nor U7262 (N_7262,N_5358,N_4945);
or U7263 (N_7263,N_3392,N_5186);
nand U7264 (N_7264,N_6013,N_4451);
or U7265 (N_7265,N_3176,N_5472);
nand U7266 (N_7266,N_4251,N_4168);
nor U7267 (N_7267,N_5297,N_3423);
xor U7268 (N_7268,N_4136,N_5883);
nor U7269 (N_7269,N_5198,N_4088);
or U7270 (N_7270,N_6154,N_4378);
nor U7271 (N_7271,N_5133,N_4786);
and U7272 (N_7272,N_4436,N_3576);
xnor U7273 (N_7273,N_4111,N_3930);
xnor U7274 (N_7274,N_4750,N_3952);
xor U7275 (N_7275,N_5122,N_4284);
xnor U7276 (N_7276,N_4049,N_4895);
nand U7277 (N_7277,N_3570,N_6125);
nor U7278 (N_7278,N_3145,N_5686);
and U7279 (N_7279,N_3131,N_4572);
xnor U7280 (N_7280,N_3375,N_5674);
nor U7281 (N_7281,N_5083,N_4187);
nand U7282 (N_7282,N_3686,N_4556);
xnor U7283 (N_7283,N_4594,N_5136);
or U7284 (N_7284,N_3888,N_4351);
nor U7285 (N_7285,N_3797,N_5149);
xnor U7286 (N_7286,N_5648,N_4684);
nor U7287 (N_7287,N_3569,N_3180);
and U7288 (N_7288,N_3466,N_3939);
nand U7289 (N_7289,N_3365,N_6162);
and U7290 (N_7290,N_5866,N_5597);
or U7291 (N_7291,N_3384,N_3514);
or U7292 (N_7292,N_6187,N_3425);
xor U7293 (N_7293,N_4215,N_3434);
nand U7294 (N_7294,N_4296,N_4394);
or U7295 (N_7295,N_4586,N_3876);
xnor U7296 (N_7296,N_4194,N_4666);
nor U7297 (N_7297,N_6039,N_5504);
nand U7298 (N_7298,N_3735,N_4116);
or U7299 (N_7299,N_5171,N_3832);
xnor U7300 (N_7300,N_4169,N_4484);
and U7301 (N_7301,N_3974,N_3435);
nor U7302 (N_7302,N_4330,N_5887);
and U7303 (N_7303,N_4022,N_5118);
and U7304 (N_7304,N_4910,N_4867);
nor U7305 (N_7305,N_5555,N_3995);
nand U7306 (N_7306,N_4865,N_4152);
and U7307 (N_7307,N_3416,N_5011);
or U7308 (N_7308,N_4311,N_3922);
nand U7309 (N_7309,N_3927,N_5572);
or U7310 (N_7310,N_5942,N_5565);
and U7311 (N_7311,N_5752,N_5826);
nand U7312 (N_7312,N_3750,N_4500);
nor U7313 (N_7313,N_4355,N_4153);
or U7314 (N_7314,N_5029,N_4191);
and U7315 (N_7315,N_5376,N_5283);
and U7316 (N_7316,N_4200,N_5500);
nand U7317 (N_7317,N_5285,N_5238);
xor U7318 (N_7318,N_4065,N_4804);
xor U7319 (N_7319,N_4745,N_5215);
and U7320 (N_7320,N_3971,N_5138);
nor U7321 (N_7321,N_5511,N_5246);
nor U7322 (N_7322,N_4147,N_5937);
nor U7323 (N_7323,N_4223,N_5541);
xnor U7324 (N_7324,N_4938,N_4494);
xor U7325 (N_7325,N_4748,N_4964);
nor U7326 (N_7326,N_6159,N_5901);
or U7327 (N_7327,N_3679,N_4559);
or U7328 (N_7328,N_3302,N_5766);
xnor U7329 (N_7329,N_3505,N_6113);
xnor U7330 (N_7330,N_3682,N_4854);
and U7331 (N_7331,N_5925,N_3852);
xor U7332 (N_7332,N_5064,N_5474);
nand U7333 (N_7333,N_5643,N_4332);
nand U7334 (N_7334,N_3937,N_4697);
nor U7335 (N_7335,N_5182,N_4825);
nor U7336 (N_7336,N_4951,N_5456);
and U7337 (N_7337,N_3808,N_5519);
nand U7338 (N_7338,N_5513,N_3211);
nand U7339 (N_7339,N_4317,N_5521);
and U7340 (N_7340,N_3326,N_3921);
nor U7341 (N_7341,N_6099,N_5270);
or U7342 (N_7342,N_4740,N_6120);
or U7343 (N_7343,N_3510,N_5623);
nor U7344 (N_7344,N_5146,N_5446);
and U7345 (N_7345,N_3716,N_4077);
or U7346 (N_7346,N_5673,N_3281);
or U7347 (N_7347,N_5714,N_4851);
xor U7348 (N_7348,N_6182,N_4370);
and U7349 (N_7349,N_4567,N_5022);
xnor U7350 (N_7350,N_5744,N_3753);
nand U7351 (N_7351,N_4776,N_4599);
xnor U7352 (N_7352,N_5663,N_4226);
or U7353 (N_7353,N_4480,N_4047);
xnor U7354 (N_7354,N_6168,N_5951);
nand U7355 (N_7355,N_4547,N_3396);
xnor U7356 (N_7356,N_5101,N_4597);
xor U7357 (N_7357,N_3908,N_5031);
xor U7358 (N_7358,N_5310,N_3762);
or U7359 (N_7359,N_5007,N_3248);
nor U7360 (N_7360,N_4491,N_3185);
nand U7361 (N_7361,N_5650,N_5764);
xnor U7362 (N_7362,N_4023,N_3696);
xor U7363 (N_7363,N_6140,N_4878);
nand U7364 (N_7364,N_4212,N_3907);
xor U7365 (N_7365,N_5139,N_6246);
and U7366 (N_7366,N_4642,N_3568);
and U7367 (N_7367,N_4905,N_4610);
nor U7368 (N_7368,N_3523,N_4010);
nor U7369 (N_7369,N_4265,N_3333);
and U7370 (N_7370,N_6200,N_3562);
and U7371 (N_7371,N_3565,N_6225);
xor U7372 (N_7372,N_4444,N_5037);
or U7373 (N_7373,N_3966,N_5191);
nor U7374 (N_7374,N_3172,N_4975);
and U7375 (N_7375,N_5342,N_3827);
and U7376 (N_7376,N_4562,N_4440);
nand U7377 (N_7377,N_5129,N_4050);
and U7378 (N_7378,N_4248,N_5469);
xor U7379 (N_7379,N_3940,N_4234);
or U7380 (N_7380,N_3798,N_3205);
nor U7381 (N_7381,N_6046,N_3192);
xor U7382 (N_7382,N_5880,N_5455);
and U7383 (N_7383,N_5867,N_5986);
and U7384 (N_7384,N_5523,N_4409);
nor U7385 (N_7385,N_5105,N_5340);
nand U7386 (N_7386,N_3606,N_4595);
and U7387 (N_7387,N_5444,N_3264);
nand U7388 (N_7388,N_5039,N_4829);
nor U7389 (N_7389,N_3945,N_3395);
and U7390 (N_7390,N_3323,N_4245);
or U7391 (N_7391,N_5391,N_5879);
xor U7392 (N_7392,N_4071,N_3900);
nor U7393 (N_7393,N_3931,N_3698);
nand U7394 (N_7394,N_3254,N_5356);
xnor U7395 (N_7395,N_5657,N_5496);
nand U7396 (N_7396,N_4636,N_5323);
and U7397 (N_7397,N_3729,N_4872);
or U7398 (N_7398,N_5525,N_5200);
xnor U7399 (N_7399,N_5343,N_5081);
nor U7400 (N_7400,N_4054,N_4685);
and U7401 (N_7401,N_4193,N_5160);
or U7402 (N_7402,N_4425,N_3664);
and U7403 (N_7403,N_5652,N_6080);
nor U7404 (N_7404,N_5558,N_4026);
nor U7405 (N_7405,N_6230,N_3454);
or U7406 (N_7406,N_4362,N_3978);
xnor U7407 (N_7407,N_5577,N_4286);
and U7408 (N_7408,N_5589,N_4558);
nor U7409 (N_7409,N_4601,N_3313);
and U7410 (N_7410,N_4983,N_4707);
nand U7411 (N_7411,N_4124,N_4859);
nand U7412 (N_7412,N_4079,N_4095);
xor U7413 (N_7413,N_3367,N_3151);
and U7414 (N_7414,N_3860,N_5091);
or U7415 (N_7415,N_3325,N_3732);
nand U7416 (N_7416,N_4376,N_5322);
nand U7417 (N_7417,N_3461,N_5838);
xor U7418 (N_7418,N_5386,N_4415);
or U7419 (N_7419,N_6135,N_4887);
and U7420 (N_7420,N_4877,N_4477);
and U7421 (N_7421,N_5716,N_5345);
nand U7422 (N_7422,N_4857,N_3883);
xnor U7423 (N_7423,N_4359,N_3314);
and U7424 (N_7424,N_3493,N_5830);
nor U7425 (N_7425,N_3938,N_3179);
or U7426 (N_7426,N_6229,N_5799);
nand U7427 (N_7427,N_3536,N_5371);
nand U7428 (N_7428,N_5113,N_3707);
and U7429 (N_7429,N_5442,N_5221);
xor U7430 (N_7430,N_4794,N_3583);
or U7431 (N_7431,N_4033,N_3640);
and U7432 (N_7432,N_5018,N_6249);
or U7433 (N_7433,N_3204,N_3444);
or U7434 (N_7434,N_4602,N_4126);
nor U7435 (N_7435,N_4496,N_4792);
xor U7436 (N_7436,N_6244,N_4810);
nor U7437 (N_7437,N_5344,N_5195);
or U7438 (N_7438,N_3224,N_3132);
and U7439 (N_7439,N_4453,N_4159);
nand U7440 (N_7440,N_3420,N_6193);
or U7441 (N_7441,N_4382,N_4080);
xnor U7442 (N_7442,N_3751,N_5816);
xor U7443 (N_7443,N_5373,N_4694);
xor U7444 (N_7444,N_3351,N_5162);
and U7445 (N_7445,N_5983,N_5806);
nand U7446 (N_7446,N_3142,N_6093);
or U7447 (N_7447,N_5204,N_4120);
xnor U7448 (N_7448,N_3342,N_5664);
xor U7449 (N_7449,N_3977,N_5084);
or U7450 (N_7450,N_3206,N_5503);
nor U7451 (N_7451,N_3164,N_3265);
xnor U7452 (N_7452,N_3747,N_4338);
nand U7453 (N_7453,N_3774,N_3134);
and U7454 (N_7454,N_5188,N_4391);
or U7455 (N_7455,N_4674,N_3418);
xor U7456 (N_7456,N_4166,N_5672);
nand U7457 (N_7457,N_3524,N_5539);
or U7458 (N_7458,N_4253,N_3691);
and U7459 (N_7459,N_6121,N_3728);
nand U7460 (N_7460,N_4059,N_5248);
nand U7461 (N_7461,N_4817,N_3639);
or U7462 (N_7462,N_4352,N_4836);
xor U7463 (N_7463,N_4428,N_4539);
and U7464 (N_7464,N_5028,N_4007);
and U7465 (N_7465,N_5603,N_4868);
or U7466 (N_7466,N_5294,N_3409);
xnor U7467 (N_7467,N_5151,N_4003);
or U7468 (N_7468,N_5366,N_3203);
nand U7469 (N_7469,N_3706,N_5036);
or U7470 (N_7470,N_4861,N_4769);
nand U7471 (N_7471,N_5605,N_4906);
nor U7472 (N_7472,N_6021,N_4345);
or U7473 (N_7473,N_5699,N_5429);
nand U7474 (N_7474,N_6088,N_5368);
nor U7475 (N_7475,N_5899,N_5825);
or U7476 (N_7476,N_3765,N_5585);
and U7477 (N_7477,N_3756,N_4489);
nor U7478 (N_7478,N_5476,N_5017);
xnor U7479 (N_7479,N_4907,N_5336);
nand U7480 (N_7480,N_5991,N_3554);
and U7481 (N_7481,N_4552,N_5406);
xnor U7482 (N_7482,N_5231,N_5163);
nand U7483 (N_7483,N_3399,N_5380);
xor U7484 (N_7484,N_4335,N_5670);
and U7485 (N_7485,N_4979,N_4778);
and U7486 (N_7486,N_4717,N_5630);
nor U7487 (N_7487,N_6108,N_4363);
and U7488 (N_7488,N_3837,N_5213);
or U7489 (N_7489,N_5464,N_6208);
nor U7490 (N_7490,N_3904,N_4827);
and U7491 (N_7491,N_4365,N_4921);
xor U7492 (N_7492,N_3666,N_4982);
or U7493 (N_7493,N_6042,N_5751);
and U7494 (N_7494,N_5401,N_3668);
nor U7495 (N_7495,N_3382,N_6165);
nand U7496 (N_7496,N_6218,N_5052);
or U7497 (N_7497,N_6151,N_4664);
nor U7498 (N_7498,N_5592,N_5306);
and U7499 (N_7499,N_4435,N_4640);
and U7500 (N_7500,N_3849,N_5685);
xnor U7501 (N_7501,N_6069,N_6231);
or U7502 (N_7502,N_4716,N_4691);
or U7503 (N_7503,N_3522,N_4342);
or U7504 (N_7504,N_4188,N_3249);
nor U7505 (N_7505,N_5962,N_6186);
nor U7506 (N_7506,N_3250,N_4506);
or U7507 (N_7507,N_6074,N_3393);
or U7508 (N_7508,N_5473,N_3942);
or U7509 (N_7509,N_3445,N_6205);
nor U7510 (N_7510,N_5046,N_5931);
nor U7511 (N_7511,N_6112,N_5375);
nand U7512 (N_7512,N_4165,N_3408);
or U7513 (N_7513,N_5621,N_4343);
and U7514 (N_7514,N_3541,N_5364);
xnor U7515 (N_7515,N_5502,N_3299);
and U7516 (N_7516,N_5295,N_5452);
and U7517 (N_7517,N_3247,N_4850);
xor U7518 (N_7518,N_3654,N_5719);
or U7519 (N_7519,N_5183,N_5608);
or U7520 (N_7520,N_4112,N_3438);
nor U7521 (N_7521,N_5148,N_4589);
and U7522 (N_7522,N_5893,N_4293);
xnor U7523 (N_7523,N_4959,N_5661);
nor U7524 (N_7524,N_3778,N_3242);
and U7525 (N_7525,N_3596,N_4530);
nor U7526 (N_7526,N_4693,N_3262);
or U7527 (N_7527,N_4171,N_3586);
nor U7528 (N_7528,N_4855,N_5635);
nand U7529 (N_7529,N_6219,N_4161);
xnor U7530 (N_7530,N_6152,N_6047);
nor U7531 (N_7531,N_3782,N_3377);
and U7532 (N_7532,N_6094,N_3186);
nand U7533 (N_7533,N_3156,N_4063);
nor U7534 (N_7534,N_5065,N_4081);
nand U7535 (N_7535,N_5156,N_4392);
and U7536 (N_7536,N_5374,N_4805);
xor U7537 (N_7537,N_5278,N_3737);
nand U7538 (N_7538,N_5467,N_4329);
nand U7539 (N_7539,N_3521,N_3552);
or U7540 (N_7540,N_4600,N_5613);
xor U7541 (N_7541,N_5054,N_3556);
or U7542 (N_7542,N_3388,N_3530);
nand U7543 (N_7543,N_4746,N_5043);
and U7544 (N_7544,N_3195,N_5798);
nor U7545 (N_7545,N_5057,N_4624);
and U7546 (N_7546,N_5153,N_4783);
nand U7547 (N_7547,N_5069,N_3579);
nor U7548 (N_7548,N_5726,N_5732);
nor U7549 (N_7549,N_4006,N_3560);
nand U7550 (N_7550,N_4622,N_5050);
and U7551 (N_7551,N_5564,N_4585);
nand U7552 (N_7552,N_3133,N_3891);
xor U7553 (N_7553,N_4438,N_5707);
nor U7554 (N_7554,N_4140,N_4821);
or U7555 (N_7555,N_5728,N_5021);
and U7556 (N_7556,N_5264,N_5756);
and U7557 (N_7557,N_4474,N_6109);
or U7558 (N_7558,N_3231,N_5677);
nand U7559 (N_7559,N_4837,N_3129);
xnor U7560 (N_7560,N_5389,N_5746);
nand U7561 (N_7561,N_5812,N_5777);
and U7562 (N_7562,N_4630,N_3790);
or U7563 (N_7563,N_5228,N_4937);
nand U7564 (N_7564,N_5973,N_4696);
or U7565 (N_7565,N_3513,N_4627);
nor U7566 (N_7566,N_5277,N_3525);
xor U7567 (N_7567,N_5518,N_4537);
nand U7568 (N_7568,N_4957,N_4875);
and U7569 (N_7569,N_5463,N_4670);
nor U7570 (N_7570,N_5953,N_6022);
nor U7571 (N_7571,N_3279,N_3245);
xnor U7572 (N_7572,N_3817,N_5255);
nand U7573 (N_7573,N_5834,N_5569);
or U7574 (N_7574,N_5848,N_5025);
and U7575 (N_7575,N_6006,N_5754);
nor U7576 (N_7576,N_6214,N_5403);
or U7577 (N_7577,N_5436,N_4879);
nor U7578 (N_7578,N_5012,N_3687);
nor U7579 (N_7579,N_5831,N_4683);
xor U7580 (N_7580,N_5369,N_5124);
and U7581 (N_7581,N_4297,N_4467);
xnor U7582 (N_7582,N_4952,N_5638);
and U7583 (N_7583,N_6067,N_6035);
nand U7584 (N_7584,N_5229,N_5024);
xnor U7585 (N_7585,N_5710,N_4287);
and U7586 (N_7586,N_3405,N_4313);
xnor U7587 (N_7587,N_5176,N_5435);
nor U7588 (N_7588,N_4502,N_4074);
xor U7589 (N_7589,N_4492,N_3766);
and U7590 (N_7590,N_5742,N_5410);
and U7591 (N_7591,N_3486,N_3307);
nand U7592 (N_7592,N_5488,N_3462);
nor U7593 (N_7593,N_4532,N_4145);
nor U7594 (N_7594,N_4347,N_4897);
or U7595 (N_7595,N_4569,N_5911);
xnor U7596 (N_7596,N_3693,N_5789);
and U7597 (N_7597,N_4324,N_4739);
nor U7598 (N_7598,N_4184,N_5797);
or U7599 (N_7599,N_5303,N_4623);
nand U7600 (N_7600,N_3763,N_3184);
nor U7601 (N_7601,N_4550,N_5535);
or U7602 (N_7602,N_5851,N_4239);
nand U7603 (N_7603,N_4252,N_4962);
nor U7604 (N_7604,N_4334,N_6195);
nor U7605 (N_7605,N_6038,N_4189);
xnor U7606 (N_7606,N_3949,N_4485);
and U7607 (N_7607,N_3689,N_4369);
or U7608 (N_7608,N_3835,N_6242);
or U7609 (N_7609,N_5721,N_5384);
and U7610 (N_7610,N_5959,N_5016);
or U7611 (N_7611,N_3809,N_4679);
nand U7612 (N_7612,N_4841,N_5568);
nor U7613 (N_7613,N_3519,N_5471);
nor U7614 (N_7614,N_4659,N_4583);
or U7615 (N_7615,N_5289,N_4459);
nand U7616 (N_7616,N_4974,N_3531);
nand U7617 (N_7617,N_5857,N_4260);
nand U7618 (N_7618,N_4816,N_3328);
and U7619 (N_7619,N_5923,N_3677);
or U7620 (N_7620,N_5194,N_4195);
nor U7621 (N_7621,N_5590,N_5835);
or U7622 (N_7622,N_6235,N_4201);
and U7623 (N_7623,N_4174,N_4511);
xor U7624 (N_7624,N_6212,N_4109);
nor U7625 (N_7625,N_5320,N_5128);
or U7626 (N_7626,N_5980,N_4824);
or U7627 (N_7627,N_3667,N_4765);
and U7628 (N_7628,N_4495,N_5337);
and U7629 (N_7629,N_5547,N_6228);
or U7630 (N_7630,N_6148,N_5892);
nor U7631 (N_7631,N_3873,N_5662);
nor U7632 (N_7632,N_3476,N_4766);
and U7633 (N_7633,N_4997,N_3631);
and U7634 (N_7634,N_4430,N_5679);
nor U7635 (N_7635,N_3366,N_5207);
or U7636 (N_7636,N_3235,N_5676);
xnor U7637 (N_7637,N_4301,N_3740);
xor U7638 (N_7638,N_6017,N_4690);
xor U7639 (N_7639,N_4702,N_5956);
xor U7640 (N_7640,N_5891,N_3504);
and U7641 (N_7641,N_5847,N_5448);
and U7642 (N_7642,N_5606,N_5954);
nor U7643 (N_7643,N_5404,N_4871);
xnor U7644 (N_7644,N_5738,N_3630);
xnor U7645 (N_7645,N_4912,N_3658);
or U7646 (N_7646,N_3655,N_5120);
or U7647 (N_7647,N_3294,N_5387);
nand U7648 (N_7648,N_3663,N_5778);
nand U7649 (N_7649,N_5461,N_3812);
nand U7650 (N_7650,N_3785,N_3306);
and U7651 (N_7651,N_4896,N_3700);
nor U7652 (N_7652,N_5976,N_5929);
or U7653 (N_7653,N_3571,N_4407);
nand U7654 (N_7654,N_5302,N_3589);
nor U7655 (N_7655,N_4157,N_4584);
xor U7656 (N_7656,N_3614,N_5846);
nand U7657 (N_7657,N_3506,N_6157);
xor U7658 (N_7658,N_5974,N_5361);
xnor U7659 (N_7659,N_5563,N_5276);
and U7660 (N_7660,N_3473,N_4035);
and U7661 (N_7661,N_4259,N_4134);
nand U7662 (N_7662,N_3550,N_3290);
or U7663 (N_7663,N_4123,N_3260);
and U7664 (N_7664,N_4170,N_5201);
nand U7665 (N_7665,N_3507,N_4181);
xnor U7666 (N_7666,N_4823,N_3669);
nand U7667 (N_7667,N_3372,N_5184);
or U7668 (N_7668,N_5655,N_4349);
and U7669 (N_7669,N_3315,N_5412);
and U7670 (N_7670,N_5527,N_3277);
or U7671 (N_7671,N_3373,N_3657);
xnor U7672 (N_7672,N_5898,N_3529);
nand U7673 (N_7673,N_5002,N_5108);
nor U7674 (N_7674,N_5705,N_4762);
or U7675 (N_7675,N_5324,N_4466);
and U7676 (N_7676,N_5363,N_6199);
and U7677 (N_7677,N_6025,N_4437);
and U7678 (N_7678,N_5154,N_4046);
nand U7679 (N_7679,N_4256,N_3954);
xnor U7680 (N_7680,N_3656,N_6223);
nand U7681 (N_7681,N_5147,N_4880);
and U7682 (N_7682,N_3720,N_4692);
nand U7683 (N_7683,N_3225,N_3770);
and U7684 (N_7684,N_4862,N_5348);
nand U7685 (N_7685,N_4321,N_4231);
and U7686 (N_7686,N_3708,N_4427);
xnor U7687 (N_7687,N_5528,N_4784);
or U7688 (N_7688,N_4535,N_5402);
nor U7689 (N_7689,N_3495,N_3327);
and U7690 (N_7690,N_3548,N_4336);
xnor U7691 (N_7691,N_4507,N_4320);
xor U7692 (N_7692,N_6102,N_3853);
and U7693 (N_7693,N_4943,N_4757);
or U7694 (N_7694,N_5284,N_3545);
nor U7695 (N_7695,N_4759,N_4210);
and U7696 (N_7696,N_5102,N_5765);
or U7697 (N_7697,N_4873,N_4386);
nor U7698 (N_7698,N_5293,N_4486);
and U7699 (N_7699,N_6216,N_4478);
nor U7700 (N_7700,N_3155,N_5536);
and U7701 (N_7701,N_4403,N_4385);
nor U7702 (N_7702,N_4110,N_5217);
xor U7703 (N_7703,N_3898,N_5383);
or U7704 (N_7704,N_3948,N_3221);
xor U7705 (N_7705,N_5693,N_6172);
nor U7706 (N_7706,N_4450,N_5952);
xor U7707 (N_7707,N_5353,N_3238);
or U7708 (N_7708,N_5058,N_4860);
or U7709 (N_7709,N_5750,N_4852);
nand U7710 (N_7710,N_3612,N_5724);
nand U7711 (N_7711,N_5301,N_4443);
or U7712 (N_7712,N_3638,N_5654);
xnor U7713 (N_7713,N_3567,N_5273);
nand U7714 (N_7714,N_4605,N_3772);
and U7715 (N_7715,N_3228,N_3157);
nand U7716 (N_7716,N_5400,N_3301);
or U7717 (N_7717,N_3880,N_5554);
nor U7718 (N_7718,N_5850,N_5056);
nand U7719 (N_7719,N_4476,N_3683);
nor U7720 (N_7720,N_5996,N_3503);
nand U7721 (N_7721,N_5550,N_5330);
nor U7722 (N_7722,N_4908,N_3144);
and U7723 (N_7723,N_3999,N_4563);
and U7724 (N_7724,N_4025,N_4045);
and U7725 (N_7725,N_4972,N_5351);
and U7726 (N_7726,N_5331,N_5703);
and U7727 (N_7727,N_5421,N_3175);
and U7728 (N_7728,N_4883,N_3573);
nor U7729 (N_7729,N_3345,N_5910);
or U7730 (N_7730,N_3430,N_6171);
xnor U7731 (N_7731,N_5678,N_6247);
or U7732 (N_7732,N_5115,N_5450);
xor U7733 (N_7733,N_3136,N_4842);
or U7734 (N_7734,N_3441,N_5669);
xnor U7735 (N_7735,N_3881,N_4028);
nor U7736 (N_7736,N_4763,N_5915);
nand U7737 (N_7737,N_3202,N_3726);
and U7738 (N_7738,N_3551,N_5731);
nand U7739 (N_7739,N_3487,N_3575);
xnor U7740 (N_7740,N_6054,N_4812);
and U7741 (N_7741,N_4066,N_4714);
nor U7742 (N_7742,N_6114,N_6138);
or U7743 (N_7743,N_5230,N_4283);
and U7744 (N_7744,N_3581,N_6206);
xnor U7745 (N_7745,N_4800,N_3886);
or U7746 (N_7746,N_5372,N_5241);
nor U7747 (N_7747,N_4893,N_4946);
nor U7748 (N_7748,N_4593,N_3143);
nand U7749 (N_7749,N_3354,N_6184);
or U7750 (N_7750,N_5552,N_6150);
nand U7751 (N_7751,N_4104,N_4963);
and U7752 (N_7752,N_5938,N_5205);
nor U7753 (N_7753,N_5849,N_3498);
or U7754 (N_7754,N_5912,N_4944);
or U7755 (N_7755,N_4353,N_3335);
nand U7756 (N_7756,N_5256,N_5758);
nor U7757 (N_7757,N_3226,N_5116);
or U7758 (N_7758,N_5202,N_6005);
or U7759 (N_7759,N_4911,N_6213);
nand U7760 (N_7760,N_3652,N_3932);
and U7761 (N_7761,N_4510,N_5394);
xnor U7762 (N_7762,N_6149,N_5445);
or U7763 (N_7763,N_5908,N_5859);
or U7764 (N_7764,N_3215,N_4037);
or U7765 (N_7765,N_4671,N_4135);
nand U7766 (N_7766,N_5810,N_6197);
or U7767 (N_7767,N_5943,N_4680);
nand U7768 (N_7768,N_5468,N_6133);
and U7769 (N_7769,N_4609,N_4419);
nand U7770 (N_7770,N_3347,N_4086);
nor U7771 (N_7771,N_5208,N_5033);
and U7772 (N_7772,N_3783,N_4932);
or U7773 (N_7773,N_3516,N_3928);
nand U7774 (N_7774,N_5786,N_5969);
and U7775 (N_7775,N_3863,N_4651);
nand U7776 (N_7776,N_5047,N_3734);
or U7777 (N_7777,N_4236,N_4497);
and U7778 (N_7778,N_4224,N_5267);
and U7779 (N_7779,N_3532,N_6238);
and U7780 (N_7780,N_5103,N_3749);
nand U7781 (N_7781,N_4061,N_5921);
xnor U7782 (N_7782,N_3981,N_3946);
xor U7783 (N_7783,N_3160,N_3378);
xnor U7784 (N_7784,N_5093,N_4929);
nor U7785 (N_7785,N_5060,N_4255);
nor U7786 (N_7786,N_3621,N_6176);
and U7787 (N_7787,N_5610,N_5187);
xor U7788 (N_7788,N_6226,N_4304);
nor U7789 (N_7789,N_4667,N_4501);
nor U7790 (N_7790,N_3760,N_4639);
and U7791 (N_7791,N_4961,N_5395);
xor U7792 (N_7792,N_3447,N_4084);
or U7793 (N_7793,N_3178,N_3810);
or U7794 (N_7794,N_4488,N_3141);
xor U7795 (N_7795,N_3182,N_3472);
or U7796 (N_7796,N_5030,N_3719);
nor U7797 (N_7797,N_3130,N_3251);
nor U7798 (N_7798,N_4675,N_3440);
or U7799 (N_7799,N_5177,N_5258);
nand U7800 (N_7800,N_6191,N_5633);
or U7801 (N_7801,N_3647,N_5325);
or U7802 (N_7802,N_3403,N_6192);
nand U7803 (N_7803,N_6058,N_4340);
nand U7804 (N_7804,N_5173,N_4009);
or U7805 (N_7805,N_4885,N_3660);
nor U7806 (N_7806,N_4162,N_3816);
or U7807 (N_7807,N_3861,N_4275);
or U7808 (N_7808,N_5586,N_3941);
nand U7809 (N_7809,N_3190,N_6043);
nand U7810 (N_7810,N_5863,N_5981);
and U7811 (N_7811,N_5454,N_5414);
nor U7812 (N_7812,N_4934,N_3933);
nand U7813 (N_7813,N_3661,N_3392);
and U7814 (N_7814,N_4500,N_5241);
nand U7815 (N_7815,N_5630,N_3690);
nor U7816 (N_7816,N_3493,N_4112);
xnor U7817 (N_7817,N_4625,N_5263);
or U7818 (N_7818,N_6060,N_4855);
or U7819 (N_7819,N_3303,N_4474);
nand U7820 (N_7820,N_4831,N_4020);
nor U7821 (N_7821,N_6181,N_5889);
nand U7822 (N_7822,N_4635,N_4324);
and U7823 (N_7823,N_3708,N_3920);
or U7824 (N_7824,N_5301,N_4217);
or U7825 (N_7825,N_3211,N_5667);
xor U7826 (N_7826,N_6136,N_4663);
or U7827 (N_7827,N_5877,N_4418);
xor U7828 (N_7828,N_4094,N_3141);
and U7829 (N_7829,N_5974,N_4733);
or U7830 (N_7830,N_6132,N_4274);
xor U7831 (N_7831,N_5683,N_4249);
or U7832 (N_7832,N_3675,N_4749);
xnor U7833 (N_7833,N_3765,N_4948);
xnor U7834 (N_7834,N_4604,N_3662);
xor U7835 (N_7835,N_3991,N_5531);
and U7836 (N_7836,N_5322,N_6215);
nand U7837 (N_7837,N_3781,N_4698);
or U7838 (N_7838,N_5114,N_4082);
and U7839 (N_7839,N_4579,N_5465);
and U7840 (N_7840,N_4384,N_3378);
nand U7841 (N_7841,N_3382,N_4597);
nor U7842 (N_7842,N_5162,N_4135);
nand U7843 (N_7843,N_4618,N_5030);
and U7844 (N_7844,N_3934,N_4768);
or U7845 (N_7845,N_4041,N_5212);
xnor U7846 (N_7846,N_6191,N_6117);
or U7847 (N_7847,N_4570,N_5937);
nand U7848 (N_7848,N_3978,N_6033);
and U7849 (N_7849,N_5051,N_3575);
or U7850 (N_7850,N_3204,N_5538);
nor U7851 (N_7851,N_3590,N_3626);
nand U7852 (N_7852,N_6244,N_5176);
nand U7853 (N_7853,N_4172,N_4931);
nor U7854 (N_7854,N_4100,N_5265);
nand U7855 (N_7855,N_5407,N_6073);
nand U7856 (N_7856,N_4322,N_3143);
or U7857 (N_7857,N_5386,N_5091);
nor U7858 (N_7858,N_5666,N_3856);
nor U7859 (N_7859,N_5314,N_4556);
nor U7860 (N_7860,N_4967,N_4592);
xor U7861 (N_7861,N_4230,N_4303);
xnor U7862 (N_7862,N_4543,N_3208);
or U7863 (N_7863,N_5017,N_4876);
or U7864 (N_7864,N_3407,N_3784);
xnor U7865 (N_7865,N_3488,N_3616);
xor U7866 (N_7866,N_5995,N_4412);
nor U7867 (N_7867,N_5044,N_6160);
or U7868 (N_7868,N_4997,N_4294);
or U7869 (N_7869,N_5738,N_5175);
nand U7870 (N_7870,N_3377,N_5013);
nor U7871 (N_7871,N_6160,N_5792);
xor U7872 (N_7872,N_3609,N_4589);
and U7873 (N_7873,N_3715,N_3335);
and U7874 (N_7874,N_4404,N_3658);
or U7875 (N_7875,N_4745,N_3947);
xor U7876 (N_7876,N_5971,N_5398);
xnor U7877 (N_7877,N_5488,N_4151);
nor U7878 (N_7878,N_5582,N_3931);
nand U7879 (N_7879,N_5948,N_5504);
xor U7880 (N_7880,N_4703,N_3290);
xor U7881 (N_7881,N_4828,N_4267);
xnor U7882 (N_7882,N_4484,N_5246);
nor U7883 (N_7883,N_5359,N_4335);
and U7884 (N_7884,N_4362,N_4200);
nor U7885 (N_7885,N_3600,N_3466);
nor U7886 (N_7886,N_4469,N_6119);
nand U7887 (N_7887,N_3318,N_5353);
and U7888 (N_7888,N_4448,N_5106);
nor U7889 (N_7889,N_5378,N_5937);
and U7890 (N_7890,N_3691,N_3215);
nor U7891 (N_7891,N_4512,N_3446);
and U7892 (N_7892,N_4174,N_5102);
or U7893 (N_7893,N_3626,N_3886);
xor U7894 (N_7894,N_6048,N_5350);
xor U7895 (N_7895,N_3235,N_5518);
and U7896 (N_7896,N_4536,N_4486);
nand U7897 (N_7897,N_4508,N_3422);
nor U7898 (N_7898,N_5332,N_5761);
and U7899 (N_7899,N_3365,N_4648);
xor U7900 (N_7900,N_4471,N_3343);
nand U7901 (N_7901,N_4797,N_3146);
nand U7902 (N_7902,N_3179,N_5353);
nand U7903 (N_7903,N_4339,N_5963);
and U7904 (N_7904,N_5823,N_5374);
xnor U7905 (N_7905,N_3812,N_5952);
and U7906 (N_7906,N_5419,N_5810);
nor U7907 (N_7907,N_4130,N_4309);
nand U7908 (N_7908,N_3754,N_4452);
nand U7909 (N_7909,N_5203,N_3920);
or U7910 (N_7910,N_5286,N_3685);
nor U7911 (N_7911,N_5032,N_6221);
and U7912 (N_7912,N_3529,N_6182);
nor U7913 (N_7913,N_3644,N_4807);
and U7914 (N_7914,N_3710,N_3497);
nand U7915 (N_7915,N_6010,N_5161);
nor U7916 (N_7916,N_4091,N_4556);
nand U7917 (N_7917,N_5439,N_3974);
nor U7918 (N_7918,N_6061,N_6163);
or U7919 (N_7919,N_3193,N_3933);
xnor U7920 (N_7920,N_4415,N_3914);
xor U7921 (N_7921,N_3579,N_4947);
or U7922 (N_7922,N_4633,N_6185);
xor U7923 (N_7923,N_5405,N_3305);
nor U7924 (N_7924,N_3126,N_3396);
or U7925 (N_7925,N_4383,N_4676);
nand U7926 (N_7926,N_4995,N_3435);
or U7927 (N_7927,N_4083,N_5005);
nand U7928 (N_7928,N_5866,N_5233);
xor U7929 (N_7929,N_5038,N_4147);
nor U7930 (N_7930,N_5843,N_4319);
and U7931 (N_7931,N_3312,N_5379);
nor U7932 (N_7932,N_4640,N_3980);
nor U7933 (N_7933,N_5515,N_5680);
or U7934 (N_7934,N_5737,N_4121);
nand U7935 (N_7935,N_3659,N_5795);
or U7936 (N_7936,N_3895,N_5332);
nand U7937 (N_7937,N_6139,N_6211);
or U7938 (N_7938,N_5536,N_5182);
and U7939 (N_7939,N_6094,N_4002);
or U7940 (N_7940,N_4151,N_4910);
or U7941 (N_7941,N_3672,N_3151);
nand U7942 (N_7942,N_4229,N_4885);
and U7943 (N_7943,N_3703,N_3533);
nand U7944 (N_7944,N_3379,N_5915);
xor U7945 (N_7945,N_3596,N_6186);
xnor U7946 (N_7946,N_6106,N_5188);
nor U7947 (N_7947,N_4291,N_3628);
nor U7948 (N_7948,N_6117,N_6085);
nor U7949 (N_7949,N_3187,N_3364);
nand U7950 (N_7950,N_3783,N_3986);
xor U7951 (N_7951,N_5717,N_4118);
and U7952 (N_7952,N_5509,N_5678);
nor U7953 (N_7953,N_5853,N_3552);
nor U7954 (N_7954,N_6236,N_5681);
xor U7955 (N_7955,N_3461,N_3694);
or U7956 (N_7956,N_4812,N_4187);
and U7957 (N_7957,N_4234,N_3674);
and U7958 (N_7958,N_4097,N_5509);
or U7959 (N_7959,N_3265,N_5182);
xor U7960 (N_7960,N_3423,N_3711);
or U7961 (N_7961,N_3242,N_5800);
and U7962 (N_7962,N_5599,N_5943);
or U7963 (N_7963,N_5276,N_3860);
or U7964 (N_7964,N_5304,N_5496);
nor U7965 (N_7965,N_5341,N_3872);
nor U7966 (N_7966,N_4481,N_5142);
or U7967 (N_7967,N_4622,N_4203);
xor U7968 (N_7968,N_5799,N_4712);
or U7969 (N_7969,N_3186,N_3645);
or U7970 (N_7970,N_5543,N_6242);
nand U7971 (N_7971,N_4310,N_4808);
nor U7972 (N_7972,N_5658,N_4167);
and U7973 (N_7973,N_3970,N_4194);
xor U7974 (N_7974,N_5594,N_4042);
nand U7975 (N_7975,N_4065,N_3217);
xnor U7976 (N_7976,N_5369,N_3258);
nand U7977 (N_7977,N_3443,N_4569);
nand U7978 (N_7978,N_4312,N_3786);
nand U7979 (N_7979,N_3294,N_4652);
nor U7980 (N_7980,N_5916,N_3474);
or U7981 (N_7981,N_5091,N_3886);
or U7982 (N_7982,N_3312,N_6247);
and U7983 (N_7983,N_4169,N_5456);
nor U7984 (N_7984,N_3270,N_3341);
and U7985 (N_7985,N_4656,N_4790);
or U7986 (N_7986,N_4622,N_5907);
and U7987 (N_7987,N_5758,N_3391);
nand U7988 (N_7988,N_4696,N_4246);
or U7989 (N_7989,N_5770,N_6088);
xor U7990 (N_7990,N_3832,N_3547);
nor U7991 (N_7991,N_6115,N_5740);
and U7992 (N_7992,N_5430,N_5380);
or U7993 (N_7993,N_3383,N_5315);
or U7994 (N_7994,N_4345,N_4838);
xor U7995 (N_7995,N_4771,N_4554);
nor U7996 (N_7996,N_4174,N_5226);
xnor U7997 (N_7997,N_5065,N_4770);
or U7998 (N_7998,N_5983,N_5661);
and U7999 (N_7999,N_4147,N_4936);
nor U8000 (N_8000,N_3886,N_5424);
nand U8001 (N_8001,N_5984,N_3244);
nand U8002 (N_8002,N_3397,N_4752);
or U8003 (N_8003,N_4892,N_5185);
and U8004 (N_8004,N_3957,N_5264);
and U8005 (N_8005,N_5814,N_5899);
and U8006 (N_8006,N_4887,N_4204);
nor U8007 (N_8007,N_4145,N_4153);
or U8008 (N_8008,N_5870,N_4141);
nand U8009 (N_8009,N_3384,N_5804);
nor U8010 (N_8010,N_4710,N_5291);
xor U8011 (N_8011,N_3599,N_3502);
or U8012 (N_8012,N_5512,N_3489);
and U8013 (N_8013,N_4436,N_5393);
and U8014 (N_8014,N_5757,N_6167);
xnor U8015 (N_8015,N_4682,N_5557);
or U8016 (N_8016,N_4594,N_5498);
nor U8017 (N_8017,N_5122,N_4013);
or U8018 (N_8018,N_3694,N_4300);
xnor U8019 (N_8019,N_5263,N_5302);
nor U8020 (N_8020,N_6015,N_5938);
nand U8021 (N_8021,N_3886,N_5163);
xor U8022 (N_8022,N_4078,N_5562);
and U8023 (N_8023,N_5405,N_3496);
or U8024 (N_8024,N_4106,N_3282);
nand U8025 (N_8025,N_5675,N_4251);
xnor U8026 (N_8026,N_5596,N_3173);
or U8027 (N_8027,N_6130,N_5419);
nor U8028 (N_8028,N_3467,N_3235);
nand U8029 (N_8029,N_4615,N_5171);
and U8030 (N_8030,N_5247,N_3213);
and U8031 (N_8031,N_3993,N_5703);
nand U8032 (N_8032,N_3202,N_3206);
nand U8033 (N_8033,N_5170,N_6015);
xor U8034 (N_8034,N_4370,N_5872);
and U8035 (N_8035,N_5872,N_3932);
and U8036 (N_8036,N_5849,N_3772);
and U8037 (N_8037,N_4157,N_3650);
or U8038 (N_8038,N_5195,N_5333);
or U8039 (N_8039,N_4290,N_3966);
nor U8040 (N_8040,N_4333,N_3518);
nor U8041 (N_8041,N_3884,N_3550);
nor U8042 (N_8042,N_3323,N_3519);
xnor U8043 (N_8043,N_5019,N_5510);
xor U8044 (N_8044,N_4583,N_3403);
or U8045 (N_8045,N_3804,N_5669);
nand U8046 (N_8046,N_5869,N_3619);
nor U8047 (N_8047,N_5353,N_3308);
nand U8048 (N_8048,N_5926,N_6183);
nand U8049 (N_8049,N_4439,N_5576);
nand U8050 (N_8050,N_4188,N_5955);
or U8051 (N_8051,N_5857,N_4786);
nor U8052 (N_8052,N_5020,N_5189);
nor U8053 (N_8053,N_3432,N_4301);
and U8054 (N_8054,N_5276,N_4000);
or U8055 (N_8055,N_4144,N_3972);
or U8056 (N_8056,N_4136,N_4866);
and U8057 (N_8057,N_3956,N_4812);
nor U8058 (N_8058,N_6038,N_3259);
nand U8059 (N_8059,N_4467,N_3149);
and U8060 (N_8060,N_3476,N_5491);
nand U8061 (N_8061,N_4202,N_5222);
nand U8062 (N_8062,N_6079,N_6217);
and U8063 (N_8063,N_4667,N_5688);
or U8064 (N_8064,N_5380,N_5841);
xor U8065 (N_8065,N_4542,N_3321);
or U8066 (N_8066,N_3838,N_3754);
or U8067 (N_8067,N_4179,N_4042);
or U8068 (N_8068,N_3773,N_3596);
or U8069 (N_8069,N_4620,N_4045);
nand U8070 (N_8070,N_4292,N_5950);
and U8071 (N_8071,N_4210,N_5337);
nor U8072 (N_8072,N_5468,N_4644);
xor U8073 (N_8073,N_3190,N_3148);
nor U8074 (N_8074,N_3126,N_4400);
nor U8075 (N_8075,N_4560,N_3507);
or U8076 (N_8076,N_5159,N_5038);
and U8077 (N_8077,N_5389,N_5767);
nor U8078 (N_8078,N_3878,N_4548);
nand U8079 (N_8079,N_3371,N_3360);
xnor U8080 (N_8080,N_4895,N_5519);
and U8081 (N_8081,N_4707,N_3323);
and U8082 (N_8082,N_3437,N_5719);
nor U8083 (N_8083,N_4231,N_5447);
nand U8084 (N_8084,N_3964,N_4443);
or U8085 (N_8085,N_4961,N_5282);
and U8086 (N_8086,N_3698,N_5347);
nand U8087 (N_8087,N_5897,N_5005);
and U8088 (N_8088,N_3509,N_4329);
or U8089 (N_8089,N_5760,N_4758);
xnor U8090 (N_8090,N_3888,N_3463);
and U8091 (N_8091,N_3804,N_3200);
or U8092 (N_8092,N_3996,N_5921);
xnor U8093 (N_8093,N_5549,N_4561);
and U8094 (N_8094,N_6025,N_3153);
or U8095 (N_8095,N_4740,N_4078);
and U8096 (N_8096,N_5320,N_5622);
xnor U8097 (N_8097,N_3613,N_3916);
xor U8098 (N_8098,N_5970,N_4195);
nor U8099 (N_8099,N_4675,N_4022);
and U8100 (N_8100,N_5054,N_4007);
nand U8101 (N_8101,N_5856,N_3392);
and U8102 (N_8102,N_6187,N_3299);
or U8103 (N_8103,N_5490,N_4338);
nor U8104 (N_8104,N_4664,N_5669);
nor U8105 (N_8105,N_4193,N_3357);
nand U8106 (N_8106,N_4376,N_4261);
nand U8107 (N_8107,N_5922,N_5633);
and U8108 (N_8108,N_4586,N_4911);
and U8109 (N_8109,N_3279,N_4672);
and U8110 (N_8110,N_4223,N_5859);
and U8111 (N_8111,N_6010,N_3825);
nor U8112 (N_8112,N_3211,N_4816);
or U8113 (N_8113,N_5914,N_5794);
nand U8114 (N_8114,N_5926,N_3423);
nand U8115 (N_8115,N_5013,N_5491);
nand U8116 (N_8116,N_3129,N_4843);
or U8117 (N_8117,N_4311,N_4374);
nor U8118 (N_8118,N_3758,N_4157);
xor U8119 (N_8119,N_5166,N_4114);
or U8120 (N_8120,N_3767,N_5159);
nand U8121 (N_8121,N_5301,N_6067);
and U8122 (N_8122,N_3868,N_3769);
xnor U8123 (N_8123,N_5080,N_3495);
nand U8124 (N_8124,N_4047,N_4893);
nand U8125 (N_8125,N_4203,N_4318);
xor U8126 (N_8126,N_5466,N_5986);
or U8127 (N_8127,N_5925,N_4176);
and U8128 (N_8128,N_5201,N_5964);
xor U8129 (N_8129,N_4372,N_4397);
xnor U8130 (N_8130,N_3380,N_3804);
nand U8131 (N_8131,N_4445,N_4960);
nand U8132 (N_8132,N_4494,N_6034);
or U8133 (N_8133,N_5750,N_5628);
and U8134 (N_8134,N_4651,N_3801);
or U8135 (N_8135,N_6226,N_4324);
xnor U8136 (N_8136,N_4845,N_4906);
xor U8137 (N_8137,N_5226,N_3723);
nand U8138 (N_8138,N_3867,N_5990);
or U8139 (N_8139,N_3714,N_5508);
nand U8140 (N_8140,N_4776,N_3741);
or U8141 (N_8141,N_3461,N_4473);
and U8142 (N_8142,N_6205,N_4321);
or U8143 (N_8143,N_5415,N_3130);
or U8144 (N_8144,N_5640,N_5202);
nor U8145 (N_8145,N_4334,N_4994);
and U8146 (N_8146,N_4368,N_3856);
or U8147 (N_8147,N_5636,N_5621);
xnor U8148 (N_8148,N_5777,N_3770);
xnor U8149 (N_8149,N_3807,N_5991);
nor U8150 (N_8150,N_3330,N_3517);
xor U8151 (N_8151,N_4979,N_3621);
and U8152 (N_8152,N_6242,N_3673);
or U8153 (N_8153,N_4883,N_5858);
or U8154 (N_8154,N_6165,N_3405);
nor U8155 (N_8155,N_5460,N_5849);
nand U8156 (N_8156,N_4811,N_5536);
xnor U8157 (N_8157,N_5860,N_4363);
nor U8158 (N_8158,N_3169,N_3656);
nand U8159 (N_8159,N_4678,N_4984);
and U8160 (N_8160,N_3538,N_5522);
nand U8161 (N_8161,N_6203,N_4106);
and U8162 (N_8162,N_3126,N_3723);
xor U8163 (N_8163,N_3616,N_3609);
or U8164 (N_8164,N_5229,N_3596);
nand U8165 (N_8165,N_4828,N_5609);
or U8166 (N_8166,N_5382,N_3686);
nor U8167 (N_8167,N_4163,N_3215);
and U8168 (N_8168,N_4875,N_3129);
nor U8169 (N_8169,N_3312,N_6204);
nand U8170 (N_8170,N_4172,N_4058);
and U8171 (N_8171,N_4306,N_5752);
xnor U8172 (N_8172,N_3207,N_3311);
or U8173 (N_8173,N_3784,N_3942);
xor U8174 (N_8174,N_4817,N_4065);
nor U8175 (N_8175,N_3125,N_3493);
nor U8176 (N_8176,N_4467,N_6015);
xnor U8177 (N_8177,N_3504,N_4051);
and U8178 (N_8178,N_3341,N_5474);
and U8179 (N_8179,N_5715,N_5526);
nand U8180 (N_8180,N_4685,N_4892);
xnor U8181 (N_8181,N_4455,N_4984);
or U8182 (N_8182,N_3259,N_4065);
and U8183 (N_8183,N_5423,N_4915);
xnor U8184 (N_8184,N_5244,N_4370);
nor U8185 (N_8185,N_4179,N_4622);
and U8186 (N_8186,N_5577,N_5809);
and U8187 (N_8187,N_4565,N_5038);
nand U8188 (N_8188,N_3870,N_3665);
xnor U8189 (N_8189,N_3130,N_4614);
and U8190 (N_8190,N_4611,N_4261);
nand U8191 (N_8191,N_4298,N_3786);
or U8192 (N_8192,N_3901,N_4921);
xor U8193 (N_8193,N_4691,N_6060);
nor U8194 (N_8194,N_5305,N_5201);
xnor U8195 (N_8195,N_5994,N_3530);
xor U8196 (N_8196,N_4544,N_3852);
or U8197 (N_8197,N_5861,N_4481);
nand U8198 (N_8198,N_4135,N_3465);
xor U8199 (N_8199,N_4251,N_4696);
nand U8200 (N_8200,N_4685,N_5374);
xnor U8201 (N_8201,N_4752,N_3411);
and U8202 (N_8202,N_3445,N_3849);
or U8203 (N_8203,N_4076,N_5239);
nand U8204 (N_8204,N_5035,N_5827);
xnor U8205 (N_8205,N_5439,N_3920);
or U8206 (N_8206,N_3682,N_4778);
nand U8207 (N_8207,N_6134,N_4565);
nand U8208 (N_8208,N_4983,N_4808);
xnor U8209 (N_8209,N_3549,N_6134);
nand U8210 (N_8210,N_6129,N_5188);
and U8211 (N_8211,N_4685,N_5644);
xor U8212 (N_8212,N_6144,N_4313);
nand U8213 (N_8213,N_5111,N_3275);
or U8214 (N_8214,N_4750,N_3692);
and U8215 (N_8215,N_3938,N_5474);
or U8216 (N_8216,N_4293,N_3161);
or U8217 (N_8217,N_6219,N_3145);
nor U8218 (N_8218,N_3560,N_3715);
nor U8219 (N_8219,N_4833,N_5620);
nor U8220 (N_8220,N_5783,N_4528);
and U8221 (N_8221,N_3415,N_3941);
or U8222 (N_8222,N_6234,N_6141);
nor U8223 (N_8223,N_4602,N_5235);
xor U8224 (N_8224,N_3381,N_5248);
and U8225 (N_8225,N_5914,N_3638);
and U8226 (N_8226,N_3834,N_5262);
or U8227 (N_8227,N_4741,N_4626);
and U8228 (N_8228,N_5895,N_3992);
and U8229 (N_8229,N_5112,N_4264);
or U8230 (N_8230,N_6021,N_3360);
xnor U8231 (N_8231,N_4060,N_3305);
nor U8232 (N_8232,N_4854,N_5066);
and U8233 (N_8233,N_6139,N_3308);
or U8234 (N_8234,N_4345,N_5083);
nor U8235 (N_8235,N_3787,N_3305);
nand U8236 (N_8236,N_3924,N_4784);
or U8237 (N_8237,N_5972,N_3519);
xor U8238 (N_8238,N_5787,N_3744);
and U8239 (N_8239,N_6237,N_3785);
nand U8240 (N_8240,N_5512,N_3804);
or U8241 (N_8241,N_4071,N_3875);
nor U8242 (N_8242,N_3624,N_5073);
nand U8243 (N_8243,N_4121,N_3710);
nor U8244 (N_8244,N_3309,N_5031);
nor U8245 (N_8245,N_5131,N_3353);
and U8246 (N_8246,N_5642,N_4767);
nor U8247 (N_8247,N_6117,N_3620);
nand U8248 (N_8248,N_4404,N_3595);
or U8249 (N_8249,N_3450,N_4150);
or U8250 (N_8250,N_4878,N_4056);
nor U8251 (N_8251,N_5653,N_5216);
xor U8252 (N_8252,N_3802,N_5611);
xnor U8253 (N_8253,N_5922,N_5801);
nand U8254 (N_8254,N_5404,N_4550);
xor U8255 (N_8255,N_4648,N_3508);
or U8256 (N_8256,N_3908,N_4156);
or U8257 (N_8257,N_5270,N_4493);
nand U8258 (N_8258,N_3181,N_3595);
nor U8259 (N_8259,N_5140,N_3317);
or U8260 (N_8260,N_4446,N_3792);
or U8261 (N_8261,N_5999,N_5354);
nor U8262 (N_8262,N_6017,N_4109);
and U8263 (N_8263,N_4725,N_3723);
or U8264 (N_8264,N_6179,N_3253);
xor U8265 (N_8265,N_5071,N_4917);
nor U8266 (N_8266,N_3917,N_4071);
xnor U8267 (N_8267,N_5288,N_5601);
xnor U8268 (N_8268,N_3813,N_5308);
nor U8269 (N_8269,N_5781,N_3227);
or U8270 (N_8270,N_6175,N_4476);
and U8271 (N_8271,N_3280,N_5994);
xor U8272 (N_8272,N_5179,N_5465);
or U8273 (N_8273,N_3502,N_3376);
nand U8274 (N_8274,N_5022,N_4268);
and U8275 (N_8275,N_5302,N_5053);
xnor U8276 (N_8276,N_3135,N_5522);
xnor U8277 (N_8277,N_4651,N_6157);
nand U8278 (N_8278,N_4449,N_6247);
nand U8279 (N_8279,N_3455,N_6101);
nor U8280 (N_8280,N_3823,N_4204);
and U8281 (N_8281,N_5720,N_4276);
nor U8282 (N_8282,N_6124,N_3430);
xnor U8283 (N_8283,N_5032,N_5203);
nand U8284 (N_8284,N_5499,N_5688);
and U8285 (N_8285,N_4488,N_3187);
nand U8286 (N_8286,N_5408,N_3436);
xor U8287 (N_8287,N_3671,N_4211);
and U8288 (N_8288,N_5311,N_4071);
nand U8289 (N_8289,N_5045,N_3696);
xor U8290 (N_8290,N_5374,N_5092);
nand U8291 (N_8291,N_4586,N_3786);
nand U8292 (N_8292,N_4852,N_5863);
or U8293 (N_8293,N_3640,N_5142);
and U8294 (N_8294,N_5064,N_4863);
nand U8295 (N_8295,N_5298,N_4205);
xor U8296 (N_8296,N_4739,N_4222);
and U8297 (N_8297,N_5062,N_6196);
nor U8298 (N_8298,N_4605,N_5943);
xnor U8299 (N_8299,N_5520,N_5761);
nor U8300 (N_8300,N_5923,N_3514);
xnor U8301 (N_8301,N_5883,N_5531);
or U8302 (N_8302,N_3654,N_4466);
and U8303 (N_8303,N_3967,N_3620);
nand U8304 (N_8304,N_3226,N_4982);
or U8305 (N_8305,N_4161,N_4712);
nand U8306 (N_8306,N_4114,N_3171);
or U8307 (N_8307,N_4032,N_3326);
or U8308 (N_8308,N_3861,N_5665);
nor U8309 (N_8309,N_3830,N_5409);
xnor U8310 (N_8310,N_5019,N_5554);
nor U8311 (N_8311,N_3373,N_3668);
or U8312 (N_8312,N_5559,N_3589);
and U8313 (N_8313,N_5405,N_5706);
nor U8314 (N_8314,N_6006,N_4399);
and U8315 (N_8315,N_4412,N_5626);
nor U8316 (N_8316,N_3649,N_4592);
xor U8317 (N_8317,N_4749,N_4947);
xnor U8318 (N_8318,N_5923,N_4125);
or U8319 (N_8319,N_5857,N_3771);
or U8320 (N_8320,N_4116,N_3411);
or U8321 (N_8321,N_5385,N_5650);
nor U8322 (N_8322,N_6136,N_4126);
xor U8323 (N_8323,N_5865,N_3929);
xor U8324 (N_8324,N_4129,N_3876);
nor U8325 (N_8325,N_4968,N_3262);
nand U8326 (N_8326,N_4873,N_5442);
and U8327 (N_8327,N_3471,N_5793);
xor U8328 (N_8328,N_4193,N_5390);
nand U8329 (N_8329,N_4192,N_5340);
nand U8330 (N_8330,N_4960,N_5150);
xor U8331 (N_8331,N_5847,N_3324);
nor U8332 (N_8332,N_4578,N_4744);
xor U8333 (N_8333,N_3598,N_4019);
nor U8334 (N_8334,N_3960,N_4068);
and U8335 (N_8335,N_3575,N_3649);
and U8336 (N_8336,N_6230,N_5872);
or U8337 (N_8337,N_4579,N_6247);
nand U8338 (N_8338,N_6164,N_5205);
and U8339 (N_8339,N_3371,N_6113);
nor U8340 (N_8340,N_4258,N_3604);
nor U8341 (N_8341,N_3757,N_5569);
or U8342 (N_8342,N_4009,N_3918);
xor U8343 (N_8343,N_5915,N_3276);
or U8344 (N_8344,N_5147,N_3881);
or U8345 (N_8345,N_4585,N_4756);
or U8346 (N_8346,N_4567,N_3795);
and U8347 (N_8347,N_4761,N_5716);
nand U8348 (N_8348,N_6090,N_5361);
and U8349 (N_8349,N_5795,N_5344);
and U8350 (N_8350,N_6194,N_5040);
nor U8351 (N_8351,N_3184,N_5473);
and U8352 (N_8352,N_4008,N_4165);
nand U8353 (N_8353,N_4597,N_4141);
xor U8354 (N_8354,N_4497,N_4310);
nor U8355 (N_8355,N_4249,N_5898);
nand U8356 (N_8356,N_3571,N_3559);
xnor U8357 (N_8357,N_4298,N_4781);
and U8358 (N_8358,N_5740,N_5378);
xnor U8359 (N_8359,N_4470,N_4675);
nand U8360 (N_8360,N_4712,N_5929);
nor U8361 (N_8361,N_5361,N_5806);
or U8362 (N_8362,N_5185,N_5043);
nand U8363 (N_8363,N_5505,N_5355);
xnor U8364 (N_8364,N_5395,N_3723);
and U8365 (N_8365,N_4514,N_4290);
or U8366 (N_8366,N_5747,N_5685);
xor U8367 (N_8367,N_5602,N_3841);
and U8368 (N_8368,N_5798,N_4727);
nor U8369 (N_8369,N_3732,N_5304);
xor U8370 (N_8370,N_3170,N_4277);
or U8371 (N_8371,N_6047,N_5348);
nor U8372 (N_8372,N_4249,N_6063);
nor U8373 (N_8373,N_4128,N_4760);
nand U8374 (N_8374,N_5529,N_5739);
xor U8375 (N_8375,N_6181,N_4071);
nand U8376 (N_8376,N_3531,N_4448);
and U8377 (N_8377,N_3569,N_5208);
or U8378 (N_8378,N_6110,N_4605);
xnor U8379 (N_8379,N_6229,N_5132);
nor U8380 (N_8380,N_3415,N_3206);
nor U8381 (N_8381,N_5206,N_3853);
nand U8382 (N_8382,N_3441,N_4583);
and U8383 (N_8383,N_5554,N_5260);
nand U8384 (N_8384,N_5430,N_3908);
and U8385 (N_8385,N_4204,N_3201);
and U8386 (N_8386,N_4443,N_6083);
xor U8387 (N_8387,N_3535,N_3235);
xor U8388 (N_8388,N_5392,N_4099);
nand U8389 (N_8389,N_5702,N_4216);
and U8390 (N_8390,N_4991,N_3739);
nand U8391 (N_8391,N_6150,N_5678);
nor U8392 (N_8392,N_3794,N_3910);
or U8393 (N_8393,N_5434,N_5805);
and U8394 (N_8394,N_5188,N_4648);
xnor U8395 (N_8395,N_5101,N_5019);
nand U8396 (N_8396,N_5542,N_3532);
nand U8397 (N_8397,N_4010,N_4463);
or U8398 (N_8398,N_5217,N_3761);
or U8399 (N_8399,N_5784,N_5192);
xor U8400 (N_8400,N_5678,N_3834);
nand U8401 (N_8401,N_4160,N_5116);
xnor U8402 (N_8402,N_4666,N_4418);
nor U8403 (N_8403,N_5311,N_5627);
xnor U8404 (N_8404,N_6044,N_5620);
xor U8405 (N_8405,N_5007,N_5357);
xor U8406 (N_8406,N_5086,N_5060);
nand U8407 (N_8407,N_4673,N_4648);
nor U8408 (N_8408,N_5137,N_3349);
or U8409 (N_8409,N_3307,N_4454);
or U8410 (N_8410,N_4552,N_4083);
xor U8411 (N_8411,N_4607,N_3200);
or U8412 (N_8412,N_5920,N_6060);
and U8413 (N_8413,N_5039,N_4116);
nand U8414 (N_8414,N_3197,N_4304);
and U8415 (N_8415,N_3467,N_3250);
nor U8416 (N_8416,N_3150,N_3972);
xor U8417 (N_8417,N_5236,N_5839);
nor U8418 (N_8418,N_4277,N_3788);
and U8419 (N_8419,N_3519,N_3364);
or U8420 (N_8420,N_4139,N_4816);
nand U8421 (N_8421,N_5648,N_5981);
or U8422 (N_8422,N_5999,N_6188);
and U8423 (N_8423,N_3958,N_3843);
and U8424 (N_8424,N_3457,N_5576);
xor U8425 (N_8425,N_4781,N_6233);
and U8426 (N_8426,N_6003,N_3837);
xor U8427 (N_8427,N_3671,N_3865);
nor U8428 (N_8428,N_3852,N_5286);
and U8429 (N_8429,N_3848,N_5346);
or U8430 (N_8430,N_5230,N_4653);
nor U8431 (N_8431,N_3786,N_5554);
xnor U8432 (N_8432,N_3347,N_3137);
or U8433 (N_8433,N_4284,N_5287);
xor U8434 (N_8434,N_4197,N_5937);
nor U8435 (N_8435,N_5201,N_3750);
and U8436 (N_8436,N_5565,N_5027);
nor U8437 (N_8437,N_6055,N_3432);
or U8438 (N_8438,N_3427,N_3675);
or U8439 (N_8439,N_3890,N_5080);
or U8440 (N_8440,N_5864,N_3462);
and U8441 (N_8441,N_5222,N_3150);
and U8442 (N_8442,N_3412,N_4227);
nand U8443 (N_8443,N_5188,N_4227);
xor U8444 (N_8444,N_3341,N_3379);
or U8445 (N_8445,N_5182,N_3215);
or U8446 (N_8446,N_4116,N_4656);
and U8447 (N_8447,N_6018,N_5306);
or U8448 (N_8448,N_5096,N_6002);
or U8449 (N_8449,N_4085,N_5474);
and U8450 (N_8450,N_3141,N_5794);
xor U8451 (N_8451,N_4223,N_5781);
or U8452 (N_8452,N_5396,N_4811);
or U8453 (N_8453,N_4338,N_4846);
nor U8454 (N_8454,N_4303,N_4069);
nand U8455 (N_8455,N_5828,N_5193);
xnor U8456 (N_8456,N_4018,N_5338);
nand U8457 (N_8457,N_4505,N_4320);
and U8458 (N_8458,N_5605,N_4758);
or U8459 (N_8459,N_5980,N_5758);
or U8460 (N_8460,N_3428,N_4080);
or U8461 (N_8461,N_4565,N_3961);
or U8462 (N_8462,N_5332,N_3767);
xnor U8463 (N_8463,N_5329,N_5192);
nor U8464 (N_8464,N_5908,N_3173);
or U8465 (N_8465,N_5666,N_6246);
nor U8466 (N_8466,N_4466,N_5644);
xnor U8467 (N_8467,N_5670,N_5517);
xor U8468 (N_8468,N_3336,N_4917);
or U8469 (N_8469,N_3242,N_4153);
nand U8470 (N_8470,N_5699,N_4807);
and U8471 (N_8471,N_4437,N_5839);
nand U8472 (N_8472,N_6024,N_3523);
xor U8473 (N_8473,N_4580,N_3585);
nand U8474 (N_8474,N_3234,N_3610);
xor U8475 (N_8475,N_5851,N_4927);
and U8476 (N_8476,N_4526,N_3986);
xnor U8477 (N_8477,N_5080,N_5229);
nand U8478 (N_8478,N_4983,N_4918);
xnor U8479 (N_8479,N_5133,N_3740);
and U8480 (N_8480,N_3812,N_5658);
or U8481 (N_8481,N_5710,N_3464);
nand U8482 (N_8482,N_4235,N_5805);
xor U8483 (N_8483,N_4667,N_5223);
and U8484 (N_8484,N_4108,N_4002);
xnor U8485 (N_8485,N_3209,N_4310);
nand U8486 (N_8486,N_4157,N_3250);
or U8487 (N_8487,N_3623,N_5796);
and U8488 (N_8488,N_5175,N_5808);
xnor U8489 (N_8489,N_4061,N_4612);
nor U8490 (N_8490,N_3206,N_3275);
or U8491 (N_8491,N_4942,N_3939);
xnor U8492 (N_8492,N_5473,N_5039);
and U8493 (N_8493,N_4798,N_4450);
xor U8494 (N_8494,N_3548,N_6193);
and U8495 (N_8495,N_5803,N_3337);
and U8496 (N_8496,N_3384,N_5801);
and U8497 (N_8497,N_5236,N_3145);
nor U8498 (N_8498,N_3304,N_3601);
and U8499 (N_8499,N_5581,N_4052);
xor U8500 (N_8500,N_4567,N_3241);
xnor U8501 (N_8501,N_4799,N_5485);
or U8502 (N_8502,N_5947,N_5219);
nor U8503 (N_8503,N_5887,N_4043);
xor U8504 (N_8504,N_6228,N_3902);
and U8505 (N_8505,N_4841,N_6114);
xnor U8506 (N_8506,N_3271,N_5958);
nor U8507 (N_8507,N_5070,N_6245);
or U8508 (N_8508,N_3475,N_3183);
nor U8509 (N_8509,N_3803,N_5334);
or U8510 (N_8510,N_5320,N_5846);
and U8511 (N_8511,N_4113,N_5923);
nand U8512 (N_8512,N_4046,N_5932);
xnor U8513 (N_8513,N_4203,N_4538);
or U8514 (N_8514,N_5383,N_4642);
nand U8515 (N_8515,N_4380,N_6221);
or U8516 (N_8516,N_5823,N_4606);
nand U8517 (N_8517,N_3564,N_3601);
nor U8518 (N_8518,N_5347,N_3876);
and U8519 (N_8519,N_4757,N_5512);
nor U8520 (N_8520,N_4556,N_4847);
nand U8521 (N_8521,N_4045,N_3735);
and U8522 (N_8522,N_4949,N_5298);
nor U8523 (N_8523,N_4805,N_3825);
and U8524 (N_8524,N_3176,N_4504);
xor U8525 (N_8525,N_3378,N_3613);
nand U8526 (N_8526,N_5999,N_4902);
nand U8527 (N_8527,N_4069,N_6035);
nor U8528 (N_8528,N_6155,N_3705);
nand U8529 (N_8529,N_3230,N_5725);
and U8530 (N_8530,N_5759,N_4242);
xnor U8531 (N_8531,N_4134,N_5290);
nand U8532 (N_8532,N_4252,N_4801);
and U8533 (N_8533,N_6215,N_5253);
nor U8534 (N_8534,N_3221,N_6043);
and U8535 (N_8535,N_4646,N_5509);
nand U8536 (N_8536,N_3893,N_4568);
nor U8537 (N_8537,N_4720,N_6192);
xor U8538 (N_8538,N_5528,N_5191);
nand U8539 (N_8539,N_4220,N_3784);
and U8540 (N_8540,N_5464,N_3339);
or U8541 (N_8541,N_3376,N_4360);
nand U8542 (N_8542,N_3537,N_5006);
nor U8543 (N_8543,N_5128,N_3669);
nor U8544 (N_8544,N_3929,N_6034);
or U8545 (N_8545,N_6213,N_3839);
nor U8546 (N_8546,N_4233,N_4890);
nor U8547 (N_8547,N_3802,N_5901);
nor U8548 (N_8548,N_4120,N_3187);
or U8549 (N_8549,N_4240,N_5657);
xnor U8550 (N_8550,N_3162,N_6038);
nand U8551 (N_8551,N_4572,N_3162);
nand U8552 (N_8552,N_4038,N_5285);
nand U8553 (N_8553,N_5246,N_4395);
nand U8554 (N_8554,N_5301,N_5057);
nand U8555 (N_8555,N_3790,N_5376);
and U8556 (N_8556,N_4994,N_5327);
xnor U8557 (N_8557,N_3903,N_3501);
nand U8558 (N_8558,N_5761,N_3708);
or U8559 (N_8559,N_3181,N_4253);
nand U8560 (N_8560,N_3535,N_4481);
xnor U8561 (N_8561,N_4448,N_3527);
xor U8562 (N_8562,N_5952,N_5019);
xnor U8563 (N_8563,N_4246,N_5698);
and U8564 (N_8564,N_3614,N_4840);
nor U8565 (N_8565,N_3569,N_4111);
and U8566 (N_8566,N_3654,N_3775);
xnor U8567 (N_8567,N_5361,N_4222);
or U8568 (N_8568,N_4556,N_4799);
xnor U8569 (N_8569,N_5525,N_3429);
or U8570 (N_8570,N_5112,N_5116);
or U8571 (N_8571,N_4781,N_5941);
nand U8572 (N_8572,N_3416,N_5549);
xnor U8573 (N_8573,N_5413,N_3275);
or U8574 (N_8574,N_5177,N_3357);
xnor U8575 (N_8575,N_3490,N_3305);
or U8576 (N_8576,N_5774,N_5631);
nor U8577 (N_8577,N_3165,N_4036);
or U8578 (N_8578,N_5755,N_3679);
nand U8579 (N_8579,N_4149,N_5982);
or U8580 (N_8580,N_5982,N_3240);
xor U8581 (N_8581,N_4467,N_5056);
nor U8582 (N_8582,N_4620,N_3880);
xor U8583 (N_8583,N_3378,N_4613);
nand U8584 (N_8584,N_5459,N_3226);
and U8585 (N_8585,N_5828,N_5699);
nand U8586 (N_8586,N_3579,N_4873);
and U8587 (N_8587,N_4947,N_3754);
nand U8588 (N_8588,N_4561,N_5416);
and U8589 (N_8589,N_3257,N_4815);
nand U8590 (N_8590,N_3479,N_3202);
xor U8591 (N_8591,N_3453,N_3835);
xor U8592 (N_8592,N_3411,N_4088);
and U8593 (N_8593,N_3470,N_5537);
nor U8594 (N_8594,N_3883,N_4048);
xnor U8595 (N_8595,N_5986,N_5395);
nand U8596 (N_8596,N_5775,N_5061);
nand U8597 (N_8597,N_6168,N_4945);
and U8598 (N_8598,N_4096,N_3746);
nand U8599 (N_8599,N_5285,N_4478);
and U8600 (N_8600,N_3213,N_6211);
nor U8601 (N_8601,N_4617,N_3726);
or U8602 (N_8602,N_3813,N_4659);
xnor U8603 (N_8603,N_5099,N_6037);
nand U8604 (N_8604,N_5686,N_5309);
nand U8605 (N_8605,N_4788,N_5322);
xnor U8606 (N_8606,N_4087,N_3703);
or U8607 (N_8607,N_4195,N_5580);
nor U8608 (N_8608,N_6148,N_5456);
and U8609 (N_8609,N_3649,N_5637);
xnor U8610 (N_8610,N_5945,N_3979);
nand U8611 (N_8611,N_5665,N_4302);
nor U8612 (N_8612,N_4215,N_6161);
xor U8613 (N_8613,N_5422,N_5989);
or U8614 (N_8614,N_6215,N_3579);
nor U8615 (N_8615,N_6018,N_4278);
xnor U8616 (N_8616,N_5542,N_6219);
nor U8617 (N_8617,N_3836,N_3892);
xor U8618 (N_8618,N_5496,N_6015);
xor U8619 (N_8619,N_3748,N_4183);
xnor U8620 (N_8620,N_6152,N_5703);
or U8621 (N_8621,N_5423,N_5155);
xnor U8622 (N_8622,N_5372,N_4160);
nor U8623 (N_8623,N_5579,N_4510);
xor U8624 (N_8624,N_5622,N_3588);
xor U8625 (N_8625,N_3487,N_4748);
nand U8626 (N_8626,N_3824,N_5347);
nand U8627 (N_8627,N_3402,N_6152);
or U8628 (N_8628,N_3375,N_5572);
xnor U8629 (N_8629,N_5644,N_5538);
nand U8630 (N_8630,N_6047,N_4435);
nor U8631 (N_8631,N_3467,N_3549);
xnor U8632 (N_8632,N_5382,N_3653);
nand U8633 (N_8633,N_5585,N_4334);
or U8634 (N_8634,N_5380,N_4098);
nand U8635 (N_8635,N_3198,N_5960);
and U8636 (N_8636,N_4681,N_5882);
xnor U8637 (N_8637,N_4198,N_5009);
xor U8638 (N_8638,N_5928,N_4126);
and U8639 (N_8639,N_6117,N_4203);
nor U8640 (N_8640,N_4249,N_5553);
or U8641 (N_8641,N_5903,N_4531);
xnor U8642 (N_8642,N_5022,N_4096);
or U8643 (N_8643,N_5675,N_3242);
or U8644 (N_8644,N_5880,N_3223);
and U8645 (N_8645,N_4279,N_5565);
nand U8646 (N_8646,N_5049,N_3500);
nand U8647 (N_8647,N_5566,N_3556);
nor U8648 (N_8648,N_4500,N_3346);
nand U8649 (N_8649,N_3909,N_3605);
nand U8650 (N_8650,N_4990,N_5189);
nor U8651 (N_8651,N_3392,N_3244);
xor U8652 (N_8652,N_4280,N_5632);
or U8653 (N_8653,N_6053,N_4751);
nor U8654 (N_8654,N_5813,N_4871);
and U8655 (N_8655,N_4634,N_6045);
xor U8656 (N_8656,N_5792,N_3212);
or U8657 (N_8657,N_3849,N_4842);
nand U8658 (N_8658,N_5667,N_4518);
or U8659 (N_8659,N_3447,N_4783);
and U8660 (N_8660,N_6093,N_4304);
xor U8661 (N_8661,N_4858,N_4976);
and U8662 (N_8662,N_5400,N_3511);
nand U8663 (N_8663,N_5859,N_5076);
nand U8664 (N_8664,N_3966,N_4606);
nor U8665 (N_8665,N_4152,N_4346);
and U8666 (N_8666,N_5464,N_4511);
and U8667 (N_8667,N_3168,N_5218);
xor U8668 (N_8668,N_4898,N_3451);
and U8669 (N_8669,N_4513,N_3333);
or U8670 (N_8670,N_3551,N_3436);
xor U8671 (N_8671,N_4605,N_4012);
nand U8672 (N_8672,N_4106,N_4897);
nand U8673 (N_8673,N_5133,N_3542);
nand U8674 (N_8674,N_4981,N_5446);
or U8675 (N_8675,N_4753,N_3655);
and U8676 (N_8676,N_5475,N_5180);
nand U8677 (N_8677,N_5510,N_5528);
or U8678 (N_8678,N_4287,N_3496);
and U8679 (N_8679,N_6227,N_5524);
and U8680 (N_8680,N_4672,N_6003);
xor U8681 (N_8681,N_5091,N_5411);
and U8682 (N_8682,N_4966,N_4665);
or U8683 (N_8683,N_4376,N_4439);
and U8684 (N_8684,N_3437,N_3610);
nor U8685 (N_8685,N_4054,N_5059);
xor U8686 (N_8686,N_3416,N_4591);
and U8687 (N_8687,N_5449,N_5388);
or U8688 (N_8688,N_3278,N_5152);
or U8689 (N_8689,N_5023,N_5594);
nor U8690 (N_8690,N_4290,N_3196);
nor U8691 (N_8691,N_5456,N_5233);
nand U8692 (N_8692,N_4697,N_4190);
xnor U8693 (N_8693,N_4557,N_4790);
nand U8694 (N_8694,N_5137,N_5761);
and U8695 (N_8695,N_6061,N_5176);
or U8696 (N_8696,N_5082,N_6061);
xor U8697 (N_8697,N_4500,N_5641);
xnor U8698 (N_8698,N_4750,N_5877);
or U8699 (N_8699,N_5350,N_5785);
nand U8700 (N_8700,N_3840,N_3935);
or U8701 (N_8701,N_5713,N_5711);
nor U8702 (N_8702,N_4567,N_4721);
nor U8703 (N_8703,N_5706,N_3263);
xnor U8704 (N_8704,N_4615,N_4211);
or U8705 (N_8705,N_4565,N_6093);
or U8706 (N_8706,N_6225,N_3212);
or U8707 (N_8707,N_5587,N_6149);
nand U8708 (N_8708,N_5607,N_3895);
nand U8709 (N_8709,N_6153,N_6035);
or U8710 (N_8710,N_5607,N_5230);
and U8711 (N_8711,N_3240,N_3203);
nand U8712 (N_8712,N_4723,N_6034);
or U8713 (N_8713,N_4579,N_3268);
nor U8714 (N_8714,N_5315,N_5035);
nand U8715 (N_8715,N_5165,N_5019);
nand U8716 (N_8716,N_4100,N_5834);
nor U8717 (N_8717,N_4296,N_3502);
and U8718 (N_8718,N_4399,N_5686);
xnor U8719 (N_8719,N_3634,N_4870);
or U8720 (N_8720,N_4547,N_3812);
xor U8721 (N_8721,N_6067,N_4070);
nand U8722 (N_8722,N_3448,N_3173);
and U8723 (N_8723,N_5086,N_5421);
and U8724 (N_8724,N_5629,N_5071);
and U8725 (N_8725,N_5130,N_3849);
nand U8726 (N_8726,N_3270,N_3671);
nor U8727 (N_8727,N_4201,N_4918);
or U8728 (N_8728,N_4046,N_6186);
or U8729 (N_8729,N_3685,N_3232);
and U8730 (N_8730,N_3230,N_4722);
or U8731 (N_8731,N_3733,N_6006);
nand U8732 (N_8732,N_4170,N_3207);
xnor U8733 (N_8733,N_4149,N_4419);
nor U8734 (N_8734,N_4766,N_5405);
xor U8735 (N_8735,N_5649,N_5303);
nor U8736 (N_8736,N_5137,N_5829);
xor U8737 (N_8737,N_3740,N_3941);
nor U8738 (N_8738,N_5547,N_5244);
or U8739 (N_8739,N_5195,N_4453);
or U8740 (N_8740,N_4110,N_3669);
or U8741 (N_8741,N_4432,N_5000);
nand U8742 (N_8742,N_5227,N_4073);
xor U8743 (N_8743,N_4922,N_5124);
nand U8744 (N_8744,N_3413,N_4641);
or U8745 (N_8745,N_3820,N_4715);
nor U8746 (N_8746,N_4990,N_3253);
or U8747 (N_8747,N_3476,N_3680);
nand U8748 (N_8748,N_4975,N_4317);
and U8749 (N_8749,N_4526,N_4788);
xnor U8750 (N_8750,N_5689,N_5761);
nor U8751 (N_8751,N_4481,N_3943);
and U8752 (N_8752,N_3988,N_3411);
xnor U8753 (N_8753,N_3987,N_5469);
xor U8754 (N_8754,N_5434,N_3602);
and U8755 (N_8755,N_5739,N_3666);
xnor U8756 (N_8756,N_5528,N_4551);
nand U8757 (N_8757,N_3181,N_6005);
or U8758 (N_8758,N_5131,N_3191);
nor U8759 (N_8759,N_5632,N_5395);
xnor U8760 (N_8760,N_4462,N_5990);
or U8761 (N_8761,N_5381,N_4930);
or U8762 (N_8762,N_4676,N_3796);
nor U8763 (N_8763,N_4849,N_6072);
or U8764 (N_8764,N_5313,N_5044);
nor U8765 (N_8765,N_5211,N_3437);
or U8766 (N_8766,N_4260,N_5830);
or U8767 (N_8767,N_4100,N_5809);
nor U8768 (N_8768,N_3792,N_4836);
and U8769 (N_8769,N_5240,N_4762);
or U8770 (N_8770,N_3484,N_5857);
xnor U8771 (N_8771,N_4035,N_4284);
or U8772 (N_8772,N_4127,N_4396);
and U8773 (N_8773,N_4720,N_4277);
nand U8774 (N_8774,N_5052,N_3743);
nor U8775 (N_8775,N_5723,N_5987);
or U8776 (N_8776,N_4680,N_5985);
nand U8777 (N_8777,N_3803,N_5074);
and U8778 (N_8778,N_5586,N_3454);
and U8779 (N_8779,N_3755,N_4766);
or U8780 (N_8780,N_5347,N_4227);
xnor U8781 (N_8781,N_5594,N_3939);
and U8782 (N_8782,N_6078,N_5967);
nand U8783 (N_8783,N_5594,N_5582);
nand U8784 (N_8784,N_5560,N_5984);
or U8785 (N_8785,N_3417,N_4900);
nand U8786 (N_8786,N_3981,N_4209);
xor U8787 (N_8787,N_4197,N_5780);
and U8788 (N_8788,N_6239,N_3724);
xnor U8789 (N_8789,N_3774,N_6018);
or U8790 (N_8790,N_5302,N_5422);
xor U8791 (N_8791,N_4247,N_5852);
nor U8792 (N_8792,N_4653,N_6136);
and U8793 (N_8793,N_5707,N_6009);
and U8794 (N_8794,N_3376,N_5407);
nor U8795 (N_8795,N_5859,N_6024);
nand U8796 (N_8796,N_6159,N_4388);
xnor U8797 (N_8797,N_3269,N_4321);
or U8798 (N_8798,N_3908,N_4263);
or U8799 (N_8799,N_5476,N_4494);
xor U8800 (N_8800,N_3242,N_5085);
nor U8801 (N_8801,N_4967,N_3680);
or U8802 (N_8802,N_6023,N_5390);
or U8803 (N_8803,N_3731,N_3589);
xor U8804 (N_8804,N_4339,N_5561);
or U8805 (N_8805,N_5800,N_5946);
xnor U8806 (N_8806,N_5489,N_5956);
xor U8807 (N_8807,N_4333,N_3760);
xnor U8808 (N_8808,N_5170,N_4435);
nor U8809 (N_8809,N_3609,N_6024);
or U8810 (N_8810,N_3129,N_5196);
and U8811 (N_8811,N_5939,N_5336);
nor U8812 (N_8812,N_3947,N_4138);
and U8813 (N_8813,N_5163,N_5506);
or U8814 (N_8814,N_4145,N_3465);
nor U8815 (N_8815,N_5647,N_5401);
nand U8816 (N_8816,N_4069,N_5577);
nor U8817 (N_8817,N_5746,N_4395);
nor U8818 (N_8818,N_4654,N_3931);
and U8819 (N_8819,N_4140,N_6096);
and U8820 (N_8820,N_3159,N_4529);
nand U8821 (N_8821,N_4526,N_3613);
nor U8822 (N_8822,N_6171,N_6193);
xor U8823 (N_8823,N_3882,N_5763);
nand U8824 (N_8824,N_6142,N_5375);
xor U8825 (N_8825,N_3311,N_4395);
and U8826 (N_8826,N_4873,N_4449);
and U8827 (N_8827,N_3519,N_4820);
nor U8828 (N_8828,N_3309,N_5941);
nor U8829 (N_8829,N_3334,N_5096);
xor U8830 (N_8830,N_5980,N_5988);
xor U8831 (N_8831,N_3481,N_5732);
nor U8832 (N_8832,N_3206,N_3773);
nand U8833 (N_8833,N_6171,N_6216);
nor U8834 (N_8834,N_4170,N_3151);
nor U8835 (N_8835,N_6197,N_3851);
nand U8836 (N_8836,N_5889,N_3667);
or U8837 (N_8837,N_5742,N_6049);
xor U8838 (N_8838,N_3846,N_3295);
or U8839 (N_8839,N_4302,N_6210);
or U8840 (N_8840,N_5473,N_5208);
and U8841 (N_8841,N_5620,N_4149);
and U8842 (N_8842,N_3624,N_6213);
nor U8843 (N_8843,N_4767,N_5929);
nor U8844 (N_8844,N_3167,N_6077);
nor U8845 (N_8845,N_4970,N_4634);
xnor U8846 (N_8846,N_6241,N_4796);
xor U8847 (N_8847,N_3541,N_3443);
nand U8848 (N_8848,N_5672,N_5317);
nor U8849 (N_8849,N_6033,N_5847);
or U8850 (N_8850,N_6163,N_4818);
and U8851 (N_8851,N_5037,N_6014);
or U8852 (N_8852,N_6185,N_5096);
nand U8853 (N_8853,N_5593,N_3227);
nand U8854 (N_8854,N_4351,N_4663);
and U8855 (N_8855,N_5851,N_4144);
nand U8856 (N_8856,N_4347,N_3357);
xnor U8857 (N_8857,N_3151,N_5163);
xor U8858 (N_8858,N_5896,N_3184);
and U8859 (N_8859,N_5019,N_4987);
nand U8860 (N_8860,N_4859,N_3828);
and U8861 (N_8861,N_4474,N_5750);
nand U8862 (N_8862,N_4306,N_6161);
and U8863 (N_8863,N_3991,N_5595);
nor U8864 (N_8864,N_4412,N_5335);
or U8865 (N_8865,N_4280,N_4334);
or U8866 (N_8866,N_5900,N_3411);
or U8867 (N_8867,N_4172,N_3699);
and U8868 (N_8868,N_4405,N_4522);
nand U8869 (N_8869,N_4491,N_4925);
nor U8870 (N_8870,N_5905,N_5738);
and U8871 (N_8871,N_4777,N_6132);
and U8872 (N_8872,N_4606,N_5425);
or U8873 (N_8873,N_5131,N_3948);
nand U8874 (N_8874,N_5855,N_3444);
and U8875 (N_8875,N_3626,N_5907);
nand U8876 (N_8876,N_5787,N_5521);
xnor U8877 (N_8877,N_3422,N_4464);
xor U8878 (N_8878,N_4702,N_5590);
xor U8879 (N_8879,N_5174,N_5704);
xor U8880 (N_8880,N_4200,N_6026);
nand U8881 (N_8881,N_5858,N_5098);
and U8882 (N_8882,N_5535,N_3265);
xnor U8883 (N_8883,N_4354,N_4988);
nor U8884 (N_8884,N_3723,N_3405);
and U8885 (N_8885,N_5820,N_3490);
or U8886 (N_8886,N_3591,N_5787);
nor U8887 (N_8887,N_6229,N_4459);
and U8888 (N_8888,N_3785,N_4019);
and U8889 (N_8889,N_3467,N_4686);
xnor U8890 (N_8890,N_4253,N_6234);
xor U8891 (N_8891,N_4750,N_5026);
nor U8892 (N_8892,N_4481,N_4341);
or U8893 (N_8893,N_3686,N_5823);
xor U8894 (N_8894,N_4300,N_5627);
and U8895 (N_8895,N_5973,N_4627);
or U8896 (N_8896,N_5786,N_3215);
xnor U8897 (N_8897,N_3411,N_3211);
xor U8898 (N_8898,N_6187,N_4271);
nand U8899 (N_8899,N_4459,N_4608);
xnor U8900 (N_8900,N_5264,N_5051);
or U8901 (N_8901,N_5117,N_5393);
nand U8902 (N_8902,N_3428,N_4917);
nand U8903 (N_8903,N_6174,N_3678);
nand U8904 (N_8904,N_3243,N_6160);
nand U8905 (N_8905,N_4692,N_5145);
xor U8906 (N_8906,N_4312,N_4139);
xnor U8907 (N_8907,N_6057,N_5677);
xor U8908 (N_8908,N_4995,N_5344);
nor U8909 (N_8909,N_5966,N_4167);
nand U8910 (N_8910,N_5192,N_4483);
and U8911 (N_8911,N_4697,N_3750);
or U8912 (N_8912,N_3679,N_6029);
or U8913 (N_8913,N_3676,N_5373);
nor U8914 (N_8914,N_3978,N_5362);
xnor U8915 (N_8915,N_5535,N_4368);
and U8916 (N_8916,N_4178,N_5119);
or U8917 (N_8917,N_5807,N_4791);
and U8918 (N_8918,N_3527,N_4231);
xor U8919 (N_8919,N_5474,N_4788);
or U8920 (N_8920,N_3246,N_4152);
nor U8921 (N_8921,N_6048,N_3698);
xnor U8922 (N_8922,N_3904,N_3758);
nand U8923 (N_8923,N_4437,N_3272);
or U8924 (N_8924,N_4305,N_5325);
nor U8925 (N_8925,N_6080,N_3696);
xor U8926 (N_8926,N_5796,N_5860);
nor U8927 (N_8927,N_3210,N_6102);
nor U8928 (N_8928,N_5648,N_4121);
nor U8929 (N_8929,N_4488,N_3421);
nor U8930 (N_8930,N_4088,N_3408);
nand U8931 (N_8931,N_4161,N_4467);
nor U8932 (N_8932,N_3785,N_5086);
or U8933 (N_8933,N_6061,N_6178);
xor U8934 (N_8934,N_3447,N_3810);
nor U8935 (N_8935,N_4940,N_4946);
nor U8936 (N_8936,N_4452,N_6190);
xnor U8937 (N_8937,N_5037,N_4043);
xnor U8938 (N_8938,N_5915,N_5518);
or U8939 (N_8939,N_3129,N_3498);
nand U8940 (N_8940,N_3621,N_5611);
xor U8941 (N_8941,N_3424,N_5640);
and U8942 (N_8942,N_5362,N_4166);
or U8943 (N_8943,N_5142,N_4755);
nor U8944 (N_8944,N_6179,N_4446);
xor U8945 (N_8945,N_3985,N_4571);
and U8946 (N_8946,N_4513,N_4755);
nor U8947 (N_8947,N_3248,N_4151);
xnor U8948 (N_8948,N_4925,N_3905);
xor U8949 (N_8949,N_4268,N_4310);
and U8950 (N_8950,N_3931,N_5892);
and U8951 (N_8951,N_5320,N_3168);
nand U8952 (N_8952,N_4484,N_4090);
or U8953 (N_8953,N_4094,N_5299);
xor U8954 (N_8954,N_3585,N_5681);
nor U8955 (N_8955,N_4014,N_4789);
and U8956 (N_8956,N_4474,N_4921);
xor U8957 (N_8957,N_3832,N_3700);
or U8958 (N_8958,N_3536,N_3214);
nor U8959 (N_8959,N_6136,N_4674);
xor U8960 (N_8960,N_5337,N_4563);
xor U8961 (N_8961,N_5390,N_4330);
nand U8962 (N_8962,N_3624,N_5017);
and U8963 (N_8963,N_6045,N_4157);
nor U8964 (N_8964,N_4325,N_5889);
nand U8965 (N_8965,N_4211,N_5854);
nor U8966 (N_8966,N_4665,N_3999);
nand U8967 (N_8967,N_5033,N_4333);
and U8968 (N_8968,N_4928,N_3239);
nand U8969 (N_8969,N_4727,N_5835);
xnor U8970 (N_8970,N_3742,N_4373);
nor U8971 (N_8971,N_6183,N_5226);
or U8972 (N_8972,N_4681,N_4363);
and U8973 (N_8973,N_4786,N_3216);
xnor U8974 (N_8974,N_4214,N_5796);
and U8975 (N_8975,N_3660,N_3517);
and U8976 (N_8976,N_6115,N_5558);
nand U8977 (N_8977,N_5788,N_5387);
or U8978 (N_8978,N_3346,N_5130);
or U8979 (N_8979,N_3228,N_4864);
nand U8980 (N_8980,N_6061,N_3944);
and U8981 (N_8981,N_3641,N_4939);
nand U8982 (N_8982,N_6070,N_5538);
xnor U8983 (N_8983,N_3142,N_4883);
or U8984 (N_8984,N_6106,N_6184);
and U8985 (N_8985,N_4347,N_6168);
nor U8986 (N_8986,N_3344,N_3381);
and U8987 (N_8987,N_5651,N_4696);
nor U8988 (N_8988,N_3324,N_4461);
or U8989 (N_8989,N_3847,N_3591);
xnor U8990 (N_8990,N_5861,N_3316);
and U8991 (N_8991,N_5673,N_5420);
xor U8992 (N_8992,N_5429,N_3521);
or U8993 (N_8993,N_3411,N_4897);
or U8994 (N_8994,N_5104,N_5039);
xor U8995 (N_8995,N_3716,N_3309);
nand U8996 (N_8996,N_4564,N_3718);
and U8997 (N_8997,N_4118,N_6117);
nor U8998 (N_8998,N_6038,N_3147);
or U8999 (N_8999,N_3208,N_5776);
xor U9000 (N_9000,N_3732,N_3554);
or U9001 (N_9001,N_3941,N_3917);
or U9002 (N_9002,N_3458,N_4320);
nor U9003 (N_9003,N_4500,N_5981);
and U9004 (N_9004,N_3898,N_5626);
and U9005 (N_9005,N_4067,N_4812);
and U9006 (N_9006,N_3863,N_3841);
nor U9007 (N_9007,N_4124,N_6235);
nor U9008 (N_9008,N_3147,N_5711);
nand U9009 (N_9009,N_3390,N_4549);
or U9010 (N_9010,N_4117,N_4945);
and U9011 (N_9011,N_3683,N_3617);
nand U9012 (N_9012,N_4526,N_5294);
xor U9013 (N_9013,N_4749,N_4449);
nor U9014 (N_9014,N_3506,N_4555);
nand U9015 (N_9015,N_3706,N_5422);
nor U9016 (N_9016,N_3727,N_4996);
or U9017 (N_9017,N_4482,N_3821);
or U9018 (N_9018,N_5733,N_5263);
and U9019 (N_9019,N_3655,N_5714);
or U9020 (N_9020,N_5565,N_5537);
nand U9021 (N_9021,N_4971,N_3410);
or U9022 (N_9022,N_5125,N_3342);
xnor U9023 (N_9023,N_3178,N_4642);
or U9024 (N_9024,N_4635,N_3612);
nor U9025 (N_9025,N_5361,N_4804);
or U9026 (N_9026,N_4802,N_5705);
and U9027 (N_9027,N_4713,N_3152);
nor U9028 (N_9028,N_4952,N_3167);
or U9029 (N_9029,N_6093,N_5608);
xor U9030 (N_9030,N_3632,N_5163);
and U9031 (N_9031,N_5712,N_4572);
nand U9032 (N_9032,N_3823,N_3860);
and U9033 (N_9033,N_4635,N_3438);
nor U9034 (N_9034,N_3773,N_5098);
and U9035 (N_9035,N_6080,N_4879);
or U9036 (N_9036,N_4575,N_5476);
xnor U9037 (N_9037,N_4969,N_4854);
or U9038 (N_9038,N_6209,N_3331);
and U9039 (N_9039,N_3872,N_6129);
nor U9040 (N_9040,N_5283,N_5212);
nand U9041 (N_9041,N_4929,N_3853);
nand U9042 (N_9042,N_4497,N_4298);
or U9043 (N_9043,N_3710,N_4117);
nand U9044 (N_9044,N_5116,N_4436);
or U9045 (N_9045,N_3308,N_5040);
nor U9046 (N_9046,N_5023,N_5937);
xnor U9047 (N_9047,N_5726,N_3189);
nand U9048 (N_9048,N_4550,N_4199);
xnor U9049 (N_9049,N_4953,N_4639);
nor U9050 (N_9050,N_4371,N_3508);
or U9051 (N_9051,N_5697,N_4542);
nand U9052 (N_9052,N_5584,N_5107);
nand U9053 (N_9053,N_4555,N_5584);
xnor U9054 (N_9054,N_4093,N_4977);
xor U9055 (N_9055,N_6015,N_4382);
nor U9056 (N_9056,N_4851,N_4382);
nand U9057 (N_9057,N_6225,N_4568);
nand U9058 (N_9058,N_3823,N_3740);
or U9059 (N_9059,N_3404,N_5139);
or U9060 (N_9060,N_4296,N_3244);
and U9061 (N_9061,N_5532,N_4896);
nand U9062 (N_9062,N_6155,N_5104);
xor U9063 (N_9063,N_4129,N_3212);
or U9064 (N_9064,N_5072,N_3945);
nand U9065 (N_9065,N_5199,N_5331);
nand U9066 (N_9066,N_3791,N_4920);
or U9067 (N_9067,N_5161,N_3688);
nand U9068 (N_9068,N_5744,N_5594);
or U9069 (N_9069,N_5383,N_3920);
nand U9070 (N_9070,N_5822,N_3809);
and U9071 (N_9071,N_3183,N_4103);
nor U9072 (N_9072,N_5101,N_5163);
xnor U9073 (N_9073,N_5778,N_5616);
nor U9074 (N_9074,N_4732,N_3538);
and U9075 (N_9075,N_3413,N_3543);
or U9076 (N_9076,N_5864,N_4619);
and U9077 (N_9077,N_3541,N_5455);
xnor U9078 (N_9078,N_4018,N_4175);
nand U9079 (N_9079,N_5160,N_4163);
nor U9080 (N_9080,N_4870,N_4908);
and U9081 (N_9081,N_5665,N_4864);
or U9082 (N_9082,N_4511,N_4649);
nand U9083 (N_9083,N_4680,N_3427);
nor U9084 (N_9084,N_3429,N_4730);
and U9085 (N_9085,N_4042,N_5161);
xnor U9086 (N_9086,N_5050,N_4807);
nand U9087 (N_9087,N_4643,N_4588);
or U9088 (N_9088,N_5451,N_5618);
xor U9089 (N_9089,N_5360,N_4959);
or U9090 (N_9090,N_6041,N_4443);
nor U9091 (N_9091,N_3251,N_6064);
and U9092 (N_9092,N_3699,N_3631);
and U9093 (N_9093,N_5440,N_4702);
nor U9094 (N_9094,N_3404,N_3971);
nand U9095 (N_9095,N_5379,N_5836);
xnor U9096 (N_9096,N_3565,N_3861);
or U9097 (N_9097,N_3506,N_4348);
xor U9098 (N_9098,N_6137,N_4402);
xnor U9099 (N_9099,N_5075,N_3441);
or U9100 (N_9100,N_5338,N_5282);
nand U9101 (N_9101,N_4867,N_4145);
xor U9102 (N_9102,N_4449,N_3350);
or U9103 (N_9103,N_3515,N_5117);
and U9104 (N_9104,N_4888,N_3741);
xnor U9105 (N_9105,N_4690,N_5783);
and U9106 (N_9106,N_5413,N_5785);
and U9107 (N_9107,N_5205,N_6146);
and U9108 (N_9108,N_4654,N_5423);
and U9109 (N_9109,N_6003,N_4623);
or U9110 (N_9110,N_3996,N_6015);
nor U9111 (N_9111,N_4798,N_6048);
xor U9112 (N_9112,N_5399,N_5767);
or U9113 (N_9113,N_5826,N_3809);
and U9114 (N_9114,N_5534,N_4333);
or U9115 (N_9115,N_4784,N_5760);
or U9116 (N_9116,N_3627,N_4264);
nor U9117 (N_9117,N_4020,N_5409);
or U9118 (N_9118,N_5622,N_3980);
nand U9119 (N_9119,N_5113,N_5325);
or U9120 (N_9120,N_5680,N_5467);
nor U9121 (N_9121,N_4916,N_3347);
xnor U9122 (N_9122,N_4562,N_6157);
nand U9123 (N_9123,N_3888,N_5997);
or U9124 (N_9124,N_4762,N_3319);
or U9125 (N_9125,N_3770,N_5488);
xnor U9126 (N_9126,N_4429,N_3453);
or U9127 (N_9127,N_3476,N_4265);
nor U9128 (N_9128,N_4095,N_3282);
nand U9129 (N_9129,N_5302,N_4664);
and U9130 (N_9130,N_5134,N_6190);
nor U9131 (N_9131,N_5494,N_5352);
or U9132 (N_9132,N_4234,N_5986);
and U9133 (N_9133,N_4515,N_4876);
and U9134 (N_9134,N_5876,N_4054);
and U9135 (N_9135,N_3275,N_5356);
nor U9136 (N_9136,N_5779,N_3455);
xnor U9137 (N_9137,N_4957,N_3867);
nor U9138 (N_9138,N_3722,N_3511);
nand U9139 (N_9139,N_5459,N_6097);
and U9140 (N_9140,N_4002,N_3445);
or U9141 (N_9141,N_4095,N_5231);
and U9142 (N_9142,N_5056,N_3645);
nand U9143 (N_9143,N_4170,N_3345);
and U9144 (N_9144,N_3343,N_4059);
nor U9145 (N_9145,N_5504,N_4436);
nand U9146 (N_9146,N_4330,N_6184);
xor U9147 (N_9147,N_4525,N_4276);
nand U9148 (N_9148,N_4457,N_4475);
xor U9149 (N_9149,N_3227,N_4189);
and U9150 (N_9150,N_5455,N_5135);
and U9151 (N_9151,N_4020,N_5976);
xor U9152 (N_9152,N_5056,N_5439);
or U9153 (N_9153,N_4969,N_5597);
or U9154 (N_9154,N_5749,N_3854);
nor U9155 (N_9155,N_3267,N_3316);
nor U9156 (N_9156,N_5469,N_5854);
nor U9157 (N_9157,N_6101,N_5430);
xnor U9158 (N_9158,N_5628,N_4597);
or U9159 (N_9159,N_3356,N_3462);
and U9160 (N_9160,N_4976,N_5652);
nand U9161 (N_9161,N_3213,N_6168);
xor U9162 (N_9162,N_5526,N_3154);
or U9163 (N_9163,N_5094,N_6091);
nand U9164 (N_9164,N_3821,N_6181);
nand U9165 (N_9165,N_5458,N_4356);
and U9166 (N_9166,N_4855,N_4093);
and U9167 (N_9167,N_4063,N_4764);
nor U9168 (N_9168,N_4644,N_3187);
and U9169 (N_9169,N_3144,N_5445);
nand U9170 (N_9170,N_3977,N_4117);
or U9171 (N_9171,N_4374,N_3653);
or U9172 (N_9172,N_3789,N_3938);
nand U9173 (N_9173,N_4831,N_3393);
nand U9174 (N_9174,N_3563,N_3522);
or U9175 (N_9175,N_3592,N_3416);
nor U9176 (N_9176,N_5102,N_6036);
or U9177 (N_9177,N_5829,N_3826);
nand U9178 (N_9178,N_5708,N_5108);
nand U9179 (N_9179,N_5479,N_4505);
nor U9180 (N_9180,N_5865,N_3826);
nor U9181 (N_9181,N_6107,N_3684);
or U9182 (N_9182,N_3873,N_4403);
and U9183 (N_9183,N_5804,N_3222);
nand U9184 (N_9184,N_4036,N_5029);
or U9185 (N_9185,N_4189,N_4019);
nor U9186 (N_9186,N_4716,N_3678);
and U9187 (N_9187,N_5940,N_4356);
or U9188 (N_9188,N_4827,N_4061);
nor U9189 (N_9189,N_4956,N_3744);
nor U9190 (N_9190,N_4231,N_5887);
xor U9191 (N_9191,N_6243,N_4905);
xnor U9192 (N_9192,N_4545,N_4892);
nor U9193 (N_9193,N_3589,N_4492);
xor U9194 (N_9194,N_5535,N_3567);
nor U9195 (N_9195,N_5143,N_3171);
nand U9196 (N_9196,N_5081,N_3470);
or U9197 (N_9197,N_4634,N_6042);
nand U9198 (N_9198,N_5599,N_4149);
xnor U9199 (N_9199,N_3505,N_5795);
and U9200 (N_9200,N_4311,N_3822);
nor U9201 (N_9201,N_5045,N_5623);
xor U9202 (N_9202,N_4410,N_5466);
nor U9203 (N_9203,N_4507,N_5508);
or U9204 (N_9204,N_4826,N_3522);
or U9205 (N_9205,N_3921,N_4035);
or U9206 (N_9206,N_4488,N_5765);
and U9207 (N_9207,N_5489,N_3723);
xnor U9208 (N_9208,N_5009,N_4244);
nand U9209 (N_9209,N_3847,N_5653);
nand U9210 (N_9210,N_6069,N_4305);
or U9211 (N_9211,N_3803,N_5780);
or U9212 (N_9212,N_5002,N_3212);
nor U9213 (N_9213,N_3261,N_3157);
xnor U9214 (N_9214,N_4964,N_4104);
nor U9215 (N_9215,N_3547,N_4695);
xnor U9216 (N_9216,N_3951,N_3632);
nand U9217 (N_9217,N_3990,N_4405);
and U9218 (N_9218,N_3993,N_5595);
nand U9219 (N_9219,N_5222,N_4768);
and U9220 (N_9220,N_3553,N_3501);
nand U9221 (N_9221,N_3699,N_3561);
nand U9222 (N_9222,N_5057,N_5889);
xor U9223 (N_9223,N_5815,N_3760);
nor U9224 (N_9224,N_4176,N_3395);
nor U9225 (N_9225,N_5487,N_5760);
or U9226 (N_9226,N_4339,N_5596);
or U9227 (N_9227,N_4452,N_5842);
xnor U9228 (N_9228,N_6151,N_5088);
and U9229 (N_9229,N_4179,N_3339);
and U9230 (N_9230,N_3254,N_4165);
nor U9231 (N_9231,N_5896,N_3725);
nor U9232 (N_9232,N_3994,N_4913);
nand U9233 (N_9233,N_4804,N_5059);
xor U9234 (N_9234,N_3590,N_4154);
or U9235 (N_9235,N_4760,N_6225);
and U9236 (N_9236,N_6098,N_5268);
xor U9237 (N_9237,N_5067,N_5717);
nand U9238 (N_9238,N_5559,N_4723);
xor U9239 (N_9239,N_4683,N_3723);
nand U9240 (N_9240,N_5718,N_3574);
or U9241 (N_9241,N_5846,N_4574);
or U9242 (N_9242,N_4347,N_4383);
nor U9243 (N_9243,N_5461,N_5121);
or U9244 (N_9244,N_3214,N_3460);
and U9245 (N_9245,N_4127,N_5678);
nand U9246 (N_9246,N_4077,N_3278);
and U9247 (N_9247,N_4283,N_4798);
nor U9248 (N_9248,N_4501,N_4885);
or U9249 (N_9249,N_4186,N_3665);
and U9250 (N_9250,N_3215,N_6108);
nand U9251 (N_9251,N_4521,N_5334);
nor U9252 (N_9252,N_4842,N_3604);
nor U9253 (N_9253,N_4523,N_3856);
nand U9254 (N_9254,N_4680,N_5655);
xnor U9255 (N_9255,N_4947,N_4914);
and U9256 (N_9256,N_3707,N_4643);
nand U9257 (N_9257,N_3865,N_3788);
or U9258 (N_9258,N_4184,N_4639);
nand U9259 (N_9259,N_3234,N_4639);
nor U9260 (N_9260,N_4867,N_6132);
and U9261 (N_9261,N_4849,N_4519);
nor U9262 (N_9262,N_5411,N_4921);
xnor U9263 (N_9263,N_5861,N_3663);
and U9264 (N_9264,N_5615,N_4319);
nand U9265 (N_9265,N_5736,N_4069);
or U9266 (N_9266,N_3901,N_4228);
nor U9267 (N_9267,N_4888,N_5420);
xor U9268 (N_9268,N_6101,N_5558);
nor U9269 (N_9269,N_6070,N_4373);
nor U9270 (N_9270,N_3134,N_5042);
xnor U9271 (N_9271,N_5981,N_3345);
and U9272 (N_9272,N_5035,N_4945);
xnor U9273 (N_9273,N_3581,N_4555);
nand U9274 (N_9274,N_5753,N_5761);
xnor U9275 (N_9275,N_3609,N_5204);
and U9276 (N_9276,N_6223,N_4904);
nand U9277 (N_9277,N_3444,N_4512);
nor U9278 (N_9278,N_5975,N_5013);
nor U9279 (N_9279,N_5514,N_4043);
nand U9280 (N_9280,N_4946,N_4697);
xor U9281 (N_9281,N_3986,N_5289);
xnor U9282 (N_9282,N_3992,N_5781);
nor U9283 (N_9283,N_5964,N_3934);
nor U9284 (N_9284,N_5678,N_3601);
or U9285 (N_9285,N_3616,N_4050);
nand U9286 (N_9286,N_5515,N_4504);
and U9287 (N_9287,N_4579,N_3269);
or U9288 (N_9288,N_4428,N_4291);
nor U9289 (N_9289,N_4657,N_4498);
nor U9290 (N_9290,N_3455,N_6070);
xor U9291 (N_9291,N_3345,N_3889);
nor U9292 (N_9292,N_3321,N_4737);
xnor U9293 (N_9293,N_5976,N_4780);
or U9294 (N_9294,N_6022,N_5721);
and U9295 (N_9295,N_5179,N_3256);
nand U9296 (N_9296,N_5413,N_3776);
and U9297 (N_9297,N_4256,N_3484);
or U9298 (N_9298,N_5151,N_4262);
xnor U9299 (N_9299,N_5413,N_5938);
xnor U9300 (N_9300,N_4995,N_5562);
nand U9301 (N_9301,N_4134,N_3890);
nand U9302 (N_9302,N_5243,N_4966);
xor U9303 (N_9303,N_3628,N_3588);
nand U9304 (N_9304,N_6213,N_4210);
and U9305 (N_9305,N_5614,N_5567);
nand U9306 (N_9306,N_4284,N_3281);
nand U9307 (N_9307,N_4490,N_4656);
or U9308 (N_9308,N_5159,N_4156);
or U9309 (N_9309,N_4595,N_5195);
xor U9310 (N_9310,N_4733,N_5569);
xor U9311 (N_9311,N_4213,N_3507);
or U9312 (N_9312,N_4448,N_4387);
or U9313 (N_9313,N_4071,N_4775);
nand U9314 (N_9314,N_5354,N_4107);
and U9315 (N_9315,N_5165,N_3964);
nor U9316 (N_9316,N_6248,N_5585);
xor U9317 (N_9317,N_3309,N_5463);
or U9318 (N_9318,N_5383,N_4225);
nor U9319 (N_9319,N_3686,N_4029);
nand U9320 (N_9320,N_4404,N_6084);
and U9321 (N_9321,N_3689,N_4820);
and U9322 (N_9322,N_3900,N_3908);
nand U9323 (N_9323,N_4196,N_5100);
nor U9324 (N_9324,N_3975,N_3515);
nor U9325 (N_9325,N_4889,N_6152);
or U9326 (N_9326,N_3831,N_5301);
nor U9327 (N_9327,N_4829,N_4511);
nor U9328 (N_9328,N_4374,N_4623);
xor U9329 (N_9329,N_3339,N_5327);
nand U9330 (N_9330,N_3957,N_4339);
nand U9331 (N_9331,N_4736,N_4263);
nor U9332 (N_9332,N_3347,N_4415);
xnor U9333 (N_9333,N_5442,N_4485);
or U9334 (N_9334,N_3268,N_4364);
and U9335 (N_9335,N_3324,N_4045);
xnor U9336 (N_9336,N_3905,N_6134);
or U9337 (N_9337,N_3201,N_5828);
nor U9338 (N_9338,N_6101,N_4505);
nor U9339 (N_9339,N_6185,N_5267);
nand U9340 (N_9340,N_4005,N_4865);
and U9341 (N_9341,N_6176,N_4517);
xnor U9342 (N_9342,N_3233,N_5593);
nand U9343 (N_9343,N_6032,N_4000);
xor U9344 (N_9344,N_5477,N_5330);
and U9345 (N_9345,N_5670,N_5484);
or U9346 (N_9346,N_6052,N_4922);
or U9347 (N_9347,N_3678,N_4955);
nand U9348 (N_9348,N_5088,N_6206);
xor U9349 (N_9349,N_3590,N_4042);
xor U9350 (N_9350,N_3671,N_5242);
nor U9351 (N_9351,N_3958,N_4600);
and U9352 (N_9352,N_3326,N_3506);
xnor U9353 (N_9353,N_4643,N_3612);
and U9354 (N_9354,N_3739,N_5966);
nand U9355 (N_9355,N_5968,N_6174);
or U9356 (N_9356,N_5235,N_4686);
nand U9357 (N_9357,N_4305,N_5433);
nand U9358 (N_9358,N_4972,N_4821);
xor U9359 (N_9359,N_3449,N_3633);
and U9360 (N_9360,N_3245,N_5409);
nand U9361 (N_9361,N_3907,N_4366);
nor U9362 (N_9362,N_3374,N_4746);
nor U9363 (N_9363,N_5965,N_5971);
or U9364 (N_9364,N_3172,N_4303);
nor U9365 (N_9365,N_6074,N_3844);
nor U9366 (N_9366,N_3641,N_5598);
nand U9367 (N_9367,N_4108,N_3338);
xnor U9368 (N_9368,N_5094,N_3312);
nand U9369 (N_9369,N_5144,N_4919);
xnor U9370 (N_9370,N_5586,N_4755);
and U9371 (N_9371,N_4764,N_5064);
and U9372 (N_9372,N_3528,N_5225);
and U9373 (N_9373,N_4479,N_5529);
nand U9374 (N_9374,N_6077,N_4943);
or U9375 (N_9375,N_6970,N_7052);
xor U9376 (N_9376,N_6989,N_6565);
nor U9377 (N_9377,N_8256,N_7347);
or U9378 (N_9378,N_7433,N_8126);
nor U9379 (N_9379,N_7521,N_6526);
or U9380 (N_9380,N_6991,N_7951);
nor U9381 (N_9381,N_6608,N_6457);
nand U9382 (N_9382,N_7535,N_8516);
nor U9383 (N_9383,N_8506,N_7050);
nor U9384 (N_9384,N_8578,N_9197);
nand U9385 (N_9385,N_8370,N_6821);
and U9386 (N_9386,N_6403,N_7306);
xnor U9387 (N_9387,N_6997,N_7839);
nand U9388 (N_9388,N_9179,N_6424);
xnor U9389 (N_9389,N_8858,N_7658);
and U9390 (N_9390,N_7810,N_7972);
or U9391 (N_9391,N_8231,N_8441);
and U9392 (N_9392,N_7547,N_7943);
or U9393 (N_9393,N_7320,N_7073);
nor U9394 (N_9394,N_6305,N_9107);
or U9395 (N_9395,N_8605,N_7388);
or U9396 (N_9396,N_6472,N_7575);
nor U9397 (N_9397,N_6840,N_8208);
xor U9398 (N_9398,N_7471,N_7754);
and U9399 (N_9399,N_8016,N_8435);
or U9400 (N_9400,N_6292,N_8127);
and U9401 (N_9401,N_7265,N_7363);
or U9402 (N_9402,N_7768,N_7239);
and U9403 (N_9403,N_8650,N_8010);
nor U9404 (N_9404,N_6841,N_8012);
and U9405 (N_9405,N_7713,N_6889);
nand U9406 (N_9406,N_7967,N_8270);
or U9407 (N_9407,N_6916,N_8026);
or U9408 (N_9408,N_8508,N_6771);
nand U9409 (N_9409,N_9183,N_8096);
nand U9410 (N_9410,N_9041,N_7062);
and U9411 (N_9411,N_7715,N_7984);
nor U9412 (N_9412,N_6559,N_8389);
or U9413 (N_9413,N_9206,N_6700);
xor U9414 (N_9414,N_7534,N_8613);
or U9415 (N_9415,N_7877,N_7409);
xnor U9416 (N_9416,N_8303,N_7036);
nand U9417 (N_9417,N_8369,N_7915);
xor U9418 (N_9418,N_7725,N_8897);
nand U9419 (N_9419,N_6844,N_9029);
nand U9420 (N_9420,N_8192,N_8057);
or U9421 (N_9421,N_6571,N_8986);
and U9422 (N_9422,N_9344,N_8065);
or U9423 (N_9423,N_8299,N_8220);
nand U9424 (N_9424,N_6733,N_9028);
nor U9425 (N_9425,N_6585,N_9103);
nand U9426 (N_9426,N_6256,N_7517);
xor U9427 (N_9427,N_8950,N_7743);
nor U9428 (N_9428,N_7757,N_9118);
or U9429 (N_9429,N_8836,N_6389);
xor U9430 (N_9430,N_9262,N_7790);
nand U9431 (N_9431,N_6765,N_7490);
xnor U9432 (N_9432,N_7702,N_8527);
or U9433 (N_9433,N_6373,N_7663);
or U9434 (N_9434,N_8367,N_7950);
nand U9435 (N_9435,N_8839,N_8318);
or U9436 (N_9436,N_7598,N_8904);
nand U9437 (N_9437,N_7314,N_9355);
nand U9438 (N_9438,N_9369,N_6544);
nand U9439 (N_9439,N_7304,N_8482);
xor U9440 (N_9440,N_7612,N_9132);
xnor U9441 (N_9441,N_9190,N_8088);
and U9442 (N_9442,N_7910,N_6774);
nor U9443 (N_9443,N_7188,N_7551);
nand U9444 (N_9444,N_6802,N_6390);
or U9445 (N_9445,N_8619,N_6607);
or U9446 (N_9446,N_8624,N_6393);
or U9447 (N_9447,N_6582,N_9311);
nor U9448 (N_9448,N_8463,N_7643);
nor U9449 (N_9449,N_7220,N_6461);
xnor U9450 (N_9450,N_8887,N_7580);
nor U9451 (N_9451,N_7684,N_7311);
xor U9452 (N_9452,N_8908,N_7396);
or U9453 (N_9453,N_9181,N_8432);
nand U9454 (N_9454,N_8414,N_7690);
and U9455 (N_9455,N_6353,N_7708);
nand U9456 (N_9456,N_8522,N_6745);
and U9457 (N_9457,N_8067,N_7548);
and U9458 (N_9458,N_9034,N_7406);
xor U9459 (N_9459,N_7894,N_6254);
nor U9460 (N_9460,N_7461,N_8959);
or U9461 (N_9461,N_8981,N_7432);
or U9462 (N_9462,N_8562,N_8309);
nor U9463 (N_9463,N_8938,N_8147);
xnor U9464 (N_9464,N_7722,N_6614);
nand U9465 (N_9465,N_8680,N_8278);
and U9466 (N_9466,N_7288,N_6788);
nor U9467 (N_9467,N_7519,N_8968);
nand U9468 (N_9468,N_7329,N_7402);
and U9469 (N_9469,N_8448,N_6799);
nor U9470 (N_9470,N_8829,N_9076);
nand U9471 (N_9471,N_8780,N_8891);
xor U9472 (N_9472,N_7589,N_7358);
xnor U9473 (N_9473,N_9020,N_9175);
nor U9474 (N_9474,N_8238,N_7023);
nand U9475 (N_9475,N_8329,N_8461);
and U9476 (N_9476,N_6302,N_7908);
and U9477 (N_9477,N_6801,N_7555);
or U9478 (N_9478,N_6708,N_6832);
nor U9479 (N_9479,N_7446,N_7227);
and U9480 (N_9480,N_6674,N_7544);
and U9481 (N_9481,N_7980,N_8116);
nor U9482 (N_9482,N_6739,N_6994);
nor U9483 (N_9483,N_7451,N_9298);
and U9484 (N_9484,N_6428,N_7107);
xor U9485 (N_9485,N_6271,N_6906);
nor U9486 (N_9486,N_6812,N_9343);
and U9487 (N_9487,N_9053,N_6400);
nor U9488 (N_9488,N_7818,N_7405);
nand U9489 (N_9489,N_7136,N_9300);
and U9490 (N_9490,N_9224,N_7398);
nor U9491 (N_9491,N_9297,N_7862);
or U9492 (N_9492,N_8323,N_7775);
nor U9493 (N_9493,N_6993,N_7918);
xor U9494 (N_9494,N_6817,N_8315);
nor U9495 (N_9495,N_6318,N_8085);
xnor U9496 (N_9496,N_7841,N_6646);
and U9497 (N_9497,N_7459,N_6277);
xnor U9498 (N_9498,N_7070,N_8027);
and U9499 (N_9499,N_8269,N_9160);
nand U9500 (N_9500,N_7428,N_8159);
nor U9501 (N_9501,N_8852,N_9372);
nor U9502 (N_9502,N_8856,N_8226);
or U9503 (N_9503,N_8433,N_7099);
nand U9504 (N_9504,N_7009,N_9255);
and U9505 (N_9505,N_6877,N_8348);
and U9506 (N_9506,N_6554,N_7816);
or U9507 (N_9507,N_6550,N_6787);
and U9508 (N_9508,N_8091,N_7112);
or U9509 (N_9509,N_8087,N_9258);
or U9510 (N_9510,N_6866,N_8290);
and U9511 (N_9511,N_8342,N_9239);
or U9512 (N_9512,N_8951,N_7527);
xor U9513 (N_9513,N_9229,N_6705);
and U9514 (N_9514,N_8177,N_7282);
and U9515 (N_9515,N_9205,N_6820);
or U9516 (N_9516,N_7257,N_8014);
nand U9517 (N_9517,N_7254,N_8265);
nor U9518 (N_9518,N_8036,N_8563);
nand U9519 (N_9519,N_8374,N_7148);
nand U9520 (N_9520,N_6307,N_8148);
nor U9521 (N_9521,N_7292,N_7305);
or U9522 (N_9522,N_7732,N_9138);
and U9523 (N_9523,N_8292,N_8074);
xor U9524 (N_9524,N_6931,N_8927);
and U9525 (N_9525,N_8687,N_6426);
nor U9526 (N_9526,N_7939,N_8121);
or U9527 (N_9527,N_8102,N_6322);
or U9528 (N_9528,N_8417,N_8412);
and U9529 (N_9529,N_7120,N_8330);
and U9530 (N_9530,N_7701,N_6859);
xor U9531 (N_9531,N_8577,N_6609);
and U9532 (N_9532,N_8281,N_6885);
or U9533 (N_9533,N_7932,N_8449);
and U9534 (N_9534,N_8550,N_6464);
xnor U9535 (N_9535,N_8013,N_8149);
or U9536 (N_9536,N_6943,N_9188);
nor U9537 (N_9537,N_7577,N_7380);
and U9538 (N_9538,N_6896,N_9358);
or U9539 (N_9539,N_9238,N_7024);
and U9540 (N_9540,N_6498,N_7889);
nor U9541 (N_9541,N_6502,N_9135);
nor U9542 (N_9542,N_6706,N_6427);
or U9543 (N_9543,N_7210,N_6589);
nand U9544 (N_9544,N_9125,N_7677);
nand U9545 (N_9545,N_7049,N_6932);
and U9546 (N_9546,N_8795,N_7770);
nand U9547 (N_9547,N_7455,N_9222);
xor U9548 (N_9548,N_7840,N_8545);
xnor U9549 (N_9549,N_6783,N_8287);
nand U9550 (N_9550,N_8728,N_8967);
xnor U9551 (N_9551,N_8398,N_8403);
and U9552 (N_9552,N_8109,N_7977);
xor U9553 (N_9553,N_8353,N_8125);
or U9554 (N_9554,N_7376,N_7198);
xor U9555 (N_9555,N_8289,N_6267);
and U9556 (N_9556,N_9352,N_7742);
and U9557 (N_9557,N_9346,N_8168);
or U9558 (N_9558,N_6386,N_8727);
nor U9559 (N_9559,N_8978,N_6779);
nand U9560 (N_9560,N_8068,N_6772);
xor U9561 (N_9561,N_6310,N_8646);
xor U9562 (N_9562,N_8870,N_6450);
xnor U9563 (N_9563,N_8260,N_6722);
or U9564 (N_9564,N_8296,N_8800);
nor U9565 (N_9565,N_8692,N_7445);
or U9566 (N_9566,N_7130,N_6874);
nand U9567 (N_9567,N_7844,N_7161);
nand U9568 (N_9568,N_6637,N_7243);
xor U9569 (N_9569,N_6830,N_8133);
nand U9570 (N_9570,N_6304,N_8247);
xnor U9571 (N_9571,N_8561,N_8002);
and U9572 (N_9572,N_8751,N_6444);
xor U9573 (N_9573,N_7875,N_7258);
xor U9574 (N_9574,N_6378,N_8718);
nand U9575 (N_9575,N_8962,N_7072);
and U9576 (N_9576,N_8612,N_7786);
and U9577 (N_9577,N_8537,N_6561);
nor U9578 (N_9578,N_6639,N_8783);
xor U9579 (N_9579,N_8314,N_7595);
nor U9580 (N_9580,N_9214,N_8975);
nand U9581 (N_9581,N_7805,N_7156);
nor U9582 (N_9582,N_8379,N_7484);
nand U9583 (N_9583,N_8570,N_8475);
xnor U9584 (N_9584,N_8976,N_6795);
nor U9585 (N_9585,N_9072,N_6456);
nor U9586 (N_9586,N_6953,N_8110);
nor U9587 (N_9587,N_9147,N_7689);
xnor U9588 (N_9588,N_7730,N_6417);
nand U9589 (N_9589,N_6868,N_6837);
or U9590 (N_9590,N_7695,N_7229);
and U9591 (N_9591,N_7522,N_6928);
nand U9592 (N_9592,N_8693,N_7675);
xor U9593 (N_9593,N_9231,N_7105);
and U9594 (N_9594,N_8726,N_6591);
or U9595 (N_9595,N_7495,N_7221);
nor U9596 (N_9596,N_9130,N_9023);
xor U9597 (N_9597,N_6748,N_7182);
or U9598 (N_9598,N_7041,N_7942);
xor U9599 (N_9599,N_6915,N_6769);
or U9600 (N_9600,N_6429,N_7191);
xor U9601 (N_9601,N_7529,N_8305);
nand U9602 (N_9602,N_8668,N_7546);
xor U9603 (N_9603,N_6368,N_7435);
xor U9604 (N_9604,N_9292,N_7333);
nand U9605 (N_9605,N_6335,N_6734);
xor U9606 (N_9606,N_6881,N_6296);
nor U9607 (N_9607,N_6852,N_7491);
nor U9608 (N_9608,N_7679,N_8006);
nand U9609 (N_9609,N_8437,N_6621);
xor U9610 (N_9610,N_7170,N_7625);
or U9611 (N_9611,N_7033,N_8682);
nand U9612 (N_9612,N_8551,N_7671);
nor U9613 (N_9613,N_9254,N_8798);
xnor U9614 (N_9614,N_9095,N_7566);
nand U9615 (N_9615,N_8890,N_6553);
and U9616 (N_9616,N_7332,N_8984);
xnor U9617 (N_9617,N_6491,N_9054);
or U9618 (N_9618,N_7798,N_8411);
nor U9619 (N_9619,N_7113,N_7357);
or U9620 (N_9620,N_6983,N_7879);
and U9621 (N_9621,N_8332,N_8038);
and U9622 (N_9622,N_9289,N_8529);
xor U9623 (N_9623,N_9021,N_7056);
nand U9624 (N_9624,N_9275,N_7134);
nand U9625 (N_9625,N_8106,N_7848);
nor U9626 (N_9626,N_6898,N_6675);
nand U9627 (N_9627,N_7460,N_7454);
or U9628 (N_9628,N_8644,N_6873);
and U9629 (N_9629,N_7241,N_7694);
nand U9630 (N_9630,N_8215,N_6807);
nor U9631 (N_9631,N_9320,N_6397);
nor U9632 (N_9632,N_7525,N_8966);
or U9633 (N_9633,N_7814,N_8567);
and U9634 (N_9634,N_6670,N_6616);
or U9635 (N_9635,N_9245,N_8846);
or U9636 (N_9636,N_9265,N_7583);
or U9637 (N_9637,N_8430,N_7307);
or U9638 (N_9638,N_8917,N_8213);
nor U9639 (N_9639,N_7321,N_7652);
nor U9640 (N_9640,N_8381,N_6694);
nand U9641 (N_9641,N_7334,N_8320);
or U9642 (N_9642,N_8474,N_7738);
and U9643 (N_9643,N_8672,N_6262);
and U9644 (N_9644,N_8029,N_8883);
nand U9645 (N_9645,N_6252,N_7882);
and U9646 (N_9646,N_6793,N_8053);
nor U9647 (N_9647,N_8408,N_7610);
xor U9648 (N_9648,N_6366,N_7385);
or U9649 (N_9649,N_8046,N_7956);
nand U9650 (N_9650,N_8351,N_8054);
nor U9651 (N_9651,N_8392,N_9000);
nor U9652 (N_9652,N_9060,N_6319);
or U9653 (N_9653,N_9003,N_8399);
or U9654 (N_9654,N_8872,N_8997);
and U9655 (N_9655,N_8770,N_6336);
or U9656 (N_9656,N_8600,N_7739);
or U9657 (N_9657,N_8180,N_7801);
nor U9658 (N_9658,N_7408,N_8214);
and U9659 (N_9659,N_7181,N_7955);
or U9660 (N_9660,N_8443,N_6798);
or U9661 (N_9661,N_8191,N_8140);
and U9662 (N_9662,N_7237,N_8349);
and U9663 (N_9663,N_9074,N_7791);
xor U9664 (N_9664,N_8530,N_6510);
nor U9665 (N_9665,N_8813,N_7760);
nor U9666 (N_9666,N_8120,N_6941);
or U9667 (N_9667,N_8945,N_6937);
xor U9668 (N_9668,N_8297,N_7604);
nand U9669 (N_9669,N_6405,N_8683);
or U9670 (N_9670,N_7046,N_7693);
or U9671 (N_9671,N_8676,N_9194);
or U9672 (N_9672,N_7174,N_7236);
and U9673 (N_9673,N_8009,N_8113);
xor U9674 (N_9674,N_7748,N_7717);
xor U9675 (N_9675,N_6693,N_8244);
or U9676 (N_9676,N_7395,N_8902);
nand U9677 (N_9677,N_6263,N_9221);
and U9678 (N_9678,N_7820,N_8181);
xor U9679 (N_9679,N_6908,N_7800);
and U9680 (N_9680,N_7883,N_8509);
nand U9681 (N_9681,N_7920,N_7361);
xor U9682 (N_9682,N_8769,N_7963);
xnor U9683 (N_9683,N_7999,N_8937);
xor U9684 (N_9684,N_7971,N_9088);
nor U9685 (N_9685,N_9014,N_7531);
xnor U9686 (N_9686,N_8434,N_9007);
xor U9687 (N_9687,N_9022,N_8920);
nor U9688 (N_9688,N_7602,N_6938);
nand U9689 (N_9689,N_8584,N_6831);
xor U9690 (N_9690,N_6264,N_8341);
xnor U9691 (N_9691,N_8531,N_6914);
and U9692 (N_9692,N_7470,N_6580);
or U9693 (N_9693,N_8190,N_6986);
xor U9694 (N_9694,N_9235,N_6392);
xnor U9695 (N_9695,N_8631,N_7520);
nor U9696 (N_9696,N_8785,N_6624);
nand U9697 (N_9697,N_8943,N_8973);
and U9698 (N_9698,N_7208,N_7144);
nand U9699 (N_9699,N_8576,N_6724);
nor U9700 (N_9700,N_8055,N_9167);
nor U9701 (N_9701,N_7988,N_8729);
and U9702 (N_9702,N_8024,N_7620);
or U9703 (N_9703,N_8716,N_9069);
nand U9704 (N_9704,N_8402,N_6568);
nand U9705 (N_9705,N_7897,N_7947);
nor U9706 (N_9706,N_6268,N_7945);
or U9707 (N_9707,N_7765,N_9274);
xor U9708 (N_9708,N_7084,N_9329);
nor U9709 (N_9709,N_9256,N_9087);
and U9710 (N_9710,N_8581,N_8542);
xor U9711 (N_9711,N_6473,N_6488);
or U9712 (N_9712,N_9001,N_7680);
nor U9713 (N_9713,N_7735,N_8094);
nand U9714 (N_9714,N_7092,N_6261);
and U9715 (N_9715,N_8099,N_8788);
nand U9716 (N_9716,N_7167,N_6570);
nand U9717 (N_9717,N_8456,N_7186);
and U9718 (N_9718,N_7886,N_6363);
nand U9719 (N_9719,N_7344,N_7507);
or U9720 (N_9720,N_6757,N_6376);
xor U9721 (N_9721,N_8607,N_6564);
and U9722 (N_9722,N_8525,N_7256);
and U9723 (N_9723,N_8655,N_7606);
or U9724 (N_9724,N_8665,N_8784);
nand U9725 (N_9725,N_7280,N_8538);
nor U9726 (N_9726,N_6423,N_9127);
and U9727 (N_9727,N_6442,N_7086);
nand U9728 (N_9728,N_7506,N_7633);
nand U9729 (N_9729,N_6250,N_6809);
or U9730 (N_9730,N_7763,N_8480);
nor U9731 (N_9731,N_9064,N_8257);
nand U9732 (N_9732,N_8926,N_8589);
nor U9733 (N_9733,N_7532,N_8383);
nor U9734 (N_9734,N_8130,N_6573);
and U9735 (N_9735,N_9108,N_6518);
and U9736 (N_9736,N_7636,N_7345);
nand U9737 (N_9737,N_8949,N_9178);
nor U9738 (N_9738,N_8558,N_9185);
or U9739 (N_9739,N_7493,N_9144);
and U9740 (N_9740,N_6810,N_6800);
and U9741 (N_9741,N_6851,N_8160);
nor U9742 (N_9742,N_8464,N_8850);
xnor U9743 (N_9743,N_8272,N_6715);
xor U9744 (N_9744,N_7071,N_6576);
nor U9745 (N_9745,N_7869,N_7803);
and U9746 (N_9746,N_9247,N_8156);
or U9747 (N_9747,N_8178,N_8071);
and U9748 (N_9748,N_7199,N_6910);
and U9749 (N_9749,N_7326,N_6729);
xnor U9750 (N_9750,N_7603,N_8965);
xor U9751 (N_9751,N_6952,N_6834);
nand U9752 (N_9752,N_9038,N_6445);
nand U9753 (N_9753,N_7691,N_6432);
nand U9754 (N_9754,N_8944,N_7704);
nand U9755 (N_9755,N_6773,N_6301);
nor U9756 (N_9756,N_9191,N_6947);
nand U9757 (N_9757,N_9211,N_6628);
nand U9758 (N_9758,N_6719,N_6477);
nor U9759 (N_9759,N_7218,N_7660);
and U9760 (N_9760,N_6543,N_7838);
and U9761 (N_9761,N_7245,N_6449);
nor U9762 (N_9762,N_7211,N_9075);
or U9763 (N_9763,N_8371,N_6777);
and U9764 (N_9764,N_7876,N_7027);
xnor U9765 (N_9765,N_6468,N_9286);
xnor U9766 (N_9766,N_8812,N_6383);
nor U9767 (N_9767,N_8235,N_9137);
nor U9768 (N_9768,N_8117,N_8892);
or U9769 (N_9769,N_7152,N_7489);
or U9770 (N_9770,N_6805,N_7362);
or U9771 (N_9771,N_7251,N_9171);
nand U9772 (N_9772,N_9315,N_8360);
nor U9773 (N_9773,N_8819,N_8947);
and U9774 (N_9774,N_7647,N_8462);
xor U9775 (N_9775,N_8285,N_7697);
and U9776 (N_9776,N_7543,N_7346);
and U9777 (N_9777,N_6845,N_9249);
and U9778 (N_9778,N_6667,N_9362);
nand U9779 (N_9779,N_6594,N_8263);
and U9780 (N_9780,N_6326,N_8789);
nor U9781 (N_9781,N_8521,N_7442);
and U9782 (N_9782,N_8999,N_6826);
nor U9783 (N_9783,N_7412,N_7809);
nor U9784 (N_9784,N_6982,N_8514);
and U9785 (N_9785,N_8877,N_8152);
and U9786 (N_9786,N_9328,N_9264);
xnor U9787 (N_9787,N_7976,N_8439);
nor U9788 (N_9788,N_9105,N_6630);
nor U9789 (N_9789,N_6520,N_7119);
xnor U9790 (N_9790,N_8206,N_7067);
xor U9791 (N_9791,N_6521,N_7673);
or U9792 (N_9792,N_6925,N_8750);
xor U9793 (N_9793,N_7145,N_6285);
nor U9794 (N_9794,N_6598,N_7540);
and U9795 (N_9795,N_7802,N_6406);
or U9796 (N_9796,N_8598,N_8782);
or U9797 (N_9797,N_9078,N_8141);
nor U9798 (N_9798,N_7002,N_7638);
nor U9799 (N_9799,N_8566,N_8466);
nor U9800 (N_9800,N_6590,N_6360);
nand U9801 (N_9801,N_8834,N_6725);
and U9802 (N_9802,N_7271,N_8145);
xor U9803 (N_9803,N_8188,N_8405);
nand U9804 (N_9804,N_6934,N_7858);
or U9805 (N_9805,N_7749,N_7808);
nand U9806 (N_9806,N_7094,N_7389);
nor U9807 (N_9807,N_9187,N_6981);
nor U9808 (N_9808,N_7761,N_8478);
xnor U9809 (N_9809,N_8195,N_6505);
xnor U9810 (N_9810,N_7659,N_6574);
or U9811 (N_9811,N_9192,N_8520);
nand U9812 (N_9812,N_8988,N_7505);
and U9813 (N_9813,N_6610,N_6901);
and U9814 (N_9814,N_7857,N_7822);
xnor U9815 (N_9815,N_8889,N_7157);
nand U9816 (N_9816,N_6944,N_7449);
xor U9817 (N_9817,N_7642,N_7275);
and U9818 (N_9818,N_7514,N_8990);
nor U9819 (N_9819,N_6340,N_7232);
xnor U9820 (N_9820,N_6897,N_9252);
xnor U9821 (N_9821,N_7905,N_8946);
nor U9822 (N_9822,N_7965,N_8445);
xor U9823 (N_9823,N_6471,N_7752);
or U9824 (N_9824,N_9036,N_6888);
or U9825 (N_9825,N_7404,N_7424);
xnor U9826 (N_9826,N_8479,N_6465);
nand U9827 (N_9827,N_8450,N_6287);
or U9828 (N_9828,N_8543,N_6726);
nor U9829 (N_9829,N_7795,N_6882);
and U9830 (N_9830,N_7121,N_6635);
nor U9831 (N_9831,N_9120,N_8234);
nor U9832 (N_9832,N_7095,N_8991);
or U9833 (N_9833,N_8752,N_8875);
and U9834 (N_9834,N_8239,N_9314);
or U9835 (N_9835,N_7244,N_8051);
and U9836 (N_9836,N_7515,N_6718);
xor U9837 (N_9837,N_7213,N_7194);
nand U9838 (N_9838,N_8579,N_6454);
nor U9839 (N_9839,N_8034,N_7758);
or U9840 (N_9840,N_7954,N_7437);
nor U9841 (N_9841,N_6509,N_8699);
xnor U9842 (N_9842,N_6525,N_7931);
nor U9843 (N_9843,N_6824,N_9334);
xor U9844 (N_9844,N_6819,N_9032);
nor U9845 (N_9845,N_8721,N_7327);
and U9846 (N_9846,N_7526,N_7622);
and U9847 (N_9847,N_7196,N_7202);
xor U9848 (N_9848,N_8922,N_7709);
nor U9849 (N_9849,N_7681,N_7200);
nand U9850 (N_9850,N_7175,N_7026);
nor U9851 (N_9851,N_9345,N_7193);
nand U9852 (N_9852,N_9004,N_7981);
and U9853 (N_9853,N_6902,N_6522);
nand U9854 (N_9854,N_8841,N_6459);
or U9855 (N_9855,N_7089,N_6391);
and U9856 (N_9856,N_6593,N_7578);
or U9857 (N_9857,N_7590,N_7093);
or U9858 (N_9858,N_8523,N_7537);
and U9859 (N_9859,N_8809,N_8778);
xor U9860 (N_9860,N_6741,N_8838);
or U9861 (N_9861,N_8736,N_9272);
nand U9862 (N_9862,N_6968,N_7350);
and U9863 (N_9863,N_6462,N_8686);
nand U9864 (N_9864,N_7287,N_6778);
xnor U9865 (N_9865,N_6999,N_7594);
and U9866 (N_9866,N_8730,N_8048);
or U9867 (N_9867,N_8958,N_7911);
nor U9868 (N_9868,N_8703,N_6766);
nand U9869 (N_9869,N_6927,N_7368);
nor U9870 (N_9870,N_7055,N_6723);
nor U9871 (N_9871,N_8105,N_8316);
nor U9872 (N_9872,N_6316,N_7315);
nor U9873 (N_9873,N_8483,N_9037);
or U9874 (N_9874,N_7541,N_6499);
or U9875 (N_9875,N_8503,N_6364);
xor U9876 (N_9876,N_7452,N_7846);
xnor U9877 (N_9877,N_6453,N_6415);
xnor U9878 (N_9878,N_6697,N_8867);
or U9879 (N_9879,N_8669,N_8063);
or U9880 (N_9880,N_9295,N_7630);
nand U9881 (N_9881,N_6344,N_8821);
nand U9882 (N_9882,N_7466,N_7946);
or U9883 (N_9883,N_7895,N_7478);
and U9884 (N_9884,N_6649,N_8108);
and U9885 (N_9885,N_7366,N_9267);
and U9886 (N_9886,N_6286,N_9098);
and U9887 (N_9887,N_6290,N_7925);
or U9888 (N_9888,N_8884,N_6780);
nor U9889 (N_9889,N_9109,N_7599);
xnor U9890 (N_9890,N_8336,N_8617);
nor U9891 (N_9891,N_8232,N_7994);
and U9892 (N_9892,N_8842,N_6679);
and U9893 (N_9893,N_6822,N_8851);
nor U9894 (N_9894,N_6992,N_9101);
or U9895 (N_9895,N_7860,N_9006);
xor U9896 (N_9896,N_8324,N_9136);
nor U9897 (N_9897,N_6904,N_8725);
nor U9898 (N_9898,N_6848,N_9073);
and U9899 (N_9899,N_8095,N_7140);
xnor U9900 (N_9900,N_6379,N_7836);
and U9901 (N_9901,N_7153,N_7160);
or U9902 (N_9902,N_9335,N_6698);
nor U9903 (N_9903,N_7195,N_9308);
or U9904 (N_9904,N_8555,N_8781);
nor U9905 (N_9905,N_7785,N_8761);
and U9906 (N_9906,N_6654,N_7135);
and U9907 (N_9907,N_8069,N_8447);
xnor U9908 (N_9908,N_7444,N_7898);
and U9909 (N_9909,N_6517,N_6660);
or U9910 (N_9910,N_7664,N_7300);
and U9911 (N_9911,N_9047,N_6496);
nor U9912 (N_9912,N_8128,N_7169);
nand U9913 (N_9913,N_6681,N_6349);
and U9914 (N_9914,N_9112,N_8240);
xnor U9915 (N_9915,N_7118,N_8322);
nor U9916 (N_9916,N_6878,N_8203);
and U9917 (N_9917,N_7295,N_7128);
or U9918 (N_9918,N_7019,N_8657);
nand U9919 (N_9919,N_7267,N_8086);
and U9920 (N_9920,N_8899,N_8334);
or U9921 (N_9921,N_7631,N_7777);
nor U9922 (N_9922,N_8107,N_6601);
xnor U9923 (N_9923,N_9157,N_7386);
nand U9924 (N_9924,N_8608,N_7783);
xor U9925 (N_9925,N_7823,N_7081);
nand U9926 (N_9926,N_9097,N_8974);
xor U9927 (N_9927,N_7392,N_7774);
xor U9928 (N_9928,N_7276,N_7228);
nand U9929 (N_9929,N_6343,N_8539);
and U9930 (N_9930,N_8039,N_6659);
and U9931 (N_9931,N_6892,N_9261);
and U9932 (N_9932,N_7274,N_7917);
nor U9933 (N_9933,N_7958,N_8419);
and U9934 (N_9934,N_7780,N_8259);
nand U9935 (N_9935,N_7640,N_9042);
and U9936 (N_9936,N_8136,N_7427);
and U9937 (N_9937,N_8460,N_7252);
nand U9938 (N_9938,N_7807,N_7183);
nor U9939 (N_9939,N_6644,N_8066);
or U9940 (N_9940,N_6838,N_7789);
xor U9941 (N_9941,N_6548,N_6480);
xor U9942 (N_9942,N_8252,N_8873);
nand U9943 (N_9943,N_6519,N_7331);
nand U9944 (N_9944,N_8745,N_7676);
or U9945 (N_9945,N_7813,N_8254);
or U9946 (N_9946,N_7685,N_8942);
xnor U9947 (N_9947,N_8266,N_8878);
nor U9948 (N_9948,N_7114,N_6476);
xor U9949 (N_9949,N_6662,N_7013);
and U9950 (N_9950,N_9146,N_9019);
or U9951 (N_9951,N_8654,N_7063);
or U9952 (N_9952,N_7762,N_6361);
nand U9953 (N_9953,N_6926,N_8407);
nand U9954 (N_9954,N_8413,N_7080);
nor U9955 (N_9955,N_7400,N_8355);
nand U9956 (N_9956,N_7234,N_7117);
and U9957 (N_9957,N_7421,N_7097);
or U9958 (N_9958,N_8723,N_7277);
and U9959 (N_9959,N_8596,N_7687);
and U9960 (N_9960,N_6437,N_7716);
xnor U9961 (N_9961,N_6864,N_6358);
xnor U9962 (N_9962,N_6586,N_9198);
xnor U9963 (N_9963,N_8092,N_7264);
or U9964 (N_9964,N_9326,N_7581);
nor U9965 (N_9965,N_7045,N_9133);
xor U9966 (N_9966,N_7644,N_9296);
or U9967 (N_9967,N_8817,N_6900);
or U9968 (N_9968,N_8688,N_6996);
xnor U9969 (N_9969,N_7083,N_7989);
nor U9970 (N_9970,N_7974,N_7782);
xnor U9971 (N_9971,N_8642,N_8993);
nor U9972 (N_9972,N_8298,N_9357);
xnor U9973 (N_9973,N_6751,N_7667);
xor U9974 (N_9974,N_8910,N_7504);
and U9975 (N_9975,N_6651,N_7012);
or U9976 (N_9976,N_7718,N_9143);
and U9977 (N_9977,N_6818,N_8440);
nor U9978 (N_9978,N_8896,N_7465);
and U9979 (N_9979,N_9177,N_6854);
nand U9980 (N_9980,N_6833,N_7563);
and U9981 (N_9981,N_7149,N_7711);
nor U9982 (N_9982,N_8713,N_8429);
nor U9983 (N_9983,N_7596,N_7440);
or U9984 (N_9984,N_7492,N_8603);
and U9985 (N_9985,N_9280,N_7057);
and U9986 (N_9986,N_7370,N_9307);
xor U9987 (N_9987,N_6713,N_8345);
nand U9988 (N_9988,N_6678,N_7082);
xor U9989 (N_9989,N_8708,N_7008);
xnor U9990 (N_9990,N_7884,N_7616);
nand U9991 (N_9991,N_8532,N_7413);
or U9992 (N_9992,N_8459,N_8758);
and U9993 (N_9993,N_8914,N_8187);
and U9994 (N_9994,N_8465,N_6270);
xnor U9995 (N_9995,N_7896,N_6792);
or U9996 (N_9996,N_6388,N_7137);
or U9997 (N_9997,N_8643,N_8473);
nand U9998 (N_9998,N_7666,N_7438);
or U9999 (N_9999,N_7289,N_8925);
xor U10000 (N_10000,N_9070,N_7078);
or U10001 (N_10001,N_9318,N_8866);
and U10002 (N_10002,N_8909,N_8489);
xnor U10003 (N_10003,N_8743,N_9067);
or U10004 (N_10004,N_6746,N_8007);
xnor U10005 (N_10005,N_9119,N_8673);
and U10006 (N_10006,N_8056,N_8797);
nor U10007 (N_10007,N_8000,N_8248);
nand U10008 (N_10008,N_7011,N_8755);
or U10009 (N_10009,N_9354,N_8649);
nand U10010 (N_10010,N_8043,N_8313);
xnor U10011 (N_10011,N_8295,N_6419);
or U10012 (N_10012,N_7255,N_7374);
or U10013 (N_10013,N_8470,N_6321);
nor U10014 (N_10014,N_6860,N_8157);
or U10015 (N_10015,N_7731,N_6375);
and U10016 (N_10016,N_7048,N_7230);
or U10017 (N_10017,N_8933,N_8559);
nor U10018 (N_10018,N_8634,N_8241);
nor U10019 (N_10019,N_8327,N_7556);
nor U10020 (N_10020,N_7674,N_7284);
nand U10021 (N_10021,N_6727,N_6796);
xnor U10022 (N_10022,N_8495,N_7554);
xor U10023 (N_10023,N_7605,N_8662);
nor U10024 (N_10024,N_8201,N_8319);
or U10025 (N_10025,N_8622,N_8580);
nand U10026 (N_10026,N_6876,N_8142);
and U10027 (N_10027,N_8825,N_7190);
nand U10028 (N_10028,N_7559,N_9330);
nor U10029 (N_10029,N_8376,N_8217);
nand U10030 (N_10030,N_8956,N_8501);
nand U10031 (N_10031,N_8112,N_6869);
or U10032 (N_10032,N_7434,N_8200);
nor U10033 (N_10033,N_8363,N_8172);
nand U10034 (N_10034,N_6493,N_6730);
xnor U10035 (N_10035,N_8528,N_8079);
and U10036 (N_10036,N_7426,N_6786);
and U10037 (N_10037,N_7907,N_6420);
or U10038 (N_10038,N_6919,N_6372);
nor U10039 (N_10039,N_7337,N_9218);
and U10040 (N_10040,N_8620,N_8895);
or U10041 (N_10041,N_7253,N_9159);
xor U10042 (N_10042,N_7611,N_7871);
nor U10043 (N_10043,N_8481,N_6815);
nor U10044 (N_10044,N_8396,N_6696);
xnor U10045 (N_10045,N_8385,N_6922);
and U10046 (N_10046,N_9251,N_8765);
xor U10047 (N_10047,N_8767,N_6281);
xnor U10048 (N_10048,N_6377,N_6974);
nand U10049 (N_10049,N_6418,N_9291);
and U10050 (N_10050,N_6404,N_7155);
nand U10051 (N_10051,N_7863,N_8223);
or U10052 (N_10052,N_6940,N_8898);
xor U10053 (N_10053,N_9094,N_6298);
nand U10054 (N_10054,N_9057,N_6448);
nand U10055 (N_10055,N_6463,N_7131);
and U10056 (N_10056,N_8651,N_7819);
and U10057 (N_10057,N_8490,N_8209);
nor U10058 (N_10058,N_8572,N_8101);
or U10059 (N_10059,N_8815,N_6865);
or U10060 (N_10060,N_8533,N_9260);
or U10061 (N_10061,N_6625,N_8685);
nor U10062 (N_10062,N_6421,N_8557);
nand U10063 (N_10063,N_6622,N_7767);
and U10064 (N_10064,N_6850,N_7510);
or U10065 (N_10065,N_7508,N_9363);
and U10066 (N_10066,N_9174,N_8982);
nand U10067 (N_10067,N_7164,N_6425);
and U10068 (N_10068,N_8282,N_7924);
nand U10069 (N_10069,N_6895,N_8444);
xnor U10070 (N_10070,N_6942,N_6359);
or U10071 (N_10071,N_8575,N_9026);
xor U10072 (N_10072,N_8498,N_7729);
nand U10073 (N_10073,N_7909,N_6566);
nor U10074 (N_10074,N_8100,N_8306);
nand U10075 (N_10075,N_7375,N_8386);
nand U10076 (N_10076,N_9361,N_6253);
and U10077 (N_10077,N_8564,N_7180);
and U10078 (N_10078,N_7051,N_7032);
nand U10079 (N_10079,N_7558,N_6374);
and U10080 (N_10080,N_6760,N_8837);
or U10081 (N_10081,N_7867,N_6863);
nand U10082 (N_10082,N_7872,N_6367);
xnor U10083 (N_10083,N_7987,N_7034);
or U10084 (N_10084,N_7224,N_6494);
or U10085 (N_10085,N_6835,N_7868);
or U10086 (N_10086,N_8425,N_8707);
and U10087 (N_10087,N_7624,N_7015);
nor U10088 (N_10088,N_7582,N_6699);
xor U10089 (N_10089,N_6627,N_6470);
nand U10090 (N_10090,N_8274,N_6655);
nor U10091 (N_10091,N_7591,N_9209);
or U10092 (N_10092,N_7085,N_9046);
nor U10093 (N_10093,N_6440,N_8969);
nand U10094 (N_10094,N_6556,N_6977);
and U10095 (N_10095,N_8423,N_7668);
or U10096 (N_10096,N_7000,N_8020);
xnor U10097 (N_10097,N_7318,N_6289);
nand U10098 (N_10098,N_7574,N_6853);
and U10099 (N_10099,N_7453,N_7539);
xnor U10100 (N_10100,N_9360,N_8636);
and U10101 (N_10101,N_9359,N_6551);
nor U10102 (N_10102,N_6251,N_8840);
and U10103 (N_10103,N_9084,N_9093);
nand U10104 (N_10104,N_7054,N_6643);
or U10105 (N_10105,N_8169,N_8830);
and U10106 (N_10106,N_8512,N_6611);
or U10107 (N_10107,N_6846,N_7609);
nand U10108 (N_10108,N_8488,N_9011);
and U10109 (N_10109,N_7850,N_8931);
nor U10110 (N_10110,N_6666,N_9364);
nand U10111 (N_10111,N_6605,N_7189);
xor U10112 (N_10112,N_9012,N_8772);
nand U10113 (N_10113,N_9154,N_6907);
and U10114 (N_10114,N_7003,N_8083);
and U10115 (N_10115,N_8625,N_7076);
xor U10116 (N_10116,N_6911,N_8985);
xnor U10117 (N_10117,N_6782,N_6484);
or U10118 (N_10118,N_8953,N_7422);
nand U10119 (N_10119,N_8775,N_9319);
and U10120 (N_10120,N_7291,N_6879);
nor U10121 (N_10121,N_7443,N_8394);
and U10122 (N_10122,N_6728,N_8497);
and U10123 (N_10123,N_8616,N_7903);
nand U10124 (N_10124,N_7755,N_6370);
xor U10125 (N_10125,N_7719,N_9050);
nand U10126 (N_10126,N_8496,N_6704);
nor U10127 (N_10127,N_8080,N_8216);
xor U10128 (N_10128,N_7720,N_8511);
or U10129 (N_10129,N_9337,N_8869);
or U10130 (N_10130,N_6758,N_7518);
nor U10131 (N_10131,N_6339,N_6744);
nor U10132 (N_10132,N_8719,N_8361);
xnor U10133 (N_10133,N_7593,N_8243);
nor U10134 (N_10134,N_6530,N_8224);
and U10135 (N_10135,N_6857,N_6775);
xnor U10136 (N_10136,N_9336,N_8081);
nor U10137 (N_10137,N_8197,N_8747);
nand U10138 (N_10138,N_8378,N_7017);
nor U10139 (N_10139,N_6273,N_6711);
or U10140 (N_10140,N_9024,N_7930);
or U10141 (N_10141,N_7621,N_6754);
or U10142 (N_10142,N_6294,N_6768);
nand U10143 (N_10143,N_6313,N_7835);
and U10144 (N_10144,N_7217,N_8179);
nand U10145 (N_10145,N_8720,N_8111);
xnor U10146 (N_10146,N_7330,N_8811);
and U10147 (N_10147,N_8033,N_6460);
xor U10148 (N_10148,N_7655,N_8641);
nor U10149 (N_10149,N_7832,N_7250);
nand U10150 (N_10150,N_7516,N_8995);
and U10151 (N_10151,N_7325,N_9082);
and U10152 (N_10152,N_7407,N_7926);
xor U10153 (N_10153,N_7627,N_9250);
and U10154 (N_10154,N_8731,N_8050);
or U10155 (N_10155,N_7439,N_7127);
and U10156 (N_10156,N_6396,N_6430);
xnor U10157 (N_10157,N_9186,N_7746);
nand U10158 (N_10158,N_7323,N_7317);
or U10159 (N_10159,N_8135,N_7565);
or U10160 (N_10160,N_8675,N_9002);
xnor U10161 (N_10161,N_7035,N_7401);
xor U10162 (N_10162,N_9035,N_6529);
nor U10163 (N_10163,N_6816,N_7151);
nand U10164 (N_10164,N_7420,N_6511);
and U10165 (N_10165,N_6691,N_7106);
or U10166 (N_10166,N_8932,N_7686);
and U10167 (N_10167,N_6720,N_8739);
xnor U10168 (N_10168,N_6894,N_6811);
or U10169 (N_10169,N_6921,N_9031);
xor U10170 (N_10170,N_9052,N_8996);
nor U10171 (N_10171,N_8515,N_9096);
xnor U10172 (N_10172,N_9215,N_6870);
nor U10173 (N_10173,N_8796,N_7069);
nor U10174 (N_10174,N_9148,N_6276);
nand U10175 (N_10175,N_6749,N_7975);
nor U10176 (N_10176,N_7571,N_6599);
and U10177 (N_10177,N_6752,N_7959);
nor U10178 (N_10178,N_7861,N_6303);
nand U10179 (N_10179,N_7178,N_6626);
nand U10180 (N_10180,N_7298,N_6532);
xor U10181 (N_10181,N_8546,N_6676);
xor U10182 (N_10182,N_9104,N_8186);
and U10183 (N_10183,N_8544,N_7586);
nor U10184 (N_10184,N_8491,N_6858);
nand U10185 (N_10185,N_8365,N_7260);
nor U10186 (N_10186,N_9086,N_7792);
and U10187 (N_10187,N_7561,N_7771);
nor U10188 (N_10188,N_8167,N_6883);
nor U10189 (N_10189,N_7949,N_8541);
nor U10190 (N_10190,N_8694,N_8420);
and U10191 (N_10191,N_8387,N_7379);
nor U10192 (N_10192,N_8929,N_7597);
nor U10193 (N_10193,N_6962,N_9066);
or U10194 (N_10194,N_7833,N_7387);
nor U10195 (N_10195,N_6849,N_8326);
or U10196 (N_10196,N_7968,N_8590);
and U10197 (N_10197,N_9071,N_7530);
nor U10198 (N_10198,N_7302,N_7969);
xor U10199 (N_10199,N_7812,N_8714);
nand U10200 (N_10200,N_7166,N_7885);
and U10201 (N_10201,N_6652,N_6855);
nand U10202 (N_10202,N_7111,N_7087);
nor U10203 (N_10203,N_8382,N_8114);
xnor U10204 (N_10204,N_9324,N_8640);
and U10205 (N_10205,N_8131,N_7005);
or U10206 (N_10206,N_6534,N_6504);
and U10207 (N_10207,N_8712,N_9102);
and U10208 (N_10208,N_8471,N_6886);
and U10209 (N_10209,N_9055,N_7560);
and U10210 (N_10210,N_7781,N_7740);
and U10211 (N_10211,N_6411,N_7286);
nor U10212 (N_10212,N_8930,N_9100);
nand U10213 (N_10213,N_7623,N_6936);
nor U10214 (N_10214,N_8552,N_9241);
nor U10215 (N_10215,N_6946,N_7096);
or U10216 (N_10216,N_8912,N_7238);
xor U10217 (N_10217,N_7913,N_6362);
xnor U10218 (N_10218,N_8182,N_8689);
nand U10219 (N_10219,N_9236,N_8279);
and U10220 (N_10220,N_8146,N_8587);
nand U10221 (N_10221,N_6329,N_7626);
or U10222 (N_10222,N_8886,N_6481);
nor U10223 (N_10223,N_7854,N_8210);
and U10224 (N_10224,N_7787,N_7416);
or U10225 (N_10225,N_9009,N_8705);
nand U10226 (N_10226,N_7497,N_6967);
and U10227 (N_10227,N_6827,N_6455);
nor U10228 (N_10228,N_8507,N_6689);
or U10229 (N_10229,N_7456,N_6618);
xor U10230 (N_10230,N_8679,N_7741);
nand U10231 (N_10231,N_7874,N_6764);
xnor U10232 (N_10232,N_7573,N_6956);
nand U10233 (N_10233,N_7901,N_7403);
nor U10234 (N_10234,N_6929,N_8777);
or U10235 (N_10235,N_8588,N_8923);
nor U10236 (N_10236,N_8410,N_8632);
xor U10237 (N_10237,N_8614,N_8900);
or U10238 (N_10238,N_9044,N_7588);
and U10239 (N_10239,N_9244,N_8442);
nor U10240 (N_10240,N_8031,N_7893);
nand U10241 (N_10241,N_6978,N_9294);
xor U10242 (N_10242,N_8828,N_7485);
and U10243 (N_10243,N_7728,N_8582);
or U10244 (N_10244,N_6664,N_9243);
or U10245 (N_10245,N_8583,N_6508);
nor U10246 (N_10246,N_6558,N_7637);
or U10247 (N_10247,N_8911,N_7310);
xor U10248 (N_10248,N_6291,N_7273);
and U10249 (N_10249,N_8183,N_6309);
xnor U10250 (N_10250,N_6685,N_8661);
xor U10251 (N_10251,N_8236,N_8115);
or U10252 (N_10252,N_6913,N_7769);
xnor U10253 (N_10253,N_8766,N_7158);
nor U10254 (N_10254,N_7570,N_7494);
nand U10255 (N_10255,N_6541,N_9152);
and U10256 (N_10256,N_7572,N_6763);
nor U10257 (N_10257,N_7297,N_7724);
and U10258 (N_10258,N_9008,N_7486);
nor U10259 (N_10259,N_7928,N_7390);
and U10260 (N_10260,N_8594,N_8005);
and U10261 (N_10261,N_6653,N_7821);
nand U10262 (N_10262,N_9173,N_7146);
nor U10263 (N_10263,N_8807,N_8760);
and U10264 (N_10264,N_8011,N_8344);
or U10265 (N_10265,N_7382,N_7242);
nor U10266 (N_10266,N_9321,N_7142);
xnor U10267 (N_10267,N_8741,N_8704);
nand U10268 (N_10268,N_6474,N_6959);
nand U10269 (N_10269,N_8173,N_9176);
and U10270 (N_10270,N_8853,N_8484);
or U10271 (N_10271,N_7100,N_7088);
and U10272 (N_10272,N_7147,N_7263);
nor U10273 (N_10273,N_7248,N_7568);
nor U10274 (N_10274,N_6512,N_8390);
nor U10275 (N_10275,N_6347,N_7348);
xnor U10276 (N_10276,N_9204,N_6955);
xnor U10277 (N_10277,N_7914,N_8103);
and U10278 (N_10278,N_7103,N_8623);
and U10279 (N_10279,N_8779,N_9049);
nand U10280 (N_10280,N_9220,N_7383);
nand U10281 (N_10281,N_8059,N_7124);
and U10282 (N_10282,N_6923,N_7615);
nand U10283 (N_10283,N_7483,N_8658);
nor U10284 (N_10284,N_7873,N_7764);
xnor U10285 (N_10285,N_8072,N_7025);
and U10286 (N_10286,N_6684,N_7617);
xnor U10287 (N_10287,N_6829,N_6808);
nor U10288 (N_10288,N_7759,N_8162);
xnor U10289 (N_10289,N_8844,N_8202);
nor U10290 (N_10290,N_7776,N_7240);
or U10291 (N_10291,N_7500,N_8368);
and U10292 (N_10292,N_8418,N_8025);
nand U10293 (N_10293,N_6617,N_7648);
xnor U10294 (N_10294,N_8690,N_7628);
or U10295 (N_10295,N_7231,N_8913);
nor U10296 (N_10296,N_8291,N_6714);
nor U10297 (N_10297,N_6806,N_8994);
or U10298 (N_10298,N_7044,N_7613);
and U10299 (N_10299,N_6297,N_9068);
nor U10300 (N_10300,N_7579,N_7632);
nand U10301 (N_10301,N_7498,N_8848);
and U10302 (N_10302,N_9219,N_7921);
nand U10303 (N_10303,N_9283,N_6973);
and U10304 (N_10304,N_8166,N_9025);
nor U10305 (N_10305,N_7934,N_7109);
or U10306 (N_10306,N_8684,N_8571);
nor U10307 (N_10307,N_7859,N_6402);
nor U10308 (N_10308,N_8288,N_8849);
nand U10309 (N_10309,N_9323,N_9117);
xor U10310 (N_10310,N_8855,N_8753);
nor U10311 (N_10311,N_6323,N_6657);
xor U10312 (N_10312,N_6976,N_9124);
nand U10313 (N_10313,N_9123,N_6750);
xnor U10314 (N_10314,N_8280,N_8277);
nor U10315 (N_10315,N_6710,N_7293);
and U10316 (N_10316,N_7074,N_6514);
or U10317 (N_10317,N_9145,N_6579);
nand U10318 (N_10318,N_6575,N_8275);
nor U10319 (N_10319,N_8862,N_8230);
nor U10320 (N_10320,N_8377,N_8122);
nand U10321 (N_10321,N_9253,N_7487);
xnor U10322 (N_10322,N_8827,N_9121);
nor U10323 (N_10323,N_7699,N_7335);
xnor U10324 (N_10324,N_8652,N_8251);
and U10325 (N_10325,N_6433,N_8864);
nand U10326 (N_10326,N_6671,N_9126);
or U10327 (N_10327,N_7503,N_9165);
and U10328 (N_10328,N_8762,N_8404);
nor U10329 (N_10329,N_6540,N_7944);
and U10330 (N_10330,N_6535,N_8307);
and U10331 (N_10331,N_7973,N_7817);
nand U10332 (N_10332,N_8472,N_8776);
or U10333 (N_10333,N_7212,N_8637);
nor U10334 (N_10334,N_7102,N_7018);
and U10335 (N_10335,N_7653,N_7745);
or U10336 (N_10336,N_8276,N_7513);
nor U10337 (N_10337,N_8395,N_8163);
nor U10338 (N_10338,N_8343,N_6490);
or U10339 (N_10339,N_7747,N_6743);
xor U10340 (N_10340,N_7834,N_7123);
and U10341 (N_10341,N_9246,N_7294);
xnor U10342 (N_10342,N_9083,N_6269);
xor U10343 (N_10343,N_7618,N_8628);
or U10344 (N_10344,N_7962,N_8304);
nor U10345 (N_10345,N_8356,N_8816);
nand U10346 (N_10346,N_7132,N_8293);
and U10347 (N_10347,N_7501,N_6563);
or U10348 (N_10348,N_6288,N_9302);
or U10349 (N_10349,N_8040,N_7162);
and U10350 (N_10350,N_6260,N_6731);
nand U10351 (N_10351,N_7998,N_6979);
and U10352 (N_10352,N_6299,N_9201);
nor U10353 (N_10353,N_7794,N_6567);
nand U10354 (N_10354,N_6538,N_9149);
xnor U10355 (N_10355,N_7480,N_9271);
and U10356 (N_10356,N_8194,N_8018);
or U10357 (N_10357,N_9090,N_7650);
and U10358 (N_10358,N_8346,N_8331);
or U10359 (N_10359,N_7473,N_6692);
nor U10360 (N_10360,N_7163,N_7996);
or U10361 (N_10361,N_7864,N_6642);
nand U10362 (N_10362,N_7635,N_6912);
and U10363 (N_10363,N_8219,N_6656);
or U10364 (N_10364,N_8602,N_6972);
xnor U10365 (N_10365,N_7477,N_7843);
and U10366 (N_10366,N_8526,N_9242);
nor U10367 (N_10367,N_9248,N_8022);
xnor U10368 (N_10368,N_7550,N_8283);
xor U10369 (N_10369,N_9140,N_6891);
nor U10370 (N_10370,N_8409,N_9208);
and U10371 (N_10371,N_8458,N_6545);
and U10372 (N_10372,N_6790,N_6542);
xor U10373 (N_10373,N_7662,N_6495);
or U10374 (N_10374,N_6702,N_7259);
xor U10375 (N_10375,N_6409,N_7845);
nand U10376 (N_10376,N_7837,N_8357);
xor U10377 (N_10377,N_7233,N_7952);
or U10378 (N_10378,N_9351,N_6823);
nor U10379 (N_10379,N_8773,N_6804);
or U10380 (N_10380,N_8328,N_8222);
and U10381 (N_10381,N_8648,N_8451);
nor U10382 (N_10382,N_6416,N_6686);
nand U10383 (N_10383,N_9216,N_7177);
xor U10384 (N_10384,N_7734,N_6332);
or U10385 (N_10385,N_8948,N_8754);
xnor U10386 (N_10386,N_7475,N_9015);
and U10387 (N_10387,N_8818,N_7793);
xnor U10388 (N_10388,N_6524,N_8001);
nor U10389 (N_10389,N_6439,N_6515);
xor U10390 (N_10390,N_8534,N_9301);
nor U10391 (N_10391,N_8681,N_9278);
nand U10392 (N_10392,N_9189,N_8058);
or U10393 (N_10393,N_8626,N_9268);
xor U10394 (N_10394,N_8258,N_6716);
xor U10395 (N_10395,N_8903,N_6501);
nand U10396 (N_10396,N_7904,N_6814);
nand U10397 (N_10397,N_7060,N_9116);
and U10398 (N_10398,N_7528,N_8335);
nor U10399 (N_10399,N_8810,N_8198);
or U10400 (N_10400,N_8401,N_8064);
xnor U10401 (N_10401,N_7219,N_8715);
nor U10402 (N_10402,N_7683,N_7283);
nand U10403 (N_10403,N_7353,N_6507);
or U10404 (N_10404,N_7247,N_8504);
xnor U10405 (N_10405,N_8801,N_6381);
nand U10406 (N_10406,N_8954,N_9237);
nor U10407 (N_10407,N_6633,N_8452);
and U10408 (N_10408,N_9199,N_9223);
nand U10409 (N_10409,N_6683,N_8793);
nor U10410 (N_10410,N_6861,N_7538);
or U10411 (N_10411,N_8597,N_8104);
nor U10412 (N_10412,N_8757,N_7829);
nor U10413 (N_10413,N_8427,N_6707);
nand U10414 (N_10414,N_7831,N_9039);
nand U10415 (N_10415,N_8476,N_8814);
nor U10416 (N_10416,N_7463,N_8143);
nand U10417 (N_10417,N_6447,N_7235);
xnor U10418 (N_10418,N_8189,N_8924);
nand U10419 (N_10419,N_7143,N_8273);
xnor U10420 (N_10420,N_6278,N_8302);
xor U10421 (N_10421,N_7678,N_8955);
and U10422 (N_10422,N_6985,N_8170);
and U10423 (N_10423,N_8759,N_7804);
nor U10424 (N_10424,N_8097,N_9240);
and U10425 (N_10425,N_9153,N_6949);
nor U10426 (N_10426,N_6650,N_8227);
nor U10427 (N_10427,N_7122,N_7129);
nor U10428 (N_10428,N_8524,N_8246);
xnor U10429 (N_10429,N_8519,N_6735);
nor U10430 (N_10430,N_7201,N_6703);
or U10431 (N_10431,N_7639,N_7993);
and U10432 (N_10432,N_6988,N_8936);
xor U10433 (N_10433,N_7079,N_6770);
or U10434 (N_10434,N_6701,N_7796);
and U10435 (N_10435,N_7482,N_7815);
or U10436 (N_10436,N_7992,N_9325);
nand U10437 (N_10437,N_6451,N_9279);
nor U10438 (N_10438,N_8366,N_6785);
xor U10439 (N_10439,N_9156,N_6555);
or U10440 (N_10440,N_6578,N_6975);
xor U10441 (N_10441,N_9305,N_6547);
nand U10442 (N_10442,N_6905,N_6753);
xnor U10443 (N_10443,N_8696,N_9172);
nand U10444 (N_10444,N_7552,N_8630);
nand U10445 (N_10445,N_8663,N_8428);
or U10446 (N_10446,N_8171,N_6479);
and U10447 (N_10447,N_6523,N_7960);
xor U10448 (N_10448,N_7645,N_7657);
or U10449 (N_10449,N_8310,N_8446);
xnor U10450 (N_10450,N_8771,N_7929);
xnor U10451 (N_10451,N_8792,N_9368);
nand U10452 (N_10452,N_7270,N_8744);
nand U10453 (N_10453,N_8347,N_7472);
and U10454 (N_10454,N_8794,N_7646);
nor U10455 (N_10455,N_6595,N_8980);
or U10456 (N_10456,N_7425,N_8017);
or U10457 (N_10457,N_7997,N_8709);
or U10458 (N_10458,N_7040,N_9111);
nand U10459 (N_10459,N_6257,N_6328);
or U10460 (N_10460,N_9048,N_9259);
and U10461 (N_10461,N_6497,N_9373);
and U10462 (N_10462,N_8165,N_8300);
nand U10463 (N_10463,N_9063,N_6365);
or U10464 (N_10464,N_6612,N_7020);
nand U10465 (N_10465,N_6600,N_6401);
xor U10466 (N_10466,N_8225,N_6354);
nand U10467 (N_10467,N_7982,N_6569);
nor U10468 (N_10468,N_8554,N_7355);
xor U10469 (N_10469,N_8082,N_7075);
and U10470 (N_10470,N_6487,N_7414);
nor U10471 (N_10471,N_8826,N_9193);
xnor U10472 (N_10472,N_7429,N_7990);
and U10473 (N_10473,N_6537,N_6587);
nand U10474 (N_10474,N_7564,N_9327);
and U10475 (N_10475,N_6331,N_6327);
nor U10476 (N_10476,N_8664,N_8150);
nor U10477 (N_10477,N_8540,N_9131);
nor U10478 (N_10478,N_7448,N_9284);
nand U10479 (N_10479,N_7381,N_9169);
or U10480 (N_10480,N_8492,N_8132);
nand U10481 (N_10481,N_8971,N_8601);
and U10482 (N_10482,N_9040,N_8003);
nand U10483 (N_10483,N_6283,N_8406);
nand U10484 (N_10484,N_8400,N_7970);
and U10485 (N_10485,N_8915,N_8671);
nand U10486 (N_10486,N_8015,N_9207);
nand U10487 (N_10487,N_9285,N_7341);
xor U10488 (N_10488,N_6356,N_9202);
or U10489 (N_10489,N_7399,N_6839);
nand U10490 (N_10490,N_7165,N_8606);
or U10491 (N_10491,N_8786,N_7705);
or U10492 (N_10492,N_7450,N_8184);
or U10493 (N_10493,N_6506,N_8593);
and U10494 (N_10494,N_8857,N_6408);
nand U10495 (N_10495,N_6412,N_6847);
nor U10496 (N_10496,N_9217,N_6266);
nor U10497 (N_10497,N_7824,N_7592);
xnor U10498 (N_10498,N_8737,N_8049);
nand U10499 (N_10499,N_8199,N_7562);
nand U10500 (N_10500,N_7468,N_7707);
xnor U10501 (N_10501,N_6960,N_7957);
and U10502 (N_10502,N_8919,N_9347);
xor U10503 (N_10503,N_6414,N_7880);
or U10504 (N_10504,N_6489,N_8467);
or U10505 (N_10505,N_9230,N_7533);
nor U10506 (N_10506,N_8998,N_6265);
nand U10507 (N_10507,N_8656,N_6825);
nand U10508 (N_10508,N_9013,N_6306);
nand U10509 (N_10509,N_8397,N_7797);
xnor U10510 (N_10510,N_7104,N_7205);
or U10511 (N_10511,N_6312,N_7415);
nor U10512 (N_10512,N_6355,N_6413);
xnor U10513 (N_10513,N_8698,N_7006);
nor U10514 (N_10514,N_7629,N_7269);
and U10515 (N_10515,N_8831,N_6629);
xor U10516 (N_10516,N_7601,N_9062);
xor U10517 (N_10517,N_6969,N_7352);
xor U10518 (N_10518,N_8860,N_8151);
nand U10519 (N_10519,N_6311,N_6581);
nor U10520 (N_10520,N_8359,N_8863);
xor U10521 (N_10521,N_8175,N_6843);
xnor U10522 (N_10522,N_8153,N_6435);
nor U10523 (N_10523,N_9316,N_8249);
and U10524 (N_10524,N_7393,N_8424);
nand U10525 (N_10525,N_6737,N_7576);
nor U10526 (N_10526,N_8735,N_8421);
and U10527 (N_10527,N_7159,N_8787);
or U10528 (N_10528,N_8599,N_6369);
nand U10529 (N_10529,N_7536,N_6615);
nor U10530 (N_10530,N_7411,N_6293);
xor U10531 (N_10531,N_7995,N_9340);
or U10532 (N_10532,N_8261,N_8901);
nand U10533 (N_10533,N_6648,N_6755);
or U10534 (N_10534,N_6371,N_6280);
nor U10535 (N_10535,N_7737,N_7309);
or U10536 (N_10536,N_8317,N_9276);
nand U10537 (N_10537,N_8505,N_6875);
nand U10538 (N_10538,N_8041,N_8301);
xor U10539 (N_10539,N_7961,N_8393);
nor U10540 (N_10540,N_6560,N_7842);
nand U10541 (N_10541,N_8076,N_7410);
or U10542 (N_10542,N_7038,N_6385);
xor U10543 (N_10543,N_9106,N_8876);
xnor U10544 (N_10544,N_6645,N_6887);
or U10545 (N_10545,N_9203,N_8791);
nor U10546 (N_10546,N_8139,N_6352);
and U10547 (N_10547,N_8089,N_8267);
or U10548 (N_10548,N_7488,N_8245);
nand U10549 (N_10549,N_7214,N_9045);
xnor U10550 (N_10550,N_7688,N_7313);
xnor U10551 (N_10551,N_7457,N_6971);
or U10552 (N_10552,N_9233,N_6492);
xnor U10553 (N_10553,N_8957,N_7865);
and U10554 (N_10554,N_7061,N_7784);
and U10555 (N_10555,N_7986,N_9139);
nand U10556 (N_10556,N_8691,N_9058);
or U10557 (N_10557,N_9065,N_8155);
xor U10558 (N_10558,N_7133,N_8047);
and U10559 (N_10559,N_9304,N_6673);
nand U10560 (N_10560,N_7261,N_7185);
and U10561 (N_10561,N_9043,N_6980);
and U10562 (N_10562,N_8939,N_6862);
xor U10563 (N_10563,N_7014,N_8264);
and U10564 (N_10564,N_6528,N_6255);
and U10565 (N_10565,N_8560,N_9228);
or U10566 (N_10566,N_9342,N_6920);
nand U10567 (N_10567,N_7207,N_7343);
xor U10568 (N_10568,N_7811,N_8635);
and U10569 (N_10569,N_8134,N_6619);
xnor U10570 (N_10570,N_7278,N_6893);
xor U10571 (N_10571,N_8176,N_6341);
nor U10572 (N_10572,N_6939,N_8700);
nor U10573 (N_10573,N_7479,N_7206);
xnor U10574 (N_10574,N_6317,N_8426);
nor U10575 (N_10575,N_7826,N_7303);
or U10576 (N_10576,N_7827,N_6380);
nand U10577 (N_10577,N_8774,N_9180);
and U10578 (N_10578,N_6516,N_7467);
and U10579 (N_10579,N_9081,N_9338);
and U10580 (N_10580,N_6584,N_7179);
or U10581 (N_10581,N_7262,N_6736);
and U10582 (N_10582,N_9225,N_7953);
and U10583 (N_10583,N_8154,N_6539);
xnor U10584 (N_10584,N_9266,N_7126);
nand U10585 (N_10585,N_8062,N_8070);
nand U10586 (N_10586,N_9091,N_6320);
or U10587 (N_10587,N_7608,N_8952);
nor U10588 (N_10588,N_8164,N_9166);
nor U10589 (N_10589,N_6315,N_8940);
xor U10590 (N_10590,N_8865,N_7607);
or U10591 (N_10591,N_9348,N_7064);
and U10592 (N_10592,N_6350,N_6813);
and U10593 (N_10593,N_7328,N_9317);
nor U10594 (N_10594,N_7853,N_7226);
xor U10595 (N_10595,N_8373,N_6871);
xnor U10596 (N_10596,N_8610,N_8510);
and U10597 (N_10597,N_8746,N_8595);
xnor U10598 (N_10598,N_6357,N_6995);
or U10599 (N_10599,N_9270,N_7933);
xnor U10600 (N_10600,N_8732,N_7354);
nor U10601 (N_10601,N_7101,N_7847);
nand U10602 (N_10602,N_8618,N_6636);
nor U10603 (N_10603,N_8586,N_7587);
and U10604 (N_10604,N_7125,N_8667);
nor U10605 (N_10605,N_6958,N_7319);
xor U10606 (N_10606,N_9310,N_6632);
and U10607 (N_10607,N_6803,N_9163);
nor U10608 (N_10608,N_7806,N_9158);
nand U10609 (N_10609,N_6500,N_7090);
xor U10610 (N_10610,N_8591,N_7351);
xnor U10611 (N_10611,N_7299,N_8042);
nor U10612 (N_10612,N_7447,N_7779);
and U10613 (N_10613,N_8339,N_6747);
and U10614 (N_10614,N_7377,N_6482);
xor U10615 (N_10615,N_7266,N_6884);
or U10616 (N_10616,N_8742,N_7110);
nand U10617 (N_10617,N_7397,N_9227);
or U10618 (N_10618,N_7168,N_7187);
and U10619 (N_10619,N_8859,N_7171);
nor U10620 (N_10620,N_9333,N_6325);
nand U10621 (N_10621,N_7222,N_7312);
nand U10622 (N_10622,N_6483,N_8453);
nor U10623 (N_10623,N_8879,N_8989);
nor U10624 (N_10624,N_6738,N_9374);
xnor U10625 (N_10625,N_9210,N_6990);
or U10626 (N_10626,N_8861,N_6950);
nand U10627 (N_10627,N_7360,N_7744);
nand U10628 (N_10628,N_8138,N_6672);
and U10629 (N_10629,N_7855,N_8893);
nor U10630 (N_10630,N_8468,N_8118);
nand U10631 (N_10631,N_7173,N_9168);
and U10632 (N_10632,N_6513,N_8422);
and U10633 (N_10633,N_8350,N_6935);
xnor U10634 (N_10634,N_8384,N_8907);
nand U10635 (N_10635,N_6394,N_8477);
nand U10636 (N_10636,N_8854,N_7474);
and U10637 (N_10637,N_8885,N_8972);
nand U10638 (N_10638,N_7948,N_9128);
nor U10639 (N_10639,N_6469,N_8093);
or U10640 (N_10640,N_7851,N_8697);
and U10641 (N_10641,N_7878,N_8517);
nor U10642 (N_10642,N_9017,N_9200);
and U10643 (N_10643,N_7141,N_8803);
nand U10644 (N_10644,N_7001,N_8487);
or U10645 (N_10645,N_7423,N_6279);
nor U10646 (N_10646,N_9287,N_6836);
and U10647 (N_10647,N_8874,N_9313);
or U10648 (N_10648,N_7887,N_6638);
nand U10649 (N_10649,N_7856,N_6274);
and U10650 (N_10650,N_8992,N_7430);
or U10651 (N_10651,N_8174,N_7912);
xor U10652 (N_10652,N_7656,N_6346);
xor U10653 (N_10653,N_7991,N_8832);
xnor U10654 (N_10654,N_6924,N_8609);
nand U10655 (N_10655,N_8638,N_8221);
nor U10656 (N_10656,N_9170,N_8740);
and U10657 (N_10657,N_9213,N_7751);
nand U10658 (N_10658,N_7584,N_8060);
nand U10659 (N_10659,N_7004,N_6467);
nor U10660 (N_10660,N_9226,N_8882);
xnor U10661 (N_10661,N_7373,N_7937);
or U10662 (N_10662,N_8044,N_7906);
nand U10663 (N_10663,N_8237,N_7371);
xor U10664 (N_10664,N_8185,N_9332);
xnor U10665 (N_10665,N_6658,N_6422);
nor U10666 (N_10666,N_8284,N_8823);
nand U10667 (N_10667,N_6382,N_9030);
or U10668 (N_10668,N_7441,N_8928);
and U10669 (N_10669,N_8364,N_9277);
nor U10670 (N_10670,N_9273,N_8961);
xor U10671 (N_10671,N_9134,N_8934);
or U10672 (N_10672,N_7669,N_8905);
nor U10673 (N_10673,N_8037,N_8536);
and U10674 (N_10674,N_6596,N_7772);
and U10675 (N_10675,N_7600,N_7290);
nor U10676 (N_10676,N_6987,N_6759);
xnor U10677 (N_10677,N_7891,N_8659);
and U10678 (N_10678,N_9059,N_7349);
or U10679 (N_10679,N_9164,N_6963);
nand U10680 (N_10680,N_8228,N_7324);
and U10681 (N_10681,N_8553,N_8629);
nor U10682 (N_10682,N_8415,N_7308);
nand U10683 (N_10683,N_6606,N_6549);
nand U10684 (N_10684,N_7649,N_7902);
and U10685 (N_10685,N_7462,N_8008);
nand U10686 (N_10686,N_6384,N_7216);
or U10687 (N_10687,N_8124,N_8983);
nand U10688 (N_10688,N_9356,N_6300);
nand U10689 (N_10689,N_7766,N_8734);
nor U10690 (N_10690,N_9141,N_8710);
nor U10691 (N_10691,N_7339,N_8004);
nor U10692 (N_10692,N_9150,N_7549);
nand U10693 (N_10693,N_8416,N_8717);
nor U10694 (N_10694,N_6272,N_8749);
nand U10695 (N_10695,N_8763,N_7703);
nor U10696 (N_10696,N_9155,N_7010);
xor U10697 (N_10697,N_7712,N_8454);
and U10698 (N_10698,N_8242,N_7098);
nor U10699 (N_10699,N_7030,N_7007);
or U10700 (N_10700,N_6948,N_8547);
xor U10701 (N_10701,N_8970,N_7022);
nor U10702 (N_10702,N_6717,N_8518);
xnor U10703 (N_10703,N_8354,N_6441);
nand U10704 (N_10704,N_8340,N_7634);
nor U10705 (N_10705,N_8144,N_7268);
or U10706 (N_10706,N_6486,N_7059);
nand U10707 (N_10707,N_6337,N_9306);
xnor U10708 (N_10708,N_7919,N_9080);
xnor U10709 (N_10709,N_9110,N_7215);
nor U10710 (N_10710,N_8880,N_9051);
nor U10711 (N_10711,N_6828,N_6604);
nand U10712 (N_10712,N_7706,N_7756);
nand U10713 (N_10713,N_8906,N_9016);
nand U10714 (N_10714,N_8805,N_7091);
nor U10715 (N_10715,N_8548,N_7916);
and U10716 (N_10716,N_7723,N_7058);
or U10717 (N_10717,N_6613,N_7927);
xor U10718 (N_10718,N_7750,N_6767);
or U10719 (N_10719,N_7922,N_6399);
or U10720 (N_10720,N_7553,N_7436);
and U10721 (N_10721,N_7698,N_7176);
or U10722 (N_10722,N_6677,N_7394);
nor U10723 (N_10723,N_8212,N_6572);
xnor U10724 (N_10724,N_7672,N_8098);
and U10725 (N_10725,N_6903,N_7369);
nand U10726 (N_10726,N_8493,N_8738);
nand U10727 (N_10727,N_8871,N_8073);
nand U10728 (N_10728,N_8711,N_8845);
nor U10729 (N_10729,N_6665,N_8311);
nand U10730 (N_10730,N_8963,N_8084);
xor U10731 (N_10731,N_7431,N_6333);
nand U10732 (N_10732,N_8733,N_7281);
or U10733 (N_10733,N_7172,N_8358);
or U10734 (N_10734,N_7356,N_6756);
xnor U10735 (N_10735,N_7336,N_8611);
or U10736 (N_10736,N_7545,N_6712);
xnor U10737 (N_10737,N_6680,N_9353);
xnor U10738 (N_10738,N_6410,N_8824);
nor U10739 (N_10739,N_8457,N_8485);
and U10740 (N_10740,N_7068,N_7665);
nor U10741 (N_10741,N_9281,N_7301);
or U10742 (N_10742,N_6562,N_7985);
or U10743 (N_10743,N_6603,N_8916);
nor U10744 (N_10744,N_7246,N_8021);
and U10745 (N_10745,N_8960,N_8894);
xnor U10746 (N_10746,N_8702,N_8639);
and U10747 (N_10747,N_8843,N_7322);
and U10748 (N_10748,N_9331,N_7890);
xor U10749 (N_10749,N_7417,N_8833);
nor U10750 (N_10750,N_6446,N_6917);
and U10751 (N_10751,N_9122,N_9212);
nor U10752 (N_10752,N_9079,N_8977);
xnor U10753 (N_10753,N_6669,N_9061);
xnor U10754 (N_10754,N_6458,N_7499);
and U10755 (N_10755,N_6351,N_6933);
xnor U10756 (N_10756,N_7773,N_7825);
xor U10757 (N_10757,N_6557,N_7696);
nor U10758 (N_10758,N_7585,N_8161);
nand U10759 (N_10759,N_6436,N_7569);
xnor U10760 (N_10760,N_7272,N_7378);
nor U10761 (N_10761,N_7116,N_8268);
nor U10762 (N_10762,N_8250,N_6314);
nor U10763 (N_10763,N_9299,N_6330);
xor U10764 (N_10764,N_6546,N_8372);
and U10765 (N_10765,N_6761,N_8677);
or U10766 (N_10766,N_8438,N_7830);
nand U10767 (N_10767,N_9293,N_7941);
nor U10768 (N_10768,N_9196,N_8627);
xnor U10769 (N_10769,N_6434,N_8255);
nand U10770 (N_10770,N_8253,N_7509);
or U10771 (N_10771,N_6438,N_7481);
and U10772 (N_10772,N_8233,N_8592);
nor U10773 (N_10773,N_9367,N_7866);
xor U10774 (N_10774,N_7021,N_8573);
nor U10775 (N_10775,N_7641,N_8621);
nand U10776 (N_10776,N_8921,N_7710);
or U10777 (N_10777,N_7542,N_8019);
xnor U10778 (N_10778,N_7567,N_6842);
xnor U10779 (N_10779,N_9184,N_7736);
or U10780 (N_10780,N_7203,N_6640);
or U10781 (N_10781,N_6856,N_9350);
and U10782 (N_10782,N_8941,N_9234);
nor U10783 (N_10783,N_7900,N_8325);
and U10784 (N_10784,N_7209,N_8075);
or U10785 (N_10785,N_7184,N_7511);
xnor U10786 (N_10786,N_9114,N_6740);
xor U10787 (N_10787,N_8333,N_8822);
nand U10788 (N_10788,N_6984,N_9288);
and U10789 (N_10789,N_6661,N_9113);
xor U10790 (N_10790,N_6709,N_6275);
nor U10791 (N_10791,N_6527,N_8500);
nand U10792 (N_10792,N_7279,N_7983);
xnor U10793 (N_10793,N_7384,N_8799);
and U10794 (N_10794,N_8764,N_7881);
nor U10795 (N_10795,N_7979,N_8035);
and U10796 (N_10796,N_7342,N_8633);
nand U10797 (N_10797,N_7661,N_8193);
xor U10798 (N_10798,N_6342,N_6945);
xor U10799 (N_10799,N_8881,N_8802);
xnor U10800 (N_10800,N_7469,N_7721);
nand U10801 (N_10801,N_8653,N_7197);
or U10802 (N_10802,N_7852,N_9099);
and U10803 (N_10803,N_7249,N_6789);
nand U10804 (N_10804,N_7557,N_6407);
nand U10805 (N_10805,N_8129,N_8032);
xor U10806 (N_10806,N_9365,N_7619);
nor U10807 (N_10807,N_7700,N_8670);
nor U10808 (N_10808,N_8207,N_7938);
nor U10809 (N_10809,N_6466,N_8123);
and U10810 (N_10810,N_8312,N_7419);
or U10811 (N_10811,N_7966,N_7043);
or U10812 (N_10812,N_6478,N_6961);
nand U10813 (N_10813,N_8569,N_8549);
xnor U10814 (N_10814,N_6577,N_9339);
xor U10815 (N_10815,N_9269,N_7115);
or U10816 (N_10816,N_7053,N_6552);
and U10817 (N_10817,N_8808,N_8979);
nand U10818 (N_10818,N_8647,N_8090);
nor U10819 (N_10819,N_9303,N_9322);
or U10820 (N_10820,N_7692,N_7418);
nand U10821 (N_10821,N_8380,N_6583);
xnor U10822 (N_10822,N_7372,N_6308);
or U10823 (N_10823,N_6282,N_6732);
and U10824 (N_10824,N_6592,N_7139);
xnor U10825 (N_10825,N_8119,N_6641);
nand U10826 (N_10826,N_6687,N_7150);
and U10827 (N_10827,N_7849,N_8756);
nand U10828 (N_10828,N_6533,N_6431);
or U10829 (N_10829,N_8556,N_6334);
nand U10830 (N_10830,N_6784,N_6634);
and U10831 (N_10831,N_6964,N_6951);
and U10832 (N_10832,N_7651,N_7753);
xnor U10833 (N_10833,N_7936,N_8052);
xor U10834 (N_10834,N_8695,N_6794);
and U10835 (N_10835,N_8218,N_7935);
nor U10836 (N_10836,N_7066,N_6918);
nand U10837 (N_10837,N_8574,N_7923);
or U10838 (N_10838,N_7524,N_8535);
nand U10839 (N_10839,N_8701,N_9085);
nor U10840 (N_10840,N_7364,N_8486);
and U10841 (N_10841,N_8229,N_8868);
nand U10842 (N_10842,N_6663,N_6588);
or U10843 (N_10843,N_9142,N_8077);
and U10844 (N_10844,N_6503,N_6721);
xor U10845 (N_10845,N_8321,N_6395);
and U10846 (N_10846,N_9018,N_7031);
nor U10847 (N_10847,N_6867,N_8078);
nor U10848 (N_10848,N_8338,N_8678);
and U10849 (N_10849,N_6890,N_8499);
or U10850 (N_10850,N_7365,N_8431);
and U10851 (N_10851,N_6776,N_8645);
and U10852 (N_10852,N_7654,N_9010);
xor U10853 (N_10853,N_8615,N_6762);
and U10854 (N_10854,N_6668,N_8308);
nor U10855 (N_10855,N_8790,N_6742);
xor U10856 (N_10856,N_7464,N_8045);
xor U10857 (N_10857,N_7223,N_8204);
nor U10858 (N_10858,N_7778,N_6623);
nand U10859 (N_10859,N_7670,N_6295);
nor U10860 (N_10860,N_6797,N_8918);
xor U10861 (N_10861,N_8604,N_7138);
and U10862 (N_10862,N_7029,N_7016);
and U10863 (N_10863,N_8337,N_7523);
or U10864 (N_10864,N_9005,N_7964);
nor U10865 (N_10865,N_9089,N_9161);
or U10866 (N_10866,N_8388,N_8987);
nor U10867 (N_10867,N_9366,N_7512);
xnor U10868 (N_10868,N_7892,N_9257);
or U10869 (N_10869,N_8585,N_8706);
nand U10870 (N_10870,N_6398,N_6899);
or U10871 (N_10871,N_7614,N_6690);
nand U10872 (N_10872,N_9092,N_8061);
nor U10873 (N_10873,N_8935,N_7225);
and U10874 (N_10874,N_6880,N_6338);
nand U10875 (N_10875,N_8804,N_8271);
nand U10876 (N_10876,N_6695,N_8888);
and U10877 (N_10877,N_6345,N_7047);
nand U10878 (N_10878,N_8820,N_9282);
xnor U10879 (N_10879,N_6536,N_6909);
and U10880 (N_10880,N_6259,N_8835);
nand U10881 (N_10881,N_7154,N_8847);
xnor U10882 (N_10882,N_7340,N_7065);
xor U10883 (N_10883,N_7733,N_7192);
xor U10884 (N_10884,N_6930,N_8352);
and U10885 (N_10885,N_6387,N_9027);
nand U10886 (N_10886,N_7367,N_6348);
nor U10887 (N_10887,N_6781,N_8023);
nand U10888 (N_10888,N_6791,N_8028);
xnor U10889 (N_10889,N_6966,N_8502);
xnor U10890 (N_10890,N_6965,N_8806);
nor U10891 (N_10891,N_8137,N_9371);
nand U10892 (N_10892,N_8294,N_8362);
nand U10893 (N_10893,N_7502,N_9115);
and U10894 (N_10894,N_6324,N_8205);
or U10895 (N_10895,N_9033,N_7828);
nor U10896 (N_10896,N_7788,N_7726);
nor U10897 (N_10897,N_7458,N_9341);
and U10898 (N_10898,N_8211,N_9162);
and U10899 (N_10899,N_9182,N_7296);
and U10900 (N_10900,N_8964,N_8565);
nand U10901 (N_10901,N_9290,N_7682);
xor U10902 (N_10902,N_6647,N_7940);
xor U10903 (N_10903,N_8666,N_8469);
nor U10904 (N_10904,N_6682,N_6602);
nand U10905 (N_10905,N_6872,N_7108);
and U10906 (N_10906,N_8455,N_9370);
nand U10907 (N_10907,N_6443,N_7391);
nand U10908 (N_10908,N_7727,N_6485);
or U10909 (N_10909,N_7978,N_7338);
nor U10910 (N_10910,N_9077,N_9349);
or U10911 (N_10911,N_7077,N_7799);
xnor U10912 (N_10912,N_8436,N_7476);
or U10913 (N_10913,N_9056,N_9129);
nand U10914 (N_10914,N_6531,N_6954);
or U10915 (N_10915,N_8030,N_8494);
nor U10916 (N_10916,N_6284,N_8196);
and U10917 (N_10917,N_7042,N_8262);
xnor U10918 (N_10918,N_6620,N_8722);
nand U10919 (N_10919,N_7316,N_6998);
xnor U10920 (N_10920,N_8391,N_6475);
xnor U10921 (N_10921,N_9232,N_9195);
xnor U10922 (N_10922,N_8660,N_9263);
xor U10923 (N_10923,N_7037,N_8286);
nand U10924 (N_10924,N_6597,N_6452);
and U10925 (N_10925,N_7028,N_7285);
and U10926 (N_10926,N_9309,N_6258);
and U10927 (N_10927,N_7870,N_7496);
xnor U10928 (N_10928,N_8513,N_6631);
nor U10929 (N_10929,N_8158,N_7714);
nor U10930 (N_10930,N_6957,N_8568);
or U10931 (N_10931,N_8674,N_9312);
nand U10932 (N_10932,N_6688,N_7888);
nand U10933 (N_10933,N_9151,N_8724);
or U10934 (N_10934,N_7204,N_7899);
xor U10935 (N_10935,N_7039,N_8748);
nor U10936 (N_10936,N_8375,N_8768);
nand U10937 (N_10937,N_7359,N_7767);
or U10938 (N_10938,N_9073,N_7930);
or U10939 (N_10939,N_9172,N_9326);
xor U10940 (N_10940,N_9247,N_6714);
nor U10941 (N_10941,N_8148,N_7442);
nand U10942 (N_10942,N_8950,N_9122);
or U10943 (N_10943,N_7982,N_6995);
nor U10944 (N_10944,N_8130,N_7272);
nor U10945 (N_10945,N_6966,N_7453);
and U10946 (N_10946,N_8784,N_7539);
nand U10947 (N_10947,N_7783,N_6342);
xnor U10948 (N_10948,N_9158,N_7621);
or U10949 (N_10949,N_6317,N_6953);
xnor U10950 (N_10950,N_9242,N_8971);
and U10951 (N_10951,N_7092,N_7054);
nand U10952 (N_10952,N_9099,N_8296);
or U10953 (N_10953,N_8972,N_8981);
or U10954 (N_10954,N_7864,N_7891);
xnor U10955 (N_10955,N_7318,N_8618);
nor U10956 (N_10956,N_9236,N_6495);
nor U10957 (N_10957,N_8477,N_7427);
and U10958 (N_10958,N_7176,N_6535);
xnor U10959 (N_10959,N_6774,N_7025);
nand U10960 (N_10960,N_7803,N_7548);
or U10961 (N_10961,N_8228,N_7894);
or U10962 (N_10962,N_8089,N_7011);
xor U10963 (N_10963,N_9370,N_6618);
or U10964 (N_10964,N_6919,N_8877);
nor U10965 (N_10965,N_7546,N_6625);
and U10966 (N_10966,N_8401,N_6563);
xor U10967 (N_10967,N_8821,N_8692);
nand U10968 (N_10968,N_7839,N_6741);
and U10969 (N_10969,N_8129,N_8349);
or U10970 (N_10970,N_6505,N_9150);
xor U10971 (N_10971,N_6967,N_8211);
nand U10972 (N_10972,N_6820,N_6361);
and U10973 (N_10973,N_8803,N_6804);
xnor U10974 (N_10974,N_7158,N_6748);
or U10975 (N_10975,N_6438,N_7793);
nor U10976 (N_10976,N_7243,N_9214);
and U10977 (N_10977,N_8317,N_7523);
nor U10978 (N_10978,N_8583,N_8664);
or U10979 (N_10979,N_6539,N_7562);
xnor U10980 (N_10980,N_8975,N_7560);
or U10981 (N_10981,N_8751,N_7894);
nor U10982 (N_10982,N_6463,N_7168);
nand U10983 (N_10983,N_8394,N_6508);
nand U10984 (N_10984,N_8066,N_7105);
nand U10985 (N_10985,N_8565,N_8155);
or U10986 (N_10986,N_8257,N_8676);
nor U10987 (N_10987,N_9356,N_9051);
nand U10988 (N_10988,N_9235,N_7595);
xnor U10989 (N_10989,N_8349,N_7707);
nand U10990 (N_10990,N_9137,N_6377);
nor U10991 (N_10991,N_9277,N_7235);
nand U10992 (N_10992,N_7473,N_6719);
xor U10993 (N_10993,N_6930,N_9041);
nor U10994 (N_10994,N_7151,N_8882);
nor U10995 (N_10995,N_7956,N_6673);
or U10996 (N_10996,N_9176,N_7826);
xor U10997 (N_10997,N_6393,N_8262);
or U10998 (N_10998,N_7411,N_6273);
and U10999 (N_10999,N_6923,N_7497);
and U11000 (N_11000,N_9007,N_7970);
nor U11001 (N_11001,N_8385,N_8208);
xor U11002 (N_11002,N_6525,N_7493);
nand U11003 (N_11003,N_8572,N_6323);
or U11004 (N_11004,N_8216,N_7097);
or U11005 (N_11005,N_6302,N_6640);
nor U11006 (N_11006,N_7692,N_7395);
nand U11007 (N_11007,N_7734,N_8333);
nand U11008 (N_11008,N_9347,N_8971);
nor U11009 (N_11009,N_8049,N_6735);
and U11010 (N_11010,N_6360,N_6642);
nand U11011 (N_11011,N_7308,N_6555);
nand U11012 (N_11012,N_6815,N_6313);
xnor U11013 (N_11013,N_7131,N_7721);
nor U11014 (N_11014,N_8571,N_9329);
and U11015 (N_11015,N_8850,N_8270);
and U11016 (N_11016,N_8777,N_6803);
nor U11017 (N_11017,N_6373,N_7313);
nand U11018 (N_11018,N_8079,N_7307);
nor U11019 (N_11019,N_6928,N_6741);
and U11020 (N_11020,N_8890,N_7459);
or U11021 (N_11021,N_7242,N_8363);
or U11022 (N_11022,N_9141,N_6981);
and U11023 (N_11023,N_7565,N_6608);
xor U11024 (N_11024,N_7275,N_8049);
xor U11025 (N_11025,N_8520,N_8361);
and U11026 (N_11026,N_7328,N_8914);
or U11027 (N_11027,N_7341,N_7474);
and U11028 (N_11028,N_7562,N_8436);
xor U11029 (N_11029,N_7209,N_8023);
nor U11030 (N_11030,N_7578,N_8037);
nand U11031 (N_11031,N_8068,N_9267);
or U11032 (N_11032,N_8697,N_9136);
or U11033 (N_11033,N_8055,N_8527);
xnor U11034 (N_11034,N_9088,N_7013);
nor U11035 (N_11035,N_8057,N_7728);
and U11036 (N_11036,N_6451,N_7804);
and U11037 (N_11037,N_8105,N_8927);
nand U11038 (N_11038,N_7390,N_7784);
or U11039 (N_11039,N_8649,N_6633);
nor U11040 (N_11040,N_6486,N_8989);
xnor U11041 (N_11041,N_7731,N_7997);
or U11042 (N_11042,N_8643,N_7688);
or U11043 (N_11043,N_6807,N_7837);
or U11044 (N_11044,N_9125,N_6355);
nor U11045 (N_11045,N_7104,N_7605);
nor U11046 (N_11046,N_9043,N_8821);
nand U11047 (N_11047,N_7688,N_8144);
and U11048 (N_11048,N_7074,N_7279);
or U11049 (N_11049,N_6638,N_8568);
or U11050 (N_11050,N_9106,N_9138);
nand U11051 (N_11051,N_8048,N_6399);
or U11052 (N_11052,N_8040,N_6990);
or U11053 (N_11053,N_8452,N_8269);
nor U11054 (N_11054,N_8997,N_8390);
nor U11055 (N_11055,N_7933,N_7517);
and U11056 (N_11056,N_7031,N_9147);
nor U11057 (N_11057,N_7573,N_6885);
nor U11058 (N_11058,N_6317,N_8769);
xor U11059 (N_11059,N_7195,N_8186);
xor U11060 (N_11060,N_8125,N_8897);
xnor U11061 (N_11061,N_6591,N_7392);
xnor U11062 (N_11062,N_8603,N_6965);
nand U11063 (N_11063,N_7120,N_8502);
and U11064 (N_11064,N_6483,N_8029);
or U11065 (N_11065,N_9240,N_8713);
and U11066 (N_11066,N_7005,N_7408);
xnor U11067 (N_11067,N_8346,N_9146);
nor U11068 (N_11068,N_7640,N_8861);
nand U11069 (N_11069,N_6736,N_7407);
nand U11070 (N_11070,N_7193,N_7095);
or U11071 (N_11071,N_9011,N_7278);
or U11072 (N_11072,N_6473,N_9150);
and U11073 (N_11073,N_8551,N_8165);
nor U11074 (N_11074,N_7819,N_6803);
or U11075 (N_11075,N_7695,N_8300);
nand U11076 (N_11076,N_8686,N_8353);
and U11077 (N_11077,N_6554,N_6810);
and U11078 (N_11078,N_7594,N_7629);
nand U11079 (N_11079,N_8412,N_6889);
and U11080 (N_11080,N_6894,N_8403);
nor U11081 (N_11081,N_8940,N_9231);
and U11082 (N_11082,N_8739,N_8266);
nand U11083 (N_11083,N_6944,N_8531);
nor U11084 (N_11084,N_6350,N_7610);
nand U11085 (N_11085,N_7895,N_8396);
and U11086 (N_11086,N_8247,N_7394);
or U11087 (N_11087,N_7497,N_6785);
and U11088 (N_11088,N_8471,N_8745);
or U11089 (N_11089,N_8666,N_8503);
nor U11090 (N_11090,N_8317,N_7063);
xnor U11091 (N_11091,N_8269,N_8878);
nor U11092 (N_11092,N_8252,N_7512);
nor U11093 (N_11093,N_7369,N_6720);
or U11094 (N_11094,N_7971,N_6779);
or U11095 (N_11095,N_8736,N_8288);
or U11096 (N_11096,N_9247,N_9021);
xor U11097 (N_11097,N_6676,N_8726);
nor U11098 (N_11098,N_7691,N_7035);
nor U11099 (N_11099,N_6484,N_8965);
and U11100 (N_11100,N_7173,N_6691);
xnor U11101 (N_11101,N_8026,N_7667);
and U11102 (N_11102,N_8802,N_7017);
nor U11103 (N_11103,N_9147,N_6366);
nor U11104 (N_11104,N_6864,N_6819);
nor U11105 (N_11105,N_7152,N_6643);
nor U11106 (N_11106,N_6714,N_7810);
xnor U11107 (N_11107,N_7617,N_9166);
or U11108 (N_11108,N_8633,N_8637);
or U11109 (N_11109,N_8104,N_8166);
nor U11110 (N_11110,N_8780,N_7751);
and U11111 (N_11111,N_6916,N_9079);
nor U11112 (N_11112,N_7153,N_6498);
nand U11113 (N_11113,N_6666,N_7471);
or U11114 (N_11114,N_8534,N_8255);
nand U11115 (N_11115,N_6871,N_7961);
xnor U11116 (N_11116,N_8439,N_7564);
and U11117 (N_11117,N_6621,N_9245);
and U11118 (N_11118,N_8019,N_8608);
nand U11119 (N_11119,N_7334,N_8224);
xor U11120 (N_11120,N_7089,N_9149);
nor U11121 (N_11121,N_7194,N_7426);
and U11122 (N_11122,N_6372,N_7273);
nor U11123 (N_11123,N_7321,N_6339);
xor U11124 (N_11124,N_9153,N_8670);
or U11125 (N_11125,N_7798,N_8097);
xnor U11126 (N_11126,N_6951,N_8028);
xnor U11127 (N_11127,N_8588,N_7307);
nor U11128 (N_11128,N_7694,N_9288);
and U11129 (N_11129,N_7140,N_9250);
and U11130 (N_11130,N_7055,N_8304);
xnor U11131 (N_11131,N_9357,N_6300);
and U11132 (N_11132,N_8784,N_9114);
or U11133 (N_11133,N_9349,N_7205);
nor U11134 (N_11134,N_8422,N_7510);
xor U11135 (N_11135,N_7962,N_6593);
and U11136 (N_11136,N_8095,N_8524);
xor U11137 (N_11137,N_8459,N_7283);
and U11138 (N_11138,N_8286,N_7360);
xor U11139 (N_11139,N_6733,N_7141);
xnor U11140 (N_11140,N_7669,N_8687);
nor U11141 (N_11141,N_7743,N_6975);
and U11142 (N_11142,N_6274,N_8365);
and U11143 (N_11143,N_9019,N_7844);
and U11144 (N_11144,N_7325,N_8758);
and U11145 (N_11145,N_7501,N_8919);
xor U11146 (N_11146,N_7626,N_8338);
and U11147 (N_11147,N_7460,N_7505);
and U11148 (N_11148,N_6962,N_9364);
nand U11149 (N_11149,N_8897,N_7584);
nor U11150 (N_11150,N_6627,N_8272);
xnor U11151 (N_11151,N_8550,N_7463);
nand U11152 (N_11152,N_8202,N_8325);
xnor U11153 (N_11153,N_6780,N_9227);
nand U11154 (N_11154,N_7677,N_7672);
or U11155 (N_11155,N_8512,N_7337);
nand U11156 (N_11156,N_7148,N_6323);
or U11157 (N_11157,N_6509,N_6787);
or U11158 (N_11158,N_6970,N_7649);
nand U11159 (N_11159,N_7950,N_6932);
and U11160 (N_11160,N_7919,N_7097);
and U11161 (N_11161,N_6657,N_7771);
xnor U11162 (N_11162,N_8022,N_8114);
nor U11163 (N_11163,N_7480,N_8990);
nand U11164 (N_11164,N_8537,N_8442);
or U11165 (N_11165,N_7649,N_8052);
nand U11166 (N_11166,N_6904,N_7141);
nand U11167 (N_11167,N_8704,N_8410);
nor U11168 (N_11168,N_9062,N_8340);
xnor U11169 (N_11169,N_8135,N_6704);
nand U11170 (N_11170,N_6749,N_6872);
xor U11171 (N_11171,N_7531,N_8322);
xnor U11172 (N_11172,N_8215,N_9085);
nand U11173 (N_11173,N_8130,N_7834);
nor U11174 (N_11174,N_7905,N_6418);
or U11175 (N_11175,N_6781,N_8245);
xnor U11176 (N_11176,N_9203,N_8119);
and U11177 (N_11177,N_9015,N_6538);
xor U11178 (N_11178,N_7819,N_7153);
nand U11179 (N_11179,N_6281,N_7319);
nand U11180 (N_11180,N_7477,N_8045);
and U11181 (N_11181,N_6662,N_6933);
xnor U11182 (N_11182,N_8046,N_6304);
or U11183 (N_11183,N_7999,N_7411);
xnor U11184 (N_11184,N_6584,N_7070);
nor U11185 (N_11185,N_8599,N_6587);
or U11186 (N_11186,N_7010,N_8698);
or U11187 (N_11187,N_6916,N_8587);
or U11188 (N_11188,N_7282,N_8548);
and U11189 (N_11189,N_8493,N_8317);
nor U11190 (N_11190,N_8311,N_9252);
nand U11191 (N_11191,N_7803,N_6956);
nand U11192 (N_11192,N_7322,N_6387);
xnor U11193 (N_11193,N_9355,N_6274);
xor U11194 (N_11194,N_8540,N_6892);
nand U11195 (N_11195,N_6693,N_8651);
or U11196 (N_11196,N_7467,N_7301);
and U11197 (N_11197,N_6395,N_9324);
nor U11198 (N_11198,N_8179,N_8102);
nor U11199 (N_11199,N_6251,N_8532);
nand U11200 (N_11200,N_7169,N_8383);
xor U11201 (N_11201,N_7259,N_6430);
or U11202 (N_11202,N_7309,N_6475);
nor U11203 (N_11203,N_7997,N_7579);
and U11204 (N_11204,N_7980,N_7878);
and U11205 (N_11205,N_7613,N_9011);
xnor U11206 (N_11206,N_6274,N_8888);
nand U11207 (N_11207,N_8009,N_9226);
nand U11208 (N_11208,N_8715,N_7811);
xor U11209 (N_11209,N_6576,N_7372);
xor U11210 (N_11210,N_8673,N_8742);
and U11211 (N_11211,N_7844,N_8917);
and U11212 (N_11212,N_7428,N_7927);
nand U11213 (N_11213,N_7782,N_6453);
or U11214 (N_11214,N_7900,N_8305);
nor U11215 (N_11215,N_8682,N_8408);
nor U11216 (N_11216,N_8109,N_8340);
and U11217 (N_11217,N_7723,N_7006);
nor U11218 (N_11218,N_8397,N_6791);
xor U11219 (N_11219,N_6956,N_6526);
or U11220 (N_11220,N_7664,N_6951);
and U11221 (N_11221,N_6491,N_8333);
or U11222 (N_11222,N_8989,N_7516);
nor U11223 (N_11223,N_7199,N_9249);
or U11224 (N_11224,N_6552,N_8496);
nor U11225 (N_11225,N_6354,N_7703);
nand U11226 (N_11226,N_9012,N_8645);
nand U11227 (N_11227,N_7098,N_7888);
nor U11228 (N_11228,N_7186,N_8425);
xnor U11229 (N_11229,N_7351,N_9087);
and U11230 (N_11230,N_7622,N_8631);
and U11231 (N_11231,N_6651,N_9235);
nor U11232 (N_11232,N_8638,N_8990);
xnor U11233 (N_11233,N_9040,N_8748);
and U11234 (N_11234,N_8653,N_8161);
xor U11235 (N_11235,N_7421,N_6937);
or U11236 (N_11236,N_7764,N_6559);
and U11237 (N_11237,N_8124,N_8715);
nor U11238 (N_11238,N_8407,N_6485);
xnor U11239 (N_11239,N_6511,N_7998);
nor U11240 (N_11240,N_9050,N_7712);
nand U11241 (N_11241,N_6467,N_6849);
or U11242 (N_11242,N_8003,N_7640);
nor U11243 (N_11243,N_8113,N_9304);
nor U11244 (N_11244,N_8566,N_7520);
xor U11245 (N_11245,N_8917,N_7016);
nor U11246 (N_11246,N_6501,N_6598);
nor U11247 (N_11247,N_7553,N_8478);
nor U11248 (N_11248,N_8675,N_7810);
nor U11249 (N_11249,N_7751,N_8109);
and U11250 (N_11250,N_7394,N_7440);
and U11251 (N_11251,N_6641,N_6365);
nand U11252 (N_11252,N_7706,N_7134);
nor U11253 (N_11253,N_6474,N_8075);
nor U11254 (N_11254,N_6287,N_7853);
nand U11255 (N_11255,N_8646,N_9290);
xor U11256 (N_11256,N_6945,N_8022);
nor U11257 (N_11257,N_8836,N_6503);
xnor U11258 (N_11258,N_6845,N_7773);
and U11259 (N_11259,N_9156,N_8302);
or U11260 (N_11260,N_9212,N_6966);
nand U11261 (N_11261,N_6535,N_6938);
or U11262 (N_11262,N_7577,N_6894);
or U11263 (N_11263,N_6587,N_6645);
and U11264 (N_11264,N_6669,N_7174);
nand U11265 (N_11265,N_7235,N_6354);
and U11266 (N_11266,N_7943,N_6440);
and U11267 (N_11267,N_9298,N_8758);
xnor U11268 (N_11268,N_8813,N_6402);
nand U11269 (N_11269,N_6964,N_7757);
nand U11270 (N_11270,N_7314,N_7640);
nor U11271 (N_11271,N_9079,N_9116);
xor U11272 (N_11272,N_6528,N_7389);
nand U11273 (N_11273,N_9216,N_6487);
xor U11274 (N_11274,N_7277,N_6421);
nand U11275 (N_11275,N_9131,N_7741);
nor U11276 (N_11276,N_7152,N_7780);
or U11277 (N_11277,N_8532,N_8378);
or U11278 (N_11278,N_8037,N_7158);
nand U11279 (N_11279,N_7896,N_9083);
and U11280 (N_11280,N_8234,N_7501);
or U11281 (N_11281,N_8393,N_9138);
or U11282 (N_11282,N_6526,N_7161);
nand U11283 (N_11283,N_7254,N_9284);
or U11284 (N_11284,N_9084,N_8283);
and U11285 (N_11285,N_7444,N_8105);
or U11286 (N_11286,N_6649,N_8545);
or U11287 (N_11287,N_8624,N_6367);
nor U11288 (N_11288,N_9050,N_7060);
and U11289 (N_11289,N_6411,N_6335);
nand U11290 (N_11290,N_9169,N_8667);
and U11291 (N_11291,N_7427,N_6311);
and U11292 (N_11292,N_7129,N_9350);
and U11293 (N_11293,N_8263,N_8861);
nand U11294 (N_11294,N_7783,N_7991);
xnor U11295 (N_11295,N_8484,N_7552);
or U11296 (N_11296,N_7153,N_7166);
xor U11297 (N_11297,N_9035,N_6955);
and U11298 (N_11298,N_7479,N_7134);
nor U11299 (N_11299,N_6637,N_7395);
nor U11300 (N_11300,N_8034,N_7903);
nor U11301 (N_11301,N_8763,N_9160);
xnor U11302 (N_11302,N_7056,N_8424);
or U11303 (N_11303,N_8418,N_6832);
nand U11304 (N_11304,N_6307,N_9291);
nand U11305 (N_11305,N_7174,N_8976);
and U11306 (N_11306,N_8702,N_9328);
and U11307 (N_11307,N_8019,N_7057);
and U11308 (N_11308,N_8716,N_6751);
and U11309 (N_11309,N_8644,N_8429);
nand U11310 (N_11310,N_6769,N_7158);
xor U11311 (N_11311,N_6726,N_7338);
xnor U11312 (N_11312,N_7533,N_9368);
nand U11313 (N_11313,N_8791,N_7829);
xnor U11314 (N_11314,N_8659,N_8307);
xor U11315 (N_11315,N_6375,N_9020);
and U11316 (N_11316,N_7923,N_6852);
and U11317 (N_11317,N_9348,N_9158);
nor U11318 (N_11318,N_6951,N_6491);
or U11319 (N_11319,N_7950,N_8339);
nor U11320 (N_11320,N_7078,N_6579);
nor U11321 (N_11321,N_9214,N_9018);
nor U11322 (N_11322,N_6441,N_7772);
xnor U11323 (N_11323,N_7260,N_8982);
nand U11324 (N_11324,N_8533,N_8289);
and U11325 (N_11325,N_8890,N_7320);
xnor U11326 (N_11326,N_7478,N_9101);
nand U11327 (N_11327,N_6309,N_6841);
nand U11328 (N_11328,N_7951,N_6888);
xor U11329 (N_11329,N_6466,N_8398);
nor U11330 (N_11330,N_9222,N_8428);
or U11331 (N_11331,N_8263,N_7695);
nand U11332 (N_11332,N_6554,N_7839);
or U11333 (N_11333,N_8327,N_8300);
and U11334 (N_11334,N_8642,N_7172);
or U11335 (N_11335,N_8634,N_9009);
nor U11336 (N_11336,N_8976,N_7120);
and U11337 (N_11337,N_8037,N_9337);
and U11338 (N_11338,N_8820,N_8150);
xnor U11339 (N_11339,N_7671,N_7143);
and U11340 (N_11340,N_8045,N_7780);
or U11341 (N_11341,N_6864,N_7405);
xnor U11342 (N_11342,N_8609,N_6828);
xnor U11343 (N_11343,N_6336,N_8786);
xor U11344 (N_11344,N_7533,N_6394);
and U11345 (N_11345,N_8493,N_8256);
nor U11346 (N_11346,N_7786,N_6707);
nor U11347 (N_11347,N_6659,N_6955);
and U11348 (N_11348,N_7465,N_6556);
or U11349 (N_11349,N_8573,N_7299);
nand U11350 (N_11350,N_9182,N_9299);
nor U11351 (N_11351,N_7543,N_8130);
xor U11352 (N_11352,N_8857,N_6418);
and U11353 (N_11353,N_7468,N_6360);
and U11354 (N_11354,N_8296,N_7212);
nor U11355 (N_11355,N_9303,N_8922);
nor U11356 (N_11356,N_7387,N_8917);
and U11357 (N_11357,N_9323,N_9201);
nor U11358 (N_11358,N_8134,N_7474);
xor U11359 (N_11359,N_6904,N_8839);
or U11360 (N_11360,N_8451,N_8357);
or U11361 (N_11361,N_7102,N_7875);
and U11362 (N_11362,N_7052,N_8024);
nor U11363 (N_11363,N_7220,N_8707);
nor U11364 (N_11364,N_6418,N_8688);
xnor U11365 (N_11365,N_8322,N_7183);
nor U11366 (N_11366,N_6962,N_8562);
or U11367 (N_11367,N_7429,N_7611);
or U11368 (N_11368,N_6661,N_6633);
or U11369 (N_11369,N_7447,N_6959);
and U11370 (N_11370,N_6422,N_6331);
nand U11371 (N_11371,N_8406,N_7352);
nand U11372 (N_11372,N_8271,N_7345);
and U11373 (N_11373,N_7427,N_7377);
nand U11374 (N_11374,N_8429,N_8454);
or U11375 (N_11375,N_7805,N_6538);
or U11376 (N_11376,N_7367,N_6820);
and U11377 (N_11377,N_8430,N_6364);
xor U11378 (N_11378,N_7542,N_7234);
nor U11379 (N_11379,N_8098,N_6624);
or U11380 (N_11380,N_6262,N_8273);
and U11381 (N_11381,N_7154,N_8121);
or U11382 (N_11382,N_6862,N_8209);
nor U11383 (N_11383,N_9345,N_6736);
and U11384 (N_11384,N_7564,N_6481);
xor U11385 (N_11385,N_7853,N_8526);
nand U11386 (N_11386,N_7703,N_8569);
or U11387 (N_11387,N_6323,N_8315);
xnor U11388 (N_11388,N_7791,N_7876);
xor U11389 (N_11389,N_6768,N_7305);
nor U11390 (N_11390,N_7047,N_7503);
nand U11391 (N_11391,N_7641,N_8949);
xor U11392 (N_11392,N_8581,N_7191);
xor U11393 (N_11393,N_7397,N_7647);
and U11394 (N_11394,N_6776,N_7127);
and U11395 (N_11395,N_7063,N_7345);
nand U11396 (N_11396,N_8298,N_6464);
nor U11397 (N_11397,N_8086,N_8254);
nand U11398 (N_11398,N_9349,N_9356);
nand U11399 (N_11399,N_7861,N_6521);
or U11400 (N_11400,N_9143,N_8629);
and U11401 (N_11401,N_7678,N_7040);
nand U11402 (N_11402,N_6722,N_7288);
nor U11403 (N_11403,N_8364,N_8315);
xnor U11404 (N_11404,N_7611,N_8746);
or U11405 (N_11405,N_7764,N_9036);
nand U11406 (N_11406,N_7278,N_9082);
or U11407 (N_11407,N_8696,N_8361);
and U11408 (N_11408,N_6829,N_7427);
and U11409 (N_11409,N_7873,N_8007);
and U11410 (N_11410,N_6552,N_9312);
nand U11411 (N_11411,N_9246,N_7317);
xnor U11412 (N_11412,N_7145,N_8387);
nor U11413 (N_11413,N_7721,N_6914);
or U11414 (N_11414,N_8582,N_6359);
nor U11415 (N_11415,N_7332,N_7982);
xor U11416 (N_11416,N_8823,N_6379);
and U11417 (N_11417,N_8691,N_7526);
xor U11418 (N_11418,N_7108,N_8273);
nand U11419 (N_11419,N_9021,N_6958);
nor U11420 (N_11420,N_7596,N_7943);
or U11421 (N_11421,N_9328,N_7549);
xnor U11422 (N_11422,N_6760,N_6327);
or U11423 (N_11423,N_8051,N_7275);
xor U11424 (N_11424,N_8612,N_7411);
or U11425 (N_11425,N_7242,N_7919);
and U11426 (N_11426,N_6721,N_7771);
and U11427 (N_11427,N_8240,N_6618);
or U11428 (N_11428,N_6678,N_9320);
or U11429 (N_11429,N_8178,N_9105);
nor U11430 (N_11430,N_6842,N_6887);
nand U11431 (N_11431,N_7086,N_8203);
nor U11432 (N_11432,N_7703,N_7779);
nor U11433 (N_11433,N_7156,N_8245);
nor U11434 (N_11434,N_9168,N_8417);
nand U11435 (N_11435,N_8497,N_7390);
nand U11436 (N_11436,N_8659,N_8586);
and U11437 (N_11437,N_7955,N_9014);
nor U11438 (N_11438,N_6442,N_8228);
xor U11439 (N_11439,N_6364,N_8869);
xor U11440 (N_11440,N_8759,N_9236);
and U11441 (N_11441,N_7290,N_6746);
xor U11442 (N_11442,N_8387,N_6837);
nand U11443 (N_11443,N_8785,N_7539);
xor U11444 (N_11444,N_7424,N_7960);
xor U11445 (N_11445,N_8524,N_6543);
nand U11446 (N_11446,N_6467,N_7564);
and U11447 (N_11447,N_7436,N_8315);
nand U11448 (N_11448,N_9190,N_7112);
xnor U11449 (N_11449,N_8425,N_8246);
or U11450 (N_11450,N_7462,N_8651);
xor U11451 (N_11451,N_8484,N_8982);
or U11452 (N_11452,N_8956,N_8122);
or U11453 (N_11453,N_9258,N_8408);
nor U11454 (N_11454,N_6818,N_7554);
and U11455 (N_11455,N_8109,N_8798);
and U11456 (N_11456,N_8956,N_8663);
xnor U11457 (N_11457,N_6917,N_8855);
and U11458 (N_11458,N_8829,N_6312);
nor U11459 (N_11459,N_8569,N_6811);
nor U11460 (N_11460,N_6726,N_8506);
or U11461 (N_11461,N_7104,N_9258);
or U11462 (N_11462,N_9290,N_6285);
or U11463 (N_11463,N_9033,N_7791);
or U11464 (N_11464,N_8808,N_9092);
and U11465 (N_11465,N_7235,N_8677);
or U11466 (N_11466,N_9353,N_8206);
and U11467 (N_11467,N_6470,N_8124);
xor U11468 (N_11468,N_8278,N_8384);
and U11469 (N_11469,N_8145,N_7991);
xor U11470 (N_11470,N_8572,N_6313);
xnor U11471 (N_11471,N_8928,N_7349);
nor U11472 (N_11472,N_6639,N_9279);
and U11473 (N_11473,N_6996,N_8448);
and U11474 (N_11474,N_7932,N_9052);
or U11475 (N_11475,N_8816,N_7871);
nor U11476 (N_11476,N_6956,N_7512);
and U11477 (N_11477,N_6575,N_9057);
xor U11478 (N_11478,N_8952,N_7649);
or U11479 (N_11479,N_9019,N_7216);
xor U11480 (N_11480,N_6537,N_7251);
or U11481 (N_11481,N_7216,N_8392);
and U11482 (N_11482,N_9158,N_6772);
nand U11483 (N_11483,N_9263,N_8512);
nand U11484 (N_11484,N_6472,N_8361);
and U11485 (N_11485,N_8974,N_7430);
and U11486 (N_11486,N_6889,N_9298);
or U11487 (N_11487,N_9290,N_8460);
or U11488 (N_11488,N_7025,N_9150);
nand U11489 (N_11489,N_7895,N_7937);
and U11490 (N_11490,N_6935,N_9287);
nor U11491 (N_11491,N_8830,N_8219);
nor U11492 (N_11492,N_7275,N_7508);
nor U11493 (N_11493,N_7876,N_6626);
nor U11494 (N_11494,N_6915,N_7606);
xor U11495 (N_11495,N_7908,N_8499);
xor U11496 (N_11496,N_7048,N_6485);
xor U11497 (N_11497,N_7302,N_6323);
nor U11498 (N_11498,N_7270,N_6336);
and U11499 (N_11499,N_7264,N_8783);
or U11500 (N_11500,N_8758,N_6487);
or U11501 (N_11501,N_6364,N_9111);
and U11502 (N_11502,N_7120,N_7289);
or U11503 (N_11503,N_7083,N_8694);
xor U11504 (N_11504,N_7759,N_8426);
and U11505 (N_11505,N_7952,N_7004);
xnor U11506 (N_11506,N_6799,N_6784);
and U11507 (N_11507,N_6827,N_8473);
nor U11508 (N_11508,N_9122,N_8259);
nand U11509 (N_11509,N_7961,N_7988);
xnor U11510 (N_11510,N_6760,N_6858);
nand U11511 (N_11511,N_6907,N_9185);
or U11512 (N_11512,N_6448,N_8856);
and U11513 (N_11513,N_8372,N_7794);
nor U11514 (N_11514,N_8991,N_7968);
or U11515 (N_11515,N_8864,N_6537);
or U11516 (N_11516,N_8174,N_7288);
nand U11517 (N_11517,N_6527,N_7514);
and U11518 (N_11518,N_6405,N_8845);
nand U11519 (N_11519,N_9164,N_6620);
or U11520 (N_11520,N_7557,N_8488);
nand U11521 (N_11521,N_8215,N_7573);
xor U11522 (N_11522,N_9337,N_6518);
nand U11523 (N_11523,N_7360,N_8965);
nand U11524 (N_11524,N_9062,N_7704);
nor U11525 (N_11525,N_6988,N_6725);
nand U11526 (N_11526,N_7116,N_9037);
xnor U11527 (N_11527,N_8668,N_7909);
nor U11528 (N_11528,N_6772,N_8187);
xor U11529 (N_11529,N_7009,N_8959);
nor U11530 (N_11530,N_7211,N_8421);
xor U11531 (N_11531,N_7661,N_8350);
or U11532 (N_11532,N_7277,N_8520);
nand U11533 (N_11533,N_8898,N_6340);
nand U11534 (N_11534,N_9028,N_9009);
nand U11535 (N_11535,N_6624,N_8989);
nor U11536 (N_11536,N_8696,N_7628);
nor U11537 (N_11537,N_6533,N_6901);
nand U11538 (N_11538,N_8127,N_7878);
nor U11539 (N_11539,N_6705,N_9143);
nor U11540 (N_11540,N_7389,N_8098);
or U11541 (N_11541,N_7026,N_8419);
xor U11542 (N_11542,N_8606,N_7277);
and U11543 (N_11543,N_8163,N_9184);
or U11544 (N_11544,N_8346,N_8973);
and U11545 (N_11545,N_7474,N_7347);
and U11546 (N_11546,N_6657,N_8009);
nand U11547 (N_11547,N_8490,N_7503);
nor U11548 (N_11548,N_7026,N_6535);
and U11549 (N_11549,N_6290,N_7330);
and U11550 (N_11550,N_8106,N_7825);
or U11551 (N_11551,N_7833,N_6403);
and U11552 (N_11552,N_8962,N_9349);
or U11553 (N_11553,N_7882,N_6297);
or U11554 (N_11554,N_6506,N_8568);
nor U11555 (N_11555,N_7153,N_6317);
nand U11556 (N_11556,N_6865,N_9309);
nand U11557 (N_11557,N_8420,N_8652);
and U11558 (N_11558,N_9318,N_6863);
xnor U11559 (N_11559,N_8641,N_8520);
and U11560 (N_11560,N_6927,N_8041);
or U11561 (N_11561,N_7362,N_7498);
xnor U11562 (N_11562,N_8890,N_6331);
and U11563 (N_11563,N_6987,N_7032);
or U11564 (N_11564,N_8772,N_9088);
nand U11565 (N_11565,N_7121,N_9014);
nor U11566 (N_11566,N_9085,N_7586);
or U11567 (N_11567,N_9121,N_6625);
nor U11568 (N_11568,N_8140,N_6317);
or U11569 (N_11569,N_6843,N_9278);
nand U11570 (N_11570,N_7707,N_6302);
nor U11571 (N_11571,N_6478,N_9241);
nand U11572 (N_11572,N_7304,N_7133);
xnor U11573 (N_11573,N_6723,N_6913);
xor U11574 (N_11574,N_6463,N_8836);
nor U11575 (N_11575,N_8891,N_6653);
and U11576 (N_11576,N_6832,N_9301);
nor U11577 (N_11577,N_9210,N_8488);
xnor U11578 (N_11578,N_7533,N_9076);
or U11579 (N_11579,N_6951,N_8156);
and U11580 (N_11580,N_9056,N_9052);
and U11581 (N_11581,N_6496,N_7099);
or U11582 (N_11582,N_8340,N_6537);
and U11583 (N_11583,N_9065,N_8461);
nand U11584 (N_11584,N_6651,N_7866);
and U11585 (N_11585,N_8627,N_7916);
nor U11586 (N_11586,N_6777,N_8785);
or U11587 (N_11587,N_7609,N_7761);
and U11588 (N_11588,N_7211,N_8475);
xor U11589 (N_11589,N_6573,N_7303);
nand U11590 (N_11590,N_6306,N_8540);
nor U11591 (N_11591,N_7919,N_6478);
nand U11592 (N_11592,N_9309,N_6265);
nor U11593 (N_11593,N_9160,N_8826);
or U11594 (N_11594,N_6911,N_6368);
xnor U11595 (N_11595,N_8323,N_8123);
xnor U11596 (N_11596,N_6679,N_7853);
nor U11597 (N_11597,N_6906,N_6649);
and U11598 (N_11598,N_7007,N_6689);
or U11599 (N_11599,N_8866,N_7493);
and U11600 (N_11600,N_8750,N_9066);
nor U11601 (N_11601,N_7534,N_9046);
and U11602 (N_11602,N_8194,N_8107);
xnor U11603 (N_11603,N_6964,N_9021);
nor U11604 (N_11604,N_7462,N_8710);
xor U11605 (N_11605,N_9017,N_6380);
nor U11606 (N_11606,N_9118,N_8823);
xnor U11607 (N_11607,N_7116,N_7943);
and U11608 (N_11608,N_7091,N_8106);
nand U11609 (N_11609,N_6821,N_8413);
and U11610 (N_11610,N_8054,N_8690);
and U11611 (N_11611,N_6451,N_9169);
or U11612 (N_11612,N_6603,N_8010);
or U11613 (N_11613,N_6830,N_8286);
and U11614 (N_11614,N_8225,N_8629);
nor U11615 (N_11615,N_7434,N_8959);
xor U11616 (N_11616,N_7689,N_9041);
nor U11617 (N_11617,N_8907,N_9294);
nand U11618 (N_11618,N_9082,N_9271);
xor U11619 (N_11619,N_6547,N_8301);
and U11620 (N_11620,N_6505,N_9068);
xor U11621 (N_11621,N_7130,N_6291);
or U11622 (N_11622,N_8464,N_8895);
or U11623 (N_11623,N_7422,N_7313);
xor U11624 (N_11624,N_7139,N_7460);
nand U11625 (N_11625,N_7041,N_6367);
or U11626 (N_11626,N_6878,N_8097);
or U11627 (N_11627,N_8529,N_8157);
nor U11628 (N_11628,N_7504,N_8489);
or U11629 (N_11629,N_7619,N_6679);
and U11630 (N_11630,N_7549,N_8109);
or U11631 (N_11631,N_8774,N_6759);
and U11632 (N_11632,N_7401,N_8488);
nor U11633 (N_11633,N_9032,N_6962);
xor U11634 (N_11634,N_7804,N_8429);
nor U11635 (N_11635,N_7729,N_6931);
and U11636 (N_11636,N_9169,N_7203);
nand U11637 (N_11637,N_7860,N_7778);
xor U11638 (N_11638,N_7138,N_7205);
nand U11639 (N_11639,N_7920,N_7091);
or U11640 (N_11640,N_7302,N_6971);
xnor U11641 (N_11641,N_6543,N_7426);
xor U11642 (N_11642,N_8749,N_9075);
or U11643 (N_11643,N_9215,N_7317);
xor U11644 (N_11644,N_8790,N_7333);
and U11645 (N_11645,N_8857,N_6483);
nand U11646 (N_11646,N_7309,N_7749);
or U11647 (N_11647,N_6589,N_7420);
xnor U11648 (N_11648,N_6659,N_8383);
and U11649 (N_11649,N_8483,N_7893);
xor U11650 (N_11650,N_7657,N_9366);
nand U11651 (N_11651,N_6370,N_6938);
or U11652 (N_11652,N_6522,N_8167);
nor U11653 (N_11653,N_8292,N_8788);
nand U11654 (N_11654,N_6911,N_8852);
or U11655 (N_11655,N_8507,N_9336);
nand U11656 (N_11656,N_8446,N_7538);
nor U11657 (N_11657,N_6297,N_9190);
nor U11658 (N_11658,N_7933,N_9175);
nor U11659 (N_11659,N_7737,N_6979);
xnor U11660 (N_11660,N_6374,N_9255);
or U11661 (N_11661,N_7314,N_6564);
and U11662 (N_11662,N_7442,N_9027);
nand U11663 (N_11663,N_7865,N_9261);
nor U11664 (N_11664,N_7529,N_8197);
or U11665 (N_11665,N_9225,N_7193);
xor U11666 (N_11666,N_9143,N_8475);
nand U11667 (N_11667,N_6268,N_6887);
xor U11668 (N_11668,N_8570,N_6767);
or U11669 (N_11669,N_8863,N_8861);
nor U11670 (N_11670,N_7835,N_9034);
or U11671 (N_11671,N_8795,N_7217);
nand U11672 (N_11672,N_6614,N_7718);
xor U11673 (N_11673,N_7872,N_7343);
or U11674 (N_11674,N_9012,N_8579);
xnor U11675 (N_11675,N_7667,N_6408);
xor U11676 (N_11676,N_7126,N_6456);
and U11677 (N_11677,N_6624,N_8184);
nand U11678 (N_11678,N_8733,N_8653);
xor U11679 (N_11679,N_9172,N_7263);
xnor U11680 (N_11680,N_8538,N_9059);
and U11681 (N_11681,N_7681,N_8893);
and U11682 (N_11682,N_7530,N_6956);
nor U11683 (N_11683,N_7471,N_9197);
xnor U11684 (N_11684,N_8442,N_8681);
xnor U11685 (N_11685,N_7039,N_9317);
xnor U11686 (N_11686,N_6854,N_7154);
nor U11687 (N_11687,N_6746,N_6738);
nand U11688 (N_11688,N_8015,N_8625);
nand U11689 (N_11689,N_9365,N_8643);
nand U11690 (N_11690,N_8696,N_8369);
nor U11691 (N_11691,N_7193,N_6646);
nand U11692 (N_11692,N_7117,N_7442);
or U11693 (N_11693,N_9225,N_6482);
xor U11694 (N_11694,N_9069,N_7340);
nand U11695 (N_11695,N_7202,N_6921);
nor U11696 (N_11696,N_6958,N_8748);
or U11697 (N_11697,N_8331,N_9042);
or U11698 (N_11698,N_9374,N_8969);
or U11699 (N_11699,N_7613,N_7322);
and U11700 (N_11700,N_7946,N_7502);
or U11701 (N_11701,N_7528,N_8477);
xnor U11702 (N_11702,N_7066,N_8050);
xnor U11703 (N_11703,N_8572,N_9270);
xor U11704 (N_11704,N_9026,N_6994);
and U11705 (N_11705,N_7897,N_8839);
nand U11706 (N_11706,N_9062,N_8659);
nand U11707 (N_11707,N_6978,N_8417);
nand U11708 (N_11708,N_8489,N_8902);
nand U11709 (N_11709,N_7375,N_9251);
nand U11710 (N_11710,N_7329,N_7063);
nand U11711 (N_11711,N_7830,N_9236);
xor U11712 (N_11712,N_9321,N_6290);
or U11713 (N_11713,N_6623,N_8194);
nand U11714 (N_11714,N_6949,N_8183);
nor U11715 (N_11715,N_8096,N_9355);
xnor U11716 (N_11716,N_7353,N_7665);
and U11717 (N_11717,N_7125,N_8929);
xor U11718 (N_11718,N_8475,N_9234);
and U11719 (N_11719,N_7305,N_6414);
nand U11720 (N_11720,N_8448,N_6352);
and U11721 (N_11721,N_8615,N_7423);
and U11722 (N_11722,N_6671,N_6921);
and U11723 (N_11723,N_9022,N_8350);
and U11724 (N_11724,N_6904,N_8565);
or U11725 (N_11725,N_7852,N_6614);
or U11726 (N_11726,N_6951,N_9193);
or U11727 (N_11727,N_9268,N_7639);
xnor U11728 (N_11728,N_7704,N_6531);
nor U11729 (N_11729,N_8360,N_7236);
xor U11730 (N_11730,N_7491,N_8175);
or U11731 (N_11731,N_7200,N_7879);
nor U11732 (N_11732,N_8947,N_6442);
nor U11733 (N_11733,N_7044,N_8736);
and U11734 (N_11734,N_7695,N_6967);
and U11735 (N_11735,N_7541,N_8438);
or U11736 (N_11736,N_6898,N_7565);
xnor U11737 (N_11737,N_8975,N_7175);
nor U11738 (N_11738,N_7010,N_7171);
and U11739 (N_11739,N_8754,N_8498);
or U11740 (N_11740,N_6721,N_6459);
nor U11741 (N_11741,N_8173,N_9313);
or U11742 (N_11742,N_6956,N_8811);
nand U11743 (N_11743,N_8618,N_7779);
and U11744 (N_11744,N_8561,N_8346);
nor U11745 (N_11745,N_8852,N_7109);
nand U11746 (N_11746,N_8102,N_9078);
and U11747 (N_11747,N_7802,N_8443);
xnor U11748 (N_11748,N_7956,N_6497);
nand U11749 (N_11749,N_8959,N_6837);
xnor U11750 (N_11750,N_6378,N_7045);
nor U11751 (N_11751,N_6568,N_6452);
xor U11752 (N_11752,N_6462,N_6914);
nor U11753 (N_11753,N_8158,N_8269);
nor U11754 (N_11754,N_6975,N_8206);
xor U11755 (N_11755,N_7140,N_8843);
nand U11756 (N_11756,N_7925,N_8234);
and U11757 (N_11757,N_9224,N_6587);
and U11758 (N_11758,N_6535,N_8209);
or U11759 (N_11759,N_6775,N_8893);
and U11760 (N_11760,N_6614,N_6894);
nand U11761 (N_11761,N_8368,N_8732);
and U11762 (N_11762,N_9017,N_6303);
nor U11763 (N_11763,N_8894,N_6871);
nor U11764 (N_11764,N_9265,N_8884);
and U11765 (N_11765,N_8464,N_6429);
nand U11766 (N_11766,N_7005,N_7605);
nor U11767 (N_11767,N_6794,N_7286);
xnor U11768 (N_11768,N_9218,N_6619);
and U11769 (N_11769,N_8993,N_6826);
and U11770 (N_11770,N_8434,N_7670);
nand U11771 (N_11771,N_7804,N_7764);
xnor U11772 (N_11772,N_7469,N_7404);
or U11773 (N_11773,N_6510,N_7343);
nor U11774 (N_11774,N_7316,N_8856);
xor U11775 (N_11775,N_8043,N_7270);
nand U11776 (N_11776,N_8339,N_7290);
nand U11777 (N_11777,N_7994,N_7537);
or U11778 (N_11778,N_7743,N_9200);
and U11779 (N_11779,N_6448,N_8106);
nor U11780 (N_11780,N_7844,N_7770);
nand U11781 (N_11781,N_8050,N_9001);
nor U11782 (N_11782,N_8351,N_7444);
nand U11783 (N_11783,N_6408,N_6498);
or U11784 (N_11784,N_9201,N_7613);
nand U11785 (N_11785,N_6746,N_7905);
or U11786 (N_11786,N_6421,N_8609);
xnor U11787 (N_11787,N_6414,N_9031);
xnor U11788 (N_11788,N_7568,N_9026);
and U11789 (N_11789,N_8446,N_7471);
xnor U11790 (N_11790,N_7203,N_6343);
nor U11791 (N_11791,N_8601,N_9374);
or U11792 (N_11792,N_7208,N_7909);
xor U11793 (N_11793,N_6625,N_7596);
or U11794 (N_11794,N_7804,N_8868);
and U11795 (N_11795,N_8113,N_6336);
nor U11796 (N_11796,N_6913,N_7366);
or U11797 (N_11797,N_7662,N_6615);
xor U11798 (N_11798,N_6537,N_6657);
or U11799 (N_11799,N_8656,N_6947);
nor U11800 (N_11800,N_8930,N_7367);
nand U11801 (N_11801,N_6433,N_8523);
xor U11802 (N_11802,N_7458,N_7140);
nor U11803 (N_11803,N_6859,N_7671);
nor U11804 (N_11804,N_9042,N_6768);
and U11805 (N_11805,N_7233,N_6430);
xor U11806 (N_11806,N_8796,N_6417);
or U11807 (N_11807,N_8399,N_8247);
xor U11808 (N_11808,N_7755,N_8431);
nor U11809 (N_11809,N_6883,N_7601);
or U11810 (N_11810,N_6548,N_8927);
xnor U11811 (N_11811,N_6517,N_6708);
and U11812 (N_11812,N_6422,N_6877);
or U11813 (N_11813,N_9079,N_6597);
or U11814 (N_11814,N_6951,N_7283);
and U11815 (N_11815,N_8057,N_9172);
or U11816 (N_11816,N_8119,N_7654);
nor U11817 (N_11817,N_7002,N_8009);
xor U11818 (N_11818,N_8523,N_7996);
nor U11819 (N_11819,N_8756,N_6871);
nor U11820 (N_11820,N_9223,N_9091);
and U11821 (N_11821,N_6788,N_7465);
and U11822 (N_11822,N_6431,N_8603);
nand U11823 (N_11823,N_8166,N_7511);
and U11824 (N_11824,N_8820,N_8621);
nand U11825 (N_11825,N_7426,N_8905);
nor U11826 (N_11826,N_8704,N_6494);
and U11827 (N_11827,N_6689,N_9039);
nand U11828 (N_11828,N_7224,N_7999);
or U11829 (N_11829,N_9326,N_7458);
nand U11830 (N_11830,N_7922,N_9156);
nand U11831 (N_11831,N_6838,N_8888);
and U11832 (N_11832,N_8524,N_9119);
or U11833 (N_11833,N_8731,N_8829);
xor U11834 (N_11834,N_7909,N_7650);
or U11835 (N_11835,N_7862,N_6459);
and U11836 (N_11836,N_9116,N_7746);
or U11837 (N_11837,N_9259,N_8935);
and U11838 (N_11838,N_6297,N_8649);
nor U11839 (N_11839,N_7230,N_7895);
nand U11840 (N_11840,N_6426,N_6908);
xor U11841 (N_11841,N_6982,N_6811);
and U11842 (N_11842,N_8351,N_9305);
xnor U11843 (N_11843,N_8607,N_9269);
and U11844 (N_11844,N_8827,N_7422);
xor U11845 (N_11845,N_8269,N_6980);
nor U11846 (N_11846,N_7176,N_8104);
and U11847 (N_11847,N_8718,N_8653);
nor U11848 (N_11848,N_6727,N_9063);
and U11849 (N_11849,N_7319,N_7124);
xnor U11850 (N_11850,N_8371,N_6904);
nor U11851 (N_11851,N_7777,N_6705);
and U11852 (N_11852,N_7475,N_7516);
nand U11853 (N_11853,N_7429,N_7716);
xor U11854 (N_11854,N_6314,N_9290);
nor U11855 (N_11855,N_9032,N_8642);
nor U11856 (N_11856,N_7163,N_6535);
and U11857 (N_11857,N_8861,N_6690);
xnor U11858 (N_11858,N_6945,N_7391);
xnor U11859 (N_11859,N_6301,N_7854);
nor U11860 (N_11860,N_9313,N_7015);
and U11861 (N_11861,N_6921,N_7584);
or U11862 (N_11862,N_6282,N_8902);
xor U11863 (N_11863,N_9109,N_8757);
nand U11864 (N_11864,N_8480,N_6679);
nand U11865 (N_11865,N_7727,N_7289);
or U11866 (N_11866,N_9143,N_7783);
or U11867 (N_11867,N_8319,N_8593);
xnor U11868 (N_11868,N_7357,N_9214);
nand U11869 (N_11869,N_7983,N_6575);
or U11870 (N_11870,N_9260,N_9296);
nor U11871 (N_11871,N_6902,N_6769);
nand U11872 (N_11872,N_8896,N_6637);
nor U11873 (N_11873,N_7284,N_9160);
nand U11874 (N_11874,N_7216,N_8241);
and U11875 (N_11875,N_6955,N_8459);
or U11876 (N_11876,N_7335,N_8122);
and U11877 (N_11877,N_7173,N_9125);
nand U11878 (N_11878,N_8617,N_7313);
and U11879 (N_11879,N_6312,N_8201);
and U11880 (N_11880,N_6510,N_8404);
and U11881 (N_11881,N_6926,N_7988);
or U11882 (N_11882,N_6292,N_7782);
or U11883 (N_11883,N_8945,N_7189);
nor U11884 (N_11884,N_7352,N_9211);
nor U11885 (N_11885,N_6653,N_6440);
nand U11886 (N_11886,N_7947,N_7909);
or U11887 (N_11887,N_9109,N_6520);
nor U11888 (N_11888,N_9034,N_9150);
nand U11889 (N_11889,N_7280,N_8086);
nand U11890 (N_11890,N_7804,N_8765);
or U11891 (N_11891,N_6320,N_6426);
xnor U11892 (N_11892,N_7214,N_7315);
nand U11893 (N_11893,N_7401,N_7766);
nand U11894 (N_11894,N_9113,N_6464);
xor U11895 (N_11895,N_8701,N_6435);
nand U11896 (N_11896,N_9085,N_7300);
nor U11897 (N_11897,N_7290,N_8783);
nor U11898 (N_11898,N_6736,N_7779);
and U11899 (N_11899,N_7250,N_6476);
or U11900 (N_11900,N_7745,N_8193);
and U11901 (N_11901,N_7750,N_7135);
and U11902 (N_11902,N_9067,N_7630);
nor U11903 (N_11903,N_8911,N_8906);
or U11904 (N_11904,N_8904,N_6602);
nor U11905 (N_11905,N_8215,N_8062);
nand U11906 (N_11906,N_7329,N_6919);
and U11907 (N_11907,N_9131,N_8243);
nand U11908 (N_11908,N_6947,N_7780);
and U11909 (N_11909,N_7966,N_9236);
and U11910 (N_11910,N_6879,N_7226);
nand U11911 (N_11911,N_9195,N_7588);
or U11912 (N_11912,N_8647,N_6616);
or U11913 (N_11913,N_8000,N_7603);
and U11914 (N_11914,N_8585,N_9066);
nor U11915 (N_11915,N_6414,N_9347);
nor U11916 (N_11916,N_7339,N_8711);
xnor U11917 (N_11917,N_8085,N_8552);
xor U11918 (N_11918,N_8370,N_8783);
or U11919 (N_11919,N_8995,N_8707);
nor U11920 (N_11920,N_6294,N_7101);
and U11921 (N_11921,N_8571,N_6808);
and U11922 (N_11922,N_7091,N_9060);
nor U11923 (N_11923,N_6965,N_9142);
nand U11924 (N_11924,N_9270,N_6627);
and U11925 (N_11925,N_9293,N_8113);
nor U11926 (N_11926,N_6253,N_6842);
and U11927 (N_11927,N_8509,N_6683);
and U11928 (N_11928,N_7441,N_6573);
and U11929 (N_11929,N_6778,N_9053);
nand U11930 (N_11930,N_9181,N_7472);
xnor U11931 (N_11931,N_6944,N_7930);
or U11932 (N_11932,N_6947,N_6362);
xnor U11933 (N_11933,N_7321,N_9305);
xor U11934 (N_11934,N_8328,N_7740);
or U11935 (N_11935,N_8024,N_6254);
xor U11936 (N_11936,N_7739,N_7459);
and U11937 (N_11937,N_6449,N_8342);
nor U11938 (N_11938,N_8851,N_7869);
nand U11939 (N_11939,N_6619,N_7630);
xor U11940 (N_11940,N_6406,N_8807);
nor U11941 (N_11941,N_7975,N_8561);
nand U11942 (N_11942,N_7475,N_8321);
nor U11943 (N_11943,N_8590,N_9222);
nand U11944 (N_11944,N_8497,N_8135);
xnor U11945 (N_11945,N_7751,N_7727);
nand U11946 (N_11946,N_8913,N_7386);
nor U11947 (N_11947,N_7217,N_7016);
nor U11948 (N_11948,N_9148,N_7057);
or U11949 (N_11949,N_8761,N_7226);
or U11950 (N_11950,N_6957,N_7323);
nor U11951 (N_11951,N_8363,N_6659);
and U11952 (N_11952,N_8692,N_7873);
nand U11953 (N_11953,N_7801,N_8836);
and U11954 (N_11954,N_9222,N_8906);
or U11955 (N_11955,N_7913,N_6797);
or U11956 (N_11956,N_8750,N_8811);
nor U11957 (N_11957,N_8499,N_7435);
xor U11958 (N_11958,N_7399,N_8297);
and U11959 (N_11959,N_7519,N_6791);
nand U11960 (N_11960,N_7712,N_6642);
nor U11961 (N_11961,N_7551,N_7642);
xor U11962 (N_11962,N_9127,N_9180);
or U11963 (N_11963,N_9067,N_7241);
or U11964 (N_11964,N_8747,N_7624);
xnor U11965 (N_11965,N_8077,N_8444);
xnor U11966 (N_11966,N_6366,N_6553);
or U11967 (N_11967,N_6287,N_8307);
nor U11968 (N_11968,N_8839,N_7694);
or U11969 (N_11969,N_6481,N_8348);
xor U11970 (N_11970,N_8205,N_8998);
xnor U11971 (N_11971,N_8929,N_7355);
nor U11972 (N_11972,N_9250,N_7130);
nor U11973 (N_11973,N_9227,N_8043);
xnor U11974 (N_11974,N_8969,N_7344);
nor U11975 (N_11975,N_8676,N_9358);
xnor U11976 (N_11976,N_7046,N_7902);
nor U11977 (N_11977,N_8416,N_7797);
or U11978 (N_11978,N_6852,N_8382);
nand U11979 (N_11979,N_8699,N_9097);
or U11980 (N_11980,N_8105,N_6834);
nand U11981 (N_11981,N_8158,N_6497);
xnor U11982 (N_11982,N_8719,N_6928);
or U11983 (N_11983,N_7526,N_8178);
xnor U11984 (N_11984,N_8261,N_7396);
nor U11985 (N_11985,N_8946,N_9222);
or U11986 (N_11986,N_7110,N_7701);
xnor U11987 (N_11987,N_7220,N_7938);
or U11988 (N_11988,N_6823,N_9064);
nand U11989 (N_11989,N_8347,N_8452);
or U11990 (N_11990,N_7319,N_6499);
and U11991 (N_11991,N_7179,N_8809);
nand U11992 (N_11992,N_6889,N_8019);
and U11993 (N_11993,N_6305,N_9259);
or U11994 (N_11994,N_6473,N_7032);
nand U11995 (N_11995,N_7095,N_8299);
nand U11996 (N_11996,N_7519,N_7415);
nand U11997 (N_11997,N_8435,N_6737);
and U11998 (N_11998,N_9029,N_7971);
xnor U11999 (N_11999,N_7202,N_8425);
or U12000 (N_12000,N_7255,N_8185);
and U12001 (N_12001,N_7861,N_6749);
and U12002 (N_12002,N_8231,N_7960);
xnor U12003 (N_12003,N_6799,N_7167);
or U12004 (N_12004,N_6616,N_7476);
xor U12005 (N_12005,N_7377,N_8778);
xnor U12006 (N_12006,N_8222,N_8192);
nand U12007 (N_12007,N_7827,N_8390);
nand U12008 (N_12008,N_8178,N_7095);
xnor U12009 (N_12009,N_8569,N_7628);
nor U12010 (N_12010,N_6297,N_7052);
nand U12011 (N_12011,N_9020,N_6852);
nor U12012 (N_12012,N_6432,N_6824);
or U12013 (N_12013,N_7249,N_7329);
nor U12014 (N_12014,N_6422,N_9120);
nor U12015 (N_12015,N_8496,N_6294);
or U12016 (N_12016,N_6482,N_7403);
and U12017 (N_12017,N_8460,N_6455);
xnor U12018 (N_12018,N_8392,N_6775);
or U12019 (N_12019,N_9005,N_8188);
and U12020 (N_12020,N_7909,N_6484);
xnor U12021 (N_12021,N_9164,N_7998);
nand U12022 (N_12022,N_6897,N_7431);
nand U12023 (N_12023,N_7658,N_8617);
xnor U12024 (N_12024,N_8207,N_7626);
nand U12025 (N_12025,N_6529,N_6830);
nor U12026 (N_12026,N_6488,N_8642);
and U12027 (N_12027,N_7245,N_8911);
xnor U12028 (N_12028,N_8028,N_6867);
xor U12029 (N_12029,N_7965,N_9244);
nand U12030 (N_12030,N_8163,N_7809);
nor U12031 (N_12031,N_6421,N_6971);
nand U12032 (N_12032,N_8219,N_7895);
or U12033 (N_12033,N_6434,N_8720);
nand U12034 (N_12034,N_6434,N_6598);
xor U12035 (N_12035,N_7578,N_8317);
nor U12036 (N_12036,N_6444,N_8370);
xnor U12037 (N_12037,N_9341,N_7260);
xnor U12038 (N_12038,N_6753,N_8823);
and U12039 (N_12039,N_6612,N_6887);
xnor U12040 (N_12040,N_6536,N_9152);
and U12041 (N_12041,N_8372,N_8793);
nor U12042 (N_12042,N_7239,N_6928);
xor U12043 (N_12043,N_7583,N_8472);
nor U12044 (N_12044,N_9220,N_8202);
nor U12045 (N_12045,N_8676,N_6519);
xor U12046 (N_12046,N_7222,N_7163);
and U12047 (N_12047,N_6289,N_7514);
xnor U12048 (N_12048,N_6511,N_8774);
xor U12049 (N_12049,N_6552,N_9042);
nand U12050 (N_12050,N_6267,N_6293);
and U12051 (N_12051,N_7615,N_6255);
nand U12052 (N_12052,N_7805,N_7440);
xnor U12053 (N_12053,N_8426,N_7391);
nand U12054 (N_12054,N_7843,N_7249);
nor U12055 (N_12055,N_7896,N_9076);
or U12056 (N_12056,N_8515,N_6327);
nand U12057 (N_12057,N_7813,N_8758);
and U12058 (N_12058,N_6529,N_8102);
and U12059 (N_12059,N_8383,N_7722);
xnor U12060 (N_12060,N_7145,N_6726);
and U12061 (N_12061,N_7987,N_8201);
and U12062 (N_12062,N_8344,N_7922);
xnor U12063 (N_12063,N_7921,N_6300);
or U12064 (N_12064,N_9185,N_7517);
nand U12065 (N_12065,N_7857,N_8758);
xnor U12066 (N_12066,N_8933,N_6913);
nand U12067 (N_12067,N_8805,N_7513);
nor U12068 (N_12068,N_7619,N_7662);
xor U12069 (N_12069,N_7587,N_8341);
and U12070 (N_12070,N_7837,N_7911);
or U12071 (N_12071,N_8623,N_9120);
or U12072 (N_12072,N_9153,N_7791);
and U12073 (N_12073,N_7406,N_7246);
nand U12074 (N_12074,N_8189,N_8668);
nor U12075 (N_12075,N_8637,N_7484);
nand U12076 (N_12076,N_6520,N_8112);
nor U12077 (N_12077,N_7460,N_7165);
and U12078 (N_12078,N_6479,N_6452);
nand U12079 (N_12079,N_6697,N_7203);
or U12080 (N_12080,N_8730,N_8644);
and U12081 (N_12081,N_9328,N_6620);
and U12082 (N_12082,N_7066,N_6848);
xor U12083 (N_12083,N_8070,N_7588);
xor U12084 (N_12084,N_7890,N_8765);
or U12085 (N_12085,N_8321,N_8658);
nor U12086 (N_12086,N_7127,N_6520);
or U12087 (N_12087,N_8283,N_9251);
or U12088 (N_12088,N_8011,N_8288);
nand U12089 (N_12089,N_8167,N_9108);
or U12090 (N_12090,N_8117,N_7543);
nor U12091 (N_12091,N_7832,N_6272);
nand U12092 (N_12092,N_6845,N_7947);
nor U12093 (N_12093,N_7376,N_9050);
nand U12094 (N_12094,N_6451,N_9360);
xor U12095 (N_12095,N_8032,N_6585);
nand U12096 (N_12096,N_7858,N_8751);
xor U12097 (N_12097,N_9312,N_6314);
or U12098 (N_12098,N_6741,N_9252);
or U12099 (N_12099,N_9168,N_8098);
and U12100 (N_12100,N_6468,N_8363);
nor U12101 (N_12101,N_6413,N_9249);
nor U12102 (N_12102,N_7276,N_7379);
xor U12103 (N_12103,N_7071,N_7779);
or U12104 (N_12104,N_7385,N_6403);
nand U12105 (N_12105,N_8053,N_6390);
and U12106 (N_12106,N_6616,N_7431);
nor U12107 (N_12107,N_7709,N_6422);
or U12108 (N_12108,N_6876,N_6737);
and U12109 (N_12109,N_6467,N_6549);
and U12110 (N_12110,N_8139,N_8798);
or U12111 (N_12111,N_7099,N_7076);
nor U12112 (N_12112,N_6999,N_8290);
and U12113 (N_12113,N_8350,N_8659);
or U12114 (N_12114,N_8445,N_7277);
or U12115 (N_12115,N_6323,N_9350);
nor U12116 (N_12116,N_8068,N_9117);
nor U12117 (N_12117,N_7955,N_8362);
xnor U12118 (N_12118,N_6770,N_8812);
and U12119 (N_12119,N_8257,N_7188);
xor U12120 (N_12120,N_7049,N_6809);
nand U12121 (N_12121,N_9281,N_8141);
or U12122 (N_12122,N_7592,N_7379);
or U12123 (N_12123,N_6352,N_6846);
or U12124 (N_12124,N_6946,N_9307);
nor U12125 (N_12125,N_9164,N_7456);
nor U12126 (N_12126,N_7226,N_8953);
and U12127 (N_12127,N_6594,N_9199);
and U12128 (N_12128,N_6587,N_8170);
xor U12129 (N_12129,N_8856,N_8245);
nor U12130 (N_12130,N_8804,N_6723);
nand U12131 (N_12131,N_7204,N_8129);
nand U12132 (N_12132,N_7403,N_8162);
and U12133 (N_12133,N_9202,N_7391);
nand U12134 (N_12134,N_8195,N_9278);
nor U12135 (N_12135,N_7845,N_7678);
or U12136 (N_12136,N_8541,N_8475);
or U12137 (N_12137,N_8317,N_6305);
xnor U12138 (N_12138,N_8898,N_8849);
and U12139 (N_12139,N_9214,N_8279);
nand U12140 (N_12140,N_7984,N_8623);
nor U12141 (N_12141,N_7143,N_8395);
or U12142 (N_12142,N_7856,N_8745);
or U12143 (N_12143,N_6876,N_7722);
and U12144 (N_12144,N_8352,N_6834);
or U12145 (N_12145,N_8998,N_7259);
or U12146 (N_12146,N_8851,N_7742);
xnor U12147 (N_12147,N_7032,N_9068);
and U12148 (N_12148,N_6977,N_9337);
xor U12149 (N_12149,N_9250,N_7926);
or U12150 (N_12150,N_8419,N_6491);
or U12151 (N_12151,N_7616,N_7577);
and U12152 (N_12152,N_7468,N_7614);
xnor U12153 (N_12153,N_8749,N_9096);
or U12154 (N_12154,N_8272,N_7747);
nor U12155 (N_12155,N_8355,N_7695);
or U12156 (N_12156,N_9060,N_8675);
or U12157 (N_12157,N_8195,N_6724);
and U12158 (N_12158,N_8566,N_7344);
xor U12159 (N_12159,N_6661,N_6322);
or U12160 (N_12160,N_8602,N_8015);
nand U12161 (N_12161,N_9339,N_6502);
and U12162 (N_12162,N_7483,N_9070);
nand U12163 (N_12163,N_9338,N_7940);
and U12164 (N_12164,N_8565,N_8925);
or U12165 (N_12165,N_8249,N_9177);
nand U12166 (N_12166,N_7023,N_7367);
nor U12167 (N_12167,N_7186,N_7758);
and U12168 (N_12168,N_8298,N_9130);
and U12169 (N_12169,N_6810,N_7429);
xnor U12170 (N_12170,N_6809,N_7828);
nor U12171 (N_12171,N_7759,N_6467);
xnor U12172 (N_12172,N_6874,N_7527);
xor U12173 (N_12173,N_8661,N_7262);
or U12174 (N_12174,N_7966,N_6832);
or U12175 (N_12175,N_9029,N_7936);
and U12176 (N_12176,N_8678,N_7396);
and U12177 (N_12177,N_6871,N_9096);
nor U12178 (N_12178,N_7325,N_6544);
nor U12179 (N_12179,N_8298,N_7084);
nand U12180 (N_12180,N_6467,N_7311);
nand U12181 (N_12181,N_6866,N_7236);
or U12182 (N_12182,N_7939,N_8631);
nand U12183 (N_12183,N_7918,N_6275);
nand U12184 (N_12184,N_8814,N_8117);
xor U12185 (N_12185,N_6415,N_6650);
nand U12186 (N_12186,N_6398,N_7513);
or U12187 (N_12187,N_8796,N_9300);
nand U12188 (N_12188,N_9071,N_6952);
nand U12189 (N_12189,N_7696,N_8337);
or U12190 (N_12190,N_9358,N_6255);
and U12191 (N_12191,N_8708,N_8093);
xnor U12192 (N_12192,N_8374,N_8999);
or U12193 (N_12193,N_7968,N_6782);
nand U12194 (N_12194,N_7813,N_6403);
xnor U12195 (N_12195,N_9084,N_7594);
or U12196 (N_12196,N_7680,N_7143);
nand U12197 (N_12197,N_9227,N_7231);
or U12198 (N_12198,N_8700,N_8174);
or U12199 (N_12199,N_9012,N_7329);
nand U12200 (N_12200,N_8794,N_7483);
nand U12201 (N_12201,N_6526,N_6338);
nand U12202 (N_12202,N_7890,N_7904);
nand U12203 (N_12203,N_6587,N_8351);
nor U12204 (N_12204,N_6888,N_8403);
or U12205 (N_12205,N_7896,N_6740);
nand U12206 (N_12206,N_7005,N_9103);
xnor U12207 (N_12207,N_9007,N_7032);
nand U12208 (N_12208,N_8552,N_7072);
and U12209 (N_12209,N_6942,N_6622);
nor U12210 (N_12210,N_8600,N_8723);
and U12211 (N_12211,N_6709,N_8981);
and U12212 (N_12212,N_6289,N_9279);
nand U12213 (N_12213,N_6345,N_9293);
nor U12214 (N_12214,N_6253,N_6320);
xnor U12215 (N_12215,N_8006,N_8445);
or U12216 (N_12216,N_8174,N_9163);
or U12217 (N_12217,N_8637,N_8758);
and U12218 (N_12218,N_7917,N_6740);
xnor U12219 (N_12219,N_8490,N_6898);
xnor U12220 (N_12220,N_6454,N_6453);
and U12221 (N_12221,N_7898,N_7186);
or U12222 (N_12222,N_7788,N_7317);
nand U12223 (N_12223,N_9203,N_6456);
or U12224 (N_12224,N_7725,N_7105);
xor U12225 (N_12225,N_8212,N_6739);
nand U12226 (N_12226,N_6614,N_9190);
and U12227 (N_12227,N_6628,N_6993);
and U12228 (N_12228,N_7403,N_7106);
or U12229 (N_12229,N_8553,N_6997);
xor U12230 (N_12230,N_7099,N_8838);
nor U12231 (N_12231,N_6335,N_8416);
xor U12232 (N_12232,N_8244,N_8439);
nand U12233 (N_12233,N_7223,N_9075);
or U12234 (N_12234,N_8703,N_7891);
and U12235 (N_12235,N_7997,N_7683);
nor U12236 (N_12236,N_7166,N_7235);
or U12237 (N_12237,N_7217,N_6468);
and U12238 (N_12238,N_8130,N_7795);
nand U12239 (N_12239,N_7100,N_6637);
or U12240 (N_12240,N_8036,N_7385);
nand U12241 (N_12241,N_6433,N_7640);
or U12242 (N_12242,N_8448,N_8511);
xnor U12243 (N_12243,N_8723,N_8309);
nand U12244 (N_12244,N_8721,N_7351);
xnor U12245 (N_12245,N_8582,N_9071);
nand U12246 (N_12246,N_9032,N_7317);
nor U12247 (N_12247,N_7203,N_7293);
xor U12248 (N_12248,N_8832,N_8369);
or U12249 (N_12249,N_8985,N_8853);
xor U12250 (N_12250,N_8328,N_7984);
or U12251 (N_12251,N_7921,N_7896);
or U12252 (N_12252,N_7171,N_7799);
nand U12253 (N_12253,N_7949,N_8441);
nor U12254 (N_12254,N_9009,N_7938);
nor U12255 (N_12255,N_8218,N_8972);
nand U12256 (N_12256,N_6368,N_8914);
nor U12257 (N_12257,N_6529,N_7841);
nand U12258 (N_12258,N_8039,N_7294);
or U12259 (N_12259,N_7402,N_6949);
nor U12260 (N_12260,N_7198,N_6589);
xnor U12261 (N_12261,N_8431,N_7428);
nor U12262 (N_12262,N_8261,N_8037);
or U12263 (N_12263,N_8233,N_7497);
and U12264 (N_12264,N_9239,N_6795);
or U12265 (N_12265,N_6391,N_7319);
xor U12266 (N_12266,N_6415,N_8662);
nand U12267 (N_12267,N_6905,N_8035);
or U12268 (N_12268,N_7495,N_6818);
or U12269 (N_12269,N_7606,N_8893);
nand U12270 (N_12270,N_8117,N_9330);
and U12271 (N_12271,N_6440,N_7740);
xnor U12272 (N_12272,N_6344,N_9368);
nor U12273 (N_12273,N_7970,N_8061);
xor U12274 (N_12274,N_8601,N_7988);
nand U12275 (N_12275,N_6402,N_8107);
or U12276 (N_12276,N_8661,N_7771);
nand U12277 (N_12277,N_8500,N_6792);
nand U12278 (N_12278,N_9064,N_8295);
xor U12279 (N_12279,N_7947,N_6874);
nand U12280 (N_12280,N_8287,N_7260);
or U12281 (N_12281,N_9283,N_7042);
xnor U12282 (N_12282,N_7121,N_9002);
nand U12283 (N_12283,N_9044,N_6295);
or U12284 (N_12284,N_6350,N_7699);
nand U12285 (N_12285,N_6568,N_8124);
or U12286 (N_12286,N_7270,N_9145);
and U12287 (N_12287,N_7265,N_8157);
nand U12288 (N_12288,N_6983,N_8847);
or U12289 (N_12289,N_6586,N_8719);
xnor U12290 (N_12290,N_7538,N_7383);
or U12291 (N_12291,N_8681,N_6395);
nor U12292 (N_12292,N_8731,N_8857);
and U12293 (N_12293,N_8651,N_6391);
or U12294 (N_12294,N_6650,N_8416);
xnor U12295 (N_12295,N_7579,N_7279);
xnor U12296 (N_12296,N_8487,N_7078);
nor U12297 (N_12297,N_7816,N_7083);
and U12298 (N_12298,N_8399,N_7889);
nor U12299 (N_12299,N_8197,N_6267);
nand U12300 (N_12300,N_7269,N_7897);
or U12301 (N_12301,N_8201,N_7345);
xnor U12302 (N_12302,N_7402,N_8444);
xnor U12303 (N_12303,N_6530,N_7178);
nor U12304 (N_12304,N_6319,N_7095);
or U12305 (N_12305,N_8453,N_7079);
and U12306 (N_12306,N_8727,N_9268);
nand U12307 (N_12307,N_7289,N_8219);
nand U12308 (N_12308,N_6471,N_7930);
nor U12309 (N_12309,N_7398,N_6344);
nand U12310 (N_12310,N_6736,N_7619);
or U12311 (N_12311,N_8981,N_7380);
and U12312 (N_12312,N_6280,N_7789);
or U12313 (N_12313,N_9127,N_9322);
and U12314 (N_12314,N_8125,N_7044);
xor U12315 (N_12315,N_7891,N_7071);
and U12316 (N_12316,N_6297,N_8210);
nor U12317 (N_12317,N_9078,N_8606);
and U12318 (N_12318,N_7249,N_7652);
nand U12319 (N_12319,N_8199,N_8632);
nor U12320 (N_12320,N_7070,N_7371);
nor U12321 (N_12321,N_9080,N_8123);
and U12322 (N_12322,N_6314,N_8216);
xnor U12323 (N_12323,N_8706,N_8965);
nor U12324 (N_12324,N_6590,N_7581);
or U12325 (N_12325,N_7246,N_8297);
or U12326 (N_12326,N_9190,N_7811);
xor U12327 (N_12327,N_6424,N_7323);
nand U12328 (N_12328,N_9052,N_6729);
nand U12329 (N_12329,N_7058,N_7646);
and U12330 (N_12330,N_6543,N_7275);
nand U12331 (N_12331,N_9160,N_6777);
nor U12332 (N_12332,N_8801,N_7715);
xnor U12333 (N_12333,N_8629,N_7149);
xor U12334 (N_12334,N_8003,N_7997);
nand U12335 (N_12335,N_7681,N_6815);
and U12336 (N_12336,N_9025,N_7847);
nor U12337 (N_12337,N_9224,N_6973);
xnor U12338 (N_12338,N_6916,N_8801);
and U12339 (N_12339,N_8111,N_6706);
nor U12340 (N_12340,N_8023,N_7339);
xnor U12341 (N_12341,N_6358,N_8697);
and U12342 (N_12342,N_8039,N_7381);
or U12343 (N_12343,N_8176,N_6869);
nand U12344 (N_12344,N_6908,N_8922);
nand U12345 (N_12345,N_8997,N_8882);
or U12346 (N_12346,N_8611,N_6432);
or U12347 (N_12347,N_8258,N_7531);
nor U12348 (N_12348,N_6928,N_7704);
and U12349 (N_12349,N_8062,N_6420);
nand U12350 (N_12350,N_6363,N_7314);
or U12351 (N_12351,N_7166,N_8728);
xnor U12352 (N_12352,N_6444,N_6632);
or U12353 (N_12353,N_6300,N_8986);
nand U12354 (N_12354,N_8244,N_9015);
or U12355 (N_12355,N_7017,N_7363);
or U12356 (N_12356,N_7306,N_9155);
xnor U12357 (N_12357,N_9076,N_6574);
and U12358 (N_12358,N_9071,N_7313);
nand U12359 (N_12359,N_8759,N_8559);
nor U12360 (N_12360,N_7806,N_7825);
nand U12361 (N_12361,N_7035,N_9047);
nand U12362 (N_12362,N_6250,N_6574);
and U12363 (N_12363,N_7452,N_7036);
nor U12364 (N_12364,N_6946,N_7938);
nor U12365 (N_12365,N_7188,N_8417);
and U12366 (N_12366,N_6878,N_7793);
xor U12367 (N_12367,N_6654,N_7003);
or U12368 (N_12368,N_7023,N_6637);
xnor U12369 (N_12369,N_9040,N_6772);
and U12370 (N_12370,N_8867,N_8951);
or U12371 (N_12371,N_6380,N_8465);
nand U12372 (N_12372,N_9230,N_8111);
or U12373 (N_12373,N_7958,N_7467);
or U12374 (N_12374,N_9058,N_8442);
nor U12375 (N_12375,N_8502,N_9075);
or U12376 (N_12376,N_9215,N_8607);
nand U12377 (N_12377,N_8212,N_8967);
xnor U12378 (N_12378,N_9127,N_6323);
or U12379 (N_12379,N_6471,N_7767);
nor U12380 (N_12380,N_7485,N_8063);
nand U12381 (N_12381,N_8081,N_7052);
or U12382 (N_12382,N_8332,N_7851);
or U12383 (N_12383,N_9138,N_9178);
nand U12384 (N_12384,N_9028,N_6671);
nor U12385 (N_12385,N_8612,N_9008);
xor U12386 (N_12386,N_6849,N_6846);
xor U12387 (N_12387,N_7678,N_6937);
nand U12388 (N_12388,N_8990,N_7073);
nor U12389 (N_12389,N_7167,N_8426);
and U12390 (N_12390,N_8067,N_8982);
nand U12391 (N_12391,N_8626,N_7707);
xor U12392 (N_12392,N_7786,N_9356);
nor U12393 (N_12393,N_7252,N_6537);
xor U12394 (N_12394,N_7694,N_6744);
xnor U12395 (N_12395,N_6385,N_7792);
or U12396 (N_12396,N_9145,N_6891);
xor U12397 (N_12397,N_6809,N_7756);
or U12398 (N_12398,N_7487,N_7663);
nor U12399 (N_12399,N_8761,N_6794);
nand U12400 (N_12400,N_8068,N_6743);
and U12401 (N_12401,N_7533,N_6371);
nor U12402 (N_12402,N_7843,N_7110);
nand U12403 (N_12403,N_9088,N_6330);
nand U12404 (N_12404,N_7945,N_7665);
xnor U12405 (N_12405,N_8136,N_8325);
or U12406 (N_12406,N_8029,N_8878);
nor U12407 (N_12407,N_6812,N_8274);
xnor U12408 (N_12408,N_8867,N_8037);
and U12409 (N_12409,N_7919,N_7587);
and U12410 (N_12410,N_7197,N_8100);
nand U12411 (N_12411,N_6252,N_8404);
and U12412 (N_12412,N_8293,N_7529);
and U12413 (N_12413,N_8291,N_9144);
and U12414 (N_12414,N_8825,N_7761);
xor U12415 (N_12415,N_6370,N_7010);
or U12416 (N_12416,N_6622,N_8291);
xnor U12417 (N_12417,N_8331,N_6546);
nand U12418 (N_12418,N_6270,N_7358);
or U12419 (N_12419,N_7466,N_9149);
or U12420 (N_12420,N_7365,N_6507);
nand U12421 (N_12421,N_9141,N_7052);
nand U12422 (N_12422,N_8818,N_6547);
nand U12423 (N_12423,N_7657,N_7476);
xor U12424 (N_12424,N_8599,N_6689);
and U12425 (N_12425,N_7061,N_7031);
nor U12426 (N_12426,N_8541,N_6959);
or U12427 (N_12427,N_8695,N_8779);
and U12428 (N_12428,N_9263,N_9096);
nand U12429 (N_12429,N_7830,N_8195);
xnor U12430 (N_12430,N_6299,N_8246);
or U12431 (N_12431,N_7225,N_9250);
nor U12432 (N_12432,N_6922,N_8763);
xor U12433 (N_12433,N_7898,N_7222);
or U12434 (N_12434,N_8362,N_6951);
or U12435 (N_12435,N_8054,N_8285);
xor U12436 (N_12436,N_9162,N_9247);
xor U12437 (N_12437,N_6680,N_7787);
or U12438 (N_12438,N_7638,N_7273);
nand U12439 (N_12439,N_8249,N_8326);
or U12440 (N_12440,N_6330,N_8297);
nand U12441 (N_12441,N_9186,N_6513);
and U12442 (N_12442,N_6501,N_7774);
and U12443 (N_12443,N_8610,N_7377);
nor U12444 (N_12444,N_7343,N_7179);
or U12445 (N_12445,N_6331,N_8606);
nor U12446 (N_12446,N_6540,N_6632);
and U12447 (N_12447,N_7278,N_6582);
xor U12448 (N_12448,N_6364,N_7619);
nand U12449 (N_12449,N_8744,N_9347);
nand U12450 (N_12450,N_8727,N_8910);
xnor U12451 (N_12451,N_6601,N_6618);
xnor U12452 (N_12452,N_7033,N_8041);
xor U12453 (N_12453,N_8758,N_8206);
xor U12454 (N_12454,N_7096,N_8146);
xor U12455 (N_12455,N_8247,N_8297);
nor U12456 (N_12456,N_8566,N_6760);
xnor U12457 (N_12457,N_8291,N_8056);
nor U12458 (N_12458,N_7723,N_8285);
nor U12459 (N_12459,N_7435,N_7816);
xor U12460 (N_12460,N_8726,N_9296);
nor U12461 (N_12461,N_6798,N_8811);
and U12462 (N_12462,N_7331,N_7198);
nor U12463 (N_12463,N_8940,N_8442);
nand U12464 (N_12464,N_7755,N_8594);
or U12465 (N_12465,N_7973,N_6400);
nor U12466 (N_12466,N_7384,N_6729);
or U12467 (N_12467,N_7633,N_7162);
nor U12468 (N_12468,N_6941,N_6921);
and U12469 (N_12469,N_8260,N_6336);
or U12470 (N_12470,N_6805,N_9164);
nor U12471 (N_12471,N_7899,N_7807);
xor U12472 (N_12472,N_8563,N_7873);
nand U12473 (N_12473,N_6567,N_7667);
nand U12474 (N_12474,N_7081,N_7362);
or U12475 (N_12475,N_8802,N_7939);
and U12476 (N_12476,N_7681,N_6441);
and U12477 (N_12477,N_7429,N_6396);
or U12478 (N_12478,N_8503,N_8017);
xnor U12479 (N_12479,N_7297,N_8943);
or U12480 (N_12480,N_6479,N_8599);
or U12481 (N_12481,N_6946,N_7929);
and U12482 (N_12482,N_6488,N_9092);
nand U12483 (N_12483,N_7413,N_8074);
and U12484 (N_12484,N_7091,N_6413);
nor U12485 (N_12485,N_8957,N_9207);
and U12486 (N_12486,N_6546,N_7088);
nor U12487 (N_12487,N_7577,N_7638);
nand U12488 (N_12488,N_6644,N_9088);
xnor U12489 (N_12489,N_6917,N_7757);
or U12490 (N_12490,N_6423,N_7967);
xnor U12491 (N_12491,N_6586,N_6826);
or U12492 (N_12492,N_6614,N_6453);
or U12493 (N_12493,N_6915,N_8053);
or U12494 (N_12494,N_7201,N_7974);
nor U12495 (N_12495,N_6971,N_8713);
xor U12496 (N_12496,N_9024,N_8341);
nor U12497 (N_12497,N_8841,N_6545);
and U12498 (N_12498,N_6379,N_6346);
nor U12499 (N_12499,N_8833,N_8080);
and U12500 (N_12500,N_11310,N_11768);
nor U12501 (N_12501,N_12146,N_9626);
or U12502 (N_12502,N_12166,N_12394);
nand U12503 (N_12503,N_10492,N_11252);
nor U12504 (N_12504,N_10167,N_10681);
nand U12505 (N_12505,N_11592,N_11492);
nor U12506 (N_12506,N_11861,N_9982);
nor U12507 (N_12507,N_9765,N_11260);
and U12508 (N_12508,N_10738,N_10408);
xor U12509 (N_12509,N_12110,N_11179);
nor U12510 (N_12510,N_9970,N_10468);
nor U12511 (N_12511,N_11964,N_10355);
or U12512 (N_12512,N_10773,N_9994);
nor U12513 (N_12513,N_10353,N_11421);
nor U12514 (N_12514,N_9962,N_11636);
xnor U12515 (N_12515,N_10657,N_10760);
nand U12516 (N_12516,N_11984,N_11199);
xnor U12517 (N_12517,N_10515,N_9717);
nand U12518 (N_12518,N_11056,N_11404);
nor U12519 (N_12519,N_10821,N_9439);
nand U12520 (N_12520,N_11731,N_11878);
nor U12521 (N_12521,N_11496,N_10002);
nor U12522 (N_12522,N_11844,N_12201);
and U12523 (N_12523,N_12019,N_11190);
nor U12524 (N_12524,N_11746,N_11045);
and U12525 (N_12525,N_11267,N_10146);
and U12526 (N_12526,N_11792,N_9771);
or U12527 (N_12527,N_11967,N_11330);
or U12528 (N_12528,N_12046,N_11809);
nand U12529 (N_12529,N_11426,N_9732);
or U12530 (N_12530,N_9404,N_12317);
nor U12531 (N_12531,N_10229,N_11978);
nand U12532 (N_12532,N_11687,N_9813);
and U12533 (N_12533,N_11667,N_12349);
or U12534 (N_12534,N_12112,N_9617);
or U12535 (N_12535,N_10252,N_9903);
xnor U12536 (N_12536,N_11917,N_11424);
or U12537 (N_12537,N_10351,N_12385);
or U12538 (N_12538,N_12375,N_9990);
and U12539 (N_12539,N_11901,N_12173);
nor U12540 (N_12540,N_12359,N_10494);
and U12541 (N_12541,N_9898,N_9575);
xor U12542 (N_12542,N_11897,N_10193);
or U12543 (N_12543,N_12072,N_9953);
or U12544 (N_12544,N_12495,N_10795);
nor U12545 (N_12545,N_12236,N_11293);
nor U12546 (N_12546,N_12003,N_9777);
and U12547 (N_12547,N_9787,N_10427);
xor U12548 (N_12548,N_11631,N_11627);
xor U12549 (N_12549,N_11651,N_12132);
nor U12550 (N_12550,N_10385,N_11756);
and U12551 (N_12551,N_10847,N_12439);
or U12552 (N_12552,N_10715,N_10251);
or U12553 (N_12553,N_9552,N_10861);
xnor U12554 (N_12554,N_11405,N_12223);
nor U12555 (N_12555,N_11970,N_10317);
nand U12556 (N_12556,N_11287,N_10166);
xor U12557 (N_12557,N_11245,N_11171);
nand U12558 (N_12558,N_9479,N_9750);
xor U12559 (N_12559,N_11112,N_10663);
nand U12560 (N_12560,N_12164,N_12256);
xnor U12561 (N_12561,N_12078,N_11590);
nand U12562 (N_12562,N_9545,N_11139);
xor U12563 (N_12563,N_11383,N_11923);
or U12564 (N_12564,N_10384,N_9614);
nand U12565 (N_12565,N_9497,N_11536);
or U12566 (N_12566,N_11581,N_11758);
and U12567 (N_12567,N_11838,N_9389);
and U12568 (N_12568,N_11381,N_10344);
and U12569 (N_12569,N_12446,N_12417);
xor U12570 (N_12570,N_10813,N_9837);
and U12571 (N_12571,N_9972,N_9939);
or U12572 (N_12572,N_10839,N_11356);
xor U12573 (N_12573,N_10890,N_11824);
nor U12574 (N_12574,N_10886,N_12272);
or U12575 (N_12575,N_11541,N_12020);
nand U12576 (N_12576,N_10018,N_10354);
or U12577 (N_12577,N_11888,N_12497);
nand U12578 (N_12578,N_12270,N_10441);
or U12579 (N_12579,N_12355,N_10213);
or U12580 (N_12580,N_12190,N_10017);
nand U12581 (N_12581,N_9658,N_9757);
nor U12582 (N_12582,N_9387,N_11064);
nand U12583 (N_12583,N_9843,N_10706);
and U12584 (N_12584,N_9555,N_11392);
and U12585 (N_12585,N_10841,N_12343);
nand U12586 (N_12586,N_11800,N_10238);
or U12587 (N_12587,N_12029,N_10459);
nor U12588 (N_12588,N_10770,N_11725);
or U12589 (N_12589,N_12154,N_9593);
or U12590 (N_12590,N_10872,N_10169);
xnor U12591 (N_12591,N_11476,N_11050);
xnor U12592 (N_12592,N_11240,N_11580);
nor U12593 (N_12593,N_11157,N_10114);
nand U12594 (N_12594,N_10832,N_10330);
nand U12595 (N_12595,N_12198,N_10179);
xor U12596 (N_12596,N_10652,N_9580);
or U12597 (N_12597,N_10658,N_11202);
and U12598 (N_12598,N_9768,N_11443);
or U12599 (N_12599,N_10424,N_10495);
and U12600 (N_12600,N_12010,N_10226);
nand U12601 (N_12601,N_11596,N_10570);
and U12602 (N_12602,N_10382,N_11027);
or U12603 (N_12603,N_12360,N_9861);
nor U12604 (N_12604,N_12025,N_10519);
nand U12605 (N_12605,N_11936,N_11924);
or U12606 (N_12606,N_11830,N_10371);
or U12607 (N_12607,N_10331,N_10616);
xor U12608 (N_12608,N_11434,N_9952);
nand U12609 (N_12609,N_10635,N_9654);
and U12610 (N_12610,N_10374,N_10324);
nand U12611 (N_12611,N_11301,N_10110);
xor U12612 (N_12612,N_10048,N_11207);
and U12613 (N_12613,N_11938,N_10664);
xnor U12614 (N_12614,N_10129,N_11894);
nand U12615 (N_12615,N_9902,N_11140);
nand U12616 (N_12616,N_10969,N_9803);
nor U12617 (N_12617,N_11610,N_11122);
nand U12618 (N_12618,N_9503,N_12278);
or U12619 (N_12619,N_9834,N_9859);
nand U12620 (N_12620,N_11604,N_12109);
xnor U12621 (N_12621,N_9657,N_10360);
nor U12622 (N_12622,N_11311,N_10144);
or U12623 (N_12623,N_10381,N_11686);
nor U12624 (N_12624,N_10119,N_10921);
or U12625 (N_12625,N_9685,N_11527);
xor U12626 (N_12626,N_11132,N_12231);
xnor U12627 (N_12627,N_12042,N_11819);
nor U12628 (N_12628,N_11125,N_12426);
and U12629 (N_12629,N_9499,N_12149);
xor U12630 (N_12630,N_9738,N_12208);
or U12631 (N_12631,N_9416,N_10091);
nand U12632 (N_12632,N_10923,N_9496);
and U12633 (N_12633,N_9909,N_9844);
nor U12634 (N_12634,N_11795,N_10417);
nand U12635 (N_12635,N_12318,N_9550);
or U12636 (N_12636,N_10970,N_11210);
nand U12637 (N_12637,N_11298,N_10465);
nand U12638 (N_12638,N_11224,N_10599);
xnor U12639 (N_12639,N_10206,N_12066);
or U12640 (N_12640,N_11235,N_9621);
nor U12641 (N_12641,N_11365,N_9398);
or U12642 (N_12642,N_9381,N_11441);
xnor U12643 (N_12643,N_12136,N_9882);
nand U12644 (N_12644,N_9831,N_10488);
nand U12645 (N_12645,N_10490,N_11371);
nor U12646 (N_12646,N_10009,N_10183);
or U12647 (N_12647,N_11200,N_11254);
nand U12648 (N_12648,N_12247,N_12291);
nand U12649 (N_12649,N_11562,N_9904);
nand U12650 (N_12650,N_12393,N_9470);
and U12651 (N_12651,N_10755,N_10780);
xor U12652 (N_12652,N_11312,N_11788);
nand U12653 (N_12653,N_11811,N_12391);
or U12654 (N_12654,N_12415,N_12427);
and U12655 (N_12655,N_12371,N_11832);
xor U12656 (N_12656,N_12444,N_10916);
nor U12657 (N_12657,N_11760,N_11347);
and U12658 (N_12658,N_10059,N_10551);
nor U12659 (N_12659,N_9977,N_9566);
or U12660 (N_12660,N_11712,N_10863);
xor U12661 (N_12661,N_11632,N_9463);
xnor U12662 (N_12662,N_12303,N_10801);
or U12663 (N_12663,N_11063,N_12306);
xor U12664 (N_12664,N_10025,N_11074);
and U12665 (N_12665,N_12101,N_9937);
and U12666 (N_12666,N_9529,N_10837);
nand U12667 (N_12667,N_10212,N_9438);
and U12668 (N_12668,N_9824,N_12021);
nor U12669 (N_12669,N_10240,N_12044);
xor U12670 (N_12670,N_12163,N_9933);
nor U12671 (N_12671,N_10020,N_11719);
or U12672 (N_12672,N_11715,N_10033);
nor U12673 (N_12673,N_10973,N_11412);
or U12674 (N_12674,N_11639,N_12048);
nor U12675 (N_12675,N_11448,N_11089);
and U12676 (N_12676,N_12027,N_9609);
xnor U12677 (N_12677,N_9734,N_10207);
or U12678 (N_12678,N_9516,N_10138);
nor U12679 (N_12679,N_11509,N_10516);
nand U12680 (N_12680,N_9967,N_11574);
xnor U12681 (N_12681,N_10511,N_11995);
and U12682 (N_12682,N_10527,N_10989);
xnor U12683 (N_12683,N_10369,N_9758);
nand U12684 (N_12684,N_10693,N_10953);
nand U12685 (N_12685,N_9660,N_10822);
xnor U12686 (N_12686,N_12353,N_9860);
and U12687 (N_12687,N_11048,N_12222);
xnor U12688 (N_12688,N_12412,N_12480);
and U12689 (N_12689,N_11619,N_11913);
nand U12690 (N_12690,N_10577,N_9969);
or U12691 (N_12691,N_10194,N_11021);
nor U12692 (N_12692,N_10312,N_9945);
or U12693 (N_12693,N_11902,N_11078);
and U12694 (N_12694,N_10493,N_10477);
nor U12695 (N_12695,N_11357,N_12437);
xor U12696 (N_12696,N_9987,N_9696);
and U12697 (N_12697,N_12000,N_10137);
or U12698 (N_12698,N_11262,N_12159);
and U12699 (N_12699,N_12059,N_10941);
nand U12700 (N_12700,N_9810,N_9726);
nand U12701 (N_12701,N_11378,N_9931);
or U12702 (N_12702,N_11152,N_10729);
nand U12703 (N_12703,N_10076,N_9506);
nand U12704 (N_12704,N_10753,N_10977);
and U12705 (N_12705,N_9647,N_11602);
or U12706 (N_12706,N_12230,N_10092);
or U12707 (N_12707,N_11095,N_11415);
and U12708 (N_12708,N_10036,N_11129);
nand U12709 (N_12709,N_11937,N_11400);
and U12710 (N_12710,N_11163,N_12344);
and U12711 (N_12711,N_9790,N_9454);
or U12712 (N_12712,N_10675,N_12142);
nor U12713 (N_12713,N_10241,N_11308);
xnor U12714 (N_12714,N_11316,N_9797);
nand U12715 (N_12715,N_10710,N_11722);
nand U12716 (N_12716,N_10122,N_11628);
nor U12717 (N_12717,N_11454,N_9441);
nor U12718 (N_12718,N_12499,N_10603);
xor U12719 (N_12719,N_10406,N_11588);
nor U12720 (N_12720,N_11119,N_11845);
and U12721 (N_12721,N_11219,N_10636);
nand U12722 (N_12722,N_11263,N_12399);
and U12723 (N_12723,N_11382,N_9636);
xnor U12724 (N_12724,N_12482,N_10994);
or U12725 (N_12725,N_10812,N_12177);
xor U12726 (N_12726,N_9427,N_12365);
or U12727 (N_12727,N_10906,N_12470);
nand U12728 (N_12728,N_10972,N_10161);
nor U12729 (N_12729,N_11759,N_10793);
xor U12730 (N_12730,N_9851,N_12477);
or U12731 (N_12731,N_9395,N_11281);
or U12732 (N_12732,N_12148,N_10667);
and U12733 (N_12733,N_10638,N_12220);
nand U12734 (N_12734,N_9853,N_10718);
nor U12735 (N_12735,N_11960,N_9542);
nor U12736 (N_12736,N_10368,N_10387);
and U12737 (N_12737,N_11749,N_10961);
nor U12738 (N_12738,N_11080,N_12491);
and U12739 (N_12739,N_11905,N_9527);
or U12740 (N_12740,N_10688,N_9639);
nand U12741 (N_12741,N_10261,N_10806);
xor U12742 (N_12742,N_11184,N_10031);
nand U12743 (N_12743,N_9820,N_10329);
or U12744 (N_12744,N_9783,N_10210);
and U12745 (N_12745,N_10402,N_11803);
nand U12746 (N_12746,N_11437,N_12176);
and U12747 (N_12747,N_12382,N_9822);
nand U12748 (N_12748,N_10538,N_10247);
xnor U12749 (N_12749,N_10524,N_9975);
nor U12750 (N_12750,N_9737,N_9914);
xor U12751 (N_12751,N_11319,N_9947);
nor U12752 (N_12752,N_10560,N_11497);
and U12753 (N_12753,N_11368,N_12257);
nand U12754 (N_12754,N_10304,N_10691);
nor U12755 (N_12755,N_12238,N_12418);
or U12756 (N_12756,N_12174,N_11669);
and U12757 (N_12757,N_9541,N_9469);
and U12758 (N_12758,N_10559,N_11133);
and U12759 (N_12759,N_11997,N_9623);
nor U12760 (N_12760,N_10101,N_10080);
or U12761 (N_12761,N_12341,N_10816);
or U12762 (N_12762,N_12065,N_11284);
nand U12763 (N_12763,N_10339,N_11762);
nor U12764 (N_12764,N_12161,N_9996);
or U12765 (N_12765,N_12410,N_9465);
nor U12766 (N_12766,N_9386,N_11061);
and U12767 (N_12767,N_9729,N_11695);
or U12768 (N_12768,N_12199,N_10584);
nor U12769 (N_12769,N_12056,N_9983);
and U12770 (N_12770,N_11881,N_10587);
nand U12771 (N_12771,N_10192,N_10163);
xor U12772 (N_12772,N_11721,N_10974);
or U12773 (N_12773,N_11170,N_12305);
and U12774 (N_12774,N_10833,N_10319);
xnor U12775 (N_12775,N_10649,N_10692);
and U12776 (N_12776,N_11868,N_11648);
or U12777 (N_12777,N_12041,N_11507);
nor U12778 (N_12778,N_10964,N_11673);
xor U12779 (N_12779,N_12331,N_9608);
or U12780 (N_12780,N_10798,N_9408);
nand U12781 (N_12781,N_11802,N_9974);
nor U12782 (N_12782,N_10637,N_10852);
and U12783 (N_12783,N_11005,N_12235);
nor U12784 (N_12784,N_10563,N_10513);
xor U12785 (N_12785,N_9943,N_11575);
and U12786 (N_12786,N_11586,N_12323);
and U12787 (N_12787,N_10997,N_11854);
nand U12788 (N_12788,N_9895,N_11601);
nor U12789 (N_12789,N_12478,N_10932);
or U12790 (N_12790,N_10361,N_10958);
nor U12791 (N_12791,N_10771,N_10178);
or U12792 (N_12792,N_12366,N_11908);
nand U12793 (N_12793,N_9677,N_12196);
or U12794 (N_12794,N_12339,N_9718);
nand U12795 (N_12795,N_11991,N_12189);
xnor U12796 (N_12796,N_9815,N_11833);
nand U12797 (N_12797,N_9752,N_10472);
or U12798 (N_12798,N_12435,N_9727);
xnor U12799 (N_12799,N_10660,N_12336);
or U12800 (N_12800,N_11754,N_10090);
nor U12801 (N_12801,N_11023,N_9396);
and U12802 (N_12802,N_10934,N_11556);
or U12803 (N_12803,N_10013,N_9418);
nor U12804 (N_12804,N_10032,N_10149);
and U12805 (N_12805,N_11962,N_11547);
or U12806 (N_12806,N_12368,N_10722);
nor U12807 (N_12807,N_11295,N_11083);
nor U12808 (N_12808,N_10774,N_9587);
xor U12809 (N_12809,N_11972,N_12404);
nor U12810 (N_12810,N_10897,N_11369);
or U12811 (N_12811,N_10626,N_12119);
nand U12812 (N_12812,N_11644,N_11035);
and U12813 (N_12813,N_9410,N_10030);
nand U12814 (N_12814,N_11930,N_9606);
nor U12815 (N_12815,N_10297,N_9518);
and U12816 (N_12816,N_9502,N_11573);
xnor U12817 (N_12817,N_11621,N_10040);
or U12818 (N_12818,N_11253,N_9709);
nor U12819 (N_12819,N_11032,N_10920);
nor U12820 (N_12820,N_12152,N_10666);
nand U12821 (N_12821,N_11390,N_11103);
and U12822 (N_12822,N_10234,N_12475);
xor U12823 (N_12823,N_11856,N_12097);
nand U12824 (N_12824,N_9514,N_9672);
nor U12825 (N_12825,N_11677,N_10151);
nor U12826 (N_12826,N_11320,N_11151);
or U12827 (N_12827,N_10265,N_11247);
or U12828 (N_12828,N_10271,N_9434);
or U12829 (N_12829,N_10136,N_9809);
or U12830 (N_12830,N_11939,N_9468);
and U12831 (N_12831,N_11422,N_12012);
and U12832 (N_12832,N_10437,N_10873);
and U12833 (N_12833,N_12186,N_12147);
nor U12834 (N_12834,N_10089,N_11511);
nor U12835 (N_12835,N_11694,N_10725);
nand U12836 (N_12836,N_11217,N_11506);
or U12837 (N_12837,N_11515,N_10249);
and U12838 (N_12838,N_9383,N_11654);
nor U12839 (N_12839,N_11613,N_11790);
nand U12840 (N_12840,N_10855,N_11727);
nand U12841 (N_12841,N_10095,N_11623);
xor U12842 (N_12842,N_10126,N_10338);
nor U12843 (N_12843,N_9807,N_11579);
xnor U12844 (N_12844,N_9792,N_9489);
xor U12845 (N_12845,N_10731,N_10346);
or U12846 (N_12846,N_11716,N_10087);
xnor U12847 (N_12847,N_11265,N_10109);
nor U12848 (N_12848,N_12358,N_11209);
nor U12849 (N_12849,N_11438,N_12087);
nand U12850 (N_12850,N_11161,N_10254);
and U12851 (N_12851,N_11469,N_11060);
nor U12852 (N_12852,N_10436,N_10517);
xnor U12853 (N_12853,N_10086,N_10836);
xor U12854 (N_12854,N_10094,N_11659);
and U12855 (N_12855,N_11912,N_11791);
xor U12856 (N_12856,N_12288,N_11011);
nand U12857 (N_12857,N_10829,N_11531);
and U12858 (N_12858,N_10888,N_11965);
or U12859 (N_12859,N_10274,N_11085);
and U12860 (N_12860,N_11110,N_12320);
and U12861 (N_12861,N_9946,N_12485);
nor U12862 (N_12862,N_10913,N_12311);
nor U12863 (N_12863,N_10118,N_11812);
or U12864 (N_12864,N_11289,N_12325);
nor U12865 (N_12865,N_10805,N_9573);
and U12866 (N_12866,N_11020,N_9451);
xnor U12867 (N_12867,N_12348,N_10278);
and U12868 (N_12868,N_10819,N_11823);
or U12869 (N_12869,N_11570,N_10799);
nand U12870 (N_12870,N_11387,N_10593);
nand U12871 (N_12871,N_9918,N_10775);
nand U12872 (N_12872,N_10676,N_10552);
nor U12873 (N_12873,N_12076,N_10003);
xnor U12874 (N_12874,N_11261,N_11180);
or U12875 (N_12875,N_9694,N_12004);
or U12876 (N_12876,N_10108,N_10765);
xnor U12877 (N_12877,N_9589,N_11377);
or U12878 (N_12878,N_9452,N_10464);
nand U12879 (N_12879,N_10909,N_9669);
nor U12880 (N_12880,N_12383,N_11560);
nand U12881 (N_12881,N_11314,N_12096);
xor U12882 (N_12882,N_11741,N_9444);
or U12883 (N_12883,N_10980,N_11933);
xnor U12884 (N_12884,N_10661,N_11872);
and U12885 (N_12885,N_10543,N_11037);
or U12886 (N_12886,N_10242,N_11680);
or U12887 (N_12887,N_12049,N_11007);
nor U12888 (N_12888,N_11701,N_11237);
and U12889 (N_12889,N_12034,N_11429);
nand U12890 (N_12890,N_12063,N_11693);
nor U12891 (N_12891,N_10139,N_9965);
and U12892 (N_12892,N_12217,N_10102);
nand U12893 (N_12893,N_10605,N_11408);
or U12894 (N_12894,N_12127,N_10742);
nor U12895 (N_12895,N_9845,N_9908);
nand U12896 (N_12896,N_9548,N_11512);
nand U12897 (N_12897,N_10011,N_10945);
or U12898 (N_12898,N_10630,N_10991);
xnor U12899 (N_12899,N_11798,N_10902);
xor U12900 (N_12900,N_10128,N_12293);
xor U12901 (N_12901,N_11843,N_11544);
or U12902 (N_12902,N_9684,N_12229);
nand U12903 (N_12903,N_12484,N_10150);
or U12904 (N_12904,N_9776,N_12023);
xnor U12905 (N_12905,N_10984,N_10215);
or U12906 (N_12906,N_11523,N_12030);
nand U12907 (N_12907,N_12055,N_11624);
or U12908 (N_12908,N_9435,N_9675);
xor U12909 (N_12909,N_12225,N_12018);
nor U12910 (N_12910,N_12007,N_10827);
and U12911 (N_12911,N_11649,N_12141);
or U12912 (N_12912,N_9838,N_10534);
nor U12913 (N_12913,N_11156,N_10066);
nand U12914 (N_12914,N_12354,N_11257);
nand U12915 (N_12915,N_9793,N_9932);
nand U12916 (N_12916,N_9498,N_11473);
nor U12917 (N_12917,N_10860,N_11134);
nand U12918 (N_12918,N_12304,N_10684);
or U12919 (N_12919,N_11399,N_10356);
nor U12920 (N_12920,N_12455,N_11545);
nor U12921 (N_12921,N_10255,N_11196);
and U12922 (N_12922,N_10550,N_12295);
xnor U12923 (N_12923,N_11166,N_11700);
or U12924 (N_12924,N_10895,N_9764);
nor U12925 (N_12925,N_9693,N_11044);
and U12926 (N_12926,N_9984,N_10619);
nand U12927 (N_12927,N_12273,N_10220);
or U12928 (N_12928,N_12264,N_10768);
xnor U12929 (N_12929,N_9920,N_10907);
nand U12930 (N_12930,N_9999,N_10365);
or U12931 (N_12931,N_9708,N_12054);
and U12932 (N_12932,N_11425,N_11491);
nor U12933 (N_12933,N_10883,N_11793);
nand U12934 (N_12934,N_12315,N_11774);
and U12935 (N_12935,N_11211,N_10620);
and U12936 (N_12936,N_10628,N_10335);
nor U12937 (N_12937,N_10522,N_10737);
and U12938 (N_12938,N_12466,N_10558);
xnor U12939 (N_12939,N_9665,N_12342);
and U12940 (N_12940,N_9642,N_9585);
nor U12941 (N_12941,N_10687,N_11940);
or U12942 (N_12942,N_9687,N_11489);
or U12943 (N_12943,N_10792,N_9781);
xor U12944 (N_12944,N_10327,N_10290);
and U12945 (N_12945,N_9811,N_11676);
or U12946 (N_12946,N_10549,N_11230);
and U12947 (N_12947,N_10993,N_11911);
nor U12948 (N_12948,N_12259,N_11641);
and U12949 (N_12949,N_11634,N_9714);
xnor U12950 (N_12950,N_10411,N_9655);
and U12951 (N_12951,N_11919,N_9868);
and U12952 (N_12952,N_9716,N_11124);
xnor U12953 (N_12953,N_9886,N_9462);
nand U12954 (N_12954,N_10208,N_9806);
xor U12955 (N_12955,N_11094,N_11130);
nand U12956 (N_12956,N_10508,N_9505);
xnor U12957 (N_12957,N_11892,N_10221);
and U12958 (N_12958,N_10745,N_10789);
or U12959 (N_12959,N_12175,N_11777);
nor U12960 (N_12960,N_10815,N_10176);
nand U12961 (N_12961,N_12134,N_9571);
nor U12962 (N_12962,N_11431,N_12363);
or U12963 (N_12963,N_11986,N_10954);
nor U12964 (N_12964,N_11079,N_11447);
nand U12965 (N_12965,N_10951,N_11728);
nor U12966 (N_12966,N_9588,N_12274);
xor U12967 (N_12967,N_11640,N_10211);
xnor U12968 (N_12968,N_12024,N_12431);
and U12969 (N_12969,N_10198,N_11228);
or U12970 (N_12970,N_10950,N_12079);
xor U12971 (N_12971,N_11865,N_11461);
xnor U12972 (N_12972,N_12170,N_12125);
xor U12973 (N_12973,N_9681,N_11691);
nand U12974 (N_12974,N_10099,N_11084);
and U12975 (N_12975,N_11055,N_10287);
nand U12976 (N_12976,N_9485,N_11532);
nand U12977 (N_12977,N_10712,N_9961);
nand U12978 (N_12978,N_9486,N_12100);
nand U12979 (N_12979,N_10900,N_9938);
xor U12980 (N_12980,N_11384,N_11630);
or U12981 (N_12981,N_11916,N_11625);
or U12982 (N_12982,N_9579,N_10732);
or U12983 (N_12983,N_10267,N_11780);
nand U12984 (N_12984,N_11784,N_10303);
or U12985 (N_12985,N_11565,N_10853);
nor U12986 (N_12986,N_9653,N_10250);
nand U12987 (N_12987,N_10960,N_11873);
nand U12988 (N_12988,N_9988,N_11309);
nor U12989 (N_12989,N_10432,N_9712);
nor U12990 (N_12990,N_10153,N_9992);
nor U12991 (N_12991,N_10343,N_11842);
or U12992 (N_12992,N_11290,N_12215);
or U12993 (N_12993,N_10574,N_11775);
xor U12994 (N_12994,N_9459,N_11041);
xnor U12995 (N_12995,N_11818,N_11717);
xor U12996 (N_12996,N_10797,N_10764);
nand U12997 (N_12997,N_9905,N_12233);
and U12998 (N_12998,N_10689,N_11550);
xor U12999 (N_12999,N_10352,N_12302);
and U13000 (N_13000,N_11336,N_10502);
nand U13001 (N_13001,N_11520,N_9774);
or U13002 (N_13002,N_12035,N_9644);
or U13003 (N_13003,N_10088,N_11358);
or U13004 (N_13004,N_10834,N_9976);
xor U13005 (N_13005,N_11225,N_10542);
xor U13006 (N_13006,N_10785,N_12145);
xnor U13007 (N_13007,N_11147,N_10435);
nand U13008 (N_13008,N_11409,N_12219);
xor U13009 (N_13009,N_12316,N_12471);
xnor U13010 (N_13010,N_9724,N_10125);
or U13011 (N_13011,N_9888,N_12118);
nor U13012 (N_13012,N_9564,N_9877);
nand U13013 (N_13013,N_11485,N_10740);
xnor U13014 (N_13014,N_9679,N_11113);
nand U13015 (N_13015,N_12406,N_10810);
nor U13016 (N_13016,N_11971,N_11340);
and U13017 (N_13017,N_11286,N_12330);
or U13018 (N_13018,N_9874,N_10189);
and U13019 (N_13019,N_12088,N_11435);
xnor U13020 (N_13020,N_10864,N_10772);
nand U13021 (N_13021,N_9620,N_12081);
and U13022 (N_13022,N_11205,N_10948);
or U13023 (N_13023,N_9730,N_11571);
nand U13024 (N_13024,N_10724,N_9826);
and U13025 (N_13025,N_11296,N_10359);
and U13026 (N_13026,N_12252,N_10899);
or U13027 (N_13027,N_11836,N_11373);
or U13028 (N_13028,N_12129,N_12299);
and U13029 (N_13029,N_12227,N_9513);
or U13030 (N_13030,N_10751,N_9786);
or U13031 (N_13031,N_10564,N_12237);
xnor U13032 (N_13032,N_9912,N_9896);
xnor U13033 (N_13033,N_10389,N_10320);
nor U13034 (N_13034,N_11197,N_12188);
and U13035 (N_13035,N_10401,N_9667);
nand U13036 (N_13036,N_11470,N_9950);
nand U13037 (N_13037,N_9481,N_10315);
nor U13038 (N_13038,N_11370,N_11615);
nor U13039 (N_13039,N_11943,N_9958);
nor U13040 (N_13040,N_11877,N_12414);
xor U13041 (N_13041,N_10116,N_10568);
and U13042 (N_13042,N_11549,N_12413);
or U13043 (N_13043,N_11698,N_12373);
xnor U13044 (N_13044,N_9414,N_11255);
nor U13045 (N_13045,N_11729,N_9867);
nor U13046 (N_13046,N_11004,N_11510);
nand U13047 (N_13047,N_10288,N_11839);
nor U13048 (N_13048,N_9501,N_11009);
or U13049 (N_13049,N_9478,N_11226);
nor U13050 (N_13050,N_10342,N_10719);
and U13051 (N_13051,N_10674,N_11900);
or U13052 (N_13052,N_12390,N_9923);
nor U13053 (N_13053,N_12440,N_11189);
and U13054 (N_13054,N_9466,N_9409);
and U13055 (N_13055,N_10978,N_10763);
xnor U13056 (N_13056,N_11517,N_9663);
and U13057 (N_13057,N_11039,N_10143);
or U13058 (N_13058,N_10380,N_9735);
xor U13059 (N_13059,N_10607,N_10079);
nand U13060 (N_13060,N_9865,N_10824);
and U13061 (N_13061,N_12103,N_11380);
and U13062 (N_13062,N_11073,N_11018);
nor U13063 (N_13063,N_11605,N_10172);
xor U13064 (N_13064,N_11963,N_10748);
or U13065 (N_13065,N_12490,N_12267);
nand U13066 (N_13066,N_10825,N_11805);
xnor U13067 (N_13067,N_11505,N_9855);
and U13068 (N_13068,N_12073,N_9406);
or U13069 (N_13069,N_11589,N_9741);
or U13070 (N_13070,N_10956,N_11072);
nor U13071 (N_13071,N_11471,N_11097);
and U13072 (N_13072,N_11062,N_12398);
xor U13073 (N_13073,N_11402,N_11862);
xor U13074 (N_13074,N_11558,N_10243);
xnor U13075 (N_13075,N_10300,N_9785);
nor U13076 (N_13076,N_10237,N_11778);
and U13077 (N_13077,N_12139,N_10140);
and U13078 (N_13078,N_9966,N_10705);
xnor U13079 (N_13079,N_10627,N_9830);
nand U13080 (N_13080,N_11002,N_11251);
and U13081 (N_13081,N_9629,N_11776);
xor U13082 (N_13082,N_12493,N_10182);
nand U13083 (N_13083,N_10246,N_10608);
and U13084 (N_13084,N_10540,N_11087);
nor U13085 (N_13085,N_9906,N_9713);
nor U13086 (N_13086,N_10418,N_10633);
and U13087 (N_13087,N_10811,N_12184);
xor U13088 (N_13088,N_11633,N_10245);
nand U13089 (N_13089,N_11393,N_9563);
nor U13090 (N_13090,N_12322,N_11884);
xor U13091 (N_13091,N_9832,N_11444);
nand U13092 (N_13092,N_10328,N_9728);
xnor U13093 (N_13093,N_12294,N_9704);
nand U13094 (N_13094,N_11564,N_10007);
nor U13095 (N_13095,N_11763,N_9535);
nor U13096 (N_13096,N_9989,N_9847);
or U13097 (N_13097,N_9568,N_11597);
xnor U13098 (N_13098,N_11671,N_10188);
nand U13099 (N_13099,N_10392,N_12338);
nand U13100 (N_13100,N_11487,N_10008);
nand U13101 (N_13101,N_11460,N_11724);
and U13102 (N_13102,N_9530,N_10842);
or U13103 (N_13103,N_12182,N_10512);
or U13104 (N_13104,N_12472,N_11707);
xor U13105 (N_13105,N_10308,N_12172);
and U13106 (N_13106,N_12494,N_10701);
and U13107 (N_13107,N_9887,N_10881);
xnor U13108 (N_13108,N_12280,N_11898);
xor U13109 (N_13109,N_11241,N_11076);
or U13110 (N_13110,N_11000,N_9449);
xor U13111 (N_13111,N_10391,N_9490);
nor U13112 (N_13112,N_10316,N_10530);
and U13113 (N_13113,N_10141,N_10685);
nor U13114 (N_13114,N_9583,N_9523);
or U13115 (N_13115,N_10565,N_9460);
xor U13116 (N_13116,N_10407,N_12062);
xor U13117 (N_13117,N_12448,N_11566);
or U13118 (N_13118,N_11012,N_10622);
nor U13119 (N_13119,N_10130,N_10145);
nor U13120 (N_13120,N_10349,N_12327);
and U13121 (N_13121,N_11351,N_9507);
xnor U13122 (N_13122,N_12452,N_12445);
xor U13123 (N_13123,N_10393,N_11675);
nor U13124 (N_13124,N_10999,N_9413);
nor U13125 (N_13125,N_12454,N_9423);
and U13126 (N_13126,N_11584,N_11706);
nand U13127 (N_13127,N_9691,N_10400);
nor U13128 (N_13128,N_9808,N_11266);
xor U13129 (N_13129,N_9656,N_10634);
or U13130 (N_13130,N_11742,N_10518);
nand U13131 (N_13131,N_10606,N_10282);
nor U13132 (N_13132,N_12395,N_12191);
or U13133 (N_13133,N_11519,N_9572);
or U13134 (N_13134,N_10618,N_10286);
nand U13135 (N_13135,N_9562,N_11121);
nand U13136 (N_13136,N_10023,N_10922);
and U13137 (N_13137,N_9736,N_10939);
and U13138 (N_13138,N_11910,N_11374);
nand U13139 (N_13139,N_10784,N_11445);
and U13140 (N_13140,N_10443,N_11502);
nand U13141 (N_13141,N_10445,N_11066);
nand U13142 (N_13142,N_12290,N_9784);
nor U13143 (N_13143,N_11993,N_11944);
nand U13144 (N_13144,N_11490,N_10302);
nand U13145 (N_13145,N_10383,N_9775);
xor U13146 (N_13146,N_10874,N_11465);
and U13147 (N_13147,N_9697,N_9884);
or U13148 (N_13148,N_10016,N_11244);
or U13149 (N_13149,N_10154,N_9699);
and U13150 (N_13150,N_12094,N_11028);
nor U13151 (N_13151,N_10397,N_11022);
nor U13152 (N_13152,N_11394,N_10065);
nand U13153 (N_13153,N_11981,N_12137);
nand U13154 (N_13154,N_12422,N_10609);
xnor U13155 (N_13155,N_12386,N_10041);
nor U13156 (N_13156,N_11065,N_11242);
or U13157 (N_13157,N_10276,N_10690);
xor U13158 (N_13158,N_9881,N_10697);
nor U13159 (N_13159,N_12085,N_11733);
nand U13160 (N_13160,N_11459,N_11879);
nand U13161 (N_13161,N_9430,N_10656);
nand U13162 (N_13162,N_10295,N_11771);
and U13163 (N_13163,N_11123,N_11477);
or U13164 (N_13164,N_10230,N_11413);
and U13165 (N_13165,N_9377,N_9511);
xor U13166 (N_13166,N_11723,N_12181);
and U13167 (N_13167,N_12289,N_9698);
xor U13168 (N_13168,N_11591,N_11516);
or U13169 (N_13169,N_10379,N_12300);
or U13170 (N_13170,N_12441,N_10943);
xor U13171 (N_13171,N_11650,N_10127);
nand U13172 (N_13172,N_9533,N_10778);
nand U13173 (N_13173,N_12180,N_11464);
xor U13174 (N_13174,N_9772,N_9625);
and U13175 (N_13175,N_9690,N_12038);
or U13176 (N_13176,N_10337,N_11472);
and U13177 (N_13177,N_9911,N_12401);
and U13178 (N_13178,N_11105,N_10802);
nor U13179 (N_13179,N_9648,N_11482);
nor U13180 (N_13180,N_9447,N_11785);
xnor U13181 (N_13181,N_11332,N_10851);
or U13182 (N_13182,N_11683,N_11710);
xor U13183 (N_13183,N_10067,N_10452);
and U13184 (N_13184,N_9598,N_10395);
xnor U13185 (N_13185,N_9848,N_11840);
and U13186 (N_13186,N_11607,N_10394);
or U13187 (N_13187,N_11204,N_10758);
nand U13188 (N_13188,N_12266,N_11533);
or U13189 (N_13189,N_10362,N_11849);
nand U13190 (N_13190,N_9683,N_9742);
nand U13191 (N_13191,N_12436,N_11643);
and U13192 (N_13192,N_11100,N_10485);
xor U13193 (N_13193,N_11876,N_12242);
nand U13194 (N_13194,N_9828,N_10546);
nor U13195 (N_13195,N_10037,N_11427);
nand U13196 (N_13196,N_11029,N_12151);
nor U13197 (N_13197,N_12167,N_12057);
and U13198 (N_13198,N_10294,N_10233);
or U13199 (N_13199,N_10072,N_11755);
xor U13200 (N_13200,N_10562,N_12369);
nor U13201 (N_13201,N_9475,N_10501);
xnor U13202 (N_13202,N_11344,N_11026);
or U13203 (N_13203,N_9964,N_10496);
nand U13204 (N_13204,N_10882,N_9852);
or U13205 (N_13205,N_11874,N_12389);
nor U13206 (N_13206,N_11428,N_10191);
nor U13207 (N_13207,N_9424,N_9643);
nand U13208 (N_13208,N_9531,N_10591);
and U13209 (N_13209,N_11155,N_9917);
nor U13210 (N_13210,N_11668,N_9417);
nand U13211 (N_13211,N_10200,N_10318);
xnor U13212 (N_13212,N_10981,N_11337);
xor U13213 (N_13213,N_9484,N_11744);
xor U13214 (N_13214,N_12387,N_9666);
xor U13215 (N_13215,N_12321,N_10340);
xor U13216 (N_13216,N_11137,N_10878);
xor U13217 (N_13217,N_12086,N_9601);
or U13218 (N_13218,N_11272,N_9525);
or U13219 (N_13219,N_9885,N_9559);
nand U13220 (N_13220,N_11019,N_11585);
xnor U13221 (N_13221,N_11106,N_11609);
nor U13222 (N_13222,N_11522,N_10019);
xnor U13223 (N_13223,N_11885,N_9464);
nor U13224 (N_13224,N_11734,N_12489);
and U13225 (N_13225,N_10750,N_9791);
and U13226 (N_13226,N_11355,N_10111);
and U13227 (N_13227,N_10937,N_9763);
or U13228 (N_13228,N_11869,N_9613);
nand U13229 (N_13229,N_10592,N_9605);
and U13230 (N_13230,N_9600,N_11820);
or U13231 (N_13231,N_9913,N_10248);
nor U13232 (N_13232,N_10537,N_11761);
nand U13233 (N_13233,N_11183,N_10112);
nand U13234 (N_13234,N_11001,N_11276);
nor U13235 (N_13235,N_10378,N_9532);
nand U13236 (N_13236,N_10484,N_9747);
nand U13237 (N_13237,N_9456,N_10203);
and U13238 (N_13238,N_11846,N_11666);
or U13239 (N_13239,N_12047,N_9749);
and U13240 (N_13240,N_9591,N_10082);
and U13241 (N_13241,N_11304,N_9397);
nor U13242 (N_13242,N_11857,N_9801);
and U13243 (N_13243,N_10001,N_11420);
xor U13244 (N_13244,N_11154,N_12037);
or U13245 (N_13245,N_11030,N_10846);
xnor U13246 (N_13246,N_12407,N_12271);
nor U13247 (N_13247,N_9816,N_9634);
nand U13248 (N_13248,N_10925,N_9940);
and U13249 (N_13249,N_9431,N_11587);
and U13250 (N_13250,N_12352,N_11462);
xor U13251 (N_13251,N_11326,N_11864);
xnor U13252 (N_13252,N_10859,N_10790);
and U13253 (N_13253,N_11576,N_12424);
and U13254 (N_13254,N_11388,N_10942);
nand U13255 (N_13255,N_10580,N_11787);
nand U13256 (N_13256,N_11069,N_12014);
xnor U13257 (N_13257,N_11203,N_11614);
and U13258 (N_13258,N_9524,N_10236);
xor U13259 (N_13259,N_12430,N_10450);
nand U13260 (N_13260,N_11081,N_10505);
nor U13261 (N_13261,N_10840,N_12265);
nor U13262 (N_13262,N_10307,N_11274);
nand U13263 (N_13263,N_9403,N_10024);
nor U13264 (N_13264,N_9676,N_9633);
and U13265 (N_13265,N_10100,N_11847);
and U13266 (N_13266,N_11208,N_10769);
or U13267 (N_13267,N_10952,N_10651);
nand U13268 (N_13268,N_11222,N_9680);
xor U13269 (N_13269,N_9759,N_10844);
and U13270 (N_13270,N_12192,N_11976);
nand U13271 (N_13271,N_10747,N_11973);
and U13272 (N_13272,N_12108,N_11529);
nand U13273 (N_13273,N_10456,N_11297);
xnor U13274 (N_13274,N_9762,N_9951);
xor U13275 (N_13275,N_10280,N_9858);
xnor U13276 (N_13276,N_10955,N_12200);
xnor U13277 (N_13277,N_10227,N_10914);
and U13278 (N_13278,N_11740,N_9840);
and U13279 (N_13279,N_9515,N_12488);
nor U13280 (N_13280,N_11417,N_10463);
and U13281 (N_13281,N_9659,N_10646);
or U13282 (N_13282,N_10244,N_9378);
nor U13283 (N_13283,N_9570,N_10727);
and U13284 (N_13284,N_10097,N_10413);
nand U13285 (N_13285,N_12397,N_9703);
nand U13286 (N_13286,N_10415,N_12367);
nor U13287 (N_13287,N_10442,N_12450);
or U13288 (N_13288,N_9870,N_10869);
and U13289 (N_13289,N_11303,N_12350);
nor U13290 (N_13290,N_9671,N_10694);
nor U13291 (N_13291,N_9554,N_9731);
nor U13292 (N_13292,N_10322,N_10078);
nor U13293 (N_13293,N_11096,N_10293);
xnor U13294 (N_13294,N_9706,N_12263);
nand U13295 (N_13295,N_12070,N_11238);
nand U13296 (N_13296,N_10268,N_11736);
nor U13297 (N_13297,N_10621,N_10615);
or U13298 (N_13298,N_10818,N_11172);
nor U13299 (N_13299,N_10683,N_9873);
nand U13300 (N_13300,N_11323,N_9610);
xnor U13301 (N_13301,N_10131,N_10077);
xnor U13302 (N_13302,N_9935,N_9997);
xor U13303 (N_13303,N_12032,N_9412);
nor U13304 (N_13304,N_11751,N_11498);
nor U13305 (N_13305,N_11889,N_10184);
and U13306 (N_13306,N_11049,N_9476);
and U13307 (N_13307,N_10850,N_10256);
nand U13308 (N_13308,N_10366,N_10004);
xor U13309 (N_13309,N_12140,N_11831);
and U13310 (N_13310,N_11227,N_11955);
xor U13311 (N_13311,N_12400,N_11169);
nor U13312 (N_13312,N_11681,N_12005);
xnor U13313 (N_13313,N_10430,N_12421);
nand U13314 (N_13314,N_11953,N_10735);
or U13315 (N_13315,N_10848,N_11379);
nand U13316 (N_13316,N_12429,N_9537);
nor U13317 (N_13317,N_9823,N_12239);
and U13318 (N_13318,N_11834,N_11629);
or U13319 (N_13319,N_9504,N_11730);
and U13320 (N_13320,N_9862,N_10601);
and U13321 (N_13321,N_10650,N_10323);
xor U13322 (N_13322,N_9517,N_10572);
or U13323 (N_13323,N_10269,N_11015);
nor U13324 (N_13324,N_10677,N_9959);
xnor U13325 (N_13325,N_10754,N_10056);
xor U13326 (N_13326,N_9382,N_12210);
or U13327 (N_13327,N_11612,N_11212);
and U13328 (N_13328,N_9544,N_10481);
or U13329 (N_13329,N_9993,N_10604);
xor U13330 (N_13330,N_11120,N_10263);
or U13331 (N_13331,N_12016,N_9957);
xnor U13332 (N_13332,N_10301,N_9528);
or U13333 (N_13333,N_11150,N_11363);
nand U13334 (N_13334,N_9753,N_12179);
or U13335 (N_13335,N_12089,N_12337);
nand U13336 (N_13336,N_11875,N_10190);
nand U13337 (N_13337,N_11966,N_10433);
nand U13338 (N_13338,N_12009,N_11361);
nand U13339 (N_13339,N_10927,N_12104);
nand U13340 (N_13340,N_9922,N_10967);
and U13341 (N_13341,N_12202,N_11352);
nor U13342 (N_13342,N_12115,N_10305);
nor U13343 (N_13343,N_11737,N_10556);
and U13344 (N_13344,N_9986,N_11925);
xnor U13345 (N_13345,N_9422,N_11848);
or U13346 (N_13346,N_9553,N_9875);
nand U13347 (N_13347,N_11099,N_10473);
nand U13348 (N_13348,N_12361,N_9878);
nor U13349 (N_13349,N_10707,N_10639);
nand U13350 (N_13350,N_9819,N_9442);
and U13351 (N_13351,N_9615,N_11952);
nor U13352 (N_13352,N_9433,N_11718);
and U13353 (N_13353,N_10930,N_9746);
and U13354 (N_13354,N_11299,N_12377);
nor U13355 (N_13355,N_12253,N_9437);
or U13356 (N_13356,N_10216,N_9649);
xor U13357 (N_13357,N_10232,N_11595);
or U13358 (N_13358,N_11752,N_10998);
nor U13359 (N_13359,N_11269,N_12226);
or U13360 (N_13360,N_11111,N_9622);
xor U13361 (N_13361,N_10982,N_12039);
nor U13362 (N_13362,N_11185,N_11040);
xnor U13363 (N_13363,N_11054,N_12248);
xor U13364 (N_13364,N_12357,N_9930);
or U13365 (N_13365,N_9627,N_10835);
and U13366 (N_13366,N_12077,N_11221);
nand U13367 (N_13367,N_11167,N_11239);
and U13368 (N_13368,N_10310,N_10893);
xor U13369 (N_13369,N_10466,N_10061);
or U13370 (N_13370,N_12183,N_9637);
nand U13371 (N_13371,N_11975,N_10022);
nor U13372 (N_13372,N_10005,N_11201);
or U13373 (N_13373,N_10321,N_12095);
or U13374 (N_13374,N_9471,N_10849);
or U13375 (N_13375,N_9651,N_11770);
or U13376 (N_13376,N_12255,N_11249);
nor U13377 (N_13377,N_11852,N_11941);
xnor U13378 (N_13378,N_11514,N_11264);
nor U13379 (N_13379,N_12434,N_12458);
nand U13380 (N_13380,N_10047,N_12051);
nor U13381 (N_13381,N_10357,N_11705);
or U13382 (N_13382,N_11542,N_9522);
nor U13383 (N_13383,N_10050,N_11983);
or U13384 (N_13384,N_9866,N_11546);
nor U13385 (N_13385,N_11599,N_12133);
or U13386 (N_13386,N_10367,N_9492);
xnor U13387 (N_13387,N_11679,N_11896);
nor U13388 (N_13388,N_10983,N_11277);
or U13389 (N_13389,N_11929,N_9711);
nor U13390 (N_13390,N_11593,N_11292);
nor U13391 (N_13391,N_12474,N_9978);
xor U13392 (N_13392,N_11530,N_11567);
or U13393 (N_13393,N_11662,N_11333);
or U13394 (N_13394,N_9802,N_12282);
nand U13395 (N_13395,N_11014,N_10533);
nand U13396 (N_13396,N_10390,N_11713);
nor U13397 (N_13397,N_9682,N_10197);
or U13398 (N_13398,N_10553,N_11503);
or U13399 (N_13399,N_12276,N_11726);
or U13400 (N_13400,N_10877,N_10063);
nand U13401 (N_13401,N_11977,N_12473);
and U13402 (N_13402,N_11158,N_11215);
xor U13403 (N_13403,N_12283,N_9521);
or U13404 (N_13404,N_10929,N_12212);
nor U13405 (N_13405,N_11807,N_9799);
xor U13406 (N_13406,N_12351,N_10901);
nor U13407 (N_13407,N_9692,N_11653);
nand U13408 (N_13408,N_11345,N_11540);
or U13409 (N_13409,N_11216,N_10201);
xor U13410 (N_13410,N_11302,N_9445);
and U13411 (N_13411,N_10617,N_11036);
nor U13412 (N_13412,N_11895,N_9457);
nor U13413 (N_13413,N_10168,N_9547);
xor U13414 (N_13414,N_10535,N_10239);
and U13415 (N_13415,N_12487,N_12314);
and U13416 (N_13416,N_10585,N_9400);
or U13417 (N_13417,N_10205,N_9602);
and U13418 (N_13418,N_11501,N_11479);
and U13419 (N_13419,N_11948,N_9805);
nor U13420 (N_13420,N_12102,N_11367);
nor U13421 (N_13421,N_12447,N_12187);
nor U13422 (N_13422,N_11350,N_11223);
nor U13423 (N_13423,N_11816,N_9520);
nand U13424 (N_13424,N_11213,N_11890);
xor U13425 (N_13425,N_11478,N_11606);
and U13426 (N_13426,N_11979,N_9551);
and U13427 (N_13427,N_10776,N_11764);
nor U13428 (N_13428,N_10106,N_10348);
nor U13429 (N_13429,N_9384,N_10723);
and U13430 (N_13430,N_9611,N_10096);
and U13431 (N_13431,N_11871,N_9919);
nand U13432 (N_13432,N_10414,N_11034);
nor U13433 (N_13433,N_10170,N_9394);
nand U13434 (N_13434,N_10403,N_11622);
and U13435 (N_13435,N_10347,N_11535);
xnor U13436 (N_13436,N_10071,N_9899);
xnor U13437 (N_13437,N_11288,N_10557);
xnor U13438 (N_13438,N_11969,N_12214);
and U13439 (N_13439,N_9854,N_11273);
or U13440 (N_13440,N_11414,N_12017);
xor U13441 (N_13441,N_10966,N_10074);
or U13442 (N_13442,N_9876,N_12120);
nor U13443 (N_13443,N_11093,N_9796);
nand U13444 (N_13444,N_12185,N_9872);
nand U13445 (N_13445,N_11346,N_11126);
xnor U13446 (N_13446,N_11646,N_11070);
or U13447 (N_13447,N_11672,N_11837);
and U13448 (N_13448,N_9458,N_11985);
and U13449 (N_13449,N_11682,N_12013);
nor U13450 (N_13450,N_10665,N_11810);
nor U13451 (N_13451,N_11829,N_11248);
or U13452 (N_13452,N_11739,N_10273);
nor U13453 (N_13453,N_10306,N_10831);
or U13454 (N_13454,N_12130,N_9739);
and U13455 (N_13455,N_9897,N_9821);
or U13456 (N_13456,N_11165,N_11457);
nor U13457 (N_13457,N_11067,N_10672);
or U13458 (N_13458,N_9695,N_9494);
nand U13459 (N_13459,N_11982,N_10704);
xor U13460 (N_13460,N_10444,N_10165);
xnor U13461 (N_13461,N_11258,N_11789);
xnor U13462 (N_13462,N_10489,N_12254);
xor U13463 (N_13463,N_12128,N_10596);
or U13464 (N_13464,N_11362,N_9436);
xor U13465 (N_13465,N_10046,N_10332);
nand U13466 (N_13466,N_10284,N_9443);
xnor U13467 (N_13467,N_11699,N_12092);
nor U13468 (N_13468,N_11071,N_9710);
xor U13469 (N_13469,N_12310,N_12168);
nor U13470 (N_13470,N_9871,N_11142);
nand U13471 (N_13471,N_11951,N_10142);
nor U13472 (N_13472,N_11559,N_12457);
and U13473 (N_13473,N_11696,N_9577);
xor U13474 (N_13474,N_10613,N_9733);
xor U13475 (N_13475,N_10115,N_9755);
xor U13476 (N_13476,N_10043,N_11186);
and U13477 (N_13477,N_9778,N_10093);
nor U13478 (N_13478,N_11321,N_11006);
or U13479 (N_13479,N_9510,N_10673);
xor U13480 (N_13480,N_10217,N_12022);
nor U13481 (N_13481,N_12249,N_10068);
or U13482 (N_13482,N_11317,N_11270);
nor U13483 (N_13483,N_10285,N_11658);
or U13484 (N_13484,N_9842,N_12453);
nor U13485 (N_13485,N_11194,N_9894);
nand U13486 (N_13486,N_12071,N_10373);
and U13487 (N_13487,N_12498,N_11091);
or U13488 (N_13488,N_11141,N_9849);
nor U13489 (N_13489,N_9429,N_12218);
and U13490 (N_13490,N_11950,N_9581);
or U13491 (N_13491,N_9380,N_9971);
nand U13492 (N_13492,N_9599,N_11794);
nor U13493 (N_13493,N_11611,N_10132);
and U13494 (N_13494,N_11449,N_10214);
xnor U13495 (N_13495,N_10590,N_9745);
or U13496 (N_13496,N_11175,N_10686);
or U13497 (N_13497,N_12052,N_10412);
and U13498 (N_13498,N_9388,N_10070);
or U13499 (N_13499,N_11486,N_12432);
nor U13500 (N_13500,N_11508,N_10423);
or U13501 (N_13501,N_9839,N_12036);
and U13502 (N_13502,N_9624,N_12411);
nor U13503 (N_13503,N_9582,N_12213);
or U13504 (N_13504,N_12379,N_9596);
nor U13505 (N_13505,N_11195,N_11551);
or U13506 (N_13506,N_12308,N_10264);
nor U13507 (N_13507,N_10471,N_9766);
or U13508 (N_13508,N_10042,N_9991);
nor U13509 (N_13509,N_10181,N_12374);
nor U13510 (N_13510,N_10892,N_10104);
nand U13511 (N_13511,N_12116,N_11116);
or U13512 (N_13512,N_11543,N_10026);
nand U13513 (N_13513,N_12193,N_11766);
and U13514 (N_13514,N_11961,N_9814);
nand U13515 (N_13515,N_11750,N_9576);
or U13516 (N_13516,N_12328,N_11518);
xnor U13517 (N_13517,N_9827,N_11665);
or U13518 (N_13518,N_11206,N_10259);
xnor U13519 (N_13519,N_12111,N_10470);
nand U13520 (N_13520,N_10800,N_9817);
and U13521 (N_13521,N_9954,N_12107);
nand U13522 (N_13522,N_10600,N_11555);
or U13523 (N_13523,N_10180,N_9488);
nand U13524 (N_13524,N_11703,N_11674);
nor U13525 (N_13525,N_10903,N_10313);
xnor U13526 (N_13526,N_10021,N_10503);
xnor U13527 (N_13527,N_10862,N_11813);
xor U13528 (N_13528,N_11886,N_11364);
nand U13529 (N_13529,N_10398,N_11814);
and U13530 (N_13530,N_11500,N_11475);
xor U13531 (N_13531,N_10739,N_10451);
nand U13532 (N_13532,N_9428,N_10529);
nand U13533 (N_13533,N_11114,N_10885);
nand U13534 (N_13534,N_12460,N_10345);
xnor U13535 (N_13535,N_11024,N_10475);
nor U13536 (N_13536,N_10573,N_11467);
nand U13537 (N_13537,N_12313,N_12241);
and U13538 (N_13538,N_10257,N_10000);
and U13539 (N_13539,N_10438,N_9721);
or U13540 (N_13540,N_9702,N_11821);
and U13541 (N_13541,N_10555,N_10235);
nand U13542 (N_13542,N_11757,N_12245);
nand U13543 (N_13543,N_10915,N_10155);
nor U13544 (N_13544,N_10098,N_10889);
nand U13545 (N_13545,N_11403,N_9812);
xnor U13546 (N_13546,N_12334,N_11327);
and U13547 (N_13547,N_10720,N_11678);
or U13548 (N_13548,N_11046,N_12456);
xnor U13549 (N_13549,N_9619,N_11104);
or U13550 (N_13550,N_11945,N_11411);
or U13551 (N_13551,N_12476,N_11569);
or U13552 (N_13552,N_11131,N_10579);
xnor U13553 (N_13553,N_11148,N_10350);
or U13554 (N_13554,N_11841,N_10817);
nand U13555 (N_13555,N_10124,N_10260);
nor U13556 (N_13556,N_10058,N_12246);
or U13557 (N_13557,N_9942,N_11934);
xor U13558 (N_13558,N_10514,N_11554);
xor U13559 (N_13559,N_9925,N_11655);
and U13560 (N_13560,N_12043,N_12451);
and U13561 (N_13561,N_11484,N_10057);
and U13562 (N_13562,N_10497,N_10917);
nand U13563 (N_13563,N_10363,N_10756);
nor U13564 (N_13564,N_11583,N_10299);
nand U13565 (N_13565,N_11863,N_9616);
nor U13566 (N_13566,N_10777,N_12296);
xor U13567 (N_13567,N_10162,N_10583);
xnor U13568 (N_13568,N_10578,N_11537);
nand U13569 (N_13569,N_9963,N_12376);
xor U13570 (N_13570,N_11689,N_12496);
nand U13571 (N_13571,N_10879,N_9722);
nor U13572 (N_13572,N_11521,N_12465);
or U13573 (N_13573,N_9391,N_10734);
xor U13574 (N_13574,N_9590,N_11068);
xor U13575 (N_13575,N_9688,N_11504);
nor U13576 (N_13576,N_10988,N_11025);
xnor U13577 (N_13577,N_11372,N_11458);
xnor U13578 (N_13578,N_9740,N_10222);
nor U13579 (N_13579,N_10642,N_11899);
xor U13580 (N_13580,N_9756,N_10963);
nor U13581 (N_13581,N_11870,N_9375);
nor U13582 (N_13582,N_10314,N_10870);
xnor U13583 (N_13583,N_10614,N_9453);
nand U13584 (N_13584,N_12105,N_9472);
xor U13585 (N_13585,N_12228,N_11534);
or U13586 (N_13586,N_9829,N_11440);
nand U13587 (N_13587,N_12001,N_11136);
nor U13588 (N_13588,N_12098,N_10121);
nand U13589 (N_13589,N_10419,N_10759);
or U13590 (N_13590,N_10199,N_9770);
and U13591 (N_13591,N_10668,N_11456);
and U13592 (N_13592,N_11801,N_12058);
xor U13593 (N_13593,N_11488,N_10164);
and U13594 (N_13594,N_9652,N_10509);
nand U13595 (N_13595,N_12309,N_9618);
or U13596 (N_13596,N_11300,N_12240);
xor U13597 (N_13597,N_11198,N_9385);
nor U13598 (N_13598,N_11453,N_11697);
nor U13599 (N_13599,N_12143,N_10453);
nor U13600 (N_13600,N_10460,N_10854);
or U13601 (N_13601,N_9421,N_10289);
and U13602 (N_13602,N_11557,N_10113);
or U13603 (N_13603,N_11638,N_12158);
and U13604 (N_13604,N_12346,N_10440);
xnor U13605 (N_13605,N_9929,N_10986);
and U13606 (N_13606,N_10364,N_9960);
nand U13607 (N_13607,N_10548,N_10298);
and U13608 (N_13608,N_10039,N_10947);
and U13609 (N_13609,N_10678,N_10898);
xor U13610 (N_13610,N_9536,N_12075);
and U13611 (N_13611,N_10586,N_10062);
xor U13612 (N_13612,N_9586,N_9857);
xnor U13613 (N_13613,N_9512,N_9402);
xnor U13614 (N_13614,N_10160,N_10679);
nor U13615 (N_13615,N_12204,N_12467);
xnor U13616 (N_13616,N_9924,N_11906);
nand U13617 (N_13617,N_12464,N_11109);
nor U13618 (N_13618,N_10641,N_10052);
and U13619 (N_13619,N_10926,N_11092);
and U13620 (N_13620,N_12402,N_10541);
xor U13621 (N_13621,N_10653,N_10857);
nor U13622 (N_13622,N_10231,N_11942);
or U13623 (N_13623,N_10487,N_11341);
and U13624 (N_13624,N_12031,N_11256);
nor U13625 (N_13625,N_11915,N_11958);
xnor U13626 (N_13626,N_11375,N_12340);
nand U13627 (N_13627,N_10726,N_11031);
and U13628 (N_13628,N_12074,N_12197);
xnor U13629 (N_13629,N_10277,N_12138);
nand U13630 (N_13630,N_10084,N_10372);
or U13631 (N_13631,N_9635,N_10370);
xnor U13632 (N_13632,N_9574,N_9744);
or U13633 (N_13633,N_11003,N_11128);
nand U13634 (N_13634,N_10736,N_9891);
nor U13635 (N_13635,N_9420,N_12416);
nand U13636 (N_13636,N_10447,N_10702);
xor U13637 (N_13637,N_11192,N_11149);
nand U13638 (N_13638,N_10743,N_9879);
nand U13639 (N_13639,N_11781,N_9662);
nor U13640 (N_13640,N_9467,N_10334);
xor U13641 (N_13641,N_10698,N_10147);
xor U13642 (N_13642,N_10987,N_11626);
xor U13643 (N_13643,N_12131,N_9565);
nand U13644 (N_13644,N_10520,N_11059);
nor U13645 (N_13645,N_10595,N_9973);
and U13646 (N_13646,N_11101,N_12312);
nand U13647 (N_13647,N_10728,N_9595);
xor U13648 (N_13648,N_10386,N_11118);
xor U13649 (N_13649,N_11107,N_10410);
and U13650 (N_13650,N_10976,N_9473);
or U13651 (N_13651,N_11188,N_9594);
and U13652 (N_13652,N_10721,N_10134);
or U13653 (N_13653,N_12279,N_11767);
nor U13654 (N_13654,N_12216,N_10467);
nor U13655 (N_13655,N_11528,N_9934);
nand U13656 (N_13656,N_11474,N_10228);
nand U13657 (N_13657,N_12083,N_10253);
or U13658 (N_13658,N_10204,N_11466);
or U13659 (N_13659,N_10843,N_10526);
nor U13660 (N_13660,N_12205,N_10575);
nand U13661 (N_13661,N_9549,N_12347);
nor U13662 (N_13662,N_9850,N_12463);
nand U13663 (N_13663,N_11921,N_10949);
or U13664 (N_13664,N_10935,N_9968);
xnor U13665 (N_13665,N_10376,N_11946);
or U13666 (N_13666,N_9916,N_12378);
nor U13667 (N_13667,N_9638,N_10012);
nand U13668 (N_13668,N_10809,N_10266);
nor U13669 (N_13669,N_10597,N_12002);
xnor U13670 (N_13670,N_10845,N_10786);
nand U13671 (N_13671,N_12126,N_11135);
nor U13672 (N_13672,N_10283,N_9461);
xor U13673 (N_13673,N_11008,N_11082);
xnor U13674 (N_13674,N_10910,N_11745);
nand U13675 (N_13675,N_10428,N_12362);
or U13676 (N_13676,N_11418,N_9864);
and U13677 (N_13677,N_10654,N_12319);
xnor U13678 (N_13678,N_9927,N_10547);
and U13679 (N_13679,N_11138,N_11765);
nand U13680 (N_13680,N_11828,N_11893);
xnor U13681 (N_13681,N_11620,N_10625);
nor U13682 (N_13682,N_10594,N_10054);
xnor U13683 (N_13683,N_10388,N_12124);
or U13684 (N_13684,N_11259,N_12372);
and U13685 (N_13685,N_10196,N_12117);
nor U13686 (N_13686,N_10120,N_9780);
or U13687 (N_13687,N_12461,N_9645);
nor U13688 (N_13688,N_9543,N_11797);
and U13689 (N_13689,N_10659,N_11086);
nor U13690 (N_13690,N_12203,N_10730);
xor U13691 (N_13691,N_9632,N_11600);
xor U13692 (N_13692,N_9509,N_10865);
xnor U13693 (N_13693,N_11656,N_12329);
nor U13694 (N_13694,N_11617,N_11013);
and U13695 (N_13695,N_11782,N_11271);
and U13696 (N_13696,N_11989,N_10060);
nor U13697 (N_13697,N_9835,N_9455);
or U13698 (N_13698,N_11176,N_12090);
and U13699 (N_13699,N_10296,N_11173);
and U13700 (N_13700,N_11246,N_10938);
nand U13701 (N_13701,N_11957,N_9450);
nand U13702 (N_13702,N_11480,N_9794);
and U13703 (N_13703,N_11075,N_9640);
nand U13704 (N_13704,N_10038,N_12425);
xnor U13705 (N_13705,N_9701,N_11391);
nand U13706 (N_13706,N_12285,N_10478);
nor U13707 (N_13707,N_9751,N_10968);
nor U13708 (N_13708,N_10461,N_11160);
and U13709 (N_13709,N_10741,N_10744);
xor U13710 (N_13710,N_11283,N_11598);
or U13711 (N_13711,N_11548,N_11354);
xnor U13712 (N_13712,N_10700,N_9789);
xor U13713 (N_13713,N_10135,N_11214);
or U13714 (N_13714,N_11360,N_11294);
nor U13715 (N_13715,N_11720,N_12028);
nand U13716 (N_13716,N_11278,N_10224);
and U13717 (N_13717,N_10051,N_10944);
and U13718 (N_13718,N_9558,N_11513);
nand U13719 (N_13719,N_11880,N_12113);
nand U13720 (N_13720,N_10326,N_11410);
or U13721 (N_13721,N_9748,N_11732);
and U13722 (N_13722,N_9560,N_12403);
xnor U13723 (N_13723,N_11783,N_11927);
or U13724 (N_13724,N_12156,N_10894);
nand U13725 (N_13725,N_9725,N_11366);
nor U13726 (N_13726,N_10405,N_11250);
or U13727 (N_13727,N_10434,N_9664);
or U13728 (N_13728,N_11275,N_9440);
nand U13729 (N_13729,N_11637,N_11714);
xor U13730 (N_13730,N_10175,N_10598);
or U13731 (N_13731,N_10107,N_11181);
or U13732 (N_13732,N_9700,N_11827);
nor U13733 (N_13733,N_10174,N_10908);
and U13734 (N_13734,N_9641,N_11279);
nand U13735 (N_13735,N_12405,N_10711);
xor U13736 (N_13736,N_10588,N_11928);
or U13737 (N_13737,N_10523,N_9419);
xor U13738 (N_13738,N_11561,N_12396);
or U13739 (N_13739,N_11779,N_10791);
xor U13740 (N_13740,N_10924,N_11153);
nor U13741 (N_13741,N_12040,N_11416);
nor U13742 (N_13742,N_10640,N_12169);
or U13743 (N_13743,N_11324,N_12153);
xor U13744 (N_13744,N_10504,N_11243);
and U13745 (N_13745,N_12449,N_11603);
nand U13746 (N_13746,N_11996,N_9979);
nand U13747 (N_13747,N_12392,N_11954);
nand U13748 (N_13748,N_10539,N_11349);
xnor U13749 (N_13749,N_10766,N_11077);
or U13750 (N_13750,N_11102,N_11088);
and U13751 (N_13751,N_9944,N_10576);
and U13752 (N_13752,N_11376,N_9767);
nand U13753 (N_13753,N_10045,N_10933);
or U13754 (N_13754,N_11033,N_10919);
nand U13755 (N_13755,N_9928,N_10507);
and U13756 (N_13756,N_10185,N_9936);
nand U13757 (N_13757,N_11850,N_11684);
or U13758 (N_13758,N_10029,N_12364);
nand U13759 (N_13759,N_11234,N_9519);
xnor U13760 (N_13760,N_9393,N_10757);
nor U13761 (N_13761,N_11495,N_12121);
xor U13762 (N_13762,N_9426,N_10965);
and U13763 (N_13763,N_11882,N_12053);
xnor U13764 (N_13764,N_9631,N_10871);
and U13765 (N_13765,N_10454,N_11907);
and U13766 (N_13766,N_10695,N_11052);
and U13767 (N_13767,N_9604,N_10610);
xor U13768 (N_13768,N_9399,N_11858);
xnor U13769 (N_13769,N_9800,N_9483);
nor U13770 (N_13770,N_12068,N_12442);
xnor U13771 (N_13771,N_11926,N_10957);
xnor U13772 (N_13772,N_11735,N_12082);
or U13773 (N_13773,N_12443,N_10936);
xnor U13774 (N_13774,N_11043,N_9592);
xnor U13775 (N_13775,N_12084,N_12165);
and U13776 (N_13776,N_11483,N_9487);
nand U13777 (N_13777,N_10887,N_9980);
or U13778 (N_13778,N_11748,N_12298);
nor U13779 (N_13779,N_11949,N_10426);
nand U13780 (N_13780,N_11164,N_12479);
and U13781 (N_13781,N_11236,N_10336);
nand U13782 (N_13782,N_10644,N_10186);
nor U13783 (N_13783,N_11563,N_9646);
nor U13784 (N_13784,N_11090,N_9900);
xnor U13785 (N_13785,N_10446,N_12281);
xor U13786 (N_13786,N_11115,N_9448);
xor U13787 (N_13787,N_12150,N_11577);
or U13788 (N_13788,N_10680,N_11162);
nand U13789 (N_13789,N_11914,N_11051);
and U13790 (N_13790,N_10876,N_10571);
nand U13791 (N_13791,N_10044,N_11494);
xor U13792 (N_13792,N_10746,N_10581);
and U13793 (N_13793,N_10971,N_11038);
xor U13794 (N_13794,N_9825,N_11178);
nand U13795 (N_13795,N_10959,N_11994);
nor U13796 (N_13796,N_10975,N_11947);
and U13797 (N_13797,N_11652,N_11335);
nor U13798 (N_13798,N_11956,N_12224);
nor U13799 (N_13799,N_10708,N_9892);
and U13800 (N_13800,N_11017,N_10510);
and U13801 (N_13801,N_10567,N_10803);
xor U13802 (N_13802,N_10035,N_9743);
nand U13803 (N_13803,N_9673,N_10469);
xor U13804 (N_13804,N_11338,N_11329);
xor U13805 (N_13805,N_9760,N_10623);
xor U13806 (N_13806,N_11851,N_12144);
or U13807 (N_13807,N_12301,N_10611);
nand U13808 (N_13808,N_11572,N_9556);
or U13809 (N_13809,N_9500,N_11568);
xor U13810 (N_13810,N_9668,N_9493);
nand U13811 (N_13811,N_10449,N_9995);
and U13812 (N_13812,N_10814,N_9798);
and U13813 (N_13813,N_10670,N_11385);
or U13814 (N_13814,N_9956,N_12419);
xnor U13815 (N_13815,N_12433,N_11229);
xnor U13816 (N_13816,N_9534,N_11218);
nor U13817 (N_13817,N_11974,N_11702);
nand U13818 (N_13818,N_10717,N_10781);
and U13819 (N_13819,N_10482,N_11708);
nand U13820 (N_13820,N_12060,N_11860);
xnor U13821 (N_13821,N_11999,N_10498);
nor U13822 (N_13822,N_11285,N_9491);
xnor U13823 (N_13823,N_12160,N_10632);
xnor U13824 (N_13824,N_10377,N_10117);
nand U13825 (N_13825,N_11191,N_11891);
or U13826 (N_13826,N_11932,N_12356);
nor U13827 (N_13827,N_9846,N_11578);
or U13828 (N_13828,N_10399,N_11322);
or U13829 (N_13829,N_10931,N_11193);
or U13830 (N_13830,N_11738,N_10828);
nor U13831 (N_13831,N_11968,N_10292);
nor U13832 (N_13832,N_10476,N_9495);
nand U13833 (N_13833,N_10714,N_10544);
nor U13834 (N_13834,N_11451,N_11468);
nor U13835 (N_13835,N_11826,N_11430);
or U13836 (N_13836,N_10448,N_10422);
nand U13837 (N_13837,N_11396,N_10823);
nand U13838 (N_13838,N_9678,N_11058);
or U13839 (N_13839,N_9715,N_10962);
or U13840 (N_13840,N_9480,N_12292);
nand U13841 (N_13841,N_9880,N_9769);
nor U13842 (N_13842,N_10421,N_10195);
xnor U13843 (N_13843,N_9376,N_12155);
nand U13844 (N_13844,N_10462,N_11232);
and U13845 (N_13845,N_11835,N_10866);
nor U13846 (N_13846,N_11436,N_10027);
or U13847 (N_13847,N_10545,N_10554);
nor U13848 (N_13848,N_9926,N_11442);
xnor U13849 (N_13849,N_12093,N_12370);
nor U13850 (N_13850,N_9856,N_12207);
and U13851 (N_13851,N_12307,N_10083);
nor U13852 (N_13852,N_11524,N_11455);
xor U13853 (N_13853,N_12015,N_12286);
nor U13854 (N_13854,N_12135,N_11315);
or U13855 (N_13855,N_9546,N_10275);
or U13856 (N_13856,N_11887,N_12469);
xor U13857 (N_13857,N_11688,N_9392);
nand U13858 (N_13858,N_10699,N_11990);
xor U13859 (N_13859,N_10696,N_11931);
nor U13860 (N_13860,N_10279,N_12262);
or U13861 (N_13861,N_12459,N_11446);
nand U13862 (N_13862,N_10569,N_11328);
nor U13863 (N_13863,N_11903,N_11853);
nand U13864 (N_13864,N_9405,N_10281);
and U13865 (N_13865,N_10566,N_9569);
nand U13866 (N_13866,N_9661,N_11231);
nor U13867 (N_13867,N_12195,N_12297);
nand U13868 (N_13868,N_11804,N_11538);
nor U13869 (N_13869,N_9597,N_10645);
xor U13870 (N_13870,N_11525,N_10064);
xor U13871 (N_13871,N_11291,N_9567);
or U13872 (N_13872,N_9425,N_10779);
xor U13873 (N_13873,N_11657,N_12008);
xnor U13874 (N_13874,N_11493,N_9883);
nand U13875 (N_13875,N_11647,N_11552);
xor U13876 (N_13876,N_10053,N_10055);
or U13877 (N_13877,N_12114,N_11042);
or U13878 (N_13878,N_10995,N_9477);
xnor U13879 (N_13879,N_11127,N_10655);
or U13880 (N_13880,N_11920,N_12250);
xnor U13881 (N_13881,N_11822,N_9482);
xnor U13882 (N_13882,N_10582,N_9561);
nor U13883 (N_13883,N_11661,N_11670);
nand U13884 (N_13884,N_10500,N_11539);
or U13885 (N_13885,N_10396,N_9379);
nand U13886 (N_13886,N_11772,N_10270);
or U13887 (N_13887,N_12335,N_10589);
xnor U13888 (N_13888,N_9804,N_10171);
nor U13889 (N_13889,N_10479,N_11704);
and U13890 (N_13890,N_9818,N_10528);
and U13891 (N_13891,N_12438,N_11144);
nor U13892 (N_13892,N_11342,N_9540);
nor U13893 (N_13893,N_10486,N_10103);
or U13894 (N_13894,N_10458,N_9720);
nand U13895 (N_13895,N_9941,N_9612);
xnor U13896 (N_13896,N_10209,N_10474);
and U13897 (N_13897,N_11334,N_9788);
or U13898 (N_13898,N_11343,N_11280);
nor U13899 (N_13899,N_9893,N_10752);
nor U13900 (N_13900,N_10177,N_9754);
xnor U13901 (N_13901,N_10612,N_12171);
nor U13902 (N_13902,N_10807,N_11747);
nor U13903 (N_13903,N_9474,N_10979);
and U13904 (N_13904,N_10429,N_11859);
nand U13905 (N_13905,N_10992,N_10034);
xor U13906 (N_13906,N_12122,N_11690);
or U13907 (N_13907,N_11146,N_11016);
nand U13908 (N_13908,N_10709,N_10891);
xor U13909 (N_13909,N_11177,N_10783);
xnor U13910 (N_13910,N_10996,N_10716);
and U13911 (N_13911,N_10258,N_10311);
nand U13912 (N_13912,N_12106,N_10457);
nor U13913 (N_13913,N_11594,N_10911);
or U13914 (N_13914,N_11318,N_10808);
or U13915 (N_13915,N_10375,N_12045);
nor U13916 (N_13916,N_11799,N_12157);
nor U13917 (N_13917,N_10416,N_12381);
xor U13918 (N_13918,N_10262,N_11481);
xor U13919 (N_13919,N_10425,N_10990);
nand U13920 (N_13920,N_9538,N_11182);
nand U13921 (N_13921,N_10905,N_10671);
and U13922 (N_13922,N_11608,N_11935);
nor U13923 (N_13923,N_11855,N_10431);
xnor U13924 (N_13924,N_12123,N_12269);
xnor U13925 (N_13925,N_11306,N_10830);
nand U13926 (N_13926,N_10918,N_10291);
nor U13927 (N_13927,N_9907,N_10309);
nor U13928 (N_13928,N_9779,N_11057);
nor U13929 (N_13929,N_9411,N_12050);
nand U13930 (N_13930,N_10272,N_10525);
or U13931 (N_13931,N_10105,N_10794);
nand U13932 (N_13932,N_10325,N_12388);
nor U13933 (N_13933,N_11313,N_12011);
nand U13934 (N_13934,N_10787,N_11526);
xor U13935 (N_13935,N_10409,N_10647);
nand U13936 (N_13936,N_11117,N_10713);
or U13937 (N_13937,N_11010,N_9526);
and U13938 (N_13938,N_11159,N_12324);
nor U13939 (N_13939,N_9761,N_11743);
or U13940 (N_13940,N_10133,N_11867);
and U13941 (N_13941,N_10796,N_9869);
nand U13942 (N_13942,N_11268,N_11909);
xor U13943 (N_13943,N_10531,N_11463);
nor U13944 (N_13944,N_9773,N_10856);
and U13945 (N_13945,N_10069,N_10733);
xnor U13946 (N_13946,N_12243,N_9628);
xnor U13947 (N_13947,N_12080,N_10404);
or U13948 (N_13948,N_11452,N_10820);
xnor U13949 (N_13949,N_12332,N_10223);
xnor U13950 (N_13950,N_11047,N_10858);
nand U13951 (N_13951,N_11922,N_10123);
or U13952 (N_13952,N_11786,N_10158);
nor U13953 (N_13953,N_11353,N_12275);
nor U13954 (N_13954,N_11769,N_10081);
nand U13955 (N_13955,N_11108,N_10420);
nand U13956 (N_13956,N_11618,N_10767);
or U13957 (N_13957,N_9841,N_10912);
xor U13958 (N_13958,N_10075,N_12026);
or U13959 (N_13959,N_11307,N_12420);
and U13960 (N_13960,N_10904,N_9401);
or U13961 (N_13961,N_10602,N_10506);
or U13962 (N_13962,N_12268,N_12232);
or U13963 (N_13963,N_12384,N_11645);
xor U13964 (N_13964,N_11663,N_10662);
nand U13965 (N_13965,N_9949,N_11389);
or U13966 (N_13966,N_10940,N_10521);
or U13967 (N_13967,N_10480,N_12260);
and U13968 (N_13968,N_11174,N_10085);
xor U13969 (N_13969,N_10762,N_10455);
and U13970 (N_13970,N_10669,N_11616);
and U13971 (N_13971,N_11439,N_11918);
and U13972 (N_13972,N_11806,N_11187);
or U13973 (N_13973,N_9390,N_12333);
xor U13974 (N_13974,N_9670,N_10880);
nand U13975 (N_13975,N_11664,N_12234);
nor U13976 (N_13976,N_10985,N_9689);
or U13977 (N_13977,N_11450,N_11904);
or U13978 (N_13978,N_10015,N_12178);
nand U13979 (N_13979,N_11808,N_9782);
xor U13980 (N_13980,N_9981,N_11433);
nor U13981 (N_13981,N_12194,N_10804);
and U13982 (N_13982,N_11992,N_11098);
and U13983 (N_13983,N_10838,N_10532);
nand U13984 (N_13984,N_11325,N_11339);
xor U13985 (N_13985,N_10187,N_11282);
and U13986 (N_13986,N_12428,N_10202);
nand U13987 (N_13987,N_9557,N_12206);
nor U13988 (N_13988,N_12061,N_12261);
nand U13989 (N_13989,N_11305,N_10928);
nor U13990 (N_13990,N_12287,N_12258);
xnor U13991 (N_13991,N_10073,N_10749);
xnor U13992 (N_13992,N_12006,N_12162);
and U13993 (N_13993,N_12326,N_10703);
nor U13994 (N_13994,N_10225,N_12409);
and U13995 (N_13995,N_10782,N_9446);
xnor U13996 (N_13996,N_12408,N_12221);
xnor U13997 (N_13997,N_9432,N_9863);
or U13998 (N_13998,N_9707,N_12064);
or U13999 (N_13999,N_10682,N_9705);
xor U14000 (N_14000,N_12211,N_10946);
nand U14001 (N_14001,N_9539,N_9415);
and U14002 (N_14002,N_11642,N_9833);
and U14003 (N_14003,N_11709,N_11980);
and U14004 (N_14004,N_9603,N_11685);
or U14005 (N_14005,N_11825,N_9998);
xnor U14006 (N_14006,N_12069,N_12486);
xor U14007 (N_14007,N_12380,N_9955);
nor U14008 (N_14008,N_10156,N_10884);
nand U14009 (N_14009,N_10010,N_11553);
nor U14010 (N_14010,N_11401,N_11397);
or U14011 (N_14011,N_11432,N_10624);
nor U14012 (N_14012,N_11796,N_9584);
nand U14013 (N_14013,N_11331,N_12251);
or U14014 (N_14014,N_12483,N_10049);
nand U14015 (N_14015,N_9630,N_10499);
nor U14016 (N_14016,N_10536,N_10152);
xnor U14017 (N_14017,N_12067,N_11817);
or U14018 (N_14018,N_10491,N_10218);
or U14019 (N_14019,N_10028,N_11883);
nand U14020 (N_14020,N_11406,N_11998);
or U14021 (N_14021,N_10761,N_9407);
xor U14022 (N_14022,N_11815,N_11398);
nand U14023 (N_14023,N_11582,N_12462);
nor U14024 (N_14024,N_12284,N_12033);
and U14025 (N_14025,N_11753,N_10643);
xnor U14026 (N_14026,N_10868,N_10173);
nor U14027 (N_14027,N_11233,N_11773);
nand U14028 (N_14028,N_9795,N_10148);
nor U14029 (N_14029,N_12492,N_10826);
nor U14030 (N_14030,N_12099,N_9508);
nand U14031 (N_14031,N_9948,N_9910);
nand U14032 (N_14032,N_11987,N_10159);
or U14033 (N_14033,N_9674,N_11395);
or U14034 (N_14034,N_11168,N_10483);
and U14035 (N_14035,N_11220,N_12244);
nand U14036 (N_14036,N_9686,N_11660);
xnor U14037 (N_14037,N_10631,N_11419);
or U14038 (N_14038,N_9719,N_9921);
or U14039 (N_14039,N_10439,N_12209);
nand U14040 (N_14040,N_10867,N_10358);
nand U14041 (N_14041,N_10219,N_10561);
and U14042 (N_14042,N_11143,N_10006);
or U14043 (N_14043,N_9901,N_11711);
xor U14044 (N_14044,N_10896,N_12481);
nand U14045 (N_14045,N_12091,N_12468);
xnor U14046 (N_14046,N_10014,N_10333);
nand U14047 (N_14047,N_11692,N_9985);
nand U14048 (N_14048,N_11348,N_10648);
xor U14049 (N_14049,N_10875,N_9607);
xor U14050 (N_14050,N_11359,N_10788);
and U14051 (N_14051,N_9889,N_9578);
xnor U14052 (N_14052,N_11988,N_12423);
nand U14053 (N_14053,N_10341,N_11407);
nor U14054 (N_14054,N_9836,N_11053);
and U14055 (N_14055,N_12277,N_9723);
and U14056 (N_14056,N_9650,N_9915);
and U14057 (N_14057,N_11386,N_10629);
xnor U14058 (N_14058,N_12345,N_11423);
and U14059 (N_14059,N_9890,N_11499);
nor U14060 (N_14060,N_11635,N_11866);
or U14061 (N_14061,N_11145,N_11959);
and U14062 (N_14062,N_10157,N_12072);
nand U14063 (N_14063,N_10623,N_10977);
xor U14064 (N_14064,N_11125,N_9967);
xor U14065 (N_14065,N_12208,N_12177);
xnor U14066 (N_14066,N_10833,N_10396);
nor U14067 (N_14067,N_9440,N_10682);
xnor U14068 (N_14068,N_9771,N_9713);
nor U14069 (N_14069,N_12136,N_10312);
nand U14070 (N_14070,N_10480,N_12408);
and U14071 (N_14071,N_11404,N_12096);
and U14072 (N_14072,N_11286,N_9498);
and U14073 (N_14073,N_11008,N_10043);
or U14074 (N_14074,N_12443,N_9992);
xor U14075 (N_14075,N_10455,N_11488);
nor U14076 (N_14076,N_9953,N_10871);
xor U14077 (N_14077,N_11619,N_11250);
and U14078 (N_14078,N_12439,N_12155);
xor U14079 (N_14079,N_11280,N_10002);
xor U14080 (N_14080,N_9733,N_11567);
nor U14081 (N_14081,N_11977,N_11966);
or U14082 (N_14082,N_12112,N_10939);
xnor U14083 (N_14083,N_10392,N_10562);
xnor U14084 (N_14084,N_10730,N_10557);
nor U14085 (N_14085,N_11818,N_9678);
or U14086 (N_14086,N_12112,N_9793);
nor U14087 (N_14087,N_10498,N_12414);
nand U14088 (N_14088,N_11914,N_12270);
or U14089 (N_14089,N_9757,N_11525);
nor U14090 (N_14090,N_10005,N_10389);
nor U14091 (N_14091,N_12346,N_12196);
nor U14092 (N_14092,N_11446,N_12191);
nor U14093 (N_14093,N_9680,N_10675);
or U14094 (N_14094,N_10092,N_10445);
and U14095 (N_14095,N_9770,N_11908);
and U14096 (N_14096,N_9754,N_10012);
xor U14097 (N_14097,N_9890,N_10301);
nor U14098 (N_14098,N_9707,N_12194);
or U14099 (N_14099,N_10713,N_11005);
and U14100 (N_14100,N_11342,N_12001);
or U14101 (N_14101,N_11577,N_12487);
xor U14102 (N_14102,N_11716,N_11627);
or U14103 (N_14103,N_10613,N_11828);
and U14104 (N_14104,N_12235,N_12183);
nand U14105 (N_14105,N_10187,N_12411);
and U14106 (N_14106,N_11049,N_10193);
nor U14107 (N_14107,N_11892,N_9685);
nor U14108 (N_14108,N_11087,N_9432);
xnor U14109 (N_14109,N_11813,N_11105);
or U14110 (N_14110,N_9409,N_12463);
nor U14111 (N_14111,N_12043,N_10359);
or U14112 (N_14112,N_11274,N_11150);
xnor U14113 (N_14113,N_11360,N_10090);
and U14114 (N_14114,N_11660,N_11674);
nor U14115 (N_14115,N_10279,N_10356);
xnor U14116 (N_14116,N_10160,N_10763);
xor U14117 (N_14117,N_11568,N_11445);
nor U14118 (N_14118,N_10633,N_9565);
nand U14119 (N_14119,N_10245,N_10671);
nand U14120 (N_14120,N_9510,N_10292);
and U14121 (N_14121,N_10967,N_10597);
or U14122 (N_14122,N_11769,N_10197);
nor U14123 (N_14123,N_12266,N_9382);
xor U14124 (N_14124,N_9420,N_9478);
xor U14125 (N_14125,N_11186,N_10708);
nor U14126 (N_14126,N_10296,N_9403);
nand U14127 (N_14127,N_10053,N_11966);
xnor U14128 (N_14128,N_10731,N_10511);
nand U14129 (N_14129,N_9459,N_9430);
and U14130 (N_14130,N_10320,N_11909);
and U14131 (N_14131,N_9556,N_10439);
xor U14132 (N_14132,N_10974,N_9979);
nor U14133 (N_14133,N_10850,N_10632);
and U14134 (N_14134,N_10819,N_11402);
nor U14135 (N_14135,N_12112,N_9591);
or U14136 (N_14136,N_11175,N_9526);
and U14137 (N_14137,N_10902,N_9561);
nand U14138 (N_14138,N_10985,N_11708);
and U14139 (N_14139,N_9890,N_11448);
or U14140 (N_14140,N_11625,N_11369);
or U14141 (N_14141,N_9725,N_10331);
xnor U14142 (N_14142,N_11245,N_11022);
nor U14143 (N_14143,N_9841,N_10168);
nor U14144 (N_14144,N_9407,N_12409);
or U14145 (N_14145,N_11647,N_11719);
xnor U14146 (N_14146,N_10091,N_9534);
nor U14147 (N_14147,N_9722,N_10285);
nor U14148 (N_14148,N_10673,N_10962);
or U14149 (N_14149,N_10426,N_10259);
or U14150 (N_14150,N_9639,N_9412);
and U14151 (N_14151,N_9878,N_11145);
and U14152 (N_14152,N_9914,N_11247);
nand U14153 (N_14153,N_11564,N_10180);
or U14154 (N_14154,N_10053,N_11036);
xnor U14155 (N_14155,N_10413,N_9910);
nor U14156 (N_14156,N_11409,N_10552);
nand U14157 (N_14157,N_10412,N_11265);
nor U14158 (N_14158,N_9829,N_11311);
nor U14159 (N_14159,N_9573,N_11423);
nand U14160 (N_14160,N_9408,N_11306);
or U14161 (N_14161,N_10870,N_10097);
and U14162 (N_14162,N_10243,N_11149);
xor U14163 (N_14163,N_10295,N_11343);
xnor U14164 (N_14164,N_11953,N_11531);
or U14165 (N_14165,N_11092,N_11319);
or U14166 (N_14166,N_11234,N_10206);
nor U14167 (N_14167,N_10816,N_10009);
nor U14168 (N_14168,N_10410,N_12181);
and U14169 (N_14169,N_10211,N_11224);
nor U14170 (N_14170,N_11083,N_10460);
nand U14171 (N_14171,N_10920,N_10023);
nor U14172 (N_14172,N_10683,N_10364);
or U14173 (N_14173,N_11082,N_11805);
nand U14174 (N_14174,N_9550,N_10095);
xnor U14175 (N_14175,N_10914,N_9933);
xor U14176 (N_14176,N_10333,N_9471);
nand U14177 (N_14177,N_10163,N_10279);
and U14178 (N_14178,N_10645,N_12024);
xor U14179 (N_14179,N_10839,N_11090);
or U14180 (N_14180,N_10652,N_9521);
nor U14181 (N_14181,N_12116,N_10680);
nor U14182 (N_14182,N_11432,N_11172);
nand U14183 (N_14183,N_11325,N_9934);
nand U14184 (N_14184,N_10337,N_11644);
xor U14185 (N_14185,N_9516,N_11925);
nand U14186 (N_14186,N_9745,N_10147);
xor U14187 (N_14187,N_10240,N_12325);
nor U14188 (N_14188,N_10510,N_9912);
xnor U14189 (N_14189,N_12101,N_10821);
nand U14190 (N_14190,N_12376,N_10870);
nand U14191 (N_14191,N_11306,N_11282);
xnor U14192 (N_14192,N_10175,N_12418);
and U14193 (N_14193,N_10409,N_10385);
nor U14194 (N_14194,N_11795,N_10753);
xnor U14195 (N_14195,N_11358,N_11838);
nand U14196 (N_14196,N_11805,N_12422);
or U14197 (N_14197,N_10084,N_10366);
or U14198 (N_14198,N_11301,N_12437);
and U14199 (N_14199,N_9514,N_11647);
xor U14200 (N_14200,N_10490,N_10586);
and U14201 (N_14201,N_10886,N_9793);
nor U14202 (N_14202,N_9826,N_11953);
nor U14203 (N_14203,N_10421,N_9990);
and U14204 (N_14204,N_10670,N_12216);
and U14205 (N_14205,N_12116,N_10975);
nand U14206 (N_14206,N_11852,N_10370);
nand U14207 (N_14207,N_10296,N_10186);
nor U14208 (N_14208,N_12422,N_11050);
and U14209 (N_14209,N_10356,N_11517);
and U14210 (N_14210,N_9809,N_12214);
nor U14211 (N_14211,N_10119,N_11758);
and U14212 (N_14212,N_10260,N_11382);
and U14213 (N_14213,N_9854,N_11118);
nand U14214 (N_14214,N_11666,N_12094);
xor U14215 (N_14215,N_10109,N_10627);
or U14216 (N_14216,N_11205,N_11305);
and U14217 (N_14217,N_10334,N_11014);
nand U14218 (N_14218,N_11675,N_9514);
nor U14219 (N_14219,N_11798,N_10613);
and U14220 (N_14220,N_12255,N_11890);
and U14221 (N_14221,N_10941,N_10799);
nand U14222 (N_14222,N_10989,N_11641);
nor U14223 (N_14223,N_9462,N_9781);
nor U14224 (N_14224,N_12178,N_12058);
xnor U14225 (N_14225,N_11636,N_12112);
nand U14226 (N_14226,N_12173,N_12383);
xor U14227 (N_14227,N_10713,N_11780);
or U14228 (N_14228,N_12205,N_12238);
or U14229 (N_14229,N_10214,N_11367);
or U14230 (N_14230,N_9949,N_10295);
or U14231 (N_14231,N_11692,N_9923);
and U14232 (N_14232,N_11954,N_11321);
or U14233 (N_14233,N_10887,N_11777);
nor U14234 (N_14234,N_12254,N_10374);
nand U14235 (N_14235,N_12375,N_10960);
nor U14236 (N_14236,N_10496,N_11394);
nor U14237 (N_14237,N_12296,N_10153);
and U14238 (N_14238,N_10792,N_12348);
and U14239 (N_14239,N_9639,N_11383);
and U14240 (N_14240,N_10543,N_12176);
or U14241 (N_14241,N_10294,N_12019);
or U14242 (N_14242,N_10707,N_11171);
or U14243 (N_14243,N_11756,N_10552);
nor U14244 (N_14244,N_12438,N_10815);
and U14245 (N_14245,N_10518,N_10793);
and U14246 (N_14246,N_9521,N_10141);
and U14247 (N_14247,N_9917,N_11719);
nor U14248 (N_14248,N_10516,N_10114);
or U14249 (N_14249,N_10106,N_12434);
or U14250 (N_14250,N_11258,N_11573);
xor U14251 (N_14251,N_11121,N_11632);
and U14252 (N_14252,N_9773,N_11991);
and U14253 (N_14253,N_11057,N_11839);
and U14254 (N_14254,N_9802,N_11931);
xor U14255 (N_14255,N_9833,N_9810);
and U14256 (N_14256,N_11819,N_11301);
nor U14257 (N_14257,N_12024,N_11963);
and U14258 (N_14258,N_11458,N_10643);
and U14259 (N_14259,N_10939,N_11912);
nor U14260 (N_14260,N_12121,N_12311);
or U14261 (N_14261,N_9700,N_11682);
xor U14262 (N_14262,N_9531,N_11318);
xnor U14263 (N_14263,N_9685,N_11070);
and U14264 (N_14264,N_9812,N_10252);
or U14265 (N_14265,N_11561,N_11299);
nor U14266 (N_14266,N_10295,N_10901);
nor U14267 (N_14267,N_11433,N_11790);
nand U14268 (N_14268,N_9716,N_11606);
nand U14269 (N_14269,N_9520,N_10197);
or U14270 (N_14270,N_10513,N_10496);
or U14271 (N_14271,N_11668,N_11486);
nor U14272 (N_14272,N_11498,N_11272);
and U14273 (N_14273,N_10564,N_12320);
and U14274 (N_14274,N_11317,N_9442);
xnor U14275 (N_14275,N_9692,N_10349);
or U14276 (N_14276,N_10265,N_11769);
xor U14277 (N_14277,N_11453,N_9533);
or U14278 (N_14278,N_9940,N_10123);
and U14279 (N_14279,N_9758,N_10387);
or U14280 (N_14280,N_9553,N_10184);
nand U14281 (N_14281,N_11908,N_10920);
or U14282 (N_14282,N_10619,N_11810);
xor U14283 (N_14283,N_9661,N_11203);
and U14284 (N_14284,N_10924,N_11788);
and U14285 (N_14285,N_10938,N_9497);
xor U14286 (N_14286,N_9748,N_12249);
and U14287 (N_14287,N_10599,N_10270);
nand U14288 (N_14288,N_11719,N_10994);
nand U14289 (N_14289,N_11507,N_9468);
xor U14290 (N_14290,N_9510,N_11659);
nand U14291 (N_14291,N_10275,N_11824);
xor U14292 (N_14292,N_11985,N_10114);
nor U14293 (N_14293,N_12189,N_9793);
and U14294 (N_14294,N_10579,N_9502);
and U14295 (N_14295,N_11252,N_11099);
nor U14296 (N_14296,N_10253,N_11785);
or U14297 (N_14297,N_10181,N_9993);
and U14298 (N_14298,N_10601,N_11796);
and U14299 (N_14299,N_12229,N_12462);
or U14300 (N_14300,N_9957,N_10309);
and U14301 (N_14301,N_11913,N_11453);
nand U14302 (N_14302,N_11688,N_9526);
and U14303 (N_14303,N_11231,N_10449);
or U14304 (N_14304,N_11372,N_10653);
and U14305 (N_14305,N_9873,N_12155);
or U14306 (N_14306,N_9489,N_11759);
or U14307 (N_14307,N_11173,N_10790);
nor U14308 (N_14308,N_12027,N_9459);
and U14309 (N_14309,N_10416,N_11286);
or U14310 (N_14310,N_10992,N_9671);
and U14311 (N_14311,N_10402,N_10358);
or U14312 (N_14312,N_10879,N_10265);
nand U14313 (N_14313,N_9772,N_9850);
and U14314 (N_14314,N_11305,N_9696);
and U14315 (N_14315,N_11913,N_11859);
and U14316 (N_14316,N_10347,N_11046);
nor U14317 (N_14317,N_11367,N_11134);
nand U14318 (N_14318,N_10445,N_10883);
or U14319 (N_14319,N_9451,N_12480);
nand U14320 (N_14320,N_9919,N_11864);
xor U14321 (N_14321,N_12151,N_12186);
xnor U14322 (N_14322,N_11174,N_10029);
and U14323 (N_14323,N_10717,N_10197);
nand U14324 (N_14324,N_10943,N_10568);
nor U14325 (N_14325,N_11645,N_9539);
and U14326 (N_14326,N_9469,N_12385);
xnor U14327 (N_14327,N_9845,N_10807);
nor U14328 (N_14328,N_9819,N_10015);
nor U14329 (N_14329,N_12127,N_10411);
and U14330 (N_14330,N_11938,N_10530);
or U14331 (N_14331,N_10629,N_12032);
or U14332 (N_14332,N_11492,N_11888);
nand U14333 (N_14333,N_12261,N_11657);
or U14334 (N_14334,N_9930,N_11009);
nor U14335 (N_14335,N_12436,N_11115);
and U14336 (N_14336,N_9908,N_12321);
nor U14337 (N_14337,N_11102,N_11037);
or U14338 (N_14338,N_12016,N_9623);
xnor U14339 (N_14339,N_11661,N_12000);
nor U14340 (N_14340,N_11163,N_10523);
xor U14341 (N_14341,N_10834,N_11611);
or U14342 (N_14342,N_10927,N_11512);
and U14343 (N_14343,N_11529,N_11618);
nand U14344 (N_14344,N_10378,N_11493);
and U14345 (N_14345,N_11167,N_9981);
nor U14346 (N_14346,N_10913,N_10741);
nor U14347 (N_14347,N_9564,N_9816);
and U14348 (N_14348,N_11342,N_9454);
or U14349 (N_14349,N_11278,N_11442);
nor U14350 (N_14350,N_12317,N_11023);
nand U14351 (N_14351,N_9621,N_11769);
and U14352 (N_14352,N_11127,N_12038);
nor U14353 (N_14353,N_10717,N_9525);
nand U14354 (N_14354,N_12085,N_9689);
and U14355 (N_14355,N_9579,N_9479);
nor U14356 (N_14356,N_11016,N_9616);
nor U14357 (N_14357,N_9391,N_12122);
nor U14358 (N_14358,N_9909,N_10371);
or U14359 (N_14359,N_12278,N_10219);
nor U14360 (N_14360,N_10431,N_12351);
and U14361 (N_14361,N_11069,N_12436);
nand U14362 (N_14362,N_10241,N_11193);
or U14363 (N_14363,N_12306,N_11006);
nor U14364 (N_14364,N_11032,N_11552);
and U14365 (N_14365,N_9513,N_9682);
nand U14366 (N_14366,N_11130,N_9698);
nor U14367 (N_14367,N_11895,N_12067);
xor U14368 (N_14368,N_12017,N_9564);
or U14369 (N_14369,N_9727,N_11957);
nand U14370 (N_14370,N_10886,N_10889);
nand U14371 (N_14371,N_11734,N_11508);
nor U14372 (N_14372,N_12136,N_9781);
nand U14373 (N_14373,N_11916,N_11722);
xnor U14374 (N_14374,N_12058,N_9639);
xor U14375 (N_14375,N_10979,N_10437);
and U14376 (N_14376,N_10599,N_9751);
and U14377 (N_14377,N_9382,N_10532);
nor U14378 (N_14378,N_11395,N_10990);
or U14379 (N_14379,N_11129,N_10709);
and U14380 (N_14380,N_11868,N_9523);
xor U14381 (N_14381,N_9850,N_10942);
nor U14382 (N_14382,N_10106,N_10416);
nand U14383 (N_14383,N_11443,N_10778);
and U14384 (N_14384,N_12017,N_9548);
nand U14385 (N_14385,N_10663,N_11692);
nand U14386 (N_14386,N_11618,N_10472);
nor U14387 (N_14387,N_11149,N_10893);
nand U14388 (N_14388,N_11086,N_9738);
xor U14389 (N_14389,N_10832,N_11651);
or U14390 (N_14390,N_11363,N_11241);
or U14391 (N_14391,N_10454,N_9657);
or U14392 (N_14392,N_11161,N_11780);
nor U14393 (N_14393,N_10188,N_10918);
nand U14394 (N_14394,N_12043,N_9439);
nor U14395 (N_14395,N_9971,N_10230);
or U14396 (N_14396,N_10739,N_10424);
nand U14397 (N_14397,N_11695,N_9901);
nand U14398 (N_14398,N_11174,N_10442);
and U14399 (N_14399,N_11374,N_10648);
and U14400 (N_14400,N_11434,N_9961);
and U14401 (N_14401,N_10667,N_11250);
and U14402 (N_14402,N_11785,N_12358);
or U14403 (N_14403,N_9907,N_11422);
nor U14404 (N_14404,N_10132,N_11050);
nand U14405 (N_14405,N_9762,N_11875);
and U14406 (N_14406,N_11934,N_11359);
xor U14407 (N_14407,N_9794,N_9805);
and U14408 (N_14408,N_11419,N_10501);
xor U14409 (N_14409,N_10350,N_11475);
nand U14410 (N_14410,N_10980,N_11173);
and U14411 (N_14411,N_11637,N_12408);
nor U14412 (N_14412,N_12023,N_9733);
or U14413 (N_14413,N_11420,N_10250);
or U14414 (N_14414,N_11653,N_11730);
nand U14415 (N_14415,N_12373,N_10408);
xnor U14416 (N_14416,N_10420,N_12484);
or U14417 (N_14417,N_12081,N_11918);
xnor U14418 (N_14418,N_11313,N_12382);
xor U14419 (N_14419,N_9702,N_10732);
or U14420 (N_14420,N_10624,N_9444);
xnor U14421 (N_14421,N_9477,N_9709);
xor U14422 (N_14422,N_10746,N_9695);
and U14423 (N_14423,N_10174,N_10425);
or U14424 (N_14424,N_10247,N_11205);
xnor U14425 (N_14425,N_9537,N_10649);
xnor U14426 (N_14426,N_10818,N_11495);
and U14427 (N_14427,N_10530,N_11766);
nand U14428 (N_14428,N_11542,N_11297);
and U14429 (N_14429,N_9707,N_11785);
nor U14430 (N_14430,N_12360,N_9385);
and U14431 (N_14431,N_9463,N_10098);
or U14432 (N_14432,N_11058,N_9851);
nand U14433 (N_14433,N_12221,N_10314);
xor U14434 (N_14434,N_11704,N_12425);
nand U14435 (N_14435,N_11026,N_10951);
nor U14436 (N_14436,N_10979,N_9747);
nand U14437 (N_14437,N_10605,N_10515);
or U14438 (N_14438,N_11740,N_10926);
or U14439 (N_14439,N_9902,N_9811);
or U14440 (N_14440,N_12052,N_12194);
xnor U14441 (N_14441,N_11301,N_10762);
nor U14442 (N_14442,N_11688,N_10657);
xnor U14443 (N_14443,N_11048,N_11399);
nand U14444 (N_14444,N_9737,N_12173);
xor U14445 (N_14445,N_11223,N_10209);
nand U14446 (N_14446,N_9950,N_11101);
xor U14447 (N_14447,N_11535,N_10881);
or U14448 (N_14448,N_10025,N_10428);
nor U14449 (N_14449,N_11596,N_9433);
nand U14450 (N_14450,N_10562,N_11766);
nor U14451 (N_14451,N_10003,N_11553);
xor U14452 (N_14452,N_10283,N_11792);
or U14453 (N_14453,N_9915,N_10468);
or U14454 (N_14454,N_10324,N_11127);
or U14455 (N_14455,N_10474,N_12213);
nand U14456 (N_14456,N_11557,N_10704);
nor U14457 (N_14457,N_10534,N_11431);
or U14458 (N_14458,N_10044,N_9755);
and U14459 (N_14459,N_9507,N_9998);
and U14460 (N_14460,N_9799,N_10180);
nand U14461 (N_14461,N_10316,N_9778);
xor U14462 (N_14462,N_11240,N_11462);
and U14463 (N_14463,N_11510,N_10329);
xor U14464 (N_14464,N_10086,N_11713);
or U14465 (N_14465,N_10476,N_12026);
nor U14466 (N_14466,N_11643,N_10752);
xnor U14467 (N_14467,N_11489,N_11281);
nor U14468 (N_14468,N_11537,N_11445);
xnor U14469 (N_14469,N_11028,N_12495);
nor U14470 (N_14470,N_11443,N_10887);
nand U14471 (N_14471,N_11942,N_12138);
xnor U14472 (N_14472,N_11155,N_9378);
nor U14473 (N_14473,N_12441,N_9859);
or U14474 (N_14474,N_10273,N_10129);
xor U14475 (N_14475,N_10085,N_11248);
nor U14476 (N_14476,N_10416,N_11389);
or U14477 (N_14477,N_11370,N_9880);
or U14478 (N_14478,N_10436,N_9919);
or U14479 (N_14479,N_9901,N_10101);
xnor U14480 (N_14480,N_11959,N_11218);
xor U14481 (N_14481,N_9907,N_12146);
xor U14482 (N_14482,N_9472,N_11777);
nor U14483 (N_14483,N_10907,N_11529);
xor U14484 (N_14484,N_11213,N_11796);
nand U14485 (N_14485,N_12136,N_11770);
and U14486 (N_14486,N_10863,N_10355);
and U14487 (N_14487,N_10360,N_10668);
or U14488 (N_14488,N_10365,N_11351);
nor U14489 (N_14489,N_9616,N_11696);
xnor U14490 (N_14490,N_12083,N_11599);
nor U14491 (N_14491,N_12132,N_12485);
xnor U14492 (N_14492,N_9802,N_9650);
nand U14493 (N_14493,N_11541,N_11543);
xor U14494 (N_14494,N_9576,N_10058);
xor U14495 (N_14495,N_12074,N_9638);
or U14496 (N_14496,N_9427,N_10250);
or U14497 (N_14497,N_12248,N_10907);
nor U14498 (N_14498,N_10163,N_10017);
and U14499 (N_14499,N_10382,N_9513);
or U14500 (N_14500,N_12091,N_11283);
nand U14501 (N_14501,N_10289,N_12293);
or U14502 (N_14502,N_10863,N_11543);
and U14503 (N_14503,N_10948,N_9526);
or U14504 (N_14504,N_10780,N_10845);
xor U14505 (N_14505,N_10554,N_12245);
or U14506 (N_14506,N_12421,N_11083);
or U14507 (N_14507,N_10651,N_11914);
or U14508 (N_14508,N_10448,N_10993);
and U14509 (N_14509,N_9635,N_11016);
nand U14510 (N_14510,N_10975,N_10300);
and U14511 (N_14511,N_12164,N_11456);
or U14512 (N_14512,N_11549,N_9588);
xor U14513 (N_14513,N_11341,N_9684);
xor U14514 (N_14514,N_11276,N_12105);
xor U14515 (N_14515,N_10960,N_11713);
and U14516 (N_14516,N_9894,N_10471);
and U14517 (N_14517,N_9743,N_11006);
xnor U14518 (N_14518,N_11503,N_10129);
xor U14519 (N_14519,N_10482,N_9535);
and U14520 (N_14520,N_9664,N_10091);
nor U14521 (N_14521,N_11657,N_12338);
or U14522 (N_14522,N_10968,N_10817);
xnor U14523 (N_14523,N_10004,N_9453);
and U14524 (N_14524,N_10266,N_10093);
xor U14525 (N_14525,N_11701,N_11293);
and U14526 (N_14526,N_11755,N_11002);
nor U14527 (N_14527,N_10182,N_11658);
nand U14528 (N_14528,N_10246,N_11024);
and U14529 (N_14529,N_11641,N_9475);
xor U14530 (N_14530,N_12109,N_11606);
nand U14531 (N_14531,N_10023,N_10786);
and U14532 (N_14532,N_12055,N_10309);
nor U14533 (N_14533,N_10460,N_10283);
or U14534 (N_14534,N_9413,N_11865);
nand U14535 (N_14535,N_10329,N_11369);
xor U14536 (N_14536,N_9385,N_11553);
xor U14537 (N_14537,N_11787,N_10579);
nor U14538 (N_14538,N_10071,N_11952);
xor U14539 (N_14539,N_10401,N_12437);
xnor U14540 (N_14540,N_11175,N_10019);
nand U14541 (N_14541,N_11755,N_12415);
or U14542 (N_14542,N_9723,N_10004);
nor U14543 (N_14543,N_12066,N_12221);
xnor U14544 (N_14544,N_11885,N_11961);
nor U14545 (N_14545,N_11737,N_9989);
xnor U14546 (N_14546,N_10371,N_12335);
and U14547 (N_14547,N_11156,N_11775);
xnor U14548 (N_14548,N_9434,N_12206);
and U14549 (N_14549,N_12470,N_11107);
nand U14550 (N_14550,N_12100,N_10094);
and U14551 (N_14551,N_12019,N_9454);
and U14552 (N_14552,N_11511,N_10886);
and U14553 (N_14553,N_9805,N_12449);
xor U14554 (N_14554,N_10364,N_10075);
xnor U14555 (N_14555,N_12253,N_11656);
nand U14556 (N_14556,N_12239,N_11510);
xnor U14557 (N_14557,N_11190,N_11109);
nand U14558 (N_14558,N_9676,N_9440);
or U14559 (N_14559,N_9782,N_11399);
xor U14560 (N_14560,N_12318,N_11607);
nor U14561 (N_14561,N_11849,N_11269);
and U14562 (N_14562,N_10366,N_9386);
and U14563 (N_14563,N_9948,N_9878);
and U14564 (N_14564,N_10854,N_10703);
nand U14565 (N_14565,N_11494,N_9474);
xnor U14566 (N_14566,N_12019,N_10614);
nand U14567 (N_14567,N_10446,N_9809);
and U14568 (N_14568,N_12153,N_9926);
nor U14569 (N_14569,N_9387,N_11462);
or U14570 (N_14570,N_10929,N_9787);
xor U14571 (N_14571,N_9614,N_9975);
or U14572 (N_14572,N_12061,N_11308);
nand U14573 (N_14573,N_12066,N_9732);
nand U14574 (N_14574,N_11706,N_11671);
nand U14575 (N_14575,N_12083,N_11034);
and U14576 (N_14576,N_10785,N_10543);
nand U14577 (N_14577,N_11629,N_11998);
nor U14578 (N_14578,N_12439,N_12324);
nor U14579 (N_14579,N_9923,N_11172);
nor U14580 (N_14580,N_11923,N_11644);
or U14581 (N_14581,N_10486,N_11779);
and U14582 (N_14582,N_12334,N_10725);
or U14583 (N_14583,N_11853,N_9690);
and U14584 (N_14584,N_10996,N_11330);
xnor U14585 (N_14585,N_12035,N_11669);
xnor U14586 (N_14586,N_9518,N_11714);
nor U14587 (N_14587,N_10200,N_12491);
or U14588 (N_14588,N_9571,N_10406);
nand U14589 (N_14589,N_9644,N_12159);
or U14590 (N_14590,N_11192,N_12179);
nor U14591 (N_14591,N_10257,N_11064);
or U14592 (N_14592,N_9440,N_10039);
nand U14593 (N_14593,N_9839,N_10614);
nor U14594 (N_14594,N_10572,N_9713);
xnor U14595 (N_14595,N_11309,N_10901);
and U14596 (N_14596,N_10117,N_10552);
and U14597 (N_14597,N_9962,N_9879);
and U14598 (N_14598,N_11120,N_12237);
and U14599 (N_14599,N_11566,N_11440);
and U14600 (N_14600,N_10203,N_12029);
nand U14601 (N_14601,N_11571,N_11047);
nand U14602 (N_14602,N_10787,N_11297);
xnor U14603 (N_14603,N_11859,N_11862);
or U14604 (N_14604,N_11523,N_10270);
xor U14605 (N_14605,N_11528,N_11742);
or U14606 (N_14606,N_11246,N_12360);
and U14607 (N_14607,N_11331,N_12340);
or U14608 (N_14608,N_10849,N_12096);
and U14609 (N_14609,N_10069,N_11880);
nor U14610 (N_14610,N_9707,N_10864);
or U14611 (N_14611,N_12387,N_10623);
nand U14612 (N_14612,N_9903,N_12221);
nor U14613 (N_14613,N_11603,N_10003);
nand U14614 (N_14614,N_11276,N_10504);
or U14615 (N_14615,N_12107,N_12355);
nand U14616 (N_14616,N_11670,N_10555);
or U14617 (N_14617,N_10947,N_12365);
nor U14618 (N_14618,N_10549,N_12300);
or U14619 (N_14619,N_9407,N_9971);
nand U14620 (N_14620,N_11031,N_9614);
nor U14621 (N_14621,N_11258,N_11694);
xnor U14622 (N_14622,N_11424,N_11279);
and U14623 (N_14623,N_10304,N_10734);
nand U14624 (N_14624,N_10750,N_11458);
or U14625 (N_14625,N_11928,N_9687);
nand U14626 (N_14626,N_9422,N_10143);
nor U14627 (N_14627,N_11148,N_11815);
or U14628 (N_14628,N_11897,N_11439);
and U14629 (N_14629,N_12322,N_9639);
nor U14630 (N_14630,N_11947,N_10270);
xor U14631 (N_14631,N_10256,N_11971);
nand U14632 (N_14632,N_10320,N_10607);
nor U14633 (N_14633,N_10825,N_11386);
xor U14634 (N_14634,N_12137,N_10378);
or U14635 (N_14635,N_11380,N_11283);
or U14636 (N_14636,N_9929,N_12067);
xnor U14637 (N_14637,N_11129,N_10793);
xnor U14638 (N_14638,N_9659,N_11524);
or U14639 (N_14639,N_10400,N_11234);
nand U14640 (N_14640,N_11839,N_9400);
nand U14641 (N_14641,N_11069,N_11886);
and U14642 (N_14642,N_11666,N_11235);
xor U14643 (N_14643,N_11879,N_10951);
or U14644 (N_14644,N_9611,N_11158);
and U14645 (N_14645,N_11546,N_9540);
nand U14646 (N_14646,N_9574,N_11928);
xnor U14647 (N_14647,N_11428,N_11339);
nand U14648 (N_14648,N_9687,N_12270);
nor U14649 (N_14649,N_11579,N_12016);
xor U14650 (N_14650,N_11269,N_10847);
nand U14651 (N_14651,N_11620,N_10977);
nand U14652 (N_14652,N_10797,N_10021);
nor U14653 (N_14653,N_10452,N_10727);
and U14654 (N_14654,N_10723,N_10730);
or U14655 (N_14655,N_10021,N_9895);
or U14656 (N_14656,N_10524,N_11577);
and U14657 (N_14657,N_9880,N_9650);
or U14658 (N_14658,N_10141,N_9676);
and U14659 (N_14659,N_9560,N_9744);
xor U14660 (N_14660,N_12100,N_11594);
nand U14661 (N_14661,N_11749,N_9735);
or U14662 (N_14662,N_10962,N_9901);
nor U14663 (N_14663,N_11162,N_11378);
and U14664 (N_14664,N_12469,N_12338);
or U14665 (N_14665,N_10734,N_11859);
xor U14666 (N_14666,N_12009,N_9882);
nor U14667 (N_14667,N_12355,N_9928);
or U14668 (N_14668,N_12021,N_11444);
xor U14669 (N_14669,N_11667,N_12145);
nor U14670 (N_14670,N_11002,N_9785);
or U14671 (N_14671,N_9795,N_10767);
nor U14672 (N_14672,N_12396,N_11189);
nand U14673 (N_14673,N_9875,N_10236);
or U14674 (N_14674,N_11630,N_10980);
nor U14675 (N_14675,N_11442,N_11860);
nand U14676 (N_14676,N_10787,N_9483);
or U14677 (N_14677,N_9833,N_9698);
and U14678 (N_14678,N_12373,N_10034);
nor U14679 (N_14679,N_10213,N_11584);
nor U14680 (N_14680,N_9489,N_9474);
or U14681 (N_14681,N_9842,N_12288);
nand U14682 (N_14682,N_11358,N_10590);
nor U14683 (N_14683,N_9943,N_10769);
nand U14684 (N_14684,N_10218,N_12189);
or U14685 (N_14685,N_11318,N_9430);
nand U14686 (N_14686,N_9909,N_10168);
nor U14687 (N_14687,N_9725,N_9917);
nand U14688 (N_14688,N_10111,N_10080);
nor U14689 (N_14689,N_11064,N_11180);
and U14690 (N_14690,N_11667,N_9992);
or U14691 (N_14691,N_11578,N_11542);
nor U14692 (N_14692,N_11435,N_10602);
xnor U14693 (N_14693,N_11589,N_9376);
or U14694 (N_14694,N_9800,N_12191);
xor U14695 (N_14695,N_11310,N_10712);
nor U14696 (N_14696,N_11436,N_10399);
and U14697 (N_14697,N_9681,N_10818);
or U14698 (N_14698,N_11805,N_9506);
xor U14699 (N_14699,N_11739,N_12426);
and U14700 (N_14700,N_10923,N_12220);
nor U14701 (N_14701,N_12363,N_10113);
nor U14702 (N_14702,N_10559,N_9608);
and U14703 (N_14703,N_11747,N_10821);
nand U14704 (N_14704,N_10275,N_10543);
and U14705 (N_14705,N_11054,N_9888);
nor U14706 (N_14706,N_10660,N_11244);
xor U14707 (N_14707,N_10684,N_9772);
xor U14708 (N_14708,N_10310,N_12145);
and U14709 (N_14709,N_9734,N_11851);
nor U14710 (N_14710,N_11847,N_12355);
or U14711 (N_14711,N_9518,N_11497);
nor U14712 (N_14712,N_11983,N_11907);
xor U14713 (N_14713,N_9659,N_9993);
xnor U14714 (N_14714,N_10003,N_11180);
nor U14715 (N_14715,N_10521,N_11658);
or U14716 (N_14716,N_10347,N_11293);
or U14717 (N_14717,N_11171,N_9839);
and U14718 (N_14718,N_12364,N_10819);
and U14719 (N_14719,N_10459,N_11628);
or U14720 (N_14720,N_9981,N_10191);
nand U14721 (N_14721,N_9735,N_9386);
xor U14722 (N_14722,N_11868,N_10707);
nor U14723 (N_14723,N_11779,N_10051);
nand U14724 (N_14724,N_11340,N_10169);
xor U14725 (N_14725,N_10292,N_10748);
or U14726 (N_14726,N_10625,N_10394);
nand U14727 (N_14727,N_10069,N_10329);
nor U14728 (N_14728,N_10430,N_11666);
xnor U14729 (N_14729,N_12001,N_12323);
or U14730 (N_14730,N_10294,N_9904);
nand U14731 (N_14731,N_10452,N_12064);
and U14732 (N_14732,N_12296,N_11946);
xnor U14733 (N_14733,N_10676,N_11741);
nand U14734 (N_14734,N_11941,N_12106);
or U14735 (N_14735,N_10412,N_9748);
xor U14736 (N_14736,N_12128,N_12295);
or U14737 (N_14737,N_9643,N_10497);
xor U14738 (N_14738,N_11908,N_11518);
nor U14739 (N_14739,N_10679,N_11315);
xnor U14740 (N_14740,N_11674,N_10779);
nand U14741 (N_14741,N_10334,N_9442);
nand U14742 (N_14742,N_10359,N_11191);
nand U14743 (N_14743,N_11825,N_11743);
and U14744 (N_14744,N_10337,N_10845);
nand U14745 (N_14745,N_10346,N_12162);
nand U14746 (N_14746,N_11237,N_9902);
or U14747 (N_14747,N_9812,N_12219);
or U14748 (N_14748,N_10873,N_11202);
nor U14749 (N_14749,N_9853,N_10131);
nand U14750 (N_14750,N_9855,N_9534);
nor U14751 (N_14751,N_12285,N_10043);
nor U14752 (N_14752,N_10853,N_12178);
xor U14753 (N_14753,N_11096,N_11178);
or U14754 (N_14754,N_10340,N_11341);
and U14755 (N_14755,N_11171,N_9919);
or U14756 (N_14756,N_12241,N_9623);
nand U14757 (N_14757,N_11449,N_10706);
or U14758 (N_14758,N_9658,N_12336);
xor U14759 (N_14759,N_10352,N_10125);
nor U14760 (N_14760,N_10214,N_10141);
nand U14761 (N_14761,N_9551,N_9661);
and U14762 (N_14762,N_11077,N_11537);
xor U14763 (N_14763,N_9696,N_10139);
and U14764 (N_14764,N_12212,N_10208);
and U14765 (N_14765,N_12398,N_11201);
nor U14766 (N_14766,N_10158,N_10933);
and U14767 (N_14767,N_11941,N_11721);
or U14768 (N_14768,N_11697,N_10756);
xnor U14769 (N_14769,N_12069,N_9391);
nand U14770 (N_14770,N_12331,N_10694);
and U14771 (N_14771,N_12447,N_9811);
nor U14772 (N_14772,N_11881,N_10866);
nand U14773 (N_14773,N_11838,N_9795);
xnor U14774 (N_14774,N_11711,N_11255);
and U14775 (N_14775,N_10472,N_12413);
nor U14776 (N_14776,N_10255,N_10677);
or U14777 (N_14777,N_12401,N_12058);
or U14778 (N_14778,N_10955,N_12094);
nand U14779 (N_14779,N_10866,N_10551);
nor U14780 (N_14780,N_10652,N_10326);
and U14781 (N_14781,N_12474,N_12316);
nand U14782 (N_14782,N_9678,N_10820);
and U14783 (N_14783,N_10547,N_10625);
nor U14784 (N_14784,N_11683,N_9580);
or U14785 (N_14785,N_10424,N_10026);
nand U14786 (N_14786,N_12049,N_12091);
nand U14787 (N_14787,N_10811,N_11346);
xnor U14788 (N_14788,N_12040,N_9894);
xnor U14789 (N_14789,N_11080,N_11525);
xor U14790 (N_14790,N_11944,N_9614);
xor U14791 (N_14791,N_12469,N_10352);
or U14792 (N_14792,N_12280,N_10283);
or U14793 (N_14793,N_12079,N_12252);
nor U14794 (N_14794,N_10933,N_10277);
and U14795 (N_14795,N_10583,N_10902);
nor U14796 (N_14796,N_9425,N_9741);
nand U14797 (N_14797,N_9674,N_11643);
xor U14798 (N_14798,N_11137,N_10977);
or U14799 (N_14799,N_11187,N_9413);
nand U14800 (N_14800,N_11622,N_11974);
nand U14801 (N_14801,N_10736,N_10643);
or U14802 (N_14802,N_12380,N_11683);
nand U14803 (N_14803,N_9832,N_10575);
and U14804 (N_14804,N_10885,N_9956);
and U14805 (N_14805,N_11431,N_11364);
or U14806 (N_14806,N_10515,N_12070);
nand U14807 (N_14807,N_11830,N_11019);
nor U14808 (N_14808,N_10711,N_10749);
nand U14809 (N_14809,N_11083,N_11036);
nor U14810 (N_14810,N_11253,N_9957);
xor U14811 (N_14811,N_10913,N_9703);
or U14812 (N_14812,N_9635,N_10577);
or U14813 (N_14813,N_12400,N_10661);
nor U14814 (N_14814,N_10291,N_11142);
nor U14815 (N_14815,N_9822,N_11175);
or U14816 (N_14816,N_10427,N_11992);
and U14817 (N_14817,N_9847,N_12254);
nand U14818 (N_14818,N_11459,N_9849);
or U14819 (N_14819,N_9583,N_11751);
or U14820 (N_14820,N_10019,N_10311);
nand U14821 (N_14821,N_9921,N_12375);
nor U14822 (N_14822,N_11346,N_12007);
nand U14823 (N_14823,N_11855,N_10524);
xnor U14824 (N_14824,N_10456,N_11614);
xor U14825 (N_14825,N_9808,N_11538);
nor U14826 (N_14826,N_11769,N_12232);
or U14827 (N_14827,N_9461,N_11556);
nand U14828 (N_14828,N_11532,N_11244);
and U14829 (N_14829,N_10990,N_11346);
nand U14830 (N_14830,N_10635,N_11472);
nor U14831 (N_14831,N_10761,N_11360);
or U14832 (N_14832,N_9916,N_12112);
xor U14833 (N_14833,N_12122,N_12292);
and U14834 (N_14834,N_9956,N_11441);
and U14835 (N_14835,N_11040,N_11636);
nor U14836 (N_14836,N_11975,N_12002);
and U14837 (N_14837,N_9701,N_12050);
xor U14838 (N_14838,N_12105,N_11720);
nor U14839 (N_14839,N_9916,N_10935);
nor U14840 (N_14840,N_11126,N_11941);
nand U14841 (N_14841,N_12199,N_11467);
or U14842 (N_14842,N_11677,N_11547);
xnor U14843 (N_14843,N_10096,N_11631);
or U14844 (N_14844,N_11865,N_11649);
nor U14845 (N_14845,N_10550,N_9825);
xor U14846 (N_14846,N_12151,N_10128);
and U14847 (N_14847,N_9985,N_10575);
nor U14848 (N_14848,N_10096,N_9579);
xor U14849 (N_14849,N_10966,N_11561);
nor U14850 (N_14850,N_11873,N_9939);
or U14851 (N_14851,N_10778,N_11899);
and U14852 (N_14852,N_12338,N_10481);
xnor U14853 (N_14853,N_11627,N_12308);
nor U14854 (N_14854,N_9732,N_10703);
nor U14855 (N_14855,N_11597,N_10542);
xnor U14856 (N_14856,N_11995,N_11066);
xor U14857 (N_14857,N_12423,N_10650);
nor U14858 (N_14858,N_11379,N_11503);
and U14859 (N_14859,N_10581,N_12494);
or U14860 (N_14860,N_9380,N_10055);
nor U14861 (N_14861,N_10053,N_11069);
and U14862 (N_14862,N_9867,N_12340);
or U14863 (N_14863,N_11754,N_9769);
and U14864 (N_14864,N_11792,N_10423);
nor U14865 (N_14865,N_10063,N_12420);
and U14866 (N_14866,N_10506,N_10747);
or U14867 (N_14867,N_10262,N_10638);
nand U14868 (N_14868,N_12392,N_10260);
nand U14869 (N_14869,N_11844,N_11407);
or U14870 (N_14870,N_11279,N_11923);
or U14871 (N_14871,N_10470,N_11301);
or U14872 (N_14872,N_11250,N_10973);
and U14873 (N_14873,N_10699,N_11500);
xor U14874 (N_14874,N_10966,N_10909);
xor U14875 (N_14875,N_10075,N_11568);
or U14876 (N_14876,N_10777,N_9588);
nor U14877 (N_14877,N_11327,N_9900);
and U14878 (N_14878,N_9698,N_10261);
or U14879 (N_14879,N_12082,N_11708);
nand U14880 (N_14880,N_9699,N_9695);
nand U14881 (N_14881,N_12217,N_10658);
xnor U14882 (N_14882,N_11590,N_11572);
and U14883 (N_14883,N_9816,N_9837);
xnor U14884 (N_14884,N_9751,N_9741);
xor U14885 (N_14885,N_10213,N_11788);
nand U14886 (N_14886,N_10832,N_11649);
and U14887 (N_14887,N_11021,N_10750);
nor U14888 (N_14888,N_10241,N_11929);
or U14889 (N_14889,N_12457,N_11566);
xor U14890 (N_14890,N_11847,N_11074);
or U14891 (N_14891,N_12293,N_11017);
nor U14892 (N_14892,N_9654,N_10212);
or U14893 (N_14893,N_12449,N_11551);
or U14894 (N_14894,N_12163,N_10711);
nor U14895 (N_14895,N_10784,N_9804);
or U14896 (N_14896,N_12287,N_11729);
nor U14897 (N_14897,N_11340,N_11687);
nor U14898 (N_14898,N_12389,N_9877);
nand U14899 (N_14899,N_11189,N_9736);
nor U14900 (N_14900,N_9643,N_9947);
nand U14901 (N_14901,N_10296,N_12163);
xnor U14902 (N_14902,N_10949,N_9861);
xnor U14903 (N_14903,N_10432,N_10019);
or U14904 (N_14904,N_11073,N_9528);
and U14905 (N_14905,N_11090,N_9628);
xnor U14906 (N_14906,N_11034,N_12104);
nand U14907 (N_14907,N_9680,N_9931);
and U14908 (N_14908,N_10022,N_9864);
and U14909 (N_14909,N_11492,N_11335);
or U14910 (N_14910,N_12367,N_10765);
nor U14911 (N_14911,N_12471,N_12322);
nand U14912 (N_14912,N_12447,N_10623);
or U14913 (N_14913,N_10180,N_10160);
or U14914 (N_14914,N_10375,N_12367);
nor U14915 (N_14915,N_9569,N_12060);
or U14916 (N_14916,N_10706,N_12219);
xor U14917 (N_14917,N_10663,N_10590);
nand U14918 (N_14918,N_11054,N_12428);
and U14919 (N_14919,N_11294,N_11044);
nand U14920 (N_14920,N_9387,N_10482);
nor U14921 (N_14921,N_11133,N_12329);
and U14922 (N_14922,N_11734,N_11421);
nor U14923 (N_14923,N_11304,N_9402);
and U14924 (N_14924,N_12091,N_12260);
nor U14925 (N_14925,N_11626,N_11635);
or U14926 (N_14926,N_10898,N_11983);
xor U14927 (N_14927,N_9551,N_9424);
nand U14928 (N_14928,N_10523,N_11515);
or U14929 (N_14929,N_11256,N_11727);
and U14930 (N_14930,N_10581,N_10220);
nor U14931 (N_14931,N_10766,N_10961);
or U14932 (N_14932,N_11631,N_11536);
or U14933 (N_14933,N_10045,N_10243);
or U14934 (N_14934,N_10547,N_12091);
nand U14935 (N_14935,N_10402,N_11264);
or U14936 (N_14936,N_10897,N_11673);
or U14937 (N_14937,N_11640,N_10509);
nand U14938 (N_14938,N_11894,N_9672);
xor U14939 (N_14939,N_11994,N_10946);
and U14940 (N_14940,N_11930,N_11555);
nor U14941 (N_14941,N_11895,N_10967);
xnor U14942 (N_14942,N_10515,N_10010);
xor U14943 (N_14943,N_10056,N_10936);
xor U14944 (N_14944,N_11261,N_10106);
xnor U14945 (N_14945,N_12008,N_9992);
or U14946 (N_14946,N_10493,N_10443);
nor U14947 (N_14947,N_10443,N_11866);
xnor U14948 (N_14948,N_12356,N_9496);
nor U14949 (N_14949,N_11274,N_11077);
nand U14950 (N_14950,N_11037,N_10000);
and U14951 (N_14951,N_9702,N_9658);
and U14952 (N_14952,N_10732,N_10324);
and U14953 (N_14953,N_9983,N_11308);
and U14954 (N_14954,N_10113,N_11007);
and U14955 (N_14955,N_11768,N_12389);
and U14956 (N_14956,N_10100,N_9827);
xor U14957 (N_14957,N_9437,N_10491);
or U14958 (N_14958,N_10504,N_10269);
xor U14959 (N_14959,N_10157,N_9631);
xor U14960 (N_14960,N_11727,N_10597);
nand U14961 (N_14961,N_9886,N_9864);
or U14962 (N_14962,N_12217,N_10040);
nand U14963 (N_14963,N_11053,N_11431);
nand U14964 (N_14964,N_10681,N_11465);
xor U14965 (N_14965,N_11225,N_11426);
nand U14966 (N_14966,N_9817,N_11236);
nand U14967 (N_14967,N_10490,N_10913);
and U14968 (N_14968,N_12386,N_10574);
or U14969 (N_14969,N_9396,N_10077);
and U14970 (N_14970,N_11983,N_9502);
or U14971 (N_14971,N_10013,N_12283);
xor U14972 (N_14972,N_9515,N_11215);
xor U14973 (N_14973,N_11257,N_9800);
nor U14974 (N_14974,N_9384,N_10750);
nor U14975 (N_14975,N_11162,N_12066);
nor U14976 (N_14976,N_11364,N_10240);
xnor U14977 (N_14977,N_11715,N_11726);
or U14978 (N_14978,N_11466,N_11075);
nand U14979 (N_14979,N_11222,N_12433);
nand U14980 (N_14980,N_12137,N_9698);
and U14981 (N_14981,N_9760,N_11763);
xor U14982 (N_14982,N_12495,N_10655);
nand U14983 (N_14983,N_11814,N_9478);
nor U14984 (N_14984,N_12447,N_10247);
xnor U14985 (N_14985,N_11300,N_10490);
nand U14986 (N_14986,N_12015,N_10169);
nand U14987 (N_14987,N_10345,N_11532);
xor U14988 (N_14988,N_10619,N_11543);
and U14989 (N_14989,N_9536,N_9785);
and U14990 (N_14990,N_10311,N_12488);
or U14991 (N_14991,N_12265,N_12269);
nor U14992 (N_14992,N_9950,N_10393);
nor U14993 (N_14993,N_9951,N_10449);
xor U14994 (N_14994,N_12426,N_11192);
nand U14995 (N_14995,N_10570,N_9855);
nor U14996 (N_14996,N_9598,N_10433);
and U14997 (N_14997,N_10999,N_10953);
or U14998 (N_14998,N_9646,N_10497);
nand U14999 (N_14999,N_10361,N_11756);
and U15000 (N_15000,N_12293,N_11896);
or U15001 (N_15001,N_12206,N_11901);
xor U15002 (N_15002,N_10136,N_11701);
or U15003 (N_15003,N_10808,N_10841);
or U15004 (N_15004,N_11553,N_9702);
and U15005 (N_15005,N_11729,N_9518);
or U15006 (N_15006,N_9749,N_9861);
or U15007 (N_15007,N_10744,N_10880);
nor U15008 (N_15008,N_10894,N_9409);
xnor U15009 (N_15009,N_9645,N_9694);
or U15010 (N_15010,N_11787,N_10984);
and U15011 (N_15011,N_9712,N_11402);
nor U15012 (N_15012,N_11157,N_10823);
or U15013 (N_15013,N_12182,N_10595);
xor U15014 (N_15014,N_10894,N_11780);
nand U15015 (N_15015,N_10042,N_10082);
or U15016 (N_15016,N_11270,N_11718);
and U15017 (N_15017,N_10925,N_11895);
or U15018 (N_15018,N_10029,N_10676);
xnor U15019 (N_15019,N_10634,N_9755);
nand U15020 (N_15020,N_9706,N_9666);
nand U15021 (N_15021,N_10522,N_9473);
and U15022 (N_15022,N_10884,N_11607);
and U15023 (N_15023,N_11655,N_9984);
or U15024 (N_15024,N_10750,N_12188);
or U15025 (N_15025,N_9736,N_11085);
xor U15026 (N_15026,N_11700,N_11919);
and U15027 (N_15027,N_10118,N_10538);
xnor U15028 (N_15028,N_9823,N_11675);
nand U15029 (N_15029,N_12399,N_10373);
and U15030 (N_15030,N_12041,N_10490);
or U15031 (N_15031,N_9906,N_10295);
xnor U15032 (N_15032,N_10181,N_11981);
and U15033 (N_15033,N_11951,N_10615);
or U15034 (N_15034,N_10904,N_10987);
nand U15035 (N_15035,N_11981,N_9760);
nand U15036 (N_15036,N_11511,N_11934);
nor U15037 (N_15037,N_12153,N_9404);
or U15038 (N_15038,N_10285,N_11729);
xnor U15039 (N_15039,N_11717,N_10848);
and U15040 (N_15040,N_10670,N_10269);
nand U15041 (N_15041,N_12242,N_11411);
nand U15042 (N_15042,N_10110,N_12264);
nor U15043 (N_15043,N_9553,N_12251);
xor U15044 (N_15044,N_10897,N_12483);
and U15045 (N_15045,N_11373,N_11150);
and U15046 (N_15046,N_9383,N_9420);
and U15047 (N_15047,N_10531,N_9935);
nand U15048 (N_15048,N_11806,N_12035);
xnor U15049 (N_15049,N_10603,N_10421);
or U15050 (N_15050,N_11972,N_12368);
and U15051 (N_15051,N_10153,N_10787);
nor U15052 (N_15052,N_9861,N_11010);
nand U15053 (N_15053,N_10788,N_10649);
or U15054 (N_15054,N_9504,N_12331);
xnor U15055 (N_15055,N_11657,N_10761);
or U15056 (N_15056,N_11744,N_11682);
nand U15057 (N_15057,N_10045,N_9403);
or U15058 (N_15058,N_12153,N_9803);
and U15059 (N_15059,N_10586,N_11324);
nand U15060 (N_15060,N_10748,N_12198);
nand U15061 (N_15061,N_11532,N_11457);
xnor U15062 (N_15062,N_12313,N_10313);
nand U15063 (N_15063,N_10396,N_9465);
xnor U15064 (N_15064,N_11870,N_12031);
or U15065 (N_15065,N_10155,N_11003);
nand U15066 (N_15066,N_11237,N_11668);
nand U15067 (N_15067,N_11275,N_11766);
and U15068 (N_15068,N_12034,N_12386);
nand U15069 (N_15069,N_11860,N_10095);
nor U15070 (N_15070,N_12058,N_11100);
nand U15071 (N_15071,N_11004,N_10495);
or U15072 (N_15072,N_9897,N_9537);
xnor U15073 (N_15073,N_9914,N_10649);
nand U15074 (N_15074,N_11466,N_10775);
nand U15075 (N_15075,N_11037,N_11482);
nand U15076 (N_15076,N_12030,N_9486);
nand U15077 (N_15077,N_9410,N_10534);
and U15078 (N_15078,N_10378,N_9647);
nand U15079 (N_15079,N_9718,N_12237);
nand U15080 (N_15080,N_11307,N_9731);
xnor U15081 (N_15081,N_11466,N_10575);
xnor U15082 (N_15082,N_11252,N_9815);
or U15083 (N_15083,N_12026,N_9658);
nand U15084 (N_15084,N_11547,N_11668);
or U15085 (N_15085,N_10995,N_11792);
nand U15086 (N_15086,N_11672,N_11387);
or U15087 (N_15087,N_12421,N_11787);
nor U15088 (N_15088,N_12292,N_11019);
nor U15089 (N_15089,N_11953,N_11483);
or U15090 (N_15090,N_10851,N_10573);
or U15091 (N_15091,N_11982,N_10826);
nor U15092 (N_15092,N_9746,N_10883);
and U15093 (N_15093,N_9588,N_12428);
xnor U15094 (N_15094,N_12359,N_11304);
nor U15095 (N_15095,N_11470,N_10817);
xnor U15096 (N_15096,N_12179,N_12431);
and U15097 (N_15097,N_11985,N_11813);
nand U15098 (N_15098,N_11561,N_11603);
nand U15099 (N_15099,N_10028,N_12107);
or U15100 (N_15100,N_11959,N_12042);
nand U15101 (N_15101,N_11592,N_10211);
nor U15102 (N_15102,N_11071,N_12426);
or U15103 (N_15103,N_10837,N_10192);
and U15104 (N_15104,N_9769,N_10977);
nand U15105 (N_15105,N_11084,N_11008);
and U15106 (N_15106,N_10256,N_10761);
nand U15107 (N_15107,N_11129,N_10402);
nor U15108 (N_15108,N_11532,N_11954);
and U15109 (N_15109,N_10047,N_10471);
nand U15110 (N_15110,N_10876,N_10944);
or U15111 (N_15111,N_10255,N_9883);
xor U15112 (N_15112,N_11084,N_10804);
or U15113 (N_15113,N_10168,N_10820);
nor U15114 (N_15114,N_10225,N_10654);
nand U15115 (N_15115,N_11050,N_10955);
nor U15116 (N_15116,N_10214,N_12283);
and U15117 (N_15117,N_11010,N_11948);
xnor U15118 (N_15118,N_10732,N_12192);
nor U15119 (N_15119,N_12168,N_12274);
and U15120 (N_15120,N_10839,N_11364);
nand U15121 (N_15121,N_10120,N_11146);
or U15122 (N_15122,N_10833,N_9590);
nor U15123 (N_15123,N_10540,N_10191);
and U15124 (N_15124,N_12291,N_10082);
and U15125 (N_15125,N_10206,N_10654);
nor U15126 (N_15126,N_11094,N_9754);
and U15127 (N_15127,N_9514,N_9872);
nor U15128 (N_15128,N_10808,N_11132);
xnor U15129 (N_15129,N_11828,N_10375);
xnor U15130 (N_15130,N_10040,N_12005);
or U15131 (N_15131,N_11174,N_11771);
nand U15132 (N_15132,N_11181,N_9967);
and U15133 (N_15133,N_10674,N_12154);
or U15134 (N_15134,N_11197,N_10296);
nor U15135 (N_15135,N_9560,N_11116);
or U15136 (N_15136,N_11577,N_10723);
and U15137 (N_15137,N_11868,N_11473);
or U15138 (N_15138,N_11354,N_9689);
xor U15139 (N_15139,N_12215,N_11642);
or U15140 (N_15140,N_11076,N_11639);
nor U15141 (N_15141,N_12353,N_9713);
and U15142 (N_15142,N_11450,N_12030);
or U15143 (N_15143,N_11904,N_10038);
nand U15144 (N_15144,N_11590,N_9853);
nand U15145 (N_15145,N_9955,N_9554);
nor U15146 (N_15146,N_11470,N_11147);
or U15147 (N_15147,N_9425,N_11851);
nor U15148 (N_15148,N_12317,N_9627);
xnor U15149 (N_15149,N_10633,N_10793);
nand U15150 (N_15150,N_10080,N_10803);
and U15151 (N_15151,N_12174,N_11399);
and U15152 (N_15152,N_10460,N_11415);
or U15153 (N_15153,N_9782,N_12162);
and U15154 (N_15154,N_10610,N_10298);
or U15155 (N_15155,N_11221,N_10644);
nor U15156 (N_15156,N_11730,N_11518);
xnor U15157 (N_15157,N_12277,N_10815);
xnor U15158 (N_15158,N_11160,N_11652);
and U15159 (N_15159,N_9722,N_11854);
or U15160 (N_15160,N_10632,N_11055);
or U15161 (N_15161,N_10951,N_11838);
or U15162 (N_15162,N_12476,N_11553);
nor U15163 (N_15163,N_11764,N_10369);
nor U15164 (N_15164,N_12046,N_11627);
xor U15165 (N_15165,N_9393,N_10535);
and U15166 (N_15166,N_10992,N_9431);
nor U15167 (N_15167,N_11664,N_11413);
nor U15168 (N_15168,N_9676,N_9409);
xor U15169 (N_15169,N_11615,N_9735);
nor U15170 (N_15170,N_9588,N_11652);
or U15171 (N_15171,N_9379,N_11765);
or U15172 (N_15172,N_9400,N_11448);
and U15173 (N_15173,N_10061,N_10718);
nand U15174 (N_15174,N_10290,N_9528);
xor U15175 (N_15175,N_11131,N_12002);
and U15176 (N_15176,N_10127,N_9896);
and U15177 (N_15177,N_11627,N_10593);
xor U15178 (N_15178,N_10586,N_10018);
nand U15179 (N_15179,N_11777,N_9457);
nor U15180 (N_15180,N_11858,N_10466);
xnor U15181 (N_15181,N_12323,N_11633);
nand U15182 (N_15182,N_12220,N_12147);
nand U15183 (N_15183,N_12146,N_11356);
nand U15184 (N_15184,N_10940,N_11692);
xnor U15185 (N_15185,N_11372,N_11674);
nor U15186 (N_15186,N_10988,N_10327);
nor U15187 (N_15187,N_10057,N_11799);
and U15188 (N_15188,N_10297,N_9704);
xnor U15189 (N_15189,N_11269,N_10351);
nor U15190 (N_15190,N_12292,N_11203);
xor U15191 (N_15191,N_11282,N_9821);
nor U15192 (N_15192,N_10083,N_11491);
and U15193 (N_15193,N_12269,N_11025);
xor U15194 (N_15194,N_10770,N_10262);
or U15195 (N_15195,N_12216,N_10150);
xor U15196 (N_15196,N_11333,N_9548);
nor U15197 (N_15197,N_10533,N_10059);
nor U15198 (N_15198,N_10041,N_10416);
nand U15199 (N_15199,N_9389,N_11519);
nor U15200 (N_15200,N_11900,N_11282);
xnor U15201 (N_15201,N_11638,N_11224);
nor U15202 (N_15202,N_9886,N_10314);
nand U15203 (N_15203,N_11691,N_11345);
xnor U15204 (N_15204,N_10077,N_11175);
xnor U15205 (N_15205,N_9956,N_11259);
nor U15206 (N_15206,N_12214,N_10254);
nor U15207 (N_15207,N_9676,N_11500);
or U15208 (N_15208,N_11744,N_10281);
nand U15209 (N_15209,N_11491,N_9481);
xor U15210 (N_15210,N_11552,N_10187);
nor U15211 (N_15211,N_9608,N_11490);
nor U15212 (N_15212,N_10926,N_9890);
nor U15213 (N_15213,N_11836,N_11981);
nand U15214 (N_15214,N_11911,N_12179);
and U15215 (N_15215,N_12381,N_9463);
nand U15216 (N_15216,N_12018,N_11888);
and U15217 (N_15217,N_10587,N_11087);
nor U15218 (N_15218,N_11400,N_12434);
nor U15219 (N_15219,N_10514,N_11433);
nand U15220 (N_15220,N_11732,N_11779);
and U15221 (N_15221,N_12091,N_11540);
and U15222 (N_15222,N_11611,N_12044);
and U15223 (N_15223,N_10531,N_12102);
and U15224 (N_15224,N_10096,N_10886);
xnor U15225 (N_15225,N_11478,N_10983);
nand U15226 (N_15226,N_11715,N_12475);
and U15227 (N_15227,N_11016,N_11613);
nor U15228 (N_15228,N_10859,N_11121);
nor U15229 (N_15229,N_9975,N_11258);
nor U15230 (N_15230,N_12042,N_10936);
nor U15231 (N_15231,N_11918,N_10937);
nand U15232 (N_15232,N_10654,N_11310);
nand U15233 (N_15233,N_12476,N_12135);
and U15234 (N_15234,N_9784,N_12466);
or U15235 (N_15235,N_10622,N_10136);
or U15236 (N_15236,N_12383,N_11141);
nor U15237 (N_15237,N_10962,N_10761);
xor U15238 (N_15238,N_12488,N_10243);
nand U15239 (N_15239,N_11643,N_10177);
xor U15240 (N_15240,N_9437,N_9547);
nand U15241 (N_15241,N_10437,N_12079);
or U15242 (N_15242,N_10647,N_12024);
and U15243 (N_15243,N_11198,N_11990);
nand U15244 (N_15244,N_10808,N_10533);
or U15245 (N_15245,N_10644,N_11220);
or U15246 (N_15246,N_10446,N_11594);
or U15247 (N_15247,N_10315,N_11366);
nor U15248 (N_15248,N_10110,N_10381);
xnor U15249 (N_15249,N_12486,N_10524);
and U15250 (N_15250,N_12218,N_11350);
xor U15251 (N_15251,N_9908,N_10276);
and U15252 (N_15252,N_10938,N_12111);
xnor U15253 (N_15253,N_9588,N_11906);
nor U15254 (N_15254,N_10030,N_10051);
and U15255 (N_15255,N_10870,N_10416);
or U15256 (N_15256,N_11168,N_10081);
or U15257 (N_15257,N_12371,N_11881);
nand U15258 (N_15258,N_10357,N_12230);
and U15259 (N_15259,N_11060,N_10949);
nand U15260 (N_15260,N_11869,N_9928);
xnor U15261 (N_15261,N_10132,N_9897);
or U15262 (N_15262,N_12172,N_10044);
nand U15263 (N_15263,N_11659,N_12181);
nand U15264 (N_15264,N_10885,N_11147);
or U15265 (N_15265,N_12263,N_12464);
nand U15266 (N_15266,N_11051,N_10631);
nor U15267 (N_15267,N_10242,N_9519);
nand U15268 (N_15268,N_11836,N_11041);
or U15269 (N_15269,N_10648,N_10888);
nor U15270 (N_15270,N_10321,N_12097);
and U15271 (N_15271,N_11455,N_9984);
or U15272 (N_15272,N_10255,N_12246);
or U15273 (N_15273,N_11193,N_11516);
xor U15274 (N_15274,N_10009,N_9859);
nor U15275 (N_15275,N_12458,N_12280);
and U15276 (N_15276,N_11460,N_11468);
and U15277 (N_15277,N_11363,N_11742);
nand U15278 (N_15278,N_9681,N_11023);
nand U15279 (N_15279,N_10454,N_11915);
nor U15280 (N_15280,N_10700,N_10907);
and U15281 (N_15281,N_11824,N_9975);
nor U15282 (N_15282,N_11869,N_11521);
xnor U15283 (N_15283,N_9753,N_11291);
or U15284 (N_15284,N_10618,N_10529);
and U15285 (N_15285,N_10529,N_9827);
nor U15286 (N_15286,N_9722,N_10662);
xor U15287 (N_15287,N_9422,N_12081);
xor U15288 (N_15288,N_10365,N_10723);
xnor U15289 (N_15289,N_10660,N_12007);
nor U15290 (N_15290,N_9481,N_11198);
nand U15291 (N_15291,N_9552,N_11459);
nor U15292 (N_15292,N_9789,N_10147);
xnor U15293 (N_15293,N_11862,N_11527);
and U15294 (N_15294,N_11656,N_12001);
nand U15295 (N_15295,N_11066,N_10347);
xnor U15296 (N_15296,N_11195,N_10289);
or U15297 (N_15297,N_10924,N_11920);
or U15298 (N_15298,N_11851,N_10864);
and U15299 (N_15299,N_9406,N_12277);
and U15300 (N_15300,N_11006,N_10170);
xnor U15301 (N_15301,N_10676,N_10846);
xor U15302 (N_15302,N_11255,N_9832);
nand U15303 (N_15303,N_12219,N_9790);
nand U15304 (N_15304,N_10471,N_10476);
and U15305 (N_15305,N_11669,N_9676);
nor U15306 (N_15306,N_12370,N_10313);
or U15307 (N_15307,N_11628,N_10581);
or U15308 (N_15308,N_12292,N_11298);
nor U15309 (N_15309,N_12316,N_11543);
and U15310 (N_15310,N_11586,N_12093);
and U15311 (N_15311,N_9649,N_11044);
xor U15312 (N_15312,N_11428,N_11466);
nor U15313 (N_15313,N_11950,N_9382);
xor U15314 (N_15314,N_12055,N_11428);
or U15315 (N_15315,N_11576,N_12219);
xnor U15316 (N_15316,N_10073,N_10127);
xnor U15317 (N_15317,N_9387,N_9861);
and U15318 (N_15318,N_12049,N_11482);
xor U15319 (N_15319,N_11413,N_11106);
nand U15320 (N_15320,N_10396,N_10010);
and U15321 (N_15321,N_10185,N_9565);
or U15322 (N_15322,N_10786,N_12301);
or U15323 (N_15323,N_9508,N_11843);
nand U15324 (N_15324,N_10216,N_10899);
xor U15325 (N_15325,N_9415,N_11811);
and U15326 (N_15326,N_9582,N_9589);
xor U15327 (N_15327,N_9694,N_12259);
nand U15328 (N_15328,N_10817,N_11883);
nand U15329 (N_15329,N_9656,N_11251);
nand U15330 (N_15330,N_11092,N_11969);
nor U15331 (N_15331,N_10203,N_10840);
and U15332 (N_15332,N_12197,N_10431);
or U15333 (N_15333,N_10998,N_10713);
nor U15334 (N_15334,N_9434,N_12087);
or U15335 (N_15335,N_12333,N_12409);
nand U15336 (N_15336,N_10274,N_10520);
xnor U15337 (N_15337,N_12479,N_10790);
nand U15338 (N_15338,N_12368,N_9722);
nor U15339 (N_15339,N_10684,N_10968);
nand U15340 (N_15340,N_10463,N_9485);
nor U15341 (N_15341,N_11729,N_11053);
and U15342 (N_15342,N_9984,N_12147);
and U15343 (N_15343,N_12251,N_11338);
nor U15344 (N_15344,N_12308,N_12138);
nor U15345 (N_15345,N_10784,N_10857);
or U15346 (N_15346,N_10661,N_10054);
nor U15347 (N_15347,N_11470,N_11339);
and U15348 (N_15348,N_11382,N_11525);
or U15349 (N_15349,N_12231,N_9938);
nor U15350 (N_15350,N_11292,N_10557);
nor U15351 (N_15351,N_10237,N_10222);
or U15352 (N_15352,N_11242,N_9855);
nor U15353 (N_15353,N_10048,N_11140);
nand U15354 (N_15354,N_11141,N_10005);
nor U15355 (N_15355,N_12365,N_9965);
nand U15356 (N_15356,N_9534,N_12099);
nand U15357 (N_15357,N_10874,N_10535);
xnor U15358 (N_15358,N_9666,N_10633);
or U15359 (N_15359,N_12289,N_12235);
or U15360 (N_15360,N_10839,N_10860);
nand U15361 (N_15361,N_9879,N_10366);
xnor U15362 (N_15362,N_11346,N_12314);
nor U15363 (N_15363,N_11012,N_10009);
nand U15364 (N_15364,N_10802,N_10004);
nor U15365 (N_15365,N_10500,N_10423);
nor U15366 (N_15366,N_11293,N_11366);
nand U15367 (N_15367,N_10124,N_11641);
nand U15368 (N_15368,N_11721,N_11298);
and U15369 (N_15369,N_11704,N_10003);
or U15370 (N_15370,N_11667,N_11291);
xor U15371 (N_15371,N_10274,N_9741);
nand U15372 (N_15372,N_9425,N_9679);
nand U15373 (N_15373,N_12098,N_11431);
nand U15374 (N_15374,N_11594,N_10238);
or U15375 (N_15375,N_9518,N_12119);
and U15376 (N_15376,N_10306,N_10711);
nand U15377 (N_15377,N_10792,N_11981);
nor U15378 (N_15378,N_12195,N_11562);
or U15379 (N_15379,N_10024,N_10894);
xnor U15380 (N_15380,N_9528,N_10392);
nor U15381 (N_15381,N_11598,N_11499);
nor U15382 (N_15382,N_9807,N_9863);
nor U15383 (N_15383,N_11897,N_12053);
nor U15384 (N_15384,N_11723,N_9382);
xor U15385 (N_15385,N_12260,N_10633);
xor U15386 (N_15386,N_10258,N_9734);
nand U15387 (N_15387,N_9738,N_11885);
nand U15388 (N_15388,N_11523,N_10567);
xnor U15389 (N_15389,N_10319,N_11284);
and U15390 (N_15390,N_11001,N_10951);
nor U15391 (N_15391,N_11736,N_9836);
nor U15392 (N_15392,N_10730,N_10403);
or U15393 (N_15393,N_11994,N_10072);
xor U15394 (N_15394,N_11154,N_12083);
xor U15395 (N_15395,N_9908,N_10399);
and U15396 (N_15396,N_11743,N_11294);
xor U15397 (N_15397,N_11728,N_12096);
nor U15398 (N_15398,N_11237,N_11313);
or U15399 (N_15399,N_10628,N_9883);
nor U15400 (N_15400,N_10895,N_12256);
nor U15401 (N_15401,N_11052,N_10116);
nand U15402 (N_15402,N_9963,N_11950);
xor U15403 (N_15403,N_10955,N_10814);
or U15404 (N_15404,N_9957,N_11990);
and U15405 (N_15405,N_10846,N_10812);
or U15406 (N_15406,N_9617,N_12046);
nor U15407 (N_15407,N_9967,N_12143);
nand U15408 (N_15408,N_10970,N_9943);
and U15409 (N_15409,N_9635,N_9790);
or U15410 (N_15410,N_12246,N_9991);
xor U15411 (N_15411,N_11109,N_11519);
xor U15412 (N_15412,N_10773,N_9422);
xnor U15413 (N_15413,N_9615,N_10461);
and U15414 (N_15414,N_10009,N_11814);
xnor U15415 (N_15415,N_11470,N_11043);
xnor U15416 (N_15416,N_12056,N_10753);
nand U15417 (N_15417,N_10173,N_12263);
nand U15418 (N_15418,N_10363,N_11845);
nand U15419 (N_15419,N_11795,N_10394);
or U15420 (N_15420,N_10805,N_9723);
nand U15421 (N_15421,N_10192,N_11620);
nor U15422 (N_15422,N_10804,N_10545);
xor U15423 (N_15423,N_11342,N_11057);
or U15424 (N_15424,N_9582,N_10554);
or U15425 (N_15425,N_9685,N_11350);
xor U15426 (N_15426,N_10489,N_10752);
or U15427 (N_15427,N_12072,N_11919);
or U15428 (N_15428,N_10312,N_10755);
and U15429 (N_15429,N_11888,N_10399);
nand U15430 (N_15430,N_10100,N_11288);
nor U15431 (N_15431,N_11613,N_11498);
xor U15432 (N_15432,N_11820,N_10718);
or U15433 (N_15433,N_9781,N_10953);
or U15434 (N_15434,N_11743,N_10655);
or U15435 (N_15435,N_11019,N_12005);
nor U15436 (N_15436,N_11419,N_9769);
and U15437 (N_15437,N_12324,N_9779);
and U15438 (N_15438,N_10019,N_10711);
and U15439 (N_15439,N_11795,N_11401);
or U15440 (N_15440,N_10714,N_11031);
nor U15441 (N_15441,N_11780,N_11603);
and U15442 (N_15442,N_11106,N_9415);
xor U15443 (N_15443,N_10463,N_10376);
xor U15444 (N_15444,N_11426,N_10799);
and U15445 (N_15445,N_10225,N_10680);
nor U15446 (N_15446,N_9974,N_10627);
or U15447 (N_15447,N_10707,N_11420);
nor U15448 (N_15448,N_10780,N_12262);
xor U15449 (N_15449,N_10560,N_10184);
nand U15450 (N_15450,N_10057,N_11526);
xor U15451 (N_15451,N_10495,N_9716);
and U15452 (N_15452,N_10443,N_11724);
nor U15453 (N_15453,N_10855,N_10754);
xor U15454 (N_15454,N_10617,N_10272);
and U15455 (N_15455,N_11538,N_10127);
or U15456 (N_15456,N_9908,N_10948);
nor U15457 (N_15457,N_11819,N_9773);
and U15458 (N_15458,N_10401,N_11370);
and U15459 (N_15459,N_12259,N_10759);
nand U15460 (N_15460,N_11126,N_10551);
nand U15461 (N_15461,N_10808,N_10899);
nand U15462 (N_15462,N_10586,N_12244);
or U15463 (N_15463,N_11677,N_10758);
nor U15464 (N_15464,N_12277,N_10014);
nor U15465 (N_15465,N_9573,N_11565);
nand U15466 (N_15466,N_11772,N_11301);
or U15467 (N_15467,N_11088,N_9580);
nand U15468 (N_15468,N_11425,N_9636);
xnor U15469 (N_15469,N_10187,N_10622);
and U15470 (N_15470,N_10145,N_11475);
and U15471 (N_15471,N_12124,N_10026);
and U15472 (N_15472,N_9905,N_11663);
nor U15473 (N_15473,N_9928,N_9434);
or U15474 (N_15474,N_12241,N_11727);
and U15475 (N_15475,N_11965,N_10179);
nor U15476 (N_15476,N_11213,N_9593);
nor U15477 (N_15477,N_11654,N_10992);
xnor U15478 (N_15478,N_12309,N_12082);
nand U15479 (N_15479,N_10601,N_10404);
nor U15480 (N_15480,N_12268,N_9641);
xor U15481 (N_15481,N_10042,N_10797);
or U15482 (N_15482,N_10979,N_9869);
nand U15483 (N_15483,N_9880,N_9744);
nor U15484 (N_15484,N_9938,N_11141);
nor U15485 (N_15485,N_11438,N_11232);
nor U15486 (N_15486,N_11108,N_10973);
nor U15487 (N_15487,N_12323,N_11835);
and U15488 (N_15488,N_9624,N_11525);
nand U15489 (N_15489,N_10393,N_11033);
xor U15490 (N_15490,N_9677,N_12059);
and U15491 (N_15491,N_9679,N_11747);
and U15492 (N_15492,N_9658,N_10082);
or U15493 (N_15493,N_12128,N_12270);
xor U15494 (N_15494,N_10836,N_12407);
xnor U15495 (N_15495,N_11445,N_10740);
nand U15496 (N_15496,N_11203,N_11747);
and U15497 (N_15497,N_10213,N_11874);
or U15498 (N_15498,N_11121,N_11950);
or U15499 (N_15499,N_11167,N_10935);
nand U15500 (N_15500,N_10339,N_9394);
nor U15501 (N_15501,N_12300,N_10202);
nand U15502 (N_15502,N_11472,N_9668);
xor U15503 (N_15503,N_10654,N_11076);
nor U15504 (N_15504,N_11670,N_9403);
nor U15505 (N_15505,N_9431,N_10107);
xnor U15506 (N_15506,N_12342,N_11797);
or U15507 (N_15507,N_12166,N_9476);
xnor U15508 (N_15508,N_11314,N_12060);
or U15509 (N_15509,N_10707,N_9815);
or U15510 (N_15510,N_9770,N_10294);
and U15511 (N_15511,N_11245,N_10196);
or U15512 (N_15512,N_11650,N_9634);
nand U15513 (N_15513,N_10398,N_10113);
and U15514 (N_15514,N_12045,N_11345);
nor U15515 (N_15515,N_11653,N_10673);
nor U15516 (N_15516,N_9420,N_10446);
and U15517 (N_15517,N_11735,N_12431);
nand U15518 (N_15518,N_9494,N_11394);
nor U15519 (N_15519,N_11838,N_10255);
or U15520 (N_15520,N_11543,N_10930);
xnor U15521 (N_15521,N_9782,N_12104);
nand U15522 (N_15522,N_11891,N_10779);
nand U15523 (N_15523,N_10828,N_9897);
and U15524 (N_15524,N_10709,N_11299);
xnor U15525 (N_15525,N_10957,N_12101);
and U15526 (N_15526,N_9663,N_9911);
xnor U15527 (N_15527,N_10264,N_10863);
nand U15528 (N_15528,N_9657,N_11501);
xor U15529 (N_15529,N_12022,N_9938);
nor U15530 (N_15530,N_10185,N_9876);
or U15531 (N_15531,N_12367,N_10064);
nor U15532 (N_15532,N_10033,N_11313);
xor U15533 (N_15533,N_10411,N_12325);
xnor U15534 (N_15534,N_12022,N_10187);
nor U15535 (N_15535,N_12063,N_11221);
and U15536 (N_15536,N_10591,N_10544);
nor U15537 (N_15537,N_11220,N_11138);
and U15538 (N_15538,N_9970,N_10517);
nand U15539 (N_15539,N_12156,N_10511);
xnor U15540 (N_15540,N_10551,N_9528);
xor U15541 (N_15541,N_9945,N_11643);
xnor U15542 (N_15542,N_12420,N_9476);
and U15543 (N_15543,N_11016,N_12194);
or U15544 (N_15544,N_10424,N_10468);
and U15545 (N_15545,N_12171,N_12303);
or U15546 (N_15546,N_10750,N_9681);
nor U15547 (N_15547,N_11422,N_11690);
nand U15548 (N_15548,N_9526,N_10253);
xor U15549 (N_15549,N_11612,N_10848);
or U15550 (N_15550,N_9556,N_12001);
nand U15551 (N_15551,N_10664,N_10449);
xor U15552 (N_15552,N_9780,N_10106);
and U15553 (N_15553,N_9927,N_9975);
nand U15554 (N_15554,N_11425,N_11438);
nor U15555 (N_15555,N_11459,N_10956);
nand U15556 (N_15556,N_11795,N_9996);
xor U15557 (N_15557,N_12060,N_10804);
xnor U15558 (N_15558,N_9873,N_10300);
or U15559 (N_15559,N_10838,N_10401);
nand U15560 (N_15560,N_10548,N_10540);
nand U15561 (N_15561,N_10781,N_10808);
nor U15562 (N_15562,N_10829,N_12370);
and U15563 (N_15563,N_9804,N_11780);
and U15564 (N_15564,N_11070,N_10448);
nand U15565 (N_15565,N_9854,N_9704);
nand U15566 (N_15566,N_11104,N_9972);
or U15567 (N_15567,N_9601,N_10766);
xnor U15568 (N_15568,N_11294,N_12164);
and U15569 (N_15569,N_11314,N_10592);
xnor U15570 (N_15570,N_9752,N_11202);
xor U15571 (N_15571,N_10216,N_11476);
and U15572 (N_15572,N_12057,N_9528);
nor U15573 (N_15573,N_11821,N_10755);
nor U15574 (N_15574,N_10291,N_9994);
nand U15575 (N_15575,N_10692,N_11288);
nor U15576 (N_15576,N_11567,N_9887);
or U15577 (N_15577,N_10561,N_10250);
nor U15578 (N_15578,N_11700,N_9401);
nand U15579 (N_15579,N_11388,N_9903);
nand U15580 (N_15580,N_11034,N_11144);
xnor U15581 (N_15581,N_12157,N_9838);
and U15582 (N_15582,N_10254,N_9686);
nor U15583 (N_15583,N_12067,N_10567);
nand U15584 (N_15584,N_9983,N_9407);
xnor U15585 (N_15585,N_11053,N_10176);
nand U15586 (N_15586,N_11233,N_10129);
nand U15587 (N_15587,N_9664,N_10263);
nand U15588 (N_15588,N_10757,N_11700);
nand U15589 (N_15589,N_10271,N_10770);
nand U15590 (N_15590,N_11727,N_10386);
xnor U15591 (N_15591,N_11813,N_10934);
nor U15592 (N_15592,N_9703,N_9429);
nor U15593 (N_15593,N_10502,N_9694);
or U15594 (N_15594,N_11837,N_11627);
xnor U15595 (N_15595,N_9379,N_9828);
nor U15596 (N_15596,N_12227,N_12178);
or U15597 (N_15597,N_9807,N_10683);
or U15598 (N_15598,N_11878,N_10529);
nor U15599 (N_15599,N_11260,N_10375);
and U15600 (N_15600,N_9972,N_11847);
or U15601 (N_15601,N_10099,N_12143);
xnor U15602 (N_15602,N_12234,N_10315);
nand U15603 (N_15603,N_10576,N_11930);
xor U15604 (N_15604,N_11159,N_9793);
and U15605 (N_15605,N_11899,N_11415);
nand U15606 (N_15606,N_10806,N_10807);
nor U15607 (N_15607,N_11288,N_9900);
nor U15608 (N_15608,N_11831,N_12274);
nor U15609 (N_15609,N_9675,N_9482);
or U15610 (N_15610,N_9909,N_9920);
and U15611 (N_15611,N_11984,N_11856);
nand U15612 (N_15612,N_11935,N_9637);
or U15613 (N_15613,N_11410,N_9553);
or U15614 (N_15614,N_11846,N_11298);
xor U15615 (N_15615,N_10473,N_12479);
and U15616 (N_15616,N_11267,N_10957);
nand U15617 (N_15617,N_9968,N_11756);
or U15618 (N_15618,N_12499,N_11111);
or U15619 (N_15619,N_12015,N_10978);
nand U15620 (N_15620,N_9709,N_10356);
and U15621 (N_15621,N_10600,N_10385);
or U15622 (N_15622,N_9765,N_10609);
nand U15623 (N_15623,N_9415,N_11660);
nand U15624 (N_15624,N_11722,N_11837);
xnor U15625 (N_15625,N_13439,N_14401);
or U15626 (N_15626,N_14887,N_13143);
and U15627 (N_15627,N_14524,N_15477);
or U15628 (N_15628,N_13026,N_14538);
nand U15629 (N_15629,N_13000,N_13263);
nor U15630 (N_15630,N_13607,N_15085);
nor U15631 (N_15631,N_15252,N_13481);
xnor U15632 (N_15632,N_13810,N_15219);
nor U15633 (N_15633,N_14807,N_14329);
and U15634 (N_15634,N_14744,N_13198);
and U15635 (N_15635,N_14178,N_12666);
xnor U15636 (N_15636,N_13638,N_14209);
xor U15637 (N_15637,N_15262,N_15323);
nand U15638 (N_15638,N_14537,N_13862);
and U15639 (N_15639,N_12570,N_12942);
nor U15640 (N_15640,N_14233,N_14529);
nor U15641 (N_15641,N_14005,N_15023);
and U15642 (N_15642,N_14086,N_13657);
xnor U15643 (N_15643,N_15165,N_12653);
or U15644 (N_15644,N_15485,N_14669);
nor U15645 (N_15645,N_15601,N_13521);
or U15646 (N_15646,N_13108,N_14316);
and U15647 (N_15647,N_13393,N_14013);
or U15648 (N_15648,N_13658,N_15494);
and U15649 (N_15649,N_13881,N_13330);
nor U15650 (N_15650,N_13407,N_13970);
or U15651 (N_15651,N_15435,N_13113);
nand U15652 (N_15652,N_13733,N_15375);
and U15653 (N_15653,N_15205,N_12893);
xnor U15654 (N_15654,N_13270,N_15214);
nor U15655 (N_15655,N_13751,N_14254);
and U15656 (N_15656,N_14126,N_13338);
nor U15657 (N_15657,N_15381,N_14167);
and U15658 (N_15658,N_13559,N_14014);
nor U15659 (N_15659,N_14639,N_13792);
xor U15660 (N_15660,N_12650,N_13651);
and U15661 (N_15661,N_14407,N_15519);
and U15662 (N_15662,N_14196,N_13546);
nand U15663 (N_15663,N_13323,N_14393);
and U15664 (N_15664,N_13560,N_15233);
xor U15665 (N_15665,N_15571,N_15129);
nor U15666 (N_15666,N_12609,N_15545);
xor U15667 (N_15667,N_14593,N_13401);
nand U15668 (N_15668,N_13177,N_15208);
or U15669 (N_15669,N_14979,N_14957);
nand U15670 (N_15670,N_13427,N_13642);
xor U15671 (N_15671,N_14309,N_14478);
nand U15672 (N_15672,N_13660,N_14519);
and U15673 (N_15673,N_14285,N_14442);
or U15674 (N_15674,N_14745,N_12999);
xor U15675 (N_15675,N_14720,N_15569);
xnor U15676 (N_15676,N_12784,N_12847);
nand U15677 (N_15677,N_13618,N_15296);
and U15678 (N_15678,N_14997,N_12800);
or U15679 (N_15679,N_13626,N_15617);
xnor U15680 (N_15680,N_13024,N_13085);
nand U15681 (N_15681,N_14444,N_15125);
and U15682 (N_15682,N_12689,N_13948);
xnor U15683 (N_15683,N_14873,N_14378);
or U15684 (N_15684,N_12756,N_14037);
or U15685 (N_15685,N_13678,N_14068);
and U15686 (N_15686,N_12521,N_13919);
or U15687 (N_15687,N_12972,N_13193);
or U15688 (N_15688,N_14334,N_14166);
or U15689 (N_15689,N_13372,N_12757);
nor U15690 (N_15690,N_12662,N_14203);
nor U15691 (N_15691,N_14297,N_13692);
nand U15692 (N_15692,N_14644,N_14643);
xor U15693 (N_15693,N_13708,N_14119);
and U15694 (N_15694,N_13191,N_13971);
and U15695 (N_15695,N_15605,N_12714);
or U15696 (N_15696,N_13664,N_12811);
or U15697 (N_15697,N_14223,N_12952);
nor U15698 (N_15698,N_15552,N_13368);
nand U15699 (N_15699,N_15489,N_13687);
or U15700 (N_15700,N_15027,N_14604);
nor U15701 (N_15701,N_12926,N_15495);
or U15702 (N_15702,N_13284,N_13420);
nand U15703 (N_15703,N_13851,N_12629);
nand U15704 (N_15704,N_13452,N_13963);
nor U15705 (N_15705,N_15531,N_13227);
or U15706 (N_15706,N_15015,N_15578);
xnor U15707 (N_15707,N_15326,N_14208);
or U15708 (N_15708,N_14279,N_14243);
or U15709 (N_15709,N_14805,N_14383);
or U15710 (N_15710,N_12635,N_14556);
nor U15711 (N_15711,N_12815,N_14812);
or U15712 (N_15712,N_14139,N_15157);
and U15713 (N_15713,N_13916,N_14433);
and U15714 (N_15714,N_13679,N_15022);
xor U15715 (N_15715,N_12956,N_15332);
xor U15716 (N_15716,N_13869,N_14295);
and U15717 (N_15717,N_13899,N_14082);
nand U15718 (N_15718,N_15091,N_14883);
nor U15719 (N_15719,N_14271,N_14814);
nand U15720 (N_15720,N_12613,N_13415);
xnor U15721 (N_15721,N_13867,N_14753);
xnor U15722 (N_15722,N_14311,N_12920);
nor U15723 (N_15723,N_12979,N_13097);
xnor U15724 (N_15724,N_13265,N_13115);
nor U15725 (N_15725,N_12987,N_12580);
and U15726 (N_15726,N_13671,N_15436);
nand U15727 (N_15727,N_14722,N_14616);
nor U15728 (N_15728,N_13061,N_12673);
nand U15729 (N_15729,N_14029,N_14924);
nor U15730 (N_15730,N_15378,N_15450);
nor U15731 (N_15731,N_14354,N_14965);
or U15732 (N_15732,N_15538,N_13170);
nand U15733 (N_15733,N_12789,N_12581);
nand U15734 (N_15734,N_14041,N_13922);
nor U15735 (N_15735,N_14816,N_13553);
nor U15736 (N_15736,N_13595,N_12870);
and U15737 (N_15737,N_15272,N_14933);
or U15738 (N_15738,N_14259,N_12592);
nand U15739 (N_15739,N_14040,N_13258);
or U15740 (N_15740,N_12879,N_13539);
nand U15741 (N_15741,N_14100,N_14060);
and U15742 (N_15742,N_15056,N_13842);
and U15743 (N_15743,N_14776,N_15146);
or U15744 (N_15744,N_15393,N_14423);
nor U15745 (N_15745,N_12659,N_13823);
xor U15746 (N_15746,N_13296,N_14467);
xor U15747 (N_15747,N_14567,N_12993);
or U15748 (N_15748,N_15028,N_14514);
nand U15749 (N_15749,N_13160,N_13925);
xnor U15750 (N_15750,N_14622,N_12769);
or U15751 (N_15751,N_13850,N_12888);
and U15752 (N_15752,N_14098,N_14505);
nand U15753 (N_15753,N_13759,N_14080);
nor U15754 (N_15754,N_12701,N_13474);
or U15755 (N_15755,N_12908,N_13279);
and U15756 (N_15756,N_12686,N_12755);
or U15757 (N_15757,N_14735,N_14661);
or U15758 (N_15758,N_15528,N_13798);
nor U15759 (N_15759,N_12643,N_13503);
and U15760 (N_15760,N_13527,N_12572);
or U15761 (N_15761,N_14688,N_13321);
or U15762 (N_15762,N_13286,N_13659);
xor U15763 (N_15763,N_14863,N_14509);
and U15764 (N_15764,N_14594,N_13973);
nor U15765 (N_15765,N_15583,N_14332);
nor U15766 (N_15766,N_12700,N_13102);
nor U15767 (N_15767,N_13755,N_13051);
nand U15768 (N_15768,N_14437,N_14135);
xnor U15769 (N_15769,N_13366,N_13103);
and U15770 (N_15770,N_14762,N_14857);
xor U15771 (N_15771,N_15213,N_15101);
nor U15772 (N_15772,N_14278,N_15620);
nand U15773 (N_15773,N_12568,N_15461);
nor U15774 (N_15774,N_13545,N_14304);
or U15775 (N_15775,N_15425,N_13905);
nor U15776 (N_15776,N_14012,N_13721);
nand U15777 (N_15777,N_14230,N_13735);
and U15778 (N_15778,N_13073,N_14881);
xor U15779 (N_15779,N_15610,N_13932);
nor U15780 (N_15780,N_12895,N_13267);
nor U15781 (N_15781,N_14472,N_14637);
nand U15782 (N_15782,N_15216,N_13730);
or U15783 (N_15783,N_14697,N_15422);
and U15784 (N_15784,N_14928,N_13579);
xnor U15785 (N_15785,N_12837,N_15224);
nor U15786 (N_15786,N_13358,N_15618);
xor U15787 (N_15787,N_13463,N_13734);
or U15788 (N_15788,N_14084,N_14947);
or U15789 (N_15789,N_15033,N_14199);
and U15790 (N_15790,N_13133,N_13602);
nor U15791 (N_15791,N_12709,N_13859);
xor U15792 (N_15792,N_14460,N_12692);
xnor U15793 (N_15793,N_15453,N_14303);
nor U15794 (N_15794,N_12678,N_12937);
nand U15795 (N_15795,N_15162,N_14476);
xnor U15796 (N_15796,N_13610,N_14206);
nand U15797 (N_15797,N_14930,N_13641);
or U15798 (N_15798,N_15548,N_12736);
xnor U15799 (N_15799,N_13081,N_15234);
nand U15800 (N_15800,N_13383,N_13957);
nand U15801 (N_15801,N_14090,N_15590);
or U15802 (N_15802,N_15096,N_13257);
nor U15803 (N_15803,N_13414,N_14482);
or U15804 (N_15804,N_13192,N_14314);
or U15805 (N_15805,N_13036,N_14019);
or U15806 (N_15806,N_14999,N_15555);
nand U15807 (N_15807,N_12681,N_15562);
and U15808 (N_15808,N_14520,N_12634);
and U15809 (N_15809,N_14511,N_13001);
and U15810 (N_15810,N_14531,N_13886);
nor U15811 (N_15811,N_15225,N_13964);
and U15812 (N_15812,N_14038,N_14020);
nor U15813 (N_15813,N_14063,N_13966);
nand U15814 (N_15814,N_15361,N_14061);
or U15815 (N_15815,N_14749,N_12916);
and U15816 (N_15816,N_15034,N_14764);
nand U15817 (N_15817,N_14907,N_14974);
and U15818 (N_15818,N_13322,N_13513);
nor U15819 (N_15819,N_13978,N_14198);
nor U15820 (N_15820,N_14569,N_14559);
and U15821 (N_15821,N_12564,N_14351);
nor U15822 (N_15822,N_12781,N_14092);
xnor U15823 (N_15823,N_15557,N_14898);
or U15824 (N_15824,N_12991,N_13608);
nand U15825 (N_15825,N_14077,N_13235);
and U15826 (N_15826,N_12642,N_13337);
and U15827 (N_15827,N_14612,N_13077);
and U15828 (N_15828,N_13013,N_14961);
xnor U15829 (N_15829,N_12886,N_13132);
and U15830 (N_15830,N_14513,N_14789);
nor U15831 (N_15831,N_14874,N_15313);
or U15832 (N_15832,N_12799,N_14544);
nand U15833 (N_15833,N_13316,N_12896);
and U15834 (N_15834,N_14220,N_13057);
nor U15835 (N_15835,N_14436,N_15051);
nand U15836 (N_15836,N_12721,N_13448);
nor U15837 (N_15837,N_15054,N_14809);
or U15838 (N_15838,N_14318,N_14684);
nand U15839 (N_15839,N_14496,N_13949);
nand U15840 (N_15840,N_14871,N_14694);
xnor U15841 (N_15841,N_12667,N_14824);
nand U15842 (N_15842,N_13391,N_13845);
nor U15843 (N_15843,N_15181,N_14668);
nand U15844 (N_15844,N_15389,N_12880);
or U15845 (N_15845,N_14676,N_15044);
or U15846 (N_15846,N_15065,N_14959);
xor U15847 (N_15847,N_12626,N_14258);
and U15848 (N_15848,N_14530,N_13529);
nor U15849 (N_15849,N_14911,N_13390);
and U15850 (N_15850,N_14186,N_15151);
and U15851 (N_15851,N_13083,N_14667);
xnor U15852 (N_15852,N_13697,N_15001);
nor U15853 (N_15853,N_15619,N_13885);
or U15854 (N_15854,N_13939,N_15532);
and U15855 (N_15855,N_14611,N_15246);
nand U15856 (N_15856,N_14076,N_14360);
or U15857 (N_15857,N_15182,N_12892);
or U15858 (N_15858,N_13802,N_15149);
nor U15859 (N_15859,N_12695,N_14692);
nand U15860 (N_15860,N_12812,N_12531);
nor U15861 (N_15861,N_14937,N_14189);
xor U15862 (N_15862,N_15573,N_14811);
or U15863 (N_15863,N_13161,N_12929);
nand U15864 (N_15864,N_13066,N_12860);
xor U15865 (N_15865,N_14369,N_13389);
and U15866 (N_15866,N_13351,N_14103);
xnor U15867 (N_15867,N_14382,N_14570);
nor U15868 (N_15868,N_13185,N_13451);
nor U15869 (N_15869,N_13022,N_12873);
or U15870 (N_15870,N_12992,N_13433);
nor U15871 (N_15871,N_12541,N_14147);
nor U15872 (N_15872,N_15241,N_14630);
nand U15873 (N_15873,N_13590,N_14112);
and U15874 (N_15874,N_15404,N_13682);
and U15875 (N_15875,N_14728,N_14244);
and U15876 (N_15876,N_13134,N_12522);
xor U15877 (N_15877,N_15206,N_15097);
or U15878 (N_15878,N_15077,N_12618);
nor U15879 (N_15879,N_14758,N_12851);
and U15880 (N_15880,N_15322,N_14024);
or U15881 (N_15881,N_14845,N_12923);
nor U15882 (N_15882,N_13172,N_13281);
nor U15883 (N_15883,N_12676,N_12788);
nand U15884 (N_15884,N_13801,N_14867);
xnor U15885 (N_15885,N_13982,N_13774);
nand U15886 (N_15886,N_13847,N_13226);
nor U15887 (N_15887,N_12682,N_14497);
or U15888 (N_15888,N_14249,N_13526);
nand U15889 (N_15889,N_13731,N_13570);
or U15890 (N_15890,N_12932,N_13770);
or U15891 (N_15891,N_15576,N_12770);
and U15892 (N_15892,N_13897,N_15328);
xor U15893 (N_15893,N_13476,N_14308);
xnor U15894 (N_15894,N_13450,N_13558);
or U15895 (N_15895,N_15368,N_14836);
or U15896 (N_15896,N_13969,N_14057);
or U15897 (N_15897,N_15265,N_12761);
nor U15898 (N_15898,N_15533,N_13187);
nand U15899 (N_15899,N_12834,N_15259);
or U15900 (N_15900,N_15093,N_14225);
nor U15901 (N_15901,N_14251,N_12985);
and U15902 (N_15902,N_14118,N_13574);
xnor U15903 (N_15903,N_13411,N_14335);
and U15904 (N_15904,N_13631,N_14282);
or U15905 (N_15905,N_12945,N_13662);
and U15906 (N_15906,N_13706,N_12619);
nand U15907 (N_15907,N_14227,N_14575);
nand U15908 (N_15908,N_13466,N_14647);
nand U15909 (N_15909,N_13713,N_12658);
xor U15910 (N_15910,N_15372,N_14266);
or U15911 (N_15911,N_14333,N_13856);
nor U15912 (N_15912,N_15602,N_13345);
nand U15913 (N_15913,N_12625,N_13153);
xor U15914 (N_15914,N_12906,N_14331);
or U15915 (N_15915,N_14588,N_13917);
and U15916 (N_15916,N_15142,N_13099);
nand U15917 (N_15917,N_14671,N_13750);
xor U15918 (N_15918,N_15579,N_15064);
xnor U15919 (N_15919,N_14840,N_14847);
nand U15920 (N_15920,N_13581,N_14218);
xor U15921 (N_15921,N_14365,N_13870);
nand U15922 (N_15922,N_15179,N_13566);
xnor U15923 (N_15923,N_13266,N_15577);
and U15924 (N_15924,N_14821,N_13627);
and U15925 (N_15925,N_15115,N_12545);
xor U15926 (N_15926,N_15408,N_12639);
nor U15927 (N_15927,N_15013,N_13309);
or U15928 (N_15928,N_15544,N_14434);
and U15929 (N_15929,N_15462,N_12567);
nor U15930 (N_15930,N_15396,N_14348);
xnor U15931 (N_15931,N_15426,N_13512);
and U15932 (N_15932,N_12790,N_13815);
and U15933 (N_15933,N_14507,N_13923);
nor U15934 (N_15934,N_13577,N_13274);
and U15935 (N_15935,N_12930,N_14670);
nor U15936 (N_15936,N_13457,N_12914);
nor U15937 (N_15937,N_14522,N_13645);
and U15938 (N_15938,N_14344,N_14817);
nor U15939 (N_15939,N_15572,N_13853);
nor U15940 (N_15940,N_13069,N_13008);
nor U15941 (N_15941,N_13540,N_13354);
nand U15942 (N_15942,N_13264,N_13091);
and U15943 (N_15943,N_13222,N_13269);
nor U15944 (N_15944,N_13890,N_12713);
nor U15945 (N_15945,N_13501,N_12708);
nand U15946 (N_15946,N_13704,N_14499);
nor U15947 (N_15947,N_13929,N_14173);
nand U15948 (N_15948,N_12868,N_13328);
and U15949 (N_15949,N_13533,N_15133);
nand U15950 (N_15950,N_12954,N_13883);
nor U15951 (N_15951,N_12752,N_13055);
nor U15952 (N_15952,N_12696,N_13686);
and U15953 (N_15953,N_12586,N_13882);
nand U15954 (N_15954,N_14168,N_12772);
nor U15955 (N_15955,N_14016,N_14835);
or U15956 (N_15956,N_15419,N_15291);
and U15957 (N_15957,N_14034,N_15243);
and U15958 (N_15958,N_14778,N_12728);
and U15959 (N_15959,N_14006,N_14690);
or U15960 (N_15960,N_14958,N_14886);
nand U15961 (N_15961,N_14700,N_14602);
nand U15962 (N_15962,N_12501,N_15043);
xor U15963 (N_15963,N_15014,N_14281);
and U15964 (N_15964,N_13100,N_15180);
nand U15965 (N_15965,N_14204,N_14683);
xor U15966 (N_15966,N_13280,N_14440);
nand U15967 (N_15967,N_13889,N_14754);
and U15968 (N_15968,N_14919,N_12960);
nor U15969 (N_15969,N_14272,N_14158);
nand U15970 (N_15970,N_15428,N_13443);
or U15971 (N_15971,N_14326,N_14806);
nor U15972 (N_15972,N_15148,N_15209);
nor U15973 (N_15973,N_14490,N_12943);
or U15974 (N_15974,N_13173,N_15460);
and U15975 (N_15975,N_14641,N_15276);
nand U15976 (N_15976,N_13833,N_14384);
nand U15977 (N_15977,N_14414,N_14783);
or U15978 (N_15978,N_12632,N_14459);
nor U15979 (N_15979,N_15607,N_13146);
and U15980 (N_15980,N_13873,N_13783);
and U15981 (N_15981,N_12884,N_14302);
xnor U15982 (N_15982,N_12502,N_14404);
nor U15983 (N_15983,N_12711,N_14398);
nand U15984 (N_15984,N_15052,N_14108);
nand U15985 (N_15985,N_13648,N_12824);
nand U15986 (N_15986,N_15401,N_15502);
nand U15987 (N_15987,N_15581,N_14070);
nand U15988 (N_15988,N_13837,N_13646);
xnor U15989 (N_15989,N_13199,N_14441);
nor U15990 (N_15990,N_14317,N_13903);
nor U15991 (N_15991,N_14897,N_13991);
nand U15992 (N_15992,N_13405,N_14978);
xnor U15993 (N_15993,N_15138,N_13567);
xnor U15994 (N_15994,N_13760,N_13287);
and U15995 (N_15995,N_12746,N_13586);
or U15996 (N_15996,N_14381,N_14572);
nor U15997 (N_15997,N_13084,N_14983);
nor U15998 (N_15998,N_13339,N_13117);
or U15999 (N_15999,N_12699,N_15000);
nand U16000 (N_16000,N_13497,N_14457);
or U16001 (N_16001,N_14051,N_13934);
or U16002 (N_16002,N_13406,N_14923);
or U16003 (N_16003,N_13872,N_15456);
or U16004 (N_16004,N_14212,N_14768);
nor U16005 (N_16005,N_13454,N_15513);
nor U16006 (N_16006,N_12691,N_12743);
or U16007 (N_16007,N_14844,N_15364);
nor U16008 (N_16008,N_15273,N_15311);
and U16009 (N_16009,N_13650,N_12876);
nand U16010 (N_16010,N_13749,N_12814);
and U16011 (N_16011,N_14386,N_15038);
xnor U16012 (N_16012,N_14548,N_12633);
or U16013 (N_16013,N_14165,N_15437);
and U16014 (N_16014,N_15307,N_13125);
xor U16015 (N_16015,N_12583,N_12543);
or U16016 (N_16016,N_13067,N_15459);
and U16017 (N_16017,N_13254,N_14798);
or U16018 (N_16018,N_15238,N_15338);
nor U16019 (N_16019,N_13860,N_15210);
and U16020 (N_16020,N_12971,N_14663);
and U16021 (N_16021,N_14732,N_14132);
or U16022 (N_16022,N_13275,N_15277);
xor U16023 (N_16023,N_12842,N_14918);
nand U16024 (N_16024,N_15183,N_14955);
and U16025 (N_16025,N_13907,N_14445);
nand U16026 (N_16026,N_13998,N_14842);
nor U16027 (N_16027,N_13362,N_13259);
xnor U16028 (N_16028,N_12602,N_12684);
nand U16029 (N_16029,N_12882,N_14127);
nand U16030 (N_16030,N_13805,N_13725);
nor U16031 (N_16031,N_13348,N_15228);
or U16032 (N_16032,N_15127,N_14179);
or U16033 (N_16033,N_12938,N_15229);
nor U16034 (N_16034,N_14884,N_15248);
nor U16035 (N_16035,N_12671,N_14665);
nand U16036 (N_16036,N_14938,N_13129);
nor U16037 (N_16037,N_15195,N_13344);
nor U16038 (N_16038,N_15122,N_13643);
xnor U16039 (N_16039,N_13285,N_14320);
or U16040 (N_16040,N_13688,N_13863);
xor U16041 (N_16041,N_15455,N_13828);
and U16042 (N_16042,N_14833,N_13892);
xnor U16043 (N_16043,N_13060,N_13156);
nor U16044 (N_16044,N_14658,N_14736);
or U16045 (N_16045,N_14096,N_14280);
nor U16046 (N_16046,N_13297,N_13569);
xor U16047 (N_16047,N_13848,N_12516);
xnor U16048 (N_16048,N_12959,N_14679);
nor U16049 (N_16049,N_15119,N_15624);
nor U16050 (N_16050,N_12672,N_13206);
nand U16051 (N_16051,N_14231,N_14944);
nand U16052 (N_16052,N_14053,N_14546);
nand U16053 (N_16053,N_12883,N_14673);
xor U16054 (N_16054,N_15141,N_15221);
or U16055 (N_16055,N_15342,N_15185);
xor U16056 (N_16056,N_14257,N_15287);
nor U16057 (N_16057,N_14095,N_12566);
nand U16058 (N_16058,N_14562,N_14325);
or U16059 (N_16059,N_13087,N_13082);
and U16060 (N_16060,N_14042,N_12900);
or U16061 (N_16061,N_14422,N_13661);
and U16062 (N_16062,N_15104,N_15433);
nor U16063 (N_16063,N_12702,N_13542);
nor U16064 (N_16064,N_12912,N_13397);
or U16065 (N_16065,N_13467,N_13684);
xnor U16066 (N_16066,N_13655,N_14370);
nand U16067 (N_16067,N_13176,N_14599);
xor U16068 (N_16068,N_12969,N_13827);
nand U16069 (N_16069,N_14138,N_12948);
or U16070 (N_16070,N_12795,N_15175);
nand U16071 (N_16071,N_12950,N_13728);
nor U16072 (N_16072,N_15463,N_12760);
nor U16073 (N_16073,N_12511,N_14312);
and U16074 (N_16074,N_12525,N_14337);
nand U16075 (N_16075,N_15199,N_14343);
nor U16076 (N_16076,N_13238,N_15440);
or U16077 (N_16077,N_14977,N_14859);
xor U16078 (N_16078,N_14693,N_14703);
nand U16079 (N_16079,N_14150,N_15534);
xnor U16080 (N_16080,N_13909,N_15008);
or U16081 (N_16081,N_15343,N_15187);
and U16082 (N_16082,N_15334,N_13895);
and U16083 (N_16083,N_13044,N_14960);
nor U16084 (N_16084,N_13928,N_13753);
nor U16085 (N_16085,N_13906,N_13288);
xnor U16086 (N_16086,N_14526,N_13814);
or U16087 (N_16087,N_15400,N_15042);
and U16088 (N_16088,N_13311,N_15524);
xnor U16089 (N_16089,N_15503,N_14431);
nor U16090 (N_16090,N_15299,N_15444);
or U16091 (N_16091,N_13294,N_13633);
nor U16092 (N_16092,N_13628,N_14319);
and U16093 (N_16093,N_12648,N_13699);
and U16094 (N_16094,N_15212,N_15472);
and U16095 (N_16095,N_14116,N_12820);
nor U16096 (N_16096,N_14675,N_13130);
and U16097 (N_16097,N_13380,N_15196);
nand U16098 (N_16098,N_13653,N_12890);
or U16099 (N_16099,N_14408,N_12745);
or U16100 (N_16100,N_14525,N_15082);
nand U16101 (N_16101,N_12638,N_13032);
nor U16102 (N_16102,N_15554,N_15188);
nand U16103 (N_16103,N_15025,N_14253);
xnor U16104 (N_16104,N_14448,N_12517);
nand U16105 (N_16105,N_14267,N_14195);
xor U16106 (N_16106,N_13891,N_15611);
nor U16107 (N_16107,N_14839,N_14626);
nor U16108 (N_16108,N_13575,N_15121);
nor U16109 (N_16109,N_13544,N_13681);
or U16110 (N_16110,N_15349,N_12835);
xnor U16111 (N_16111,N_14583,N_14188);
nand U16112 (N_16112,N_14099,N_15110);
nand U16113 (N_16113,N_13983,N_13635);
nand U16114 (N_16114,N_12569,N_13379);
nand U16115 (N_16115,N_13028,N_12909);
xor U16116 (N_16116,N_13896,N_12933);
and U16117 (N_16117,N_13394,N_15376);
nor U16118 (N_16118,N_12897,N_14430);
nor U16119 (N_16119,N_15107,N_13487);
nand U16120 (N_16120,N_13412,N_13262);
nor U16121 (N_16121,N_13722,N_13727);
and U16122 (N_16122,N_13711,N_15580);
and U16123 (N_16123,N_14174,N_13200);
and U16124 (N_16124,N_14341,N_14355);
or U16125 (N_16125,N_13268,N_14517);
xnor U16126 (N_16126,N_13843,N_14356);
and U16127 (N_16127,N_14409,N_15264);
nand U16128 (N_16128,N_14790,N_13346);
nor U16129 (N_16129,N_12867,N_13385);
and U16130 (N_16130,N_14032,N_13398);
nand U16131 (N_16131,N_14777,N_13114);
xor U16132 (N_16132,N_13795,N_14200);
nor U16133 (N_16133,N_13764,N_14518);
nor U16134 (N_16134,N_13817,N_14951);
or U16135 (N_16135,N_12965,N_14904);
and U16136 (N_16136,N_15220,N_12610);
nor U16137 (N_16137,N_12796,N_12845);
nand U16138 (N_16138,N_13548,N_12825);
nand U16139 (N_16139,N_14908,N_13428);
and U16140 (N_16140,N_13696,N_14299);
xor U16141 (N_16141,N_15194,N_14794);
and U16142 (N_16142,N_14549,N_13246);
xnor U16143 (N_16143,N_12652,N_13167);
nand U16144 (N_16144,N_12533,N_12742);
or U16145 (N_16145,N_14412,N_13625);
nand U16146 (N_16146,N_15442,N_13811);
xor U16147 (N_16147,N_14201,N_13413);
xor U16148 (N_16148,N_15080,N_12839);
xor U16149 (N_16149,N_15321,N_14916);
nand U16150 (N_16150,N_15161,N_15046);
and U16151 (N_16151,N_14862,N_15410);
nand U16152 (N_16152,N_13705,N_14653);
nor U16153 (N_16153,N_13952,N_14171);
nor U16154 (N_16154,N_15575,N_13968);
and U16155 (N_16155,N_14477,N_13942);
nand U16156 (N_16156,N_14160,N_14504);
nand U16157 (N_16157,N_13493,N_13152);
xor U16158 (N_16158,N_12660,N_14535);
xnor U16159 (N_16159,N_12921,N_13355);
xor U16160 (N_16160,N_14330,N_15488);
nor U16161 (N_16161,N_14192,N_13690);
and U16162 (N_16162,N_13276,N_13852);
xnor U16163 (N_16163,N_15090,N_12765);
nand U16164 (N_16164,N_13056,N_13058);
or U16165 (N_16165,N_15539,N_12718);
nand U16166 (N_16166,N_13701,N_12739);
nor U16167 (N_16167,N_14153,N_15447);
xnor U16168 (N_16168,N_15594,N_14725);
or U16169 (N_16169,N_12687,N_12924);
nand U16170 (N_16170,N_12616,N_13273);
xor U16171 (N_16171,N_15612,N_12574);
and U16172 (N_16172,N_14941,N_13603);
and U16173 (N_16173,N_13104,N_14446);
or U16174 (N_16174,N_15475,N_12553);
nor U16175 (N_16175,N_13218,N_14632);
and U16176 (N_16176,N_13021,N_15471);
nor U16177 (N_16177,N_15414,N_14065);
or U16178 (N_16178,N_15048,N_15144);
or U16179 (N_16179,N_13007,N_14432);
or U16180 (N_16180,N_15566,N_14101);
and U16181 (N_16181,N_15339,N_12726);
and U16182 (N_16182,N_14963,N_13040);
or U16183 (N_16183,N_14403,N_13619);
and U16184 (N_16184,N_14241,N_12600);
nand U16185 (N_16185,N_13155,N_15067);
or U16186 (N_16186,N_14394,N_12665);
xor U16187 (N_16187,N_13480,N_12838);
xor U16188 (N_16188,N_12715,N_14888);
nor U16189 (N_16189,N_13496,N_13434);
and U16190 (N_16190,N_15130,N_12970);
or U16191 (N_16191,N_13148,N_13748);
nor U16192 (N_16192,N_15109,N_15016);
nand U16193 (N_16193,N_12877,N_12606);
nand U16194 (N_16194,N_12955,N_12657);
or U16195 (N_16195,N_12554,N_15173);
and U16196 (N_16196,N_15235,N_15306);
nor U16197 (N_16197,N_12622,N_13486);
and U16198 (N_16198,N_14376,N_15390);
and U16199 (N_16199,N_15398,N_15247);
xnor U16200 (N_16200,N_14636,N_15423);
and U16201 (N_16201,N_12595,N_12866);
xor U16202 (N_16202,N_14691,N_14868);
nor U16203 (N_16203,N_13261,N_14808);
or U16204 (N_16204,N_14110,N_12826);
or U16205 (N_16205,N_15516,N_13913);
xor U16206 (N_16206,N_15546,N_13151);
or U16207 (N_16207,N_12663,N_13421);
and U16208 (N_16208,N_14831,N_15371);
or U16209 (N_16209,N_13255,N_13849);
nand U16210 (N_16210,N_14552,N_12514);
xor U16211 (N_16211,N_14869,N_15526);
and U16212 (N_16212,N_15584,N_13675);
nand U16213 (N_16213,N_14751,N_14287);
and U16214 (N_16214,N_14717,N_14727);
and U16215 (N_16215,N_13857,N_13776);
nand U16216 (N_16216,N_15542,N_12768);
nand U16217 (N_16217,N_15120,N_13030);
or U16218 (N_16218,N_15498,N_13124);
nand U16219 (N_16219,N_13791,N_14193);
nor U16220 (N_16220,N_14143,N_15047);
nand U16221 (N_16221,N_15399,N_12584);
nand U16222 (N_16222,N_14347,N_13303);
nor U16223 (N_16223,N_13184,N_15509);
or U16224 (N_16224,N_13378,N_14498);
nor U16225 (N_16225,N_13110,N_14071);
xnor U16226 (N_16226,N_15394,N_12806);
nor U16227 (N_16227,N_13556,N_13752);
xnor U16228 (N_16228,N_13741,N_14891);
xnor U16229 (N_16229,N_15511,N_15478);
and U16230 (N_16230,N_13777,N_13479);
xnor U16231 (N_16231,N_12850,N_15164);
and U16232 (N_16232,N_14182,N_15010);
nand U16233 (N_16233,N_14169,N_15039);
or U16234 (N_16234,N_13367,N_13819);
nand U16235 (N_16235,N_14607,N_14137);
or U16236 (N_16236,N_15154,N_13636);
nand U16237 (N_16237,N_12749,N_12697);
xor U16238 (N_16238,N_15615,N_13914);
and U16239 (N_16239,N_13236,N_14741);
xnor U16240 (N_16240,N_15284,N_14055);
or U16241 (N_16241,N_12631,N_13622);
xnor U16242 (N_16242,N_12744,N_13213);
and U16243 (N_16243,N_15049,N_15072);
nor U16244 (N_16244,N_13455,N_13518);
nor U16245 (N_16245,N_13012,N_14846);
xor U16246 (N_16246,N_14493,N_12777);
or U16247 (N_16247,N_13336,N_14115);
nand U16248 (N_16248,N_14113,N_12939);
or U16249 (N_16249,N_15582,N_14810);
and U16250 (N_16250,N_13880,N_13601);
and U16251 (N_16251,N_15452,N_14146);
and U16252 (N_16252,N_13157,N_13388);
xor U16253 (N_16253,N_14827,N_13981);
nand U16254 (N_16254,N_14131,N_13918);
nor U16255 (N_16255,N_14952,N_12940);
and U16256 (N_16256,N_13089,N_15029);
xor U16257 (N_16257,N_13782,N_15257);
nand U16258 (N_16258,N_14033,N_14263);
and U16259 (N_16259,N_13219,N_14002);
xnor U16260 (N_16260,N_12983,N_15005);
or U16261 (N_16261,N_12670,N_13600);
nand U16262 (N_16262,N_13300,N_14942);
or U16263 (N_16263,N_14264,N_14540);
nand U16264 (N_16264,N_15327,N_14989);
nand U16265 (N_16265,N_14129,N_14515);
nand U16266 (N_16266,N_14852,N_15166);
and U16267 (N_16267,N_14453,N_14739);
and U16268 (N_16268,N_13576,N_13637);
or U16269 (N_16269,N_14417,N_13994);
nand U16270 (N_16270,N_14428,N_13465);
xor U16271 (N_16271,N_13371,N_13985);
xnor U16272 (N_16272,N_15438,N_13471);
or U16273 (N_16273,N_12578,N_14781);
nor U16274 (N_16274,N_15347,N_13584);
nand U16275 (N_16275,N_14133,N_15324);
nor U16276 (N_16276,N_15230,N_14948);
nor U16277 (N_16277,N_13502,N_15551);
xnor U16278 (N_16278,N_14416,N_15026);
or U16279 (N_16279,N_14981,N_15032);
and U16280 (N_16280,N_15126,N_14551);
and U16281 (N_16281,N_12830,N_15315);
nor U16282 (N_16282,N_12646,N_14731);
nor U16283 (N_16283,N_15134,N_13538);
nor U16284 (N_16284,N_14242,N_15270);
or U16285 (N_16285,N_13940,N_14424);
xor U16286 (N_16286,N_15504,N_12764);
nand U16287 (N_16287,N_14721,N_13788);
nand U16288 (N_16288,N_14976,N_13315);
xnor U16289 (N_16289,N_15204,N_14211);
and U16290 (N_16290,N_12904,N_13972);
nand U16291 (N_16291,N_13865,N_14687);
or U16292 (N_16292,N_13984,N_13054);
xor U16293 (N_16293,N_13204,N_14579);
xor U16294 (N_16294,N_13014,N_14813);
xnor U16295 (N_16295,N_13327,N_13834);
and U16296 (N_16296,N_14420,N_14734);
nand U16297 (N_16297,N_13435,N_14191);
xor U16298 (N_16298,N_14469,N_12949);
and U16299 (N_16299,N_12524,N_13506);
nand U16300 (N_16300,N_14323,N_14111);
nor U16301 (N_16301,N_15609,N_12716);
xor U16302 (N_16302,N_13947,N_13042);
xor U16303 (N_16303,N_15083,N_14818);
nand U16304 (N_16304,N_15574,N_15603);
nor U16305 (N_16305,N_14121,N_14648);
and U16306 (N_16306,N_13020,N_15231);
and U16307 (N_16307,N_13440,N_13095);
nor U16308 (N_16308,N_14392,N_14094);
nand U16309 (N_16309,N_13900,N_13763);
nor U16310 (N_16310,N_14576,N_15226);
or U16311 (N_16311,N_13019,N_15379);
and U16312 (N_16312,N_14825,N_13350);
and U16313 (N_16313,N_13965,N_15530);
or U16314 (N_16314,N_14608,N_14239);
or U16315 (N_16315,N_13612,N_14389);
nor U16316 (N_16316,N_14617,N_13846);
xor U16317 (N_16317,N_13441,N_15556);
nor U16318 (N_16318,N_13820,N_14738);
and U16319 (N_16319,N_12863,N_14291);
xnor U16320 (N_16320,N_14373,N_12951);
xor U16321 (N_16321,N_15318,N_14761);
nor U16322 (N_16322,N_13096,N_15508);
xor U16323 (N_16323,N_13340,N_14710);
nor U16324 (N_16324,N_12500,N_13768);
or U16325 (N_16325,N_14255,N_14695);
or U16326 (N_16326,N_13400,N_13762);
and U16327 (N_16327,N_14197,N_13511);
nand U16328 (N_16328,N_13587,N_14589);
or U16329 (N_16329,N_15333,N_12591);
nand U16330 (N_16330,N_15178,N_13772);
nor U16331 (N_16331,N_14899,N_15606);
nand U16332 (N_16332,N_12732,N_14350);
or U16333 (N_16333,N_14380,N_14050);
xnor U16334 (N_16334,N_14595,N_13025);
xnor U16335 (N_16335,N_15421,N_13404);
xnor U16336 (N_16336,N_14503,N_14621);
or U16337 (N_16337,N_13065,N_12859);
and U16338 (N_16338,N_14949,N_14229);
xnor U16339 (N_16339,N_13048,N_14140);
and U16340 (N_16340,N_12792,N_13494);
xnor U16341 (N_16341,N_15087,N_14596);
and U16342 (N_16342,N_12656,N_15331);
or U16343 (N_16343,N_13106,N_13508);
nand U16344 (N_16344,N_15518,N_14163);
nor U16345 (N_16345,N_13531,N_12751);
xnor U16346 (N_16346,N_14048,N_13011);
or U16347 (N_16347,N_13205,N_15486);
and U16348 (N_16348,N_15062,N_14853);
xor U16349 (N_16349,N_14685,N_13754);
and U16350 (N_16350,N_13243,N_13784);
and U16351 (N_16351,N_14971,N_15176);
or U16352 (N_16352,N_15037,N_13382);
nor U16353 (N_16353,N_15024,N_12750);
nor U16354 (N_16354,N_15537,N_15068);
nor U16355 (N_16355,N_14510,N_13879);
nand U16356 (N_16356,N_15377,N_12589);
and U16357 (N_16357,N_15497,N_13432);
nor U16358 (N_16358,N_13597,N_12775);
nand U16359 (N_16359,N_14920,N_14296);
or U16360 (N_16360,N_13668,N_13700);
nand U16361 (N_16361,N_15329,N_12693);
and U16362 (N_16362,N_12723,N_13962);
and U16363 (N_16363,N_12808,N_13424);
nand U16364 (N_16364,N_12623,N_13396);
or U16365 (N_16365,N_14729,N_14353);
and U16366 (N_16366,N_14574,N_14454);
nor U16367 (N_16367,N_13809,N_15300);
nand U16368 (N_16368,N_15449,N_13431);
or U16369 (N_16369,N_12535,N_13789);
nor U16370 (N_16370,N_14927,N_15527);
or U16371 (N_16371,N_12651,N_14418);
xnor U16372 (N_16372,N_12786,N_13363);
or U16373 (N_16373,N_14067,N_14774);
and U16374 (N_16374,N_15310,N_15283);
nand U16375 (N_16375,N_15198,N_12519);
xor U16376 (N_16376,N_14702,N_13333);
xnor U16377 (N_16377,N_13685,N_14106);
nor U16378 (N_16378,N_15070,N_15457);
or U16379 (N_16379,N_14305,N_12549);
nor U16380 (N_16380,N_13825,N_13469);
xor U16381 (N_16381,N_14322,N_13568);
xnor U16382 (N_16382,N_14021,N_13464);
xor U16383 (N_16383,N_13159,N_15169);
nor U16384 (N_16384,N_13670,N_12936);
xor U16385 (N_16385,N_14760,N_14144);
or U16386 (N_16386,N_13855,N_13374);
nor U16387 (N_16387,N_15622,N_13483);
and U16388 (N_16388,N_13009,N_13472);
or U16389 (N_16389,N_14368,N_14072);
and U16390 (N_16390,N_13644,N_15261);
and U16391 (N_16391,N_14349,N_14052);
xor U16392 (N_16392,N_13256,N_12573);
xnor U16393 (N_16393,N_13005,N_14180);
and U16394 (N_16394,N_15587,N_12773);
and U16395 (N_16395,N_15105,N_15215);
xnor U16396 (N_16396,N_14117,N_15063);
and U16397 (N_16397,N_14284,N_15145);
or U16398 (N_16398,N_14185,N_13992);
nand U16399 (N_16399,N_13376,N_15491);
nand U16400 (N_16400,N_14536,N_13695);
or U16401 (N_16401,N_15102,N_14913);
and U16402 (N_16402,N_14560,N_13990);
nand U16403 (N_16403,N_13131,N_13996);
nor U16404 (N_16404,N_14719,N_14625);
and U16405 (N_16405,N_12982,N_14605);
or U16406 (N_16406,N_12731,N_15369);
nor U16407 (N_16407,N_15158,N_14892);
xnor U16408 (N_16408,N_14795,N_13373);
or U16409 (N_16409,N_13233,N_14838);
xor U16410 (N_16410,N_13485,N_14964);
nor U16411 (N_16411,N_15484,N_13669);
nor U16412 (N_16412,N_15623,N_13063);
or U16413 (N_16413,N_12894,N_14338);
or U16414 (N_16414,N_13169,N_13514);
xor U16415 (N_16415,N_14026,N_13523);
and U16416 (N_16416,N_13976,N_13596);
nor U16417 (N_16417,N_13482,N_15568);
or U16418 (N_16418,N_13239,N_13179);
and U16419 (N_16419,N_14987,N_14802);
or U16420 (N_16420,N_14372,N_12597);
and U16421 (N_16421,N_13580,N_15561);
and U16422 (N_16422,N_15170,N_12762);
or U16423 (N_16423,N_14364,N_14164);
nor U16424 (N_16424,N_14120,N_15030);
nand U16425 (N_16425,N_14584,N_14896);
or U16426 (N_16426,N_12539,N_13935);
xor U16427 (N_16427,N_12853,N_13384);
or U16428 (N_16428,N_13168,N_14290);
and U16429 (N_16429,N_12922,N_15432);
or U16430 (N_16430,N_13715,N_14228);
nand U16431 (N_16431,N_15439,N_12803);
nand U16432 (N_16432,N_15366,N_13723);
or U16433 (N_16433,N_14190,N_14088);
nand U16434 (N_16434,N_12710,N_15469);
and U16435 (N_16435,N_13746,N_13334);
xor U16436 (N_16436,N_14619,N_13877);
and U16437 (N_16437,N_13841,N_14967);
xor U16438 (N_16438,N_13186,N_14357);
and U16439 (N_16439,N_15147,N_12996);
and U16440 (N_16440,N_12857,N_14468);
nand U16441 (N_16441,N_15237,N_15222);
or U16442 (N_16442,N_14945,N_13813);
and U16443 (N_16443,N_13740,N_15600);
xor U16444 (N_16444,N_13611,N_13050);
nand U16445 (N_16445,N_15429,N_13901);
or U16446 (N_16446,N_15445,N_13111);
or U16447 (N_16447,N_15294,N_14170);
nor U16448 (N_16448,N_15564,N_14793);
or U16449 (N_16449,N_13445,N_14485);
nand U16450 (N_16450,N_13370,N_13317);
or U16451 (N_16451,N_12813,N_13446);
and U16452 (N_16452,N_13426,N_14419);
or U16453 (N_16453,N_13301,N_15057);
and U16454 (N_16454,N_14706,N_13515);
nand U16455 (N_16455,N_13773,N_12717);
or U16456 (N_16456,N_15373,N_13375);
or U16457 (N_16457,N_13033,N_12783);
or U16458 (N_16458,N_13799,N_14585);
xor U16459 (N_16459,N_14826,N_14936);
xnor U16460 (N_16460,N_14301,N_13326);
xnor U16461 (N_16461,N_13979,N_13766);
or U16462 (N_16462,N_12644,N_12754);
nand U16463 (N_16463,N_14915,N_14620);
nand U16464 (N_16464,N_15289,N_12727);
nor U16465 (N_16465,N_13150,N_14953);
or U16466 (N_16466,N_14324,N_14162);
and U16467 (N_16467,N_14860,N_15108);
and U16468 (N_16468,N_13041,N_14078);
nor U16469 (N_16469,N_15055,N_15352);
or U16470 (N_16470,N_12964,N_15360);
nor U16471 (N_16471,N_15416,N_13241);
xor U16472 (N_16472,N_14262,N_14235);
nor U16473 (N_16473,N_13174,N_13999);
or U16474 (N_16474,N_13228,N_14699);
nand U16475 (N_16475,N_14962,N_15567);
or U16476 (N_16476,N_14837,N_14256);
nand U16477 (N_16477,N_12989,N_12780);
nand U16478 (N_16478,N_13663,N_14726);
nand U16479 (N_16479,N_13499,N_14232);
or U16480 (N_16480,N_14779,N_15468);
and U16481 (N_16481,N_13598,N_14488);
nor U16482 (N_16482,N_12801,N_15374);
xor U16483 (N_16483,N_15249,N_15499);
nor U16484 (N_16484,N_14815,N_13800);
nand U16485 (N_16485,N_14849,N_15586);
or U16486 (N_16486,N_15505,N_13242);
and U16487 (N_16487,N_14850,N_13027);
xnor U16488 (N_16488,N_13838,N_13490);
xnor U16489 (N_16489,N_13894,N_13223);
xnor U16490 (N_16490,N_12628,N_12874);
and U16491 (N_16491,N_14787,N_14597);
nor U16492 (N_16492,N_14628,N_15207);
nand U16493 (N_16493,N_14415,N_12599);
nor U16494 (N_16494,N_14363,N_15483);
nand U16495 (N_16495,N_14159,N_13093);
or U16496 (N_16496,N_14481,N_13456);
nand U16497 (N_16497,N_14609,N_14361);
nor U16498 (N_16498,N_12911,N_15506);
xnor U16499 (N_16499,N_13283,N_14894);
xnor U16500 (N_16500,N_13416,N_14775);
xnor U16501 (N_16501,N_15314,N_15454);
and U16502 (N_16502,N_15036,N_12582);
and U16503 (N_16503,N_14307,N_12607);
nor U16504 (N_16504,N_15239,N_15160);
and U16505 (N_16505,N_14247,N_14240);
xor U16506 (N_16506,N_12729,N_13831);
nor U16507 (N_16507,N_14782,N_15099);
and U16508 (N_16508,N_13673,N_14829);
nand U16509 (N_16509,N_15391,N_12875);
or U16510 (N_16510,N_14083,N_14205);
nor U16511 (N_16511,N_12577,N_12907);
nor U16512 (N_16512,N_14759,N_12931);
or U16513 (N_16513,N_15358,N_13120);
or U16514 (N_16514,N_14752,N_12998);
xnor U16515 (N_16515,N_13530,N_15558);
nor U16516 (N_16516,N_13563,N_14207);
xor U16517 (N_16517,N_15593,N_14045);
and U16518 (N_16518,N_13458,N_14889);
xor U16519 (N_16519,N_14610,N_13158);
and U16520 (N_16520,N_14929,N_15559);
xor U16521 (N_16521,N_13953,N_14615);
xor U16522 (N_16522,N_12529,N_13904);
and U16523 (N_16523,N_13977,N_14273);
xnor U16524 (N_16524,N_13162,N_14934);
and U16525 (N_16525,N_12680,N_13588);
nor U16526 (N_16526,N_14921,N_12505);
nand U16527 (N_16527,N_13975,N_13554);
or U16528 (N_16528,N_15223,N_14172);
nor U16529 (N_16529,N_14784,N_13541);
or U16530 (N_16530,N_15382,N_15050);
nor U16531 (N_16531,N_15521,N_13190);
xor U16532 (N_16532,N_12854,N_15386);
or U16533 (N_16533,N_13757,N_14025);
or U16534 (N_16534,N_13402,N_13196);
or U16535 (N_16535,N_12967,N_14992);
and U16536 (N_16536,N_12563,N_13491);
nand U16537 (N_16537,N_15297,N_13778);
or U16538 (N_16538,N_13995,N_13332);
nor U16539 (N_16539,N_12994,N_13342);
or U16540 (N_16540,N_13039,N_12828);
xnor U16541 (N_16541,N_14219,N_14606);
and U16542 (N_16542,N_12797,N_14480);
or U16543 (N_16543,N_13149,N_14145);
xor U16544 (N_16544,N_12774,N_13535);
nor U16545 (N_16545,N_13532,N_13209);
nand U16546 (N_16546,N_13874,N_14712);
and U16547 (N_16547,N_15319,N_15201);
nand U16548 (N_16548,N_12829,N_14049);
nand U16549 (N_16549,N_15172,N_13534);
nor U16550 (N_16550,N_12858,N_13092);
xor U16551 (N_16551,N_14800,N_13214);
and U16552 (N_16552,N_15565,N_15302);
and U16553 (N_16553,N_14823,N_14656);
nor U16554 (N_16554,N_13509,N_13797);
or U16555 (N_16555,N_13986,N_14270);
or U16556 (N_16556,N_15443,N_12641);
xnor U16557 (N_16557,N_13839,N_13826);
xnor U16558 (N_16558,N_13703,N_13068);
and U16559 (N_16559,N_12794,N_14105);
or U16560 (N_16560,N_14737,N_15599);
xnor U16561 (N_16561,N_14339,N_15285);
nand U16562 (N_16562,N_14527,N_15512);
nand U16563 (N_16563,N_13565,N_12995);
nor U16564 (N_16564,N_15434,N_12590);
nor U16565 (N_16565,N_13666,N_13647);
and U16566 (N_16566,N_14176,N_12548);
nand U16567 (N_16567,N_13616,N_14755);
nand U16568 (N_16568,N_14031,N_15388);
and U16569 (N_16569,N_14968,N_14402);
or U16570 (N_16570,N_13924,N_13832);
nand U16571 (N_16571,N_14848,N_15301);
nor U16572 (N_16572,N_14834,N_14385);
and U16573 (N_16573,N_14939,N_13858);
xor U16574 (N_16574,N_12507,N_15293);
nand U16575 (N_16575,N_12741,N_13887);
or U16576 (N_16576,N_14500,N_15430);
xnor U16577 (N_16577,N_13178,N_13987);
or U16578 (N_16578,N_15415,N_14545);
nand U16579 (N_16579,N_12630,N_15348);
or U16580 (N_16580,N_13549,N_14028);
and U16581 (N_16581,N_13249,N_12818);
nor U16582 (N_16582,N_13381,N_14059);
nor U16583 (N_16583,N_13387,N_12862);
or U16584 (N_16584,N_14214,N_14893);
nand U16585 (N_16585,N_12627,N_12869);
nor U16586 (N_16586,N_13944,N_14565);
or U16587 (N_16587,N_14773,N_12840);
or U16588 (N_16588,N_12706,N_13229);
nor U16589 (N_16589,N_13052,N_12707);
and U16590 (N_16590,N_15004,N_15591);
nand U16591 (N_16591,N_13599,N_14039);
or U16592 (N_16592,N_13253,N_13793);
nand U16593 (N_16593,N_14104,N_14508);
and U16594 (N_16594,N_15066,N_13743);
nor U16595 (N_16595,N_14306,N_13306);
xor U16596 (N_16596,N_15094,N_14359);
xor U16597 (N_16597,N_14400,N_13070);
and U16598 (N_16598,N_14582,N_14678);
nand U16599 (N_16599,N_14375,N_14494);
nor U16600 (N_16600,N_15150,N_14011);
nand U16601 (N_16601,N_15608,N_14705);
nand U16602 (N_16602,N_15100,N_14922);
nand U16603 (N_16603,N_13557,N_12988);
and U16604 (N_16604,N_14988,N_13489);
or U16605 (N_16605,N_13997,N_14489);
and U16606 (N_16606,N_14586,N_14856);
and U16607 (N_16607,N_15103,N_15387);
xnor U16608 (N_16608,N_13830,N_13232);
and U16609 (N_16609,N_13744,N_13926);
or U16610 (N_16610,N_13654,N_14561);
nand U16611 (N_16611,N_13047,N_15308);
xnor U16612 (N_16612,N_15267,N_14547);
nand U16613 (N_16613,N_13429,N_14184);
or U16614 (N_16614,N_15465,N_13015);
and U16615 (N_16615,N_15031,N_13551);
xnor U16616 (N_16616,N_14566,N_15193);
or U16617 (N_16617,N_14788,N_15095);
or U16618 (N_16618,N_12976,N_14906);
and U16619 (N_16619,N_13488,N_14558);
nand U16620 (N_16620,N_13079,N_14069);
or U16621 (N_16621,N_13277,N_13796);
nand U16622 (N_16622,N_13034,N_14073);
nor U16623 (N_16623,N_12787,N_14878);
or U16624 (N_16624,N_14023,N_12968);
nand U16625 (N_16625,N_13955,N_13197);
and U16626 (N_16626,N_13353,N_14202);
nand U16627 (N_16627,N_12690,N_15474);
and U16628 (N_16628,N_14785,N_14022);
xor U16629 (N_16629,N_13908,N_13078);
and U16630 (N_16630,N_13194,N_15541);
nor U16631 (N_16631,N_14474,N_14747);
xnor U16632 (N_16632,N_15549,N_14666);
xnor U16633 (N_16633,N_14340,N_13299);
nor U16634 (N_16634,N_12925,N_14577);
nand U16635 (N_16635,N_13691,N_14443);
nand U16636 (N_16636,N_15589,N_15128);
or U16637 (N_16637,N_14635,N_12685);
and U16638 (N_16638,N_12973,N_14954);
and U16639 (N_16639,N_14124,N_12506);
nand U16640 (N_16640,N_13002,N_15616);
nand U16641 (N_16641,N_14932,N_13364);
or U16642 (N_16642,N_13623,N_15520);
nor U16643 (N_16643,N_12819,N_15550);
or U16644 (N_16644,N_14555,N_14054);
xnor U16645 (N_16645,N_14940,N_14194);
nand U16646 (N_16646,N_15547,N_15041);
and U16647 (N_16647,N_13689,N_14455);
nor U16648 (N_16648,N_15191,N_15363);
nor U16649 (N_16649,N_13098,N_12928);
nand U16650 (N_16650,N_14075,N_13195);
and U16651 (N_16651,N_14395,N_14646);
nor U16652 (N_16652,N_13438,N_15271);
nand U16653 (N_16653,N_12733,N_14564);
xnor U16654 (N_16654,N_12604,N_13803);
and U16655 (N_16655,N_13208,N_14152);
or U16656 (N_16656,N_15114,N_12748);
or U16657 (N_16657,N_15045,N_14533);
or U16658 (N_16658,N_13461,N_13127);
nand U16659 (N_16659,N_13624,N_12503);
nand U16660 (N_16660,N_12538,N_12547);
and U16661 (N_16661,N_13956,N_14265);
xor U16662 (N_16662,N_13442,N_12878);
xor U16663 (N_16663,N_14058,N_12552);
and U16664 (N_16664,N_14970,N_14379);
nand U16665 (N_16665,N_14876,N_12941);
or U16666 (N_16666,N_14461,N_12821);
nand U16667 (N_16667,N_12585,N_13714);
and U16668 (N_16668,N_12605,N_12865);
nand U16669 (N_16669,N_14512,N_13278);
nand U16670 (N_16670,N_13395,N_14634);
or U16671 (N_16671,N_15492,N_13961);
nor U16672 (N_16672,N_14177,N_12612);
nand U16673 (N_16673,N_14765,N_14000);
nand U16674 (N_16674,N_13680,N_13386);
or U16675 (N_16675,N_15418,N_12704);
xnor U16676 (N_16676,N_13787,N_12537);
nand U16677 (N_16677,N_14405,N_14458);
xnor U16678 (N_16678,N_13758,N_15106);
and U16679 (N_16679,N_15522,N_13447);
or U16680 (N_16680,N_13225,N_14864);
and U16681 (N_16681,N_12881,N_15197);
and U16682 (N_16682,N_14010,N_13677);
nand U16683 (N_16683,N_15135,N_14450);
xor U16684 (N_16684,N_14841,N_13144);
xor U16685 (N_16685,N_15501,N_14723);
and U16686 (N_16686,N_14429,N_15427);
or U16687 (N_16687,N_15292,N_14342);
nor U16688 (N_16688,N_14733,N_15325);
and U16689 (N_16689,N_13365,N_15286);
or U16690 (N_16690,N_13674,N_12822);
and U16691 (N_16691,N_15081,N_15529);
nor U16692 (N_16692,N_13181,N_15058);
nor U16693 (N_16693,N_15132,N_13310);
nand U16694 (N_16694,N_13630,N_12601);
or U16695 (N_16695,N_12621,N_15242);
nor U16696 (N_16696,N_15476,N_15407);
and U16697 (N_16697,N_15035,N_15490);
xnor U16698 (N_16698,N_15078,N_13166);
xor U16699 (N_16699,N_15614,N_14130);
nor U16700 (N_16700,N_14931,N_14128);
xnor U16701 (N_16701,N_13207,N_14449);
xnor U16702 (N_16702,N_14956,N_15018);
xor U16703 (N_16703,N_15304,N_12561);
and U16704 (N_16704,N_14623,N_12540);
xor U16705 (N_16705,N_15098,N_15409);
or U16706 (N_16706,N_13683,N_15266);
nand U16707 (N_16707,N_14107,N_14289);
and U16708 (N_16708,N_15448,N_14581);
and U16709 (N_16709,N_14681,N_13076);
and U16710 (N_16710,N_14631,N_14470);
xnor U16711 (N_16711,N_12640,N_12645);
nor U16712 (N_16712,N_15053,N_14114);
and U16713 (N_16713,N_15006,N_12515);
nor U16714 (N_16714,N_13812,N_12836);
and U16715 (N_16715,N_14554,N_13171);
xor U16716 (N_16716,N_12817,N_15060);
and U16717 (N_16717,N_14707,N_14008);
nor U16718 (N_16718,N_13477,N_15493);
nor U16719 (N_16719,N_15357,N_13059);
xnor U16720 (N_16720,N_14221,N_15186);
nand U16721 (N_16721,N_14413,N_14649);
or U16722 (N_16722,N_14248,N_13875);
or U16723 (N_16723,N_15021,N_13888);
and U16724 (N_16724,N_14064,N_12719);
nor U16725 (N_16725,N_15288,N_14277);
nor U16726 (N_16726,N_13201,N_13417);
xnor U16727 (N_16727,N_13272,N_14300);
xor U16728 (N_16728,N_13943,N_14125);
and U16729 (N_16729,N_13094,N_14274);
or U16730 (N_16730,N_12852,N_14677);
nand U16731 (N_16731,N_12649,N_14686);
xor U16732 (N_16732,N_14662,N_14148);
xor U16733 (N_16733,N_14123,N_13304);
or U16734 (N_16734,N_13765,N_15084);
or U16735 (N_16735,N_15137,N_15507);
nor U16736 (N_16736,N_15232,N_12889);
or U16737 (N_16737,N_12809,N_13516);
and U16738 (N_16738,N_13119,N_12887);
nand U16739 (N_16739,N_13308,N_13958);
and U16740 (N_16740,N_12603,N_14655);
or U16741 (N_16741,N_12575,N_13305);
xor U16742 (N_16742,N_13088,N_15017);
nand U16743 (N_16743,N_15515,N_12946);
or U16744 (N_16744,N_12724,N_12778);
or U16745 (N_16745,N_13356,N_15217);
nor U16746 (N_16746,N_14791,N_13128);
nor U16747 (N_16747,N_14492,N_12902);
or U16748 (N_16748,N_14780,N_14642);
nand U16749 (N_16749,N_15203,N_12978);
or U16750 (N_16750,N_15479,N_15256);
or U16751 (N_16751,N_14855,N_14756);
nand U16752 (N_16752,N_14245,N_12832);
or U16753 (N_16753,N_13123,N_14495);
or U16754 (N_16754,N_13302,N_14286);
nor U16755 (N_16755,N_15337,N_13617);
nand U16756 (N_16756,N_14427,N_12798);
nand U16757 (N_16757,N_13240,N_15245);
xor U16758 (N_16758,N_15406,N_13927);
nor U16759 (N_16759,N_12705,N_15190);
nand U16760 (N_16760,N_14486,N_14528);
nor U16761 (N_16761,N_15316,N_15116);
xor U16762 (N_16762,N_15553,N_12816);
xor U16763 (N_16763,N_14321,N_13319);
xor U16764 (N_16764,N_15251,N_14328);
nor U16765 (N_16765,N_13248,N_15019);
or U16766 (N_16766,N_12722,N_13462);
or U16767 (N_16767,N_15510,N_14410);
or U16768 (N_16768,N_13164,N_14740);
and U16769 (N_16769,N_13967,N_14015);
and U16770 (N_16770,N_14757,N_12674);
xnor U16771 (N_16771,N_14633,N_13180);
xnor U16772 (N_16772,N_13314,N_13739);
or U16773 (N_16773,N_12508,N_14465);
nand U16774 (N_16774,N_13665,N_13116);
or U16775 (N_16775,N_12737,N_12617);
nor U16776 (N_16776,N_14079,N_14543);
nand U16777 (N_16777,N_13220,N_13543);
nor U16778 (N_16778,N_14027,N_15131);
and U16779 (N_16779,N_13418,N_14366);
nor U16780 (N_16780,N_14645,N_14007);
xor U16781 (N_16781,N_13282,N_14534);
nand U16782 (N_16782,N_12980,N_13821);
nand U16783 (N_16783,N_14651,N_14882);
nand U16784 (N_16784,N_12984,N_13524);
or U16785 (N_16785,N_15500,N_14613);
or U16786 (N_16786,N_15496,N_13425);
and U16787 (N_16787,N_14087,N_14716);
nor U16788 (N_16788,N_15353,N_14313);
nor U16789 (N_16789,N_12846,N_14769);
and U16790 (N_16790,N_12791,N_15168);
nor U16791 (N_16791,N_13915,N_15340);
nor U16792 (N_16792,N_14943,N_15069);
nor U16793 (N_16793,N_14903,N_14294);
nand U16794 (N_16794,N_14995,N_12654);
and U16795 (N_16795,N_13938,N_12885);
and U16796 (N_16796,N_13640,N_13605);
and U16797 (N_16797,N_14820,N_14238);
or U16798 (N_16798,N_12620,N_13247);
nor U16799 (N_16799,N_13737,N_13844);
or U16800 (N_16800,N_14771,N_15007);
nor U16801 (N_16801,N_12725,N_13064);
nand U16802 (N_16802,N_13357,N_15124);
xnor U16803 (N_16803,N_14592,N_14713);
and U16804 (N_16804,N_12771,N_15295);
or U16805 (N_16805,N_14870,N_12849);
nand U16806 (N_16806,N_12637,N_14996);
xor U16807 (N_16807,N_14149,N_13252);
and U16808 (N_16808,N_14288,N_13719);
nand U16809 (N_16809,N_12523,N_13215);
nand U16810 (N_16810,N_13453,N_13583);
nand U16811 (N_16811,N_13399,N_14796);
xnor U16812 (N_16812,N_12917,N_14283);
or U16813 (N_16813,N_14832,N_13552);
and U16814 (N_16814,N_13080,N_12831);
nor U16815 (N_16815,N_13053,N_13369);
xor U16816 (N_16816,N_15525,N_14399);
xnor U16817 (N_16817,N_12827,N_14017);
or U16818 (N_16818,N_14362,N_14590);
nor U16819 (N_16819,N_14091,N_12712);
nor U16820 (N_16820,N_13718,N_12957);
or U16821 (N_16821,N_14521,N_12655);
or U16822 (N_16822,N_13140,N_14452);
nor U16823 (N_16823,N_12614,N_13676);
or U16824 (N_16824,N_13522,N_15303);
or U16825 (N_16825,N_14917,N_13604);
or U16826 (N_16826,N_12918,N_12555);
or U16827 (N_16827,N_15383,N_13410);
xor U16828 (N_16828,N_13038,N_15086);
and U16829 (N_16829,N_14652,N_14425);
nor U16830 (N_16830,N_12738,N_14004);
and U16831 (N_16831,N_12947,N_13136);
nor U16832 (N_16832,N_15003,N_14659);
nand U16833 (N_16833,N_15092,N_14345);
or U16834 (N_16834,N_12864,N_12758);
or U16835 (N_16835,N_12669,N_15079);
nand U16836 (N_16836,N_14122,N_13824);
xnor U16837 (N_16837,N_13592,N_13260);
and U16838 (N_16838,N_14175,N_13946);
or U16839 (N_16839,N_12735,N_14990);
and U16840 (N_16840,N_13993,N_13517);
xnor U16841 (N_16841,N_14352,N_14601);
xor U16842 (N_16842,N_13893,N_12802);
xnor U16843 (N_16843,N_14614,N_13769);
nand U16844 (N_16844,N_14479,N_12913);
and U16845 (N_16845,N_15481,N_12785);
nor U16846 (N_16846,N_13536,N_13325);
or U16847 (N_16847,N_13836,N_15480);
or U16848 (N_16848,N_12823,N_12679);
and U16849 (N_16849,N_13107,N_12759);
nand U16850 (N_16850,N_13652,N_13495);
and U16851 (N_16851,N_13898,N_15189);
xnor U16852 (N_16852,N_13591,N_13589);
and U16853 (N_16853,N_15362,N_12734);
xnor U16854 (N_16854,N_15395,N_15260);
nor U16855 (N_16855,N_14036,N_15543);
or U16856 (N_16856,N_12587,N_14346);
or U16857 (N_16857,N_14600,N_15585);
xnor U16858 (N_16858,N_14154,N_13738);
xnor U16859 (N_16859,N_14252,N_14463);
and U16860 (N_16860,N_15536,N_14501);
nand U16861 (N_16861,N_14292,N_13183);
or U16862 (N_16862,N_15139,N_15143);
xor U16863 (N_16863,N_14550,N_12518);
nor U16864 (N_16864,N_14044,N_14704);
and U16865 (N_16865,N_13840,N_13921);
or U16866 (N_16866,N_14865,N_14447);
and U16867 (N_16867,N_15088,N_14390);
xnor U16868 (N_16868,N_15163,N_13188);
nor U16869 (N_16869,N_15258,N_14912);
and U16870 (N_16870,N_14772,N_12953);
or U16871 (N_16871,N_14799,N_14475);
nor U16872 (N_16872,N_13910,N_14975);
or U16873 (N_16873,N_14298,N_12542);
nor U16874 (N_16874,N_13594,N_14993);
or U16875 (N_16875,N_15061,N_15464);
xnor U16876 (N_16876,N_14743,N_12975);
nor U16877 (N_16877,N_14910,N_12509);
xor U16878 (N_16878,N_15441,N_13564);
nor U16879 (N_16879,N_13312,N_14532);
and U16880 (N_16880,N_15263,N_13289);
xor U16881 (N_16881,N_12776,N_14935);
nand U16882 (N_16882,N_15588,N_13202);
nand U16883 (N_16883,N_13571,N_14629);
xor U16884 (N_16884,N_14657,N_14066);
or U16885 (N_16885,N_13175,N_12527);
nand U16886 (N_16886,N_14696,N_14682);
nand U16887 (N_16887,N_15411,N_13437);
and U16888 (N_16888,N_13343,N_13016);
xor U16889 (N_16889,N_13112,N_13075);
nand U16890 (N_16890,N_13141,N_13537);
or U16891 (N_16891,N_15384,N_14701);
and U16892 (N_16892,N_14998,N_15356);
nand U16893 (N_16893,N_14746,N_14819);
nor U16894 (N_16894,N_14969,N_13756);
nand U16895 (N_16895,N_13436,N_15397);
nand U16896 (N_16896,N_14081,N_15350);
and U16897 (N_16897,N_13717,N_15317);
xor U16898 (N_16898,N_13716,N_13613);
nor U16899 (N_16899,N_13475,N_14714);
xor U16900 (N_16900,N_15071,N_12544);
nand U16901 (N_16901,N_13212,N_13912);
xnor U16902 (N_16902,N_13422,N_14315);
nor U16903 (N_16903,N_15540,N_13292);
nand U16904 (N_16904,N_12526,N_13726);
and U16905 (N_16905,N_12698,N_13736);
nor U16906 (N_16906,N_13216,N_13505);
and U16907 (N_16907,N_13101,N_15009);
nand U16908 (N_16908,N_15020,N_14718);
nor U16909 (N_16909,N_14056,N_14097);
or U16910 (N_16910,N_13331,N_15514);
and U16911 (N_16911,N_13988,N_13629);
or U16912 (N_16912,N_13419,N_13023);
xnor U16913 (N_16913,N_14830,N_13902);
nand U16914 (N_16914,N_12576,N_13712);
or U16915 (N_16915,N_15153,N_12510);
and U16916 (N_16916,N_12833,N_14900);
nand U16917 (N_16917,N_15118,N_15482);
xnor U16918 (N_16918,N_13614,N_12596);
nand U16919 (N_16919,N_12915,N_15250);
nor U16920 (N_16920,N_13444,N_12551);
nor U16921 (N_16921,N_12935,N_15112);
nand U16922 (N_16922,N_14925,N_14624);
and U16923 (N_16923,N_15192,N_15298);
xor U16924 (N_16924,N_13118,N_15282);
or U16925 (N_16925,N_14367,N_13237);
xor U16926 (N_16926,N_14009,N_13667);
nor U16927 (N_16927,N_13313,N_13632);
and U16928 (N_16928,N_12513,N_14926);
and U16929 (N_16929,N_15604,N_15002);
nand U16930 (N_16930,N_13989,N_12997);
and U16931 (N_16931,N_15413,N_13780);
xnor U16932 (N_16932,N_12856,N_13271);
xor U16933 (N_16933,N_15405,N_14822);
nand U16934 (N_16934,N_14801,N_13307);
nor U16935 (N_16935,N_14102,N_15424);
nor U16936 (N_16936,N_15470,N_12891);
nor U16937 (N_16937,N_13043,N_14261);
nor U16938 (N_16938,N_14156,N_13500);
and U16939 (N_16939,N_15227,N_15336);
and U16940 (N_16940,N_13320,N_13290);
and U16941 (N_16941,N_13449,N_13649);
xnor U16942 (N_16942,N_14587,N_14984);
nand U16943 (N_16943,N_14293,N_13786);
or U16944 (N_16944,N_14866,N_14843);
nand U16945 (N_16945,N_15240,N_15451);
nand U16946 (N_16946,N_13504,N_12562);
nand U16947 (N_16947,N_12805,N_14222);
and U16948 (N_16948,N_13520,N_15458);
nor U16949 (N_16949,N_14539,N_14872);
xnor U16950 (N_16950,N_13210,N_13029);
nor U16951 (N_16951,N_13498,N_13049);
or U16952 (N_16952,N_15174,N_13615);
or U16953 (N_16953,N_12703,N_13693);
xnor U16954 (N_16954,N_12683,N_12871);
xnor U16955 (N_16955,N_13430,N_14391);
or U16956 (N_16956,N_13349,N_13138);
nor U16957 (N_16957,N_14435,N_14210);
nor U16958 (N_16958,N_13707,N_15211);
and U16959 (N_16959,N_14043,N_13147);
nor U16960 (N_16960,N_13470,N_14895);
or U16961 (N_16961,N_14161,N_14358);
nand U16962 (N_16962,N_14327,N_12919);
and U16963 (N_16963,N_14650,N_14483);
xnor U16964 (N_16964,N_14861,N_14750);
or U16965 (N_16965,N_13403,N_15596);
xor U16966 (N_16966,N_14542,N_14260);
and U16967 (N_16967,N_14973,N_15123);
nor U16968 (N_16968,N_14858,N_14541);
nand U16969 (N_16969,N_14062,N_12843);
nand U16970 (N_16970,N_15011,N_13804);
and U16971 (N_16971,N_12740,N_13291);
xor U16972 (N_16972,N_12720,N_14466);
and U16973 (N_16973,N_15320,N_13578);
nand U16974 (N_16974,N_13911,N_12898);
nor U16975 (N_16975,N_13182,N_14664);
nor U16976 (N_16976,N_15344,N_14155);
and U16977 (N_16977,N_12675,N_12668);
xnor U16978 (N_16978,N_15268,N_13071);
and U16979 (N_16979,N_13974,N_13298);
xnor U16980 (N_16980,N_13829,N_12694);
nor U16981 (N_16981,N_13861,N_15171);
nand U16982 (N_16982,N_13742,N_14991);
or U16983 (N_16983,N_13950,N_15253);
xor U16984 (N_16984,N_13621,N_13392);
xor U16985 (N_16985,N_13408,N_13672);
xor U16986 (N_16986,N_13230,N_13572);
xor U16987 (N_16987,N_13747,N_14226);
nor U16988 (N_16988,N_14914,N_13868);
nor U16989 (N_16989,N_14141,N_14877);
nor U16990 (N_16990,N_14966,N_13217);
xnor U16991 (N_16991,N_13361,N_14438);
nor U16992 (N_16992,N_13224,N_12782);
xnor U16993 (N_16993,N_14901,N_13937);
or U16994 (N_16994,N_14089,N_14557);
or U16995 (N_16995,N_14268,N_14689);
nand U16996 (N_16996,N_14573,N_15279);
xnor U16997 (N_16997,N_13959,N_15156);
xor U16998 (N_16998,N_14618,N_15517);
nand U16999 (N_16999,N_14804,N_14151);
nor U17000 (N_17000,N_15089,N_15403);
and U17001 (N_17001,N_14234,N_14181);
and U17002 (N_17002,N_15351,N_13231);
or U17003 (N_17003,N_14471,N_13593);
xnor U17004 (N_17004,N_14698,N_13980);
nand U17005 (N_17005,N_12793,N_13785);
xnor U17006 (N_17006,N_15309,N_12861);
xor U17007 (N_17007,N_13062,N_14603);
nor U17008 (N_17008,N_14487,N_15523);
nand U17009 (N_17009,N_14134,N_13694);
and U17010 (N_17010,N_14578,N_15040);
and U17011 (N_17011,N_14236,N_12560);
nor U17012 (N_17012,N_15184,N_14213);
xor U17013 (N_17013,N_12810,N_14516);
or U17014 (N_17014,N_13139,N_14421);
nand U17015 (N_17015,N_14627,N_14484);
xor U17016 (N_17016,N_12963,N_12536);
nor U17017 (N_17017,N_13423,N_13468);
or U17018 (N_17018,N_13006,N_15598);
and U17019 (N_17019,N_14276,N_14563);
xor U17020 (N_17020,N_15563,N_14986);
nor U17021 (N_17021,N_13460,N_14885);
nor U17022 (N_17022,N_15385,N_13547);
nor U17023 (N_17023,N_15359,N_14250);
nor U17024 (N_17024,N_14909,N_15012);
nor U17025 (N_17025,N_13808,N_14074);
and U17026 (N_17026,N_13347,N_13709);
or U17027 (N_17027,N_15370,N_13360);
nor U17028 (N_17028,N_12504,N_14371);
xnor U17029 (N_17029,N_13359,N_13293);
and U17030 (N_17030,N_14142,N_13931);
nand U17031 (N_17031,N_12753,N_14709);
and U17032 (N_17032,N_13761,N_13550);
nor U17033 (N_17033,N_14828,N_13245);
or U17034 (N_17034,N_12624,N_15269);
or U17035 (N_17035,N_12528,N_13004);
and U17036 (N_17036,N_12981,N_13951);
and U17037 (N_17037,N_13745,N_14217);
or U17038 (N_17038,N_15244,N_13010);
and U17039 (N_17039,N_15167,N_13035);
and U17040 (N_17040,N_14397,N_13250);
or U17041 (N_17041,N_12962,N_15155);
xor U17042 (N_17042,N_13876,N_12593);
nor U17043 (N_17043,N_13639,N_13318);
nand U17044 (N_17044,N_15355,N_15254);
xor U17045 (N_17045,N_13945,N_14035);
xnor U17046 (N_17046,N_13822,N_15330);
nor U17047 (N_17047,N_14715,N_12598);
and U17048 (N_17048,N_14792,N_14406);
nor U17049 (N_17049,N_12910,N_14985);
and U17050 (N_17050,N_13775,N_13045);
nand U17051 (N_17051,N_14724,N_14473);
and U17052 (N_17052,N_13018,N_13620);
xnor U17053 (N_17053,N_13606,N_13854);
nand U17054 (N_17054,N_14875,N_12974);
xnor U17055 (N_17055,N_15420,N_14890);
nand U17056 (N_17056,N_13352,N_15281);
nor U17057 (N_17057,N_15076,N_12520);
and U17058 (N_17058,N_14640,N_14553);
or U17059 (N_17059,N_13031,N_14047);
or U17060 (N_17060,N_15354,N_12899);
xor U17061 (N_17061,N_13335,N_14269);
or U17062 (N_17062,N_14742,N_13507);
xnor U17063 (N_17063,N_13779,N_12688);
nand U17064 (N_17064,N_13807,N_15380);
nand U17065 (N_17065,N_12534,N_13295);
xnor U17066 (N_17066,N_13154,N_15140);
nand U17067 (N_17067,N_15075,N_13930);
and U17068 (N_17068,N_12677,N_14396);
or U17069 (N_17069,N_13484,N_13562);
nor U17070 (N_17070,N_12594,N_14030);
nand U17071 (N_17071,N_13941,N_13920);
nand U17072 (N_17072,N_15466,N_12767);
nand U17073 (N_17073,N_15392,N_15613);
and U17074 (N_17074,N_14786,N_12546);
xnor U17075 (N_17075,N_14377,N_13519);
nor U17076 (N_17076,N_14224,N_13459);
nand U17077 (N_17077,N_13724,N_14660);
or U17078 (N_17078,N_12763,N_12557);
or U17079 (N_17079,N_14216,N_14748);
and U17080 (N_17080,N_13037,N_12855);
xor U17081 (N_17081,N_15473,N_13165);
or U17082 (N_17082,N_15305,N_15467);
nor U17083 (N_17083,N_14902,N_15341);
nand U17084 (N_17084,N_14591,N_15560);
and U17085 (N_17085,N_14980,N_14880);
nor U17086 (N_17086,N_13072,N_15367);
and U17087 (N_17087,N_13781,N_14568);
xor U17088 (N_17088,N_14946,N_15346);
or U17089 (N_17089,N_13767,N_14046);
and U17090 (N_17090,N_14803,N_12766);
and U17091 (N_17091,N_12556,N_12661);
xor U17092 (N_17092,N_12636,N_13135);
nor U17093 (N_17093,N_14523,N_12841);
nand U17094 (N_17094,N_15113,N_14246);
and U17095 (N_17095,N_15345,N_13871);
xnor U17096 (N_17096,N_13573,N_15335);
and U17097 (N_17097,N_15595,N_15487);
and U17098 (N_17098,N_14879,N_14215);
nand U17099 (N_17099,N_13478,N_14464);
or U17100 (N_17100,N_12588,N_13341);
nand U17101 (N_17101,N_12558,N_15278);
nand U17102 (N_17102,N_15255,N_13555);
and U17103 (N_17103,N_13074,N_12565);
or U17104 (N_17104,N_13234,N_14502);
nor U17105 (N_17105,N_13003,N_14654);
or U17106 (N_17106,N_13211,N_12966);
and U17107 (N_17107,N_12611,N_14763);
nand U17108 (N_17108,N_15412,N_13203);
nand U17109 (N_17109,N_14730,N_12550);
xor U17110 (N_17110,N_12608,N_15402);
xor U17111 (N_17111,N_14994,N_14456);
and U17112 (N_17112,N_13510,N_15365);
xnor U17113 (N_17113,N_13017,N_14003);
and U17114 (N_17114,N_13609,N_14598);
nor U17115 (N_17115,N_13525,N_14387);
and U17116 (N_17116,N_15202,N_13528);
nand U17117 (N_17117,N_13954,N_13121);
nor U17118 (N_17118,N_14109,N_12944);
and U17119 (N_17119,N_15417,N_14770);
nor U17120 (N_17120,N_13244,N_13790);
and U17121 (N_17121,N_14680,N_14571);
or U17122 (N_17122,N_14157,N_15535);
and U17123 (N_17123,N_14972,N_12905);
and U17124 (N_17124,N_13409,N_12872);
nor U17125 (N_17125,N_12532,N_13582);
and U17126 (N_17126,N_15074,N_14001);
xnor U17127 (N_17127,N_13086,N_13933);
or U17128 (N_17128,N_13145,N_12571);
nor U17129 (N_17129,N_14439,N_13818);
or U17130 (N_17130,N_12664,N_13864);
or U17131 (N_17131,N_15312,N_14237);
nand U17132 (N_17132,N_12961,N_13105);
xor U17133 (N_17133,N_14708,N_15159);
xnor U17134 (N_17134,N_13142,N_13473);
xor U17135 (N_17135,N_15236,N_12647);
xor U17136 (N_17136,N_14854,N_13585);
or U17137 (N_17137,N_12807,N_12986);
nand U17138 (N_17138,N_12530,N_13866);
nand U17139 (N_17139,N_13046,N_13163);
nor U17140 (N_17140,N_14187,N_14766);
xnor U17141 (N_17141,N_15570,N_13634);
nand U17142 (N_17142,N_15621,N_13729);
or U17143 (N_17143,N_14797,N_14711);
xnor U17144 (N_17144,N_15117,N_14767);
or U17145 (N_17145,N_15446,N_14085);
nor U17146 (N_17146,N_15152,N_13732);
and U17147 (N_17147,N_13492,N_14275);
and U17148 (N_17148,N_13221,N_13324);
nand U17149 (N_17149,N_13122,N_13251);
and U17150 (N_17150,N_14018,N_13835);
and U17151 (N_17151,N_13878,N_13816);
nor U17152 (N_17152,N_15136,N_14905);
nand U17153 (N_17153,N_14451,N_12844);
and U17154 (N_17154,N_12779,N_12512);
nor U17155 (N_17155,N_15431,N_12804);
nand U17156 (N_17156,N_15290,N_13771);
nand U17157 (N_17157,N_13884,N_12848);
xnor U17158 (N_17158,N_14411,N_15280);
xnor U17159 (N_17159,N_13561,N_15111);
xor U17160 (N_17160,N_14491,N_13698);
or U17161 (N_17161,N_15200,N_14426);
nand U17162 (N_17162,N_14310,N_14638);
nand U17163 (N_17163,N_13109,N_15177);
xnor U17164 (N_17164,N_12958,N_13090);
or U17165 (N_17165,N_12730,N_13960);
nor U17166 (N_17166,N_13329,N_15073);
and U17167 (N_17167,N_14336,N_14506);
and U17168 (N_17168,N_13656,N_12927);
nor U17169 (N_17169,N_12747,N_14982);
nor U17170 (N_17170,N_13702,N_14374);
and U17171 (N_17171,N_12934,N_15597);
and U17172 (N_17172,N_14462,N_15059);
xnor U17173 (N_17173,N_13137,N_13189);
xnor U17174 (N_17174,N_14183,N_15275);
and U17175 (N_17175,N_14674,N_13794);
or U17176 (N_17176,N_14580,N_14136);
and U17177 (N_17177,N_12903,N_12559);
xor U17178 (N_17178,N_14851,N_12977);
and U17179 (N_17179,N_13806,N_13720);
nand U17180 (N_17180,N_14950,N_12990);
and U17181 (N_17181,N_14672,N_14093);
and U17182 (N_17182,N_15218,N_12579);
nand U17183 (N_17183,N_14388,N_15274);
nor U17184 (N_17184,N_13377,N_12615);
and U17185 (N_17185,N_12901,N_15592);
xnor U17186 (N_17186,N_13710,N_13126);
and U17187 (N_17187,N_13936,N_12566);
nand U17188 (N_17188,N_15161,N_15345);
nor U17189 (N_17189,N_13163,N_14582);
and U17190 (N_17190,N_14820,N_12557);
and U17191 (N_17191,N_14749,N_14231);
and U17192 (N_17192,N_14580,N_15472);
and U17193 (N_17193,N_13243,N_15441);
and U17194 (N_17194,N_15208,N_12732);
nand U17195 (N_17195,N_14362,N_14115);
and U17196 (N_17196,N_13775,N_14103);
and U17197 (N_17197,N_13191,N_13355);
and U17198 (N_17198,N_12830,N_12926);
nor U17199 (N_17199,N_12756,N_15300);
and U17200 (N_17200,N_14435,N_14380);
and U17201 (N_17201,N_13507,N_13056);
xnor U17202 (N_17202,N_15056,N_15569);
nor U17203 (N_17203,N_13601,N_13096);
nor U17204 (N_17204,N_14779,N_13516);
xnor U17205 (N_17205,N_12990,N_13180);
nand U17206 (N_17206,N_15351,N_13286);
xor U17207 (N_17207,N_15596,N_15001);
nand U17208 (N_17208,N_15330,N_14749);
nor U17209 (N_17209,N_15291,N_14007);
or U17210 (N_17210,N_15585,N_14903);
xnor U17211 (N_17211,N_14109,N_15081);
xnor U17212 (N_17212,N_14938,N_14329);
or U17213 (N_17213,N_12504,N_14065);
or U17214 (N_17214,N_14852,N_12683);
xnor U17215 (N_17215,N_13601,N_13824);
nor U17216 (N_17216,N_14915,N_14169);
nor U17217 (N_17217,N_15264,N_13521);
nand U17218 (N_17218,N_14363,N_13047);
nor U17219 (N_17219,N_14417,N_15113);
nand U17220 (N_17220,N_13199,N_13428);
or U17221 (N_17221,N_13827,N_13957);
and U17222 (N_17222,N_14930,N_15067);
and U17223 (N_17223,N_15088,N_13844);
or U17224 (N_17224,N_13999,N_13411);
and U17225 (N_17225,N_15233,N_12804);
nand U17226 (N_17226,N_14017,N_15393);
nor U17227 (N_17227,N_13285,N_14935);
and U17228 (N_17228,N_14965,N_12868);
nand U17229 (N_17229,N_13808,N_13326);
nor U17230 (N_17230,N_14093,N_12516);
and U17231 (N_17231,N_13038,N_14860);
nor U17232 (N_17232,N_14705,N_14986);
and U17233 (N_17233,N_15475,N_13139);
or U17234 (N_17234,N_13938,N_15048);
nand U17235 (N_17235,N_13327,N_12574);
nand U17236 (N_17236,N_13681,N_14091);
and U17237 (N_17237,N_13906,N_15122);
and U17238 (N_17238,N_14032,N_12956);
xnor U17239 (N_17239,N_12697,N_14930);
nand U17240 (N_17240,N_13848,N_12566);
or U17241 (N_17241,N_14374,N_15408);
xnor U17242 (N_17242,N_15607,N_13221);
and U17243 (N_17243,N_14600,N_13767);
and U17244 (N_17244,N_15201,N_13479);
and U17245 (N_17245,N_12799,N_13736);
nor U17246 (N_17246,N_14184,N_14418);
or U17247 (N_17247,N_13243,N_14524);
or U17248 (N_17248,N_15331,N_13790);
xor U17249 (N_17249,N_14121,N_15178);
xnor U17250 (N_17250,N_12569,N_14092);
nor U17251 (N_17251,N_13573,N_15569);
or U17252 (N_17252,N_12711,N_13803);
xnor U17253 (N_17253,N_15580,N_14771);
nand U17254 (N_17254,N_14583,N_15206);
nand U17255 (N_17255,N_14814,N_15198);
xnor U17256 (N_17256,N_14128,N_12840);
and U17257 (N_17257,N_15171,N_12588);
nor U17258 (N_17258,N_12748,N_14247);
xor U17259 (N_17259,N_15121,N_14852);
and U17260 (N_17260,N_13208,N_13897);
nand U17261 (N_17261,N_14761,N_14299);
xor U17262 (N_17262,N_14903,N_14974);
or U17263 (N_17263,N_14853,N_12668);
and U17264 (N_17264,N_14082,N_12861);
xor U17265 (N_17265,N_13965,N_13008);
or U17266 (N_17266,N_15624,N_13388);
nor U17267 (N_17267,N_13859,N_14344);
nand U17268 (N_17268,N_14021,N_12701);
or U17269 (N_17269,N_13750,N_14967);
nor U17270 (N_17270,N_14413,N_13494);
or U17271 (N_17271,N_14721,N_14762);
nand U17272 (N_17272,N_12770,N_14586);
and U17273 (N_17273,N_13221,N_14865);
or U17274 (N_17274,N_14499,N_15282);
nand U17275 (N_17275,N_14071,N_13102);
nand U17276 (N_17276,N_14275,N_14879);
or U17277 (N_17277,N_14932,N_14576);
and U17278 (N_17278,N_12887,N_15182);
xnor U17279 (N_17279,N_13645,N_13343);
and U17280 (N_17280,N_14978,N_13087);
or U17281 (N_17281,N_14701,N_14193);
xnor U17282 (N_17282,N_12679,N_15186);
xnor U17283 (N_17283,N_13125,N_15293);
and U17284 (N_17284,N_13782,N_14313);
xor U17285 (N_17285,N_15215,N_14738);
nand U17286 (N_17286,N_14008,N_14761);
nor U17287 (N_17287,N_12929,N_15110);
or U17288 (N_17288,N_15059,N_15371);
nand U17289 (N_17289,N_14197,N_12545);
nand U17290 (N_17290,N_13551,N_14364);
xnor U17291 (N_17291,N_14519,N_15411);
or U17292 (N_17292,N_13462,N_12864);
nor U17293 (N_17293,N_12569,N_15604);
and U17294 (N_17294,N_15508,N_15380);
and U17295 (N_17295,N_12801,N_14440);
or U17296 (N_17296,N_12519,N_15601);
nor U17297 (N_17297,N_12826,N_14025);
nand U17298 (N_17298,N_14031,N_14424);
nand U17299 (N_17299,N_14534,N_12981);
or U17300 (N_17300,N_12685,N_14766);
nand U17301 (N_17301,N_14433,N_14882);
and U17302 (N_17302,N_15109,N_14417);
nand U17303 (N_17303,N_14911,N_13840);
nor U17304 (N_17304,N_13833,N_14210);
nand U17305 (N_17305,N_12765,N_14907);
nand U17306 (N_17306,N_14452,N_15570);
or U17307 (N_17307,N_14725,N_15481);
or U17308 (N_17308,N_15013,N_13609);
or U17309 (N_17309,N_12673,N_12907);
or U17310 (N_17310,N_13630,N_14333);
and U17311 (N_17311,N_12882,N_13696);
nor U17312 (N_17312,N_15597,N_15138);
or U17313 (N_17313,N_15266,N_15200);
and U17314 (N_17314,N_13566,N_13082);
xor U17315 (N_17315,N_15388,N_14862);
and U17316 (N_17316,N_13149,N_14119);
nor U17317 (N_17317,N_12949,N_13078);
nor U17318 (N_17318,N_13550,N_14516);
xor U17319 (N_17319,N_14796,N_12737);
and U17320 (N_17320,N_14751,N_13166);
nand U17321 (N_17321,N_15214,N_15618);
nor U17322 (N_17322,N_15514,N_14281);
nor U17323 (N_17323,N_13955,N_12611);
or U17324 (N_17324,N_14081,N_13797);
and U17325 (N_17325,N_13001,N_14502);
and U17326 (N_17326,N_14365,N_15089);
or U17327 (N_17327,N_14745,N_13906);
nor U17328 (N_17328,N_15118,N_15319);
or U17329 (N_17329,N_15512,N_12885);
nor U17330 (N_17330,N_13322,N_15471);
nor U17331 (N_17331,N_14668,N_15271);
nand U17332 (N_17332,N_14151,N_14997);
nor U17333 (N_17333,N_14974,N_14549);
or U17334 (N_17334,N_14323,N_12639);
and U17335 (N_17335,N_14750,N_15079);
nand U17336 (N_17336,N_14817,N_13885);
or U17337 (N_17337,N_14381,N_13714);
and U17338 (N_17338,N_14545,N_13191);
or U17339 (N_17339,N_13985,N_14735);
and U17340 (N_17340,N_13938,N_13353);
xor U17341 (N_17341,N_14948,N_14676);
or U17342 (N_17342,N_14392,N_15397);
and U17343 (N_17343,N_12600,N_12777);
and U17344 (N_17344,N_15040,N_13878);
xor U17345 (N_17345,N_14591,N_12692);
and U17346 (N_17346,N_15226,N_13692);
nand U17347 (N_17347,N_13122,N_12669);
xnor U17348 (N_17348,N_15126,N_12556);
xor U17349 (N_17349,N_13723,N_13063);
or U17350 (N_17350,N_14817,N_15012);
xor U17351 (N_17351,N_14675,N_12985);
and U17352 (N_17352,N_13340,N_15468);
xnor U17353 (N_17353,N_13293,N_15459);
xnor U17354 (N_17354,N_14097,N_13155);
nor U17355 (N_17355,N_15504,N_15094);
nor U17356 (N_17356,N_13079,N_13912);
and U17357 (N_17357,N_12939,N_14559);
nand U17358 (N_17358,N_15550,N_13784);
xnor U17359 (N_17359,N_15544,N_15265);
xnor U17360 (N_17360,N_13866,N_13279);
or U17361 (N_17361,N_12622,N_12698);
or U17362 (N_17362,N_14951,N_13091);
nand U17363 (N_17363,N_14705,N_15448);
or U17364 (N_17364,N_13949,N_13910);
and U17365 (N_17365,N_14495,N_13738);
or U17366 (N_17366,N_13520,N_15299);
and U17367 (N_17367,N_14415,N_13061);
or U17368 (N_17368,N_12646,N_12551);
xor U17369 (N_17369,N_15621,N_13126);
or U17370 (N_17370,N_12941,N_15307);
xnor U17371 (N_17371,N_13764,N_14220);
and U17372 (N_17372,N_15577,N_14158);
xor U17373 (N_17373,N_14075,N_13465);
xor U17374 (N_17374,N_14207,N_14455);
or U17375 (N_17375,N_14646,N_14327);
nor U17376 (N_17376,N_12532,N_13881);
xor U17377 (N_17377,N_13268,N_12865);
nor U17378 (N_17378,N_14670,N_15226);
nor U17379 (N_17379,N_14178,N_15085);
and U17380 (N_17380,N_12813,N_15604);
and U17381 (N_17381,N_15083,N_13244);
nand U17382 (N_17382,N_15278,N_15106);
xnor U17383 (N_17383,N_12996,N_14526);
and U17384 (N_17384,N_13306,N_15094);
or U17385 (N_17385,N_14809,N_14832);
or U17386 (N_17386,N_13005,N_14194);
or U17387 (N_17387,N_13139,N_12720);
and U17388 (N_17388,N_15171,N_15268);
and U17389 (N_17389,N_15514,N_12501);
or U17390 (N_17390,N_13224,N_12715);
and U17391 (N_17391,N_12734,N_15301);
nor U17392 (N_17392,N_15292,N_14477);
and U17393 (N_17393,N_15055,N_13840);
nor U17394 (N_17394,N_12740,N_14000);
nor U17395 (N_17395,N_14526,N_14295);
and U17396 (N_17396,N_13715,N_13755);
or U17397 (N_17397,N_13246,N_15440);
or U17398 (N_17398,N_14088,N_15447);
and U17399 (N_17399,N_14490,N_14726);
or U17400 (N_17400,N_14925,N_13845);
nand U17401 (N_17401,N_12660,N_15096);
or U17402 (N_17402,N_12599,N_14748);
and U17403 (N_17403,N_13334,N_13775);
nor U17404 (N_17404,N_14820,N_15408);
nor U17405 (N_17405,N_14876,N_15451);
or U17406 (N_17406,N_14958,N_13106);
and U17407 (N_17407,N_13682,N_14435);
or U17408 (N_17408,N_12940,N_14945);
nand U17409 (N_17409,N_13408,N_15314);
nand U17410 (N_17410,N_15328,N_13625);
nor U17411 (N_17411,N_13734,N_15566);
and U17412 (N_17412,N_15323,N_14838);
and U17413 (N_17413,N_14984,N_13878);
nor U17414 (N_17414,N_15065,N_13349);
xor U17415 (N_17415,N_12511,N_13339);
nor U17416 (N_17416,N_14215,N_13746);
xor U17417 (N_17417,N_13970,N_14518);
xor U17418 (N_17418,N_15160,N_14699);
nor U17419 (N_17419,N_13032,N_14427);
nand U17420 (N_17420,N_15320,N_15193);
and U17421 (N_17421,N_13451,N_12964);
xor U17422 (N_17422,N_14454,N_13021);
or U17423 (N_17423,N_14431,N_15523);
and U17424 (N_17424,N_12718,N_13218);
nor U17425 (N_17425,N_13299,N_12744);
or U17426 (N_17426,N_13829,N_13129);
nor U17427 (N_17427,N_12595,N_14557);
and U17428 (N_17428,N_14656,N_15357);
xnor U17429 (N_17429,N_15571,N_12865);
nand U17430 (N_17430,N_14192,N_14791);
nand U17431 (N_17431,N_14286,N_13537);
nor U17432 (N_17432,N_13458,N_15021);
and U17433 (N_17433,N_14543,N_14882);
and U17434 (N_17434,N_12555,N_12659);
xor U17435 (N_17435,N_15322,N_15566);
nand U17436 (N_17436,N_14812,N_13004);
and U17437 (N_17437,N_12829,N_13181);
xnor U17438 (N_17438,N_14970,N_13161);
nor U17439 (N_17439,N_14376,N_13647);
xnor U17440 (N_17440,N_15113,N_14606);
or U17441 (N_17441,N_14311,N_13029);
or U17442 (N_17442,N_12557,N_13748);
nor U17443 (N_17443,N_14534,N_13072);
nand U17444 (N_17444,N_12554,N_15534);
nor U17445 (N_17445,N_14852,N_14230);
xnor U17446 (N_17446,N_14122,N_15421);
and U17447 (N_17447,N_12505,N_13083);
xnor U17448 (N_17448,N_12520,N_13781);
nand U17449 (N_17449,N_12683,N_14716);
or U17450 (N_17450,N_13483,N_14476);
and U17451 (N_17451,N_14782,N_13528);
nor U17452 (N_17452,N_15268,N_13103);
or U17453 (N_17453,N_14905,N_13011);
nor U17454 (N_17454,N_14845,N_13720);
nor U17455 (N_17455,N_15005,N_14262);
nor U17456 (N_17456,N_15190,N_13768);
xor U17457 (N_17457,N_14157,N_14382);
or U17458 (N_17458,N_14732,N_14435);
nor U17459 (N_17459,N_12719,N_13221);
nor U17460 (N_17460,N_14914,N_13132);
and U17461 (N_17461,N_15427,N_14445);
nand U17462 (N_17462,N_15381,N_13125);
and U17463 (N_17463,N_14090,N_14077);
and U17464 (N_17464,N_12667,N_14361);
and U17465 (N_17465,N_13966,N_12679);
nor U17466 (N_17466,N_12868,N_12974);
nor U17467 (N_17467,N_14261,N_14127);
or U17468 (N_17468,N_14938,N_13302);
and U17469 (N_17469,N_14832,N_14257);
nand U17470 (N_17470,N_14135,N_14625);
and U17471 (N_17471,N_14299,N_14643);
and U17472 (N_17472,N_13195,N_13214);
nand U17473 (N_17473,N_15440,N_15159);
and U17474 (N_17474,N_12803,N_13343);
or U17475 (N_17475,N_12826,N_12590);
and U17476 (N_17476,N_13628,N_12612);
or U17477 (N_17477,N_13941,N_15488);
nand U17478 (N_17478,N_13742,N_13724);
and U17479 (N_17479,N_14938,N_13253);
or U17480 (N_17480,N_14595,N_15609);
nand U17481 (N_17481,N_14325,N_15405);
nor U17482 (N_17482,N_15145,N_15460);
or U17483 (N_17483,N_14432,N_15603);
xnor U17484 (N_17484,N_13168,N_13471);
nand U17485 (N_17485,N_12670,N_15315);
or U17486 (N_17486,N_14505,N_15083);
nand U17487 (N_17487,N_14826,N_14349);
or U17488 (N_17488,N_14389,N_12981);
or U17489 (N_17489,N_14672,N_13952);
and U17490 (N_17490,N_13117,N_14798);
nor U17491 (N_17491,N_14197,N_14644);
and U17492 (N_17492,N_13165,N_15205);
and U17493 (N_17493,N_15408,N_14581);
or U17494 (N_17494,N_14485,N_12953);
and U17495 (N_17495,N_13085,N_14107);
or U17496 (N_17496,N_12860,N_14808);
nand U17497 (N_17497,N_15020,N_13755);
xnor U17498 (N_17498,N_15331,N_12609);
xor U17499 (N_17499,N_15594,N_14937);
and U17500 (N_17500,N_14264,N_13798);
xor U17501 (N_17501,N_14192,N_12928);
nand U17502 (N_17502,N_14531,N_15009);
or U17503 (N_17503,N_12596,N_13616);
and U17504 (N_17504,N_14265,N_13036);
or U17505 (N_17505,N_15336,N_13273);
nor U17506 (N_17506,N_13453,N_14148);
or U17507 (N_17507,N_12565,N_15209);
and U17508 (N_17508,N_13522,N_13385);
xor U17509 (N_17509,N_13165,N_13270);
nor U17510 (N_17510,N_13165,N_15385);
nand U17511 (N_17511,N_14519,N_14020);
nor U17512 (N_17512,N_13264,N_14106);
or U17513 (N_17513,N_13155,N_15266);
or U17514 (N_17514,N_14418,N_15133);
and U17515 (N_17515,N_14760,N_14640);
xnor U17516 (N_17516,N_15507,N_14099);
xnor U17517 (N_17517,N_13917,N_14574);
nand U17518 (N_17518,N_12788,N_14660);
nor U17519 (N_17519,N_12506,N_15324);
xor U17520 (N_17520,N_13707,N_14698);
or U17521 (N_17521,N_12678,N_14485);
xnor U17522 (N_17522,N_13181,N_15236);
and U17523 (N_17523,N_15534,N_14796);
and U17524 (N_17524,N_14145,N_14687);
and U17525 (N_17525,N_13162,N_14253);
or U17526 (N_17526,N_15128,N_15169);
and U17527 (N_17527,N_14043,N_12598);
and U17528 (N_17528,N_14846,N_12851);
or U17529 (N_17529,N_15394,N_13109);
or U17530 (N_17530,N_15251,N_14467);
and U17531 (N_17531,N_14324,N_13763);
nand U17532 (N_17532,N_14887,N_12774);
xor U17533 (N_17533,N_13695,N_12916);
nor U17534 (N_17534,N_15562,N_14680);
or U17535 (N_17535,N_13072,N_13275);
nor U17536 (N_17536,N_12596,N_14953);
nand U17537 (N_17537,N_13210,N_13040);
xor U17538 (N_17538,N_13733,N_13008);
nand U17539 (N_17539,N_13329,N_15349);
or U17540 (N_17540,N_13791,N_13514);
and U17541 (N_17541,N_14064,N_14641);
and U17542 (N_17542,N_13417,N_15247);
nor U17543 (N_17543,N_13367,N_15491);
xor U17544 (N_17544,N_13198,N_14870);
nand U17545 (N_17545,N_15342,N_12522);
nand U17546 (N_17546,N_14881,N_14619);
nor U17547 (N_17547,N_13269,N_14084);
nand U17548 (N_17548,N_13488,N_14169);
nor U17549 (N_17549,N_15484,N_14847);
and U17550 (N_17550,N_13712,N_14897);
nor U17551 (N_17551,N_15484,N_13006);
xnor U17552 (N_17552,N_14575,N_14484);
xor U17553 (N_17553,N_15548,N_15269);
and U17554 (N_17554,N_13575,N_14610);
xnor U17555 (N_17555,N_13768,N_13728);
nand U17556 (N_17556,N_14876,N_13492);
nand U17557 (N_17557,N_13321,N_14289);
xnor U17558 (N_17558,N_15151,N_14826);
nand U17559 (N_17559,N_13645,N_13139);
xnor U17560 (N_17560,N_15393,N_14713);
nand U17561 (N_17561,N_15352,N_13838);
nor U17562 (N_17562,N_12912,N_14370);
nor U17563 (N_17563,N_14258,N_15498);
xor U17564 (N_17564,N_14698,N_14831);
nand U17565 (N_17565,N_13474,N_13097);
or U17566 (N_17566,N_13077,N_14381);
or U17567 (N_17567,N_14730,N_15506);
and U17568 (N_17568,N_15618,N_15592);
or U17569 (N_17569,N_15504,N_13605);
nand U17570 (N_17570,N_14711,N_12613);
xor U17571 (N_17571,N_14143,N_13453);
or U17572 (N_17572,N_12780,N_15221);
nand U17573 (N_17573,N_13610,N_13043);
or U17574 (N_17574,N_12987,N_14775);
nand U17575 (N_17575,N_13623,N_13382);
and U17576 (N_17576,N_15209,N_13197);
nor U17577 (N_17577,N_13993,N_12853);
or U17578 (N_17578,N_12904,N_15093);
nand U17579 (N_17579,N_13849,N_15318);
nor U17580 (N_17580,N_12961,N_15402);
nor U17581 (N_17581,N_13887,N_12966);
or U17582 (N_17582,N_13206,N_15452);
nand U17583 (N_17583,N_14209,N_12541);
xnor U17584 (N_17584,N_14225,N_14456);
nor U17585 (N_17585,N_14817,N_13191);
and U17586 (N_17586,N_14008,N_15231);
nor U17587 (N_17587,N_13586,N_13518);
and U17588 (N_17588,N_14121,N_15119);
nand U17589 (N_17589,N_14787,N_14682);
xor U17590 (N_17590,N_13807,N_15094);
nor U17591 (N_17591,N_12604,N_15548);
xor U17592 (N_17592,N_13199,N_13423);
xnor U17593 (N_17593,N_14004,N_13941);
nor U17594 (N_17594,N_14581,N_15052);
and U17595 (N_17595,N_14380,N_15568);
or U17596 (N_17596,N_14597,N_14261);
xnor U17597 (N_17597,N_15286,N_13786);
or U17598 (N_17598,N_14431,N_13904);
nor U17599 (N_17599,N_14339,N_15278);
or U17600 (N_17600,N_14427,N_13363);
xor U17601 (N_17601,N_15624,N_13739);
nand U17602 (N_17602,N_13042,N_14202);
and U17603 (N_17603,N_14425,N_12541);
nand U17604 (N_17604,N_14097,N_14357);
xor U17605 (N_17605,N_13236,N_13320);
or U17606 (N_17606,N_14736,N_14860);
nor U17607 (N_17607,N_13136,N_15307);
xnor U17608 (N_17608,N_15509,N_14051);
and U17609 (N_17609,N_13755,N_14883);
nand U17610 (N_17610,N_14933,N_14583);
nand U17611 (N_17611,N_12764,N_13830);
or U17612 (N_17612,N_15611,N_14740);
and U17613 (N_17613,N_13933,N_14000);
or U17614 (N_17614,N_14419,N_12974);
and U17615 (N_17615,N_15118,N_13115);
or U17616 (N_17616,N_13617,N_14866);
nand U17617 (N_17617,N_14083,N_15537);
nor U17618 (N_17618,N_15484,N_15431);
xor U17619 (N_17619,N_13674,N_15418);
or U17620 (N_17620,N_12682,N_12962);
xnor U17621 (N_17621,N_14747,N_14187);
nor U17622 (N_17622,N_15192,N_13191);
nor U17623 (N_17623,N_14574,N_12906);
nor U17624 (N_17624,N_13796,N_13631);
nor U17625 (N_17625,N_14971,N_15190);
and U17626 (N_17626,N_15336,N_13178);
or U17627 (N_17627,N_14164,N_15375);
nand U17628 (N_17628,N_13513,N_14352);
nor U17629 (N_17629,N_13799,N_15512);
nor U17630 (N_17630,N_15165,N_15449);
nor U17631 (N_17631,N_13219,N_13471);
nor U17632 (N_17632,N_13880,N_13841);
nor U17633 (N_17633,N_13443,N_12554);
xnor U17634 (N_17634,N_13897,N_12939);
or U17635 (N_17635,N_12662,N_13033);
xor U17636 (N_17636,N_13284,N_13101);
and U17637 (N_17637,N_13318,N_13245);
xnor U17638 (N_17638,N_14137,N_14739);
xor U17639 (N_17639,N_12766,N_13209);
and U17640 (N_17640,N_13425,N_14550);
and U17641 (N_17641,N_15592,N_13597);
nor U17642 (N_17642,N_12805,N_12597);
nand U17643 (N_17643,N_13971,N_14190);
and U17644 (N_17644,N_15288,N_13706);
xor U17645 (N_17645,N_13260,N_13403);
xor U17646 (N_17646,N_12752,N_13156);
nand U17647 (N_17647,N_15227,N_14979);
or U17648 (N_17648,N_12756,N_12935);
nor U17649 (N_17649,N_13783,N_14333);
xnor U17650 (N_17650,N_13991,N_14665);
xor U17651 (N_17651,N_12668,N_12793);
nand U17652 (N_17652,N_14063,N_14375);
nand U17653 (N_17653,N_13272,N_15562);
and U17654 (N_17654,N_14902,N_12818);
nor U17655 (N_17655,N_13478,N_15386);
and U17656 (N_17656,N_13357,N_13414);
and U17657 (N_17657,N_12652,N_12968);
or U17658 (N_17658,N_15371,N_12727);
nand U17659 (N_17659,N_12590,N_13447);
or U17660 (N_17660,N_15208,N_12961);
xnor U17661 (N_17661,N_15197,N_12695);
nand U17662 (N_17662,N_14678,N_12915);
or U17663 (N_17663,N_14930,N_13650);
xor U17664 (N_17664,N_14277,N_13445);
or U17665 (N_17665,N_13806,N_13608);
nor U17666 (N_17666,N_14300,N_13037);
nand U17667 (N_17667,N_14809,N_14123);
xor U17668 (N_17668,N_15191,N_14709);
nor U17669 (N_17669,N_14830,N_15052);
xor U17670 (N_17670,N_13178,N_12923);
nor U17671 (N_17671,N_12957,N_15062);
xor U17672 (N_17672,N_12989,N_15543);
xor U17673 (N_17673,N_15249,N_14788);
nand U17674 (N_17674,N_15604,N_15579);
nor U17675 (N_17675,N_14193,N_13467);
or U17676 (N_17676,N_14567,N_13560);
and U17677 (N_17677,N_12945,N_13202);
nand U17678 (N_17678,N_13101,N_13562);
nand U17679 (N_17679,N_13865,N_15287);
or U17680 (N_17680,N_15045,N_14953);
nand U17681 (N_17681,N_14532,N_15560);
or U17682 (N_17682,N_15148,N_13061);
and U17683 (N_17683,N_13380,N_13850);
xnor U17684 (N_17684,N_13367,N_14543);
nand U17685 (N_17685,N_14011,N_14009);
nand U17686 (N_17686,N_14896,N_15470);
or U17687 (N_17687,N_15241,N_13427);
xnor U17688 (N_17688,N_15606,N_15264);
or U17689 (N_17689,N_13357,N_14143);
and U17690 (N_17690,N_14787,N_14911);
nor U17691 (N_17691,N_13734,N_14032);
or U17692 (N_17692,N_13997,N_14380);
and U17693 (N_17693,N_15108,N_12644);
and U17694 (N_17694,N_13152,N_13427);
and U17695 (N_17695,N_14230,N_15007);
or U17696 (N_17696,N_15123,N_14503);
and U17697 (N_17697,N_14724,N_15354);
and U17698 (N_17698,N_13830,N_13397);
and U17699 (N_17699,N_12627,N_13997);
or U17700 (N_17700,N_13813,N_13162);
and U17701 (N_17701,N_13271,N_13551);
xor U17702 (N_17702,N_14562,N_14164);
or U17703 (N_17703,N_14655,N_15022);
and U17704 (N_17704,N_12953,N_12601);
and U17705 (N_17705,N_14056,N_13984);
or U17706 (N_17706,N_12674,N_13180);
or U17707 (N_17707,N_14399,N_12530);
nand U17708 (N_17708,N_15460,N_13301);
nand U17709 (N_17709,N_14990,N_15208);
xnor U17710 (N_17710,N_14337,N_14341);
xnor U17711 (N_17711,N_13631,N_12694);
or U17712 (N_17712,N_13780,N_13407);
and U17713 (N_17713,N_13410,N_13117);
and U17714 (N_17714,N_12636,N_12606);
or U17715 (N_17715,N_14348,N_12545);
xnor U17716 (N_17716,N_15367,N_12657);
or U17717 (N_17717,N_14056,N_14006);
nand U17718 (N_17718,N_12956,N_13448);
xnor U17719 (N_17719,N_13226,N_15606);
or U17720 (N_17720,N_13575,N_14052);
and U17721 (N_17721,N_13625,N_12804);
xor U17722 (N_17722,N_15020,N_13851);
nor U17723 (N_17723,N_12961,N_12524);
and U17724 (N_17724,N_15524,N_12569);
nor U17725 (N_17725,N_13318,N_15394);
nor U17726 (N_17726,N_13087,N_14174);
nor U17727 (N_17727,N_14046,N_15119);
nand U17728 (N_17728,N_12690,N_13768);
nand U17729 (N_17729,N_12614,N_13932);
nor U17730 (N_17730,N_15179,N_13390);
and U17731 (N_17731,N_13633,N_13104);
nand U17732 (N_17732,N_14848,N_12633);
xor U17733 (N_17733,N_14602,N_14507);
or U17734 (N_17734,N_14221,N_15425);
or U17735 (N_17735,N_15052,N_15186);
xnor U17736 (N_17736,N_14176,N_12986);
or U17737 (N_17737,N_13709,N_14487);
xor U17738 (N_17738,N_14763,N_14266);
nand U17739 (N_17739,N_15537,N_13437);
nor U17740 (N_17740,N_14398,N_12667);
and U17741 (N_17741,N_14714,N_14150);
or U17742 (N_17742,N_14421,N_15475);
nand U17743 (N_17743,N_13533,N_13603);
xnor U17744 (N_17744,N_15376,N_14027);
or U17745 (N_17745,N_14187,N_13179);
and U17746 (N_17746,N_12625,N_14819);
nor U17747 (N_17747,N_13994,N_12973);
and U17748 (N_17748,N_12673,N_15226);
or U17749 (N_17749,N_13941,N_13756);
or U17750 (N_17750,N_14903,N_14970);
nor U17751 (N_17751,N_13453,N_15412);
xor U17752 (N_17752,N_13582,N_13408);
nor U17753 (N_17753,N_12814,N_12630);
nand U17754 (N_17754,N_14783,N_14921);
nor U17755 (N_17755,N_14819,N_14732);
and U17756 (N_17756,N_14022,N_14624);
and U17757 (N_17757,N_13586,N_12775);
nor U17758 (N_17758,N_14038,N_15041);
nor U17759 (N_17759,N_13250,N_14227);
and U17760 (N_17760,N_12939,N_13825);
and U17761 (N_17761,N_12748,N_12502);
nand U17762 (N_17762,N_15434,N_14512);
nand U17763 (N_17763,N_12938,N_14173);
nand U17764 (N_17764,N_14087,N_14640);
nand U17765 (N_17765,N_13799,N_14246);
nor U17766 (N_17766,N_14657,N_15007);
nand U17767 (N_17767,N_14928,N_14576);
or U17768 (N_17768,N_14107,N_13772);
and U17769 (N_17769,N_14879,N_14178);
nor U17770 (N_17770,N_15347,N_14208);
nand U17771 (N_17771,N_12566,N_14675);
or U17772 (N_17772,N_15414,N_14887);
or U17773 (N_17773,N_15534,N_15135);
and U17774 (N_17774,N_14147,N_12941);
xnor U17775 (N_17775,N_13043,N_14545);
nand U17776 (N_17776,N_15121,N_14275);
nor U17777 (N_17777,N_14808,N_13688);
xor U17778 (N_17778,N_14343,N_13355);
and U17779 (N_17779,N_13992,N_12655);
or U17780 (N_17780,N_12684,N_13437);
nand U17781 (N_17781,N_13562,N_12934);
or U17782 (N_17782,N_14543,N_12504);
and U17783 (N_17783,N_13876,N_14553);
and U17784 (N_17784,N_14462,N_14595);
nand U17785 (N_17785,N_13514,N_13590);
nor U17786 (N_17786,N_13502,N_15024);
xnor U17787 (N_17787,N_14776,N_14101);
and U17788 (N_17788,N_15472,N_13916);
nand U17789 (N_17789,N_15431,N_13668);
nand U17790 (N_17790,N_15593,N_14435);
nand U17791 (N_17791,N_12755,N_13380);
nor U17792 (N_17792,N_14460,N_13776);
xor U17793 (N_17793,N_12573,N_14688);
and U17794 (N_17794,N_13880,N_15549);
or U17795 (N_17795,N_13174,N_14201);
nand U17796 (N_17796,N_14531,N_13779);
and U17797 (N_17797,N_12517,N_12676);
or U17798 (N_17798,N_13942,N_13450);
nand U17799 (N_17799,N_15372,N_13728);
nor U17800 (N_17800,N_14662,N_13468);
and U17801 (N_17801,N_15243,N_12656);
or U17802 (N_17802,N_13662,N_14252);
nor U17803 (N_17803,N_15513,N_15059);
xor U17804 (N_17804,N_13342,N_14615);
nand U17805 (N_17805,N_14279,N_14322);
and U17806 (N_17806,N_13419,N_13689);
nor U17807 (N_17807,N_15586,N_13037);
nand U17808 (N_17808,N_13963,N_12892);
xor U17809 (N_17809,N_14197,N_14303);
nand U17810 (N_17810,N_14851,N_12776);
and U17811 (N_17811,N_13910,N_13642);
xnor U17812 (N_17812,N_15592,N_12993);
and U17813 (N_17813,N_14992,N_13822);
and U17814 (N_17814,N_13595,N_14837);
nor U17815 (N_17815,N_15522,N_13577);
nand U17816 (N_17816,N_13994,N_15341);
or U17817 (N_17817,N_15171,N_15050);
nor U17818 (N_17818,N_14385,N_13475);
or U17819 (N_17819,N_14885,N_15464);
nor U17820 (N_17820,N_12799,N_14082);
or U17821 (N_17821,N_13163,N_13100);
or U17822 (N_17822,N_13189,N_13272);
or U17823 (N_17823,N_13204,N_13007);
and U17824 (N_17824,N_12833,N_13820);
and U17825 (N_17825,N_12811,N_12682);
nand U17826 (N_17826,N_13495,N_14867);
or U17827 (N_17827,N_14509,N_13800);
and U17828 (N_17828,N_12959,N_15120);
xnor U17829 (N_17829,N_13879,N_12636);
or U17830 (N_17830,N_13207,N_15508);
xor U17831 (N_17831,N_14582,N_14987);
and U17832 (N_17832,N_13882,N_15137);
and U17833 (N_17833,N_15562,N_12943);
and U17834 (N_17834,N_14440,N_15598);
and U17835 (N_17835,N_13671,N_14423);
nand U17836 (N_17836,N_12942,N_15344);
nor U17837 (N_17837,N_12968,N_12732);
nor U17838 (N_17838,N_14040,N_14073);
xor U17839 (N_17839,N_12628,N_15214);
xnor U17840 (N_17840,N_14293,N_13986);
nor U17841 (N_17841,N_15303,N_14849);
nand U17842 (N_17842,N_14646,N_12823);
xnor U17843 (N_17843,N_12767,N_14692);
nor U17844 (N_17844,N_13079,N_14824);
or U17845 (N_17845,N_13924,N_13731);
or U17846 (N_17846,N_14001,N_15503);
nor U17847 (N_17847,N_15255,N_14921);
or U17848 (N_17848,N_12619,N_15112);
or U17849 (N_17849,N_12552,N_14807);
and U17850 (N_17850,N_15282,N_14247);
nor U17851 (N_17851,N_12650,N_15136);
or U17852 (N_17852,N_14643,N_14480);
nor U17853 (N_17853,N_14671,N_14431);
and U17854 (N_17854,N_14729,N_14134);
or U17855 (N_17855,N_13531,N_13234);
nand U17856 (N_17856,N_13804,N_14132);
nand U17857 (N_17857,N_15338,N_14773);
nand U17858 (N_17858,N_14037,N_12897);
and U17859 (N_17859,N_14811,N_14160);
nor U17860 (N_17860,N_14809,N_13503);
and U17861 (N_17861,N_14175,N_13425);
nand U17862 (N_17862,N_15236,N_13124);
or U17863 (N_17863,N_12608,N_12539);
or U17864 (N_17864,N_12836,N_12636);
nor U17865 (N_17865,N_15588,N_13407);
and U17866 (N_17866,N_15108,N_14994);
nor U17867 (N_17867,N_15274,N_13653);
xor U17868 (N_17868,N_14353,N_13399);
nor U17869 (N_17869,N_14468,N_12801);
nand U17870 (N_17870,N_14461,N_12806);
nor U17871 (N_17871,N_14038,N_13117);
xnor U17872 (N_17872,N_14588,N_13933);
nor U17873 (N_17873,N_13205,N_14118);
xor U17874 (N_17874,N_12757,N_13969);
nor U17875 (N_17875,N_13024,N_12775);
or U17876 (N_17876,N_14814,N_15057);
and U17877 (N_17877,N_13527,N_14415);
or U17878 (N_17878,N_13148,N_14788);
nor U17879 (N_17879,N_13674,N_14049);
xnor U17880 (N_17880,N_13919,N_14563);
xnor U17881 (N_17881,N_13331,N_12598);
xnor U17882 (N_17882,N_14667,N_14937);
nand U17883 (N_17883,N_13867,N_13333);
and U17884 (N_17884,N_14480,N_12893);
nand U17885 (N_17885,N_13591,N_13938);
nor U17886 (N_17886,N_14975,N_13548);
xor U17887 (N_17887,N_14011,N_12866);
and U17888 (N_17888,N_12904,N_15095);
nor U17889 (N_17889,N_13800,N_13667);
xor U17890 (N_17890,N_13981,N_12988);
and U17891 (N_17891,N_13286,N_15567);
or U17892 (N_17892,N_14396,N_12519);
nand U17893 (N_17893,N_14187,N_14326);
nand U17894 (N_17894,N_14135,N_13596);
nand U17895 (N_17895,N_14014,N_15418);
and U17896 (N_17896,N_14190,N_12631);
or U17897 (N_17897,N_13068,N_14613);
and U17898 (N_17898,N_14746,N_15380);
nor U17899 (N_17899,N_14187,N_14051);
xnor U17900 (N_17900,N_13230,N_13015);
nor U17901 (N_17901,N_12728,N_14256);
nor U17902 (N_17902,N_13381,N_13005);
or U17903 (N_17903,N_13925,N_13473);
xor U17904 (N_17904,N_15606,N_12926);
xnor U17905 (N_17905,N_12915,N_14676);
and U17906 (N_17906,N_13954,N_14678);
or U17907 (N_17907,N_13072,N_12610);
xnor U17908 (N_17908,N_15093,N_13502);
nor U17909 (N_17909,N_13890,N_14885);
xor U17910 (N_17910,N_15051,N_12587);
nand U17911 (N_17911,N_14640,N_13182);
xnor U17912 (N_17912,N_14699,N_15205);
nor U17913 (N_17913,N_13349,N_14283);
nor U17914 (N_17914,N_15066,N_14377);
nand U17915 (N_17915,N_15241,N_13634);
or U17916 (N_17916,N_14103,N_15146);
and U17917 (N_17917,N_13693,N_15264);
or U17918 (N_17918,N_14088,N_15588);
and U17919 (N_17919,N_15457,N_14301);
or U17920 (N_17920,N_14256,N_15030);
or U17921 (N_17921,N_14087,N_15287);
and U17922 (N_17922,N_14742,N_14365);
nor U17923 (N_17923,N_12533,N_12804);
and U17924 (N_17924,N_13316,N_14411);
or U17925 (N_17925,N_14601,N_13952);
or U17926 (N_17926,N_13574,N_13459);
nor U17927 (N_17927,N_14152,N_12844);
nor U17928 (N_17928,N_15135,N_12630);
nand U17929 (N_17929,N_14772,N_13920);
or U17930 (N_17930,N_14344,N_14174);
xor U17931 (N_17931,N_12967,N_14326);
nand U17932 (N_17932,N_15087,N_13037);
and U17933 (N_17933,N_13382,N_13391);
nor U17934 (N_17934,N_14702,N_15444);
and U17935 (N_17935,N_13730,N_13010);
nor U17936 (N_17936,N_14081,N_13628);
nor U17937 (N_17937,N_15271,N_14971);
and U17938 (N_17938,N_13956,N_13358);
xnor U17939 (N_17939,N_12741,N_15251);
xor U17940 (N_17940,N_13649,N_15311);
or U17941 (N_17941,N_15065,N_15135);
and U17942 (N_17942,N_14899,N_14617);
or U17943 (N_17943,N_13656,N_14973);
and U17944 (N_17944,N_15277,N_13562);
nand U17945 (N_17945,N_13134,N_15425);
or U17946 (N_17946,N_13118,N_14645);
xnor U17947 (N_17947,N_14760,N_15322);
and U17948 (N_17948,N_15185,N_14805);
and U17949 (N_17949,N_14708,N_13772);
nand U17950 (N_17950,N_13505,N_15206);
and U17951 (N_17951,N_14065,N_13609);
or U17952 (N_17952,N_14485,N_13639);
and U17953 (N_17953,N_14064,N_13282);
and U17954 (N_17954,N_12676,N_13783);
or U17955 (N_17955,N_13623,N_14047);
and U17956 (N_17956,N_14956,N_14427);
xor U17957 (N_17957,N_13696,N_12544);
nand U17958 (N_17958,N_13189,N_12775);
or U17959 (N_17959,N_13794,N_15080);
xor U17960 (N_17960,N_13731,N_13545);
nor U17961 (N_17961,N_15120,N_12688);
and U17962 (N_17962,N_12996,N_13044);
nand U17963 (N_17963,N_13066,N_13318);
nor U17964 (N_17964,N_13055,N_14355);
xnor U17965 (N_17965,N_14264,N_13785);
and U17966 (N_17966,N_13185,N_14651);
nand U17967 (N_17967,N_12977,N_14208);
nor U17968 (N_17968,N_13293,N_14364);
or U17969 (N_17969,N_14613,N_15531);
and U17970 (N_17970,N_13756,N_14731);
nand U17971 (N_17971,N_12529,N_12979);
nand U17972 (N_17972,N_14751,N_15140);
and U17973 (N_17973,N_15166,N_13083);
or U17974 (N_17974,N_12532,N_13745);
nand U17975 (N_17975,N_14584,N_12750);
nand U17976 (N_17976,N_14296,N_14144);
nor U17977 (N_17977,N_14631,N_13754);
xor U17978 (N_17978,N_13203,N_13552);
xor U17979 (N_17979,N_14823,N_15129);
nand U17980 (N_17980,N_12860,N_12828);
and U17981 (N_17981,N_15012,N_14857);
or U17982 (N_17982,N_14811,N_14703);
and U17983 (N_17983,N_14938,N_14092);
or U17984 (N_17984,N_13302,N_12836);
and U17985 (N_17985,N_14484,N_13366);
nand U17986 (N_17986,N_15103,N_12907);
nor U17987 (N_17987,N_15302,N_15023);
nand U17988 (N_17988,N_13187,N_13218);
xnor U17989 (N_17989,N_13218,N_13494);
nand U17990 (N_17990,N_14180,N_15097);
nor U17991 (N_17991,N_14807,N_14098);
nor U17992 (N_17992,N_15616,N_12553);
nand U17993 (N_17993,N_13318,N_13271);
and U17994 (N_17994,N_14579,N_12686);
nor U17995 (N_17995,N_12920,N_14771);
nor U17996 (N_17996,N_13743,N_14943);
and U17997 (N_17997,N_15256,N_14904);
nor U17998 (N_17998,N_15259,N_13469);
xnor U17999 (N_17999,N_14239,N_13040);
nor U18000 (N_18000,N_13514,N_14788);
xnor U18001 (N_18001,N_14163,N_12602);
or U18002 (N_18002,N_14869,N_15176);
or U18003 (N_18003,N_14099,N_14378);
nor U18004 (N_18004,N_15333,N_14092);
or U18005 (N_18005,N_14470,N_13744);
and U18006 (N_18006,N_15291,N_14499);
nor U18007 (N_18007,N_12584,N_12649);
nand U18008 (N_18008,N_14567,N_13606);
xor U18009 (N_18009,N_14489,N_14895);
nand U18010 (N_18010,N_13216,N_14289);
nor U18011 (N_18011,N_13851,N_13654);
or U18012 (N_18012,N_15523,N_14528);
nor U18013 (N_18013,N_15087,N_15259);
nand U18014 (N_18014,N_15534,N_15315);
nor U18015 (N_18015,N_15407,N_15446);
xor U18016 (N_18016,N_14716,N_13310);
nand U18017 (N_18017,N_13974,N_15624);
nand U18018 (N_18018,N_13333,N_14447);
or U18019 (N_18019,N_14166,N_13452);
or U18020 (N_18020,N_12796,N_14528);
or U18021 (N_18021,N_15327,N_15047);
or U18022 (N_18022,N_13936,N_15606);
or U18023 (N_18023,N_13974,N_13063);
nand U18024 (N_18024,N_14839,N_15577);
or U18025 (N_18025,N_12820,N_13478);
nor U18026 (N_18026,N_13586,N_13104);
nand U18027 (N_18027,N_14234,N_12682);
and U18028 (N_18028,N_13232,N_13678);
nor U18029 (N_18029,N_12952,N_14905);
and U18030 (N_18030,N_14822,N_13335);
or U18031 (N_18031,N_12941,N_13437);
nor U18032 (N_18032,N_15604,N_12612);
and U18033 (N_18033,N_14816,N_14087);
nand U18034 (N_18034,N_13558,N_15186);
nand U18035 (N_18035,N_14282,N_15577);
nor U18036 (N_18036,N_13600,N_15574);
and U18037 (N_18037,N_13310,N_13724);
nor U18038 (N_18038,N_15104,N_13857);
nand U18039 (N_18039,N_14004,N_12775);
xnor U18040 (N_18040,N_15360,N_14161);
nand U18041 (N_18041,N_12891,N_13153);
nor U18042 (N_18042,N_14822,N_15450);
and U18043 (N_18043,N_12718,N_12996);
xor U18044 (N_18044,N_15379,N_14292);
xnor U18045 (N_18045,N_12705,N_13559);
nor U18046 (N_18046,N_15266,N_15286);
nor U18047 (N_18047,N_12854,N_14695);
xnor U18048 (N_18048,N_15436,N_13523);
nand U18049 (N_18049,N_12887,N_13483);
or U18050 (N_18050,N_14236,N_14534);
nand U18051 (N_18051,N_13445,N_14330);
nor U18052 (N_18052,N_12869,N_13277);
and U18053 (N_18053,N_15259,N_13536);
nand U18054 (N_18054,N_14308,N_12620);
xor U18055 (N_18055,N_14740,N_13590);
xnor U18056 (N_18056,N_15402,N_15005);
nand U18057 (N_18057,N_15456,N_14408);
xor U18058 (N_18058,N_15474,N_14186);
or U18059 (N_18059,N_12993,N_13798);
and U18060 (N_18060,N_12757,N_15594);
nand U18061 (N_18061,N_13191,N_13821);
nand U18062 (N_18062,N_14902,N_15226);
and U18063 (N_18063,N_14811,N_14549);
nor U18064 (N_18064,N_12966,N_13774);
xor U18065 (N_18065,N_12976,N_14864);
xnor U18066 (N_18066,N_14028,N_14632);
nand U18067 (N_18067,N_14205,N_13958);
or U18068 (N_18068,N_14257,N_14413);
and U18069 (N_18069,N_15215,N_13002);
xor U18070 (N_18070,N_12702,N_14840);
nand U18071 (N_18071,N_14007,N_12562);
xor U18072 (N_18072,N_13456,N_13704);
nand U18073 (N_18073,N_12508,N_12561);
nor U18074 (N_18074,N_12691,N_14451);
or U18075 (N_18075,N_15283,N_15462);
nand U18076 (N_18076,N_14848,N_12520);
and U18077 (N_18077,N_13507,N_15097);
or U18078 (N_18078,N_13950,N_12694);
or U18079 (N_18079,N_14595,N_15518);
nor U18080 (N_18080,N_14281,N_12973);
or U18081 (N_18081,N_14486,N_13727);
nor U18082 (N_18082,N_15455,N_15550);
nor U18083 (N_18083,N_14153,N_13502);
and U18084 (N_18084,N_14082,N_14460);
or U18085 (N_18085,N_12540,N_15580);
nor U18086 (N_18086,N_13615,N_15436);
or U18087 (N_18087,N_14816,N_13273);
and U18088 (N_18088,N_15336,N_14249);
or U18089 (N_18089,N_14369,N_13553);
and U18090 (N_18090,N_14096,N_15199);
and U18091 (N_18091,N_13084,N_15432);
xnor U18092 (N_18092,N_15012,N_12553);
and U18093 (N_18093,N_15507,N_13468);
xor U18094 (N_18094,N_13185,N_14813);
nor U18095 (N_18095,N_12608,N_15377);
nand U18096 (N_18096,N_14908,N_14956);
nand U18097 (N_18097,N_14755,N_14094);
nand U18098 (N_18098,N_14873,N_13841);
nor U18099 (N_18099,N_14370,N_13912);
or U18100 (N_18100,N_15238,N_15289);
nand U18101 (N_18101,N_13632,N_12670);
and U18102 (N_18102,N_15129,N_12988);
or U18103 (N_18103,N_12681,N_12913);
xor U18104 (N_18104,N_12861,N_14497);
xor U18105 (N_18105,N_15313,N_14555);
nor U18106 (N_18106,N_15493,N_13475);
or U18107 (N_18107,N_13360,N_14658);
and U18108 (N_18108,N_12782,N_12777);
nor U18109 (N_18109,N_12848,N_14570);
xor U18110 (N_18110,N_12860,N_14732);
nor U18111 (N_18111,N_13164,N_15416);
and U18112 (N_18112,N_14554,N_15126);
or U18113 (N_18113,N_13993,N_14600);
nor U18114 (N_18114,N_15063,N_13745);
nor U18115 (N_18115,N_14526,N_14716);
and U18116 (N_18116,N_13746,N_15553);
xnor U18117 (N_18117,N_13452,N_15031);
and U18118 (N_18118,N_13824,N_14497);
xnor U18119 (N_18119,N_15098,N_13375);
nand U18120 (N_18120,N_14110,N_14573);
nor U18121 (N_18121,N_14133,N_12847);
and U18122 (N_18122,N_12662,N_14995);
or U18123 (N_18123,N_14236,N_14568);
or U18124 (N_18124,N_13757,N_13575);
and U18125 (N_18125,N_12573,N_13749);
nand U18126 (N_18126,N_14302,N_12989);
nor U18127 (N_18127,N_13052,N_12513);
nor U18128 (N_18128,N_15485,N_13053);
xnor U18129 (N_18129,N_13725,N_13698);
xor U18130 (N_18130,N_14404,N_15281);
nor U18131 (N_18131,N_13975,N_15023);
xnor U18132 (N_18132,N_14453,N_12775);
xor U18133 (N_18133,N_14166,N_13846);
nand U18134 (N_18134,N_15518,N_14153);
xor U18135 (N_18135,N_14181,N_14871);
nor U18136 (N_18136,N_14982,N_13682);
and U18137 (N_18137,N_13138,N_15605);
nand U18138 (N_18138,N_15081,N_13824);
or U18139 (N_18139,N_13165,N_13473);
or U18140 (N_18140,N_14903,N_15083);
nor U18141 (N_18141,N_13530,N_15147);
xnor U18142 (N_18142,N_14054,N_14466);
xnor U18143 (N_18143,N_12907,N_15548);
or U18144 (N_18144,N_15604,N_12977);
nor U18145 (N_18145,N_13085,N_13158);
or U18146 (N_18146,N_14955,N_13414);
nand U18147 (N_18147,N_12799,N_15087);
xnor U18148 (N_18148,N_15068,N_14043);
and U18149 (N_18149,N_12995,N_14065);
or U18150 (N_18150,N_14890,N_13876);
nand U18151 (N_18151,N_15428,N_13545);
and U18152 (N_18152,N_13895,N_12884);
and U18153 (N_18153,N_14996,N_13286);
or U18154 (N_18154,N_14347,N_15372);
or U18155 (N_18155,N_13213,N_12814);
and U18156 (N_18156,N_13821,N_14039);
nor U18157 (N_18157,N_13245,N_14410);
xnor U18158 (N_18158,N_15558,N_13681);
nor U18159 (N_18159,N_13916,N_13548);
nor U18160 (N_18160,N_15510,N_13771);
nor U18161 (N_18161,N_15563,N_13542);
nor U18162 (N_18162,N_14975,N_15584);
and U18163 (N_18163,N_13956,N_12670);
or U18164 (N_18164,N_15559,N_13145);
and U18165 (N_18165,N_14962,N_14873);
nor U18166 (N_18166,N_13419,N_15517);
nor U18167 (N_18167,N_14274,N_13022);
and U18168 (N_18168,N_14445,N_12943);
or U18169 (N_18169,N_14286,N_13607);
xor U18170 (N_18170,N_13166,N_12594);
or U18171 (N_18171,N_14553,N_13499);
nor U18172 (N_18172,N_14203,N_13191);
or U18173 (N_18173,N_13140,N_15586);
or U18174 (N_18174,N_15338,N_12802);
nand U18175 (N_18175,N_13773,N_14985);
and U18176 (N_18176,N_13436,N_15296);
nor U18177 (N_18177,N_14695,N_14156);
xor U18178 (N_18178,N_14090,N_12504);
and U18179 (N_18179,N_15367,N_15009);
and U18180 (N_18180,N_15222,N_13320);
nand U18181 (N_18181,N_14934,N_13257);
and U18182 (N_18182,N_15496,N_13159);
and U18183 (N_18183,N_14234,N_14291);
xor U18184 (N_18184,N_12516,N_12659);
or U18185 (N_18185,N_14678,N_12550);
nand U18186 (N_18186,N_13864,N_12871);
nand U18187 (N_18187,N_14399,N_15142);
xnor U18188 (N_18188,N_12791,N_14528);
nand U18189 (N_18189,N_14790,N_13551);
nand U18190 (N_18190,N_14672,N_14756);
xor U18191 (N_18191,N_13927,N_14434);
nor U18192 (N_18192,N_13810,N_14855);
or U18193 (N_18193,N_14643,N_12715);
or U18194 (N_18194,N_13702,N_13528);
nand U18195 (N_18195,N_13523,N_13800);
and U18196 (N_18196,N_15367,N_13390);
and U18197 (N_18197,N_15089,N_12688);
nor U18198 (N_18198,N_14005,N_14808);
xnor U18199 (N_18199,N_14982,N_13686);
or U18200 (N_18200,N_15012,N_15586);
or U18201 (N_18201,N_13396,N_13652);
xnor U18202 (N_18202,N_13518,N_13609);
or U18203 (N_18203,N_14601,N_14225);
nor U18204 (N_18204,N_13943,N_13101);
nand U18205 (N_18205,N_13483,N_14479);
nor U18206 (N_18206,N_14876,N_12875);
nand U18207 (N_18207,N_14130,N_14784);
xor U18208 (N_18208,N_15210,N_15425);
or U18209 (N_18209,N_13838,N_15019);
and U18210 (N_18210,N_12603,N_15526);
and U18211 (N_18211,N_14006,N_14587);
xor U18212 (N_18212,N_14056,N_13735);
xor U18213 (N_18213,N_15285,N_12818);
nor U18214 (N_18214,N_14312,N_14270);
xor U18215 (N_18215,N_12920,N_15513);
xor U18216 (N_18216,N_13547,N_13982);
nor U18217 (N_18217,N_12639,N_13290);
nor U18218 (N_18218,N_13638,N_12837);
nand U18219 (N_18219,N_12791,N_13876);
nand U18220 (N_18220,N_14333,N_14806);
nor U18221 (N_18221,N_14389,N_15247);
and U18222 (N_18222,N_13240,N_14265);
xor U18223 (N_18223,N_13463,N_14702);
nor U18224 (N_18224,N_13738,N_13162);
nor U18225 (N_18225,N_12993,N_14395);
xor U18226 (N_18226,N_14607,N_12713);
nand U18227 (N_18227,N_14822,N_12533);
and U18228 (N_18228,N_13033,N_13014);
and U18229 (N_18229,N_14950,N_14365);
nor U18230 (N_18230,N_15345,N_13507);
xor U18231 (N_18231,N_14461,N_15335);
or U18232 (N_18232,N_15238,N_14051);
xnor U18233 (N_18233,N_14447,N_12899);
xor U18234 (N_18234,N_14257,N_12710);
nor U18235 (N_18235,N_15318,N_13464);
xnor U18236 (N_18236,N_13030,N_14780);
nor U18237 (N_18237,N_15534,N_13201);
nor U18238 (N_18238,N_12674,N_13574);
or U18239 (N_18239,N_13990,N_12715);
or U18240 (N_18240,N_15276,N_13139);
nand U18241 (N_18241,N_15331,N_12969);
xnor U18242 (N_18242,N_14647,N_15179);
and U18243 (N_18243,N_13848,N_15024);
and U18244 (N_18244,N_15035,N_15218);
nand U18245 (N_18245,N_15524,N_13051);
or U18246 (N_18246,N_15377,N_13833);
nand U18247 (N_18247,N_12520,N_15061);
and U18248 (N_18248,N_12589,N_12534);
and U18249 (N_18249,N_14941,N_13911);
xnor U18250 (N_18250,N_12801,N_15373);
nand U18251 (N_18251,N_13604,N_14697);
nor U18252 (N_18252,N_12965,N_14543);
and U18253 (N_18253,N_12560,N_15429);
or U18254 (N_18254,N_15306,N_13526);
nor U18255 (N_18255,N_15326,N_14670);
nand U18256 (N_18256,N_12956,N_13447);
nor U18257 (N_18257,N_13323,N_14800);
nor U18258 (N_18258,N_14656,N_14698);
xor U18259 (N_18259,N_13394,N_15090);
nand U18260 (N_18260,N_14335,N_15003);
or U18261 (N_18261,N_13981,N_15598);
or U18262 (N_18262,N_14127,N_15110);
and U18263 (N_18263,N_13705,N_14628);
xnor U18264 (N_18264,N_14763,N_15129);
and U18265 (N_18265,N_14059,N_13173);
nor U18266 (N_18266,N_12751,N_14359);
nor U18267 (N_18267,N_14761,N_14194);
nand U18268 (N_18268,N_12997,N_14528);
and U18269 (N_18269,N_12929,N_14406);
or U18270 (N_18270,N_13529,N_14088);
xor U18271 (N_18271,N_13158,N_12852);
nand U18272 (N_18272,N_14898,N_13168);
nor U18273 (N_18273,N_14848,N_14583);
nand U18274 (N_18274,N_13095,N_12553);
or U18275 (N_18275,N_12796,N_13288);
or U18276 (N_18276,N_15350,N_13420);
nand U18277 (N_18277,N_14260,N_13175);
and U18278 (N_18278,N_13613,N_13774);
and U18279 (N_18279,N_12906,N_13349);
and U18280 (N_18280,N_15563,N_15584);
or U18281 (N_18281,N_13677,N_12917);
nor U18282 (N_18282,N_13893,N_12756);
nor U18283 (N_18283,N_14050,N_13023);
and U18284 (N_18284,N_13573,N_13314);
xnor U18285 (N_18285,N_12513,N_13398);
and U18286 (N_18286,N_12946,N_14035);
xnor U18287 (N_18287,N_13291,N_13879);
and U18288 (N_18288,N_14914,N_15603);
and U18289 (N_18289,N_12888,N_13978);
xnor U18290 (N_18290,N_14895,N_13132);
xor U18291 (N_18291,N_13942,N_14180);
nand U18292 (N_18292,N_12846,N_13258);
xor U18293 (N_18293,N_14207,N_12522);
or U18294 (N_18294,N_14738,N_15128);
and U18295 (N_18295,N_14890,N_13107);
nor U18296 (N_18296,N_13386,N_14032);
and U18297 (N_18297,N_12902,N_14642);
xnor U18298 (N_18298,N_14727,N_14899);
xnor U18299 (N_18299,N_13103,N_15369);
and U18300 (N_18300,N_12814,N_14068);
nand U18301 (N_18301,N_14634,N_15360);
or U18302 (N_18302,N_15437,N_13212);
nor U18303 (N_18303,N_14365,N_13137);
nor U18304 (N_18304,N_13289,N_14256);
or U18305 (N_18305,N_15258,N_14322);
nor U18306 (N_18306,N_14635,N_13398);
nand U18307 (N_18307,N_14902,N_13497);
nand U18308 (N_18308,N_15082,N_13464);
nor U18309 (N_18309,N_14681,N_15113);
and U18310 (N_18310,N_14616,N_13971);
and U18311 (N_18311,N_14965,N_15419);
and U18312 (N_18312,N_14902,N_15142);
nand U18313 (N_18313,N_15358,N_15224);
and U18314 (N_18314,N_15229,N_14505);
nand U18315 (N_18315,N_14455,N_14582);
xor U18316 (N_18316,N_12996,N_14738);
or U18317 (N_18317,N_15321,N_15444);
xnor U18318 (N_18318,N_15585,N_15582);
or U18319 (N_18319,N_12984,N_12568);
or U18320 (N_18320,N_13373,N_14013);
nand U18321 (N_18321,N_13521,N_14710);
or U18322 (N_18322,N_12844,N_15052);
and U18323 (N_18323,N_13102,N_13290);
or U18324 (N_18324,N_14777,N_13165);
nor U18325 (N_18325,N_12753,N_13224);
or U18326 (N_18326,N_14217,N_14731);
and U18327 (N_18327,N_14931,N_13839);
xor U18328 (N_18328,N_13598,N_13025);
and U18329 (N_18329,N_14764,N_14796);
xor U18330 (N_18330,N_14022,N_14880);
and U18331 (N_18331,N_14226,N_13835);
or U18332 (N_18332,N_15520,N_12994);
or U18333 (N_18333,N_13881,N_13870);
nand U18334 (N_18334,N_12532,N_13453);
xor U18335 (N_18335,N_13826,N_14036);
or U18336 (N_18336,N_13321,N_15133);
nand U18337 (N_18337,N_14282,N_15619);
and U18338 (N_18338,N_14705,N_14135);
nor U18339 (N_18339,N_13178,N_14127);
xnor U18340 (N_18340,N_15490,N_14403);
nor U18341 (N_18341,N_13780,N_14731);
or U18342 (N_18342,N_14606,N_13603);
xor U18343 (N_18343,N_13026,N_15271);
nor U18344 (N_18344,N_12812,N_14888);
or U18345 (N_18345,N_12665,N_13484);
nor U18346 (N_18346,N_13159,N_13988);
and U18347 (N_18347,N_15549,N_13059);
or U18348 (N_18348,N_14936,N_13027);
nand U18349 (N_18349,N_14403,N_13227);
nand U18350 (N_18350,N_12706,N_14760);
xor U18351 (N_18351,N_13857,N_12675);
and U18352 (N_18352,N_13844,N_14629);
or U18353 (N_18353,N_15131,N_12555);
nor U18354 (N_18354,N_12722,N_14222);
xor U18355 (N_18355,N_15017,N_12812);
and U18356 (N_18356,N_15001,N_12909);
xor U18357 (N_18357,N_15234,N_14589);
or U18358 (N_18358,N_12995,N_14157);
nor U18359 (N_18359,N_13776,N_15544);
and U18360 (N_18360,N_14892,N_12656);
nor U18361 (N_18361,N_14390,N_13375);
or U18362 (N_18362,N_13925,N_12594);
and U18363 (N_18363,N_15282,N_15092);
and U18364 (N_18364,N_13915,N_13772);
nor U18365 (N_18365,N_14900,N_15306);
nor U18366 (N_18366,N_14375,N_14042);
xor U18367 (N_18367,N_14151,N_14137);
or U18368 (N_18368,N_13605,N_12557);
xor U18369 (N_18369,N_15596,N_13903);
nor U18370 (N_18370,N_12505,N_15170);
xnor U18371 (N_18371,N_15210,N_14393);
and U18372 (N_18372,N_13498,N_14110);
nor U18373 (N_18373,N_14117,N_13168);
nor U18374 (N_18374,N_15539,N_15359);
nor U18375 (N_18375,N_14234,N_13924);
nor U18376 (N_18376,N_14430,N_15291);
xnor U18377 (N_18377,N_13816,N_14733);
nand U18378 (N_18378,N_15319,N_13451);
or U18379 (N_18379,N_14768,N_12631);
xor U18380 (N_18380,N_14021,N_13420);
and U18381 (N_18381,N_14586,N_15352);
nand U18382 (N_18382,N_12689,N_14234);
and U18383 (N_18383,N_14490,N_13131);
nand U18384 (N_18384,N_14945,N_12976);
and U18385 (N_18385,N_15495,N_12760);
and U18386 (N_18386,N_13626,N_13810);
and U18387 (N_18387,N_15489,N_14947);
and U18388 (N_18388,N_13362,N_12762);
nand U18389 (N_18389,N_13156,N_14090);
or U18390 (N_18390,N_15125,N_14832);
nor U18391 (N_18391,N_12660,N_15045);
and U18392 (N_18392,N_14968,N_13500);
or U18393 (N_18393,N_12667,N_13621);
nand U18394 (N_18394,N_12549,N_13221);
xor U18395 (N_18395,N_15407,N_13077);
and U18396 (N_18396,N_13790,N_13989);
nor U18397 (N_18397,N_13407,N_13439);
nor U18398 (N_18398,N_14381,N_14983);
nand U18399 (N_18399,N_15561,N_13478);
nor U18400 (N_18400,N_13006,N_12714);
nor U18401 (N_18401,N_12597,N_12538);
and U18402 (N_18402,N_13295,N_14976);
nand U18403 (N_18403,N_12536,N_14053);
nor U18404 (N_18404,N_13377,N_12659);
nand U18405 (N_18405,N_12864,N_15139);
or U18406 (N_18406,N_13445,N_15529);
and U18407 (N_18407,N_14261,N_12588);
or U18408 (N_18408,N_13615,N_13171);
nand U18409 (N_18409,N_14365,N_15006);
nor U18410 (N_18410,N_14296,N_13725);
nor U18411 (N_18411,N_13860,N_13981);
nor U18412 (N_18412,N_12819,N_14816);
xor U18413 (N_18413,N_14909,N_15180);
and U18414 (N_18414,N_13802,N_13804);
xnor U18415 (N_18415,N_14575,N_15185);
and U18416 (N_18416,N_13777,N_14206);
nor U18417 (N_18417,N_14760,N_12858);
nor U18418 (N_18418,N_14842,N_15375);
nand U18419 (N_18419,N_15573,N_14774);
and U18420 (N_18420,N_14958,N_15381);
xor U18421 (N_18421,N_15574,N_15082);
or U18422 (N_18422,N_12649,N_13139);
or U18423 (N_18423,N_15251,N_13215);
or U18424 (N_18424,N_13966,N_13407);
and U18425 (N_18425,N_15100,N_15127);
and U18426 (N_18426,N_14434,N_12966);
nand U18427 (N_18427,N_13654,N_13186);
xnor U18428 (N_18428,N_13061,N_13985);
xnor U18429 (N_18429,N_14374,N_13192);
or U18430 (N_18430,N_12518,N_15005);
or U18431 (N_18431,N_13220,N_14696);
and U18432 (N_18432,N_13349,N_14920);
xor U18433 (N_18433,N_12848,N_13662);
or U18434 (N_18434,N_14697,N_12725);
nand U18435 (N_18435,N_15083,N_13547);
nand U18436 (N_18436,N_15174,N_14012);
nand U18437 (N_18437,N_13352,N_14565);
nor U18438 (N_18438,N_12637,N_13714);
and U18439 (N_18439,N_12573,N_14127);
nand U18440 (N_18440,N_12608,N_14984);
nand U18441 (N_18441,N_14912,N_13833);
xnor U18442 (N_18442,N_15263,N_13361);
nand U18443 (N_18443,N_14823,N_14975);
xor U18444 (N_18444,N_14512,N_14290);
and U18445 (N_18445,N_14974,N_14337);
or U18446 (N_18446,N_13002,N_15483);
and U18447 (N_18447,N_14843,N_13167);
or U18448 (N_18448,N_14519,N_14099);
nand U18449 (N_18449,N_14922,N_12501);
nand U18450 (N_18450,N_15167,N_14350);
and U18451 (N_18451,N_14670,N_13772);
and U18452 (N_18452,N_14715,N_14433);
or U18453 (N_18453,N_13906,N_12706);
or U18454 (N_18454,N_12760,N_13028);
nand U18455 (N_18455,N_14627,N_13154);
nor U18456 (N_18456,N_12965,N_15374);
nor U18457 (N_18457,N_14959,N_14381);
nor U18458 (N_18458,N_12747,N_14216);
nor U18459 (N_18459,N_14323,N_13962);
or U18460 (N_18460,N_15499,N_13186);
and U18461 (N_18461,N_12620,N_14468);
and U18462 (N_18462,N_15055,N_13612);
xor U18463 (N_18463,N_13244,N_13345);
nor U18464 (N_18464,N_12543,N_15254);
xor U18465 (N_18465,N_15492,N_15373);
or U18466 (N_18466,N_12963,N_12827);
xor U18467 (N_18467,N_14515,N_15288);
nand U18468 (N_18468,N_13196,N_13277);
nor U18469 (N_18469,N_15103,N_13487);
nor U18470 (N_18470,N_15579,N_13090);
xor U18471 (N_18471,N_14454,N_13779);
nand U18472 (N_18472,N_13871,N_13086);
xor U18473 (N_18473,N_13093,N_12740);
nor U18474 (N_18474,N_15404,N_15078);
nor U18475 (N_18475,N_15382,N_14959);
nand U18476 (N_18476,N_13475,N_15100);
and U18477 (N_18477,N_14925,N_13280);
nor U18478 (N_18478,N_13844,N_13723);
nand U18479 (N_18479,N_14305,N_13993);
nor U18480 (N_18480,N_15564,N_14559);
nand U18481 (N_18481,N_14199,N_13189);
nor U18482 (N_18482,N_12968,N_13902);
nand U18483 (N_18483,N_15440,N_12540);
and U18484 (N_18484,N_12552,N_15026);
or U18485 (N_18485,N_15174,N_15522);
xor U18486 (N_18486,N_15317,N_13615);
and U18487 (N_18487,N_14843,N_12739);
xnor U18488 (N_18488,N_15178,N_14086);
nand U18489 (N_18489,N_13796,N_12719);
and U18490 (N_18490,N_15243,N_15070);
xnor U18491 (N_18491,N_14487,N_14657);
or U18492 (N_18492,N_13349,N_13048);
nor U18493 (N_18493,N_13734,N_13626);
or U18494 (N_18494,N_12924,N_15246);
and U18495 (N_18495,N_14101,N_14481);
nor U18496 (N_18496,N_14670,N_14162);
or U18497 (N_18497,N_13352,N_15273);
nor U18498 (N_18498,N_15196,N_13016);
nor U18499 (N_18499,N_14070,N_13654);
xnor U18500 (N_18500,N_15306,N_14447);
nor U18501 (N_18501,N_13963,N_14000);
nor U18502 (N_18502,N_14520,N_14972);
nor U18503 (N_18503,N_14543,N_14168);
nand U18504 (N_18504,N_15309,N_15102);
nand U18505 (N_18505,N_13624,N_13008);
xor U18506 (N_18506,N_12806,N_12538);
or U18507 (N_18507,N_14643,N_13809);
nand U18508 (N_18508,N_14037,N_14865);
and U18509 (N_18509,N_14996,N_15512);
nor U18510 (N_18510,N_12882,N_15068);
nor U18511 (N_18511,N_13131,N_13120);
nor U18512 (N_18512,N_14830,N_14614);
or U18513 (N_18513,N_15533,N_13313);
or U18514 (N_18514,N_15324,N_13608);
nor U18515 (N_18515,N_12674,N_14201);
nand U18516 (N_18516,N_13630,N_14077);
and U18517 (N_18517,N_12564,N_13379);
or U18518 (N_18518,N_15519,N_14456);
nand U18519 (N_18519,N_15144,N_13145);
or U18520 (N_18520,N_15078,N_14233);
and U18521 (N_18521,N_15255,N_12622);
nand U18522 (N_18522,N_13455,N_14791);
nand U18523 (N_18523,N_15081,N_12524);
nand U18524 (N_18524,N_14598,N_15065);
and U18525 (N_18525,N_14495,N_12893);
nor U18526 (N_18526,N_13430,N_14084);
and U18527 (N_18527,N_15018,N_14734);
and U18528 (N_18528,N_14361,N_14329);
or U18529 (N_18529,N_15355,N_13466);
and U18530 (N_18530,N_13369,N_13826);
xnor U18531 (N_18531,N_13939,N_15034);
nand U18532 (N_18532,N_12547,N_15088);
xor U18533 (N_18533,N_15384,N_14279);
nor U18534 (N_18534,N_12577,N_15237);
nor U18535 (N_18535,N_13990,N_13238);
nand U18536 (N_18536,N_14399,N_15021);
or U18537 (N_18537,N_14841,N_13504);
xnor U18538 (N_18538,N_15328,N_15238);
nor U18539 (N_18539,N_13088,N_14554);
nand U18540 (N_18540,N_14237,N_13634);
nand U18541 (N_18541,N_14553,N_13121);
and U18542 (N_18542,N_15239,N_13921);
and U18543 (N_18543,N_13094,N_15483);
xnor U18544 (N_18544,N_14947,N_12524);
nor U18545 (N_18545,N_14538,N_15281);
or U18546 (N_18546,N_12667,N_12818);
and U18547 (N_18547,N_13739,N_14159);
xor U18548 (N_18548,N_13936,N_13525);
nand U18549 (N_18549,N_12976,N_13678);
or U18550 (N_18550,N_14504,N_14033);
and U18551 (N_18551,N_13969,N_14119);
nor U18552 (N_18552,N_13459,N_15349);
and U18553 (N_18553,N_12667,N_13963);
xor U18554 (N_18554,N_15307,N_12993);
or U18555 (N_18555,N_15399,N_13105);
and U18556 (N_18556,N_14466,N_13680);
nand U18557 (N_18557,N_13938,N_13039);
nand U18558 (N_18558,N_15373,N_14105);
and U18559 (N_18559,N_13424,N_13944);
nor U18560 (N_18560,N_14514,N_15031);
nor U18561 (N_18561,N_13912,N_14686);
and U18562 (N_18562,N_14060,N_12728);
or U18563 (N_18563,N_12535,N_13712);
and U18564 (N_18564,N_13885,N_14093);
and U18565 (N_18565,N_12934,N_13684);
or U18566 (N_18566,N_13326,N_15059);
nor U18567 (N_18567,N_13794,N_14657);
xnor U18568 (N_18568,N_15305,N_14628);
xor U18569 (N_18569,N_15335,N_13448);
or U18570 (N_18570,N_14849,N_14898);
and U18571 (N_18571,N_12847,N_13440);
and U18572 (N_18572,N_14718,N_15455);
and U18573 (N_18573,N_13448,N_13379);
nand U18574 (N_18574,N_15442,N_14630);
nor U18575 (N_18575,N_15121,N_12709);
xor U18576 (N_18576,N_13740,N_13906);
nand U18577 (N_18577,N_13550,N_13233);
nor U18578 (N_18578,N_14360,N_14180);
nand U18579 (N_18579,N_15190,N_13282);
or U18580 (N_18580,N_12981,N_15544);
xnor U18581 (N_18581,N_12671,N_14986);
nand U18582 (N_18582,N_12784,N_12518);
or U18583 (N_18583,N_13253,N_13040);
and U18584 (N_18584,N_13919,N_15412);
nor U18585 (N_18585,N_13132,N_15613);
or U18586 (N_18586,N_13859,N_13794);
xor U18587 (N_18587,N_12727,N_13068);
or U18588 (N_18588,N_12786,N_15270);
nand U18589 (N_18589,N_13482,N_13923);
and U18590 (N_18590,N_14421,N_14545);
xnor U18591 (N_18591,N_14373,N_13345);
nor U18592 (N_18592,N_15101,N_14955);
or U18593 (N_18593,N_14791,N_13644);
or U18594 (N_18594,N_13116,N_13392);
nand U18595 (N_18595,N_14863,N_13861);
nand U18596 (N_18596,N_13765,N_15276);
xor U18597 (N_18597,N_14961,N_14617);
xnor U18598 (N_18598,N_14947,N_15209);
nand U18599 (N_18599,N_13229,N_12546);
and U18600 (N_18600,N_14974,N_13307);
xor U18601 (N_18601,N_12950,N_13353);
and U18602 (N_18602,N_13581,N_13332);
nor U18603 (N_18603,N_15256,N_14962);
nor U18604 (N_18604,N_12696,N_12939);
xor U18605 (N_18605,N_13231,N_12946);
xnor U18606 (N_18606,N_13677,N_14792);
xor U18607 (N_18607,N_15386,N_14791);
and U18608 (N_18608,N_12962,N_14222);
nor U18609 (N_18609,N_13348,N_14489);
or U18610 (N_18610,N_15301,N_13244);
and U18611 (N_18611,N_12882,N_14188);
or U18612 (N_18612,N_12662,N_14953);
nor U18613 (N_18613,N_12965,N_14975);
or U18614 (N_18614,N_14020,N_13778);
nor U18615 (N_18615,N_15134,N_12710);
nand U18616 (N_18616,N_12577,N_13616);
nand U18617 (N_18617,N_13087,N_12841);
and U18618 (N_18618,N_14644,N_14965);
nand U18619 (N_18619,N_15372,N_13896);
nand U18620 (N_18620,N_13733,N_14581);
or U18621 (N_18621,N_14085,N_12759);
or U18622 (N_18622,N_14684,N_14365);
and U18623 (N_18623,N_12531,N_13714);
nor U18624 (N_18624,N_13688,N_13006);
and U18625 (N_18625,N_14563,N_14306);
nand U18626 (N_18626,N_13290,N_15158);
and U18627 (N_18627,N_15048,N_13058);
nor U18628 (N_18628,N_12839,N_14254);
or U18629 (N_18629,N_12879,N_14187);
nand U18630 (N_18630,N_12584,N_15374);
and U18631 (N_18631,N_14829,N_14362);
xor U18632 (N_18632,N_13516,N_14700);
or U18633 (N_18633,N_14554,N_13729);
and U18634 (N_18634,N_14777,N_14467);
and U18635 (N_18635,N_15236,N_15134);
or U18636 (N_18636,N_14489,N_14498);
and U18637 (N_18637,N_15433,N_15162);
nand U18638 (N_18638,N_14028,N_14338);
xnor U18639 (N_18639,N_14992,N_12682);
xnor U18640 (N_18640,N_14433,N_13012);
or U18641 (N_18641,N_13679,N_13463);
and U18642 (N_18642,N_14601,N_15497);
nor U18643 (N_18643,N_14249,N_13630);
and U18644 (N_18644,N_15194,N_14301);
nor U18645 (N_18645,N_12917,N_14456);
nand U18646 (N_18646,N_13597,N_15538);
or U18647 (N_18647,N_13372,N_13874);
xor U18648 (N_18648,N_12546,N_14644);
xnor U18649 (N_18649,N_13234,N_14324);
and U18650 (N_18650,N_14089,N_15482);
nand U18651 (N_18651,N_15194,N_12892);
nor U18652 (N_18652,N_15099,N_13431);
xnor U18653 (N_18653,N_13099,N_12922);
nand U18654 (N_18654,N_12642,N_14386);
xnor U18655 (N_18655,N_14173,N_13337);
or U18656 (N_18656,N_14212,N_12922);
xor U18657 (N_18657,N_14983,N_12899);
and U18658 (N_18658,N_13528,N_15192);
or U18659 (N_18659,N_15283,N_15157);
nor U18660 (N_18660,N_14793,N_14442);
or U18661 (N_18661,N_13327,N_13731);
or U18662 (N_18662,N_13088,N_14309);
xnor U18663 (N_18663,N_12959,N_12906);
nor U18664 (N_18664,N_14672,N_15486);
nand U18665 (N_18665,N_12970,N_13587);
nand U18666 (N_18666,N_13740,N_13398);
nand U18667 (N_18667,N_15509,N_14092);
and U18668 (N_18668,N_13586,N_15052);
nor U18669 (N_18669,N_15266,N_13510);
and U18670 (N_18670,N_15435,N_14528);
nand U18671 (N_18671,N_15287,N_13998);
and U18672 (N_18672,N_14685,N_13967);
xnor U18673 (N_18673,N_13441,N_14321);
or U18674 (N_18674,N_15129,N_14025);
xnor U18675 (N_18675,N_13843,N_14335);
and U18676 (N_18676,N_15059,N_12842);
nand U18677 (N_18677,N_13889,N_14764);
xor U18678 (N_18678,N_15566,N_14171);
or U18679 (N_18679,N_12948,N_15060);
nand U18680 (N_18680,N_12824,N_15183);
or U18681 (N_18681,N_13097,N_14038);
xor U18682 (N_18682,N_13176,N_12958);
xnor U18683 (N_18683,N_15207,N_14920);
xor U18684 (N_18684,N_14141,N_15613);
nand U18685 (N_18685,N_14766,N_15173);
and U18686 (N_18686,N_14877,N_15031);
or U18687 (N_18687,N_15117,N_12998);
nor U18688 (N_18688,N_13683,N_14887);
nand U18689 (N_18689,N_12554,N_13333);
nor U18690 (N_18690,N_13187,N_13603);
or U18691 (N_18691,N_13861,N_14427);
nor U18692 (N_18692,N_13265,N_14614);
nor U18693 (N_18693,N_13019,N_13040);
nor U18694 (N_18694,N_14980,N_15394);
nand U18695 (N_18695,N_12572,N_12768);
nand U18696 (N_18696,N_14075,N_14007);
nand U18697 (N_18697,N_14313,N_13636);
nand U18698 (N_18698,N_14428,N_13947);
xnor U18699 (N_18699,N_14100,N_15287);
or U18700 (N_18700,N_14561,N_14182);
nor U18701 (N_18701,N_12735,N_14445);
and U18702 (N_18702,N_13336,N_13113);
nor U18703 (N_18703,N_14415,N_15050);
and U18704 (N_18704,N_14795,N_14876);
or U18705 (N_18705,N_13610,N_14439);
xor U18706 (N_18706,N_14915,N_13713);
and U18707 (N_18707,N_15087,N_15473);
nor U18708 (N_18708,N_12725,N_14155);
and U18709 (N_18709,N_13705,N_13630);
and U18710 (N_18710,N_14146,N_14036);
xor U18711 (N_18711,N_13160,N_14170);
nor U18712 (N_18712,N_14122,N_13802);
and U18713 (N_18713,N_12913,N_12518);
nor U18714 (N_18714,N_15359,N_13847);
xnor U18715 (N_18715,N_13338,N_15488);
nand U18716 (N_18716,N_12944,N_13289);
nand U18717 (N_18717,N_14350,N_13863);
and U18718 (N_18718,N_13930,N_15112);
nor U18719 (N_18719,N_13356,N_13232);
and U18720 (N_18720,N_13610,N_14965);
and U18721 (N_18721,N_13894,N_14751);
or U18722 (N_18722,N_13613,N_13059);
or U18723 (N_18723,N_13535,N_14002);
nand U18724 (N_18724,N_14580,N_12531);
xor U18725 (N_18725,N_13228,N_12618);
and U18726 (N_18726,N_14854,N_12524);
or U18727 (N_18727,N_13206,N_12612);
and U18728 (N_18728,N_13802,N_15342);
or U18729 (N_18729,N_15000,N_15574);
or U18730 (N_18730,N_14402,N_13472);
nor U18731 (N_18731,N_13022,N_14806);
nor U18732 (N_18732,N_15014,N_14259);
nor U18733 (N_18733,N_14514,N_13287);
xor U18734 (N_18734,N_14170,N_15556);
nand U18735 (N_18735,N_13201,N_13816);
and U18736 (N_18736,N_13090,N_14749);
nand U18737 (N_18737,N_14392,N_13211);
nor U18738 (N_18738,N_15340,N_12745);
xnor U18739 (N_18739,N_14370,N_14033);
nor U18740 (N_18740,N_12524,N_15003);
and U18741 (N_18741,N_12904,N_15406);
nand U18742 (N_18742,N_14354,N_12556);
xnor U18743 (N_18743,N_14218,N_15135);
nand U18744 (N_18744,N_14023,N_12620);
and U18745 (N_18745,N_13075,N_13389);
xor U18746 (N_18746,N_13679,N_13274);
nand U18747 (N_18747,N_14957,N_14399);
or U18748 (N_18748,N_15196,N_13338);
nor U18749 (N_18749,N_15499,N_13329);
nand U18750 (N_18750,N_18565,N_15770);
nand U18751 (N_18751,N_15669,N_15916);
or U18752 (N_18752,N_18733,N_16562);
xor U18753 (N_18753,N_17915,N_16393);
nor U18754 (N_18754,N_18745,N_16850);
or U18755 (N_18755,N_17738,N_18187);
xnor U18756 (N_18756,N_18603,N_18705);
xor U18757 (N_18757,N_15924,N_16495);
nor U18758 (N_18758,N_18381,N_18612);
nor U18759 (N_18759,N_16711,N_15719);
or U18760 (N_18760,N_15922,N_18685);
or U18761 (N_18761,N_17778,N_17917);
nand U18762 (N_18762,N_16667,N_17544);
and U18763 (N_18763,N_17559,N_16568);
xnor U18764 (N_18764,N_15646,N_18416);
and U18765 (N_18765,N_17894,N_17398);
nand U18766 (N_18766,N_18614,N_16143);
nor U18767 (N_18767,N_16808,N_18445);
nor U18768 (N_18768,N_18472,N_16602);
xor U18769 (N_18769,N_18332,N_16512);
and U18770 (N_18770,N_17522,N_16194);
nand U18771 (N_18771,N_18376,N_17085);
nor U18772 (N_18772,N_16122,N_15845);
and U18773 (N_18773,N_16878,N_18465);
nand U18774 (N_18774,N_17172,N_16572);
xnor U18775 (N_18775,N_15988,N_15907);
xnor U18776 (N_18776,N_17184,N_16539);
nor U18777 (N_18777,N_18575,N_15807);
or U18778 (N_18778,N_17923,N_16229);
xnor U18779 (N_18779,N_18741,N_16774);
nand U18780 (N_18780,N_16396,N_18353);
and U18781 (N_18781,N_17862,N_17850);
or U18782 (N_18782,N_18667,N_17325);
and U18783 (N_18783,N_18660,N_16281);
xor U18784 (N_18784,N_18724,N_16471);
nor U18785 (N_18785,N_17821,N_15911);
or U18786 (N_18786,N_17889,N_16849);
and U18787 (N_18787,N_15681,N_18721);
or U18788 (N_18788,N_16675,N_16177);
and U18789 (N_18789,N_18483,N_16155);
nand U18790 (N_18790,N_18170,N_16172);
nand U18791 (N_18791,N_17379,N_17277);
nor U18792 (N_18792,N_16296,N_16438);
nand U18793 (N_18793,N_16875,N_16334);
xor U18794 (N_18794,N_16635,N_16534);
nand U18795 (N_18795,N_18282,N_15730);
xnor U18796 (N_18796,N_18340,N_17956);
and U18797 (N_18797,N_18456,N_17471);
or U18798 (N_18798,N_18380,N_16966);
nand U18799 (N_18799,N_18028,N_15634);
nand U18800 (N_18800,N_18108,N_18296);
nand U18801 (N_18801,N_18392,N_17273);
nor U18802 (N_18802,N_15952,N_16069);
nand U18803 (N_18803,N_16030,N_16744);
nor U18804 (N_18804,N_16307,N_16874);
and U18805 (N_18805,N_18163,N_15731);
xor U18806 (N_18806,N_16517,N_16932);
nor U18807 (N_18807,N_18396,N_18375);
or U18808 (N_18808,N_16792,N_15836);
nor U18809 (N_18809,N_16333,N_16518);
nand U18810 (N_18810,N_18540,N_15741);
nand U18811 (N_18811,N_17762,N_17620);
nand U18812 (N_18812,N_16059,N_18179);
nand U18813 (N_18813,N_15991,N_16825);
and U18814 (N_18814,N_17008,N_18084);
or U18815 (N_18815,N_15860,N_17390);
xor U18816 (N_18816,N_17797,N_17427);
or U18817 (N_18817,N_16599,N_17100);
or U18818 (N_18818,N_16315,N_18434);
and U18819 (N_18819,N_16713,N_16452);
nand U18820 (N_18820,N_15961,N_16513);
xnor U18821 (N_18821,N_16592,N_17053);
xor U18822 (N_18822,N_17310,N_16530);
xor U18823 (N_18823,N_16862,N_18387);
nand U18824 (N_18824,N_17510,N_16482);
and U18825 (N_18825,N_16734,N_16113);
nor U18826 (N_18826,N_17947,N_17927);
or U18827 (N_18827,N_17959,N_17474);
xnor U18828 (N_18828,N_16945,N_16853);
nand U18829 (N_18829,N_16654,N_18219);
nand U18830 (N_18830,N_17918,N_17714);
xor U18831 (N_18831,N_17105,N_16662);
and U18832 (N_18832,N_16048,N_17384);
and U18833 (N_18833,N_16876,N_17609);
and U18834 (N_18834,N_17642,N_16695);
nand U18835 (N_18835,N_17146,N_17148);
nor U18836 (N_18836,N_18127,N_16623);
and U18837 (N_18837,N_18176,N_15673);
xor U18838 (N_18838,N_18089,N_17088);
xnor U18839 (N_18839,N_17244,N_18671);
or U18840 (N_18840,N_16532,N_16802);
nor U18841 (N_18841,N_17176,N_18617);
nand U18842 (N_18842,N_18659,N_16724);
nand U18843 (N_18843,N_18645,N_15931);
or U18844 (N_18844,N_16410,N_16103);
or U18845 (N_18845,N_16392,N_16362);
and U18846 (N_18846,N_17162,N_17689);
or U18847 (N_18847,N_16761,N_16897);
nor U18848 (N_18848,N_16598,N_18679);
xor U18849 (N_18849,N_16244,N_16644);
nand U18850 (N_18850,N_16310,N_17648);
or U18851 (N_18851,N_16264,N_17879);
nand U18852 (N_18852,N_18169,N_16573);
xnor U18853 (N_18853,N_17473,N_18528);
nand U18854 (N_18854,N_18083,N_17216);
nand U18855 (N_18855,N_16201,N_18443);
and U18856 (N_18856,N_16917,N_15917);
nor U18857 (N_18857,N_15781,N_18099);
nor U18858 (N_18858,N_17909,N_17854);
xnor U18859 (N_18859,N_18607,N_16721);
or U18860 (N_18860,N_18135,N_18501);
or U18861 (N_18861,N_17932,N_17316);
or U18862 (N_18862,N_18742,N_18735);
or U18863 (N_18863,N_18041,N_17723);
nand U18864 (N_18864,N_17577,N_16273);
nand U18865 (N_18865,N_16492,N_16961);
or U18866 (N_18866,N_17010,N_17436);
nor U18867 (N_18867,N_16274,N_17367);
or U18868 (N_18868,N_18286,N_16451);
xnor U18869 (N_18869,N_18715,N_17170);
nor U18870 (N_18870,N_18009,N_18585);
and U18871 (N_18871,N_16367,N_18520);
and U18872 (N_18872,N_18299,N_17291);
nor U18873 (N_18873,N_17371,N_17940);
xnor U18874 (N_18874,N_17394,N_17814);
nand U18875 (N_18875,N_15814,N_16004);
xor U18876 (N_18876,N_15754,N_15633);
nor U18877 (N_18877,N_16268,N_16054);
nand U18878 (N_18878,N_15829,N_16361);
nand U18879 (N_18879,N_17783,N_18466);
nor U18880 (N_18880,N_17406,N_16081);
xor U18881 (N_18881,N_15838,N_18657);
or U18882 (N_18882,N_15759,N_17449);
nand U18883 (N_18883,N_18019,N_16949);
nor U18884 (N_18884,N_16123,N_17518);
or U18885 (N_18885,N_16223,N_17054);
xor U18886 (N_18886,N_18419,N_15839);
or U18887 (N_18887,N_18577,N_15958);
nor U18888 (N_18888,N_17736,N_18251);
nand U18889 (N_18889,N_17952,N_16204);
nor U18890 (N_18890,N_16360,N_15785);
xnor U18891 (N_18891,N_18271,N_17426);
nor U18892 (N_18892,N_16319,N_16678);
nand U18893 (N_18893,N_17865,N_17327);
nand U18894 (N_18894,N_18687,N_18345);
nor U18895 (N_18895,N_17283,N_16009);
or U18896 (N_18896,N_17536,N_17167);
nor U18897 (N_18897,N_16570,N_17635);
xnor U18898 (N_18898,N_17305,N_18228);
nor U18899 (N_18899,N_17663,N_17037);
nand U18900 (N_18900,N_18648,N_15682);
nand U18901 (N_18901,N_18712,N_18067);
or U18902 (N_18902,N_17122,N_16835);
nand U18903 (N_18903,N_17207,N_16363);
nand U18904 (N_18904,N_15935,N_16869);
nor U18905 (N_18905,N_16720,N_16659);
nor U18906 (N_18906,N_16984,N_15626);
nand U18907 (N_18907,N_18634,N_16558);
nand U18908 (N_18908,N_18273,N_17684);
or U18909 (N_18909,N_16205,N_16098);
nand U18910 (N_18910,N_15908,N_16390);
or U18911 (N_18911,N_17898,N_18427);
nand U18912 (N_18912,N_17389,N_17882);
or U18913 (N_18913,N_16557,N_18235);
nand U18914 (N_18914,N_16769,N_17951);
and U18915 (N_18915,N_18018,N_17351);
nor U18916 (N_18916,N_17086,N_18482);
nor U18917 (N_18917,N_15992,N_17154);
and U18918 (N_18918,N_17653,N_16737);
and U18919 (N_18919,N_18088,N_16981);
nor U18920 (N_18920,N_18233,N_16655);
nor U18921 (N_18921,N_18126,N_16236);
xor U18922 (N_18922,N_16070,N_18319);
nand U18923 (N_18923,N_16292,N_17715);
nor U18924 (N_18924,N_17140,N_15885);
nor U18925 (N_18925,N_17751,N_15960);
and U18926 (N_18926,N_16506,N_16186);
nand U18927 (N_18927,N_15930,N_16752);
nand U18928 (N_18928,N_18312,N_16941);
nand U18929 (N_18929,N_16826,N_17571);
or U18930 (N_18930,N_16794,N_16082);
and U18931 (N_18931,N_16107,N_18452);
or U18932 (N_18932,N_17464,N_15904);
or U18933 (N_18933,N_17914,N_15756);
xor U18934 (N_18934,N_17841,N_18622);
nand U18935 (N_18935,N_16439,N_16262);
nor U18936 (N_18936,N_16339,N_18277);
xnor U18937 (N_18937,N_17247,N_16388);
and U18938 (N_18938,N_18238,N_16852);
xnor U18939 (N_18939,N_18304,N_17455);
nand U18940 (N_18940,N_16609,N_17324);
nand U18941 (N_18941,N_18439,N_17666);
or U18942 (N_18942,N_15969,N_18664);
nand U18943 (N_18943,N_18406,N_18599);
and U18944 (N_18944,N_15914,N_16096);
nand U18945 (N_18945,N_17144,N_18682);
xor U18946 (N_18946,N_18409,N_16666);
or U18947 (N_18947,N_16240,N_16957);
and U18948 (N_18948,N_18403,N_16831);
nand U18949 (N_18949,N_18477,N_17594);
and U18950 (N_18950,N_16728,N_17175);
nor U18951 (N_18951,N_17018,N_17104);
and U18952 (N_18952,N_16309,N_15787);
nand U18953 (N_18953,N_17576,N_16790);
nand U18954 (N_18954,N_17721,N_18077);
and U18955 (N_18955,N_18582,N_15693);
and U18956 (N_18956,N_18183,N_17094);
xnor U18957 (N_18957,N_18141,N_15828);
and U18958 (N_18958,N_18290,N_15708);
nor U18959 (N_18959,N_18078,N_18075);
nand U18960 (N_18960,N_17002,N_16350);
nand U18961 (N_18961,N_16158,N_15718);
or U18962 (N_18962,N_17687,N_15799);
or U18963 (N_18963,N_18531,N_17636);
xnor U18964 (N_18964,N_18087,N_15888);
nor U18965 (N_18965,N_17638,N_18719);
nand U18966 (N_18966,N_17567,N_17488);
or U18967 (N_18967,N_15998,N_18284);
nand U18968 (N_18968,N_18668,N_15674);
xor U18969 (N_18969,N_17541,N_18379);
and U18970 (N_18970,N_18226,N_18010);
xor U18971 (N_18971,N_16417,N_15967);
and U18972 (N_18972,N_16051,N_18532);
and U18973 (N_18973,N_15627,N_15773);
xor U18974 (N_18974,N_17581,N_16314);
nor U18975 (N_18975,N_15818,N_16704);
xnor U18976 (N_18976,N_17440,N_17478);
nor U18977 (N_18977,N_18543,N_15894);
and U18978 (N_18978,N_17494,N_18291);
nand U18979 (N_18979,N_17766,N_17498);
nor U18980 (N_18980,N_17268,N_16887);
nand U18981 (N_18981,N_16903,N_18385);
nor U18982 (N_18982,N_17730,N_16308);
or U18983 (N_18983,N_17239,N_16011);
nor U18984 (N_18984,N_17570,N_18508);
or U18985 (N_18985,N_18329,N_16726);
and U18986 (N_18986,N_17479,N_17454);
nor U18987 (N_18987,N_15995,N_16137);
and U18988 (N_18988,N_17514,N_16622);
nand U18989 (N_18989,N_17087,N_16284);
or U18990 (N_18990,N_16646,N_18595);
or U18991 (N_18991,N_18548,N_18196);
xnor U18992 (N_18992,N_15883,N_18637);
or U18993 (N_18993,N_18467,N_18414);
nand U18994 (N_18994,N_17366,N_17000);
nand U18995 (N_18995,N_18208,N_16370);
xnor U18996 (N_18996,N_17073,N_17156);
nand U18997 (N_18997,N_18216,N_18432);
and U18998 (N_18998,N_18529,N_16159);
or U18999 (N_18999,N_17611,N_15880);
or U19000 (N_19000,N_15690,N_15726);
nand U19001 (N_19001,N_16791,N_16649);
nand U19002 (N_19002,N_17548,N_17979);
nor U19003 (N_19003,N_17580,N_18113);
nand U19004 (N_19004,N_17853,N_17444);
xor U19005 (N_19005,N_18037,N_17465);
or U19006 (N_19006,N_16987,N_17771);
nand U19007 (N_19007,N_18317,N_18263);
and U19008 (N_19008,N_15909,N_16730);
nor U19009 (N_19009,N_17212,N_15873);
or U19010 (N_19010,N_16560,N_17859);
nand U19011 (N_19011,N_17222,N_16297);
and U19012 (N_19012,N_16776,N_18608);
and U19013 (N_19013,N_15750,N_17810);
or U19014 (N_19014,N_16813,N_17802);
or U19015 (N_19015,N_17939,N_16249);
nor U19016 (N_19016,N_17098,N_16246);
xnor U19017 (N_19017,N_16289,N_16466);
nand U19018 (N_19018,N_16252,N_16805);
xor U19019 (N_19019,N_15851,N_18642);
and U19020 (N_19020,N_17463,N_17786);
or U19021 (N_19021,N_17860,N_18635);
or U19022 (N_19022,N_17805,N_17032);
xnor U19023 (N_19023,N_17302,N_16168);
and U19024 (N_19024,N_18542,N_16010);
or U19025 (N_19025,N_17902,N_16060);
nor U19026 (N_19026,N_17065,N_18093);
nand U19027 (N_19027,N_16617,N_18541);
and U19028 (N_19028,N_18515,N_15970);
and U19029 (N_19029,N_16714,N_18649);
xnor U19030 (N_19030,N_16625,N_17339);
nor U19031 (N_19031,N_16440,N_17486);
xor U19032 (N_19032,N_17031,N_16584);
and U19033 (N_19033,N_18738,N_18578);
or U19034 (N_19034,N_17101,N_16823);
nor U19035 (N_19035,N_16651,N_17772);
and U19036 (N_19036,N_16458,N_17353);
or U19037 (N_19037,N_15810,N_17005);
or U19038 (N_19038,N_17868,N_17540);
or U19039 (N_19039,N_16605,N_15762);
and U19040 (N_19040,N_16331,N_16220);
and U19041 (N_19041,N_15921,N_16253);
nor U19042 (N_19042,N_16050,N_16196);
nor U19043 (N_19043,N_17496,N_17674);
nand U19044 (N_19044,N_16541,N_17030);
and U19045 (N_19045,N_18651,N_18220);
nand U19046 (N_19046,N_17574,N_16942);
nand U19047 (N_19047,N_16842,N_17847);
or U19048 (N_19048,N_16225,N_17705);
xor U19049 (N_19049,N_15981,N_15699);
xor U19050 (N_19050,N_15973,N_16442);
or U19051 (N_19051,N_16994,N_16407);
nor U19052 (N_19052,N_18563,N_18128);
and U19053 (N_19053,N_18436,N_17282);
nand U19054 (N_19054,N_17368,N_17241);
and U19055 (N_19055,N_18092,N_16109);
or U19056 (N_19056,N_16226,N_17832);
and U19057 (N_19057,N_18343,N_17343);
nand U19058 (N_19058,N_17198,N_17260);
and U19059 (N_19059,N_16326,N_15676);
xor U19060 (N_19060,N_17655,N_17303);
nor U19061 (N_19061,N_16279,N_16457);
or U19062 (N_19062,N_18131,N_17937);
and U19063 (N_19063,N_17147,N_17948);
and U19064 (N_19064,N_16975,N_18391);
or U19065 (N_19065,N_17664,N_16983);
nor U19066 (N_19066,N_16337,N_17127);
nand U19067 (N_19067,N_17228,N_17673);
nand U19068 (N_19068,N_18145,N_16593);
and U19069 (N_19069,N_18581,N_15653);
and U19070 (N_19070,N_16555,N_17745);
xor U19071 (N_19071,N_18181,N_15796);
xnor U19072 (N_19072,N_18285,N_15987);
and U19073 (N_19073,N_17255,N_18020);
nand U19074 (N_19074,N_16475,N_16868);
or U19075 (N_19075,N_17740,N_18460);
nor U19076 (N_19076,N_16968,N_15710);
and U19077 (N_19077,N_17102,N_16960);
xnor U19078 (N_19078,N_17110,N_17729);
nor U19079 (N_19079,N_17735,N_18034);
nand U19080 (N_19080,N_17931,N_16501);
and U19081 (N_19081,N_16369,N_18629);
xnor U19082 (N_19082,N_16321,N_16477);
nand U19083 (N_19083,N_16964,N_18232);
nand U19084 (N_19084,N_17562,N_15671);
xor U19085 (N_19085,N_16946,N_17186);
or U19086 (N_19086,N_16134,N_17409);
and U19087 (N_19087,N_18188,N_18341);
nor U19088 (N_19088,N_16432,N_15820);
nor U19089 (N_19089,N_16491,N_16312);
nand U19090 (N_19090,N_16311,N_17099);
or U19091 (N_19091,N_17043,N_17320);
nor U19092 (N_19092,N_17682,N_18154);
nor U19093 (N_19093,N_16398,N_17899);
nor U19094 (N_19094,N_17188,N_17297);
nor U19095 (N_19095,N_17448,N_17858);
xnor U19096 (N_19096,N_16828,N_16275);
nand U19097 (N_19097,N_16344,N_17820);
xor U19098 (N_19098,N_18580,N_18144);
nor U19099 (N_19099,N_18355,N_15980);
and U19100 (N_19100,N_16085,N_17380);
xor U19101 (N_19101,N_18321,N_15640);
nor U19102 (N_19102,N_17628,N_17063);
nor U19103 (N_19103,N_17192,N_18146);
nor U19104 (N_19104,N_18260,N_16610);
or U19105 (N_19105,N_17685,N_18206);
or U19106 (N_19106,N_16514,N_16446);
nand U19107 (N_19107,N_17051,N_15947);
or U19108 (N_19108,N_16986,N_17408);
nor U19109 (N_19109,N_16423,N_15985);
xor U19110 (N_19110,N_16413,N_17784);
nand U19111 (N_19111,N_18297,N_18514);
xor U19112 (N_19112,N_17141,N_18716);
xnor U19113 (N_19113,N_16147,N_18168);
or U19114 (N_19114,N_18709,N_17848);
xnor U19115 (N_19115,N_16580,N_16465);
nor U19116 (N_19116,N_17430,N_15768);
nand U19117 (N_19117,N_17259,N_17645);
xor U19118 (N_19118,N_16782,N_17139);
nand U19119 (N_19119,N_17836,N_18559);
and U19120 (N_19120,N_18522,N_17575);
or U19121 (N_19121,N_17584,N_17160);
nand U19122 (N_19122,N_18241,N_17341);
and U19123 (N_19123,N_16016,N_18691);
xnor U19124 (N_19124,N_16689,N_16306);
nor U19125 (N_19125,N_17340,N_16015);
nor U19126 (N_19126,N_16402,N_16811);
and U19127 (N_19127,N_16161,N_16211);
xnor U19128 (N_19128,N_16947,N_17790);
nand U19129 (N_19129,N_17138,N_17846);
nor U19130 (N_19130,N_15959,N_16106);
xor U19131 (N_19131,N_18513,N_17922);
or U19132 (N_19132,N_16366,N_17377);
or U19133 (N_19133,N_16703,N_16497);
nor U19134 (N_19134,N_16179,N_18111);
nor U19135 (N_19135,N_17975,N_16456);
nand U19136 (N_19136,N_18717,N_16521);
or U19137 (N_19137,N_17437,N_16634);
or U19138 (N_19138,N_17924,N_17106);
or U19139 (N_19139,N_18407,N_16207);
nand U19140 (N_19140,N_17511,N_16323);
or U19141 (N_19141,N_17028,N_16909);
xor U19142 (N_19142,N_16683,N_17202);
and U19143 (N_19143,N_16827,N_18102);
and U19144 (N_19144,N_15872,N_18695);
or U19145 (N_19145,N_16722,N_16489);
and U19146 (N_19146,N_17417,N_15629);
nand U19147 (N_19147,N_15938,N_16872);
nand U19148 (N_19148,N_16712,N_17253);
xor U19149 (N_19149,N_18229,N_15825);
and U19150 (N_19150,N_18370,N_17396);
nand U19151 (N_19151,N_16139,N_18692);
nand U19152 (N_19152,N_16812,N_17968);
and U19153 (N_19153,N_16241,N_18239);
nor U19154 (N_19154,N_17042,N_18104);
nand U19155 (N_19155,N_16049,N_17484);
nor U19156 (N_19156,N_16527,N_17811);
or U19157 (N_19157,N_17130,N_17323);
or U19158 (N_19158,N_17669,N_16858);
and U19159 (N_19159,N_16169,N_15645);
xor U19160 (N_19160,N_17719,N_16669);
and U19161 (N_19161,N_18198,N_15968);
nor U19162 (N_19162,N_15857,N_16119);
and U19163 (N_19163,N_16318,N_17203);
nand U19164 (N_19164,N_17829,N_16193);
xor U19165 (N_19165,N_18498,N_16079);
and U19166 (N_19166,N_16322,N_15650);
nor U19167 (N_19167,N_16911,N_16406);
xnor U19168 (N_19168,N_17447,N_15723);
and U19169 (N_19169,N_18358,N_18412);
nand U19170 (N_19170,N_16864,N_15950);
nor U19171 (N_19171,N_16221,N_15827);
nand U19172 (N_19172,N_16065,N_17512);
xnor U19173 (N_19173,N_17185,N_17289);
or U19174 (N_19174,N_16719,N_18476);
or U19175 (N_19175,N_18177,N_17967);
xnor U19176 (N_19176,N_16639,N_17034);
or U19177 (N_19177,N_18545,N_17617);
or U19178 (N_19178,N_18618,N_16624);
nor U19179 (N_19179,N_17331,N_18032);
nor U19180 (N_19180,N_18174,N_18624);
and U19181 (N_19181,N_16447,N_17972);
xnor U19182 (N_19182,N_18074,N_16469);
and U19183 (N_19183,N_16405,N_16877);
xor U19184 (N_19184,N_18666,N_17219);
xnor U19185 (N_19185,N_17516,N_17257);
xnor U19186 (N_19186,N_16014,N_17727);
and U19187 (N_19187,N_17634,N_16727);
or U19188 (N_19188,N_18499,N_18318);
nand U19189 (N_19189,N_17677,N_17696);
or U19190 (N_19190,N_16638,N_16755);
xnor U19191 (N_19191,N_17429,N_17928);
nor U19192 (N_19192,N_17986,N_16507);
nand U19193 (N_19193,N_17871,N_16394);
nor U19194 (N_19194,N_17606,N_18053);
and U19195 (N_19195,N_15891,N_17128);
nand U19196 (N_19196,N_18003,N_16515);
nor U19197 (N_19197,N_17549,N_18148);
and U19198 (N_19198,N_16058,N_16913);
nand U19199 (N_19199,N_17560,N_18007);
and U19200 (N_19200,N_18597,N_18413);
or U19201 (N_19201,N_16063,N_16230);
xnor U19202 (N_19202,N_17061,N_18024);
nor U19203 (N_19203,N_17622,N_17356);
nand U19204 (N_19204,N_16575,N_16800);
nand U19205 (N_19205,N_17345,N_18107);
xor U19206 (N_19206,N_17849,N_17361);
or U19207 (N_19207,N_17062,N_16594);
xor U19208 (N_19208,N_16005,N_16068);
nor U19209 (N_19209,N_17839,N_16547);
xnor U19210 (N_19210,N_16820,N_17084);
or U19211 (N_19211,N_17508,N_18085);
or U19212 (N_19212,N_17553,N_18367);
nand U19213 (N_19213,N_18424,N_15886);
nor U19214 (N_19214,N_18702,N_17369);
xor U19215 (N_19215,N_15941,N_15709);
xor U19216 (N_19216,N_18365,N_17504);
and U19217 (N_19217,N_18361,N_17249);
or U19218 (N_19218,N_16908,N_16219);
and U19219 (N_19219,N_18549,N_16787);
or U19220 (N_19220,N_17671,N_15929);
nand U19221 (N_19221,N_16444,N_18536);
nand U19222 (N_19222,N_17391,N_17025);
nand U19223 (N_19223,N_17363,N_16565);
nand U19224 (N_19224,N_16821,N_17495);
nor U19225 (N_19225,N_16243,N_17420);
or U19226 (N_19226,N_17845,N_18564);
and U19227 (N_19227,N_17813,N_17451);
nor U19228 (N_19228,N_16094,N_16191);
and U19229 (N_19229,N_17995,N_17962);
xor U19230 (N_19230,N_18002,N_17883);
nor U19231 (N_19231,N_16628,N_17887);
and U19232 (N_19232,N_18247,N_17011);
or U19233 (N_19233,N_17640,N_15808);
nor U19234 (N_19234,N_18492,N_17925);
and U19235 (N_19235,N_16443,N_17350);
nor U19236 (N_19236,N_17754,N_16329);
nor U19237 (N_19237,N_15784,N_16290);
and U19238 (N_19238,N_17411,N_17489);
and U19239 (N_19239,N_18011,N_17886);
and U19240 (N_19240,N_16053,N_15956);
or U19241 (N_19241,N_16779,N_17637);
nor U19242 (N_19242,N_15884,N_17563);
nand U19243 (N_19243,N_17415,N_17233);
nand U19244 (N_19244,N_18236,N_17068);
and U19245 (N_19245,N_17012,N_18546);
and U19246 (N_19246,N_16837,N_16162);
nor U19247 (N_19247,N_15882,N_16801);
and U19248 (N_19248,N_17382,N_15651);
nor U19249 (N_19249,N_16461,N_17372);
and U19250 (N_19250,N_16901,N_16237);
or U19251 (N_19251,N_16182,N_18446);
and U19252 (N_19252,N_15830,N_16799);
or U19253 (N_19253,N_17756,N_17878);
xor U19254 (N_19254,N_18013,N_18132);
or U19255 (N_19255,N_15996,N_18305);
or U19256 (N_19256,N_16550,N_16347);
nand U19257 (N_19257,N_15905,N_18315);
nor U19258 (N_19258,N_17976,N_18579);
and U19259 (N_19259,N_17083,N_15901);
nor U19260 (N_19260,N_16335,N_17443);
nand U19261 (N_19261,N_15746,N_17787);
xor U19262 (N_19262,N_18415,N_18661);
nor U19263 (N_19263,N_16615,N_17539);
xnor U19264 (N_19264,N_17322,N_18056);
or U19265 (N_19265,N_18221,N_16086);
xor U19266 (N_19266,N_17091,N_18440);
nand U19267 (N_19267,N_17718,N_17220);
nor U19268 (N_19268,N_17195,N_16133);
nor U19269 (N_19269,N_15926,N_16520);
xnor U19270 (N_19270,N_17610,N_18503);
nand U19271 (N_19271,N_18334,N_17402);
nand U19272 (N_19272,N_15896,N_15841);
and U19273 (N_19273,N_16476,N_17874);
and U19274 (N_19274,N_16117,N_16200);
nand U19275 (N_19275,N_16740,N_16426);
nor U19276 (N_19276,N_17501,N_15625);
xnor U19277 (N_19277,N_18491,N_17993);
and U19278 (N_19278,N_18377,N_18680);
or U19279 (N_19279,N_18098,N_16484);
nand U19280 (N_19280,N_17704,N_17621);
nor U19281 (N_19281,N_17639,N_18544);
xor U19282 (N_19282,N_16234,N_16709);
or U19283 (N_19283,N_18422,N_17658);
xor U19284 (N_19284,N_16166,N_17263);
xor U19285 (N_19285,N_17135,N_17421);
xnor U19286 (N_19286,N_16130,N_17133);
or U19287 (N_19287,N_18480,N_18004);
or U19288 (N_19288,N_17568,N_18557);
or U19289 (N_19289,N_18455,N_17572);
nand U19290 (N_19290,N_15636,N_17211);
xnor U19291 (N_19291,N_17779,N_16251);
nand U19292 (N_19292,N_17434,N_16789);
or U19293 (N_19293,N_17555,N_17881);
or U19294 (N_19294,N_17422,N_16340);
or U19295 (N_19295,N_16940,N_18119);
nor U19296 (N_19296,N_15892,N_17863);
xor U19297 (N_19297,N_17822,N_18703);
nand U19298 (N_19298,N_17056,N_16483);
xor U19299 (N_19299,N_15879,N_17374);
nor U19300 (N_19300,N_18383,N_15798);
nor U19301 (N_19301,N_17112,N_18138);
or U19302 (N_19302,N_17399,N_18309);
nand U19303 (N_19303,N_18584,N_17759);
nor U19304 (N_19304,N_17557,N_18621);
nor U19305 (N_19305,N_16008,N_18534);
xnor U19306 (N_19306,N_16295,N_16736);
xnor U19307 (N_19307,N_18014,N_17373);
nand U19308 (N_19308,N_18524,N_17393);
or U19309 (N_19309,N_18551,N_18484);
nor U19310 (N_19310,N_17903,N_17193);
nand U19311 (N_19311,N_15635,N_18046);
or U19312 (N_19312,N_15737,N_16202);
or U19313 (N_19313,N_16351,N_17129);
nor U19314 (N_19314,N_16454,N_18550);
and U19315 (N_19315,N_17294,N_18069);
or U19316 (N_19316,N_17251,N_16765);
or U19317 (N_19317,N_16338,N_17001);
or U19318 (N_19318,N_17276,N_16796);
or U19319 (N_19319,N_15953,N_18475);
xnor U19320 (N_19320,N_16250,N_18539);
nor U19321 (N_19321,N_16627,N_18294);
or U19322 (N_19322,N_16259,N_18662);
xnor U19323 (N_19323,N_17537,N_16320);
nor U19324 (N_19324,N_16601,N_16378);
nor U19325 (N_19325,N_16355,N_15815);
nand U19326 (N_19326,N_16990,N_16804);
and U19327 (N_19327,N_16563,N_15948);
and U19328 (N_19328,N_15795,N_18675);
nor U19329 (N_19329,N_17137,N_18160);
nand U19330 (N_19330,N_18091,N_17698);
nand U19331 (N_19331,N_18171,N_18275);
and U19332 (N_19332,N_17590,N_16317);
nand U19333 (N_19333,N_16995,N_17760);
or U19334 (N_19334,N_16391,N_18147);
and U19335 (N_19335,N_16834,N_16600);
and U19336 (N_19336,N_16346,N_17877);
or U19337 (N_19337,N_18478,N_16753);
and U19338 (N_19338,N_18096,N_16067);
or U19339 (N_19339,N_17908,N_17596);
or U19340 (N_19340,N_17602,N_18454);
nand U19341 (N_19341,N_18270,N_17414);
nand U19342 (N_19342,N_16265,N_17546);
nor U19343 (N_19343,N_18646,N_17485);
and U19344 (N_19344,N_17554,N_16976);
and U19345 (N_19345,N_17388,N_15794);
nand U19346 (N_19346,N_17279,N_18351);
xor U19347 (N_19347,N_18663,N_16697);
or U19348 (N_19348,N_16348,N_17985);
and U19349 (N_19349,N_16436,N_16184);
and U19350 (N_19350,N_15703,N_18325);
and U19351 (N_19351,N_15801,N_18601);
or U19352 (N_19352,N_17755,N_17123);
nor U19353 (N_19353,N_17809,N_17295);
nor U19354 (N_19354,N_16569,N_17301);
nand U19355 (N_19355,N_17788,N_15706);
and U19356 (N_19356,N_15655,N_18462);
xnor U19357 (N_19357,N_16523,N_16997);
nand U19358 (N_19358,N_18117,N_16939);
and U19359 (N_19359,N_16962,N_17768);
and U19360 (N_19360,N_17830,N_16183);
or U19361 (N_19361,N_16116,N_17970);
nor U19362 (N_19362,N_15780,N_17315);
or U19363 (N_19363,N_18708,N_15786);
nor U19364 (N_19364,N_17933,N_17288);
nand U19365 (N_19365,N_18479,N_15823);
and U19366 (N_19366,N_15881,N_18346);
or U19367 (N_19367,N_16125,N_17534);
or U19368 (N_19368,N_16871,N_17375);
or U19369 (N_19369,N_17632,N_15793);
xor U19370 (N_19370,N_16111,N_17806);
nor U19371 (N_19371,N_16090,N_16228);
or U19372 (N_19372,N_17605,N_18307);
nand U19373 (N_19373,N_16756,N_16926);
nor U19374 (N_19374,N_18185,N_16970);
nor U19375 (N_19375,N_17884,N_16349);
nor U19376 (N_19376,N_16747,N_17262);
and U19377 (N_19377,N_17900,N_16144);
or U19378 (N_19378,N_16187,N_16705);
and U19379 (N_19379,N_17204,N_16441);
nor U19380 (N_19380,N_16345,N_18213);
xnor U19381 (N_19381,N_15955,N_17524);
nor U19382 (N_19382,N_16764,N_18140);
or U19383 (N_19383,N_16694,N_16620);
nor U19384 (N_19384,N_17953,N_15667);
xnor U19385 (N_19385,N_16718,N_18337);
or U19386 (N_19386,N_18288,N_16591);
nand U19387 (N_19387,N_17826,N_15763);
or U19388 (N_19388,N_18310,N_17338);
and U19389 (N_19389,N_17081,N_17412);
xor U19390 (N_19390,N_17153,N_16822);
nor U19391 (N_19391,N_16735,N_16160);
xor U19392 (N_19392,N_18197,N_18569);
and U19393 (N_19393,N_18537,N_16368);
or U19394 (N_19394,N_18293,N_17039);
nand U19395 (N_19395,N_17551,N_17875);
xor U19396 (N_19396,N_16672,N_16809);
nand U19397 (N_19397,N_15748,N_16892);
nor U19398 (N_19398,N_16247,N_18699);
nand U19399 (N_19399,N_16922,N_18272);
xnor U19400 (N_19400,N_16676,N_18231);
nor U19401 (N_19401,N_17072,N_16216);
nand U19402 (N_19402,N_18605,N_15864);
nor U19403 (N_19403,N_16886,N_17152);
xor U19404 (N_19404,N_17381,N_16288);
or U19405 (N_19405,N_16953,N_17616);
xnor U19406 (N_19406,N_15865,N_17386);
and U19407 (N_19407,N_16112,N_16682);
nand U19408 (N_19408,N_16690,N_17773);
nor U19409 (N_19409,N_16100,N_17114);
or U19410 (N_19410,N_18079,N_16472);
or U19411 (N_19411,N_16132,N_17644);
or U19412 (N_19412,N_16332,N_18261);
xnor U19413 (N_19413,N_18129,N_16948);
and U19414 (N_19414,N_15849,N_17016);
nor U19415 (N_19415,N_17267,N_17467);
and U19416 (N_19416,N_17419,N_18049);
xnor U19417 (N_19417,N_17515,N_17633);
and U19418 (N_19418,N_15962,N_16425);
nor U19419 (N_19419,N_18114,N_17711);
nor U19420 (N_19420,N_18588,N_15720);
nand U19421 (N_19421,N_17082,N_16486);
or U19422 (N_19422,N_16841,N_18212);
nand U19423 (N_19423,N_18039,N_15889);
nor U19424 (N_19424,N_17446,N_18324);
or U19425 (N_19425,N_15663,N_17395);
nand U19426 (N_19426,N_18704,N_16896);
nor U19427 (N_19427,N_17428,N_16151);
xnor U19428 (N_19428,N_16026,N_16612);
nor U19429 (N_19429,N_16029,N_16245);
nor U19430 (N_19430,N_18535,N_15869);
or U19431 (N_19431,N_16741,N_17270);
xor U19432 (N_19432,N_18218,N_18576);
and U19433 (N_19433,N_15744,N_15918);
nand U19434 (N_19434,N_16316,N_15742);
nor U19435 (N_19435,N_18448,N_18095);
xor U19436 (N_19436,N_17182,N_18256);
xnor U19437 (N_19437,N_17035,N_17425);
xnor U19438 (N_19438,N_17799,N_16101);
nor U19439 (N_19439,N_17181,N_17392);
nor U19440 (N_19440,N_18723,N_17441);
or U19441 (N_19441,N_17245,N_18109);
nand U19442 (N_19442,N_18511,N_15711);
xnor U19443 (N_19443,N_17014,N_16938);
or U19444 (N_19444,N_17808,N_15797);
or U19445 (N_19445,N_18726,N_16924);
or U19446 (N_19446,N_17095,N_17612);
nor U19447 (N_19447,N_16596,N_15678);
nand U19448 (N_19448,N_17743,N_18433);
nor U19449 (N_19449,N_17460,N_17124);
or U19450 (N_19450,N_17661,N_15809);
xor U19451 (N_19451,N_17747,N_17466);
xnor U19452 (N_19452,N_17601,N_17248);
nand U19453 (N_19453,N_16971,N_17418);
and U19454 (N_19454,N_17458,N_16751);
and U19455 (N_19455,N_16588,N_17321);
nor U19456 (N_19456,N_17013,N_18488);
nor U19457 (N_19457,N_17701,N_18064);
xor U19458 (N_19458,N_16793,N_16870);
or U19459 (N_19459,N_16463,N_17319);
nor U19460 (N_19460,N_17991,N_17600);
nor U19461 (N_19461,N_17794,N_17142);
and U19462 (N_19462,N_16266,N_18344);
or U19463 (N_19463,N_17161,N_18610);
and U19464 (N_19464,N_15940,N_15854);
xor U19465 (N_19465,N_17397,N_18057);
and U19466 (N_19466,N_15694,N_18644);
nor U19467 (N_19467,N_18684,N_15819);
and U19468 (N_19468,N_16899,N_17483);
and U19469 (N_19469,N_18159,N_16036);
or U19470 (N_19470,N_18526,N_16817);
or U19471 (N_19471,N_17311,N_15764);
and U19472 (N_19472,N_15945,N_18647);
xor U19473 (N_19473,N_18328,N_16342);
nand U19474 (N_19474,N_16084,N_18561);
nand U19475 (N_19475,N_16963,N_15713);
or U19476 (N_19476,N_16271,N_16076);
nor U19477 (N_19477,N_15965,N_18269);
nand U19478 (N_19478,N_17974,N_16255);
nor U19479 (N_19479,N_17905,N_18749);
nor U19480 (N_19480,N_18727,N_17404);
xor U19481 (N_19481,N_16356,N_15783);
or U19482 (N_19482,N_16509,N_18530);
xor U19483 (N_19483,N_16142,N_17700);
or U19484 (N_19484,N_17020,N_18097);
nand U19485 (N_19485,N_18063,N_17579);
nand U19486 (N_19486,N_16732,N_16954);
nand U19487 (N_19487,N_16688,N_17694);
xnor U19488 (N_19488,N_16586,N_17798);
nand U19489 (N_19489,N_17789,N_15890);
xnor U19490 (N_19490,N_15897,N_16467);
or U19491 (N_19491,N_17385,N_16904);
nor U19492 (N_19492,N_15776,N_16263);
xnor U19493 (N_19493,N_16848,N_16613);
xnor U19494 (N_19494,N_17545,N_16830);
xnor U19495 (N_19495,N_16597,N_16587);
nor U19496 (N_19496,N_16260,N_16126);
xnor U19497 (N_19497,N_18435,N_16028);
or U19498 (N_19498,N_16936,N_16287);
nand U19499 (N_19499,N_17566,N_17722);
nor U19500 (N_19500,N_16267,N_17281);
or U19501 (N_19501,N_16209,N_17961);
nand U19502 (N_19502,N_18506,N_16898);
and U19503 (N_19503,N_16399,N_16571);
nor U19504 (N_19504,N_16227,N_16763);
nand U19505 (N_19505,N_18360,N_15684);
nand U19506 (N_19506,N_16385,N_16533);
nand U19507 (N_19507,N_16429,N_16498);
and U19508 (N_19508,N_18570,N_18258);
xnor U19509 (N_19509,N_18210,N_18045);
xor U19510 (N_19510,N_16066,N_16389);
nor U19511 (N_19511,N_16879,N_17869);
or U19512 (N_19512,N_18195,N_18133);
or U19513 (N_19513,N_17214,N_15990);
xnor U19514 (N_19514,N_18112,N_17732);
nand U19515 (N_19515,N_15805,N_17892);
nor U19516 (N_19516,N_15691,N_18746);
or U19517 (N_19517,N_17261,N_17984);
nor U19518 (N_19518,N_16414,N_17629);
and U19519 (N_19519,N_18266,N_16771);
or U19520 (N_19520,N_16641,N_16212);
or U19521 (N_19521,N_18178,N_18035);
nand U19522 (N_19522,N_17641,N_17044);
and U19523 (N_19523,N_15774,N_18068);
nand U19524 (N_19524,N_17221,N_17707);
nor U19525 (N_19525,N_15685,N_18554);
and U19526 (N_19526,N_18725,N_16582);
or U19527 (N_19527,N_17692,N_16528);
nor U19528 (N_19528,N_16846,N_16301);
xnor U19529 (N_19529,N_18469,N_16687);
nor U19530 (N_19530,N_18161,N_16934);
nand U19531 (N_19531,N_16900,N_17603);
nor U19532 (N_19532,N_15944,N_16170);
nand U19533 (N_19533,N_17119,N_16192);
nor U19534 (N_19534,N_16257,N_15837);
and U19535 (N_19535,N_16656,N_17529);
xnor U19536 (N_19536,N_16403,N_18224);
nand U19537 (N_19537,N_16093,N_16072);
and U19538 (N_19538,N_17365,N_17046);
or U19539 (N_19539,N_17472,N_17507);
and U19540 (N_19540,N_17089,N_16108);
or U19541 (N_19541,N_16032,N_16131);
or U19542 (N_19542,N_15734,N_16673);
xnor U19543 (N_19543,N_17912,N_17803);
or U19544 (N_19544,N_18693,N_17136);
nor U19545 (N_19545,N_15875,N_16606);
nor U19546 (N_19546,N_16604,N_17017);
nor U19547 (N_19547,N_18573,N_16832);
nor U19548 (N_19548,N_16002,N_17047);
and U19549 (N_19549,N_17159,N_17750);
and U19550 (N_19550,N_17108,N_18611);
or U19551 (N_19551,N_17819,N_16254);
xor U19552 (N_19552,N_18225,N_16075);
or U19553 (N_19553,N_15725,N_17942);
xor U19554 (N_19554,N_16680,N_15847);
and U19555 (N_19555,N_18650,N_16630);
xor U19556 (N_19556,N_17342,N_16902);
nor U19557 (N_19557,N_17651,N_15683);
and U19558 (N_19558,N_16912,N_16829);
or U19559 (N_19559,N_16450,N_16153);
or U19560 (N_19560,N_18116,N_15871);
xnor U19561 (N_19561,N_17856,N_16427);
xor U19562 (N_19562,N_15856,N_16944);
and U19563 (N_19563,N_16043,N_16743);
nand U19564 (N_19564,N_15790,N_17532);
nand U19565 (N_19565,N_18222,N_18490);
nor U19566 (N_19566,N_18423,N_15919);
xor U19567 (N_19567,N_18655,N_16665);
nand U19568 (N_19568,N_15700,N_17543);
nor U19569 (N_19569,N_15984,N_16033);
xnor U19570 (N_19570,N_17864,N_16784);
nor U19571 (N_19571,N_16551,N_15668);
or U19572 (N_19572,N_16083,N_16478);
or U19573 (N_19573,N_15649,N_18029);
and U19574 (N_19574,N_15659,N_18670);
or U19575 (N_19575,N_16773,N_17963);
xnor U19576 (N_19576,N_17509,N_18354);
nand U19577 (N_19577,N_16071,N_18393);
nor U19578 (N_19578,N_17462,N_18262);
and U19579 (N_19579,N_17383,N_18384);
xor U19580 (N_19580,N_18033,N_16748);
nand U19581 (N_19581,N_16920,N_18201);
or U19582 (N_19582,N_15979,N_16611);
or U19583 (N_19583,N_15999,N_16115);
or U19584 (N_19584,N_18106,N_16141);
nor U19585 (N_19585,N_18447,N_18347);
nor U19586 (N_19586,N_16303,N_15782);
nand U19587 (N_19587,N_18058,N_17329);
xor U19588 (N_19588,N_16993,N_18071);
nand U19589 (N_19589,N_16717,N_16857);
and U19590 (N_19590,N_16163,N_15874);
nor U19591 (N_19591,N_18348,N_18641);
nor U19592 (N_19592,N_17619,N_18583);
xnor U19593 (N_19593,N_18464,N_17150);
and U19594 (N_19594,N_15749,N_17158);
nand U19595 (N_19595,N_17936,N_18124);
and U19596 (N_19596,N_15712,N_17526);
or U19597 (N_19597,N_17378,N_18690);
or U19598 (N_19598,N_16859,N_16269);
and U19599 (N_19599,N_16102,N_17558);
xnor U19600 (N_19600,N_17265,N_17954);
xor U19601 (N_19601,N_15852,N_18026);
xor U19602 (N_19602,N_17929,N_17196);
or U19603 (N_19603,N_17019,N_17589);
nand U19604 (N_19604,N_16933,N_16419);
nor U19605 (N_19605,N_17944,N_16664);
xor U19606 (N_19606,N_15887,N_16810);
nor U19607 (N_19607,N_17503,N_17697);
xnor U19608 (N_19608,N_16725,N_16453);
nand U19609 (N_19609,N_17075,N_17238);
nand U19610 (N_19610,N_17224,N_15687);
xnor U19611 (N_19611,N_18517,N_15804);
and U19612 (N_19612,N_17835,N_18240);
xnor U19613 (N_19613,N_18598,N_16781);
nand U19614 (N_19614,N_16866,N_18070);
or U19615 (N_19615,N_16969,N_15803);
or U19616 (N_19616,N_17800,N_16803);
nor U19617 (N_19617,N_17996,N_18207);
nand U19618 (N_19618,N_16972,N_17317);
and U19619 (N_19619,N_16745,N_17183);
and U19620 (N_19620,N_18638,N_18214);
nor U19621 (N_19621,N_16300,N_18048);
xor U19622 (N_19622,N_16999,N_16175);
nor U19623 (N_19623,N_18000,N_15751);
nand U19624 (N_19624,N_15766,N_18060);
and U19625 (N_19625,N_16910,N_15925);
nor U19626 (N_19626,N_18566,N_18265);
or U19627 (N_19627,N_17066,N_17036);
nand U19628 (N_19628,N_16437,N_16642);
or U19629 (N_19629,N_16188,N_17988);
nor U19630 (N_19630,N_15631,N_18308);
or U19631 (N_19631,N_18568,N_17982);
nand U19632 (N_19632,N_16785,N_16814);
nor U19633 (N_19633,N_18055,N_18125);
and U19634 (N_19634,N_17456,N_17708);
and U19635 (N_19635,N_15648,N_17680);
and U19636 (N_19636,N_17855,N_18639);
nand U19637 (N_19637,N_16171,N_15978);
and U19638 (N_19638,N_16686,N_18606);
xnor U19639 (N_19639,N_17499,N_17726);
nor U19640 (N_19640,N_17155,N_18615);
nand U19641 (N_19641,N_16616,N_17189);
nor U19642 (N_19642,N_16401,N_17957);
and U19643 (N_19643,N_16526,N_16549);
or U19644 (N_19644,N_16699,N_18459);
and U19645 (N_19645,N_16487,N_17355);
or U19646 (N_19646,N_17926,N_18243);
nor U19647 (N_19647,N_15666,N_17876);
xnor U19648 (N_19648,N_15932,N_16775);
nor U19649 (N_19649,N_15769,N_17432);
xor U19650 (N_19650,N_18734,N_18122);
or U19651 (N_19651,N_17891,N_18356);
or U19652 (N_19652,N_15760,N_16873);
or U19653 (N_19653,N_17844,N_18298);
or U19654 (N_19654,N_15647,N_18398);
xnor U19655 (N_19655,N_16648,N_18281);
or U19656 (N_19656,N_18100,N_16923);
and U19657 (N_19657,N_17866,N_18313);
and U19658 (N_19658,N_16798,N_16353);
xor U19659 (N_19659,N_16354,N_17893);
nor U19660 (N_19660,N_15752,N_17824);
xnor U19661 (N_19661,N_17604,N_15800);
xnor U19662 (N_19662,N_16154,N_18722);
xnor U19663 (N_19663,N_17250,N_17840);
and U19664 (N_19664,N_16715,N_17780);
nand U19665 (N_19665,N_17078,N_16488);
xnor U19666 (N_19666,N_17197,N_16120);
or U19667 (N_19667,N_18729,N_16430);
xnor U19668 (N_19668,N_16124,N_17583);
or U19669 (N_19669,N_16021,N_17690);
and U19670 (N_19670,N_17439,N_17149);
nor U19671 (N_19671,N_18523,N_17271);
and U19672 (N_19672,N_17405,N_15840);
nor U19673 (N_19673,N_17459,N_18560);
or U19674 (N_19674,N_18714,N_16118);
nand U19675 (N_19675,N_18211,N_15963);
nor U19676 (N_19676,N_15972,N_17243);
and U19677 (N_19677,N_16302,N_16529);
or U19678 (N_19678,N_18250,N_16500);
and U19679 (N_19679,N_16833,N_16490);
nor U19680 (N_19680,N_15675,N_15983);
nand U19681 (N_19681,N_16382,N_16198);
and U19682 (N_19682,N_16359,N_17791);
nand U19683 (N_19683,N_16978,N_16552);
nand U19684 (N_19684,N_16698,N_17870);
xnor U19685 (N_19685,N_16328,N_16906);
nor U19686 (N_19686,N_18364,N_15698);
nor U19687 (N_19687,N_17045,N_18350);
or U19688 (N_19688,N_18507,N_16777);
nand U19689 (N_19689,N_17825,N_18217);
or U19690 (N_19690,N_16422,N_16860);
nor U19691 (N_19691,N_17607,N_16959);
nor U19692 (N_19692,N_16232,N_16738);
nand U19693 (N_19693,N_16493,N_16270);
nor U19694 (N_19694,N_18162,N_16965);
and U19695 (N_19695,N_17215,N_17178);
and U19696 (N_19696,N_18121,N_15677);
or U19697 (N_19697,N_16576,N_17096);
or U19698 (N_19698,N_16248,N_17246);
nor U19699 (N_19699,N_16428,N_16242);
and U19700 (N_19700,N_18538,N_17307);
or U19701 (N_19701,N_18103,N_17728);
nand U19702 (N_19702,N_18374,N_17695);
and U19703 (N_19703,N_17205,N_17278);
or U19704 (N_19704,N_17477,N_17646);
or U19705 (N_19705,N_16590,N_16652);
and U19706 (N_19706,N_15662,N_17333);
nand U19707 (N_19707,N_18182,N_15721);
xor U19708 (N_19708,N_17843,N_17561);
nand U19709 (N_19709,N_16840,N_17304);
and U19710 (N_19710,N_18623,N_17679);
nor U19711 (N_19711,N_18289,N_16937);
nor U19712 (N_19712,N_17592,N_16708);
xor U19713 (N_19713,N_15923,N_16626);
nand U19714 (N_19714,N_17076,N_16409);
or U19715 (N_19715,N_16485,N_16921);
nand U19716 (N_19716,N_16540,N_16371);
and U19717 (N_19717,N_15632,N_17476);
or U19718 (N_19718,N_18246,N_17872);
nand U19719 (N_19719,N_16387,N_18631);
nor U19720 (N_19720,N_18494,N_16742);
or U19721 (N_19721,N_16434,N_16589);
nand U19722 (N_19722,N_16199,N_16283);
nor U19723 (N_19723,N_18710,N_16928);
xnor U19724 (N_19724,N_18237,N_16974);
and U19725 (N_19725,N_15898,N_17435);
and U19726 (N_19726,N_18489,N_17693);
or U19727 (N_19727,N_17284,N_15866);
nor U19728 (N_19728,N_15824,N_16768);
nand U19729 (N_19729,N_17706,N_17370);
or U19730 (N_19730,N_18042,N_17519);
nand U19731 (N_19731,N_15943,N_17318);
nor U19732 (N_19732,N_16468,N_17724);
nor U19733 (N_19733,N_17423,N_18574);
and U19734 (N_19734,N_17111,N_18006);
and U19735 (N_19735,N_18043,N_15761);
xnor U19736 (N_19736,N_18301,N_17208);
nor U19737 (N_19737,N_16138,N_17746);
xor U19738 (N_19738,N_16089,N_16679);
and U19739 (N_19739,N_17989,N_16206);
nor U19740 (N_19740,N_18362,N_18153);
or U19741 (N_19741,N_17880,N_16258);
xor U19742 (N_19742,N_18101,N_17349);
and U19743 (N_19743,N_15772,N_18038);
and U19744 (N_19744,N_18626,N_16696);
nor U19745 (N_19745,N_15900,N_18322);
xor U19746 (N_19746,N_16778,N_17978);
xnor U19747 (N_19747,N_15775,N_18473);
nor U19748 (N_19748,N_18689,N_17120);
nor U19749 (N_19749,N_16967,N_16759);
nor U19750 (N_19750,N_16025,N_16327);
nand U19751 (N_19751,N_16985,N_16397);
nand U19752 (N_19752,N_17269,N_17293);
nand U19753 (N_19753,N_18399,N_16952);
or U19754 (N_19754,N_16189,N_15672);
nand U19755 (N_19755,N_18553,N_17151);
and U19756 (N_19756,N_18252,N_16460);
or U19757 (N_19757,N_16762,N_15966);
nor U19758 (N_19758,N_18081,N_16542);
xor U19759 (N_19759,N_15833,N_18155);
and U19760 (N_19760,N_16208,N_17525);
xnor U19761 (N_19761,N_17569,N_18015);
nand U19762 (N_19762,N_17334,N_18417);
or U19763 (N_19763,N_17527,N_18388);
xnor U19764 (N_19764,N_17834,N_18190);
or U19765 (N_19765,N_16019,N_18556);
xnor U19766 (N_19766,N_16505,N_16918);
nand U19767 (N_19767,N_17670,N_16754);
or U19768 (N_19768,N_17103,N_16165);
and U19769 (N_19769,N_18030,N_16156);
and U19770 (N_19770,N_16504,N_17132);
nor U19771 (N_19771,N_18203,N_15792);
or U19772 (N_19772,N_15628,N_18073);
nand U19773 (N_19773,N_15639,N_17070);
and U19774 (N_19774,N_15779,N_15777);
nor U19775 (N_19775,N_18302,N_16213);
nand U19776 (N_19776,N_18558,N_17681);
xor U19777 (N_19777,N_15643,N_16767);
xnor U19778 (N_19778,N_18139,N_16693);
xor U19779 (N_19779,N_16766,N_15863);
xor U19780 (N_19780,N_18683,N_16473);
xor U19781 (N_19781,N_16041,N_18430);
or U19782 (N_19782,N_15778,N_15707);
or U19783 (N_19783,N_17588,N_17218);
or U19784 (N_19784,N_17237,N_16022);
xor U19785 (N_19785,N_17983,N_17093);
nand U19786 (N_19786,N_16256,N_16499);
nor U19787 (N_19787,N_17236,N_18728);
and U19788 (N_19788,N_16018,N_16210);
and U19789 (N_19789,N_17157,N_18711);
or U19790 (N_19790,N_15903,N_16040);
and U19791 (N_19791,N_18521,N_17240);
nand U19792 (N_19792,N_17623,N_16819);
nor U19793 (N_19793,N_15867,N_17614);
xnor U19794 (N_19794,N_18331,N_15642);
nor U19795 (N_19795,N_15964,N_18279);
or U19796 (N_19796,N_17337,N_18592);
nor U19797 (N_19797,N_16061,N_17040);
and U19798 (N_19798,N_17782,N_18363);
nand U19799 (N_19799,N_16758,N_16007);
or U19800 (N_19800,N_16824,N_18429);
xnor U19801 (N_19801,N_17943,N_17457);
xnor U19802 (N_19802,N_18696,N_17668);
nor U19803 (N_19803,N_18357,N_17292);
or U19804 (N_19804,N_17354,N_16553);
or U19805 (N_19805,N_16178,N_17675);
xnor U19806 (N_19806,N_18352,N_18496);
xor U19807 (N_19807,N_16012,N_17765);
nor U19808 (N_19808,N_18105,N_15954);
nor U19809 (N_19809,N_16519,N_17667);
and U19810 (N_19810,N_18059,N_18444);
nor U19811 (N_19811,N_15821,N_16535);
xor U19812 (N_19812,N_18283,N_17475);
or U19813 (N_19813,N_16658,N_18199);
nand U19814 (N_19814,N_16431,N_16031);
or U19815 (N_19815,N_16895,N_18202);
nand U19816 (N_19816,N_18330,N_16129);
or U19817 (N_19817,N_17873,N_15686);
nand U19818 (N_19818,N_17796,N_17833);
nand U19819 (N_19819,N_18189,N_17533);
xor U19820 (N_19820,N_18410,N_18688);
nand U19821 (N_19821,N_17482,N_16176);
nand U19822 (N_19822,N_17958,N_17209);
and U19823 (N_19823,N_17274,N_17595);
nand U19824 (N_19824,N_16989,N_18633);
xor U19825 (N_19825,N_16286,N_16700);
or U19826 (N_19826,N_18061,N_15848);
xnor U19827 (N_19827,N_15735,N_17625);
xor U19828 (N_19828,N_15811,N_17672);
nor U19829 (N_19829,N_16148,N_17613);
and U19830 (N_19830,N_15878,N_18311);
and U19831 (N_19831,N_16786,N_17823);
and U19832 (N_19832,N_16464,N_18254);
xor U19833 (N_19833,N_17266,N_18242);
nand U19834 (N_19834,N_18386,N_17049);
or U19835 (N_19835,N_16411,N_16511);
xor U19836 (N_19836,N_17709,N_18643);
nand U19837 (N_19837,N_16770,N_17593);
nor U19838 (N_19838,N_18180,N_16496);
xnor U19839 (N_19839,N_16415,N_18316);
nand U19840 (N_19840,N_15982,N_18149);
nand U19841 (N_19841,N_15733,N_17480);
and U19842 (N_19842,N_16479,N_18486);
nand U19843 (N_19843,N_17949,N_17888);
or U19844 (N_19844,N_18016,N_15656);
nor U19845 (N_19845,N_16996,N_16706);
xnor U19846 (N_19846,N_18052,N_17015);
nor U19847 (N_19847,N_15802,N_16150);
nor U19848 (N_19848,N_17296,N_16095);
and U19849 (N_19849,N_16057,N_16980);
and U19850 (N_19850,N_15816,N_16556);
nand U19851 (N_19851,N_18425,N_16299);
xor U19852 (N_19852,N_18730,N_17973);
and U19853 (N_19853,N_17950,N_17057);
xnor U19854 (N_19854,N_18072,N_17960);
xnor U19855 (N_19855,N_16847,N_16044);
xor U19856 (N_19856,N_15853,N_18718);
or U19857 (N_19857,N_18223,N_17807);
xor U19858 (N_19858,N_16395,N_15644);
xor U19859 (N_19859,N_18602,N_17387);
or U19860 (N_19860,N_18338,N_17166);
nand U19861 (N_19861,N_17169,N_18164);
xnor U19862 (N_19862,N_15664,N_16343);
nor U19863 (N_19863,N_16578,N_16384);
or U19864 (N_19864,N_18706,N_17004);
nor U19865 (N_19865,N_17716,N_16851);
nor U19866 (N_19866,N_18748,N_16235);
nor U19867 (N_19867,N_18458,N_16671);
nor U19868 (N_19868,N_18572,N_17652);
nor U19869 (N_19869,N_16907,N_18461);
and U19870 (N_19870,N_16889,N_17438);
xor U19871 (N_19871,N_16883,N_18054);
nor U19872 (N_19872,N_16783,N_15722);
or U19873 (N_19873,N_16372,N_17521);
nor U19874 (N_19874,N_18025,N_16881);
xnor U19875 (N_19875,N_15834,N_17564);
nand U19876 (N_19876,N_18264,N_18156);
and U19877 (N_19877,N_17686,N_17744);
nand U19878 (N_19878,N_18257,N_18654);
nor U19879 (N_19879,N_16062,N_18130);
nor U19880 (N_19880,N_17225,N_18426);
nand U19881 (N_19881,N_18094,N_15927);
and U19882 (N_19882,N_17650,N_15657);
and U19883 (N_19883,N_16657,N_15716);
or U19884 (N_19884,N_18652,N_15689);
and U19885 (N_19885,N_16261,N_17048);
or U19886 (N_19886,N_17079,N_17720);
and U19887 (N_19887,N_18373,N_17190);
nand U19888 (N_19888,N_18474,N_18628);
nand U19889 (N_19889,N_16088,N_17200);
nand U19890 (N_19890,N_17631,N_17992);
nand U19891 (N_19891,N_16757,N_17702);
and U19892 (N_19892,N_17069,N_17910);
xor U19893 (N_19893,N_16420,N_18744);
nand U19894 (N_19894,N_17097,N_17309);
or U19895 (N_19895,N_18408,N_15732);
or U19896 (N_19896,N_16078,N_16525);
nor U19897 (N_19897,N_17362,N_15826);
xor U19898 (N_19898,N_16956,N_16845);
xor U19899 (N_19899,N_16645,N_18512);
and U19900 (N_19900,N_16099,N_15997);
nand U19901 (N_19901,N_17431,N_16979);
and U19902 (N_19902,N_18519,N_16863);
xnor U19903 (N_19903,N_18209,N_16684);
or U19904 (N_19904,N_16135,N_15842);
nor U19905 (N_19905,N_17731,N_17643);
or U19906 (N_19906,N_17904,N_16522);
or U19907 (N_19907,N_17657,N_15692);
xor U19908 (N_19908,N_18630,N_16746);
nor U19909 (N_19909,N_18428,N_18487);
or U19910 (N_19910,N_18253,N_17816);
or U19911 (N_19911,N_17059,N_17358);
xor U19912 (N_19912,N_17027,N_15724);
nand U19913 (N_19913,N_18495,N_18012);
and U19914 (N_19914,N_16733,N_15877);
and U19915 (N_19915,N_18632,N_18036);
xnor U19916 (N_19916,N_18594,N_16185);
xor U19917 (N_19917,N_17468,N_18259);
nand U19918 (N_19918,N_17258,N_18192);
nand U19919 (N_19919,N_16195,N_16293);
nand U19920 (N_19920,N_16238,N_17275);
or U19921 (N_19921,N_18368,N_15843);
or U19922 (N_19922,N_16055,N_16660);
or U19923 (N_19923,N_17242,N_16092);
or U19924 (N_19924,N_16574,N_18142);
nand U19925 (N_19925,N_18342,N_16073);
nor U19926 (N_19926,N_16017,N_16045);
or U19927 (N_19927,N_18420,N_18044);
xnor U19928 (N_19928,N_18369,N_17857);
nor U19929 (N_19929,N_17916,N_18674);
xnor U19930 (N_19930,N_18050,N_17582);
xor U19931 (N_19931,N_16110,N_17450);
nand U19932 (N_19932,N_15740,N_17330);
xor U19933 (N_19933,N_17712,N_15739);
nor U19934 (N_19934,N_17229,N_18274);
or U19935 (N_19935,N_16383,N_18451);
nor U19936 (N_19936,N_18134,N_16039);
xor U19937 (N_19937,N_17348,N_18470);
xnor U19938 (N_19938,N_17055,N_18062);
and U19939 (N_19939,N_17815,N_16607);
nand U19940 (N_19940,N_15855,N_16663);
xnor U19941 (N_19941,N_16380,N_16567);
nand U19942 (N_19942,N_17531,N_18021);
and U19943 (N_19943,N_16424,N_16731);
or U19944 (N_19944,N_17538,N_16797);
nor U19945 (N_19945,N_16149,N_17769);
or U19946 (N_19946,N_16324,N_15870);
or U19947 (N_19947,N_17347,N_16037);
or U19948 (N_19948,N_18497,N_18152);
and U19949 (N_19949,N_18186,N_16566);
or U19950 (N_19950,N_16313,N_17763);
nor U19951 (N_19951,N_16087,N_17742);
nor U19952 (N_19952,N_18194,N_15701);
xnor U19953 (N_19953,N_15630,N_16214);
nand U19954 (N_19954,N_16692,N_16448);
or U19955 (N_19955,N_17071,N_16404);
nand U19956 (N_19956,N_17999,N_18505);
and U19957 (N_19957,N_17921,N_17173);
and U19958 (N_19958,N_18713,N_17029);
xnor U19959 (N_19959,N_16074,N_16760);
nor U19960 (N_19960,N_18336,N_15846);
and U19961 (N_19961,N_17326,N_17256);
and U19962 (N_19962,N_16181,N_18023);
nand U19963 (N_19963,N_16916,N_17346);
nand U19964 (N_19964,N_16977,N_18739);
xor U19965 (N_19965,N_17618,N_18527);
and U19966 (N_19966,N_16632,N_17733);
nand U19967 (N_19967,N_17022,N_17781);
and U19968 (N_19968,N_18115,N_16462);
nor U19969 (N_19969,N_16203,N_17235);
nor U19970 (N_19970,N_18123,N_17753);
or U19971 (N_19971,N_16807,N_16650);
nor U19972 (N_19972,N_15641,N_18268);
and U19973 (N_19973,N_16581,N_17710);
xnor U19974 (N_19974,N_18008,N_17969);
nand U19975 (N_19975,N_17050,N_18366);
nor U19976 (N_19976,N_15975,N_15936);
nand U19977 (N_19977,N_16174,N_18627);
or U19978 (N_19978,N_16546,N_18620);
xor U19979 (N_19979,N_18698,N_16365);
nor U19980 (N_19980,N_17528,N_16435);
nor U19981 (N_19981,N_16867,N_17659);
or U19982 (N_19982,N_18658,N_17971);
nand U19983 (N_19983,N_17598,N_18335);
or U19984 (N_19984,N_17547,N_17998);
nor U19985 (N_19985,N_18625,N_16951);
or U19986 (N_19986,N_18017,N_17335);
nand U19987 (N_19987,N_18320,N_16104);
or U19988 (N_19988,N_16750,N_17442);
nand U19989 (N_19989,N_17734,N_17523);
or U19990 (N_19990,N_15743,N_17490);
nor U19991 (N_19991,N_16843,N_16865);
xnor U19992 (N_19992,N_16929,N_15934);
or U19993 (N_19993,N_18604,N_16554);
xor U19994 (N_19994,N_16931,N_16988);
or U19995 (N_19995,N_16559,N_17041);
or U19996 (N_19996,N_18378,N_15738);
xor U19997 (N_19997,N_17179,N_16614);
or U19998 (N_19998,N_17817,N_17364);
or U19999 (N_19999,N_16640,N_17287);
nor U20000 (N_20000,N_17168,N_17770);
nand U20001 (N_20001,N_18278,N_17336);
and U20002 (N_20002,N_17852,N_18300);
and U20003 (N_20003,N_18166,N_16647);
xnor U20004 (N_20004,N_17851,N_17945);
or U20005 (N_20005,N_15758,N_18204);
nand U20006 (N_20006,N_17934,N_17074);
xor U20007 (N_20007,N_17145,N_16653);
and U20008 (N_20008,N_17647,N_17792);
xnor U20009 (N_20009,N_17206,N_15654);
nand U20010 (N_20010,N_17026,N_17901);
nand U20011 (N_20011,N_17060,N_15949);
nor U20012 (N_20012,N_16818,N_15813);
nor U20013 (N_20013,N_15688,N_16815);
nand U20014 (N_20014,N_18619,N_16884);
nor U20015 (N_20015,N_17630,N_17344);
xor U20016 (N_20016,N_15913,N_18457);
xor U20017 (N_20017,N_18394,N_18395);
and U20018 (N_20018,N_17535,N_17842);
nand U20019 (N_20019,N_16855,N_15715);
and U20020 (N_20020,N_17627,N_15714);
nand U20021 (N_20021,N_16379,N_18227);
xnor U20022 (N_20022,N_17573,N_16561);
nor U20023 (N_20023,N_18234,N_18371);
or U20024 (N_20024,N_18151,N_15736);
or U20025 (N_20025,N_16633,N_16136);
nand U20026 (N_20026,N_17052,N_17761);
xor U20027 (N_20027,N_18694,N_16381);
or U20028 (N_20028,N_15915,N_17828);
nand U20029 (N_20029,N_16047,N_17502);
nand U20030 (N_20030,N_17938,N_17597);
xor U20031 (N_20031,N_17941,N_17223);
and U20032 (N_20032,N_18172,N_17300);
or U20033 (N_20033,N_15702,N_18525);
nand U20034 (N_20034,N_15727,N_18165);
nand U20035 (N_20035,N_18463,N_15806);
nand U20036 (N_20036,N_17125,N_16474);
or U20037 (N_20037,N_18747,N_18421);
nor U20038 (N_20038,N_16480,N_17911);
nor U20039 (N_20039,N_18267,N_17058);
xor U20040 (N_20040,N_17312,N_17376);
or U20041 (N_20041,N_17314,N_16545);
xor U20042 (N_20042,N_17678,N_17795);
and U20043 (N_20043,N_17946,N_15831);
xnor U20044 (N_20044,N_16716,N_18438);
or U20045 (N_20045,N_18590,N_17890);
nor U20046 (N_20046,N_18280,N_18397);
or U20047 (N_20047,N_17163,N_17935);
or U20048 (N_20048,N_16806,N_17416);
and U20049 (N_20049,N_16364,N_16543);
and U20050 (N_20050,N_17038,N_16418);
xnor U20051 (N_20051,N_16239,N_18593);
and U20052 (N_20052,N_15680,N_16277);
xnor U20053 (N_20053,N_17118,N_17177);
and U20054 (N_20054,N_18591,N_16890);
and U20055 (N_20055,N_16677,N_17691);
nand U20056 (N_20056,N_17552,N_18255);
xor U20057 (N_20057,N_16445,N_18676);
nor U20058 (N_20058,N_16629,N_16894);
and U20059 (N_20059,N_16140,N_18022);
or U20060 (N_20060,N_17308,N_16893);
and U20061 (N_20061,N_16955,N_16167);
xor U20062 (N_20062,N_18314,N_16992);
nand U20063 (N_20063,N_17306,N_16861);
nand U20064 (N_20064,N_15850,N_17491);
or U20065 (N_20065,N_15661,N_16844);
nand U20066 (N_20066,N_15696,N_17064);
or U20067 (N_20067,N_17033,N_16305);
or U20068 (N_20068,N_17107,N_16856);
nand U20069 (N_20069,N_18701,N_17896);
nor U20070 (N_20070,N_18333,N_17199);
and U20071 (N_20071,N_18405,N_18442);
or U20072 (N_20072,N_18167,N_17165);
xnor U20073 (N_20073,N_16233,N_17505);
or U20074 (N_20074,N_16723,N_17497);
nor U20075 (N_20075,N_18616,N_18303);
or U20076 (N_20076,N_17359,N_16376);
nor U20077 (N_20077,N_17837,N_16836);
or U20078 (N_20078,N_16537,N_16042);
or U20079 (N_20079,N_18441,N_17586);
or U20080 (N_20080,N_16013,N_17171);
or U20081 (N_20081,N_17109,N_17994);
xor U20082 (N_20082,N_17785,N_17683);
nand U20083 (N_20083,N_17676,N_17965);
nand U20084 (N_20084,N_16459,N_18249);
and U20085 (N_20085,N_18547,N_17077);
or U20086 (N_20086,N_15844,N_18437);
and U20087 (N_20087,N_17599,N_16914);
and U20088 (N_20088,N_16180,N_17654);
or U20089 (N_20089,N_17831,N_17210);
or U20090 (N_20090,N_17180,N_17739);
nor U20091 (N_20091,N_17699,N_16298);
and U20092 (N_20092,N_16585,N_17867);
or U20093 (N_20093,N_18700,N_16637);
xnor U20094 (N_20094,N_16373,N_17964);
and U20095 (N_20095,N_15767,N_16052);
and U20096 (N_20096,N_18047,N_17003);
nor U20097 (N_20097,N_17407,N_16218);
and U20098 (N_20098,N_18157,N_17143);
and U20099 (N_20099,N_16003,N_16538);
xor U20100 (N_20100,N_17748,N_16027);
and U20101 (N_20101,N_17469,N_17232);
nor U20102 (N_20102,N_18200,N_18740);
or U20103 (N_20103,N_18090,N_17092);
nand U20104 (N_20104,N_17445,N_16880);
and U20105 (N_20105,N_16749,N_17542);
xnor U20106 (N_20106,N_17764,N_16352);
nor U20107 (N_20107,N_16330,N_17578);
nand U20108 (N_20108,N_16408,N_17656);
nand U20109 (N_20109,N_16795,N_18359);
nor U20110 (N_20110,N_18248,N_17838);
nand U20111 (N_20111,N_17492,N_17626);
xor U20112 (N_20112,N_16729,N_17424);
or U20113 (N_20113,N_18065,N_18110);
or U20114 (N_20114,N_16006,N_17226);
xnor U20115 (N_20115,N_16636,N_16982);
xor U20116 (N_20116,N_17080,N_18502);
and U20117 (N_20117,N_16217,N_15989);
and U20118 (N_20118,N_18678,N_15679);
and U20119 (N_20119,N_15638,N_16278);
and U20120 (N_20120,N_17410,N_17725);
xor U20121 (N_20121,N_18720,N_15665);
or U20122 (N_20122,N_18120,N_16046);
nand U20123 (N_20123,N_15895,N_18418);
nor U20124 (N_20124,N_17299,N_16121);
nand U20125 (N_20125,N_15717,N_17977);
or U20126 (N_20126,N_17997,N_17990);
or U20127 (N_20127,N_16097,N_17741);
nand U20128 (N_20128,N_16608,N_16024);
xor U20129 (N_20129,N_17749,N_16788);
and U20130 (N_20130,N_18295,N_18339);
nand U20131 (N_20131,N_17403,N_15861);
nor U20132 (N_20132,N_18533,N_18031);
nand U20133 (N_20133,N_16681,N_15899);
and U20134 (N_20134,N_17230,N_17777);
xor U20135 (N_20135,N_17090,N_17116);
xor U20136 (N_20136,N_18287,N_18323);
and U20137 (N_20137,N_18737,N_16272);
nor U20138 (N_20138,N_18681,N_16000);
xnor U20139 (N_20139,N_18404,N_18086);
xor U20140 (N_20140,N_15977,N_16091);
and U20141 (N_20141,N_15789,N_16503);
and U20142 (N_20142,N_15747,N_16885);
nand U20143 (N_20143,N_17164,N_16772);
or U20144 (N_20144,N_16661,N_15876);
or U20145 (N_20145,N_17955,N_16991);
xor U20146 (N_20146,N_17660,N_17776);
nor U20147 (N_20147,N_16449,N_16433);
nor U20148 (N_20148,N_16882,N_15791);
nand U20149 (N_20149,N_18173,N_17252);
and U20150 (N_20150,N_16621,N_15705);
nor U20151 (N_20151,N_18276,N_16564);
and U20152 (N_20152,N_15755,N_16579);
xor U20153 (N_20153,N_16114,N_15832);
nor U20154 (N_20154,N_15765,N_18372);
nor U20155 (N_20155,N_17587,N_16958);
nor U20156 (N_20156,N_18400,N_17401);
or U20157 (N_20157,N_18493,N_17767);
and U20158 (N_20158,N_16034,N_16222);
or U20159 (N_20159,N_15902,N_17801);
xor U20160 (N_20160,N_18609,N_16524);
nand U20161 (N_20161,N_16357,N_17113);
xor U20162 (N_20162,N_18040,N_17006);
or U20163 (N_20163,N_15974,N_15971);
nand U20164 (N_20164,N_16508,N_18191);
xor U20165 (N_20165,N_16145,N_15788);
or U20166 (N_20166,N_17752,N_17920);
xnor U20167 (N_20167,N_16888,N_16280);
nor U20168 (N_20168,N_18743,N_18001);
xor U20169 (N_20169,N_18669,N_18450);
nand U20170 (N_20170,N_16619,N_16224);
or U20171 (N_20171,N_18150,N_15986);
nor U20172 (N_20172,N_17591,N_17481);
or U20173 (N_20173,N_16905,N_17713);
xnor U20174 (N_20174,N_15822,N_18485);
or U20175 (N_20175,N_17585,N_17453);
and U20176 (N_20176,N_16536,N_16707);
xor U20177 (N_20177,N_18587,N_16056);
nor U20178 (N_20178,N_18118,N_17980);
or U20179 (N_20179,N_16595,N_16919);
or U20180 (N_20180,N_16190,N_16702);
nand U20181 (N_20181,N_16127,N_15729);
nand U20182 (N_20182,N_15652,N_17556);
nor U20183 (N_20183,N_16915,N_15893);
nor U20184 (N_20184,N_18567,N_15660);
xnor U20185 (N_20185,N_16854,N_15817);
xnor U20186 (N_20186,N_17117,N_18402);
or U20187 (N_20187,N_16341,N_15976);
nor U20188 (N_20188,N_18516,N_16838);
or U20189 (N_20189,N_17827,N_17254);
or U20190 (N_20190,N_15928,N_17608);
and U20191 (N_20191,N_17737,N_18613);
xor U20192 (N_20192,N_16157,N_18677);
or U20193 (N_20193,N_18552,N_16739);
nand U20194 (N_20194,N_17227,N_17067);
nor U20195 (N_20195,N_15946,N_17264);
xnor U20196 (N_20196,N_18158,N_15868);
or U20197 (N_20197,N_15858,N_16374);
or U20198 (N_20198,N_16023,N_16583);
nor U20199 (N_20199,N_18193,N_16386);
nand U20200 (N_20200,N_18510,N_15835);
and U20201 (N_20201,N_16470,N_16412);
or U20202 (N_20202,N_15920,N_17487);
nor U20203 (N_20203,N_18390,N_16421);
and U20204 (N_20204,N_17433,N_18175);
xnor U20205 (N_20205,N_16325,N_17007);
xnor U20206 (N_20206,N_17624,N_18215);
nor U20207 (N_20207,N_16780,N_18665);
or U20208 (N_20208,N_16516,N_17234);
xor U20209 (N_20209,N_18431,N_16674);
or U20210 (N_20210,N_18230,N_18672);
or U20211 (N_20211,N_17649,N_17286);
and U20212 (N_20212,N_18184,N_18411);
xor U20213 (N_20213,N_17793,N_16701);
xor U20214 (N_20214,N_15658,N_18244);
nand U20215 (N_20215,N_15862,N_17126);
and U20216 (N_20216,N_17201,N_16631);
xor U20217 (N_20217,N_15993,N_15910);
nor U20218 (N_20218,N_16502,N_17818);
nand U20219 (N_20219,N_17703,N_17115);
and U20220 (N_20220,N_16710,N_15757);
nor U20221 (N_20221,N_18382,N_17861);
and U20222 (N_20222,N_15957,N_18306);
nor U20223 (N_20223,N_17231,N_18051);
xnor U20224 (N_20224,N_18292,N_18349);
or U20225 (N_20225,N_17987,N_18640);
and U20226 (N_20226,N_18326,N_17121);
and U20227 (N_20227,N_16173,N_17021);
nand U20228 (N_20228,N_15704,N_17757);
and U20229 (N_20229,N_17907,N_18707);
nand U20230 (N_20230,N_16998,N_16494);
and U20231 (N_20231,N_17530,N_17981);
or U20232 (N_20232,N_17023,N_17131);
xor U20233 (N_20233,N_16128,N_16670);
or U20234 (N_20234,N_18732,N_18327);
and U20235 (N_20235,N_16691,N_17328);
nor U20236 (N_20236,N_16282,N_18636);
or U20237 (N_20237,N_15771,N_16304);
nand U20238 (N_20238,N_15951,N_17357);
nor U20239 (N_20239,N_17493,N_16336);
xnor U20240 (N_20240,N_15753,N_17662);
nor U20241 (N_20241,N_17930,N_18066);
and U20242 (N_20242,N_16544,N_17520);
nand U20243 (N_20243,N_17812,N_18562);
or U20244 (N_20244,N_16891,N_18245);
nor U20245 (N_20245,N_17009,N_16035);
nand U20246 (N_20246,N_18205,N_18509);
and U20247 (N_20247,N_17290,N_16927);
and U20248 (N_20248,N_16548,N_18082);
xnor U20249 (N_20249,N_17758,N_16577);
nor U20250 (N_20250,N_16064,N_17897);
nor U20251 (N_20251,N_17332,N_16455);
nor U20252 (N_20252,N_16294,N_17688);
nand U20253 (N_20253,N_16531,N_15994);
nor U20254 (N_20254,N_16291,N_16973);
xnor U20255 (N_20255,N_16077,N_15937);
xnor U20256 (N_20256,N_16603,N_18137);
nand U20257 (N_20257,N_16215,N_17280);
xnor U20258 (N_20258,N_18453,N_17775);
xor U20259 (N_20259,N_16080,N_15637);
and U20260 (N_20260,N_17187,N_15933);
nand U20261 (N_20261,N_16816,N_16950);
nand U20262 (N_20262,N_16038,N_17174);
or U20263 (N_20263,N_18600,N_16020);
xnor U20264 (N_20264,N_17774,N_18555);
nand U20265 (N_20265,N_16231,N_17470);
nor U20266 (N_20266,N_18449,N_18500);
nand U20267 (N_20267,N_16276,N_16152);
and U20268 (N_20268,N_17213,N_18143);
xor U20269 (N_20269,N_17895,N_15728);
and U20270 (N_20270,N_17717,N_17885);
and U20271 (N_20271,N_17313,N_16105);
nand U20272 (N_20272,N_16839,N_17272);
nand U20273 (N_20273,N_18518,N_18731);
and U20274 (N_20274,N_17550,N_16164);
or U20275 (N_20275,N_15939,N_16197);
nor U20276 (N_20276,N_18504,N_16935);
nor U20277 (N_20277,N_18027,N_18481);
nor U20278 (N_20278,N_15912,N_17665);
nor U20279 (N_20279,N_16925,N_16146);
or U20280 (N_20280,N_18005,N_15745);
nor U20281 (N_20281,N_17285,N_15695);
nor U20282 (N_20282,N_18686,N_17517);
or U20283 (N_20283,N_18673,N_18471);
nor U20284 (N_20284,N_17217,N_18468);
nor U20285 (N_20285,N_17024,N_16400);
nor U20286 (N_20286,N_15697,N_18656);
and U20287 (N_20287,N_18136,N_16943);
xor U20288 (N_20288,N_17400,N_17804);
or U20289 (N_20289,N_17513,N_17919);
and U20290 (N_20290,N_15812,N_17966);
or U20291 (N_20291,N_15942,N_17506);
nand U20292 (N_20292,N_18389,N_16685);
xor U20293 (N_20293,N_16643,N_17134);
nand U20294 (N_20294,N_16001,N_17461);
xor U20295 (N_20295,N_17500,N_18589);
or U20296 (N_20296,N_17191,N_16375);
and U20297 (N_20297,N_17906,N_16416);
nor U20298 (N_20298,N_17615,N_18596);
or U20299 (N_20299,N_18076,N_16358);
nand U20300 (N_20300,N_15859,N_16510);
nand U20301 (N_20301,N_15670,N_18697);
or U20302 (N_20302,N_17413,N_18736);
nor U20303 (N_20303,N_16285,N_17360);
and U20304 (N_20304,N_18653,N_17298);
and U20305 (N_20305,N_16668,N_17194);
nand U20306 (N_20306,N_17352,N_18401);
and U20307 (N_20307,N_16930,N_16377);
xnor U20308 (N_20308,N_16618,N_17565);
and U20309 (N_20309,N_18586,N_18080);
xor U20310 (N_20310,N_15906,N_17452);
nor U20311 (N_20311,N_17913,N_18571);
or U20312 (N_20312,N_16481,N_15902);
nor U20313 (N_20313,N_16224,N_17158);
nand U20314 (N_20314,N_17038,N_15878);
xor U20315 (N_20315,N_15631,N_15663);
and U20316 (N_20316,N_18629,N_17778);
xor U20317 (N_20317,N_17762,N_17412);
and U20318 (N_20318,N_15885,N_15709);
nor U20319 (N_20319,N_16972,N_16832);
and U20320 (N_20320,N_17380,N_16006);
or U20321 (N_20321,N_18236,N_15919);
nor U20322 (N_20322,N_17717,N_15702);
and U20323 (N_20323,N_17266,N_16325);
nand U20324 (N_20324,N_16562,N_17893);
nand U20325 (N_20325,N_18035,N_16508);
nor U20326 (N_20326,N_18093,N_15947);
and U20327 (N_20327,N_17194,N_18143);
and U20328 (N_20328,N_16022,N_15883);
nor U20329 (N_20329,N_18468,N_17843);
xor U20330 (N_20330,N_16518,N_15917);
xnor U20331 (N_20331,N_18457,N_15935);
or U20332 (N_20332,N_15738,N_18449);
nor U20333 (N_20333,N_17376,N_16895);
xor U20334 (N_20334,N_17909,N_18189);
xor U20335 (N_20335,N_17846,N_18730);
nand U20336 (N_20336,N_16023,N_15879);
or U20337 (N_20337,N_17012,N_18358);
nand U20338 (N_20338,N_16163,N_16215);
xor U20339 (N_20339,N_15639,N_16481);
or U20340 (N_20340,N_17601,N_16735);
nand U20341 (N_20341,N_16829,N_16479);
nand U20342 (N_20342,N_16138,N_16682);
nand U20343 (N_20343,N_18065,N_18408);
and U20344 (N_20344,N_18224,N_17207);
nor U20345 (N_20345,N_16325,N_15782);
xor U20346 (N_20346,N_17448,N_16701);
and U20347 (N_20347,N_17010,N_17351);
nor U20348 (N_20348,N_16011,N_16409);
xnor U20349 (N_20349,N_16267,N_16887);
xnor U20350 (N_20350,N_16764,N_16845);
or U20351 (N_20351,N_17711,N_18130);
and U20352 (N_20352,N_16317,N_17661);
nor U20353 (N_20353,N_17016,N_15990);
nor U20354 (N_20354,N_17659,N_16799);
or U20355 (N_20355,N_16043,N_16970);
nor U20356 (N_20356,N_16890,N_18441);
and U20357 (N_20357,N_15709,N_16273);
xor U20358 (N_20358,N_17492,N_18299);
and U20359 (N_20359,N_18029,N_18687);
xor U20360 (N_20360,N_16137,N_16517);
nand U20361 (N_20361,N_17758,N_16394);
xor U20362 (N_20362,N_18337,N_18585);
and U20363 (N_20363,N_17560,N_17773);
and U20364 (N_20364,N_17227,N_17986);
xnor U20365 (N_20365,N_15857,N_16466);
nor U20366 (N_20366,N_17599,N_18407);
and U20367 (N_20367,N_17575,N_16056);
nand U20368 (N_20368,N_16622,N_18143);
xnor U20369 (N_20369,N_15774,N_17110);
nor U20370 (N_20370,N_16948,N_17659);
nand U20371 (N_20371,N_18069,N_16265);
and U20372 (N_20372,N_17283,N_17659);
and U20373 (N_20373,N_16532,N_18259);
nor U20374 (N_20374,N_17064,N_18689);
nor U20375 (N_20375,N_18362,N_18161);
and U20376 (N_20376,N_16571,N_18259);
and U20377 (N_20377,N_17060,N_17522);
or U20378 (N_20378,N_16132,N_17471);
and U20379 (N_20379,N_18400,N_17569);
nor U20380 (N_20380,N_16466,N_15729);
nand U20381 (N_20381,N_18280,N_17685);
and U20382 (N_20382,N_16307,N_18255);
nor U20383 (N_20383,N_16473,N_16510);
xor U20384 (N_20384,N_16747,N_17914);
nand U20385 (N_20385,N_15876,N_18339);
nor U20386 (N_20386,N_17892,N_16288);
nor U20387 (N_20387,N_18394,N_15638);
and U20388 (N_20388,N_16589,N_18444);
and U20389 (N_20389,N_17669,N_16040);
xnor U20390 (N_20390,N_18606,N_17965);
xor U20391 (N_20391,N_16550,N_15726);
nand U20392 (N_20392,N_17361,N_15797);
nor U20393 (N_20393,N_18517,N_17976);
nand U20394 (N_20394,N_16439,N_18469);
or U20395 (N_20395,N_18325,N_15677);
or U20396 (N_20396,N_17511,N_18068);
xor U20397 (N_20397,N_15738,N_16102);
or U20398 (N_20398,N_17583,N_16545);
or U20399 (N_20399,N_15974,N_18153);
nor U20400 (N_20400,N_15638,N_18186);
and U20401 (N_20401,N_18697,N_15829);
nor U20402 (N_20402,N_16232,N_17733);
nor U20403 (N_20403,N_16935,N_15928);
nand U20404 (N_20404,N_17407,N_17953);
and U20405 (N_20405,N_17439,N_15636);
and U20406 (N_20406,N_17890,N_16606);
nor U20407 (N_20407,N_17249,N_17313);
or U20408 (N_20408,N_17083,N_17897);
xnor U20409 (N_20409,N_16796,N_18710);
or U20410 (N_20410,N_16820,N_17912);
or U20411 (N_20411,N_17259,N_18007);
nand U20412 (N_20412,N_16106,N_15735);
xnor U20413 (N_20413,N_16471,N_16364);
or U20414 (N_20414,N_17936,N_17421);
or U20415 (N_20415,N_16555,N_18707);
nand U20416 (N_20416,N_17720,N_16881);
nand U20417 (N_20417,N_17141,N_18384);
xnor U20418 (N_20418,N_18104,N_16591);
nand U20419 (N_20419,N_16173,N_18026);
and U20420 (N_20420,N_17068,N_17679);
or U20421 (N_20421,N_16865,N_16524);
nand U20422 (N_20422,N_16009,N_17151);
or U20423 (N_20423,N_18744,N_15692);
or U20424 (N_20424,N_18727,N_17218);
or U20425 (N_20425,N_16004,N_18686);
nor U20426 (N_20426,N_16880,N_16423);
xor U20427 (N_20427,N_16219,N_17667);
nand U20428 (N_20428,N_18055,N_17430);
nor U20429 (N_20429,N_17805,N_17432);
nor U20430 (N_20430,N_16742,N_16332);
xnor U20431 (N_20431,N_18458,N_17575);
or U20432 (N_20432,N_16276,N_17715);
or U20433 (N_20433,N_18209,N_17141);
or U20434 (N_20434,N_17275,N_17130);
nor U20435 (N_20435,N_17674,N_15918);
nor U20436 (N_20436,N_16017,N_17927);
xor U20437 (N_20437,N_17042,N_18545);
xnor U20438 (N_20438,N_16726,N_15746);
or U20439 (N_20439,N_18376,N_17646);
nor U20440 (N_20440,N_17768,N_16625);
xor U20441 (N_20441,N_18282,N_15872);
nor U20442 (N_20442,N_17284,N_16694);
xor U20443 (N_20443,N_16674,N_16752);
nand U20444 (N_20444,N_15986,N_18181);
and U20445 (N_20445,N_16858,N_16199);
nor U20446 (N_20446,N_18251,N_16517);
nand U20447 (N_20447,N_15823,N_17499);
or U20448 (N_20448,N_16689,N_17023);
nor U20449 (N_20449,N_17306,N_18636);
nor U20450 (N_20450,N_18591,N_18746);
and U20451 (N_20451,N_17411,N_17932);
nor U20452 (N_20452,N_16249,N_17211);
and U20453 (N_20453,N_17153,N_17556);
nor U20454 (N_20454,N_18177,N_16027);
nor U20455 (N_20455,N_16086,N_17847);
or U20456 (N_20456,N_16206,N_17076);
and U20457 (N_20457,N_16227,N_17031);
and U20458 (N_20458,N_18190,N_16232);
or U20459 (N_20459,N_16168,N_18198);
nor U20460 (N_20460,N_16313,N_18227);
or U20461 (N_20461,N_16697,N_16684);
and U20462 (N_20462,N_15759,N_16362);
and U20463 (N_20463,N_17042,N_17915);
nor U20464 (N_20464,N_18417,N_16267);
nand U20465 (N_20465,N_16001,N_16649);
nand U20466 (N_20466,N_16030,N_18697);
nand U20467 (N_20467,N_16993,N_18316);
xnor U20468 (N_20468,N_17113,N_18174);
nor U20469 (N_20469,N_18539,N_15839);
nor U20470 (N_20470,N_16914,N_18276);
xor U20471 (N_20471,N_17549,N_17805);
and U20472 (N_20472,N_18702,N_18279);
and U20473 (N_20473,N_15676,N_16817);
nand U20474 (N_20474,N_17558,N_17145);
xor U20475 (N_20475,N_16203,N_17301);
nor U20476 (N_20476,N_17185,N_18641);
nand U20477 (N_20477,N_15844,N_18569);
nor U20478 (N_20478,N_18305,N_18053);
or U20479 (N_20479,N_16580,N_18157);
nand U20480 (N_20480,N_17134,N_16489);
and U20481 (N_20481,N_18386,N_17751);
or U20482 (N_20482,N_15838,N_18393);
and U20483 (N_20483,N_18122,N_18168);
xnor U20484 (N_20484,N_16098,N_16923);
nand U20485 (N_20485,N_17308,N_16485);
or U20486 (N_20486,N_16705,N_17616);
or U20487 (N_20487,N_16896,N_17687);
nor U20488 (N_20488,N_17696,N_17451);
and U20489 (N_20489,N_17178,N_15647);
or U20490 (N_20490,N_15800,N_15663);
or U20491 (N_20491,N_18583,N_17705);
and U20492 (N_20492,N_16072,N_16672);
and U20493 (N_20493,N_17441,N_16790);
xor U20494 (N_20494,N_17258,N_17188);
or U20495 (N_20495,N_16821,N_17973);
nand U20496 (N_20496,N_18033,N_16493);
nor U20497 (N_20497,N_15777,N_17639);
and U20498 (N_20498,N_15845,N_18741);
nand U20499 (N_20499,N_17743,N_17406);
and U20500 (N_20500,N_15980,N_15824);
and U20501 (N_20501,N_16623,N_16505);
xor U20502 (N_20502,N_15829,N_17167);
and U20503 (N_20503,N_18712,N_18089);
nand U20504 (N_20504,N_15652,N_16769);
and U20505 (N_20505,N_16228,N_17277);
and U20506 (N_20506,N_17702,N_17562);
xnor U20507 (N_20507,N_16435,N_18066);
xor U20508 (N_20508,N_15659,N_17467);
nor U20509 (N_20509,N_16089,N_16733);
and U20510 (N_20510,N_16045,N_18537);
nor U20511 (N_20511,N_16203,N_18464);
and U20512 (N_20512,N_17316,N_18004);
nor U20513 (N_20513,N_15965,N_16116);
nand U20514 (N_20514,N_16484,N_15838);
nor U20515 (N_20515,N_16651,N_15867);
nand U20516 (N_20516,N_15879,N_18147);
or U20517 (N_20517,N_17126,N_17746);
xnor U20518 (N_20518,N_16126,N_17130);
nand U20519 (N_20519,N_15637,N_16419);
xnor U20520 (N_20520,N_16633,N_17708);
or U20521 (N_20521,N_16320,N_18409);
or U20522 (N_20522,N_15752,N_16612);
or U20523 (N_20523,N_17922,N_15987);
nand U20524 (N_20524,N_16163,N_18497);
and U20525 (N_20525,N_18629,N_16059);
or U20526 (N_20526,N_18108,N_16777);
and U20527 (N_20527,N_17858,N_18677);
nor U20528 (N_20528,N_18335,N_17415);
xor U20529 (N_20529,N_16414,N_18034);
and U20530 (N_20530,N_16677,N_17854);
nor U20531 (N_20531,N_18504,N_16945);
or U20532 (N_20532,N_17560,N_18226);
nand U20533 (N_20533,N_18657,N_16306);
or U20534 (N_20534,N_15888,N_15976);
or U20535 (N_20535,N_18128,N_16448);
and U20536 (N_20536,N_15844,N_16969);
nand U20537 (N_20537,N_18401,N_16705);
nand U20538 (N_20538,N_18595,N_16513);
nand U20539 (N_20539,N_15825,N_16355);
and U20540 (N_20540,N_17120,N_18701);
nor U20541 (N_20541,N_17568,N_16172);
and U20542 (N_20542,N_15749,N_16735);
or U20543 (N_20543,N_16487,N_15631);
nor U20544 (N_20544,N_18115,N_16938);
nor U20545 (N_20545,N_16097,N_18227);
nor U20546 (N_20546,N_17037,N_17596);
and U20547 (N_20547,N_17632,N_16039);
nand U20548 (N_20548,N_17215,N_18475);
nand U20549 (N_20549,N_18455,N_17650);
nor U20550 (N_20550,N_18420,N_17737);
nor U20551 (N_20551,N_18650,N_16929);
nand U20552 (N_20552,N_17817,N_16331);
nand U20553 (N_20553,N_16025,N_17020);
nor U20554 (N_20554,N_17063,N_17456);
xor U20555 (N_20555,N_17659,N_16754);
xnor U20556 (N_20556,N_17308,N_18087);
xnor U20557 (N_20557,N_17132,N_17181);
xor U20558 (N_20558,N_16469,N_15971);
xor U20559 (N_20559,N_15783,N_16320);
nor U20560 (N_20560,N_17009,N_17604);
or U20561 (N_20561,N_17509,N_15803);
nand U20562 (N_20562,N_18429,N_15869);
xnor U20563 (N_20563,N_16737,N_16891);
nand U20564 (N_20564,N_16151,N_18695);
xnor U20565 (N_20565,N_16033,N_18656);
xor U20566 (N_20566,N_17210,N_18012);
and U20567 (N_20567,N_16220,N_18211);
and U20568 (N_20568,N_15910,N_16618);
xnor U20569 (N_20569,N_17091,N_17184);
xor U20570 (N_20570,N_17482,N_17275);
xor U20571 (N_20571,N_16680,N_17852);
and U20572 (N_20572,N_18294,N_17793);
nor U20573 (N_20573,N_17626,N_17766);
xor U20574 (N_20574,N_17475,N_18643);
and U20575 (N_20575,N_15848,N_15857);
and U20576 (N_20576,N_17250,N_16664);
and U20577 (N_20577,N_16148,N_15984);
nor U20578 (N_20578,N_18246,N_16368);
nand U20579 (N_20579,N_18523,N_15984);
nand U20580 (N_20580,N_17658,N_15693);
xnor U20581 (N_20581,N_15772,N_18490);
or U20582 (N_20582,N_15977,N_16267);
nor U20583 (N_20583,N_15840,N_18749);
nand U20584 (N_20584,N_18467,N_16444);
xnor U20585 (N_20585,N_17831,N_18423);
nor U20586 (N_20586,N_15634,N_16846);
or U20587 (N_20587,N_16468,N_16798);
nand U20588 (N_20588,N_17699,N_17484);
and U20589 (N_20589,N_16244,N_15833);
or U20590 (N_20590,N_17066,N_16545);
xnor U20591 (N_20591,N_16606,N_16391);
xor U20592 (N_20592,N_17064,N_16036);
nand U20593 (N_20593,N_18710,N_17414);
xor U20594 (N_20594,N_18556,N_16449);
xnor U20595 (N_20595,N_15840,N_15965);
and U20596 (N_20596,N_17326,N_16847);
or U20597 (N_20597,N_18109,N_18294);
nand U20598 (N_20598,N_17672,N_16007);
xor U20599 (N_20599,N_16594,N_16906);
nand U20600 (N_20600,N_17571,N_17242);
nor U20601 (N_20601,N_16656,N_18115);
or U20602 (N_20602,N_15764,N_16662);
xor U20603 (N_20603,N_17694,N_16448);
xor U20604 (N_20604,N_15763,N_17503);
and U20605 (N_20605,N_15646,N_17364);
nor U20606 (N_20606,N_18136,N_15849);
or U20607 (N_20607,N_17177,N_17459);
nor U20608 (N_20608,N_15776,N_17538);
nand U20609 (N_20609,N_17120,N_17416);
nor U20610 (N_20610,N_18444,N_16578);
nor U20611 (N_20611,N_18310,N_16364);
xor U20612 (N_20612,N_16666,N_18031);
or U20613 (N_20613,N_15921,N_17003);
nor U20614 (N_20614,N_15817,N_17859);
xnor U20615 (N_20615,N_16958,N_18067);
nor U20616 (N_20616,N_18605,N_15929);
xnor U20617 (N_20617,N_16203,N_17786);
or U20618 (N_20618,N_16542,N_18433);
nor U20619 (N_20619,N_18373,N_18506);
nor U20620 (N_20620,N_17856,N_17301);
xnor U20621 (N_20621,N_16835,N_17963);
nor U20622 (N_20622,N_16423,N_15716);
xor U20623 (N_20623,N_16751,N_18030);
or U20624 (N_20624,N_16518,N_18038);
nor U20625 (N_20625,N_17099,N_18709);
and U20626 (N_20626,N_18703,N_18426);
nand U20627 (N_20627,N_16390,N_18131);
or U20628 (N_20628,N_15755,N_17892);
nand U20629 (N_20629,N_18621,N_15760);
and U20630 (N_20630,N_18508,N_17965);
and U20631 (N_20631,N_17205,N_17654);
nor U20632 (N_20632,N_16793,N_18331);
or U20633 (N_20633,N_16301,N_18386);
nor U20634 (N_20634,N_17799,N_17368);
or U20635 (N_20635,N_15685,N_17905);
or U20636 (N_20636,N_17490,N_15681);
xnor U20637 (N_20637,N_15628,N_17840);
nor U20638 (N_20638,N_18061,N_17891);
nor U20639 (N_20639,N_18200,N_18668);
xor U20640 (N_20640,N_18499,N_18138);
or U20641 (N_20641,N_17081,N_17209);
or U20642 (N_20642,N_18705,N_15788);
xor U20643 (N_20643,N_16614,N_18632);
xnor U20644 (N_20644,N_16928,N_16301);
nor U20645 (N_20645,N_16332,N_16669);
nand U20646 (N_20646,N_16427,N_16624);
nor U20647 (N_20647,N_18535,N_17539);
or U20648 (N_20648,N_17315,N_17062);
nor U20649 (N_20649,N_15963,N_16245);
or U20650 (N_20650,N_18116,N_16538);
nand U20651 (N_20651,N_16720,N_15687);
nor U20652 (N_20652,N_17743,N_18105);
nand U20653 (N_20653,N_16800,N_17500);
or U20654 (N_20654,N_16405,N_18448);
xor U20655 (N_20655,N_18447,N_17112);
or U20656 (N_20656,N_16247,N_16979);
or U20657 (N_20657,N_16219,N_16788);
nor U20658 (N_20658,N_15877,N_18551);
nand U20659 (N_20659,N_18032,N_18711);
or U20660 (N_20660,N_17474,N_16014);
or U20661 (N_20661,N_16803,N_18185);
nand U20662 (N_20662,N_18169,N_15805);
xnor U20663 (N_20663,N_18730,N_16433);
or U20664 (N_20664,N_16457,N_16876);
and U20665 (N_20665,N_17236,N_16117);
and U20666 (N_20666,N_17449,N_15943);
and U20667 (N_20667,N_18114,N_18735);
or U20668 (N_20668,N_17867,N_16544);
xnor U20669 (N_20669,N_17680,N_17131);
and U20670 (N_20670,N_16708,N_16924);
nand U20671 (N_20671,N_16983,N_16476);
or U20672 (N_20672,N_17703,N_17500);
and U20673 (N_20673,N_15999,N_16075);
or U20674 (N_20674,N_15645,N_17370);
and U20675 (N_20675,N_15908,N_17591);
xor U20676 (N_20676,N_16800,N_16767);
nor U20677 (N_20677,N_18328,N_15801);
xor U20678 (N_20678,N_15865,N_16231);
and U20679 (N_20679,N_18173,N_16210);
xnor U20680 (N_20680,N_17127,N_18477);
nor U20681 (N_20681,N_17302,N_16870);
and U20682 (N_20682,N_18027,N_16035);
nand U20683 (N_20683,N_16950,N_16310);
and U20684 (N_20684,N_18345,N_17930);
xor U20685 (N_20685,N_18142,N_15963);
or U20686 (N_20686,N_15838,N_16367);
and U20687 (N_20687,N_17374,N_18732);
and U20688 (N_20688,N_18407,N_16510);
or U20689 (N_20689,N_16331,N_16794);
or U20690 (N_20690,N_17387,N_16538);
xor U20691 (N_20691,N_18132,N_17287);
xor U20692 (N_20692,N_18243,N_16948);
and U20693 (N_20693,N_15829,N_18217);
xor U20694 (N_20694,N_16116,N_18325);
nand U20695 (N_20695,N_17980,N_17202);
or U20696 (N_20696,N_16251,N_15722);
or U20697 (N_20697,N_16769,N_16697);
xnor U20698 (N_20698,N_18192,N_15978);
nor U20699 (N_20699,N_18005,N_17224);
nand U20700 (N_20700,N_17719,N_16150);
nand U20701 (N_20701,N_16617,N_16990);
nand U20702 (N_20702,N_18404,N_18388);
and U20703 (N_20703,N_16263,N_17097);
and U20704 (N_20704,N_16183,N_18494);
xor U20705 (N_20705,N_16243,N_18590);
or U20706 (N_20706,N_16760,N_18666);
and U20707 (N_20707,N_16398,N_15711);
xnor U20708 (N_20708,N_16395,N_15637);
or U20709 (N_20709,N_16770,N_17662);
and U20710 (N_20710,N_16178,N_18706);
nor U20711 (N_20711,N_16313,N_16412);
xnor U20712 (N_20712,N_18589,N_17386);
xor U20713 (N_20713,N_17973,N_18156);
nor U20714 (N_20714,N_16419,N_18661);
and U20715 (N_20715,N_15639,N_15787);
and U20716 (N_20716,N_18627,N_17578);
and U20717 (N_20717,N_16517,N_18384);
nand U20718 (N_20718,N_17527,N_17428);
nor U20719 (N_20719,N_16669,N_18082);
nor U20720 (N_20720,N_16641,N_17554);
or U20721 (N_20721,N_17840,N_17709);
nand U20722 (N_20722,N_17532,N_15668);
nand U20723 (N_20723,N_17735,N_16422);
nand U20724 (N_20724,N_15638,N_16440);
nor U20725 (N_20725,N_17257,N_17061);
nor U20726 (N_20726,N_16051,N_16134);
nand U20727 (N_20727,N_17017,N_15851);
xnor U20728 (N_20728,N_17566,N_18299);
nor U20729 (N_20729,N_17825,N_17550);
nor U20730 (N_20730,N_18211,N_16634);
nor U20731 (N_20731,N_17865,N_18554);
or U20732 (N_20732,N_17273,N_16163);
or U20733 (N_20733,N_18640,N_15840);
nor U20734 (N_20734,N_15855,N_18140);
or U20735 (N_20735,N_17682,N_18469);
or U20736 (N_20736,N_18394,N_17683);
nor U20737 (N_20737,N_16290,N_16249);
or U20738 (N_20738,N_15955,N_16627);
or U20739 (N_20739,N_17402,N_16625);
xnor U20740 (N_20740,N_15691,N_18307);
xor U20741 (N_20741,N_16888,N_18466);
nor U20742 (N_20742,N_15690,N_16295);
or U20743 (N_20743,N_16464,N_17691);
or U20744 (N_20744,N_17379,N_18299);
nor U20745 (N_20745,N_18185,N_17492);
and U20746 (N_20746,N_17390,N_18336);
or U20747 (N_20747,N_16045,N_18434);
nor U20748 (N_20748,N_17521,N_18086);
or U20749 (N_20749,N_15714,N_18130);
or U20750 (N_20750,N_18591,N_15672);
xnor U20751 (N_20751,N_18513,N_17649);
nand U20752 (N_20752,N_16970,N_18272);
xor U20753 (N_20753,N_18686,N_18512);
or U20754 (N_20754,N_17663,N_18407);
and U20755 (N_20755,N_16382,N_16054);
nor U20756 (N_20756,N_18333,N_17342);
and U20757 (N_20757,N_17891,N_16372);
nand U20758 (N_20758,N_18243,N_16196);
or U20759 (N_20759,N_16830,N_16190);
xnor U20760 (N_20760,N_18158,N_18252);
or U20761 (N_20761,N_16185,N_16938);
xor U20762 (N_20762,N_18214,N_18689);
nor U20763 (N_20763,N_16521,N_16251);
or U20764 (N_20764,N_17534,N_16374);
or U20765 (N_20765,N_17229,N_17247);
xor U20766 (N_20766,N_17121,N_18001);
nand U20767 (N_20767,N_18468,N_17127);
or U20768 (N_20768,N_18429,N_18562);
nand U20769 (N_20769,N_16607,N_16682);
or U20770 (N_20770,N_16644,N_17272);
xnor U20771 (N_20771,N_17016,N_16556);
and U20772 (N_20772,N_17908,N_18433);
or U20773 (N_20773,N_18542,N_18655);
or U20774 (N_20774,N_16756,N_16221);
or U20775 (N_20775,N_18039,N_17753);
and U20776 (N_20776,N_17711,N_17905);
nor U20777 (N_20777,N_18661,N_17691);
xnor U20778 (N_20778,N_18248,N_16331);
xor U20779 (N_20779,N_16966,N_17727);
nand U20780 (N_20780,N_18161,N_16919);
or U20781 (N_20781,N_18597,N_16101);
xnor U20782 (N_20782,N_17534,N_17224);
or U20783 (N_20783,N_16981,N_16018);
xnor U20784 (N_20784,N_18737,N_17482);
nand U20785 (N_20785,N_17219,N_18098);
and U20786 (N_20786,N_16084,N_16052);
or U20787 (N_20787,N_16996,N_18087);
xnor U20788 (N_20788,N_18052,N_15653);
nor U20789 (N_20789,N_17383,N_17067);
or U20790 (N_20790,N_16814,N_17031);
nor U20791 (N_20791,N_17347,N_15692);
nor U20792 (N_20792,N_17125,N_16206);
xor U20793 (N_20793,N_17949,N_17084);
xor U20794 (N_20794,N_16016,N_15825);
and U20795 (N_20795,N_16753,N_18667);
and U20796 (N_20796,N_16708,N_17379);
nor U20797 (N_20797,N_18422,N_18564);
nand U20798 (N_20798,N_18456,N_17787);
nand U20799 (N_20799,N_17422,N_17369);
or U20800 (N_20800,N_18376,N_17305);
or U20801 (N_20801,N_15870,N_17947);
xor U20802 (N_20802,N_17518,N_17337);
nand U20803 (N_20803,N_15991,N_18342);
or U20804 (N_20804,N_17420,N_17409);
or U20805 (N_20805,N_18265,N_17740);
nor U20806 (N_20806,N_16336,N_18196);
and U20807 (N_20807,N_16699,N_18545);
xor U20808 (N_20808,N_18478,N_18089);
or U20809 (N_20809,N_17911,N_17632);
nand U20810 (N_20810,N_17870,N_18495);
or U20811 (N_20811,N_17691,N_16610);
nor U20812 (N_20812,N_16353,N_16158);
or U20813 (N_20813,N_16238,N_16566);
nand U20814 (N_20814,N_17486,N_16879);
nor U20815 (N_20815,N_18208,N_18631);
xnor U20816 (N_20816,N_15826,N_17755);
or U20817 (N_20817,N_17835,N_16067);
or U20818 (N_20818,N_18407,N_15798);
and U20819 (N_20819,N_16414,N_15992);
or U20820 (N_20820,N_17844,N_16120);
xor U20821 (N_20821,N_16665,N_18044);
and U20822 (N_20822,N_17595,N_17638);
nand U20823 (N_20823,N_15901,N_18425);
nor U20824 (N_20824,N_16027,N_18618);
nor U20825 (N_20825,N_17674,N_17205);
nand U20826 (N_20826,N_15797,N_18609);
xnor U20827 (N_20827,N_18154,N_15693);
xor U20828 (N_20828,N_18323,N_18609);
xnor U20829 (N_20829,N_16766,N_16081);
nor U20830 (N_20830,N_18445,N_15804);
xor U20831 (N_20831,N_18706,N_18212);
nand U20832 (N_20832,N_16215,N_18621);
nand U20833 (N_20833,N_16731,N_16418);
nor U20834 (N_20834,N_17872,N_16331);
xor U20835 (N_20835,N_18376,N_17435);
nand U20836 (N_20836,N_17270,N_16943);
nor U20837 (N_20837,N_17911,N_16739);
nand U20838 (N_20838,N_16776,N_17576);
nand U20839 (N_20839,N_17209,N_18396);
nand U20840 (N_20840,N_16790,N_16953);
and U20841 (N_20841,N_16900,N_17601);
and U20842 (N_20842,N_16784,N_16624);
and U20843 (N_20843,N_16013,N_18179);
xor U20844 (N_20844,N_17135,N_18603);
nor U20845 (N_20845,N_16959,N_17374);
xor U20846 (N_20846,N_16831,N_17733);
nor U20847 (N_20847,N_16782,N_18367);
nor U20848 (N_20848,N_17067,N_17136);
or U20849 (N_20849,N_18509,N_18174);
or U20850 (N_20850,N_17056,N_18398);
and U20851 (N_20851,N_16793,N_16482);
xor U20852 (N_20852,N_18471,N_18273);
nor U20853 (N_20853,N_16746,N_16271);
or U20854 (N_20854,N_16334,N_17758);
and U20855 (N_20855,N_17183,N_16201);
or U20856 (N_20856,N_16258,N_16282);
or U20857 (N_20857,N_16583,N_15812);
and U20858 (N_20858,N_17263,N_16061);
or U20859 (N_20859,N_16379,N_16180);
nor U20860 (N_20860,N_16671,N_16262);
or U20861 (N_20861,N_18483,N_16343);
nand U20862 (N_20862,N_17831,N_16429);
nand U20863 (N_20863,N_17860,N_15640);
nor U20864 (N_20864,N_18208,N_16789);
nand U20865 (N_20865,N_17124,N_15795);
and U20866 (N_20866,N_15962,N_17853);
xnor U20867 (N_20867,N_16373,N_18587);
xnor U20868 (N_20868,N_17549,N_15707);
xor U20869 (N_20869,N_18636,N_17221);
nand U20870 (N_20870,N_18560,N_16464);
nand U20871 (N_20871,N_16857,N_16459);
nor U20872 (N_20872,N_18017,N_16469);
xnor U20873 (N_20873,N_18082,N_15671);
and U20874 (N_20874,N_17094,N_17255);
and U20875 (N_20875,N_17837,N_18540);
and U20876 (N_20876,N_18342,N_15994);
nor U20877 (N_20877,N_16812,N_18159);
xor U20878 (N_20878,N_17874,N_18633);
and U20879 (N_20879,N_15983,N_18464);
nor U20880 (N_20880,N_18550,N_17931);
nand U20881 (N_20881,N_16019,N_15692);
nand U20882 (N_20882,N_17961,N_15853);
xnor U20883 (N_20883,N_16836,N_17954);
nor U20884 (N_20884,N_16634,N_15625);
nand U20885 (N_20885,N_16188,N_18247);
nand U20886 (N_20886,N_18375,N_16800);
and U20887 (N_20887,N_16655,N_17595);
or U20888 (N_20888,N_16113,N_16420);
nand U20889 (N_20889,N_18150,N_17237);
and U20890 (N_20890,N_15676,N_16130);
or U20891 (N_20891,N_17913,N_16197);
xnor U20892 (N_20892,N_16938,N_18623);
xnor U20893 (N_20893,N_18002,N_18202);
or U20894 (N_20894,N_18726,N_16318);
and U20895 (N_20895,N_18286,N_15767);
nor U20896 (N_20896,N_17106,N_16198);
nand U20897 (N_20897,N_17345,N_17177);
and U20898 (N_20898,N_17212,N_17475);
or U20899 (N_20899,N_15848,N_16125);
or U20900 (N_20900,N_17785,N_17867);
xnor U20901 (N_20901,N_18041,N_18740);
xor U20902 (N_20902,N_15837,N_16607);
xnor U20903 (N_20903,N_17759,N_15758);
nand U20904 (N_20904,N_17185,N_17700);
and U20905 (N_20905,N_16442,N_17950);
nor U20906 (N_20906,N_17156,N_16833);
or U20907 (N_20907,N_16712,N_16786);
nor U20908 (N_20908,N_17818,N_17789);
nor U20909 (N_20909,N_17329,N_17668);
and U20910 (N_20910,N_16732,N_17703);
nand U20911 (N_20911,N_18320,N_16794);
xor U20912 (N_20912,N_15826,N_17541);
nand U20913 (N_20913,N_18681,N_18743);
and U20914 (N_20914,N_18405,N_18344);
nand U20915 (N_20915,N_16524,N_15828);
nand U20916 (N_20916,N_18576,N_16322);
and U20917 (N_20917,N_15838,N_17260);
nand U20918 (N_20918,N_17951,N_18359);
or U20919 (N_20919,N_15977,N_18372);
nand U20920 (N_20920,N_15961,N_17095);
or U20921 (N_20921,N_15882,N_18041);
nand U20922 (N_20922,N_16949,N_18203);
nor U20923 (N_20923,N_17097,N_15899);
and U20924 (N_20924,N_16927,N_16723);
xor U20925 (N_20925,N_18060,N_16138);
or U20926 (N_20926,N_16402,N_18380);
or U20927 (N_20927,N_16114,N_17212);
and U20928 (N_20928,N_17104,N_17597);
nor U20929 (N_20929,N_16467,N_18664);
xor U20930 (N_20930,N_15659,N_17226);
or U20931 (N_20931,N_15665,N_16072);
nor U20932 (N_20932,N_17874,N_18138);
xor U20933 (N_20933,N_17546,N_17625);
nor U20934 (N_20934,N_16358,N_16749);
nand U20935 (N_20935,N_15711,N_18108);
xor U20936 (N_20936,N_17251,N_18560);
nor U20937 (N_20937,N_17399,N_16623);
xor U20938 (N_20938,N_17751,N_17320);
xor U20939 (N_20939,N_17149,N_17310);
nor U20940 (N_20940,N_18180,N_18366);
and U20941 (N_20941,N_17449,N_16892);
or U20942 (N_20942,N_16011,N_16131);
xnor U20943 (N_20943,N_18144,N_15929);
nand U20944 (N_20944,N_16742,N_17345);
and U20945 (N_20945,N_15804,N_17429);
nand U20946 (N_20946,N_18078,N_16979);
nor U20947 (N_20947,N_17857,N_18729);
nand U20948 (N_20948,N_18187,N_16337);
and U20949 (N_20949,N_16751,N_15838);
nor U20950 (N_20950,N_17693,N_18011);
nand U20951 (N_20951,N_15902,N_15807);
xnor U20952 (N_20952,N_18681,N_17567);
xnor U20953 (N_20953,N_18731,N_18639);
nand U20954 (N_20954,N_16173,N_18049);
or U20955 (N_20955,N_16890,N_16493);
and U20956 (N_20956,N_17322,N_17204);
nand U20957 (N_20957,N_16872,N_17211);
nor U20958 (N_20958,N_18745,N_16366);
and U20959 (N_20959,N_16138,N_18744);
or U20960 (N_20960,N_16183,N_17842);
nand U20961 (N_20961,N_18465,N_18576);
nand U20962 (N_20962,N_16017,N_18575);
xnor U20963 (N_20963,N_16438,N_16194);
xor U20964 (N_20964,N_18272,N_15874);
nand U20965 (N_20965,N_16554,N_16516);
and U20966 (N_20966,N_18559,N_17744);
xor U20967 (N_20967,N_17059,N_16481);
or U20968 (N_20968,N_16812,N_18356);
nand U20969 (N_20969,N_15705,N_18088);
nand U20970 (N_20970,N_16988,N_16183);
nand U20971 (N_20971,N_16730,N_16866);
or U20972 (N_20972,N_17712,N_15670);
and U20973 (N_20973,N_18615,N_18594);
nor U20974 (N_20974,N_16844,N_18276);
nand U20975 (N_20975,N_16615,N_18134);
and U20976 (N_20976,N_15707,N_16127);
nand U20977 (N_20977,N_16840,N_15701);
or U20978 (N_20978,N_17014,N_16753);
or U20979 (N_20979,N_16891,N_17332);
or U20980 (N_20980,N_17601,N_16722);
or U20981 (N_20981,N_17572,N_15837);
or U20982 (N_20982,N_15673,N_17080);
and U20983 (N_20983,N_17404,N_17860);
and U20984 (N_20984,N_16221,N_17920);
and U20985 (N_20985,N_18306,N_16854);
or U20986 (N_20986,N_16005,N_18354);
xnor U20987 (N_20987,N_17526,N_16904);
or U20988 (N_20988,N_18259,N_15812);
nor U20989 (N_20989,N_17610,N_18436);
and U20990 (N_20990,N_17898,N_16058);
and U20991 (N_20991,N_17469,N_17882);
or U20992 (N_20992,N_16858,N_16959);
and U20993 (N_20993,N_16461,N_16164);
xnor U20994 (N_20994,N_18464,N_17224);
nor U20995 (N_20995,N_17862,N_16639);
nor U20996 (N_20996,N_17603,N_18498);
and U20997 (N_20997,N_18053,N_18683);
xnor U20998 (N_20998,N_17768,N_17812);
nor U20999 (N_20999,N_18300,N_16953);
xnor U21000 (N_21000,N_17162,N_17882);
or U21001 (N_21001,N_16849,N_16583);
nor U21002 (N_21002,N_18386,N_17358);
or U21003 (N_21003,N_15730,N_17117);
xnor U21004 (N_21004,N_18240,N_17740);
xor U21005 (N_21005,N_15708,N_17873);
xor U21006 (N_21006,N_17562,N_17043);
or U21007 (N_21007,N_17549,N_16156);
nor U21008 (N_21008,N_16405,N_17614);
nand U21009 (N_21009,N_15809,N_18737);
nand U21010 (N_21010,N_17024,N_17719);
xnor U21011 (N_21011,N_18284,N_18288);
and U21012 (N_21012,N_17026,N_18479);
or U21013 (N_21013,N_16023,N_18659);
and U21014 (N_21014,N_18600,N_15634);
xor U21015 (N_21015,N_16920,N_16721);
nor U21016 (N_21016,N_16313,N_18270);
or U21017 (N_21017,N_17825,N_18419);
or U21018 (N_21018,N_18600,N_17893);
xor U21019 (N_21019,N_17716,N_18494);
nor U21020 (N_21020,N_16247,N_18275);
and U21021 (N_21021,N_16015,N_17041);
nand U21022 (N_21022,N_18131,N_16684);
nor U21023 (N_21023,N_16114,N_16620);
xnor U21024 (N_21024,N_16692,N_17893);
nor U21025 (N_21025,N_15797,N_15747);
xor U21026 (N_21026,N_18721,N_16731);
nor U21027 (N_21027,N_18073,N_17971);
and U21028 (N_21028,N_17285,N_16747);
and U21029 (N_21029,N_17733,N_16802);
or U21030 (N_21030,N_16476,N_17070);
nor U21031 (N_21031,N_18521,N_16430);
or U21032 (N_21032,N_18438,N_15859);
nand U21033 (N_21033,N_18531,N_17713);
nor U21034 (N_21034,N_17076,N_15772);
and U21035 (N_21035,N_17180,N_16167);
nor U21036 (N_21036,N_15628,N_17935);
xnor U21037 (N_21037,N_18182,N_16149);
nor U21038 (N_21038,N_18099,N_15977);
nand U21039 (N_21039,N_17219,N_15846);
nor U21040 (N_21040,N_17066,N_16866);
or U21041 (N_21041,N_17769,N_16081);
and U21042 (N_21042,N_16895,N_17401);
xor U21043 (N_21043,N_17221,N_15633);
nor U21044 (N_21044,N_17881,N_17181);
nor U21045 (N_21045,N_17107,N_17836);
and U21046 (N_21046,N_17120,N_18387);
xnor U21047 (N_21047,N_15886,N_17695);
nand U21048 (N_21048,N_16779,N_17214);
xor U21049 (N_21049,N_18442,N_17406);
nand U21050 (N_21050,N_18111,N_16683);
xor U21051 (N_21051,N_18079,N_16612);
xnor U21052 (N_21052,N_16731,N_18456);
or U21053 (N_21053,N_16508,N_17374);
or U21054 (N_21054,N_16100,N_16624);
xnor U21055 (N_21055,N_18449,N_16760);
and U21056 (N_21056,N_15762,N_18511);
nor U21057 (N_21057,N_17736,N_16095);
or U21058 (N_21058,N_16911,N_16156);
or U21059 (N_21059,N_16870,N_18239);
and U21060 (N_21060,N_16809,N_15803);
and U21061 (N_21061,N_18005,N_15815);
and U21062 (N_21062,N_18589,N_18640);
or U21063 (N_21063,N_16763,N_18463);
xnor U21064 (N_21064,N_16010,N_15983);
xor U21065 (N_21065,N_18221,N_17379);
nor U21066 (N_21066,N_16516,N_18608);
xor U21067 (N_21067,N_16756,N_17472);
nor U21068 (N_21068,N_16244,N_16091);
nand U21069 (N_21069,N_18698,N_17925);
nand U21070 (N_21070,N_18635,N_17178);
nand U21071 (N_21071,N_18260,N_16160);
nor U21072 (N_21072,N_18702,N_18297);
nor U21073 (N_21073,N_17605,N_16774);
nor U21074 (N_21074,N_16635,N_17346);
xnor U21075 (N_21075,N_16088,N_18260);
and U21076 (N_21076,N_18041,N_18496);
and U21077 (N_21077,N_17801,N_17111);
and U21078 (N_21078,N_16968,N_17235);
xnor U21079 (N_21079,N_18746,N_15804);
nand U21080 (N_21080,N_18208,N_16841);
xnor U21081 (N_21081,N_16787,N_18034);
xor U21082 (N_21082,N_16082,N_18540);
nand U21083 (N_21083,N_16777,N_15978);
nand U21084 (N_21084,N_17027,N_17502);
and U21085 (N_21085,N_17773,N_17744);
nand U21086 (N_21086,N_18710,N_15906);
nor U21087 (N_21087,N_15891,N_16486);
nor U21088 (N_21088,N_16256,N_16850);
or U21089 (N_21089,N_17594,N_16500);
xor U21090 (N_21090,N_16903,N_17786);
nand U21091 (N_21091,N_16076,N_16253);
nand U21092 (N_21092,N_17469,N_18399);
xor U21093 (N_21093,N_15661,N_16490);
and U21094 (N_21094,N_17924,N_18324);
nand U21095 (N_21095,N_16647,N_17799);
or U21096 (N_21096,N_16822,N_16156);
xor U21097 (N_21097,N_17956,N_18321);
nand U21098 (N_21098,N_15871,N_15790);
or U21099 (N_21099,N_17454,N_18571);
nor U21100 (N_21100,N_17176,N_18431);
nor U21101 (N_21101,N_17771,N_15781);
xnor U21102 (N_21102,N_17176,N_15988);
or U21103 (N_21103,N_16062,N_15967);
nand U21104 (N_21104,N_15808,N_17698);
nor U21105 (N_21105,N_17572,N_16943);
xnor U21106 (N_21106,N_18503,N_18329);
xnor U21107 (N_21107,N_15992,N_17510);
xnor U21108 (N_21108,N_17184,N_16812);
nand U21109 (N_21109,N_16046,N_18044);
or U21110 (N_21110,N_17324,N_16443);
and U21111 (N_21111,N_17513,N_18326);
nor U21112 (N_21112,N_18539,N_18061);
nor U21113 (N_21113,N_17192,N_16498);
xnor U21114 (N_21114,N_17692,N_17401);
and U21115 (N_21115,N_17208,N_16646);
nor U21116 (N_21116,N_17250,N_16678);
nand U21117 (N_21117,N_16292,N_16619);
or U21118 (N_21118,N_15994,N_16871);
xor U21119 (N_21119,N_17115,N_16516);
xnor U21120 (N_21120,N_16286,N_18308);
nor U21121 (N_21121,N_16126,N_18308);
or U21122 (N_21122,N_18412,N_18056);
and U21123 (N_21123,N_16638,N_15824);
xnor U21124 (N_21124,N_15811,N_17608);
and U21125 (N_21125,N_17941,N_16688);
nand U21126 (N_21126,N_16705,N_15893);
xnor U21127 (N_21127,N_18650,N_16610);
and U21128 (N_21128,N_18405,N_18449);
and U21129 (N_21129,N_17647,N_16356);
nor U21130 (N_21130,N_17445,N_18713);
xor U21131 (N_21131,N_15930,N_15647);
and U21132 (N_21132,N_18609,N_17932);
or U21133 (N_21133,N_18666,N_18710);
or U21134 (N_21134,N_18709,N_17860);
nand U21135 (N_21135,N_17451,N_17060);
and U21136 (N_21136,N_17143,N_15649);
xor U21137 (N_21137,N_16625,N_18411);
and U21138 (N_21138,N_17824,N_18633);
and U21139 (N_21139,N_18446,N_17974);
nor U21140 (N_21140,N_16731,N_18201);
xnor U21141 (N_21141,N_15872,N_16323);
or U21142 (N_21142,N_15928,N_15772);
xnor U21143 (N_21143,N_17744,N_16272);
and U21144 (N_21144,N_18243,N_18533);
or U21145 (N_21145,N_15772,N_16441);
and U21146 (N_21146,N_18405,N_16856);
xnor U21147 (N_21147,N_17136,N_16153);
and U21148 (N_21148,N_15668,N_17131);
nor U21149 (N_21149,N_18427,N_18099);
nor U21150 (N_21150,N_18187,N_18194);
nor U21151 (N_21151,N_18450,N_17198);
xnor U21152 (N_21152,N_18540,N_16786);
nor U21153 (N_21153,N_15665,N_16142);
or U21154 (N_21154,N_17040,N_18401);
or U21155 (N_21155,N_17666,N_17981);
or U21156 (N_21156,N_17975,N_16728);
or U21157 (N_21157,N_17182,N_16986);
nand U21158 (N_21158,N_16923,N_15728);
nor U21159 (N_21159,N_16271,N_15683);
nor U21160 (N_21160,N_15665,N_17052);
nand U21161 (N_21161,N_16008,N_18104);
xnor U21162 (N_21162,N_18284,N_15644);
xor U21163 (N_21163,N_16479,N_16183);
or U21164 (N_21164,N_16331,N_15882);
or U21165 (N_21165,N_16739,N_18442);
nand U21166 (N_21166,N_16840,N_18198);
and U21167 (N_21167,N_16790,N_16247);
and U21168 (N_21168,N_16623,N_16581);
and U21169 (N_21169,N_18748,N_16514);
nor U21170 (N_21170,N_15745,N_16903);
nand U21171 (N_21171,N_16392,N_15909);
nor U21172 (N_21172,N_16772,N_16418);
and U21173 (N_21173,N_18154,N_16133);
xnor U21174 (N_21174,N_16896,N_18310);
or U21175 (N_21175,N_18228,N_18584);
nor U21176 (N_21176,N_16116,N_16250);
nor U21177 (N_21177,N_18004,N_17641);
nand U21178 (N_21178,N_17792,N_18169);
and U21179 (N_21179,N_16166,N_17011);
or U21180 (N_21180,N_15910,N_16345);
nand U21181 (N_21181,N_18210,N_15644);
nand U21182 (N_21182,N_18639,N_17507);
nand U21183 (N_21183,N_17921,N_17880);
xor U21184 (N_21184,N_17387,N_18197);
nor U21185 (N_21185,N_16164,N_15980);
and U21186 (N_21186,N_16673,N_17814);
nor U21187 (N_21187,N_18240,N_17510);
nor U21188 (N_21188,N_17711,N_16008);
nand U21189 (N_21189,N_18570,N_16955);
and U21190 (N_21190,N_15810,N_17278);
nor U21191 (N_21191,N_17820,N_16535);
or U21192 (N_21192,N_18480,N_16400);
or U21193 (N_21193,N_16219,N_16960);
nor U21194 (N_21194,N_16567,N_17020);
and U21195 (N_21195,N_16452,N_16308);
nand U21196 (N_21196,N_18165,N_16303);
or U21197 (N_21197,N_17817,N_18328);
and U21198 (N_21198,N_16112,N_16034);
or U21199 (N_21199,N_15873,N_18229);
xnor U21200 (N_21200,N_17298,N_15753);
or U21201 (N_21201,N_16487,N_17879);
nand U21202 (N_21202,N_18191,N_18327);
nand U21203 (N_21203,N_17868,N_17045);
and U21204 (N_21204,N_17974,N_17980);
xor U21205 (N_21205,N_17272,N_18436);
and U21206 (N_21206,N_15844,N_17000);
nand U21207 (N_21207,N_17982,N_16507);
xnor U21208 (N_21208,N_18216,N_15919);
xor U21209 (N_21209,N_16862,N_16031);
or U21210 (N_21210,N_17321,N_17296);
or U21211 (N_21211,N_16609,N_18580);
xnor U21212 (N_21212,N_16361,N_16230);
nor U21213 (N_21213,N_18414,N_15773);
or U21214 (N_21214,N_17328,N_18513);
nand U21215 (N_21215,N_18554,N_17844);
nor U21216 (N_21216,N_17820,N_16475);
nand U21217 (N_21217,N_15668,N_16169);
or U21218 (N_21218,N_16921,N_16947);
nand U21219 (N_21219,N_16598,N_16171);
nor U21220 (N_21220,N_18738,N_16378);
or U21221 (N_21221,N_17055,N_17990);
nor U21222 (N_21222,N_17833,N_15831);
nand U21223 (N_21223,N_18658,N_17098);
and U21224 (N_21224,N_17785,N_16496);
nand U21225 (N_21225,N_17761,N_16414);
and U21226 (N_21226,N_17648,N_17892);
xor U21227 (N_21227,N_18018,N_16829);
nand U21228 (N_21228,N_15830,N_18589);
or U21229 (N_21229,N_18244,N_15911);
or U21230 (N_21230,N_16261,N_17716);
or U21231 (N_21231,N_18708,N_15824);
xor U21232 (N_21232,N_17866,N_16320);
and U21233 (N_21233,N_18298,N_18680);
nor U21234 (N_21234,N_18589,N_17520);
nand U21235 (N_21235,N_16470,N_18246);
and U21236 (N_21236,N_17244,N_18176);
and U21237 (N_21237,N_17786,N_16249);
or U21238 (N_21238,N_17611,N_18162);
and U21239 (N_21239,N_18159,N_17767);
and U21240 (N_21240,N_16689,N_18310);
and U21241 (N_21241,N_18260,N_16995);
xnor U21242 (N_21242,N_16356,N_17368);
nand U21243 (N_21243,N_17124,N_16854);
or U21244 (N_21244,N_16714,N_17701);
and U21245 (N_21245,N_16415,N_18270);
nand U21246 (N_21246,N_18312,N_18146);
nor U21247 (N_21247,N_17346,N_18457);
and U21248 (N_21248,N_18099,N_18563);
and U21249 (N_21249,N_17891,N_18567);
nor U21250 (N_21250,N_17438,N_18686);
or U21251 (N_21251,N_18616,N_16298);
or U21252 (N_21252,N_15822,N_16043);
and U21253 (N_21253,N_17956,N_16687);
nand U21254 (N_21254,N_16051,N_16797);
xnor U21255 (N_21255,N_15828,N_16270);
xor U21256 (N_21256,N_17462,N_17011);
nor U21257 (N_21257,N_18565,N_16003);
xnor U21258 (N_21258,N_17028,N_16413);
xnor U21259 (N_21259,N_16019,N_16462);
and U21260 (N_21260,N_17256,N_17333);
nand U21261 (N_21261,N_16605,N_16355);
nand U21262 (N_21262,N_15976,N_17343);
and U21263 (N_21263,N_17028,N_18667);
and U21264 (N_21264,N_16890,N_16720);
or U21265 (N_21265,N_18401,N_18402);
and U21266 (N_21266,N_17643,N_15647);
or U21267 (N_21267,N_16661,N_16986);
xor U21268 (N_21268,N_17374,N_15731);
nor U21269 (N_21269,N_17059,N_15735);
xnor U21270 (N_21270,N_17732,N_16329);
nand U21271 (N_21271,N_17038,N_17709);
xnor U21272 (N_21272,N_17152,N_18545);
or U21273 (N_21273,N_17647,N_16492);
nand U21274 (N_21274,N_18170,N_17155);
xnor U21275 (N_21275,N_16115,N_16012);
xnor U21276 (N_21276,N_15821,N_16753);
nor U21277 (N_21277,N_17897,N_16981);
nand U21278 (N_21278,N_16069,N_15931);
and U21279 (N_21279,N_16313,N_18368);
xor U21280 (N_21280,N_18631,N_17419);
or U21281 (N_21281,N_15683,N_18180);
nor U21282 (N_21282,N_16805,N_17347);
xnor U21283 (N_21283,N_17063,N_17572);
xnor U21284 (N_21284,N_18361,N_16740);
nand U21285 (N_21285,N_16306,N_15856);
nand U21286 (N_21286,N_18041,N_16346);
and U21287 (N_21287,N_17667,N_16547);
or U21288 (N_21288,N_16013,N_18326);
or U21289 (N_21289,N_17190,N_17922);
nor U21290 (N_21290,N_16515,N_17798);
or U21291 (N_21291,N_16455,N_16019);
nand U21292 (N_21292,N_16294,N_16650);
nor U21293 (N_21293,N_17296,N_17195);
nand U21294 (N_21294,N_17753,N_16006);
nor U21295 (N_21295,N_16405,N_18335);
or U21296 (N_21296,N_17325,N_16306);
and U21297 (N_21297,N_16624,N_16774);
or U21298 (N_21298,N_16559,N_15737);
nor U21299 (N_21299,N_16452,N_18447);
nand U21300 (N_21300,N_18628,N_18527);
or U21301 (N_21301,N_16251,N_15832);
nand U21302 (N_21302,N_18183,N_16245);
or U21303 (N_21303,N_18309,N_18619);
nor U21304 (N_21304,N_18704,N_18614);
xnor U21305 (N_21305,N_16969,N_16926);
or U21306 (N_21306,N_16101,N_17311);
or U21307 (N_21307,N_17664,N_18194);
xnor U21308 (N_21308,N_17739,N_17086);
nor U21309 (N_21309,N_17384,N_16776);
xnor U21310 (N_21310,N_16302,N_17805);
or U21311 (N_21311,N_18509,N_17705);
nor U21312 (N_21312,N_17360,N_17079);
nand U21313 (N_21313,N_15826,N_18188);
nor U21314 (N_21314,N_18127,N_17203);
nor U21315 (N_21315,N_17719,N_16053);
nor U21316 (N_21316,N_17299,N_16788);
or U21317 (N_21317,N_17668,N_16999);
nand U21318 (N_21318,N_17559,N_15851);
xor U21319 (N_21319,N_16672,N_18660);
nand U21320 (N_21320,N_18264,N_16046);
nor U21321 (N_21321,N_15780,N_17200);
nor U21322 (N_21322,N_17177,N_18435);
xnor U21323 (N_21323,N_17715,N_18463);
or U21324 (N_21324,N_16781,N_15989);
or U21325 (N_21325,N_18235,N_18364);
xnor U21326 (N_21326,N_15868,N_17955);
and U21327 (N_21327,N_15726,N_18308);
or U21328 (N_21328,N_18557,N_15668);
nand U21329 (N_21329,N_16214,N_16083);
nand U21330 (N_21330,N_16718,N_18440);
nor U21331 (N_21331,N_16749,N_16426);
nor U21332 (N_21332,N_16701,N_16423);
nor U21333 (N_21333,N_17350,N_17365);
nor U21334 (N_21334,N_16553,N_17293);
or U21335 (N_21335,N_17388,N_17613);
xor U21336 (N_21336,N_15978,N_17091);
nor U21337 (N_21337,N_18120,N_18044);
nor U21338 (N_21338,N_18735,N_17745);
xnor U21339 (N_21339,N_16524,N_17368);
nor U21340 (N_21340,N_17161,N_16040);
nand U21341 (N_21341,N_17105,N_16653);
nor U21342 (N_21342,N_17847,N_17355);
or U21343 (N_21343,N_17985,N_16151);
xor U21344 (N_21344,N_17423,N_18324);
nor U21345 (N_21345,N_18130,N_16045);
nand U21346 (N_21346,N_15802,N_16814);
xor U21347 (N_21347,N_18693,N_16929);
nand U21348 (N_21348,N_17868,N_16114);
nor U21349 (N_21349,N_18018,N_18083);
nand U21350 (N_21350,N_17707,N_18110);
nor U21351 (N_21351,N_17362,N_16945);
or U21352 (N_21352,N_17661,N_16420);
nor U21353 (N_21353,N_15778,N_18016);
or U21354 (N_21354,N_18542,N_18632);
or U21355 (N_21355,N_16707,N_16083);
or U21356 (N_21356,N_16598,N_17082);
nor U21357 (N_21357,N_17961,N_18571);
or U21358 (N_21358,N_16407,N_17986);
and U21359 (N_21359,N_17421,N_18282);
nor U21360 (N_21360,N_17799,N_17653);
nor U21361 (N_21361,N_15968,N_16907);
and U21362 (N_21362,N_16697,N_17306);
or U21363 (N_21363,N_15728,N_18589);
nand U21364 (N_21364,N_16039,N_17261);
or U21365 (N_21365,N_16237,N_17323);
nand U21366 (N_21366,N_18686,N_16775);
nor U21367 (N_21367,N_17959,N_17906);
or U21368 (N_21368,N_16900,N_17724);
nand U21369 (N_21369,N_16397,N_17222);
nand U21370 (N_21370,N_16864,N_17873);
nand U21371 (N_21371,N_16625,N_17197);
and U21372 (N_21372,N_18385,N_17404);
or U21373 (N_21373,N_16586,N_17567);
xnor U21374 (N_21374,N_17171,N_16693);
nor U21375 (N_21375,N_18354,N_16335);
xor U21376 (N_21376,N_15835,N_17910);
and U21377 (N_21377,N_18487,N_16296);
nor U21378 (N_21378,N_17463,N_16317);
or U21379 (N_21379,N_18736,N_16086);
nand U21380 (N_21380,N_17740,N_18386);
or U21381 (N_21381,N_16152,N_17487);
xor U21382 (N_21382,N_16851,N_15678);
nand U21383 (N_21383,N_17419,N_16284);
and U21384 (N_21384,N_17468,N_16512);
or U21385 (N_21385,N_15957,N_18537);
or U21386 (N_21386,N_16973,N_17750);
xnor U21387 (N_21387,N_17120,N_17666);
xnor U21388 (N_21388,N_17093,N_16789);
and U21389 (N_21389,N_16651,N_15803);
xnor U21390 (N_21390,N_15815,N_17715);
and U21391 (N_21391,N_17633,N_18209);
nor U21392 (N_21392,N_16105,N_17454);
or U21393 (N_21393,N_16328,N_15870);
and U21394 (N_21394,N_17846,N_16460);
and U21395 (N_21395,N_17495,N_16125);
or U21396 (N_21396,N_17770,N_16835);
nand U21397 (N_21397,N_17400,N_15903);
and U21398 (N_21398,N_16773,N_17895);
nand U21399 (N_21399,N_17456,N_17853);
or U21400 (N_21400,N_15934,N_16247);
nor U21401 (N_21401,N_17429,N_18466);
or U21402 (N_21402,N_17609,N_18574);
xnor U21403 (N_21403,N_17461,N_16861);
nor U21404 (N_21404,N_18069,N_18191);
or U21405 (N_21405,N_16567,N_17537);
nand U21406 (N_21406,N_17484,N_15682);
nand U21407 (N_21407,N_18654,N_16291);
nor U21408 (N_21408,N_17521,N_17152);
xor U21409 (N_21409,N_18722,N_18492);
nor U21410 (N_21410,N_18456,N_17782);
xnor U21411 (N_21411,N_16520,N_18643);
nand U21412 (N_21412,N_17840,N_15847);
or U21413 (N_21413,N_15663,N_16167);
or U21414 (N_21414,N_16914,N_16962);
nor U21415 (N_21415,N_16793,N_16149);
or U21416 (N_21416,N_16422,N_18621);
nor U21417 (N_21417,N_16580,N_17336);
nor U21418 (N_21418,N_16596,N_18135);
nor U21419 (N_21419,N_16686,N_18224);
nor U21420 (N_21420,N_15671,N_17127);
or U21421 (N_21421,N_18598,N_15963);
and U21422 (N_21422,N_18244,N_16320);
nor U21423 (N_21423,N_15920,N_17106);
xor U21424 (N_21424,N_16127,N_17429);
xor U21425 (N_21425,N_17110,N_16220);
nor U21426 (N_21426,N_16263,N_17102);
and U21427 (N_21427,N_17937,N_16700);
nand U21428 (N_21428,N_15649,N_15830);
xnor U21429 (N_21429,N_17196,N_16099);
nand U21430 (N_21430,N_17737,N_17692);
xnor U21431 (N_21431,N_17188,N_17496);
nor U21432 (N_21432,N_16449,N_16617);
and U21433 (N_21433,N_16543,N_16456);
nor U21434 (N_21434,N_16346,N_15780);
and U21435 (N_21435,N_15835,N_17874);
and U21436 (N_21436,N_18706,N_17922);
or U21437 (N_21437,N_17267,N_18227);
nand U21438 (N_21438,N_18361,N_16553);
xnor U21439 (N_21439,N_17394,N_15799);
nor U21440 (N_21440,N_16670,N_18311);
nor U21441 (N_21441,N_18489,N_18006);
nor U21442 (N_21442,N_17488,N_16839);
xnor U21443 (N_21443,N_18649,N_16429);
nor U21444 (N_21444,N_17825,N_18304);
or U21445 (N_21445,N_18463,N_17916);
xnor U21446 (N_21446,N_17870,N_18700);
nor U21447 (N_21447,N_15887,N_17147);
xnor U21448 (N_21448,N_18342,N_17797);
xor U21449 (N_21449,N_17981,N_16897);
xor U21450 (N_21450,N_15834,N_17862);
xor U21451 (N_21451,N_18320,N_16051);
nand U21452 (N_21452,N_18427,N_16276);
or U21453 (N_21453,N_16281,N_18296);
or U21454 (N_21454,N_15829,N_15667);
and U21455 (N_21455,N_16707,N_15683);
xor U21456 (N_21456,N_16697,N_15900);
nor U21457 (N_21457,N_16491,N_17993);
nand U21458 (N_21458,N_18631,N_17381);
or U21459 (N_21459,N_18455,N_18719);
nand U21460 (N_21460,N_15828,N_16920);
nand U21461 (N_21461,N_15668,N_17848);
or U21462 (N_21462,N_18719,N_17299);
and U21463 (N_21463,N_17041,N_18160);
or U21464 (N_21464,N_17509,N_16098);
nor U21465 (N_21465,N_17987,N_18118);
nand U21466 (N_21466,N_17133,N_17809);
or U21467 (N_21467,N_17695,N_18041);
xor U21468 (N_21468,N_18148,N_16728);
xor U21469 (N_21469,N_15842,N_17691);
or U21470 (N_21470,N_17138,N_16077);
nor U21471 (N_21471,N_17964,N_15722);
or U21472 (N_21472,N_16316,N_17819);
xnor U21473 (N_21473,N_17577,N_16870);
and U21474 (N_21474,N_16474,N_16698);
xor U21475 (N_21475,N_17338,N_18513);
or U21476 (N_21476,N_18021,N_17194);
nand U21477 (N_21477,N_17234,N_16426);
or U21478 (N_21478,N_18159,N_16486);
and U21479 (N_21479,N_18056,N_16248);
and U21480 (N_21480,N_18085,N_18679);
and U21481 (N_21481,N_16462,N_16774);
and U21482 (N_21482,N_17513,N_17276);
xor U21483 (N_21483,N_16492,N_17551);
nand U21484 (N_21484,N_17680,N_17859);
nand U21485 (N_21485,N_18099,N_18063);
nor U21486 (N_21486,N_16692,N_17831);
nor U21487 (N_21487,N_15816,N_17395);
nor U21488 (N_21488,N_17352,N_17652);
and U21489 (N_21489,N_17598,N_16700);
nor U21490 (N_21490,N_16162,N_16064);
or U21491 (N_21491,N_18132,N_18590);
xnor U21492 (N_21492,N_17894,N_15924);
nor U21493 (N_21493,N_18003,N_15819);
xnor U21494 (N_21494,N_17972,N_18300);
nand U21495 (N_21495,N_16140,N_17553);
nand U21496 (N_21496,N_18465,N_17550);
xnor U21497 (N_21497,N_18284,N_15721);
nor U21498 (N_21498,N_18015,N_17583);
and U21499 (N_21499,N_18744,N_16948);
nor U21500 (N_21500,N_18685,N_16132);
nor U21501 (N_21501,N_16102,N_17950);
or U21502 (N_21502,N_16643,N_16348);
and U21503 (N_21503,N_17893,N_15680);
or U21504 (N_21504,N_18073,N_18692);
xor U21505 (N_21505,N_18162,N_17793);
and U21506 (N_21506,N_18492,N_15911);
and U21507 (N_21507,N_17148,N_16112);
xor U21508 (N_21508,N_16319,N_18183);
and U21509 (N_21509,N_18511,N_16272);
nand U21510 (N_21510,N_17971,N_16814);
or U21511 (N_21511,N_16132,N_15654);
and U21512 (N_21512,N_17995,N_16362);
and U21513 (N_21513,N_15982,N_16929);
or U21514 (N_21514,N_18529,N_17349);
xor U21515 (N_21515,N_15655,N_18374);
and U21516 (N_21516,N_17124,N_17399);
and U21517 (N_21517,N_17419,N_16073);
nor U21518 (N_21518,N_18703,N_18432);
or U21519 (N_21519,N_16083,N_18032);
or U21520 (N_21520,N_15717,N_17204);
nand U21521 (N_21521,N_16259,N_15729);
nor U21522 (N_21522,N_17902,N_16616);
nor U21523 (N_21523,N_18592,N_18631);
xor U21524 (N_21524,N_16399,N_16323);
or U21525 (N_21525,N_18143,N_17625);
and U21526 (N_21526,N_17335,N_16100);
nor U21527 (N_21527,N_15843,N_15695);
xor U21528 (N_21528,N_16465,N_15787);
nor U21529 (N_21529,N_16804,N_18193);
nand U21530 (N_21530,N_17388,N_18241);
xor U21531 (N_21531,N_16555,N_18142);
or U21532 (N_21532,N_17674,N_15844);
nor U21533 (N_21533,N_17944,N_16815);
nand U21534 (N_21534,N_17960,N_16119);
nand U21535 (N_21535,N_16208,N_15879);
and U21536 (N_21536,N_17288,N_18125);
or U21537 (N_21537,N_18508,N_18660);
xnor U21538 (N_21538,N_16178,N_16745);
and U21539 (N_21539,N_16094,N_16570);
xor U21540 (N_21540,N_16659,N_17991);
xnor U21541 (N_21541,N_15888,N_16450);
and U21542 (N_21542,N_16874,N_16516);
nor U21543 (N_21543,N_16451,N_18046);
or U21544 (N_21544,N_17126,N_16297);
xor U21545 (N_21545,N_16649,N_16584);
and U21546 (N_21546,N_16640,N_16130);
or U21547 (N_21547,N_16568,N_16326);
or U21548 (N_21548,N_18469,N_16202);
nand U21549 (N_21549,N_18650,N_17450);
nor U21550 (N_21550,N_15723,N_17734);
nand U21551 (N_21551,N_17264,N_17720);
nand U21552 (N_21552,N_16706,N_15652);
nand U21553 (N_21553,N_16472,N_17326);
or U21554 (N_21554,N_16870,N_16650);
and U21555 (N_21555,N_16876,N_17760);
nand U21556 (N_21556,N_16282,N_18540);
and U21557 (N_21557,N_17912,N_15650);
or U21558 (N_21558,N_18698,N_18550);
or U21559 (N_21559,N_16656,N_15871);
nor U21560 (N_21560,N_17543,N_18614);
or U21561 (N_21561,N_18370,N_17239);
and U21562 (N_21562,N_16983,N_17737);
nor U21563 (N_21563,N_15808,N_16839);
and U21564 (N_21564,N_18514,N_17028);
nor U21565 (N_21565,N_18566,N_17075);
nor U21566 (N_21566,N_18396,N_16337);
nor U21567 (N_21567,N_15844,N_16732);
nand U21568 (N_21568,N_17037,N_17305);
xnor U21569 (N_21569,N_16361,N_16225);
and U21570 (N_21570,N_15941,N_18320);
nor U21571 (N_21571,N_18155,N_15666);
and U21572 (N_21572,N_16016,N_15907);
nor U21573 (N_21573,N_15709,N_17846);
xnor U21574 (N_21574,N_17814,N_18029);
nand U21575 (N_21575,N_17656,N_17497);
nor U21576 (N_21576,N_15940,N_17369);
xnor U21577 (N_21577,N_15772,N_17464);
and U21578 (N_21578,N_16472,N_18068);
nand U21579 (N_21579,N_17845,N_17298);
and U21580 (N_21580,N_16091,N_17283);
nor U21581 (N_21581,N_18239,N_16651);
nor U21582 (N_21582,N_17783,N_17470);
xnor U21583 (N_21583,N_17866,N_17085);
or U21584 (N_21584,N_18448,N_18646);
nand U21585 (N_21585,N_17499,N_18681);
and U21586 (N_21586,N_17405,N_15863);
xor U21587 (N_21587,N_18030,N_16997);
and U21588 (N_21588,N_16067,N_18335);
nand U21589 (N_21589,N_17202,N_18372);
nand U21590 (N_21590,N_18696,N_15785);
and U21591 (N_21591,N_16243,N_16842);
or U21592 (N_21592,N_16419,N_18268);
or U21593 (N_21593,N_15644,N_17122);
or U21594 (N_21594,N_17166,N_18207);
xnor U21595 (N_21595,N_17564,N_16901);
or U21596 (N_21596,N_17397,N_17644);
or U21597 (N_21597,N_18554,N_16895);
xor U21598 (N_21598,N_18096,N_17372);
nand U21599 (N_21599,N_17791,N_16062);
nor U21600 (N_21600,N_18392,N_16776);
or U21601 (N_21601,N_17638,N_17495);
nor U21602 (N_21602,N_17668,N_16490);
nand U21603 (N_21603,N_17522,N_18546);
nand U21604 (N_21604,N_16773,N_17654);
or U21605 (N_21605,N_17832,N_18420);
and U21606 (N_21606,N_16048,N_18375);
and U21607 (N_21607,N_18422,N_17770);
and U21608 (N_21608,N_16888,N_16318);
xnor U21609 (N_21609,N_15880,N_17581);
nand U21610 (N_21610,N_16534,N_17419);
xnor U21611 (N_21611,N_16014,N_16370);
nor U21612 (N_21612,N_16086,N_17993);
nand U21613 (N_21613,N_17479,N_17294);
xnor U21614 (N_21614,N_18123,N_16484);
nand U21615 (N_21615,N_15845,N_15718);
or U21616 (N_21616,N_17734,N_18194);
nand U21617 (N_21617,N_15940,N_17346);
xnor U21618 (N_21618,N_18341,N_18117);
nor U21619 (N_21619,N_18175,N_17406);
or U21620 (N_21620,N_18328,N_18014);
or U21621 (N_21621,N_15702,N_16715);
or U21622 (N_21622,N_15674,N_18598);
or U21623 (N_21623,N_17193,N_17191);
nor U21624 (N_21624,N_16459,N_17374);
xor U21625 (N_21625,N_16778,N_17022);
nor U21626 (N_21626,N_17529,N_17942);
nor U21627 (N_21627,N_16878,N_15800);
and U21628 (N_21628,N_17533,N_18515);
nor U21629 (N_21629,N_17601,N_15926);
nand U21630 (N_21630,N_18456,N_17222);
nor U21631 (N_21631,N_18698,N_16881);
nand U21632 (N_21632,N_16553,N_18425);
nand U21633 (N_21633,N_16017,N_16767);
and U21634 (N_21634,N_16665,N_17325);
nor U21635 (N_21635,N_18255,N_17060);
nand U21636 (N_21636,N_16328,N_18709);
or U21637 (N_21637,N_18373,N_17256);
or U21638 (N_21638,N_18278,N_15635);
nor U21639 (N_21639,N_18207,N_16354);
and U21640 (N_21640,N_18583,N_15712);
xnor U21641 (N_21641,N_17898,N_18388);
nor U21642 (N_21642,N_17088,N_17996);
nor U21643 (N_21643,N_16015,N_17258);
or U21644 (N_21644,N_15690,N_16090);
or U21645 (N_21645,N_17111,N_18713);
nor U21646 (N_21646,N_16270,N_15903);
nand U21647 (N_21647,N_17677,N_16273);
xor U21648 (N_21648,N_18453,N_16451);
nand U21649 (N_21649,N_16626,N_17709);
xnor U21650 (N_21650,N_16902,N_15950);
xor U21651 (N_21651,N_16533,N_17294);
or U21652 (N_21652,N_17073,N_18444);
xnor U21653 (N_21653,N_17120,N_15888);
nand U21654 (N_21654,N_18290,N_18443);
nor U21655 (N_21655,N_17761,N_18449);
nor U21656 (N_21656,N_16974,N_17723);
or U21657 (N_21657,N_15917,N_17040);
or U21658 (N_21658,N_15958,N_17566);
nor U21659 (N_21659,N_18072,N_16575);
xnor U21660 (N_21660,N_15989,N_16087);
xnor U21661 (N_21661,N_16013,N_18718);
nand U21662 (N_21662,N_16361,N_17341);
xor U21663 (N_21663,N_16039,N_17881);
nor U21664 (N_21664,N_17273,N_17891);
xnor U21665 (N_21665,N_16520,N_16451);
nand U21666 (N_21666,N_17786,N_17058);
nand U21667 (N_21667,N_16767,N_16825);
nand U21668 (N_21668,N_16781,N_17932);
nand U21669 (N_21669,N_16854,N_17550);
nand U21670 (N_21670,N_16514,N_15910);
nand U21671 (N_21671,N_16217,N_16553);
nor U21672 (N_21672,N_16939,N_16197);
nand U21673 (N_21673,N_15934,N_18483);
xor U21674 (N_21674,N_16459,N_17793);
nand U21675 (N_21675,N_16268,N_16761);
nand U21676 (N_21676,N_15951,N_16797);
or U21677 (N_21677,N_16917,N_16981);
and U21678 (N_21678,N_17815,N_15886);
or U21679 (N_21679,N_16617,N_18272);
and U21680 (N_21680,N_16982,N_18625);
nand U21681 (N_21681,N_15922,N_17618);
and U21682 (N_21682,N_18667,N_16106);
xnor U21683 (N_21683,N_16474,N_18007);
or U21684 (N_21684,N_16191,N_16978);
or U21685 (N_21685,N_16347,N_16607);
nor U21686 (N_21686,N_16919,N_16473);
nor U21687 (N_21687,N_18348,N_16776);
xnor U21688 (N_21688,N_17654,N_17570);
nand U21689 (N_21689,N_16223,N_15766);
nor U21690 (N_21690,N_18397,N_17201);
xor U21691 (N_21691,N_16287,N_16062);
nor U21692 (N_21692,N_16564,N_17116);
xnor U21693 (N_21693,N_16649,N_18179);
and U21694 (N_21694,N_17214,N_16259);
or U21695 (N_21695,N_16487,N_16038);
nand U21696 (N_21696,N_16428,N_18608);
nand U21697 (N_21697,N_15786,N_16770);
or U21698 (N_21698,N_17939,N_15628);
nand U21699 (N_21699,N_15764,N_16059);
or U21700 (N_21700,N_18013,N_16564);
xnor U21701 (N_21701,N_17626,N_16342);
or U21702 (N_21702,N_16431,N_15926);
nor U21703 (N_21703,N_18165,N_17988);
or U21704 (N_21704,N_16745,N_17376);
nand U21705 (N_21705,N_18095,N_16398);
nor U21706 (N_21706,N_17159,N_16841);
xor U21707 (N_21707,N_17794,N_17101);
nor U21708 (N_21708,N_16864,N_18739);
nor U21709 (N_21709,N_18470,N_18040);
xor U21710 (N_21710,N_18500,N_18228);
nor U21711 (N_21711,N_16524,N_15829);
and U21712 (N_21712,N_15889,N_15789);
nor U21713 (N_21713,N_16901,N_17250);
or U21714 (N_21714,N_17835,N_15886);
nand U21715 (N_21715,N_15828,N_15821);
nand U21716 (N_21716,N_16147,N_16519);
nand U21717 (N_21717,N_16509,N_17241);
nand U21718 (N_21718,N_18717,N_17156);
xor U21719 (N_21719,N_16601,N_17435);
or U21720 (N_21720,N_16224,N_16695);
nand U21721 (N_21721,N_17853,N_16731);
or U21722 (N_21722,N_17264,N_17235);
xor U21723 (N_21723,N_16695,N_18049);
or U21724 (N_21724,N_16370,N_17558);
nand U21725 (N_21725,N_16044,N_16659);
nand U21726 (N_21726,N_17932,N_16088);
nor U21727 (N_21727,N_15676,N_16016);
nor U21728 (N_21728,N_18095,N_18468);
or U21729 (N_21729,N_17055,N_16627);
xnor U21730 (N_21730,N_16434,N_16543);
nand U21731 (N_21731,N_16729,N_18080);
xnor U21732 (N_21732,N_17465,N_18252);
nor U21733 (N_21733,N_17144,N_15763);
nor U21734 (N_21734,N_16692,N_16685);
nor U21735 (N_21735,N_18743,N_17898);
nor U21736 (N_21736,N_17533,N_16242);
nand U21737 (N_21737,N_16812,N_15747);
nor U21738 (N_21738,N_16810,N_17424);
xnor U21739 (N_21739,N_15694,N_15771);
xor U21740 (N_21740,N_16304,N_16664);
or U21741 (N_21741,N_16454,N_18313);
nor U21742 (N_21742,N_17638,N_17794);
or U21743 (N_21743,N_17368,N_17983);
and U21744 (N_21744,N_17860,N_16278);
and U21745 (N_21745,N_18055,N_15948);
nand U21746 (N_21746,N_16841,N_18153);
xor U21747 (N_21747,N_16290,N_17226);
nand U21748 (N_21748,N_17095,N_16693);
and U21749 (N_21749,N_18629,N_16569);
xor U21750 (N_21750,N_16522,N_17869);
xor U21751 (N_21751,N_17211,N_17794);
and U21752 (N_21752,N_17417,N_18002);
and U21753 (N_21753,N_16451,N_17615);
nor U21754 (N_21754,N_16047,N_16081);
or U21755 (N_21755,N_17469,N_15929);
nand U21756 (N_21756,N_16469,N_15894);
nor U21757 (N_21757,N_15885,N_17395);
and U21758 (N_21758,N_15844,N_18281);
or U21759 (N_21759,N_16355,N_17560);
or U21760 (N_21760,N_18660,N_18021);
nor U21761 (N_21761,N_18198,N_15753);
nor U21762 (N_21762,N_16631,N_17517);
or U21763 (N_21763,N_18160,N_16785);
xnor U21764 (N_21764,N_18560,N_16641);
or U21765 (N_21765,N_16410,N_17811);
or U21766 (N_21766,N_16667,N_16072);
nor U21767 (N_21767,N_16328,N_17558);
nor U21768 (N_21768,N_17480,N_18380);
or U21769 (N_21769,N_18322,N_15885);
nor U21770 (N_21770,N_17367,N_18561);
or U21771 (N_21771,N_17695,N_15729);
or U21772 (N_21772,N_16786,N_17486);
nor U21773 (N_21773,N_16594,N_17270);
and U21774 (N_21774,N_16971,N_16443);
nor U21775 (N_21775,N_16834,N_17438);
nand U21776 (N_21776,N_17060,N_15940);
or U21777 (N_21777,N_16664,N_17611);
and U21778 (N_21778,N_16498,N_17284);
or U21779 (N_21779,N_16264,N_18150);
xor U21780 (N_21780,N_16498,N_17896);
or U21781 (N_21781,N_16947,N_16585);
xor U21782 (N_21782,N_17908,N_18349);
xor U21783 (N_21783,N_16503,N_16574);
xor U21784 (N_21784,N_16942,N_16931);
or U21785 (N_21785,N_17573,N_18409);
or U21786 (N_21786,N_17792,N_18256);
xnor U21787 (N_21787,N_16023,N_17449);
nor U21788 (N_21788,N_16897,N_16044);
nor U21789 (N_21789,N_18618,N_15765);
nand U21790 (N_21790,N_17983,N_18433);
or U21791 (N_21791,N_17917,N_16166);
or U21792 (N_21792,N_16039,N_17558);
and U21793 (N_21793,N_18171,N_15859);
or U21794 (N_21794,N_17586,N_16582);
and U21795 (N_21795,N_18465,N_18062);
nor U21796 (N_21796,N_18155,N_18393);
nand U21797 (N_21797,N_16210,N_16529);
and U21798 (N_21798,N_18642,N_16160);
xnor U21799 (N_21799,N_16884,N_16323);
or U21800 (N_21800,N_17456,N_16489);
nand U21801 (N_21801,N_16732,N_17223);
or U21802 (N_21802,N_17294,N_17206);
or U21803 (N_21803,N_17406,N_18660);
nand U21804 (N_21804,N_15654,N_17112);
xnor U21805 (N_21805,N_16577,N_17005);
xnor U21806 (N_21806,N_17026,N_18704);
nor U21807 (N_21807,N_17527,N_17228);
or U21808 (N_21808,N_18612,N_15643);
or U21809 (N_21809,N_16780,N_16168);
xor U21810 (N_21810,N_17086,N_15928);
and U21811 (N_21811,N_17571,N_17453);
xnor U21812 (N_21812,N_17083,N_18530);
nand U21813 (N_21813,N_17258,N_15655);
or U21814 (N_21814,N_18676,N_17662);
or U21815 (N_21815,N_16837,N_16142);
nor U21816 (N_21816,N_18006,N_17487);
or U21817 (N_21817,N_17390,N_18062);
xor U21818 (N_21818,N_15637,N_16890);
nor U21819 (N_21819,N_17330,N_17242);
xor U21820 (N_21820,N_17975,N_16409);
xnor U21821 (N_21821,N_18262,N_16113);
nand U21822 (N_21822,N_16738,N_18111);
and U21823 (N_21823,N_17871,N_16990);
and U21824 (N_21824,N_18379,N_16365);
and U21825 (N_21825,N_15652,N_17109);
nor U21826 (N_21826,N_16737,N_16699);
nor U21827 (N_21827,N_18291,N_16783);
nor U21828 (N_21828,N_16869,N_17049);
xor U21829 (N_21829,N_18140,N_17008);
xnor U21830 (N_21830,N_15774,N_15648);
or U21831 (N_21831,N_17811,N_16074);
nor U21832 (N_21832,N_18529,N_17513);
and U21833 (N_21833,N_15750,N_15979);
nand U21834 (N_21834,N_16001,N_16132);
or U21835 (N_21835,N_15692,N_15679);
nand U21836 (N_21836,N_18318,N_17335);
and U21837 (N_21837,N_16756,N_15905);
nand U21838 (N_21838,N_15733,N_17551);
or U21839 (N_21839,N_18100,N_16602);
xor U21840 (N_21840,N_16565,N_16988);
and U21841 (N_21841,N_16250,N_18698);
nor U21842 (N_21842,N_16837,N_16406);
nor U21843 (N_21843,N_16255,N_17336);
nand U21844 (N_21844,N_17134,N_16224);
xnor U21845 (N_21845,N_16022,N_18289);
or U21846 (N_21846,N_17583,N_17935);
and U21847 (N_21847,N_18710,N_17785);
or U21848 (N_21848,N_16135,N_18319);
or U21849 (N_21849,N_15852,N_16411);
nor U21850 (N_21850,N_18024,N_16735);
nor U21851 (N_21851,N_16776,N_16289);
nand U21852 (N_21852,N_17357,N_16874);
or U21853 (N_21853,N_16625,N_17437);
nand U21854 (N_21854,N_17465,N_18208);
nand U21855 (N_21855,N_16329,N_17433);
nor U21856 (N_21856,N_18285,N_18184);
xnor U21857 (N_21857,N_16833,N_18280);
nor U21858 (N_21858,N_16198,N_15661);
or U21859 (N_21859,N_16706,N_18632);
or U21860 (N_21860,N_17959,N_17465);
nor U21861 (N_21861,N_16606,N_16058);
xnor U21862 (N_21862,N_16576,N_18211);
nor U21863 (N_21863,N_15984,N_17982);
or U21864 (N_21864,N_18107,N_17510);
xnor U21865 (N_21865,N_17120,N_18625);
xor U21866 (N_21866,N_18416,N_17590);
nand U21867 (N_21867,N_17924,N_18036);
and U21868 (N_21868,N_17679,N_16744);
nor U21869 (N_21869,N_17509,N_18202);
or U21870 (N_21870,N_18450,N_18688);
nand U21871 (N_21871,N_18564,N_16574);
or U21872 (N_21872,N_17138,N_17958);
xnor U21873 (N_21873,N_16585,N_18410);
nand U21874 (N_21874,N_18663,N_18112);
xnor U21875 (N_21875,N_19216,N_19566);
xnor U21876 (N_21876,N_21282,N_18863);
or U21877 (N_21877,N_20962,N_19679);
nor U21878 (N_21878,N_18912,N_19045);
and U21879 (N_21879,N_20954,N_21622);
or U21880 (N_21880,N_21199,N_19726);
and U21881 (N_21881,N_19415,N_21113);
nand U21882 (N_21882,N_19212,N_20926);
and U21883 (N_21883,N_21515,N_21647);
or U21884 (N_21884,N_21830,N_20566);
or U21885 (N_21885,N_20121,N_19981);
xnor U21886 (N_21886,N_19673,N_19464);
nor U21887 (N_21887,N_20354,N_20271);
xor U21888 (N_21888,N_21538,N_20757);
xor U21889 (N_21889,N_20139,N_21833);
nor U21890 (N_21890,N_20716,N_19780);
and U21891 (N_21891,N_21344,N_21564);
nor U21892 (N_21892,N_19739,N_21391);
nand U21893 (N_21893,N_19043,N_19366);
nand U21894 (N_21894,N_21131,N_20594);
or U21895 (N_21895,N_21571,N_20624);
xnor U21896 (N_21896,N_19141,N_20610);
nand U21897 (N_21897,N_19837,N_20433);
xor U21898 (N_21898,N_19922,N_20071);
or U21899 (N_21899,N_20491,N_20927);
nor U21900 (N_21900,N_19071,N_19625);
nand U21901 (N_21901,N_21652,N_20074);
nor U21902 (N_21902,N_20058,N_19823);
or U21903 (N_21903,N_19219,N_19574);
nand U21904 (N_21904,N_19569,N_18821);
nor U21905 (N_21905,N_21419,N_18916);
or U21906 (N_21906,N_20778,N_18816);
nor U21907 (N_21907,N_18802,N_19921);
nor U21908 (N_21908,N_20356,N_19988);
and U21909 (N_21909,N_19746,N_19388);
xnor U21910 (N_21910,N_20189,N_20267);
nand U21911 (N_21911,N_19320,N_19352);
nor U21912 (N_21912,N_20478,N_21811);
nor U21913 (N_21913,N_20761,N_21856);
nand U21914 (N_21914,N_19952,N_19736);
nor U21915 (N_21915,N_19041,N_21291);
xnor U21916 (N_21916,N_19236,N_20222);
or U21917 (N_21917,N_19325,N_21508);
and U21918 (N_21918,N_20575,N_19314);
or U21919 (N_21919,N_21500,N_21542);
or U21920 (N_21920,N_20389,N_19166);
nand U21921 (N_21921,N_20515,N_19289);
nor U21922 (N_21922,N_20488,N_19640);
nor U21923 (N_21923,N_19884,N_19067);
and U21924 (N_21924,N_21706,N_21260);
xnor U21925 (N_21925,N_21699,N_19716);
or U21926 (N_21926,N_20273,N_18873);
nand U21927 (N_21927,N_21171,N_19046);
and U21928 (N_21928,N_21208,N_18791);
or U21929 (N_21929,N_20542,N_19515);
or U21930 (N_21930,N_19907,N_20143);
and U21931 (N_21931,N_19160,N_20547);
nand U21932 (N_21932,N_21488,N_21196);
or U21933 (N_21933,N_21049,N_19529);
and U21934 (N_21934,N_20257,N_21740);
xnor U21935 (N_21935,N_20947,N_20873);
and U21936 (N_21936,N_21099,N_19465);
xnor U21937 (N_21937,N_19315,N_18985);
or U21938 (N_21938,N_21270,N_20439);
nand U21939 (N_21939,N_19117,N_20153);
nor U21940 (N_21940,N_21016,N_18855);
nand U21941 (N_21941,N_20655,N_20069);
and U21942 (N_21942,N_19942,N_21690);
xnor U21943 (N_21943,N_21333,N_21286);
nor U21944 (N_21944,N_18877,N_19389);
nand U21945 (N_21945,N_20412,N_21470);
or U21946 (N_21946,N_20463,N_20764);
nand U21947 (N_21947,N_20514,N_19001);
nand U21948 (N_21948,N_20998,N_20252);
nor U21949 (N_21949,N_19963,N_19980);
nand U21950 (N_21950,N_19728,N_20559);
or U21951 (N_21951,N_19663,N_20205);
nand U21952 (N_21952,N_21594,N_19594);
nand U21953 (N_21953,N_20835,N_20538);
or U21954 (N_21954,N_21871,N_19107);
or U21955 (N_21955,N_20051,N_21212);
xnor U21956 (N_21956,N_19124,N_20743);
or U21957 (N_21957,N_21549,N_20268);
and U21958 (N_21958,N_20017,N_21834);
nand U21959 (N_21959,N_21028,N_19047);
nor U21960 (N_21960,N_21007,N_21437);
or U21961 (N_21961,N_20129,N_20206);
and U21962 (N_21962,N_18799,N_21070);
or U21963 (N_21963,N_20936,N_20219);
xnor U21964 (N_21964,N_21742,N_19627);
xor U21965 (N_21965,N_19915,N_19059);
nor U21966 (N_21966,N_20528,N_21772);
nor U21967 (N_21967,N_20746,N_20572);
nand U21968 (N_21968,N_20885,N_19609);
nor U21969 (N_21969,N_19240,N_19493);
nor U21970 (N_21970,N_19062,N_19345);
nand U21971 (N_21971,N_21785,N_18935);
nor U21972 (N_21972,N_18865,N_20940);
and U21973 (N_21973,N_21472,N_20719);
or U21974 (N_21974,N_19094,N_19018);
nor U21975 (N_21975,N_21719,N_20907);
xnor U21976 (N_21976,N_21205,N_19154);
xnor U21977 (N_21977,N_18758,N_20086);
xnor U21978 (N_21978,N_19879,N_21401);
or U21979 (N_21979,N_20803,N_19403);
and U21980 (N_21980,N_21275,N_20380);
nor U21981 (N_21981,N_20003,N_19731);
and U21982 (N_21982,N_19308,N_21844);
nor U21983 (N_21983,N_20630,N_18807);
nor U21984 (N_21984,N_21012,N_19063);
or U21985 (N_21985,N_19483,N_20314);
or U21986 (N_21986,N_19409,N_19135);
and U21987 (N_21987,N_18796,N_18870);
xnor U21988 (N_21988,N_19101,N_19858);
and U21989 (N_21989,N_19319,N_21490);
xor U21990 (N_21990,N_20519,N_20929);
or U21991 (N_21991,N_20866,N_20647);
xnor U21992 (N_21992,N_20820,N_19178);
or U21993 (N_21993,N_21821,N_20427);
and U21994 (N_21994,N_19777,N_21238);
xnor U21995 (N_21995,N_21239,N_21584);
and U21996 (N_21996,N_21707,N_21119);
nand U21997 (N_21997,N_21602,N_20571);
nand U21998 (N_21998,N_19576,N_20725);
and U21999 (N_21999,N_19191,N_20009);
and U22000 (N_22000,N_19603,N_18993);
or U22001 (N_22001,N_19984,N_19859);
or U22002 (N_22002,N_20472,N_20251);
xnor U22003 (N_22003,N_21025,N_19740);
nand U22004 (N_22004,N_19022,N_19185);
and U22005 (N_22005,N_21739,N_20775);
or U22006 (N_22006,N_20373,N_19770);
nor U22007 (N_22007,N_20669,N_20179);
and U22008 (N_22008,N_19601,N_18771);
xor U22009 (N_22009,N_21780,N_20800);
nand U22010 (N_22010,N_19499,N_19204);
and U22011 (N_22011,N_19037,N_18806);
nand U22012 (N_22012,N_20544,N_21400);
nor U22013 (N_22013,N_21759,N_19343);
and U22014 (N_22014,N_20371,N_19151);
nand U22015 (N_22015,N_20768,N_20502);
nand U22016 (N_22016,N_21777,N_20963);
xnor U22017 (N_22017,N_20474,N_19749);
nor U22018 (N_22018,N_21676,N_21279);
nand U22019 (N_22019,N_19072,N_21321);
and U22020 (N_22020,N_21573,N_19996);
and U22021 (N_22021,N_19668,N_20014);
nor U22022 (N_22022,N_20619,N_20946);
nand U22023 (N_22023,N_20924,N_19639);
xor U22024 (N_22024,N_19895,N_19148);
or U22025 (N_22025,N_19145,N_21559);
or U22026 (N_22026,N_18756,N_18983);
nand U22027 (N_22027,N_19467,N_20638);
nor U22028 (N_22028,N_21442,N_21632);
or U22029 (N_22029,N_18876,N_21200);
nor U22030 (N_22030,N_21411,N_21203);
xnor U22031 (N_22031,N_19501,N_20229);
xnor U22032 (N_22032,N_19055,N_19142);
and U22033 (N_22033,N_19847,N_21445);
and U22034 (N_22034,N_20168,N_20413);
nor U22035 (N_22035,N_21367,N_19964);
or U22036 (N_22036,N_20847,N_19687);
xor U22037 (N_22037,N_20365,N_20902);
xnor U22038 (N_22038,N_19841,N_21713);
nor U22039 (N_22039,N_19634,N_20088);
and U22040 (N_22040,N_20280,N_19196);
nor U22041 (N_22041,N_20277,N_18891);
nand U22042 (N_22042,N_19158,N_21518);
xor U22043 (N_22043,N_21336,N_20243);
nor U22044 (N_22044,N_21292,N_21217);
and U22045 (N_22045,N_19238,N_21737);
and U22046 (N_22046,N_20374,N_20712);
and U22047 (N_22047,N_21655,N_19233);
nor U22048 (N_22048,N_18990,N_19844);
xnor U22049 (N_22049,N_20912,N_20334);
nand U22050 (N_22050,N_19245,N_19187);
nand U22051 (N_22051,N_18857,N_21278);
nand U22052 (N_22052,N_20173,N_20298);
nand U22053 (N_22053,N_21497,N_19069);
nor U22054 (N_22054,N_21779,N_19371);
nor U22055 (N_22055,N_19809,N_20990);
or U22056 (N_22056,N_21263,N_20584);
nor U22057 (N_22057,N_21194,N_20601);
nor U22058 (N_22058,N_21646,N_19806);
and U22059 (N_22059,N_20355,N_21600);
nand U22060 (N_22060,N_20932,N_19544);
xnor U22061 (N_22061,N_20958,N_20819);
and U22062 (N_22062,N_19163,N_21000);
nor U22063 (N_22063,N_21589,N_21305);
and U22064 (N_22064,N_19478,N_21587);
and U22065 (N_22065,N_20221,N_21798);
nand U22066 (N_22066,N_20417,N_19674);
and U22067 (N_22067,N_19316,N_19845);
nor U22068 (N_22068,N_20451,N_21373);
nand U22069 (N_22069,N_19102,N_18764);
xnor U22070 (N_22070,N_19384,N_19336);
or U22071 (N_22071,N_18977,N_19267);
nand U22072 (N_22072,N_21349,N_20604);
and U22073 (N_22073,N_20013,N_20392);
xor U22074 (N_22074,N_21688,N_19195);
nor U22075 (N_22075,N_20732,N_20312);
nor U22076 (N_22076,N_21628,N_19270);
or U22077 (N_22077,N_19798,N_21671);
xnor U22078 (N_22078,N_19350,N_19425);
or U22079 (N_22079,N_18963,N_19558);
and U22080 (N_22080,N_20193,N_21020);
xor U22081 (N_22081,N_20649,N_21698);
xnor U22082 (N_22082,N_20149,N_19870);
nor U22083 (N_22083,N_19608,N_20957);
nand U22084 (N_22084,N_20241,N_19817);
or U22085 (N_22085,N_20369,N_19993);
nor U22086 (N_22086,N_21635,N_21603);
nor U22087 (N_22087,N_19591,N_21301);
nand U22088 (N_22088,N_19220,N_18842);
nor U22089 (N_22089,N_20539,N_18782);
nor U22090 (N_22090,N_21145,N_21796);
xor U22091 (N_22091,N_19431,N_19500);
xnor U22092 (N_22092,N_21519,N_21074);
nor U22093 (N_22093,N_21439,N_21177);
nand U22094 (N_22094,N_20207,N_19623);
nor U22095 (N_22095,N_19581,N_20771);
nand U22096 (N_22096,N_19539,N_19670);
or U22097 (N_22097,N_20675,N_20614);
and U22098 (N_22098,N_21694,N_20201);
nor U22099 (N_22099,N_20437,N_21862);
or U22100 (N_22100,N_19508,N_19034);
nand U22101 (N_22101,N_18976,N_20845);
xnor U22102 (N_22102,N_19919,N_20471);
xor U22103 (N_22103,N_18770,N_20747);
nor U22104 (N_22104,N_20879,N_19134);
or U22105 (N_22105,N_18903,N_21040);
xor U22106 (N_22106,N_18918,N_20860);
xnor U22107 (N_22107,N_21226,N_21232);
and U22108 (N_22108,N_20646,N_21861);
and U22109 (N_22109,N_21431,N_19053);
nor U22110 (N_22110,N_21393,N_19546);
nor U22111 (N_22111,N_20813,N_20418);
nor U22112 (N_22112,N_20939,N_20052);
nand U22113 (N_22113,N_18930,N_20165);
nand U22114 (N_22114,N_21110,N_21410);
nor U22115 (N_22115,N_20075,N_18905);
xnor U22116 (N_22116,N_20503,N_21197);
or U22117 (N_22117,N_21744,N_21316);
nand U22118 (N_22118,N_19871,N_20342);
and U22119 (N_22119,N_21745,N_19560);
nand U22120 (N_22120,N_20760,N_20245);
nand U22121 (N_22121,N_20598,N_20070);
nor U22122 (N_22122,N_19104,N_20037);
xnor U22123 (N_22123,N_18845,N_21634);
or U22124 (N_22124,N_19433,N_21734);
nand U22125 (N_22125,N_20315,N_18944);
nor U22126 (N_22126,N_18755,N_21293);
nand U22127 (N_22127,N_21329,N_19678);
nand U22128 (N_22128,N_19970,N_21753);
nor U22129 (N_22129,N_21342,N_21433);
nor U22130 (N_22130,N_19265,N_21181);
nor U22131 (N_22131,N_19450,N_21152);
nor U22132 (N_22132,N_19792,N_20394);
nor U22133 (N_22133,N_20323,N_20825);
xor U22134 (N_22134,N_20035,N_18933);
and U22135 (N_22135,N_21254,N_20034);
xor U22136 (N_22136,N_19712,N_20111);
nand U22137 (N_22137,N_21331,N_19435);
xnor U22138 (N_22138,N_19900,N_21266);
nand U22139 (N_22139,N_18826,N_19635);
or U22140 (N_22140,N_21845,N_20333);
xnor U22141 (N_22141,N_19867,N_20589);
nor U22142 (N_22142,N_21044,N_20870);
nand U22143 (N_22143,N_21610,N_20203);
xnor U22144 (N_22144,N_19190,N_21220);
nor U22145 (N_22145,N_20641,N_20414);
nand U22146 (N_22146,N_19054,N_19451);
nand U22147 (N_22147,N_19514,N_20979);
nand U22148 (N_22148,N_20170,N_18934);
xnor U22149 (N_22149,N_20863,N_19972);
xnor U22150 (N_22150,N_19857,N_19751);
and U22151 (N_22151,N_18982,N_20386);
or U22152 (N_22152,N_20152,N_19214);
nor U22153 (N_22153,N_21755,N_21193);
xor U22154 (N_22154,N_19274,N_21397);
nand U22155 (N_22155,N_19688,N_18810);
or U22156 (N_22156,N_20041,N_21369);
xor U22157 (N_22157,N_19311,N_21683);
xor U22158 (N_22158,N_18894,N_20824);
and U22159 (N_22159,N_20233,N_21824);
nand U22160 (N_22160,N_19019,N_20454);
nor U22161 (N_22161,N_20192,N_21158);
or U22162 (N_22162,N_19693,N_20754);
or U22163 (N_22163,N_19702,N_19013);
or U22164 (N_22164,N_19264,N_20969);
xnor U22165 (N_22165,N_18953,N_21453);
nand U22166 (N_22166,N_21122,N_19360);
xor U22167 (N_22167,N_20795,N_19482);
or U22168 (N_22168,N_19305,N_19642);
or U22169 (N_22169,N_21170,N_20468);
nor U22170 (N_22170,N_19424,N_20141);
or U22171 (N_22171,N_19012,N_21489);
xor U22172 (N_22172,N_19174,N_19288);
and U22173 (N_22173,N_20130,N_18812);
and U22174 (N_22174,N_20884,N_18937);
or U22175 (N_22175,N_20449,N_21024);
nor U22176 (N_22176,N_19694,N_20238);
or U22177 (N_22177,N_20617,N_21823);
and U22178 (N_22178,N_21661,N_19354);
and U22179 (N_22179,N_20328,N_19027);
nand U22180 (N_22180,N_18869,N_20551);
xnor U22181 (N_22181,N_19571,N_20923);
nor U22182 (N_22182,N_21700,N_21831);
nand U22183 (N_22183,N_19815,N_19498);
or U22184 (N_22184,N_21054,N_21138);
and U22185 (N_22185,N_18835,N_20805);
nand U22186 (N_22186,N_20164,N_20626);
xor U22187 (N_22187,N_21556,N_19804);
xor U22188 (N_22188,N_19734,N_20767);
and U22189 (N_22189,N_19772,N_20574);
nor U22190 (N_22190,N_20781,N_19813);
and U22191 (N_22191,N_19721,N_19894);
and U22192 (N_22192,N_21109,N_20769);
and U22193 (N_22193,N_21667,N_19452);
or U22194 (N_22194,N_20260,N_19058);
and U22195 (N_22195,N_21580,N_21059);
nand U22196 (N_22196,N_19920,N_20270);
xor U22197 (N_22197,N_19525,N_19421);
nor U22198 (N_22198,N_21364,N_20263);
xnor U22199 (N_22199,N_21817,N_20253);
nand U22200 (N_22200,N_20115,N_20255);
or U22201 (N_22201,N_18988,N_21402);
or U22202 (N_22202,N_18750,N_20210);
nor U22203 (N_22203,N_19567,N_20853);
and U22204 (N_22204,N_21385,N_20426);
nand U22205 (N_22205,N_21427,N_19754);
xnor U22206 (N_22206,N_21674,N_19259);
xnor U22207 (N_22207,N_19292,N_19899);
or U22208 (N_22208,N_19524,N_21814);
nor U22209 (N_22209,N_19032,N_20529);
or U22210 (N_22210,N_18932,N_18851);
nor U22211 (N_22211,N_18753,N_20218);
nor U22212 (N_22212,N_21539,N_18781);
or U22213 (N_22213,N_19275,N_19437);
nand U22214 (N_22214,N_19936,N_21793);
or U22215 (N_22215,N_19671,N_20855);
nand U22216 (N_22216,N_19923,N_19955);
or U22217 (N_22217,N_20387,N_21607);
and U22218 (N_22218,N_18936,N_19494);
xnor U22219 (N_22219,N_19630,N_19973);
nand U22220 (N_22220,N_18777,N_20920);
and U22221 (N_22221,N_18757,N_19946);
nand U22222 (N_22222,N_21042,N_20516);
or U22223 (N_22223,N_20444,N_20448);
or U22224 (N_22224,N_21481,N_21459);
nor U22225 (N_22225,N_21355,N_19210);
nor U22226 (N_22226,N_21487,N_18954);
nor U22227 (N_22227,N_21710,N_20684);
nand U22228 (N_22228,N_19375,N_19050);
nor U22229 (N_22229,N_20609,N_18965);
nor U22230 (N_22230,N_21368,N_21009);
nor U22231 (N_22231,N_19913,N_19161);
or U22232 (N_22232,N_18754,N_21495);
nor U22233 (N_22233,N_20364,N_21416);
xor U22234 (N_22234,N_19802,N_21289);
and U22235 (N_22235,N_18880,N_19006);
and U22236 (N_22236,N_21435,N_19522);
or U22237 (N_22237,N_18895,N_19788);
and U22238 (N_22238,N_20868,N_18949);
and U22239 (N_22239,N_20020,N_21560);
and U22240 (N_22240,N_20687,N_20275);
xnor U22241 (N_22241,N_19617,N_19249);
nor U22242 (N_22242,N_19816,N_19468);
nand U22243 (N_22243,N_19048,N_21383);
and U22244 (N_22244,N_20317,N_19790);
and U22245 (N_22245,N_21822,N_21529);
nand U22246 (N_22246,N_19486,N_20066);
xor U22247 (N_22247,N_19561,N_20916);
nor U22248 (N_22248,N_20410,N_20223);
and U22249 (N_22249,N_21339,N_20643);
or U22250 (N_22250,N_19434,N_21684);
nor U22251 (N_22251,N_20423,N_20016);
nand U22252 (N_22252,N_20332,N_20787);
xnor U22253 (N_22253,N_19370,N_19448);
nor U22254 (N_22254,N_19897,N_19604);
or U22255 (N_22255,N_19974,N_21229);
nor U22256 (N_22256,N_19248,N_20289);
nor U22257 (N_22257,N_20612,N_21849);
nor U22258 (N_22258,N_19593,N_21108);
or U22259 (N_22259,N_20329,N_18801);
and U22260 (N_22260,N_21031,N_19812);
xor U22261 (N_22261,N_20050,N_18979);
xnor U22262 (N_22262,N_19654,N_21079);
and U22263 (N_22263,N_20082,N_19438);
xnor U22264 (N_22264,N_20385,N_19155);
nor U22265 (N_22265,N_20438,N_19898);
and U22266 (N_22266,N_21456,N_20980);
nand U22267 (N_22267,N_20199,N_18763);
and U22268 (N_22268,N_20567,N_19700);
xor U22269 (N_22269,N_20330,N_19461);
or U22270 (N_22270,N_18822,N_19906);
or U22271 (N_22271,N_21124,N_21511);
or U22272 (N_22272,N_19750,N_19224);
xnor U22273 (N_22273,N_19436,N_20948);
nor U22274 (N_22274,N_20690,N_19170);
xor U22275 (N_22275,N_21738,N_21327);
nand U22276 (N_22276,N_20276,N_19727);
nand U22277 (N_22277,N_20806,N_20299);
xor U22278 (N_22278,N_19179,N_19977);
or U22279 (N_22279,N_20228,N_19268);
or U22280 (N_22280,N_19401,N_20106);
or U22281 (N_22281,N_20319,N_20042);
nand U22282 (N_22282,N_19310,N_20024);
and U22283 (N_22283,N_20893,N_20350);
and U22284 (N_22284,N_19116,N_21866);
xor U22285 (N_22285,N_19570,N_21747);
and U22286 (N_22286,N_19535,N_19648);
xor U22287 (N_22287,N_21143,N_20309);
nor U22288 (N_22288,N_21680,N_19171);
or U22289 (N_22289,N_18760,N_18911);
nor U22290 (N_22290,N_20019,N_19412);
nor U22291 (N_22291,N_21251,N_19020);
and U22292 (N_22292,N_21283,N_18886);
nor U22293 (N_22293,N_18960,N_20959);
xnor U22294 (N_22294,N_19291,N_20000);
nand U22295 (N_22295,N_19819,N_20895);
and U22296 (N_22296,N_20933,N_18774);
nand U22297 (N_22297,N_19290,N_19175);
nor U22298 (N_22298,N_20404,N_20673);
nor U22299 (N_22299,N_20955,N_19986);
xor U22300 (N_22300,N_19380,N_21526);
and U22301 (N_22301,N_19787,N_20739);
nand U22302 (N_22302,N_19659,N_19105);
xor U22303 (N_22303,N_20021,N_21868);
nand U22304 (N_22304,N_20942,N_20125);
or U22305 (N_22305,N_21754,N_19263);
and U22306 (N_22306,N_21653,N_20466);
xnor U22307 (N_22307,N_21835,N_19198);
nor U22308 (N_22308,N_21644,N_21081);
nor U22309 (N_22309,N_20759,N_18980);
nor U22310 (N_22310,N_20496,N_20520);
xnor U22311 (N_22311,N_19606,N_21725);
nor U22312 (N_22312,N_19579,N_21235);
nand U22313 (N_22313,N_21287,N_21248);
xnor U22314 (N_22314,N_21127,N_19710);
xnor U22315 (N_22315,N_21187,N_19945);
nor U22316 (N_22316,N_19666,N_19507);
or U22317 (N_22317,N_20662,N_21163);
nor U22318 (N_22318,N_19838,N_21702);
nand U22319 (N_22319,N_19280,N_20118);
or U22320 (N_22320,N_19793,N_19033);
or U22321 (N_22321,N_20737,N_21156);
nand U22322 (N_22322,N_19475,N_19949);
and U22323 (N_22323,N_20892,N_19960);
xor U22324 (N_22324,N_19797,N_20945);
nand U22325 (N_22325,N_20861,N_21061);
xor U22326 (N_22326,N_20841,N_20660);
xor U22327 (N_22327,N_20313,N_20772);
or U22328 (N_22328,N_19778,N_21265);
nor U22329 (N_22329,N_20110,N_19615);
nand U22330 (N_22330,N_20415,N_20858);
nand U22331 (N_22331,N_20079,N_21444);
nand U22332 (N_22332,N_21568,N_19090);
nor U22333 (N_22333,N_20240,N_21210);
nand U22334 (N_22334,N_18991,N_18800);
xnor U22335 (N_22335,N_20654,N_21717);
or U22336 (N_22336,N_20212,N_21065);
xnor U22337 (N_22337,N_19260,N_21429);
nor U22338 (N_22338,N_19626,N_21673);
nand U22339 (N_22339,N_20992,N_21636);
and U22340 (N_22340,N_20005,N_19304);
and U22341 (N_22341,N_20475,N_20247);
nor U22342 (N_22342,N_21829,N_20080);
or U22343 (N_22343,N_21575,N_20310);
nand U22344 (N_22344,N_19633,N_21466);
or U22345 (N_22345,N_21298,N_19492);
or U22346 (N_22346,N_20367,N_19562);
or U22347 (N_22347,N_21478,N_21514);
nor U22348 (N_22348,N_21151,N_20621);
xor U22349 (N_22349,N_19825,N_19927);
or U22350 (N_22350,N_18843,N_19829);
or U22351 (N_22351,N_19976,N_18833);
nor U22352 (N_22352,N_20906,N_19495);
or U22353 (N_22353,N_21851,N_20311);
xnor U22354 (N_22354,N_19785,N_21469);
xor U22355 (N_22355,N_20015,N_21407);
nand U22356 (N_22356,N_20499,N_19767);
and U22357 (N_22357,N_20642,N_21102);
and U22358 (N_22358,N_21018,N_21338);
nand U22359 (N_22359,N_20620,N_20636);
and U22360 (N_22360,N_21352,N_19121);
or U22361 (N_22361,N_21148,N_21045);
nor U22362 (N_22362,N_19332,N_20065);
nor U22363 (N_22363,N_21775,N_20441);
nand U22364 (N_22364,N_20838,N_20135);
xnor U22365 (N_22365,N_20482,N_21859);
or U22366 (N_22366,N_21548,N_21379);
xnor U22367 (N_22367,N_20994,N_21084);
and U22368 (N_22368,N_20096,N_21638);
nor U22369 (N_22369,N_21366,N_19965);
and U22370 (N_22370,N_19097,N_19850);
or U22371 (N_22371,N_20047,N_20811);
nand U22372 (N_22372,N_21479,N_18943);
or U22373 (N_22373,N_20556,N_21166);
and U22374 (N_22374,N_20961,N_19223);
nor U22375 (N_22375,N_18967,N_19250);
and U22376 (N_22376,N_19177,N_20843);
and U22377 (N_22377,N_21358,N_18910);
nand U22378 (N_22378,N_18776,N_19197);
xor U22379 (N_22379,N_20379,N_21064);
and U22380 (N_22380,N_19297,N_18808);
xnor U22381 (N_22381,N_20549,N_19085);
nor U22382 (N_22382,N_19725,N_19730);
xnor U22383 (N_22383,N_21236,N_21233);
or U22384 (N_22384,N_19645,N_18892);
nand U22385 (N_22385,N_21356,N_20986);
and U22386 (N_22386,N_21693,N_20985);
or U22387 (N_22387,N_20430,N_20928);
nor U22388 (N_22388,N_20765,N_20291);
nand U22389 (N_22389,N_21408,N_20450);
and U22390 (N_22390,N_21565,N_21211);
nand U22391 (N_22391,N_20789,N_18958);
or U22392 (N_22392,N_21800,N_21718);
nand U22393 (N_22393,N_21593,N_19362);
nand U22394 (N_22394,N_20736,N_19660);
nor U22395 (N_22395,N_19327,N_20909);
nor U22396 (N_22396,N_20938,N_20629);
nand U22397 (N_22397,N_19672,N_20977);
nor U22398 (N_22398,N_20644,N_20718);
nor U22399 (N_22399,N_20160,N_19079);
xor U22400 (N_22400,N_19519,N_21313);
and U22401 (N_22401,N_19680,N_19779);
or U22402 (N_22402,N_21731,N_20651);
and U22403 (N_22403,N_19381,N_19100);
or U22404 (N_22404,N_19575,N_19622);
and U22405 (N_22405,N_21395,N_20631);
nand U22406 (N_22406,N_21643,N_21801);
nand U22407 (N_22407,N_21389,N_21010);
and U22408 (N_22408,N_19686,N_19651);
xnor U22409 (N_22409,N_19376,N_20431);
or U22410 (N_22410,N_20882,N_21206);
or U22411 (N_22411,N_20810,N_20479);
or U22412 (N_22412,N_21290,N_20406);
nand U22413 (N_22413,N_19641,N_19244);
and U22414 (N_22414,N_19657,N_19554);
and U22415 (N_22415,N_20831,N_20132);
nand U22416 (N_22416,N_21786,N_19821);
xor U22417 (N_22417,N_20011,N_20522);
and U22418 (N_22418,N_19302,N_20151);
xor U22419 (N_22419,N_18875,N_20473);
xor U22420 (N_22420,N_20973,N_20461);
nor U22421 (N_22421,N_20349,N_20623);
or U22422 (N_22422,N_20187,N_20181);
nor U22423 (N_22423,N_20557,N_19966);
xor U22424 (N_22424,N_19848,N_21847);
and U22425 (N_22425,N_20236,N_20563);
nand U22426 (N_22426,N_20258,N_20854);
nor U22427 (N_22427,N_21629,N_20045);
xor U22428 (N_22428,N_21051,N_20634);
nor U22429 (N_22429,N_19232,N_20511);
or U22430 (N_22430,N_21172,N_21726);
nor U22431 (N_22431,N_20846,N_21097);
nand U22432 (N_22432,N_19192,N_19768);
nand U22433 (N_22433,N_21001,N_18817);
nand U22434 (N_22434,N_21300,N_19056);
nand U22435 (N_22435,N_20670,N_19378);
xnor U22436 (N_22436,N_19368,N_19318);
or U22437 (N_22437,N_20733,N_20057);
or U22438 (N_22438,N_20184,N_21190);
nor U22439 (N_22439,N_19115,N_21136);
or U22440 (N_22440,N_20676,N_21813);
nor U22441 (N_22441,N_20512,N_18917);
and U22442 (N_22442,N_20320,N_20568);
or U22443 (N_22443,N_21249,N_21522);
xnor U22444 (N_22444,N_21612,N_21311);
xnor U22445 (N_22445,N_20600,N_21089);
nor U22446 (N_22446,N_19647,N_21381);
xnor U22447 (N_22447,N_20147,N_21658);
xor U22448 (N_22448,N_21665,N_19082);
and U22449 (N_22449,N_19796,N_20710);
or U22450 (N_22450,N_19109,N_21141);
nand U22451 (N_22451,N_20952,N_19078);
nand U22452 (N_22452,N_18759,N_20934);
nand U22453 (N_22453,N_19527,N_18885);
or U22454 (N_22454,N_18871,N_19281);
xor U22455 (N_22455,N_19471,N_19474);
or U22456 (N_22456,N_20083,N_20553);
or U22457 (N_22457,N_18927,N_19083);
xnor U22458 (N_22458,N_19049,N_19417);
nor U22459 (N_22459,N_21708,N_19039);
xor U22460 (N_22460,N_19074,N_21277);
xnor U22461 (N_22461,N_19392,N_19077);
or U22462 (N_22462,N_19540,N_20580);
and U22463 (N_22463,N_21198,N_18844);
or U22464 (N_22464,N_19901,N_20306);
xnor U22465 (N_22465,N_21017,N_19701);
xor U22466 (N_22466,N_20122,N_21129);
xnor U22467 (N_22467,N_19690,N_19760);
or U22468 (N_22468,N_18848,N_20840);
and U22469 (N_22469,N_21457,N_21432);
nand U22470 (N_22470,N_20971,N_19969);
nand U22471 (N_22471,N_20788,N_19510);
nand U22472 (N_22472,N_20677,N_21776);
nor U22473 (N_22473,N_21618,N_19824);
or U22474 (N_22474,N_19776,N_19278);
or U22475 (N_22475,N_21841,N_19110);
xnor U22476 (N_22476,N_20359,N_19346);
or U22477 (N_22477,N_20142,N_19735);
and U22478 (N_22478,N_19367,N_18919);
and U22479 (N_22479,N_21761,N_20061);
nand U22480 (N_22480,N_19485,N_18941);
or U22481 (N_22481,N_21464,N_21250);
nor U22482 (N_22482,N_19989,N_19762);
nor U22483 (N_22483,N_19298,N_19756);
xnor U22484 (N_22484,N_19472,N_19588);
nand U22485 (N_22485,N_19596,N_19273);
or U22486 (N_22486,N_20462,N_19051);
xor U22487 (N_22487,N_18947,N_20023);
nor U22488 (N_22488,N_19257,N_19301);
or U22489 (N_22489,N_19341,N_19460);
nor U22490 (N_22490,N_21530,N_20817);
nor U22491 (N_22491,N_20691,N_20383);
nor U22492 (N_22492,N_20628,N_20198);
xor U22493 (N_22493,N_19613,N_20543);
nor U22494 (N_22494,N_21499,N_20338);
and U22495 (N_22495,N_19893,N_20508);
or U22496 (N_22496,N_20605,N_19926);
nand U22497 (N_22497,N_20246,N_19902);
nand U22498 (N_22498,N_19511,N_19614);
and U22499 (N_22499,N_20378,N_19469);
or U22500 (N_22500,N_21224,N_19379);
xnor U22501 (N_22501,N_21626,N_20576);
xnor U22502 (N_22502,N_19328,N_21303);
xnor U22503 (N_22503,N_18914,N_21659);
or U22504 (N_22504,N_21536,N_20405);
or U22505 (N_22505,N_21021,N_21295);
and U22506 (N_22506,N_19221,N_20776);
and U22507 (N_22507,N_21764,N_19638);
xnor U22508 (N_22508,N_20352,N_21230);
nor U22509 (N_22509,N_19505,N_21624);
nor U22510 (N_22510,N_21476,N_19713);
or U22511 (N_22511,N_19753,N_20091);
and U22512 (N_22512,N_21505,N_20435);
nor U22513 (N_22513,N_19269,N_20398);
nor U22514 (N_22514,N_19143,N_20881);
nand U22515 (N_22515,N_18838,N_20650);
nor U22516 (N_22516,N_19628,N_18920);
nand U22517 (N_22517,N_19007,N_20351);
or U22518 (N_22518,N_20220,N_21090);
nand U22519 (N_22519,N_20869,N_21404);
xor U22520 (N_22520,N_18946,N_18824);
or U22521 (N_22521,N_19732,N_19583);
xnor U22522 (N_22522,N_19545,N_21832);
and U22523 (N_22523,N_19364,N_21014);
xor U22524 (N_22524,N_21043,N_18828);
and U22525 (N_22525,N_20890,N_19095);
and U22526 (N_22526,N_21566,N_21596);
or U22527 (N_22527,N_20680,N_19157);
and U22528 (N_22528,N_21465,N_19738);
nor U22529 (N_22529,N_21513,N_19287);
xnor U22530 (N_22530,N_19872,N_20044);
xor U22531 (N_22531,N_20664,N_20859);
and U22532 (N_22532,N_19029,N_21611);
and U22533 (N_22533,N_20828,N_20104);
nand U22534 (N_22534,N_20792,N_21570);
nor U22535 (N_22535,N_19140,N_19426);
nand U22536 (N_22536,N_20322,N_21361);
or U22537 (N_22537,N_21735,N_20062);
nor U22538 (N_22538,N_21852,N_21818);
nand U22539 (N_22539,N_20696,N_20325);
nand U22540 (N_22540,N_21732,N_19231);
xor U22541 (N_22541,N_19127,N_19910);
nand U22542 (N_22542,N_18925,N_21697);
nand U22543 (N_22543,N_21447,N_20183);
nand U22544 (N_22544,N_20832,N_19644);
nor U22545 (N_22545,N_21778,N_20196);
nor U22546 (N_22546,N_20648,N_19534);
nand U22547 (N_22547,N_19186,N_21869);
xnor U22548 (N_22548,N_21253,N_19948);
and U22549 (N_22549,N_20944,N_19347);
and U22550 (N_22550,N_21657,N_20603);
nor U22551 (N_22551,N_21259,N_19201);
xnor U22552 (N_22552,N_19580,N_18769);
xnor U22553 (N_22553,N_19791,N_21797);
and U22554 (N_22554,N_20033,N_19064);
or U22555 (N_22555,N_20950,N_19449);
nand U22556 (N_22556,N_18823,N_20602);
nand U22557 (N_22557,N_20372,N_20456);
nand U22558 (N_22558,N_21858,N_21183);
xor U22559 (N_22559,N_20176,N_21597);
and U22560 (N_22560,N_21615,N_21359);
nor U22561 (N_22561,N_21294,N_19103);
or U22562 (N_22562,N_20727,N_21405);
nand U22563 (N_22563,N_21532,N_20608);
nand U22564 (N_22564,N_21551,N_19133);
or U22565 (N_22565,N_21771,N_21677);
nor U22566 (N_22566,N_20874,N_20674);
nand U22567 (N_22567,N_19549,N_19789);
or U22568 (N_22568,N_19408,N_21337);
nand U22569 (N_22569,N_21325,N_18938);
and U22570 (N_22570,N_20304,N_20889);
xor U22571 (N_22571,N_20706,N_21516);
and U22572 (N_22572,N_20708,N_19480);
and U22573 (N_22573,N_19138,N_20925);
nor U22574 (N_22574,N_21174,N_20758);
nand U22575 (N_22575,N_19715,N_20595);
and U22576 (N_22576,N_21480,N_20790);
xor U22577 (N_22577,N_19399,N_20072);
xor U22578 (N_22578,N_21058,N_20865);
nand U22579 (N_22579,N_19842,N_19372);
nand U22580 (N_22580,N_19665,N_21836);
or U22581 (N_22581,N_20010,N_19987);
nand U22582 (N_22582,N_19729,N_19491);
or U22583 (N_22583,N_19429,N_19924);
nand U22584 (N_22584,N_18792,N_21703);
xor U22585 (N_22585,N_18878,N_21848);
and U22586 (N_22586,N_21791,N_21557);
nand U22587 (N_22587,N_21616,N_20144);
and U22588 (N_22588,N_20026,N_19466);
and U22589 (N_22589,N_20774,N_19276);
nand U22590 (N_22590,N_21424,N_20829);
nor U22591 (N_22591,N_21599,N_20715);
xor U22592 (N_22592,N_20067,N_20794);
nand U22593 (N_22593,N_21237,N_20428);
or U22594 (N_22594,N_21104,N_21649);
or U22595 (N_22595,N_21839,N_20388);
xnor U22596 (N_22596,N_19144,N_19188);
and U22597 (N_22597,N_19337,N_20679);
nor U22598 (N_22598,N_21134,N_18888);
xor U22599 (N_22599,N_19669,N_21668);
xnor U22600 (N_22600,N_20217,N_20699);
or U22601 (N_22601,N_19711,N_21062);
nor U22602 (N_22602,N_19254,N_20517);
and U22603 (N_22603,N_21002,N_18928);
nand U22604 (N_22604,N_21252,N_20904);
or U22605 (N_22605,N_20154,N_18989);
nor U22606 (N_22606,N_20256,N_21309);
nand U22607 (N_22607,N_20182,N_21240);
or U22608 (N_22608,N_21766,N_20396);
or U22609 (N_22609,N_20215,N_19784);
nand U22610 (N_22610,N_21363,N_21006);
and U22611 (N_22611,N_21257,N_20974);
nor U22612 (N_22612,N_21155,N_20265);
or U22613 (N_22613,N_19551,N_20162);
nand U22614 (N_22614,N_19612,N_21579);
nor U22615 (N_22615,N_19009,N_18981);
nand U22616 (N_22616,N_20740,N_21182);
and U22617 (N_22617,N_21087,N_18834);
nor U22618 (N_22618,N_20844,N_20470);
nand U22619 (N_22619,N_21838,N_21274);
xnor U22620 (N_22620,N_20195,N_20343);
xnor U22621 (N_22621,N_20108,N_21139);
and U22622 (N_22622,N_20711,N_21207);
nand U22623 (N_22623,N_18924,N_18847);
or U22624 (N_22624,N_21228,N_20523);
or U22625 (N_22625,N_21162,N_19851);
xnor U22626 (N_22626,N_20339,N_21558);
or U22627 (N_22627,N_21642,N_20487);
nand U22628 (N_22628,N_21315,N_19395);
and U22629 (N_22629,N_20877,N_19861);
nand U22630 (N_22630,N_19877,N_21510);
xor U22631 (N_22631,N_20591,N_18767);
or U22632 (N_22632,N_21630,N_20622);
xnor U22633 (N_22633,N_20688,N_21783);
xor U22634 (N_22634,N_19361,N_20966);
nand U22635 (N_22635,N_20136,N_21406);
or U22636 (N_22636,N_19030,N_19766);
nor U22637 (N_22637,N_19763,N_21748);
and U22638 (N_22638,N_19021,N_18803);
and U22639 (N_22639,N_21685,N_19307);
nor U22640 (N_22640,N_19203,N_19423);
or U22641 (N_22641,N_19330,N_20377);
xor U22642 (N_22642,N_21055,N_19456);
nand U22643 (N_22643,N_19869,N_21741);
and U22644 (N_22644,N_21036,N_20953);
xor U22645 (N_22645,N_19698,N_20053);
xnor U22646 (N_22646,N_21387,N_20002);
nor U22647 (N_22647,N_20509,N_21123);
xnor U22648 (N_22648,N_18765,N_20336);
or U22649 (N_22649,N_21306,N_20717);
nor U22650 (N_22650,N_20564,N_19876);
xor U22651 (N_22651,N_19225,N_19677);
xor U22652 (N_22652,N_21095,N_20501);
or U22653 (N_22653,N_19230,N_20411);
nand U22654 (N_22654,N_20730,N_19386);
and U22655 (N_22655,N_19600,N_21346);
nand U22656 (N_22656,N_20978,N_19572);
xor U22657 (N_22657,N_21334,N_21758);
nand U22658 (N_22658,N_21175,N_21590);
nand U22659 (N_22659,N_20536,N_20707);
and U22660 (N_22660,N_20899,N_21384);
nor U22661 (N_22661,N_19552,N_20836);
nand U22662 (N_22662,N_20318,N_21645);
xor U22663 (N_22663,N_19303,N_20852);
or U22664 (N_22664,N_21751,N_19123);
or U22665 (N_22665,N_21492,N_19661);
nand U22666 (N_22666,N_21782,N_19262);
nand U22667 (N_22667,N_21244,N_20713);
xor U22668 (N_22668,N_20300,N_19928);
nand U22669 (N_22669,N_19420,N_20324);
xor U22670 (N_22670,N_21060,N_18798);
nor U22671 (N_22671,N_19682,N_20460);
nor U22672 (N_22672,N_20618,N_21076);
and U22673 (N_22673,N_20815,N_20467);
or U22674 (N_22674,N_20588,N_20751);
or U22675 (N_22675,N_21583,N_19632);
nand U22676 (N_22676,N_19111,N_20286);
and U22677 (N_22677,N_18908,N_18901);
or U22678 (N_22678,N_21350,N_21614);
or U22679 (N_22679,N_19557,N_19093);
nand U22680 (N_22680,N_21724,N_21273);
or U22681 (N_22681,N_21621,N_21425);
or U22682 (N_22682,N_21188,N_19411);
xor U22683 (N_22683,N_20006,N_20288);
nand U22684 (N_22684,N_21809,N_21506);
or U22685 (N_22685,N_19394,N_21795);
nand U22686 (N_22686,N_20107,N_18987);
and U22687 (N_22687,N_19324,N_21242);
or U22688 (N_22688,N_19755,N_19390);
xor U22689 (N_22689,N_21072,N_20637);
and U22690 (N_22690,N_20607,N_21733);
xor U22691 (N_22691,N_18785,N_20546);
or U22692 (N_22692,N_21088,N_20700);
xnor U22693 (N_22693,N_20049,N_21153);
nor U22694 (N_22694,N_19521,N_19353);
or U22695 (N_22695,N_21052,N_18931);
xnor U22696 (N_22696,N_20697,N_21264);
and U22697 (N_22697,N_20578,N_18867);
nand U22698 (N_22698,N_19016,N_20615);
nor U22699 (N_22699,N_20274,N_21322);
xor U22700 (N_22700,N_20833,N_19227);
or U22701 (N_22701,N_19649,N_21370);
or U22702 (N_22702,N_19113,N_21872);
or U22703 (N_22703,N_20025,N_20134);
nor U22704 (N_22704,N_20521,N_21050);
nor U22705 (N_22705,N_19714,N_21606);
or U22706 (N_22706,N_20842,N_20534);
and U22707 (N_22707,N_19853,N_18853);
or U22708 (N_22708,N_19616,N_21460);
nor U22709 (N_22709,N_19504,N_19374);
and U22710 (N_22710,N_21687,N_19335);
and U22711 (N_22711,N_21810,N_20094);
nor U22712 (N_22712,N_19488,N_19933);
or U22713 (N_22713,N_20425,N_21840);
nor U22714 (N_22714,N_21867,N_20735);
or U22715 (N_22715,N_19568,N_19406);
nand U22716 (N_22716,N_20402,N_21563);
or U22717 (N_22717,N_20455,N_19026);
nand U22718 (N_22718,N_19794,N_20308);
or U22719 (N_22719,N_18836,N_20784);
nor U22720 (N_22720,N_18829,N_19496);
and U22721 (N_22721,N_19407,N_20507);
and U22722 (N_22722,N_19122,N_18913);
nor U22723 (N_22723,N_21420,N_20988);
nor U22724 (N_22724,N_19664,N_21752);
and U22725 (N_22725,N_20375,N_19042);
or U22726 (N_22726,N_21073,N_21728);
nand U22727 (N_22727,N_19293,N_20728);
nor U22728 (N_22728,N_21679,N_19132);
and U22729 (N_22729,N_19497,N_20131);
xor U22730 (N_22730,N_21005,N_21533);
nand U22731 (N_22731,N_21150,N_20616);
nor U22732 (N_22732,N_20434,N_20293);
xnor U22733 (N_22733,N_21399,N_20202);
nand U22734 (N_22734,N_19564,N_19773);
nor U22735 (N_22735,N_20921,N_19650);
or U22736 (N_22736,N_19349,N_19990);
nand U22737 (N_22737,N_19242,N_19863);
nor U22738 (N_22738,N_18783,N_18751);
or U22739 (N_22739,N_20915,N_19487);
and U22740 (N_22740,N_19811,N_20785);
and U22741 (N_22741,N_20723,N_19537);
xor U22742 (N_22742,N_19599,N_19556);
and U22743 (N_22743,N_18854,N_21314);
or U22744 (N_22744,N_20635,N_20368);
or U22745 (N_22745,N_20720,N_21843);
xor U22746 (N_22746,N_19446,N_21789);
nor U22747 (N_22747,N_21348,N_20849);
nor U22748 (N_22748,N_19031,N_20140);
nand U22749 (N_22749,N_19441,N_21142);
and U22750 (N_22750,N_20390,N_18921);
and U22751 (N_22751,N_20821,N_18898);
nand U22752 (N_22752,N_20714,N_18793);
nand U22753 (N_22753,N_19088,N_19704);
and U22754 (N_22754,N_20506,N_20495);
nor U22755 (N_22755,N_20793,N_19881);
or U22756 (N_22756,N_20224,N_19215);
or U22757 (N_22757,N_20724,N_20682);
or U22758 (N_22758,N_21496,N_21458);
nand U22759 (N_22759,N_20031,N_18929);
nand U22760 (N_22760,N_18906,N_21178);
nor U22761 (N_22761,N_21705,N_18762);
nand U22762 (N_22762,N_20541,N_21709);
or U22763 (N_22763,N_21799,N_21463);
nand U22764 (N_22764,N_19080,N_21540);
and U22765 (N_22765,N_20481,N_19807);
or U22766 (N_22766,N_19439,N_19781);
nor U22767 (N_22767,N_18752,N_19359);
or U22768 (N_22768,N_21413,N_20639);
nor U22769 (N_22769,N_19489,N_21554);
nand U22770 (N_22770,N_19369,N_18904);
nor U22771 (N_22771,N_19643,N_21116);
xor U22772 (N_22772,N_19592,N_19284);
and U22773 (N_22773,N_21461,N_21664);
xnor U22774 (N_22774,N_19416,N_21085);
nand U22775 (N_22775,N_21189,N_19911);
nand U22776 (N_22776,N_21545,N_19831);
xor U22777 (N_22777,N_19383,N_18779);
xnor U22778 (N_22778,N_20100,N_20888);
nor U22779 (N_22779,N_21234,N_21455);
xor U22780 (N_22780,N_19931,N_20445);
and U22781 (N_22781,N_20464,N_19271);
xor U22782 (N_22782,N_20996,N_21794);
or U22783 (N_22783,N_21243,N_19624);
nor U22784 (N_22784,N_19611,N_19419);
xnor U22785 (N_22785,N_20302,N_18862);
and U22786 (N_22786,N_21462,N_20087);
nand U22787 (N_22787,N_20030,N_19322);
xor U22788 (N_22788,N_19038,N_20581);
and U22789 (N_22789,N_20391,N_21736);
xor U22790 (N_22790,N_19286,N_19619);
or U22791 (N_22791,N_19629,N_21388);
or U22792 (N_22792,N_19442,N_18814);
nor U22793 (N_22793,N_21015,N_20133);
nor U22794 (N_22794,N_20659,N_20777);
nor U22795 (N_22795,N_18984,N_20227);
xor U22796 (N_22796,N_20656,N_19944);
and U22797 (N_22797,N_20880,N_20261);
or U22798 (N_22798,N_19128,N_19533);
nand U22799 (N_22799,N_19397,N_21846);
xor U22800 (N_22800,N_18926,N_20741);
and U22801 (N_22801,N_21126,N_21039);
xor U22802 (N_22802,N_20545,N_21302);
and U22803 (N_22803,N_19194,N_19356);
or U22804 (N_22804,N_21804,N_21430);
nand U22805 (N_22805,N_21269,N_21164);
and U22806 (N_22806,N_19075,N_21086);
xnor U22807 (N_22807,N_20773,N_20975);
and U22808 (N_22808,N_21689,N_20483);
xor U22809 (N_22809,N_20266,N_21398);
nor U22810 (N_22810,N_20447,N_20807);
nor U22811 (N_22811,N_20995,N_18832);
and U22812 (N_22812,N_19757,N_20382);
or U22813 (N_22813,N_19631,N_18974);
or U22814 (N_22814,N_21245,N_20208);
nand U22815 (N_22815,N_18897,N_19697);
and U22816 (N_22816,N_21770,N_19028);
xnor U22817 (N_22817,N_21578,N_20918);
xnor U22818 (N_22818,N_18780,N_20583);
nand U22819 (N_22819,N_20744,N_20169);
or U22820 (N_22820,N_21760,N_21423);
or U22821 (N_22821,N_21561,N_19180);
xor U22822 (N_22822,N_19830,N_20570);
nor U22823 (N_22823,N_21310,N_20752);
nand U22824 (N_22824,N_20126,N_21222);
and U22825 (N_22825,N_21523,N_19800);
nand U22826 (N_22826,N_21720,N_20827);
nand U22827 (N_22827,N_19656,N_19226);
nor U22828 (N_22828,N_21382,N_19285);
nor U22829 (N_22829,N_21048,N_21467);
and U22830 (N_22830,N_19119,N_18899);
and U22831 (N_22831,N_18789,N_19189);
or U22832 (N_22832,N_18998,N_20347);
nand U22833 (N_22833,N_19317,N_21815);
nor U22834 (N_22834,N_21128,N_18907);
nand U22835 (N_22835,N_21440,N_20753);
and U22836 (N_22836,N_21318,N_21179);
or U22837 (N_22837,N_20822,N_21093);
nor U22838 (N_22838,N_18831,N_21509);
nand U22839 (N_22839,N_18804,N_21223);
and U22840 (N_22840,N_20565,N_21140);
nor U22841 (N_22841,N_21426,N_20056);
nand U22842 (N_22842,N_18922,N_18915);
or U22843 (N_22843,N_19387,N_21450);
or U22844 (N_22844,N_19961,N_21850);
nand U22845 (N_22845,N_21258,N_18887);
or U22846 (N_22846,N_20407,N_21165);
xnor U22847 (N_22847,N_20376,N_19218);
or U22848 (N_22848,N_20731,N_18961);
and U22849 (N_22849,N_19833,N_21670);
or U22850 (N_22850,N_19553,N_21268);
or U22851 (N_22851,N_20158,N_19849);
nor U22852 (N_22852,N_18864,N_21047);
and U22853 (N_22853,N_19428,N_20668);
nand U22854 (N_22854,N_18852,N_20116);
or U22855 (N_22855,N_20432,N_21787);
nand U22856 (N_22856,N_20726,N_19234);
or U22857 (N_22857,N_21324,N_21101);
xor U22858 (N_22858,N_20883,N_21854);
nor U22859 (N_22859,N_20007,N_21299);
nand U22860 (N_22860,N_20174,N_21133);
nor U22861 (N_22861,N_19979,N_19676);
xnor U22862 (N_22862,N_19005,N_19555);
nand U22863 (N_22863,N_21675,N_20592);
and U22864 (N_22864,N_19843,N_19172);
or U22865 (N_22865,N_21641,N_21553);
nand U22866 (N_22866,N_19741,N_18773);
nand U22867 (N_22867,N_20497,N_21347);
xor U22868 (N_22868,N_21004,N_20327);
and U22869 (N_22869,N_19703,N_21013);
xor U22870 (N_22870,N_19803,N_20419);
or U22871 (N_22871,N_20590,N_20146);
nand U22872 (N_22872,N_21585,N_19683);
nor U22873 (N_22873,N_21527,N_18978);
nand U22874 (N_22874,N_20114,N_19193);
or U22875 (N_22875,N_20804,N_20244);
xnor U22876 (N_22876,N_20681,N_20582);
nand U22877 (N_22877,N_21191,N_19607);
nor U22878 (N_22878,N_19129,N_20178);
or U22879 (N_22879,N_19602,N_20123);
nand U22880 (N_22880,N_20055,N_20399);
xnor U22881 (N_22881,N_20839,N_21414);
nor U22882 (N_22882,N_20063,N_20120);
or U22883 (N_22883,N_21711,N_21027);
and U22884 (N_22884,N_21231,N_20027);
or U22885 (N_22885,N_21662,N_21535);
nor U22886 (N_22886,N_21715,N_21774);
nor U22887 (N_22887,N_21746,N_20667);
and U22888 (N_22888,N_18825,N_21773);
and U22889 (N_22889,N_21281,N_18966);
nand U22890 (N_22890,N_18859,N_19164);
and U22891 (N_22891,N_18766,N_20903);
xor U22892 (N_22892,N_20250,N_19675);
nor U22893 (N_22893,N_20163,N_19086);
and U22894 (N_22894,N_19477,N_20235);
xor U22895 (N_22895,N_18996,N_20200);
xor U22896 (N_22896,N_21512,N_21326);
or U22897 (N_22897,N_19885,N_19589);
nor U22898 (N_22898,N_20745,N_21083);
and U22899 (N_22899,N_21340,N_21714);
xor U22900 (N_22900,N_21763,N_19908);
nand U22901 (N_22901,N_19125,N_21098);
and U22902 (N_22902,N_21160,N_20077);
nand U22903 (N_22903,N_21304,N_20436);
xor U22904 (N_22904,N_20510,N_21053);
nand U22905 (N_22905,N_21491,N_21454);
xnor U22906 (N_22906,N_19685,N_21271);
or U22907 (N_22907,N_18951,N_21577);
and U22908 (N_22908,N_21168,N_18784);
nand U22909 (N_22909,N_20586,N_20956);
xor U22910 (N_22910,N_19358,N_19795);
and U22911 (N_22911,N_19440,N_21562);
xnor U22912 (N_22912,N_19217,N_21428);
or U22913 (N_22913,N_19706,N_21111);
xnor U22914 (N_22914,N_20038,N_19708);
nor U22915 (N_22915,N_20490,N_19520);
or U22916 (N_22916,N_20783,N_21631);
nor U22917 (N_22917,N_21873,N_21784);
nand U22918 (N_22918,N_18896,N_19782);
xor U22919 (N_22919,N_20127,N_19855);
xor U22920 (N_22920,N_18850,N_21071);
xor U22921 (N_22921,N_21105,N_20871);
or U22922 (N_22922,N_20898,N_21504);
nor U22923 (N_22923,N_19866,N_20001);
nand U22924 (N_22924,N_20585,N_20689);
and U22925 (N_22925,N_19752,N_18790);
xnor U22926 (N_22926,N_19905,N_21345);
nand U22927 (N_22927,N_21284,N_18786);
and U22928 (N_22928,N_19761,N_20734);
xor U22929 (N_22929,N_21092,N_20254);
xnor U22930 (N_22930,N_19718,N_20297);
xnor U22931 (N_22931,N_19655,N_21576);
and U22932 (N_22932,N_19239,N_21285);
nand U22933 (N_22933,N_20867,N_20480);
or U22934 (N_22934,N_19530,N_19509);
or U22935 (N_22935,N_20943,N_21820);
nand U22936 (N_22936,N_19321,N_19176);
nor U22937 (N_22937,N_19246,N_19598);
or U22938 (N_22938,N_21184,N_21768);
and U22939 (N_22939,N_21451,N_19860);
and U22940 (N_22940,N_20983,N_21161);
xor U22941 (N_22941,N_21765,N_20886);
nand U22942 (N_22942,N_18761,N_21125);
xor U22943 (N_22943,N_19938,N_21692);
and U22944 (N_22944,N_21550,N_18994);
nor U22945 (N_22945,N_20901,N_21473);
nor U22946 (N_22946,N_20442,N_20171);
or U22947 (N_22947,N_21617,N_20316);
xor U22948 (N_22948,N_20344,N_21037);
or U22949 (N_22949,N_21227,N_18995);
or U22950 (N_22950,N_20209,N_21008);
nor U22951 (N_22951,N_19743,N_20112);
and U22952 (N_22952,N_20550,N_20307);
nor U22953 (N_22953,N_19003,N_20540);
nand U22954 (N_22954,N_19834,N_19313);
nand U22955 (N_22955,N_21403,N_20922);
xnor U22956 (N_22956,N_21757,N_19342);
or U22957 (N_22957,N_19550,N_19801);
nand U22958 (N_22958,N_19889,N_21520);
xor U22959 (N_22959,N_20105,N_18768);
xor U22960 (N_22960,N_21214,N_19277);
nor U22961 (N_22961,N_20489,N_20397);
or U22962 (N_22962,N_20341,N_19253);
or U22963 (N_22963,N_21106,N_21069);
nor U22964 (N_22964,N_19213,N_20259);
nor U22965 (N_22965,N_19418,N_19506);
xnor U22966 (N_22966,N_21721,N_19954);
or U22967 (N_22967,N_20279,N_20560);
or U22968 (N_22968,N_19518,N_21591);
and U22969 (N_22969,N_19577,N_21544);
and U22970 (N_22970,N_21360,N_20791);
nor U22971 (N_22971,N_19941,N_21176);
nor U22972 (N_22972,N_19929,N_21117);
xnor U22973 (N_22973,N_20156,N_20569);
nor U22974 (N_22974,N_21648,N_21396);
or U22975 (N_22975,N_20078,N_21586);
nand U22976 (N_22976,N_19917,N_18872);
nor U22977 (N_22977,N_20180,N_21609);
and U22978 (N_22978,N_18856,N_20284);
nor U22979 (N_22979,N_21498,N_19355);
and U22980 (N_22980,N_21296,N_19573);
xnor U22981 (N_22981,N_20102,N_21096);
xnor U22982 (N_22982,N_19036,N_19925);
nand U22983 (N_22983,N_19892,N_19108);
nor U22984 (N_22984,N_19283,N_20345);
and U22985 (N_22985,N_19999,N_20353);
nor U22986 (N_22986,N_20416,N_21261);
nor U22987 (N_22987,N_18970,N_21863);
nand U22988 (N_22988,N_19978,N_18830);
or U22989 (N_22989,N_19707,N_21354);
xnor U22990 (N_22990,N_19432,N_20103);
nor U22991 (N_22991,N_19548,N_21038);
and U22992 (N_22992,N_21865,N_21828);
nand U22993 (N_22993,N_19705,N_19035);
xor U22994 (N_22994,N_19891,N_21173);
nand U22995 (N_22995,N_19888,N_20703);
or U22996 (N_22996,N_20999,N_19061);
nand U22997 (N_22997,N_21493,N_19684);
nor U22998 (N_22998,N_19447,N_20054);
or U22999 (N_22999,N_19476,N_21421);
or U23000 (N_23000,N_20305,N_20738);
or U23001 (N_23001,N_19040,N_19146);
or U23002 (N_23002,N_20672,N_19887);
and U23003 (N_23003,N_19523,N_20059);
nor U23004 (N_23004,N_19826,N_19168);
or U23005 (N_23005,N_21415,N_19081);
nand U23006 (N_23006,N_19856,N_19414);
nand U23007 (N_23007,N_21864,N_21100);
nand U23008 (N_23008,N_19839,N_20043);
xnor U23009 (N_23009,N_20204,N_21701);
nand U23010 (N_23010,N_20296,N_21503);
nand U23011 (N_23011,N_18860,N_20211);
or U23012 (N_23012,N_20694,N_20653);
and U23013 (N_23013,N_20137,N_18997);
or U23014 (N_23014,N_21035,N_20175);
nand U23015 (N_23015,N_19183,N_18794);
or U23016 (N_23016,N_19445,N_20826);
nor U23017 (N_23017,N_21241,N_19836);
xor U23018 (N_23018,N_20786,N_21418);
or U23019 (N_23019,N_19618,N_21371);
and U23020 (N_23020,N_19398,N_20763);
nand U23021 (N_23021,N_20818,N_21582);
xnor U23022 (N_23022,N_19967,N_20848);
nand U23023 (N_23023,N_20834,N_20124);
and U23024 (N_23024,N_21066,N_20997);
nand U23025 (N_23025,N_21372,N_19323);
and U23026 (N_23026,N_19076,N_21365);
and U23027 (N_23027,N_19951,N_20894);
or U23028 (N_23028,N_19333,N_18805);
and U23029 (N_23029,N_21729,N_21218);
and U23030 (N_23030,N_20360,N_20678);
nand U23031 (N_23031,N_19874,N_18939);
and U23032 (N_23032,N_19199,N_19470);
xor U23033 (N_23033,N_21202,N_21842);
or U23034 (N_23034,N_20606,N_18861);
nor U23035 (N_23035,N_21696,N_19479);
nor U23036 (N_23036,N_21672,N_21180);
and U23037 (N_23037,N_20799,N_21080);
and U23038 (N_23038,N_19247,N_20573);
nor U23039 (N_23039,N_20493,N_19822);
nor U23040 (N_23040,N_20937,N_20686);
and U23041 (N_23041,N_21640,N_21436);
nor U23042 (N_23042,N_21749,N_18820);
and U23043 (N_23043,N_19015,N_18772);
or U23044 (N_23044,N_20303,N_19914);
xnor U23045 (N_23045,N_20625,N_21482);
and U23046 (N_23046,N_21107,N_21552);
or U23047 (N_23047,N_19279,N_19089);
xnor U23048 (N_23048,N_20384,N_20249);
or U23049 (N_23049,N_20194,N_21574);
and U23050 (N_23050,N_20484,N_20526);
nand U23051 (N_23051,N_19528,N_19737);
xnor U23052 (N_23052,N_20802,N_20421);
nor U23053 (N_23053,N_21546,N_19099);
xnor U23054 (N_23054,N_19808,N_20262);
and U23055 (N_23055,N_20099,N_20657);
and U23056 (N_23056,N_19331,N_21195);
xnor U23057 (N_23057,N_21112,N_19444);
or U23058 (N_23058,N_19173,N_21485);
or U23059 (N_23059,N_19060,N_21209);
xor U23060 (N_23060,N_20084,N_19983);
nand U23061 (N_23061,N_18968,N_19865);
or U23062 (N_23062,N_19363,N_20597);
or U23063 (N_23063,N_20225,N_21029);
and U23064 (N_23064,N_20812,N_20917);
xor U23065 (N_23065,N_20213,N_19453);
nor U23066 (N_23066,N_19696,N_19266);
or U23067 (N_23067,N_18882,N_20658);
and U23068 (N_23068,N_21003,N_18797);
nor U23069 (N_23069,N_19309,N_21046);
nand U23070 (N_23070,N_20486,N_19584);
xor U23071 (N_23071,N_21034,N_19681);
nand U23072 (N_23072,N_18909,N_20008);
and U23073 (N_23073,N_18841,N_19985);
xor U23074 (N_23074,N_21788,N_19365);
nand U23075 (N_23075,N_19422,N_20809);
nor U23076 (N_23076,N_19068,N_20722);
xor U23077 (N_23077,N_20138,N_21332);
xor U23078 (N_23078,N_20537,N_19205);
and U23079 (N_23079,N_21604,N_21547);
or U23080 (N_23080,N_19689,N_19255);
and U23081 (N_23081,N_18881,N_19692);
xor U23082 (N_23082,N_19252,N_19147);
and U23083 (N_23083,N_19982,N_18900);
xor U23084 (N_23084,N_21663,N_19873);
and U23085 (N_23085,N_20900,N_19484);
or U23086 (N_23086,N_19312,N_18795);
xnor U23087 (N_23087,N_21280,N_21723);
and U23088 (N_23088,N_21501,N_20476);
nand U23089 (N_23089,N_20494,N_20457);
nor U23090 (N_23090,N_20095,N_19621);
nor U23091 (N_23091,N_21619,N_19542);
or U23092 (N_23092,N_20358,N_19840);
and U23093 (N_23093,N_21412,N_21319);
xnor U23094 (N_23094,N_19150,N_19904);
xor U23095 (N_23095,N_20048,N_20749);
xor U23096 (N_23096,N_18969,N_21262);
or U23097 (N_23097,N_20092,N_20919);
and U23098 (N_23098,N_19828,N_21588);
or U23099 (N_23099,N_19547,N_19065);
xor U23100 (N_23100,N_20278,N_21870);
and U23101 (N_23101,N_20161,N_20230);
nor U23102 (N_23102,N_21494,N_20796);
and U23103 (N_23103,N_20579,N_21608);
xnor U23104 (N_23104,N_20395,N_20167);
nor U23105 (N_23105,N_19455,N_21669);
or U23106 (N_23106,N_21078,N_21057);
nand U23107 (N_23107,N_21767,N_20705);
or U23108 (N_23108,N_20166,N_18815);
or U23109 (N_23109,N_20076,N_20692);
or U23110 (N_23110,N_20232,N_19724);
nor U23111 (N_23111,N_20548,N_19943);
nand U23112 (N_23112,N_20004,N_21130);
or U23113 (N_23113,N_18809,N_20756);
or U23114 (N_23114,N_20935,N_19410);
nor U23115 (N_23115,N_20348,N_19306);
and U23116 (N_23116,N_19968,N_19152);
or U23117 (N_23117,N_21807,N_19832);
and U23118 (N_23118,N_19958,N_21803);
nand U23119 (N_23119,N_20984,N_21605);
or U23120 (N_23120,N_21449,N_19222);
or U23121 (N_23121,N_19880,N_20346);
nor U23122 (N_23122,N_21376,N_20891);
or U23123 (N_23123,N_19997,N_20872);
or U23124 (N_23124,N_19578,N_19912);
nand U23125 (N_23125,N_21750,N_20119);
nor U23126 (N_23126,N_19430,N_21722);
or U23127 (N_23127,N_21816,N_19748);
or U23128 (N_23128,N_20469,N_19295);
nand U23129 (N_23129,N_20429,N_21353);
nand U23130 (N_23130,N_19586,N_18889);
and U23131 (N_23131,N_20721,N_20766);
nor U23132 (N_23132,N_21730,N_19251);
or U23133 (N_23133,N_21857,N_20972);
and U23134 (N_23134,N_19563,N_21790);
xor U23135 (N_23135,N_21581,N_20148);
and U23136 (N_23136,N_19382,N_21569);
nor U23137 (N_23137,N_19532,N_20527);
nor U23138 (N_23138,N_19745,N_18942);
and U23139 (N_23139,N_21247,N_20029);
or U23140 (N_23140,N_19454,N_20113);
xnor U23141 (N_23141,N_21204,N_19340);
nor U23142 (N_23142,N_19457,N_21375);
and U23143 (N_23143,N_20531,N_19165);
nor U23144 (N_23144,N_19950,N_21543);
nand U23145 (N_23145,N_18948,N_19585);
or U23146 (N_23146,N_20698,N_19181);
xor U23147 (N_23147,N_20652,N_21167);
nand U23148 (N_23148,N_21267,N_19443);
nor U23149 (N_23149,N_20155,N_18787);
and U23150 (N_23150,N_18840,N_19699);
nor U23151 (N_23151,N_21837,N_18883);
or U23152 (N_23152,N_19459,N_20226);
nor U23153 (N_23153,N_20505,N_21417);
or U23154 (N_23154,N_18868,N_21802);
and U23155 (N_23155,N_19799,N_19538);
xnor U23156 (N_23156,N_20532,N_21276);
or U23157 (N_23157,N_21620,N_20816);
nor U23158 (N_23158,N_19427,N_21335);
nor U23159 (N_23159,N_20281,N_21650);
or U23160 (N_23160,N_19709,N_19723);
nand U23161 (N_23161,N_19458,N_21067);
nand U23162 (N_23162,N_20897,N_19774);
xnor U23163 (N_23163,N_19391,N_21246);
nand U23164 (N_23164,N_19405,N_19962);
xor U23165 (N_23165,N_19139,N_20856);
nand U23166 (N_23166,N_21362,N_19597);
xor U23167 (N_23167,N_21144,N_19878);
or U23168 (N_23168,N_21537,N_19011);
xor U23169 (N_23169,N_18940,N_19256);
nand U23170 (N_23170,N_20285,N_20911);
or U23171 (N_23171,N_18957,N_21221);
xor U23172 (N_23172,N_21682,N_20290);
xnor U23173 (N_23173,N_19814,N_19744);
nand U23174 (N_23174,N_20633,N_20780);
nand U23175 (N_23175,N_20797,N_19956);
and U23176 (N_23176,N_20186,N_19092);
nor U23177 (N_23177,N_20150,N_19066);
or U23178 (N_23178,N_19258,N_19008);
or U23179 (N_23179,N_19206,N_19010);
or U23180 (N_23180,N_21256,N_20613);
or U23181 (N_23181,N_19112,N_19282);
nand U23182 (N_23182,N_19326,N_20231);
nor U23183 (N_23183,N_18890,N_18884);
nand U23184 (N_23184,N_19890,N_20340);
nor U23185 (N_23185,N_18923,N_19747);
and U23186 (N_23186,N_21434,N_20661);
and U23187 (N_23187,N_20453,N_19582);
and U23188 (N_23188,N_18811,N_19202);
or U23189 (N_23189,N_21185,N_21019);
and U23190 (N_23190,N_19742,N_19373);
nand U23191 (N_23191,N_20283,N_21855);
and U23192 (N_23192,N_19695,N_21567);
xor U23193 (N_23193,N_20965,N_18964);
nand U23194 (N_23194,N_21678,N_19073);
xor U23195 (N_23195,N_20234,N_19385);
xor U23196 (N_23196,N_20533,N_19653);
nor U23197 (N_23197,N_21769,N_20361);
or U23198 (N_23198,N_20452,N_20090);
nor U23199 (N_23199,N_19339,N_20022);
nor U23200 (N_23200,N_19875,N_20970);
or U23201 (N_23201,N_19909,N_21082);
or U23202 (N_23202,N_20012,N_19300);
xnor U23203 (N_23203,N_20742,N_19002);
xor U23204 (N_23204,N_18837,N_19759);
nand U23205 (N_23205,N_19344,N_21011);
xor U23206 (N_23206,N_21727,N_21808);
and U23207 (N_23207,N_19393,N_21386);
or U23208 (N_23208,N_21041,N_21613);
xnor U23209 (N_23209,N_21534,N_21541);
or U23210 (N_23210,N_20190,N_21157);
or U23211 (N_23211,N_19299,N_20577);
nand U23212 (N_23212,N_19211,N_19764);
nand U23213 (N_23213,N_20709,N_21394);
nor U23214 (N_23214,N_20264,N_20458);
or U23215 (N_23215,N_21806,N_19200);
nand U23216 (N_23216,N_19862,N_21623);
or U23217 (N_23217,N_19261,N_20157);
nor U23218 (N_23218,N_21474,N_20530);
nor U23219 (N_23219,N_18952,N_21443);
nor U23220 (N_23220,N_20857,N_21103);
xnor U23221 (N_23221,N_20908,N_21452);
nand U23222 (N_23222,N_20443,N_21114);
nor U23223 (N_23223,N_20993,N_21091);
and U23224 (N_23224,N_19957,N_19348);
or U23225 (N_23225,N_21288,N_18992);
or U23226 (N_23226,N_19868,N_20693);
and U23227 (N_23227,N_21378,N_20081);
and U23228 (N_23228,N_20401,N_19513);
nor U23229 (N_23229,N_19637,N_21756);
nor U23230 (N_23230,N_20593,N_20750);
xor U23231 (N_23231,N_19932,N_21022);
xnor U23232 (N_23232,N_19930,N_20036);
nor U23233 (N_23233,N_19939,N_19241);
or U23234 (N_23234,N_19131,N_19159);
nor U23235 (N_23235,N_18975,N_20337);
nor U23236 (N_23236,N_19940,N_19818);
xor U23237 (N_23237,N_19565,N_19720);
xnor U23238 (N_23238,N_21502,N_21380);
or U23239 (N_23239,N_20064,N_20513);
nand U23240 (N_23240,N_19237,N_20701);
nor U23241 (N_23241,N_19502,N_19137);
or U23242 (N_23242,N_19091,N_20159);
or U23243 (N_23243,N_20188,N_19184);
or U23244 (N_23244,N_21743,N_19130);
nand U23245 (N_23245,N_20440,N_19765);
nand U23246 (N_23246,N_20216,N_20587);
or U23247 (N_23247,N_19149,N_21691);
or U23248 (N_23248,N_21068,N_20459);
or U23249 (N_23249,N_19852,N_21525);
or U23250 (N_23250,N_19805,N_20403);
and U23251 (N_23251,N_21308,N_21695);
xor U23252 (N_23252,N_20326,N_20941);
or U23253 (N_23253,N_21094,N_19228);
nand U23254 (N_23254,N_19835,N_20683);
and U23255 (N_23255,N_18893,N_18874);
nand U23256 (N_23256,N_21192,N_20599);
and U23257 (N_23257,N_19167,N_19590);
and U23258 (N_23258,N_19595,N_20504);
or U23259 (N_23259,N_21357,N_18818);
xnor U23260 (N_23260,N_20301,N_20837);
and U23261 (N_23261,N_20500,N_20073);
nand U23262 (N_23262,N_19235,N_19636);
nand U23263 (N_23263,N_20555,N_20967);
xor U23264 (N_23264,N_19024,N_19120);
and U23265 (N_23265,N_18972,N_19896);
and U23266 (N_23266,N_19995,N_20197);
or U23267 (N_23267,N_21115,N_20239);
nor U23268 (N_23268,N_19526,N_21075);
and U23269 (N_23269,N_21149,N_18973);
and U23270 (N_23270,N_21377,N_20782);
nand U23271 (N_23271,N_20381,N_20060);
nor U23272 (N_23272,N_20645,N_21422);
xor U23273 (N_23273,N_20801,N_19272);
or U23274 (N_23274,N_19106,N_21390);
xor U23275 (N_23275,N_19207,N_20558);
or U23276 (N_23276,N_19118,N_19014);
nand U23277 (N_23277,N_21032,N_21819);
xnor U23278 (N_23278,N_20039,N_20951);
nand U23279 (N_23279,N_20191,N_18788);
or U23280 (N_23280,N_20875,N_19886);
or U23281 (N_23281,N_19169,N_20117);
nor U23282 (N_23282,N_19357,N_19329);
xnor U23283 (N_23283,N_19473,N_18879);
and U23284 (N_23284,N_20292,N_21255);
or U23285 (N_23285,N_21521,N_21827);
and U23286 (N_23286,N_20272,N_18956);
nor U23287 (N_23287,N_21812,N_20524);
nor U23288 (N_23288,N_18849,N_21517);
and U23289 (N_23289,N_21484,N_21524);
nor U23290 (N_23290,N_21033,N_19916);
nand U23291 (N_23291,N_20321,N_21312);
nor U23292 (N_23292,N_20989,N_19918);
xor U23293 (N_23293,N_19087,N_21201);
nand U23294 (N_23294,N_20640,N_20851);
or U23295 (N_23295,N_21704,N_19052);
and U23296 (N_23296,N_19937,N_21186);
or U23297 (N_23297,N_19182,N_20755);
nand U23298 (N_23298,N_21651,N_19935);
or U23299 (N_23299,N_18813,N_20535);
nor U23300 (N_23300,N_19462,N_21272);
nor U23301 (N_23301,N_19882,N_19667);
nand U23302 (N_23302,N_18950,N_21555);
or U23303 (N_23303,N_20028,N_19481);
or U23304 (N_23304,N_20331,N_19541);
or U23305 (N_23305,N_19209,N_20109);
nor U23306 (N_23306,N_18955,N_20357);
nand U23307 (N_23307,N_18945,N_19658);
nand U23308 (N_23308,N_19536,N_20552);
and U23309 (N_23309,N_19490,N_20400);
nor U23310 (N_23310,N_21030,N_19827);
or U23311 (N_23311,N_19786,N_20101);
xor U23312 (N_23312,N_21374,N_20596);
nand U23313 (N_23313,N_20287,N_21781);
nand U23314 (N_23314,N_18971,N_20762);
and U23315 (N_23315,N_21438,N_21297);
xor U23316 (N_23316,N_19400,N_19605);
nand U23317 (N_23317,N_19543,N_20981);
or U23318 (N_23318,N_21121,N_19017);
nor U23319 (N_23319,N_21137,N_20968);
or U23320 (N_23320,N_21681,N_19516);
nor U23321 (N_23321,N_20704,N_21633);
and U23322 (N_23322,N_20930,N_20779);
or U23323 (N_23323,N_19771,N_20424);
or U23324 (N_23324,N_20914,N_20446);
or U23325 (N_23325,N_20632,N_19810);
or U23326 (N_23326,N_19377,N_21486);
nand U23327 (N_23327,N_20498,N_19758);
and U23328 (N_23328,N_20976,N_20185);
nor U23329 (N_23329,N_18999,N_19243);
and U23330 (N_23330,N_21146,N_21154);
nand U23331 (N_23331,N_20949,N_21441);
nor U23332 (N_23332,N_21531,N_18846);
xor U23333 (N_23333,N_21446,N_21063);
or U23334 (N_23334,N_21598,N_19722);
and U23335 (N_23335,N_21468,N_21654);
nand U23336 (N_23336,N_19992,N_19903);
xor U23337 (N_23337,N_20878,N_20665);
and U23338 (N_23338,N_18858,N_21118);
or U23339 (N_23339,N_21225,N_19531);
nor U23340 (N_23340,N_21317,N_21625);
nor U23341 (N_23341,N_21874,N_20685);
and U23342 (N_23342,N_19229,N_18778);
nand U23343 (N_23343,N_19854,N_19998);
or U23344 (N_23344,N_21023,N_19096);
and U23345 (N_23345,N_21483,N_19587);
nor U23346 (N_23346,N_19559,N_19820);
xor U23347 (N_23347,N_19934,N_19000);
nand U23348 (N_23348,N_21792,N_20097);
nor U23349 (N_23349,N_20671,N_20611);
nand U23350 (N_23350,N_20991,N_19098);
nor U23351 (N_23351,N_19057,N_20770);
xnor U23352 (N_23352,N_20798,N_20362);
nand U23353 (N_23353,N_19717,N_20366);
nand U23354 (N_23354,N_19652,N_20046);
xnor U23355 (N_23355,N_21169,N_20695);
and U23356 (N_23356,N_19294,N_20896);
or U23357 (N_23357,N_18959,N_19136);
and U23358 (N_23358,N_21639,N_19156);
nand U23359 (N_23359,N_20876,N_21860);
xnor U23360 (N_23360,N_20862,N_20295);
or U23361 (N_23361,N_20214,N_20830);
nand U23362 (N_23362,N_21448,N_19463);
or U23363 (N_23363,N_20748,N_20128);
or U23364 (N_23364,N_20561,N_20018);
nand U23365 (N_23365,N_19953,N_20093);
nor U23366 (N_23366,N_20242,N_18839);
or U23367 (N_23367,N_20420,N_21826);
nand U23368 (N_23368,N_20964,N_20237);
and U23369 (N_23369,N_20663,N_20040);
nand U23370 (N_23370,N_20554,N_20913);
nand U23371 (N_23371,N_21627,N_19351);
and U23372 (N_23372,N_21762,N_19404);
xor U23373 (N_23373,N_21343,N_21825);
and U23374 (N_23374,N_20408,N_20850);
and U23375 (N_23375,N_20409,N_20294);
or U23376 (N_23376,N_20177,N_19402);
nor U23377 (N_23377,N_21219,N_19338);
or U23378 (N_23378,N_21351,N_19864);
and U23379 (N_23379,N_19959,N_19126);
nand U23380 (N_23380,N_19971,N_19396);
nand U23381 (N_23381,N_19413,N_18986);
and U23382 (N_23382,N_20485,N_20808);
and U23383 (N_23383,N_19991,N_19662);
nand U23384 (N_23384,N_21572,N_19162);
and U23385 (N_23385,N_19947,N_20363);
xor U23386 (N_23386,N_20666,N_18962);
xnor U23387 (N_23387,N_21307,N_18827);
and U23388 (N_23388,N_18866,N_20525);
xor U23389 (N_23389,N_21132,N_21475);
nor U23390 (N_23390,N_21323,N_20905);
and U23391 (N_23391,N_21056,N_19883);
xor U23392 (N_23392,N_20269,N_21213);
nor U23393 (N_23393,N_19646,N_21853);
nand U23394 (N_23394,N_19769,N_20864);
nand U23395 (N_23395,N_21409,N_21026);
nand U23396 (N_23396,N_19044,N_20248);
or U23397 (N_23397,N_20145,N_20098);
or U23398 (N_23398,N_19719,N_21330);
and U23399 (N_23399,N_19733,N_21656);
nand U23400 (N_23400,N_21666,N_21507);
and U23401 (N_23401,N_21716,N_21215);
or U23402 (N_23402,N_21320,N_19503);
nor U23403 (N_23403,N_19517,N_21159);
or U23404 (N_23404,N_19994,N_19153);
xor U23405 (N_23405,N_21216,N_20562);
or U23406 (N_23406,N_20982,N_20814);
nand U23407 (N_23407,N_19114,N_19691);
or U23408 (N_23408,N_21637,N_20987);
nand U23409 (N_23409,N_21528,N_19783);
nand U23410 (N_23410,N_20393,N_20729);
or U23411 (N_23411,N_19023,N_20492);
xnor U23412 (N_23412,N_21120,N_20910);
or U23413 (N_23413,N_21601,N_20370);
nand U23414 (N_23414,N_20960,N_19512);
nand U23415 (N_23415,N_21712,N_18775);
nor U23416 (N_23416,N_19975,N_21135);
nor U23417 (N_23417,N_19846,N_19610);
and U23418 (N_23418,N_20477,N_20422);
xnor U23419 (N_23419,N_19070,N_20068);
nand U23420 (N_23420,N_20089,N_21805);
nand U23421 (N_23421,N_20465,N_19334);
nand U23422 (N_23422,N_21147,N_20627);
or U23423 (N_23423,N_19296,N_19084);
xnor U23424 (N_23424,N_21595,N_20887);
and U23425 (N_23425,N_19620,N_19208);
and U23426 (N_23426,N_18902,N_20282);
xor U23427 (N_23427,N_21592,N_19025);
or U23428 (N_23428,N_21077,N_21471);
or U23429 (N_23429,N_20085,N_21686);
nor U23430 (N_23430,N_21328,N_19004);
and U23431 (N_23431,N_21341,N_20518);
nor U23432 (N_23432,N_21392,N_20172);
xnor U23433 (N_23433,N_18819,N_20032);
or U23434 (N_23434,N_20823,N_21477);
nand U23435 (N_23435,N_19775,N_20335);
nor U23436 (N_23436,N_20931,N_21660);
nand U23437 (N_23437,N_20702,N_21735);
nor U23438 (N_23438,N_19341,N_20042);
xnor U23439 (N_23439,N_20241,N_20997);
or U23440 (N_23440,N_20988,N_20519);
or U23441 (N_23441,N_19783,N_19696);
or U23442 (N_23442,N_19828,N_20811);
and U23443 (N_23443,N_21591,N_21295);
and U23444 (N_23444,N_20893,N_19067);
xor U23445 (N_23445,N_20506,N_21546);
or U23446 (N_23446,N_21432,N_21340);
xor U23447 (N_23447,N_20112,N_21472);
or U23448 (N_23448,N_20216,N_19614);
xnor U23449 (N_23449,N_21778,N_21064);
xnor U23450 (N_23450,N_21687,N_19289);
nand U23451 (N_23451,N_19944,N_19613);
nor U23452 (N_23452,N_19585,N_19264);
nor U23453 (N_23453,N_21631,N_20867);
nand U23454 (N_23454,N_19337,N_20391);
or U23455 (N_23455,N_20909,N_20400);
and U23456 (N_23456,N_18966,N_21479);
or U23457 (N_23457,N_19286,N_20155);
and U23458 (N_23458,N_21848,N_18991);
xor U23459 (N_23459,N_19123,N_21311);
nor U23460 (N_23460,N_20392,N_19856);
nor U23461 (N_23461,N_19598,N_20789);
nand U23462 (N_23462,N_20392,N_21104);
or U23463 (N_23463,N_20135,N_20430);
and U23464 (N_23464,N_21206,N_21450);
nand U23465 (N_23465,N_18791,N_19718);
or U23466 (N_23466,N_19138,N_20985);
nor U23467 (N_23467,N_19274,N_20233);
nand U23468 (N_23468,N_21577,N_20609);
and U23469 (N_23469,N_19586,N_19786);
nor U23470 (N_23470,N_21861,N_19403);
xnor U23471 (N_23471,N_19623,N_20325);
and U23472 (N_23472,N_18784,N_21656);
xor U23473 (N_23473,N_20198,N_21261);
or U23474 (N_23474,N_19580,N_21731);
xor U23475 (N_23475,N_21673,N_20709);
nand U23476 (N_23476,N_20551,N_20378);
and U23477 (N_23477,N_19647,N_19372);
or U23478 (N_23478,N_21138,N_21261);
nand U23479 (N_23479,N_21393,N_21140);
and U23480 (N_23480,N_21746,N_19338);
and U23481 (N_23481,N_20203,N_19735);
xor U23482 (N_23482,N_20103,N_20238);
or U23483 (N_23483,N_20366,N_19981);
and U23484 (N_23484,N_19284,N_21813);
or U23485 (N_23485,N_19009,N_20774);
or U23486 (N_23486,N_21354,N_20693);
xnor U23487 (N_23487,N_20633,N_20776);
nand U23488 (N_23488,N_18826,N_19996);
nand U23489 (N_23489,N_20855,N_21775);
xnor U23490 (N_23490,N_20369,N_19538);
or U23491 (N_23491,N_20611,N_19420);
xor U23492 (N_23492,N_20571,N_20575);
and U23493 (N_23493,N_19476,N_20219);
nor U23494 (N_23494,N_20166,N_20686);
and U23495 (N_23495,N_18817,N_21413);
nand U23496 (N_23496,N_21221,N_19229);
or U23497 (N_23497,N_19224,N_20783);
or U23498 (N_23498,N_19321,N_19144);
nor U23499 (N_23499,N_21001,N_20529);
and U23500 (N_23500,N_20576,N_20757);
and U23501 (N_23501,N_21866,N_20238);
and U23502 (N_23502,N_21739,N_21368);
nor U23503 (N_23503,N_20115,N_21486);
or U23504 (N_23504,N_21536,N_19737);
and U23505 (N_23505,N_18870,N_21015);
nor U23506 (N_23506,N_19253,N_21222);
nand U23507 (N_23507,N_21376,N_20450);
xor U23508 (N_23508,N_18826,N_21874);
and U23509 (N_23509,N_19579,N_19369);
nor U23510 (N_23510,N_21509,N_18775);
nor U23511 (N_23511,N_21624,N_21658);
and U23512 (N_23512,N_20560,N_19434);
nand U23513 (N_23513,N_21010,N_19836);
and U23514 (N_23514,N_21373,N_21490);
or U23515 (N_23515,N_19004,N_20135);
nand U23516 (N_23516,N_20370,N_19177);
nor U23517 (N_23517,N_20394,N_20131);
or U23518 (N_23518,N_19495,N_21708);
nand U23519 (N_23519,N_20214,N_20712);
or U23520 (N_23520,N_20962,N_21570);
and U23521 (N_23521,N_21523,N_20094);
xor U23522 (N_23522,N_21231,N_19534);
xor U23523 (N_23523,N_19505,N_18824);
and U23524 (N_23524,N_19241,N_19963);
nand U23525 (N_23525,N_20214,N_20786);
nor U23526 (N_23526,N_20891,N_20668);
or U23527 (N_23527,N_20373,N_21210);
or U23528 (N_23528,N_20778,N_20644);
xnor U23529 (N_23529,N_21655,N_19593);
nand U23530 (N_23530,N_20995,N_18800);
xor U23531 (N_23531,N_19714,N_19449);
nor U23532 (N_23532,N_21586,N_18836);
nor U23533 (N_23533,N_19235,N_21594);
xnor U23534 (N_23534,N_20130,N_21027);
nand U23535 (N_23535,N_19347,N_20140);
nand U23536 (N_23536,N_19228,N_19070);
and U23537 (N_23537,N_21339,N_21566);
nor U23538 (N_23538,N_19026,N_20263);
nand U23539 (N_23539,N_21542,N_19181);
nand U23540 (N_23540,N_21511,N_20731);
and U23541 (N_23541,N_19993,N_19784);
xnor U23542 (N_23542,N_18959,N_21344);
nor U23543 (N_23543,N_21527,N_20924);
or U23544 (N_23544,N_21862,N_19527);
xnor U23545 (N_23545,N_21377,N_21434);
nor U23546 (N_23546,N_20308,N_20829);
xor U23547 (N_23547,N_21778,N_19652);
or U23548 (N_23548,N_21236,N_20377);
nand U23549 (N_23549,N_21538,N_19563);
xnor U23550 (N_23550,N_20044,N_20926);
nor U23551 (N_23551,N_21458,N_19034);
or U23552 (N_23552,N_18921,N_20560);
nor U23553 (N_23553,N_18848,N_19102);
nor U23554 (N_23554,N_20894,N_20338);
nand U23555 (N_23555,N_19798,N_19905);
xor U23556 (N_23556,N_21041,N_21158);
and U23557 (N_23557,N_21224,N_20013);
or U23558 (N_23558,N_21176,N_20091);
nand U23559 (N_23559,N_18905,N_19264);
or U23560 (N_23560,N_19192,N_19208);
nand U23561 (N_23561,N_21002,N_19421);
or U23562 (N_23562,N_20005,N_20048);
and U23563 (N_23563,N_20717,N_21329);
nand U23564 (N_23564,N_19060,N_20516);
nand U23565 (N_23565,N_20145,N_21330);
nor U23566 (N_23566,N_19778,N_20867);
nand U23567 (N_23567,N_21633,N_21470);
and U23568 (N_23568,N_19404,N_20277);
nand U23569 (N_23569,N_20845,N_18919);
or U23570 (N_23570,N_21431,N_20877);
or U23571 (N_23571,N_19381,N_20671);
and U23572 (N_23572,N_18783,N_21250);
or U23573 (N_23573,N_19230,N_18853);
or U23574 (N_23574,N_19797,N_20772);
nand U23575 (N_23575,N_20537,N_19794);
and U23576 (N_23576,N_21141,N_19512);
xnor U23577 (N_23577,N_21454,N_19882);
xnor U23578 (N_23578,N_19973,N_21055);
or U23579 (N_23579,N_18771,N_20828);
or U23580 (N_23580,N_21738,N_20638);
xnor U23581 (N_23581,N_20933,N_20738);
nor U23582 (N_23582,N_21623,N_20664);
or U23583 (N_23583,N_20134,N_20280);
or U23584 (N_23584,N_19205,N_21100);
xnor U23585 (N_23585,N_21503,N_20798);
nand U23586 (N_23586,N_19467,N_19842);
or U23587 (N_23587,N_21086,N_20104);
nand U23588 (N_23588,N_21621,N_18901);
or U23589 (N_23589,N_20007,N_18769);
xor U23590 (N_23590,N_19373,N_20688);
nor U23591 (N_23591,N_21318,N_19241);
nand U23592 (N_23592,N_19768,N_20684);
xnor U23593 (N_23593,N_19944,N_20988);
xnor U23594 (N_23594,N_20790,N_18842);
nand U23595 (N_23595,N_20087,N_19599);
nor U23596 (N_23596,N_19580,N_21440);
and U23597 (N_23597,N_21044,N_18823);
nand U23598 (N_23598,N_20409,N_19198);
or U23599 (N_23599,N_21536,N_19516);
xnor U23600 (N_23600,N_21037,N_18803);
and U23601 (N_23601,N_20006,N_19371);
nor U23602 (N_23602,N_19032,N_18804);
xnor U23603 (N_23603,N_21050,N_21771);
nor U23604 (N_23604,N_20450,N_21499);
xnor U23605 (N_23605,N_21633,N_20869);
nand U23606 (N_23606,N_19873,N_21006);
nor U23607 (N_23607,N_19266,N_19844);
nand U23608 (N_23608,N_19320,N_19073);
xor U23609 (N_23609,N_19768,N_18885);
or U23610 (N_23610,N_21576,N_19028);
nand U23611 (N_23611,N_20568,N_20245);
or U23612 (N_23612,N_18969,N_19268);
xnor U23613 (N_23613,N_21350,N_21238);
and U23614 (N_23614,N_19858,N_21233);
or U23615 (N_23615,N_20582,N_19032);
or U23616 (N_23616,N_19400,N_21465);
nor U23617 (N_23617,N_19983,N_21298);
nand U23618 (N_23618,N_20612,N_20163);
nand U23619 (N_23619,N_20677,N_21850);
or U23620 (N_23620,N_21219,N_21327);
nor U23621 (N_23621,N_20542,N_20841);
nand U23622 (N_23622,N_21318,N_19305);
or U23623 (N_23623,N_19092,N_21407);
or U23624 (N_23624,N_18911,N_19999);
nor U23625 (N_23625,N_20379,N_21589);
or U23626 (N_23626,N_21377,N_21551);
and U23627 (N_23627,N_21150,N_18871);
and U23628 (N_23628,N_20720,N_21386);
xnor U23629 (N_23629,N_20403,N_20601);
and U23630 (N_23630,N_20394,N_19865);
or U23631 (N_23631,N_19814,N_19228);
nand U23632 (N_23632,N_21526,N_21308);
and U23633 (N_23633,N_21199,N_19686);
or U23634 (N_23634,N_19485,N_19908);
and U23635 (N_23635,N_19291,N_19010);
nor U23636 (N_23636,N_20608,N_21585);
xor U23637 (N_23637,N_20227,N_19916);
xor U23638 (N_23638,N_20420,N_20466);
or U23639 (N_23639,N_19800,N_21452);
or U23640 (N_23640,N_19362,N_21692);
and U23641 (N_23641,N_21688,N_18954);
nor U23642 (N_23642,N_20011,N_18833);
or U23643 (N_23643,N_21644,N_21168);
nor U23644 (N_23644,N_18879,N_20095);
nor U23645 (N_23645,N_19855,N_21715);
xnor U23646 (N_23646,N_20308,N_19388);
nand U23647 (N_23647,N_19516,N_21755);
or U23648 (N_23648,N_19054,N_20002);
xnor U23649 (N_23649,N_19998,N_20853);
nand U23650 (N_23650,N_20549,N_21052);
nor U23651 (N_23651,N_20546,N_20916);
or U23652 (N_23652,N_19300,N_19181);
or U23653 (N_23653,N_19977,N_21300);
nor U23654 (N_23654,N_20657,N_19138);
nor U23655 (N_23655,N_18769,N_20674);
xor U23656 (N_23656,N_21304,N_19821);
nor U23657 (N_23657,N_19847,N_20698);
xnor U23658 (N_23658,N_18886,N_21435);
xor U23659 (N_23659,N_21203,N_18962);
and U23660 (N_23660,N_19561,N_21777);
and U23661 (N_23661,N_19540,N_21542);
and U23662 (N_23662,N_19631,N_19150);
or U23663 (N_23663,N_18785,N_19096);
nand U23664 (N_23664,N_21141,N_18869);
or U23665 (N_23665,N_19549,N_19131);
or U23666 (N_23666,N_18944,N_20703);
and U23667 (N_23667,N_19475,N_21128);
nand U23668 (N_23668,N_20969,N_20072);
nor U23669 (N_23669,N_20152,N_21617);
xor U23670 (N_23670,N_20217,N_20224);
or U23671 (N_23671,N_20638,N_20682);
nor U23672 (N_23672,N_21349,N_19623);
nand U23673 (N_23673,N_20675,N_21783);
nor U23674 (N_23674,N_20298,N_21344);
nand U23675 (N_23675,N_19241,N_20974);
or U23676 (N_23676,N_20714,N_21129);
xnor U23677 (N_23677,N_20096,N_19277);
nand U23678 (N_23678,N_18873,N_21220);
xnor U23679 (N_23679,N_19845,N_19334);
and U23680 (N_23680,N_19660,N_21582);
nand U23681 (N_23681,N_20171,N_19411);
and U23682 (N_23682,N_18846,N_20430);
and U23683 (N_23683,N_19925,N_20434);
xor U23684 (N_23684,N_19719,N_18845);
and U23685 (N_23685,N_19429,N_20318);
and U23686 (N_23686,N_20103,N_19117);
or U23687 (N_23687,N_20703,N_19897);
xor U23688 (N_23688,N_20076,N_19183);
or U23689 (N_23689,N_20700,N_20176);
or U23690 (N_23690,N_21362,N_20183);
and U23691 (N_23691,N_19594,N_20457);
or U23692 (N_23692,N_19535,N_21124);
nor U23693 (N_23693,N_21342,N_19976);
or U23694 (N_23694,N_20878,N_21049);
nor U23695 (N_23695,N_21586,N_20351);
nand U23696 (N_23696,N_20620,N_20425);
xor U23697 (N_23697,N_19159,N_19345);
nor U23698 (N_23698,N_19288,N_19233);
nand U23699 (N_23699,N_18843,N_21309);
and U23700 (N_23700,N_20249,N_20906);
xnor U23701 (N_23701,N_18872,N_21338);
xnor U23702 (N_23702,N_21505,N_19913);
xor U23703 (N_23703,N_21624,N_20101);
and U23704 (N_23704,N_20149,N_19298);
xnor U23705 (N_23705,N_21816,N_20630);
xor U23706 (N_23706,N_21083,N_20158);
nand U23707 (N_23707,N_19435,N_20679);
and U23708 (N_23708,N_19910,N_21699);
and U23709 (N_23709,N_20953,N_21318);
nand U23710 (N_23710,N_20274,N_19104);
xor U23711 (N_23711,N_21445,N_20161);
nor U23712 (N_23712,N_19971,N_20060);
xor U23713 (N_23713,N_18881,N_18785);
xnor U23714 (N_23714,N_19255,N_20343);
nand U23715 (N_23715,N_20434,N_21139);
nor U23716 (N_23716,N_19149,N_20781);
and U23717 (N_23717,N_19935,N_19982);
nor U23718 (N_23718,N_19253,N_19832);
and U23719 (N_23719,N_20608,N_18765);
nand U23720 (N_23720,N_19998,N_18906);
xnor U23721 (N_23721,N_20552,N_19041);
nand U23722 (N_23722,N_21524,N_20374);
nand U23723 (N_23723,N_21126,N_20472);
or U23724 (N_23724,N_20408,N_19562);
nand U23725 (N_23725,N_20306,N_20958);
or U23726 (N_23726,N_20224,N_18869);
xor U23727 (N_23727,N_19699,N_21319);
or U23728 (N_23728,N_19900,N_19750);
nand U23729 (N_23729,N_19547,N_19630);
nor U23730 (N_23730,N_21698,N_19692);
nand U23731 (N_23731,N_19523,N_21207);
or U23732 (N_23732,N_20505,N_19737);
xnor U23733 (N_23733,N_19103,N_19325);
xnor U23734 (N_23734,N_21032,N_19061);
nor U23735 (N_23735,N_20515,N_19119);
or U23736 (N_23736,N_19130,N_20044);
nand U23737 (N_23737,N_19318,N_19514);
or U23738 (N_23738,N_21524,N_21279);
or U23739 (N_23739,N_21449,N_20281);
xnor U23740 (N_23740,N_20325,N_20007);
nand U23741 (N_23741,N_19933,N_19611);
xnor U23742 (N_23742,N_19715,N_20830);
and U23743 (N_23743,N_21337,N_20064);
nor U23744 (N_23744,N_18922,N_19881);
nor U23745 (N_23745,N_20567,N_20126);
nor U23746 (N_23746,N_20028,N_19462);
or U23747 (N_23747,N_21327,N_19287);
or U23748 (N_23748,N_19896,N_21135);
xor U23749 (N_23749,N_20724,N_20294);
nand U23750 (N_23750,N_19208,N_19327);
nor U23751 (N_23751,N_21781,N_19238);
nor U23752 (N_23752,N_21705,N_19351);
and U23753 (N_23753,N_20519,N_20472);
nand U23754 (N_23754,N_19403,N_18806);
or U23755 (N_23755,N_19345,N_21567);
nor U23756 (N_23756,N_21872,N_19382);
nand U23757 (N_23757,N_21844,N_20880);
or U23758 (N_23758,N_19890,N_20814);
and U23759 (N_23759,N_19971,N_20798);
nor U23760 (N_23760,N_20100,N_21196);
xnor U23761 (N_23761,N_20225,N_19960);
xnor U23762 (N_23762,N_20355,N_20494);
xnor U23763 (N_23763,N_19640,N_19213);
nor U23764 (N_23764,N_20140,N_20352);
xor U23765 (N_23765,N_18760,N_21063);
or U23766 (N_23766,N_19644,N_20810);
nor U23767 (N_23767,N_19459,N_21462);
and U23768 (N_23768,N_19938,N_19324);
nand U23769 (N_23769,N_19947,N_21269);
and U23770 (N_23770,N_20455,N_19014);
nand U23771 (N_23771,N_20535,N_19688);
or U23772 (N_23772,N_21260,N_21153);
or U23773 (N_23773,N_19680,N_19966);
and U23774 (N_23774,N_19443,N_18956);
nor U23775 (N_23775,N_20185,N_20507);
nand U23776 (N_23776,N_20111,N_21498);
xnor U23777 (N_23777,N_19490,N_21047);
and U23778 (N_23778,N_19525,N_21256);
or U23779 (N_23779,N_21455,N_19734);
nor U23780 (N_23780,N_20242,N_20816);
and U23781 (N_23781,N_21142,N_21465);
xnor U23782 (N_23782,N_20239,N_20461);
or U23783 (N_23783,N_20035,N_20946);
and U23784 (N_23784,N_20885,N_20741);
and U23785 (N_23785,N_20036,N_19890);
and U23786 (N_23786,N_19446,N_19427);
or U23787 (N_23787,N_18810,N_20038);
xnor U23788 (N_23788,N_19234,N_20463);
and U23789 (N_23789,N_19544,N_20532);
xor U23790 (N_23790,N_20819,N_19389);
nand U23791 (N_23791,N_19001,N_20339);
nor U23792 (N_23792,N_21341,N_19010);
or U23793 (N_23793,N_20276,N_19636);
or U23794 (N_23794,N_21489,N_19599);
and U23795 (N_23795,N_21042,N_21732);
nand U23796 (N_23796,N_18914,N_21410);
nand U23797 (N_23797,N_21041,N_20484);
xnor U23798 (N_23798,N_19484,N_21723);
xnor U23799 (N_23799,N_19385,N_19084);
nor U23800 (N_23800,N_21635,N_20939);
nand U23801 (N_23801,N_20341,N_21240);
or U23802 (N_23802,N_21750,N_20048);
nor U23803 (N_23803,N_21831,N_18900);
or U23804 (N_23804,N_19323,N_21506);
nand U23805 (N_23805,N_19397,N_19421);
nand U23806 (N_23806,N_19930,N_18874);
nand U23807 (N_23807,N_19505,N_20438);
nor U23808 (N_23808,N_20356,N_21654);
xor U23809 (N_23809,N_19999,N_21146);
nand U23810 (N_23810,N_20821,N_21685);
or U23811 (N_23811,N_21298,N_19597);
nand U23812 (N_23812,N_20989,N_21200);
nor U23813 (N_23813,N_21453,N_19566);
and U23814 (N_23814,N_21401,N_20396);
nand U23815 (N_23815,N_19886,N_19405);
nor U23816 (N_23816,N_21386,N_19984);
nor U23817 (N_23817,N_20111,N_20207);
nor U23818 (N_23818,N_19677,N_21411);
nor U23819 (N_23819,N_19825,N_19170);
nor U23820 (N_23820,N_21304,N_20748);
or U23821 (N_23821,N_21176,N_20840);
or U23822 (N_23822,N_19114,N_20113);
and U23823 (N_23823,N_20671,N_21268);
or U23824 (N_23824,N_19834,N_20222);
xnor U23825 (N_23825,N_18955,N_19442);
nor U23826 (N_23826,N_19476,N_19868);
and U23827 (N_23827,N_21100,N_19128);
nand U23828 (N_23828,N_21017,N_19930);
nand U23829 (N_23829,N_19958,N_19646);
or U23830 (N_23830,N_21823,N_20786);
xor U23831 (N_23831,N_20001,N_20302);
nand U23832 (N_23832,N_19063,N_19108);
nand U23833 (N_23833,N_20956,N_20646);
nor U23834 (N_23834,N_21409,N_19687);
xor U23835 (N_23835,N_20248,N_19016);
xnor U23836 (N_23836,N_20127,N_21147);
nand U23837 (N_23837,N_19197,N_19182);
or U23838 (N_23838,N_21315,N_20382);
and U23839 (N_23839,N_20519,N_18826);
and U23840 (N_23840,N_20998,N_19376);
nand U23841 (N_23841,N_19057,N_20375);
nor U23842 (N_23842,N_19996,N_20215);
or U23843 (N_23843,N_19124,N_20896);
or U23844 (N_23844,N_20715,N_19247);
or U23845 (N_23845,N_20911,N_21298);
nand U23846 (N_23846,N_21812,N_19010);
nor U23847 (N_23847,N_19792,N_21313);
xor U23848 (N_23848,N_18786,N_18830);
nand U23849 (N_23849,N_21769,N_21736);
and U23850 (N_23850,N_19284,N_21593);
xor U23851 (N_23851,N_20931,N_19980);
xor U23852 (N_23852,N_21688,N_21825);
nand U23853 (N_23853,N_19589,N_18996);
nand U23854 (N_23854,N_20462,N_19289);
nor U23855 (N_23855,N_21796,N_20212);
and U23856 (N_23856,N_21642,N_21332);
or U23857 (N_23857,N_21214,N_20254);
and U23858 (N_23858,N_21287,N_20138);
xnor U23859 (N_23859,N_21782,N_21386);
nand U23860 (N_23860,N_19076,N_21585);
nand U23861 (N_23861,N_20925,N_21599);
or U23862 (N_23862,N_19675,N_19825);
xor U23863 (N_23863,N_21778,N_21053);
nand U23864 (N_23864,N_20584,N_20796);
and U23865 (N_23865,N_21309,N_21628);
nand U23866 (N_23866,N_21653,N_20562);
or U23867 (N_23867,N_19216,N_19354);
nor U23868 (N_23868,N_19713,N_18939);
or U23869 (N_23869,N_18957,N_20373);
nor U23870 (N_23870,N_19285,N_21543);
nand U23871 (N_23871,N_20288,N_20889);
or U23872 (N_23872,N_19979,N_19090);
and U23873 (N_23873,N_21672,N_21071);
and U23874 (N_23874,N_19043,N_20939);
and U23875 (N_23875,N_20949,N_19947);
and U23876 (N_23876,N_20842,N_20631);
and U23877 (N_23877,N_19066,N_19934);
xor U23878 (N_23878,N_20384,N_19200);
nand U23879 (N_23879,N_20294,N_21310);
nand U23880 (N_23880,N_21339,N_20619);
nand U23881 (N_23881,N_20800,N_19396);
or U23882 (N_23882,N_21514,N_21834);
or U23883 (N_23883,N_20203,N_18937);
nor U23884 (N_23884,N_18860,N_21265);
and U23885 (N_23885,N_19160,N_19659);
and U23886 (N_23886,N_21237,N_21128);
nand U23887 (N_23887,N_20371,N_19431);
nor U23888 (N_23888,N_19409,N_20381);
and U23889 (N_23889,N_19682,N_20764);
or U23890 (N_23890,N_20704,N_20745);
nor U23891 (N_23891,N_21677,N_20345);
and U23892 (N_23892,N_19122,N_20386);
and U23893 (N_23893,N_20643,N_19536);
nand U23894 (N_23894,N_20813,N_18874);
and U23895 (N_23895,N_18901,N_20059);
or U23896 (N_23896,N_19508,N_19069);
nand U23897 (N_23897,N_20356,N_21290);
xor U23898 (N_23898,N_20021,N_21155);
and U23899 (N_23899,N_19197,N_20151);
or U23900 (N_23900,N_19146,N_21510);
nor U23901 (N_23901,N_20252,N_19184);
and U23902 (N_23902,N_20662,N_20392);
nand U23903 (N_23903,N_20850,N_21147);
nor U23904 (N_23904,N_19046,N_21863);
or U23905 (N_23905,N_20557,N_21202);
nor U23906 (N_23906,N_20699,N_19884);
and U23907 (N_23907,N_20429,N_19936);
and U23908 (N_23908,N_20708,N_19711);
nor U23909 (N_23909,N_21412,N_19015);
xor U23910 (N_23910,N_20929,N_21582);
nor U23911 (N_23911,N_21345,N_20391);
nor U23912 (N_23912,N_19608,N_21852);
and U23913 (N_23913,N_19890,N_21510);
or U23914 (N_23914,N_21594,N_19159);
or U23915 (N_23915,N_19573,N_20829);
nor U23916 (N_23916,N_20723,N_18998);
or U23917 (N_23917,N_20956,N_21572);
nand U23918 (N_23918,N_19198,N_20579);
and U23919 (N_23919,N_19489,N_19535);
or U23920 (N_23920,N_20644,N_20486);
xnor U23921 (N_23921,N_19171,N_19533);
nor U23922 (N_23922,N_20885,N_19381);
and U23923 (N_23923,N_18798,N_21004);
xor U23924 (N_23924,N_20573,N_19580);
nand U23925 (N_23925,N_19587,N_19476);
and U23926 (N_23926,N_19396,N_19579);
or U23927 (N_23927,N_20235,N_20254);
nor U23928 (N_23928,N_20912,N_21525);
or U23929 (N_23929,N_21214,N_21539);
xnor U23930 (N_23930,N_19973,N_20693);
or U23931 (N_23931,N_21634,N_19984);
or U23932 (N_23932,N_21659,N_21547);
nand U23933 (N_23933,N_20530,N_20761);
xnor U23934 (N_23934,N_19816,N_19714);
or U23935 (N_23935,N_19489,N_21361);
nand U23936 (N_23936,N_20023,N_20773);
and U23937 (N_23937,N_20312,N_20504);
nor U23938 (N_23938,N_19024,N_21470);
nand U23939 (N_23939,N_21512,N_19366);
and U23940 (N_23940,N_19434,N_21199);
nand U23941 (N_23941,N_21669,N_19893);
and U23942 (N_23942,N_20251,N_21803);
xnor U23943 (N_23943,N_21169,N_20816);
nand U23944 (N_23944,N_21134,N_19488);
and U23945 (N_23945,N_20690,N_20157);
and U23946 (N_23946,N_21561,N_19195);
xnor U23947 (N_23947,N_19071,N_20288);
or U23948 (N_23948,N_19029,N_19371);
or U23949 (N_23949,N_20338,N_19635);
and U23950 (N_23950,N_19009,N_21761);
and U23951 (N_23951,N_21552,N_19149);
nor U23952 (N_23952,N_20510,N_19725);
or U23953 (N_23953,N_21648,N_20352);
and U23954 (N_23954,N_20823,N_19262);
and U23955 (N_23955,N_21056,N_19361);
nand U23956 (N_23956,N_20621,N_21836);
and U23957 (N_23957,N_18884,N_21500);
or U23958 (N_23958,N_20756,N_19692);
or U23959 (N_23959,N_19348,N_20630);
nand U23960 (N_23960,N_20280,N_19275);
nand U23961 (N_23961,N_19970,N_19298);
xnor U23962 (N_23962,N_19357,N_20548);
xor U23963 (N_23963,N_21587,N_20909);
and U23964 (N_23964,N_20625,N_20971);
nor U23965 (N_23965,N_19639,N_21391);
and U23966 (N_23966,N_20272,N_21686);
or U23967 (N_23967,N_21331,N_20711);
nor U23968 (N_23968,N_19923,N_19121);
or U23969 (N_23969,N_21531,N_21290);
nor U23970 (N_23970,N_19790,N_21169);
nor U23971 (N_23971,N_19267,N_19441);
nand U23972 (N_23972,N_21343,N_21779);
xor U23973 (N_23973,N_20417,N_21450);
xnor U23974 (N_23974,N_19462,N_19449);
or U23975 (N_23975,N_19734,N_19935);
xnor U23976 (N_23976,N_20799,N_21498);
nand U23977 (N_23977,N_19726,N_21465);
xnor U23978 (N_23978,N_20470,N_20412);
nand U23979 (N_23979,N_18897,N_19924);
nand U23980 (N_23980,N_20905,N_19319);
nor U23981 (N_23981,N_20451,N_18915);
xnor U23982 (N_23982,N_21657,N_21665);
and U23983 (N_23983,N_19118,N_19777);
or U23984 (N_23984,N_19787,N_21485);
nor U23985 (N_23985,N_21595,N_19571);
or U23986 (N_23986,N_19666,N_20495);
and U23987 (N_23987,N_19175,N_19711);
nor U23988 (N_23988,N_18909,N_21366);
xnor U23989 (N_23989,N_19377,N_20037);
or U23990 (N_23990,N_21680,N_20264);
or U23991 (N_23991,N_20250,N_20438);
or U23992 (N_23992,N_21378,N_19279);
or U23993 (N_23993,N_19964,N_19627);
or U23994 (N_23994,N_18972,N_20638);
nand U23995 (N_23995,N_21503,N_19960);
or U23996 (N_23996,N_20022,N_19530);
xnor U23997 (N_23997,N_21508,N_19917);
nor U23998 (N_23998,N_19059,N_20463);
nand U23999 (N_23999,N_19367,N_21273);
nor U24000 (N_24000,N_21212,N_18942);
or U24001 (N_24001,N_21152,N_20050);
nand U24002 (N_24002,N_18838,N_20867);
and U24003 (N_24003,N_18871,N_20398);
nor U24004 (N_24004,N_20224,N_20108);
nand U24005 (N_24005,N_20504,N_20816);
nor U24006 (N_24006,N_20818,N_21378);
or U24007 (N_24007,N_20087,N_19868);
and U24008 (N_24008,N_19266,N_20764);
nand U24009 (N_24009,N_19588,N_19750);
or U24010 (N_24010,N_20641,N_21042);
xnor U24011 (N_24011,N_18787,N_19878);
and U24012 (N_24012,N_21812,N_20054);
nand U24013 (N_24013,N_20381,N_20718);
xor U24014 (N_24014,N_20159,N_20095);
nor U24015 (N_24015,N_21170,N_20434);
nand U24016 (N_24016,N_20774,N_19541);
nor U24017 (N_24017,N_19505,N_19592);
or U24018 (N_24018,N_21212,N_19177);
nor U24019 (N_24019,N_20999,N_20176);
nand U24020 (N_24020,N_21419,N_19959);
nor U24021 (N_24021,N_20096,N_19557);
xnor U24022 (N_24022,N_21532,N_19307);
nor U24023 (N_24023,N_21634,N_21510);
xnor U24024 (N_24024,N_21059,N_20776);
and U24025 (N_24025,N_19284,N_18998);
nor U24026 (N_24026,N_21613,N_19682);
xor U24027 (N_24027,N_19181,N_19418);
xor U24028 (N_24028,N_20400,N_20329);
nand U24029 (N_24029,N_21612,N_21244);
or U24030 (N_24030,N_18770,N_20965);
and U24031 (N_24031,N_19137,N_21160);
nor U24032 (N_24032,N_21045,N_21020);
nor U24033 (N_24033,N_19840,N_19604);
xor U24034 (N_24034,N_20722,N_19177);
or U24035 (N_24035,N_21041,N_21688);
nor U24036 (N_24036,N_20704,N_21197);
and U24037 (N_24037,N_20815,N_21094);
nand U24038 (N_24038,N_19339,N_20010);
nand U24039 (N_24039,N_20676,N_20769);
or U24040 (N_24040,N_19980,N_21764);
nand U24041 (N_24041,N_19944,N_21771);
xnor U24042 (N_24042,N_21313,N_18898);
xor U24043 (N_24043,N_19555,N_21835);
and U24044 (N_24044,N_20952,N_20696);
or U24045 (N_24045,N_21436,N_19125);
nand U24046 (N_24046,N_18980,N_20408);
nand U24047 (N_24047,N_21317,N_21434);
xor U24048 (N_24048,N_19260,N_21165);
xnor U24049 (N_24049,N_19259,N_20010);
nand U24050 (N_24050,N_19271,N_19029);
nand U24051 (N_24051,N_20155,N_19823);
and U24052 (N_24052,N_21058,N_20485);
and U24053 (N_24053,N_19552,N_18994);
nand U24054 (N_24054,N_19280,N_20347);
and U24055 (N_24055,N_20154,N_19790);
nor U24056 (N_24056,N_19955,N_19758);
or U24057 (N_24057,N_21485,N_19507);
nor U24058 (N_24058,N_20598,N_19988);
or U24059 (N_24059,N_20768,N_21868);
nor U24060 (N_24060,N_21375,N_21246);
and U24061 (N_24061,N_19236,N_19305);
and U24062 (N_24062,N_20398,N_21300);
and U24063 (N_24063,N_19893,N_21580);
xnor U24064 (N_24064,N_19032,N_19171);
nand U24065 (N_24065,N_19513,N_21600);
and U24066 (N_24066,N_18987,N_18893);
xnor U24067 (N_24067,N_19887,N_20551);
nor U24068 (N_24068,N_21562,N_21521);
and U24069 (N_24069,N_21573,N_19850);
nor U24070 (N_24070,N_21464,N_19766);
nor U24071 (N_24071,N_21293,N_20078);
or U24072 (N_24072,N_20913,N_21410);
and U24073 (N_24073,N_19960,N_19351);
nor U24074 (N_24074,N_19295,N_19259);
xor U24075 (N_24075,N_20089,N_20773);
xnor U24076 (N_24076,N_21433,N_19038);
or U24077 (N_24077,N_19078,N_20005);
xnor U24078 (N_24078,N_19503,N_20177);
nor U24079 (N_24079,N_21490,N_19166);
and U24080 (N_24080,N_19719,N_21087);
and U24081 (N_24081,N_19215,N_19264);
xor U24082 (N_24082,N_19900,N_21082);
nand U24083 (N_24083,N_19231,N_20153);
nor U24084 (N_24084,N_18794,N_19222);
nor U24085 (N_24085,N_20348,N_21128);
nor U24086 (N_24086,N_21759,N_19207);
nand U24087 (N_24087,N_21013,N_19196);
nand U24088 (N_24088,N_20829,N_20791);
nand U24089 (N_24089,N_20003,N_20096);
nand U24090 (N_24090,N_19868,N_21598);
nor U24091 (N_24091,N_20479,N_20695);
nor U24092 (N_24092,N_20917,N_21868);
or U24093 (N_24093,N_19065,N_19650);
or U24094 (N_24094,N_19959,N_21247);
xor U24095 (N_24095,N_19670,N_21135);
nand U24096 (N_24096,N_20185,N_20482);
xnor U24097 (N_24097,N_19228,N_21248);
nand U24098 (N_24098,N_18852,N_19389);
and U24099 (N_24099,N_20798,N_19117);
nand U24100 (N_24100,N_18871,N_21250);
and U24101 (N_24101,N_20620,N_19579);
and U24102 (N_24102,N_21592,N_20119);
nor U24103 (N_24103,N_18855,N_21831);
or U24104 (N_24104,N_20792,N_20384);
xor U24105 (N_24105,N_20194,N_20147);
nor U24106 (N_24106,N_20152,N_21636);
or U24107 (N_24107,N_20305,N_20379);
nand U24108 (N_24108,N_19311,N_20358);
nor U24109 (N_24109,N_21064,N_18847);
xor U24110 (N_24110,N_19096,N_19777);
and U24111 (N_24111,N_21457,N_19618);
nor U24112 (N_24112,N_19947,N_20509);
or U24113 (N_24113,N_18976,N_20633);
nor U24114 (N_24114,N_19217,N_21678);
nor U24115 (N_24115,N_21728,N_19976);
or U24116 (N_24116,N_19936,N_21457);
nor U24117 (N_24117,N_21429,N_20424);
xor U24118 (N_24118,N_21025,N_21165);
xnor U24119 (N_24119,N_20905,N_19706);
or U24120 (N_24120,N_19456,N_19611);
or U24121 (N_24121,N_21552,N_21009);
xor U24122 (N_24122,N_19918,N_20392);
xnor U24123 (N_24123,N_19031,N_18957);
nand U24124 (N_24124,N_21209,N_20983);
xor U24125 (N_24125,N_20595,N_19236);
nand U24126 (N_24126,N_21179,N_19236);
nor U24127 (N_24127,N_21342,N_19194);
or U24128 (N_24128,N_20571,N_21535);
nand U24129 (N_24129,N_20694,N_21104);
and U24130 (N_24130,N_20623,N_20096);
nor U24131 (N_24131,N_19996,N_19767);
xnor U24132 (N_24132,N_21333,N_19910);
nand U24133 (N_24133,N_20620,N_18984);
or U24134 (N_24134,N_20843,N_21686);
nand U24135 (N_24135,N_18791,N_20691);
xor U24136 (N_24136,N_18951,N_19896);
xor U24137 (N_24137,N_20769,N_21234);
xor U24138 (N_24138,N_19035,N_21344);
or U24139 (N_24139,N_20753,N_20858);
xnor U24140 (N_24140,N_19189,N_21492);
and U24141 (N_24141,N_20515,N_18821);
or U24142 (N_24142,N_19287,N_19511);
and U24143 (N_24143,N_21508,N_19992);
or U24144 (N_24144,N_21684,N_21212);
or U24145 (N_24145,N_19157,N_19681);
or U24146 (N_24146,N_20946,N_19896);
nand U24147 (N_24147,N_21169,N_21124);
xor U24148 (N_24148,N_20971,N_20416);
nand U24149 (N_24149,N_20732,N_18780);
xnor U24150 (N_24150,N_21137,N_20979);
nor U24151 (N_24151,N_19616,N_18932);
nor U24152 (N_24152,N_21110,N_19431);
xor U24153 (N_24153,N_19656,N_21183);
and U24154 (N_24154,N_19822,N_20550);
and U24155 (N_24155,N_20511,N_20124);
nor U24156 (N_24156,N_20881,N_20337);
nor U24157 (N_24157,N_20931,N_19026);
nor U24158 (N_24158,N_19862,N_21857);
nand U24159 (N_24159,N_20227,N_19051);
nor U24160 (N_24160,N_21666,N_21506);
nand U24161 (N_24161,N_18804,N_19631);
xor U24162 (N_24162,N_21322,N_21332);
nand U24163 (N_24163,N_19565,N_20064);
nor U24164 (N_24164,N_21288,N_20794);
xnor U24165 (N_24165,N_20316,N_18941);
xnor U24166 (N_24166,N_20635,N_20919);
and U24167 (N_24167,N_19775,N_20885);
and U24168 (N_24168,N_19388,N_19809);
xnor U24169 (N_24169,N_19347,N_20893);
nor U24170 (N_24170,N_19045,N_21566);
xnor U24171 (N_24171,N_21789,N_20771);
xor U24172 (N_24172,N_19710,N_21776);
nand U24173 (N_24173,N_21247,N_21338);
or U24174 (N_24174,N_19479,N_19492);
nand U24175 (N_24175,N_20096,N_19674);
xnor U24176 (N_24176,N_20983,N_19663);
xnor U24177 (N_24177,N_21851,N_20455);
and U24178 (N_24178,N_21563,N_20512);
nand U24179 (N_24179,N_20421,N_21660);
nand U24180 (N_24180,N_19625,N_21310);
nand U24181 (N_24181,N_19830,N_19702);
xor U24182 (N_24182,N_20031,N_20062);
nand U24183 (N_24183,N_19963,N_20619);
and U24184 (N_24184,N_19251,N_19395);
nand U24185 (N_24185,N_21746,N_18910);
and U24186 (N_24186,N_20843,N_19661);
xor U24187 (N_24187,N_20448,N_20542);
xnor U24188 (N_24188,N_21019,N_21501);
nand U24189 (N_24189,N_21428,N_20714);
or U24190 (N_24190,N_18885,N_21009);
nor U24191 (N_24191,N_21279,N_21833);
nand U24192 (N_24192,N_19645,N_21261);
or U24193 (N_24193,N_20887,N_20160);
xnor U24194 (N_24194,N_18752,N_21195);
xor U24195 (N_24195,N_18829,N_18794);
nor U24196 (N_24196,N_18927,N_21792);
nand U24197 (N_24197,N_20457,N_19816);
or U24198 (N_24198,N_20262,N_20631);
nor U24199 (N_24199,N_21679,N_20571);
nor U24200 (N_24200,N_20442,N_19619);
xor U24201 (N_24201,N_20862,N_21213);
or U24202 (N_24202,N_19885,N_21498);
nor U24203 (N_24203,N_18778,N_20767);
nor U24204 (N_24204,N_21187,N_20193);
nand U24205 (N_24205,N_21519,N_21722);
xor U24206 (N_24206,N_21215,N_21561);
nand U24207 (N_24207,N_21384,N_19899);
nand U24208 (N_24208,N_20482,N_19501);
xnor U24209 (N_24209,N_20931,N_19161);
or U24210 (N_24210,N_19799,N_21193);
or U24211 (N_24211,N_20153,N_21313);
and U24212 (N_24212,N_21347,N_19294);
and U24213 (N_24213,N_19364,N_20392);
nand U24214 (N_24214,N_20551,N_21821);
or U24215 (N_24215,N_21554,N_21400);
or U24216 (N_24216,N_20977,N_20708);
nor U24217 (N_24217,N_20763,N_19728);
nand U24218 (N_24218,N_21183,N_19527);
nor U24219 (N_24219,N_20150,N_19765);
nor U24220 (N_24220,N_18829,N_20811);
xnor U24221 (N_24221,N_20183,N_18954);
nand U24222 (N_24222,N_19396,N_20491);
and U24223 (N_24223,N_19627,N_19532);
nor U24224 (N_24224,N_20204,N_20521);
and U24225 (N_24225,N_21286,N_18840);
nor U24226 (N_24226,N_20555,N_20676);
or U24227 (N_24227,N_19674,N_18855);
and U24228 (N_24228,N_20792,N_20035);
or U24229 (N_24229,N_19223,N_21204);
and U24230 (N_24230,N_21428,N_18828);
nor U24231 (N_24231,N_20189,N_21454);
nand U24232 (N_24232,N_20568,N_21112);
and U24233 (N_24233,N_19574,N_21703);
or U24234 (N_24234,N_18824,N_20162);
nand U24235 (N_24235,N_19363,N_18890);
nor U24236 (N_24236,N_19104,N_20257);
xnor U24237 (N_24237,N_18932,N_20226);
nor U24238 (N_24238,N_19480,N_21199);
nand U24239 (N_24239,N_20929,N_20394);
and U24240 (N_24240,N_20745,N_20295);
xnor U24241 (N_24241,N_19738,N_20719);
and U24242 (N_24242,N_20798,N_21823);
and U24243 (N_24243,N_20876,N_20728);
or U24244 (N_24244,N_21662,N_19755);
and U24245 (N_24245,N_21739,N_20278);
nor U24246 (N_24246,N_19647,N_21104);
or U24247 (N_24247,N_19667,N_21001);
nand U24248 (N_24248,N_20445,N_20294);
and U24249 (N_24249,N_20968,N_19986);
nor U24250 (N_24250,N_19327,N_21011);
xor U24251 (N_24251,N_20943,N_21266);
and U24252 (N_24252,N_21264,N_19878);
nand U24253 (N_24253,N_19571,N_19476);
and U24254 (N_24254,N_21677,N_19457);
or U24255 (N_24255,N_20692,N_20327);
nor U24256 (N_24256,N_21589,N_21585);
xnor U24257 (N_24257,N_19182,N_20486);
and U24258 (N_24258,N_20058,N_20770);
nand U24259 (N_24259,N_21648,N_19957);
or U24260 (N_24260,N_19059,N_21597);
and U24261 (N_24261,N_20374,N_19899);
nand U24262 (N_24262,N_19286,N_21813);
nand U24263 (N_24263,N_21018,N_21429);
and U24264 (N_24264,N_19973,N_19950);
and U24265 (N_24265,N_19277,N_19201);
xor U24266 (N_24266,N_20481,N_19077);
and U24267 (N_24267,N_20102,N_20900);
nand U24268 (N_24268,N_19592,N_20528);
nand U24269 (N_24269,N_20242,N_20308);
xnor U24270 (N_24270,N_20543,N_19115);
nor U24271 (N_24271,N_18750,N_21502);
nand U24272 (N_24272,N_20018,N_21151);
nor U24273 (N_24273,N_19617,N_19439);
or U24274 (N_24274,N_19249,N_19481);
xor U24275 (N_24275,N_19211,N_21313);
or U24276 (N_24276,N_19276,N_20242);
nor U24277 (N_24277,N_19180,N_20536);
nand U24278 (N_24278,N_21303,N_20053);
xnor U24279 (N_24279,N_20855,N_20014);
nor U24280 (N_24280,N_18779,N_18826);
nand U24281 (N_24281,N_20878,N_21620);
or U24282 (N_24282,N_18760,N_19513);
nand U24283 (N_24283,N_21064,N_20883);
and U24284 (N_24284,N_19519,N_21288);
nand U24285 (N_24285,N_19887,N_19703);
or U24286 (N_24286,N_21343,N_19651);
nand U24287 (N_24287,N_20858,N_19034);
xnor U24288 (N_24288,N_19332,N_21397);
nor U24289 (N_24289,N_20665,N_21177);
nand U24290 (N_24290,N_20938,N_19722);
nor U24291 (N_24291,N_20041,N_19437);
xor U24292 (N_24292,N_19944,N_21001);
xor U24293 (N_24293,N_20659,N_19568);
nand U24294 (N_24294,N_21464,N_21114);
nor U24295 (N_24295,N_20383,N_18932);
xor U24296 (N_24296,N_21045,N_21084);
nor U24297 (N_24297,N_18999,N_18877);
nor U24298 (N_24298,N_20699,N_21852);
or U24299 (N_24299,N_20092,N_20715);
xor U24300 (N_24300,N_21691,N_18920);
nor U24301 (N_24301,N_19549,N_19848);
nor U24302 (N_24302,N_19235,N_19307);
nand U24303 (N_24303,N_19209,N_19472);
xnor U24304 (N_24304,N_21429,N_19450);
nand U24305 (N_24305,N_20039,N_20968);
or U24306 (N_24306,N_20485,N_20880);
xnor U24307 (N_24307,N_18773,N_19525);
nand U24308 (N_24308,N_19520,N_20117);
or U24309 (N_24309,N_21134,N_21268);
and U24310 (N_24310,N_20595,N_20135);
nand U24311 (N_24311,N_21556,N_21297);
and U24312 (N_24312,N_19383,N_20949);
and U24313 (N_24313,N_19025,N_20954);
nand U24314 (N_24314,N_21796,N_19741);
xor U24315 (N_24315,N_21662,N_21743);
xor U24316 (N_24316,N_19124,N_21075);
nor U24317 (N_24317,N_19831,N_21172);
and U24318 (N_24318,N_18996,N_21862);
xor U24319 (N_24319,N_18829,N_21143);
nor U24320 (N_24320,N_21376,N_20751);
xor U24321 (N_24321,N_19737,N_19177);
nor U24322 (N_24322,N_20882,N_21569);
or U24323 (N_24323,N_21022,N_21783);
nor U24324 (N_24324,N_21260,N_19670);
or U24325 (N_24325,N_20623,N_20237);
nand U24326 (N_24326,N_20237,N_21042);
xor U24327 (N_24327,N_21400,N_21208);
xnor U24328 (N_24328,N_20045,N_20593);
nor U24329 (N_24329,N_19926,N_21872);
and U24330 (N_24330,N_19779,N_19724);
and U24331 (N_24331,N_20248,N_19070);
nor U24332 (N_24332,N_20161,N_20036);
xnor U24333 (N_24333,N_20435,N_21046);
nor U24334 (N_24334,N_20097,N_20544);
and U24335 (N_24335,N_19629,N_20285);
xor U24336 (N_24336,N_19565,N_18888);
nand U24337 (N_24337,N_19699,N_18933);
nor U24338 (N_24338,N_19029,N_19665);
and U24339 (N_24339,N_18793,N_19290);
and U24340 (N_24340,N_21344,N_21345);
xor U24341 (N_24341,N_19794,N_19301);
and U24342 (N_24342,N_18976,N_19028);
nor U24343 (N_24343,N_19198,N_19064);
and U24344 (N_24344,N_20652,N_21261);
or U24345 (N_24345,N_20372,N_21115);
nor U24346 (N_24346,N_19105,N_20995);
or U24347 (N_24347,N_21391,N_19544);
xor U24348 (N_24348,N_20429,N_20367);
xor U24349 (N_24349,N_19610,N_21247);
and U24350 (N_24350,N_20799,N_21228);
xor U24351 (N_24351,N_20057,N_19741);
and U24352 (N_24352,N_21843,N_19620);
nor U24353 (N_24353,N_19769,N_19159);
and U24354 (N_24354,N_21391,N_19302);
xor U24355 (N_24355,N_21777,N_21548);
or U24356 (N_24356,N_20736,N_20197);
or U24357 (N_24357,N_21423,N_19601);
xor U24358 (N_24358,N_19799,N_19931);
or U24359 (N_24359,N_19114,N_19323);
nor U24360 (N_24360,N_21753,N_20782);
and U24361 (N_24361,N_20957,N_20129);
or U24362 (N_24362,N_18855,N_20569);
xnor U24363 (N_24363,N_19867,N_20475);
nor U24364 (N_24364,N_20802,N_20942);
xor U24365 (N_24365,N_19465,N_20640);
or U24366 (N_24366,N_19260,N_20207);
nor U24367 (N_24367,N_19467,N_19510);
or U24368 (N_24368,N_19803,N_20461);
xnor U24369 (N_24369,N_20806,N_21454);
nand U24370 (N_24370,N_21390,N_20156);
nand U24371 (N_24371,N_18996,N_20990);
and U24372 (N_24372,N_19808,N_19255);
xor U24373 (N_24373,N_20535,N_20072);
and U24374 (N_24374,N_21661,N_19186);
and U24375 (N_24375,N_20112,N_19617);
xnor U24376 (N_24376,N_21444,N_21400);
or U24377 (N_24377,N_19266,N_21024);
xor U24378 (N_24378,N_21315,N_21703);
nand U24379 (N_24379,N_20902,N_21810);
and U24380 (N_24380,N_21256,N_20383);
or U24381 (N_24381,N_20959,N_18793);
and U24382 (N_24382,N_20990,N_19550);
xnor U24383 (N_24383,N_21606,N_21447);
xnor U24384 (N_24384,N_19330,N_18789);
nor U24385 (N_24385,N_20375,N_20886);
and U24386 (N_24386,N_20560,N_20733);
or U24387 (N_24387,N_20268,N_21818);
nor U24388 (N_24388,N_18926,N_18849);
nor U24389 (N_24389,N_20842,N_20699);
and U24390 (N_24390,N_21003,N_20903);
xnor U24391 (N_24391,N_20023,N_21083);
nand U24392 (N_24392,N_18770,N_20957);
nor U24393 (N_24393,N_21741,N_19450);
or U24394 (N_24394,N_19709,N_19347);
and U24395 (N_24395,N_19451,N_21619);
xnor U24396 (N_24396,N_19516,N_21047);
nor U24397 (N_24397,N_20293,N_20440);
xor U24398 (N_24398,N_21180,N_19386);
nor U24399 (N_24399,N_19690,N_21286);
nand U24400 (N_24400,N_18972,N_20052);
or U24401 (N_24401,N_19985,N_21865);
or U24402 (N_24402,N_21060,N_21247);
xor U24403 (N_24403,N_20154,N_20331);
or U24404 (N_24404,N_19355,N_21680);
or U24405 (N_24405,N_19032,N_20662);
or U24406 (N_24406,N_20842,N_20472);
xor U24407 (N_24407,N_20499,N_19375);
and U24408 (N_24408,N_19841,N_18939);
nand U24409 (N_24409,N_19301,N_19271);
and U24410 (N_24410,N_21774,N_21469);
or U24411 (N_24411,N_20223,N_21291);
and U24412 (N_24412,N_19182,N_19344);
xnor U24413 (N_24413,N_20457,N_20550);
nand U24414 (N_24414,N_21276,N_19358);
nor U24415 (N_24415,N_19379,N_20988);
or U24416 (N_24416,N_20157,N_19154);
or U24417 (N_24417,N_21615,N_19036);
nand U24418 (N_24418,N_20024,N_19846);
and U24419 (N_24419,N_19568,N_21394);
or U24420 (N_24420,N_19437,N_21573);
nand U24421 (N_24421,N_20369,N_21241);
nor U24422 (N_24422,N_19669,N_20673);
nor U24423 (N_24423,N_21325,N_19913);
or U24424 (N_24424,N_20794,N_21842);
nor U24425 (N_24425,N_21338,N_21518);
nor U24426 (N_24426,N_20858,N_19815);
or U24427 (N_24427,N_21691,N_20546);
and U24428 (N_24428,N_20483,N_18994);
xnor U24429 (N_24429,N_20662,N_21348);
or U24430 (N_24430,N_18771,N_19796);
nor U24431 (N_24431,N_19305,N_20501);
and U24432 (N_24432,N_20227,N_19427);
xnor U24433 (N_24433,N_21018,N_19913);
nor U24434 (N_24434,N_21347,N_20937);
nand U24435 (N_24435,N_19707,N_20152);
nand U24436 (N_24436,N_20689,N_21380);
nor U24437 (N_24437,N_21154,N_20659);
or U24438 (N_24438,N_21767,N_21537);
and U24439 (N_24439,N_19919,N_21396);
nand U24440 (N_24440,N_19767,N_20597);
xnor U24441 (N_24441,N_20459,N_21438);
xnor U24442 (N_24442,N_21124,N_19327);
nor U24443 (N_24443,N_21577,N_21247);
nor U24444 (N_24444,N_21075,N_19265);
nand U24445 (N_24445,N_20597,N_21656);
xor U24446 (N_24446,N_21714,N_19587);
and U24447 (N_24447,N_21471,N_19910);
xor U24448 (N_24448,N_20715,N_19856);
or U24449 (N_24449,N_21038,N_21559);
nand U24450 (N_24450,N_19264,N_19875);
and U24451 (N_24451,N_21589,N_19199);
nand U24452 (N_24452,N_21009,N_21261);
or U24453 (N_24453,N_21377,N_18894);
xnor U24454 (N_24454,N_21318,N_21193);
nor U24455 (N_24455,N_18914,N_21198);
nand U24456 (N_24456,N_21441,N_21421);
nand U24457 (N_24457,N_18828,N_19802);
or U24458 (N_24458,N_20756,N_21841);
or U24459 (N_24459,N_21868,N_19080);
nand U24460 (N_24460,N_21448,N_21336);
xor U24461 (N_24461,N_20061,N_20293);
nor U24462 (N_24462,N_20654,N_20383);
xor U24463 (N_24463,N_19211,N_21200);
nand U24464 (N_24464,N_21240,N_20296);
and U24465 (N_24465,N_20373,N_20308);
and U24466 (N_24466,N_21300,N_20530);
and U24467 (N_24467,N_20315,N_18856);
or U24468 (N_24468,N_18846,N_20290);
nor U24469 (N_24469,N_21638,N_19056);
nand U24470 (N_24470,N_20804,N_19709);
xor U24471 (N_24471,N_19400,N_20120);
xor U24472 (N_24472,N_20492,N_19817);
xor U24473 (N_24473,N_18963,N_21618);
xnor U24474 (N_24474,N_21786,N_19371);
xor U24475 (N_24475,N_20998,N_21589);
nand U24476 (N_24476,N_21096,N_20755);
nand U24477 (N_24477,N_20761,N_19693);
xor U24478 (N_24478,N_21066,N_20995);
or U24479 (N_24479,N_18767,N_21537);
nand U24480 (N_24480,N_21506,N_20325);
nor U24481 (N_24481,N_19719,N_21504);
and U24482 (N_24482,N_20197,N_21857);
xor U24483 (N_24483,N_19572,N_19432);
nand U24484 (N_24484,N_20930,N_21427);
nor U24485 (N_24485,N_20799,N_20101);
xnor U24486 (N_24486,N_20447,N_19989);
xor U24487 (N_24487,N_20930,N_19583);
nand U24488 (N_24488,N_20848,N_19961);
and U24489 (N_24489,N_19234,N_19293);
and U24490 (N_24490,N_20071,N_18844);
and U24491 (N_24491,N_21001,N_21783);
xor U24492 (N_24492,N_21587,N_19953);
or U24493 (N_24493,N_21306,N_20483);
xor U24494 (N_24494,N_20435,N_21411);
or U24495 (N_24495,N_21087,N_18966);
xnor U24496 (N_24496,N_21817,N_20361);
nand U24497 (N_24497,N_21654,N_20289);
and U24498 (N_24498,N_20568,N_19549);
and U24499 (N_24499,N_21651,N_21018);
and U24500 (N_24500,N_20493,N_19588);
nor U24501 (N_24501,N_20027,N_20670);
xnor U24502 (N_24502,N_21013,N_21649);
and U24503 (N_24503,N_21393,N_21425);
xnor U24504 (N_24504,N_19697,N_21597);
or U24505 (N_24505,N_19625,N_19023);
nand U24506 (N_24506,N_20190,N_19420);
or U24507 (N_24507,N_21388,N_19840);
or U24508 (N_24508,N_21539,N_20613);
nor U24509 (N_24509,N_20056,N_19528);
and U24510 (N_24510,N_20598,N_21790);
nor U24511 (N_24511,N_20021,N_20438);
nor U24512 (N_24512,N_20759,N_20897);
nand U24513 (N_24513,N_21451,N_19241);
and U24514 (N_24514,N_19772,N_18870);
or U24515 (N_24515,N_21834,N_19160);
xor U24516 (N_24516,N_19349,N_19049);
xnor U24517 (N_24517,N_20107,N_18791);
or U24518 (N_24518,N_18817,N_21599);
nand U24519 (N_24519,N_21473,N_19991);
nand U24520 (N_24520,N_18829,N_20981);
xor U24521 (N_24521,N_19703,N_20800);
xor U24522 (N_24522,N_20986,N_20049);
nor U24523 (N_24523,N_20744,N_19995);
or U24524 (N_24524,N_19127,N_21249);
xor U24525 (N_24525,N_18833,N_21026);
nor U24526 (N_24526,N_20484,N_21404);
nand U24527 (N_24527,N_20035,N_19326);
or U24528 (N_24528,N_20938,N_20296);
or U24529 (N_24529,N_21216,N_21707);
or U24530 (N_24530,N_20167,N_19024);
nor U24531 (N_24531,N_20074,N_19563);
nor U24532 (N_24532,N_19531,N_19265);
nor U24533 (N_24533,N_21181,N_20471);
nor U24534 (N_24534,N_20329,N_19089);
xor U24535 (N_24535,N_21334,N_19693);
and U24536 (N_24536,N_18780,N_20117);
nand U24537 (N_24537,N_18939,N_21367);
xnor U24538 (N_24538,N_20153,N_21137);
nand U24539 (N_24539,N_21490,N_21650);
nand U24540 (N_24540,N_20771,N_19092);
and U24541 (N_24541,N_20835,N_21212);
and U24542 (N_24542,N_20943,N_19629);
xnor U24543 (N_24543,N_19291,N_19236);
xnor U24544 (N_24544,N_21513,N_20442);
or U24545 (N_24545,N_19451,N_21658);
nor U24546 (N_24546,N_19664,N_20755);
or U24547 (N_24547,N_20960,N_20081);
nor U24548 (N_24548,N_20429,N_20569);
nor U24549 (N_24549,N_20653,N_19476);
xor U24550 (N_24550,N_20321,N_20003);
or U24551 (N_24551,N_20273,N_21278);
xnor U24552 (N_24552,N_21494,N_20538);
and U24553 (N_24553,N_19504,N_19597);
xor U24554 (N_24554,N_21151,N_20456);
nand U24555 (N_24555,N_20546,N_18840);
nor U24556 (N_24556,N_19671,N_19870);
or U24557 (N_24557,N_20811,N_20583);
and U24558 (N_24558,N_21153,N_21285);
nor U24559 (N_24559,N_19782,N_19517);
or U24560 (N_24560,N_20319,N_19001);
xor U24561 (N_24561,N_19899,N_21619);
nand U24562 (N_24562,N_21121,N_20390);
and U24563 (N_24563,N_18969,N_21659);
and U24564 (N_24564,N_19390,N_19584);
nand U24565 (N_24565,N_20995,N_20045);
xnor U24566 (N_24566,N_21714,N_18787);
nand U24567 (N_24567,N_20346,N_20560);
nand U24568 (N_24568,N_20217,N_20738);
nand U24569 (N_24569,N_19921,N_20804);
and U24570 (N_24570,N_21588,N_19489);
nor U24571 (N_24571,N_20242,N_21111);
xor U24572 (N_24572,N_19320,N_20235);
nand U24573 (N_24573,N_21284,N_21161);
xnor U24574 (N_24574,N_20793,N_19711);
xor U24575 (N_24575,N_20606,N_19193);
and U24576 (N_24576,N_21824,N_20559);
or U24577 (N_24577,N_19636,N_21846);
nand U24578 (N_24578,N_20374,N_20332);
xor U24579 (N_24579,N_21230,N_20913);
and U24580 (N_24580,N_20022,N_19368);
nand U24581 (N_24581,N_19404,N_19031);
and U24582 (N_24582,N_19614,N_20681);
and U24583 (N_24583,N_20397,N_20510);
xor U24584 (N_24584,N_19593,N_19898);
and U24585 (N_24585,N_20880,N_21728);
or U24586 (N_24586,N_20681,N_19344);
xor U24587 (N_24587,N_20704,N_20675);
xnor U24588 (N_24588,N_21501,N_18921);
nor U24589 (N_24589,N_19423,N_21310);
xnor U24590 (N_24590,N_19046,N_19856);
nand U24591 (N_24591,N_19207,N_19448);
nand U24592 (N_24592,N_19477,N_18942);
nor U24593 (N_24593,N_21334,N_19686);
nor U24594 (N_24594,N_20935,N_21076);
nor U24595 (N_24595,N_21168,N_19039);
or U24596 (N_24596,N_21717,N_20523);
and U24597 (N_24597,N_19012,N_18794);
nor U24598 (N_24598,N_19774,N_21465);
nor U24599 (N_24599,N_20211,N_20634);
xor U24600 (N_24600,N_21195,N_18762);
xnor U24601 (N_24601,N_19171,N_20678);
and U24602 (N_24602,N_20531,N_21140);
xnor U24603 (N_24603,N_19319,N_21661);
nor U24604 (N_24604,N_20569,N_21780);
or U24605 (N_24605,N_21466,N_19681);
nor U24606 (N_24606,N_19240,N_19163);
or U24607 (N_24607,N_20196,N_21499);
and U24608 (N_24608,N_20812,N_21832);
and U24609 (N_24609,N_19846,N_19175);
nand U24610 (N_24610,N_20944,N_18786);
and U24611 (N_24611,N_19776,N_20392);
and U24612 (N_24612,N_19407,N_21344);
nor U24613 (N_24613,N_21865,N_19525);
nand U24614 (N_24614,N_20084,N_20446);
nand U24615 (N_24615,N_19124,N_20944);
and U24616 (N_24616,N_19267,N_20170);
nor U24617 (N_24617,N_21743,N_18885);
and U24618 (N_24618,N_21785,N_18854);
nor U24619 (N_24619,N_18960,N_21701);
or U24620 (N_24620,N_21642,N_21673);
nand U24621 (N_24621,N_19058,N_19317);
or U24622 (N_24622,N_18865,N_20874);
and U24623 (N_24623,N_19489,N_20437);
nand U24624 (N_24624,N_21465,N_21814);
nand U24625 (N_24625,N_20984,N_21843);
and U24626 (N_24626,N_19582,N_20795);
nand U24627 (N_24627,N_21729,N_21140);
and U24628 (N_24628,N_20768,N_20849);
nor U24629 (N_24629,N_20860,N_21708);
nor U24630 (N_24630,N_20284,N_20320);
and U24631 (N_24631,N_19109,N_21699);
nor U24632 (N_24632,N_18783,N_21252);
or U24633 (N_24633,N_21256,N_20344);
nor U24634 (N_24634,N_19775,N_21797);
nand U24635 (N_24635,N_19397,N_19356);
xor U24636 (N_24636,N_20321,N_20435);
and U24637 (N_24637,N_19615,N_20017);
or U24638 (N_24638,N_19599,N_21449);
or U24639 (N_24639,N_21175,N_19328);
and U24640 (N_24640,N_21095,N_18767);
xnor U24641 (N_24641,N_20607,N_20004);
xor U24642 (N_24642,N_21147,N_20018);
or U24643 (N_24643,N_19678,N_20934);
nand U24644 (N_24644,N_18865,N_21046);
nand U24645 (N_24645,N_21491,N_19452);
nand U24646 (N_24646,N_20270,N_19119);
and U24647 (N_24647,N_20443,N_20993);
xor U24648 (N_24648,N_21803,N_19559);
and U24649 (N_24649,N_21396,N_20669);
or U24650 (N_24650,N_21421,N_19034);
or U24651 (N_24651,N_20924,N_19819);
xor U24652 (N_24652,N_20570,N_21172);
and U24653 (N_24653,N_21625,N_21322);
or U24654 (N_24654,N_20984,N_19708);
nor U24655 (N_24655,N_20949,N_21417);
or U24656 (N_24656,N_19325,N_18846);
xor U24657 (N_24657,N_18818,N_21214);
nand U24658 (N_24658,N_19038,N_19145);
nand U24659 (N_24659,N_21059,N_19178);
nand U24660 (N_24660,N_20808,N_19670);
nand U24661 (N_24661,N_19829,N_20922);
and U24662 (N_24662,N_20969,N_21232);
and U24663 (N_24663,N_20124,N_19292);
nor U24664 (N_24664,N_20996,N_20810);
xnor U24665 (N_24665,N_18940,N_19859);
nand U24666 (N_24666,N_21718,N_21830);
xor U24667 (N_24667,N_20045,N_20906);
or U24668 (N_24668,N_20085,N_19494);
or U24669 (N_24669,N_19736,N_21402);
xnor U24670 (N_24670,N_18879,N_20865);
or U24671 (N_24671,N_21556,N_20010);
and U24672 (N_24672,N_19944,N_19383);
or U24673 (N_24673,N_20202,N_19613);
xor U24674 (N_24674,N_19507,N_18765);
or U24675 (N_24675,N_19383,N_20868);
xnor U24676 (N_24676,N_19104,N_19266);
xor U24677 (N_24677,N_20490,N_21252);
or U24678 (N_24678,N_19103,N_20381);
and U24679 (N_24679,N_20136,N_19653);
nor U24680 (N_24680,N_18860,N_19166);
nand U24681 (N_24681,N_20873,N_20459);
and U24682 (N_24682,N_19432,N_20070);
or U24683 (N_24683,N_21564,N_19826);
nor U24684 (N_24684,N_20813,N_21413);
nor U24685 (N_24685,N_20054,N_21149);
xor U24686 (N_24686,N_20393,N_20755);
xor U24687 (N_24687,N_19851,N_19920);
or U24688 (N_24688,N_19058,N_20938);
and U24689 (N_24689,N_20031,N_20230);
and U24690 (N_24690,N_20323,N_19440);
or U24691 (N_24691,N_18860,N_19341);
nor U24692 (N_24692,N_21425,N_20006);
nand U24693 (N_24693,N_19246,N_21321);
or U24694 (N_24694,N_20289,N_19028);
nor U24695 (N_24695,N_19235,N_20878);
and U24696 (N_24696,N_21136,N_21733);
xor U24697 (N_24697,N_19039,N_20573);
nand U24698 (N_24698,N_21160,N_20908);
or U24699 (N_24699,N_19987,N_21251);
or U24700 (N_24700,N_19603,N_21562);
and U24701 (N_24701,N_19117,N_20407);
xnor U24702 (N_24702,N_19761,N_20940);
nor U24703 (N_24703,N_20061,N_20209);
and U24704 (N_24704,N_20668,N_20434);
nand U24705 (N_24705,N_21274,N_19125);
nor U24706 (N_24706,N_21050,N_18926);
nand U24707 (N_24707,N_19797,N_21537);
xnor U24708 (N_24708,N_19776,N_18801);
nand U24709 (N_24709,N_19155,N_20241);
nor U24710 (N_24710,N_21731,N_21873);
nand U24711 (N_24711,N_20410,N_21859);
or U24712 (N_24712,N_20095,N_19877);
and U24713 (N_24713,N_20514,N_21666);
xnor U24714 (N_24714,N_20264,N_21382);
xor U24715 (N_24715,N_20652,N_21273);
and U24716 (N_24716,N_20148,N_19228);
nor U24717 (N_24717,N_18756,N_19728);
nand U24718 (N_24718,N_20957,N_18880);
xor U24719 (N_24719,N_18852,N_20589);
or U24720 (N_24720,N_20001,N_20515);
and U24721 (N_24721,N_20003,N_20179);
or U24722 (N_24722,N_20545,N_18928);
and U24723 (N_24723,N_20427,N_21681);
xnor U24724 (N_24724,N_19736,N_18773);
xor U24725 (N_24725,N_19885,N_21572);
nor U24726 (N_24726,N_21540,N_19020);
and U24727 (N_24727,N_21003,N_20404);
or U24728 (N_24728,N_21752,N_19391);
nand U24729 (N_24729,N_20317,N_19362);
and U24730 (N_24730,N_19491,N_19661);
xor U24731 (N_24731,N_20378,N_18816);
nor U24732 (N_24732,N_19260,N_21575);
or U24733 (N_24733,N_21774,N_21088);
nor U24734 (N_24734,N_20331,N_19994);
or U24735 (N_24735,N_19566,N_21115);
nor U24736 (N_24736,N_20194,N_21133);
or U24737 (N_24737,N_21662,N_20286);
nor U24738 (N_24738,N_19995,N_21592);
xnor U24739 (N_24739,N_21593,N_19104);
or U24740 (N_24740,N_19951,N_19703);
nor U24741 (N_24741,N_21413,N_19973);
or U24742 (N_24742,N_21377,N_21383);
xor U24743 (N_24743,N_21337,N_20085);
and U24744 (N_24744,N_19608,N_20171);
nand U24745 (N_24745,N_20825,N_20324);
or U24746 (N_24746,N_21532,N_19700);
xor U24747 (N_24747,N_19761,N_19975);
nor U24748 (N_24748,N_19059,N_21133);
xnor U24749 (N_24749,N_20887,N_19990);
xor U24750 (N_24750,N_19269,N_21394);
nor U24751 (N_24751,N_19663,N_21462);
nor U24752 (N_24752,N_18846,N_20434);
or U24753 (N_24753,N_20750,N_20276);
nor U24754 (N_24754,N_21659,N_20207);
and U24755 (N_24755,N_20602,N_21110);
nand U24756 (N_24756,N_21605,N_20040);
nor U24757 (N_24757,N_20361,N_20112);
nor U24758 (N_24758,N_19652,N_19666);
xnor U24759 (N_24759,N_20260,N_21806);
or U24760 (N_24760,N_21076,N_20525);
nand U24761 (N_24761,N_18847,N_18960);
or U24762 (N_24762,N_20041,N_21749);
xor U24763 (N_24763,N_20626,N_19255);
nand U24764 (N_24764,N_21807,N_21017);
nand U24765 (N_24765,N_19887,N_20710);
nand U24766 (N_24766,N_21283,N_18861);
or U24767 (N_24767,N_19720,N_19079);
nor U24768 (N_24768,N_20428,N_20963);
nor U24769 (N_24769,N_19944,N_18976);
and U24770 (N_24770,N_19184,N_19397);
or U24771 (N_24771,N_19376,N_18767);
and U24772 (N_24772,N_21459,N_19231);
nor U24773 (N_24773,N_19878,N_19448);
or U24774 (N_24774,N_21586,N_19800);
or U24775 (N_24775,N_19738,N_18867);
xor U24776 (N_24776,N_18768,N_19241);
xor U24777 (N_24777,N_18847,N_21629);
xor U24778 (N_24778,N_19271,N_20246);
nand U24779 (N_24779,N_20802,N_21633);
nor U24780 (N_24780,N_20344,N_19954);
or U24781 (N_24781,N_19312,N_19142);
and U24782 (N_24782,N_21695,N_20497);
xnor U24783 (N_24783,N_20325,N_18929);
and U24784 (N_24784,N_20657,N_19446);
nand U24785 (N_24785,N_20826,N_19534);
nor U24786 (N_24786,N_20354,N_20693);
and U24787 (N_24787,N_19096,N_19204);
or U24788 (N_24788,N_20626,N_20508);
xor U24789 (N_24789,N_20849,N_19925);
nor U24790 (N_24790,N_21478,N_19114);
nor U24791 (N_24791,N_20417,N_20892);
or U24792 (N_24792,N_20887,N_19300);
or U24793 (N_24793,N_20451,N_19550);
or U24794 (N_24794,N_19232,N_20262);
nor U24795 (N_24795,N_21838,N_18969);
xnor U24796 (N_24796,N_19760,N_19706);
nor U24797 (N_24797,N_20213,N_19976);
xnor U24798 (N_24798,N_21447,N_19777);
or U24799 (N_24799,N_20800,N_19611);
or U24800 (N_24800,N_19941,N_21290);
and U24801 (N_24801,N_20053,N_20844);
nand U24802 (N_24802,N_19202,N_21088);
nor U24803 (N_24803,N_20675,N_21338);
nand U24804 (N_24804,N_21747,N_21474);
xnor U24805 (N_24805,N_19717,N_21739);
nor U24806 (N_24806,N_18784,N_20975);
nor U24807 (N_24807,N_20807,N_19719);
and U24808 (N_24808,N_21613,N_20075);
nor U24809 (N_24809,N_21235,N_19424);
nand U24810 (N_24810,N_21165,N_20999);
nor U24811 (N_24811,N_19166,N_21753);
nor U24812 (N_24812,N_19956,N_21170);
and U24813 (N_24813,N_20593,N_19646);
xnor U24814 (N_24814,N_19687,N_18917);
nor U24815 (N_24815,N_19385,N_19119);
xor U24816 (N_24816,N_20765,N_19158);
nand U24817 (N_24817,N_21596,N_19317);
xnor U24818 (N_24818,N_20286,N_20894);
nor U24819 (N_24819,N_19634,N_19386);
nand U24820 (N_24820,N_19956,N_21346);
xor U24821 (N_24821,N_20031,N_19616);
nand U24822 (N_24822,N_20809,N_20340);
or U24823 (N_24823,N_19388,N_20160);
xor U24824 (N_24824,N_19817,N_21277);
or U24825 (N_24825,N_19255,N_20576);
nand U24826 (N_24826,N_20545,N_19322);
xnor U24827 (N_24827,N_21792,N_18853);
nor U24828 (N_24828,N_19591,N_19466);
nor U24829 (N_24829,N_21595,N_21273);
or U24830 (N_24830,N_19606,N_19669);
or U24831 (N_24831,N_18983,N_20862);
nor U24832 (N_24832,N_20363,N_21690);
or U24833 (N_24833,N_19592,N_20772);
or U24834 (N_24834,N_21286,N_18833);
and U24835 (N_24835,N_20908,N_18830);
or U24836 (N_24836,N_20859,N_20808);
and U24837 (N_24837,N_21422,N_20864);
and U24838 (N_24838,N_18887,N_21669);
and U24839 (N_24839,N_19792,N_20276);
xor U24840 (N_24840,N_19121,N_20717);
and U24841 (N_24841,N_21276,N_21082);
nand U24842 (N_24842,N_20141,N_21571);
and U24843 (N_24843,N_19106,N_19280);
and U24844 (N_24844,N_20767,N_20721);
nor U24845 (N_24845,N_20407,N_19163);
or U24846 (N_24846,N_20241,N_21733);
xor U24847 (N_24847,N_20273,N_21036);
nor U24848 (N_24848,N_21581,N_20811);
nor U24849 (N_24849,N_21004,N_19866);
nor U24850 (N_24850,N_19935,N_19090);
xor U24851 (N_24851,N_19269,N_21611);
nor U24852 (N_24852,N_20882,N_20020);
nor U24853 (N_24853,N_20702,N_20213);
nand U24854 (N_24854,N_21150,N_20827);
nand U24855 (N_24855,N_19248,N_20466);
nand U24856 (N_24856,N_19960,N_19528);
and U24857 (N_24857,N_20881,N_18948);
nor U24858 (N_24858,N_20432,N_20825);
nor U24859 (N_24859,N_21180,N_20331);
and U24860 (N_24860,N_19847,N_20396);
xnor U24861 (N_24861,N_20691,N_19619);
or U24862 (N_24862,N_19598,N_21100);
or U24863 (N_24863,N_21765,N_20467);
xnor U24864 (N_24864,N_20303,N_18754);
nor U24865 (N_24865,N_19139,N_18929);
nand U24866 (N_24866,N_21784,N_21667);
and U24867 (N_24867,N_20706,N_20423);
xor U24868 (N_24868,N_21112,N_21060);
nand U24869 (N_24869,N_19664,N_20387);
xnor U24870 (N_24870,N_19421,N_20979);
xnor U24871 (N_24871,N_19644,N_19707);
nor U24872 (N_24872,N_19824,N_19851);
and U24873 (N_24873,N_19302,N_18972);
and U24874 (N_24874,N_19198,N_19999);
and U24875 (N_24875,N_19987,N_19902);
and U24876 (N_24876,N_20843,N_20891);
nor U24877 (N_24877,N_19485,N_19395);
nor U24878 (N_24878,N_20835,N_21765);
or U24879 (N_24879,N_19656,N_20992);
or U24880 (N_24880,N_19228,N_20376);
or U24881 (N_24881,N_19641,N_19396);
or U24882 (N_24882,N_20354,N_20570);
and U24883 (N_24883,N_19857,N_18927);
nor U24884 (N_24884,N_19430,N_19230);
nand U24885 (N_24885,N_20592,N_21140);
xor U24886 (N_24886,N_20282,N_20688);
xnor U24887 (N_24887,N_21247,N_21386);
nor U24888 (N_24888,N_18957,N_19345);
or U24889 (N_24889,N_20036,N_19477);
or U24890 (N_24890,N_19784,N_19042);
nand U24891 (N_24891,N_20786,N_19461);
and U24892 (N_24892,N_18821,N_18780);
or U24893 (N_24893,N_20989,N_19208);
nor U24894 (N_24894,N_19822,N_20694);
or U24895 (N_24895,N_20092,N_20731);
or U24896 (N_24896,N_21317,N_19301);
or U24897 (N_24897,N_19320,N_19652);
nand U24898 (N_24898,N_21160,N_21564);
and U24899 (N_24899,N_21304,N_21471);
nand U24900 (N_24900,N_21397,N_21752);
nand U24901 (N_24901,N_20108,N_20037);
xor U24902 (N_24902,N_19348,N_21152);
nor U24903 (N_24903,N_19776,N_19117);
nand U24904 (N_24904,N_19815,N_21486);
xnor U24905 (N_24905,N_20035,N_19948);
nor U24906 (N_24906,N_20565,N_20023);
nor U24907 (N_24907,N_19012,N_19844);
nand U24908 (N_24908,N_20062,N_19392);
xnor U24909 (N_24909,N_21358,N_20769);
nand U24910 (N_24910,N_21597,N_20184);
nand U24911 (N_24911,N_19278,N_20238);
nor U24912 (N_24912,N_19975,N_21216);
and U24913 (N_24913,N_21685,N_19750);
nand U24914 (N_24914,N_20636,N_21781);
nand U24915 (N_24915,N_21366,N_19114);
and U24916 (N_24916,N_20460,N_20684);
and U24917 (N_24917,N_19847,N_20862);
and U24918 (N_24918,N_19808,N_19322);
nor U24919 (N_24919,N_20281,N_20389);
nor U24920 (N_24920,N_21738,N_21079);
or U24921 (N_24921,N_19411,N_20041);
and U24922 (N_24922,N_21279,N_21403);
xor U24923 (N_24923,N_18967,N_20058);
nor U24924 (N_24924,N_20661,N_20714);
nor U24925 (N_24925,N_19401,N_20857);
and U24926 (N_24926,N_19488,N_20590);
nand U24927 (N_24927,N_20753,N_21836);
nand U24928 (N_24928,N_21685,N_19669);
and U24929 (N_24929,N_20963,N_21372);
nor U24930 (N_24930,N_19273,N_19957);
and U24931 (N_24931,N_19195,N_19588);
nor U24932 (N_24932,N_21774,N_19762);
nand U24933 (N_24933,N_21684,N_19599);
nand U24934 (N_24934,N_19914,N_20262);
nand U24935 (N_24935,N_19979,N_21033);
nand U24936 (N_24936,N_20168,N_20368);
nor U24937 (N_24937,N_21296,N_21567);
xor U24938 (N_24938,N_19971,N_20990);
or U24939 (N_24939,N_19951,N_20244);
nand U24940 (N_24940,N_19428,N_20062);
xor U24941 (N_24941,N_18757,N_18995);
xor U24942 (N_24942,N_19979,N_21536);
nor U24943 (N_24943,N_21088,N_19667);
or U24944 (N_24944,N_21538,N_19084);
or U24945 (N_24945,N_19013,N_21205);
and U24946 (N_24946,N_20359,N_18966);
nor U24947 (N_24947,N_19471,N_19490);
nor U24948 (N_24948,N_20333,N_18894);
nand U24949 (N_24949,N_19346,N_21405);
xor U24950 (N_24950,N_20357,N_20942);
and U24951 (N_24951,N_21088,N_19722);
and U24952 (N_24952,N_21820,N_19901);
nor U24953 (N_24953,N_21510,N_20309);
nor U24954 (N_24954,N_18993,N_20911);
nand U24955 (N_24955,N_19508,N_20571);
or U24956 (N_24956,N_21816,N_19193);
xnor U24957 (N_24957,N_19662,N_21763);
nor U24958 (N_24958,N_20006,N_20848);
nand U24959 (N_24959,N_21562,N_20949);
xor U24960 (N_24960,N_20392,N_19390);
and U24961 (N_24961,N_21363,N_19632);
or U24962 (N_24962,N_20614,N_21453);
nor U24963 (N_24963,N_18920,N_19405);
xnor U24964 (N_24964,N_20951,N_20613);
or U24965 (N_24965,N_19476,N_20863);
nand U24966 (N_24966,N_19328,N_21675);
nor U24967 (N_24967,N_20879,N_18904);
xor U24968 (N_24968,N_21807,N_19978);
or U24969 (N_24969,N_18846,N_20084);
and U24970 (N_24970,N_19313,N_21114);
nand U24971 (N_24971,N_20663,N_19155);
and U24972 (N_24972,N_20563,N_21481);
or U24973 (N_24973,N_20198,N_21597);
or U24974 (N_24974,N_20338,N_20566);
nor U24975 (N_24975,N_20353,N_20312);
xor U24976 (N_24976,N_19540,N_21606);
and U24977 (N_24977,N_20174,N_20317);
nor U24978 (N_24978,N_19149,N_21271);
nand U24979 (N_24979,N_19798,N_19136);
and U24980 (N_24980,N_21731,N_20943);
xor U24981 (N_24981,N_20221,N_20240);
nor U24982 (N_24982,N_19712,N_20137);
nor U24983 (N_24983,N_21651,N_20127);
or U24984 (N_24984,N_20745,N_21050);
or U24985 (N_24985,N_21187,N_19474);
nor U24986 (N_24986,N_19852,N_20894);
and U24987 (N_24987,N_20269,N_21719);
nand U24988 (N_24988,N_21273,N_20545);
xor U24989 (N_24989,N_19011,N_21846);
nand U24990 (N_24990,N_20108,N_21299);
xor U24991 (N_24991,N_20141,N_20948);
nand U24992 (N_24992,N_21166,N_19946);
nand U24993 (N_24993,N_19448,N_20603);
nor U24994 (N_24994,N_19932,N_19072);
nor U24995 (N_24995,N_21833,N_19855);
or U24996 (N_24996,N_21259,N_21356);
xnor U24997 (N_24997,N_19100,N_20694);
xor U24998 (N_24998,N_20758,N_19035);
nand U24999 (N_24999,N_19063,N_20362);
or UO_0 (O_0,N_23582,N_22810);
and UO_1 (O_1,N_24190,N_22462);
or UO_2 (O_2,N_22246,N_24506);
nand UO_3 (O_3,N_23481,N_22606);
or UO_4 (O_4,N_24534,N_24782);
and UO_5 (O_5,N_23544,N_24995);
nand UO_6 (O_6,N_23320,N_23463);
nand UO_7 (O_7,N_24587,N_22902);
and UO_8 (O_8,N_22146,N_24830);
and UO_9 (O_9,N_23881,N_23500);
nor UO_10 (O_10,N_24721,N_23900);
nor UO_11 (O_11,N_23236,N_23842);
xnor UO_12 (O_12,N_21938,N_23394);
nand UO_13 (O_13,N_24529,N_22262);
xor UO_14 (O_14,N_22743,N_23462);
or UO_15 (O_15,N_23848,N_23209);
xnor UO_16 (O_16,N_22782,N_23343);
nand UO_17 (O_17,N_22125,N_22927);
or UO_18 (O_18,N_22896,N_23936);
nor UO_19 (O_19,N_23257,N_24516);
or UO_20 (O_20,N_22417,N_22383);
nand UO_21 (O_21,N_24521,N_24872);
or UO_22 (O_22,N_22047,N_22270);
nand UO_23 (O_23,N_24320,N_24442);
or UO_24 (O_24,N_22536,N_22430);
xor UO_25 (O_25,N_22991,N_23303);
nor UO_26 (O_26,N_23680,N_23069);
nand UO_27 (O_27,N_23461,N_22769);
nand UO_28 (O_28,N_24776,N_24917);
nor UO_29 (O_29,N_23150,N_22284);
nand UO_30 (O_30,N_24852,N_22106);
nor UO_31 (O_31,N_23846,N_22660);
or UO_32 (O_32,N_23888,N_22195);
xor UO_33 (O_33,N_22238,N_23005);
nand UO_34 (O_34,N_23415,N_22551);
or UO_35 (O_35,N_24282,N_24208);
nand UO_36 (O_36,N_22711,N_21988);
nor UO_37 (O_37,N_24079,N_23068);
xnor UO_38 (O_38,N_24615,N_24233);
nor UO_39 (O_39,N_21926,N_24429);
xor UO_40 (O_40,N_24346,N_24561);
or UO_41 (O_41,N_22547,N_23824);
nand UO_42 (O_42,N_24179,N_23245);
nor UO_43 (O_43,N_22318,N_24310);
xor UO_44 (O_44,N_23490,N_24185);
xnor UO_45 (O_45,N_23008,N_22103);
nor UO_46 (O_46,N_22577,N_23982);
nor UO_47 (O_47,N_23189,N_22385);
nand UO_48 (O_48,N_23618,N_22903);
or UO_49 (O_49,N_23976,N_23720);
nand UO_50 (O_50,N_23272,N_23965);
nor UO_51 (O_51,N_24189,N_24243);
nand UO_52 (O_52,N_24101,N_24726);
or UO_53 (O_53,N_22818,N_23221);
nand UO_54 (O_54,N_24862,N_22064);
and UO_55 (O_55,N_23015,N_23104);
or UO_56 (O_56,N_22330,N_24971);
or UO_57 (O_57,N_21995,N_23191);
xnor UO_58 (O_58,N_22232,N_23917);
and UO_59 (O_59,N_24137,N_22035);
nand UO_60 (O_60,N_22770,N_22981);
or UO_61 (O_61,N_23157,N_23469);
and UO_62 (O_62,N_22832,N_21900);
nand UO_63 (O_63,N_24009,N_24713);
and UO_64 (O_64,N_24296,N_23673);
or UO_65 (O_65,N_21908,N_23143);
xor UO_66 (O_66,N_22940,N_24412);
or UO_67 (O_67,N_23716,N_23704);
and UO_68 (O_68,N_23187,N_22227);
xnor UO_69 (O_69,N_22575,N_24930);
nor UO_70 (O_70,N_23207,N_23766);
or UO_71 (O_71,N_22984,N_24178);
nand UO_72 (O_72,N_22290,N_23280);
and UO_73 (O_73,N_22358,N_22972);
or UO_74 (O_74,N_24280,N_23670);
xnor UO_75 (O_75,N_23374,N_23470);
or UO_76 (O_76,N_22544,N_24460);
nor UO_77 (O_77,N_23373,N_22507);
nor UO_78 (O_78,N_22697,N_24955);
nor UO_79 (O_79,N_24389,N_22826);
nand UO_80 (O_80,N_22578,N_22734);
nor UO_81 (O_81,N_23416,N_23893);
xnor UO_82 (O_82,N_24559,N_24375);
xnor UO_83 (O_83,N_24263,N_21897);
xor UO_84 (O_84,N_23682,N_24738);
nand UO_85 (O_85,N_22677,N_22167);
and UO_86 (O_86,N_22944,N_23379);
xor UO_87 (O_87,N_23498,N_23139);
and UO_88 (O_88,N_23492,N_22432);
nor UO_89 (O_89,N_21940,N_23903);
or UO_90 (O_90,N_23753,N_21875);
nand UO_91 (O_91,N_24600,N_22532);
nor UO_92 (O_92,N_23614,N_23386);
nor UO_93 (O_93,N_24783,N_23696);
nand UO_94 (O_94,N_22825,N_23654);
and UO_95 (O_95,N_24291,N_24476);
or UO_96 (O_96,N_22219,N_23183);
nand UO_97 (O_97,N_24126,N_24212);
xnor UO_98 (O_98,N_24624,N_22929);
nor UO_99 (O_99,N_24834,N_22965);
and UO_100 (O_100,N_23140,N_24452);
or UO_101 (O_101,N_23075,N_22584);
or UO_102 (O_102,N_23676,N_22579);
and UO_103 (O_103,N_22007,N_23464);
nor UO_104 (O_104,N_22654,N_22692);
xor UO_105 (O_105,N_22977,N_24984);
nor UO_106 (O_106,N_24882,N_23220);
nor UO_107 (O_107,N_23884,N_22211);
and UO_108 (O_108,N_24215,N_23545);
xnor UO_109 (O_109,N_24145,N_22558);
nand UO_110 (O_110,N_24149,N_22694);
nor UO_111 (O_111,N_22500,N_21960);
or UO_112 (O_112,N_23080,N_23963);
nand UO_113 (O_113,N_23843,N_24261);
and UO_114 (O_114,N_22687,N_22244);
and UO_115 (O_115,N_23851,N_24068);
nand UO_116 (O_116,N_23569,N_23083);
nand UO_117 (O_117,N_23214,N_22312);
nor UO_118 (O_118,N_24949,N_22172);
or UO_119 (O_119,N_24863,N_24592);
nand UO_120 (O_120,N_22588,N_22175);
and UO_121 (O_121,N_23732,N_22846);
and UO_122 (O_122,N_23467,N_24259);
or UO_123 (O_123,N_23125,N_23928);
nand UO_124 (O_124,N_23459,N_24449);
or UO_125 (O_125,N_24200,N_23230);
or UO_126 (O_126,N_23951,N_24118);
and UO_127 (O_127,N_24318,N_23318);
and UO_128 (O_128,N_23381,N_24403);
nand UO_129 (O_129,N_24766,N_22519);
nor UO_130 (O_130,N_23938,N_22080);
or UO_131 (O_131,N_21924,N_22627);
nor UO_132 (O_132,N_23637,N_24251);
and UO_133 (O_133,N_24000,N_24513);
and UO_134 (O_134,N_24342,N_23810);
nand UO_135 (O_135,N_24509,N_22024);
or UO_136 (O_136,N_22072,N_24434);
nor UO_137 (O_137,N_22961,N_24255);
and UO_138 (O_138,N_24678,N_22267);
xor UO_139 (O_139,N_24531,N_22530);
nor UO_140 (O_140,N_22163,N_23899);
nor UO_141 (O_141,N_23585,N_22774);
and UO_142 (O_142,N_24848,N_24708);
xor UO_143 (O_143,N_24657,N_23663);
xor UO_144 (O_144,N_24188,N_23697);
and UO_145 (O_145,N_22276,N_23588);
nand UO_146 (O_146,N_22404,N_23348);
nand UO_147 (O_147,N_22116,N_23085);
or UO_148 (O_148,N_24821,N_23011);
nor UO_149 (O_149,N_22650,N_22835);
xnor UO_150 (O_150,N_23042,N_22434);
and UO_151 (O_151,N_22552,N_24025);
or UO_152 (O_152,N_24889,N_23939);
and UO_153 (O_153,N_23361,N_23084);
or UO_154 (O_154,N_22523,N_24567);
or UO_155 (O_155,N_24565,N_24809);
and UO_156 (O_156,N_22114,N_24638);
or UO_157 (O_157,N_24787,N_24269);
and UO_158 (O_158,N_24680,N_24104);
or UO_159 (O_159,N_23460,N_23602);
nor UO_160 (O_160,N_24835,N_22772);
nor UO_161 (O_161,N_24242,N_24329);
xor UO_162 (O_162,N_24122,N_24309);
nand UO_163 (O_163,N_22804,N_22973);
xnor UO_164 (O_164,N_22733,N_22741);
nand UO_165 (O_165,N_22824,N_21886);
nand UO_166 (O_166,N_22298,N_22620);
xor UO_167 (O_167,N_24945,N_23310);
and UO_168 (O_168,N_23642,N_23273);
or UO_169 (O_169,N_22648,N_22429);
or UO_170 (O_170,N_24577,N_23550);
nor UO_171 (O_171,N_22535,N_22022);
nand UO_172 (O_172,N_22249,N_24351);
nor UO_173 (O_173,N_23611,N_22468);
xor UO_174 (O_174,N_24336,N_21957);
or UO_175 (O_175,N_23711,N_23222);
or UO_176 (O_176,N_23816,N_23919);
xnor UO_177 (O_177,N_23797,N_22135);
nor UO_178 (O_178,N_21891,N_22196);
nor UO_179 (O_179,N_22967,N_22340);
and UO_180 (O_180,N_22941,N_21992);
nand UO_181 (O_181,N_22985,N_22548);
xor UO_182 (O_182,N_23118,N_24605);
nand UO_183 (O_183,N_23541,N_21906);
xor UO_184 (O_184,N_22518,N_24213);
xnor UO_185 (O_185,N_22722,N_24560);
or UO_186 (O_186,N_23163,N_24530);
nor UO_187 (O_187,N_24732,N_24859);
and UO_188 (O_188,N_22631,N_22142);
nor UO_189 (O_189,N_23981,N_22726);
nand UO_190 (O_190,N_23448,N_24793);
or UO_191 (O_191,N_23531,N_23185);
nand UO_192 (O_192,N_24866,N_22626);
nand UO_193 (O_193,N_22268,N_22282);
xnor UO_194 (O_194,N_24341,N_23046);
and UO_195 (O_195,N_23941,N_23340);
or UO_196 (O_196,N_24688,N_24220);
and UO_197 (O_197,N_24512,N_24537);
nand UO_198 (O_198,N_22107,N_24883);
or UO_199 (O_199,N_22714,N_24231);
nand UO_200 (O_200,N_23645,N_23154);
and UO_201 (O_201,N_22870,N_23420);
nand UO_202 (O_202,N_24719,N_22971);
and UO_203 (O_203,N_24723,N_24966);
and UO_204 (O_204,N_24675,N_22785);
xor UO_205 (O_205,N_24614,N_24880);
nand UO_206 (O_206,N_24364,N_22592);
nand UO_207 (O_207,N_24191,N_22455);
or UO_208 (O_208,N_23718,N_22031);
xnor UO_209 (O_209,N_22236,N_22173);
xor UO_210 (O_210,N_23418,N_24858);
nor UO_211 (O_211,N_24897,N_21981);
or UO_212 (O_212,N_22052,N_24217);
xnor UO_213 (O_213,N_24132,N_22964);
or UO_214 (O_214,N_22789,N_23999);
nand UO_215 (O_215,N_23218,N_24324);
nor UO_216 (O_216,N_23813,N_23484);
xor UO_217 (O_217,N_23653,N_23891);
nand UO_218 (O_218,N_24832,N_23821);
nor UO_219 (O_219,N_24352,N_22093);
or UO_220 (O_220,N_24807,N_24919);
or UO_221 (O_221,N_23300,N_24963);
nor UO_222 (O_222,N_24979,N_22460);
nand UO_223 (O_223,N_22729,N_24472);
nor UO_224 (O_224,N_22229,N_23054);
or UO_225 (O_225,N_21882,N_24580);
and UO_226 (O_226,N_23306,N_24900);
xor UO_227 (O_227,N_22091,N_24302);
and UO_228 (O_228,N_24174,N_24968);
nor UO_229 (O_229,N_24443,N_23477);
and UO_230 (O_230,N_22360,N_23354);
and UO_231 (O_231,N_24824,N_24958);
xor UO_232 (O_232,N_22564,N_23003);
and UO_233 (O_233,N_22038,N_22086);
xnor UO_234 (O_234,N_22928,N_22416);
xor UO_235 (O_235,N_24760,N_22843);
or UO_236 (O_236,N_24368,N_24609);
xnor UO_237 (O_237,N_24112,N_22593);
nand UO_238 (O_238,N_23093,N_23495);
nor UO_239 (O_239,N_22997,N_23170);
xor UO_240 (O_240,N_24151,N_24102);
and UO_241 (O_241,N_24353,N_22683);
and UO_242 (O_242,N_22557,N_23609);
xor UO_243 (O_243,N_23114,N_23436);
nor UO_244 (O_244,N_21979,N_23124);
nor UO_245 (O_245,N_24855,N_24991);
and UO_246 (O_246,N_23922,N_24998);
xor UO_247 (O_247,N_24407,N_24182);
and UO_248 (O_248,N_21953,N_24669);
xor UO_249 (O_249,N_21969,N_24652);
xnor UO_250 (O_250,N_23782,N_24608);
nor UO_251 (O_251,N_22983,N_23615);
xnor UO_252 (O_252,N_24907,N_24402);
or UO_253 (O_253,N_23423,N_22018);
nor UO_254 (O_254,N_22866,N_23521);
nor UO_255 (O_255,N_22303,N_24475);
nand UO_256 (O_256,N_24306,N_23535);
and UO_257 (O_257,N_22077,N_22419);
or UO_258 (O_258,N_23253,N_22780);
or UO_259 (O_259,N_22841,N_23362);
xor UO_260 (O_260,N_22747,N_23442);
nor UO_261 (O_261,N_22094,N_22757);
and UO_262 (O_262,N_23540,N_22682);
or UO_263 (O_263,N_24797,N_23587);
or UO_264 (O_264,N_23341,N_23962);
and UO_265 (O_265,N_22555,N_24695);
nand UO_266 (O_266,N_22292,N_23800);
xor UO_267 (O_267,N_24021,N_22712);
nand UO_268 (O_268,N_23978,N_23431);
nor UO_269 (O_269,N_23687,N_23798);
xnor UO_270 (O_270,N_22897,N_22815);
and UO_271 (O_271,N_24316,N_24439);
or UO_272 (O_272,N_22100,N_22321);
nand UO_273 (O_273,N_23038,N_24946);
and UO_274 (O_274,N_22124,N_23561);
nor UO_275 (O_275,N_22127,N_22475);
nor UO_276 (O_276,N_24494,N_23413);
xor UO_277 (O_277,N_24195,N_22139);
nand UO_278 (O_278,N_22589,N_24825);
and UO_279 (O_279,N_23721,N_23478);
or UO_280 (O_280,N_22948,N_23242);
and UO_281 (O_281,N_23451,N_22123);
and UO_282 (O_282,N_23044,N_23434);
nor UO_283 (O_283,N_22487,N_23421);
or UO_284 (O_284,N_23358,N_23266);
or UO_285 (O_285,N_24642,N_22698);
or UO_286 (O_286,N_22410,N_24337);
xor UO_287 (O_287,N_23094,N_24163);
or UO_288 (O_288,N_23426,N_24639);
nand UO_289 (O_289,N_22513,N_24884);
nor UO_290 (O_290,N_22912,N_22408);
xor UO_291 (O_291,N_23749,N_22936);
or UO_292 (O_292,N_24238,N_23882);
xor UO_293 (O_293,N_22433,N_23148);
and UO_294 (O_294,N_24947,N_24831);
nor UO_295 (O_295,N_24237,N_23729);
nor UO_296 (O_296,N_24794,N_23786);
nand UO_297 (O_297,N_22420,N_24066);
xor UO_298 (O_298,N_23619,N_22465);
or UO_299 (O_299,N_24078,N_21950);
and UO_300 (O_300,N_22338,N_24667);
nand UO_301 (O_301,N_24620,N_22623);
xor UO_302 (O_302,N_21942,N_22148);
nand UO_303 (O_303,N_24637,N_22006);
or UO_304 (O_304,N_22187,N_22412);
and UO_305 (O_305,N_23686,N_22349);
and UO_306 (O_306,N_22867,N_23971);
xor UO_307 (O_307,N_22688,N_23712);
or UO_308 (O_308,N_22962,N_24095);
nand UO_309 (O_309,N_22326,N_23141);
nand UO_310 (O_310,N_22915,N_23133);
xnor UO_311 (O_311,N_22406,N_23617);
or UO_312 (O_312,N_22574,N_21991);
or UO_313 (O_313,N_24970,N_24969);
or UO_314 (O_314,N_21931,N_22225);
nand UO_315 (O_315,N_22021,N_23567);
nor UO_316 (O_316,N_23244,N_23058);
and UO_317 (O_317,N_23727,N_22768);
or UO_318 (O_318,N_24350,N_23162);
and UO_319 (O_319,N_23890,N_23866);
nand UO_320 (O_320,N_22679,N_22723);
or UO_321 (O_321,N_24729,N_23465);
or UO_322 (O_322,N_22043,N_23171);
nor UO_323 (O_323,N_24127,N_22400);
nand UO_324 (O_324,N_24379,N_24583);
nor UO_325 (O_325,N_23031,N_23933);
nand UO_326 (O_326,N_24232,N_23750);
nor UO_327 (O_327,N_22339,N_23127);
nor UO_328 (O_328,N_22963,N_22386);
or UO_329 (O_329,N_24929,N_23819);
or UO_330 (O_330,N_23533,N_23814);
and UO_331 (O_331,N_23039,N_22822);
nand UO_332 (O_332,N_24249,N_22908);
xor UO_333 (O_333,N_23409,N_23623);
nor UO_334 (O_334,N_24409,N_23359);
or UO_335 (O_335,N_22158,N_24986);
nand UO_336 (O_336,N_23512,N_22279);
nor UO_337 (O_337,N_24913,N_22325);
and UO_338 (O_338,N_24377,N_22005);
nor UO_339 (O_339,N_22959,N_23053);
xor UO_340 (O_340,N_24325,N_23947);
xor UO_341 (O_341,N_21883,N_22953);
xnor UO_342 (O_342,N_23560,N_23835);
and UO_343 (O_343,N_22787,N_21922);
nand UO_344 (O_344,N_23186,N_22473);
xnor UO_345 (O_345,N_23246,N_21881);
xnor UO_346 (O_346,N_22783,N_22937);
and UO_347 (O_347,N_24211,N_22931);
nand UO_348 (O_348,N_23158,N_22201);
nor UO_349 (O_349,N_22333,N_22305);
and UO_350 (O_350,N_22664,N_23847);
xnor UO_351 (O_351,N_24557,N_24944);
xor UO_352 (O_352,N_23238,N_24845);
and UO_353 (O_353,N_23201,N_22182);
nor UO_354 (O_354,N_21955,N_22556);
or UO_355 (O_355,N_23826,N_24865);
and UO_356 (O_356,N_24728,N_24334);
xor UO_357 (O_357,N_22130,N_24796);
nor UO_358 (O_358,N_22097,N_23714);
and UO_359 (O_359,N_24481,N_22792);
nand UO_360 (O_360,N_22779,N_22840);
and UO_361 (O_361,N_22619,N_24803);
nor UO_362 (O_362,N_24706,N_23733);
or UO_363 (O_363,N_23041,N_22418);
nor UO_364 (O_364,N_23395,N_24956);
xnor UO_365 (O_365,N_23643,N_23410);
xor UO_366 (O_366,N_22008,N_22208);
nand UO_367 (O_367,N_22671,N_24414);
xor UO_368 (O_368,N_22924,N_24508);
nor UO_369 (O_369,N_22837,N_22257);
and UO_370 (O_370,N_23120,N_23926);
nor UO_371 (O_371,N_23205,N_21968);
and UO_372 (O_372,N_22736,N_24544);
nand UO_373 (O_373,N_23809,N_23601);
or UO_374 (O_374,N_22713,N_21887);
nor UO_375 (O_375,N_22105,N_22220);
nor UO_376 (O_376,N_22251,N_21983);
and UO_377 (O_377,N_23799,N_24692);
nor UO_378 (O_378,N_24067,N_23709);
and UO_379 (O_379,N_22753,N_22950);
and UO_380 (O_380,N_23770,N_24720);
nor UO_381 (O_381,N_22666,N_23992);
nand UO_382 (O_382,N_24463,N_23401);
and UO_383 (O_383,N_24367,N_23159);
xnor UO_384 (O_384,N_23649,N_23674);
or UO_385 (O_385,N_22381,N_23959);
xor UO_386 (O_386,N_23989,N_21949);
or UO_387 (O_387,N_22719,N_22868);
nor UO_388 (O_388,N_23472,N_23378);
or UO_389 (O_389,N_22501,N_23063);
nor UO_390 (O_390,N_22724,N_23677);
xnor UO_391 (O_391,N_24461,N_22474);
nand UO_392 (O_392,N_23631,N_21996);
xor UO_393 (O_393,N_24558,N_24745);
xnor UO_394 (O_394,N_23744,N_22044);
xor UO_395 (O_395,N_24550,N_24063);
nand UO_396 (O_396,N_22287,N_22533);
nor UO_397 (O_397,N_24349,N_22147);
or UO_398 (O_398,N_22934,N_23412);
nand UO_399 (O_399,N_24586,N_22058);
or UO_400 (O_400,N_22765,N_23513);
nor UO_401 (O_401,N_23055,N_24433);
and UO_402 (O_402,N_24480,N_24636);
nor UO_403 (O_403,N_23871,N_22054);
or UO_404 (O_404,N_23497,N_23350);
xor UO_405 (O_405,N_23153,N_22335);
and UO_406 (O_406,N_24203,N_22570);
nor UO_407 (O_407,N_23281,N_24146);
nand UO_408 (O_408,N_23731,N_24626);
or UO_409 (O_409,N_24418,N_23224);
nand UO_410 (O_410,N_22884,N_22013);
nand UO_411 (O_411,N_24993,N_24596);
nor UO_412 (O_412,N_24003,N_23398);
or UO_413 (O_413,N_23433,N_23592);
nor UO_414 (O_414,N_24131,N_21905);
and UO_415 (O_415,N_24286,N_22856);
or UO_416 (O_416,N_24023,N_23249);
nand UO_417 (O_417,N_23262,N_24585);
nor UO_418 (O_418,N_23748,N_24933);
nor UO_419 (O_419,N_23593,N_22443);
nor UO_420 (O_420,N_24701,N_21963);
nand UO_421 (O_421,N_23324,N_22379);
and UO_422 (O_422,N_24885,N_23877);
and UO_423 (O_423,N_22176,N_23471);
and UO_424 (O_424,N_23261,N_22426);
nand UO_425 (O_425,N_23265,N_22876);
nor UO_426 (O_426,N_24967,N_22730);
and UO_427 (O_427,N_24500,N_23268);
xnor UO_428 (O_428,N_24028,N_22459);
and UO_429 (O_429,N_24864,N_24789);
nor UO_430 (O_430,N_24854,N_23511);
or UO_431 (O_431,N_24523,N_24058);
nor UO_432 (O_432,N_23504,N_24214);
and UO_433 (O_433,N_24814,N_22362);
and UO_434 (O_434,N_23216,N_22169);
or UO_435 (O_435,N_24496,N_23510);
xnor UO_436 (O_436,N_24510,N_22252);
or UO_437 (O_437,N_22390,N_23286);
and UO_438 (O_438,N_23563,N_24002);
or UO_439 (O_439,N_24380,N_24974);
xor UO_440 (O_440,N_24641,N_22447);
nand UO_441 (O_441,N_23297,N_22636);
nor UO_442 (O_442,N_24750,N_22760);
and UO_443 (O_443,N_24493,N_24454);
and UO_444 (O_444,N_22471,N_23954);
nor UO_445 (O_445,N_22717,N_23640);
or UO_446 (O_446,N_21934,N_23918);
nand UO_447 (O_447,N_22545,N_22088);
xor UO_448 (O_448,N_23344,N_22670);
xor UO_449 (O_449,N_23940,N_23708);
or UO_450 (O_450,N_23970,N_23458);
or UO_451 (O_451,N_23876,N_22301);
nand UO_452 (O_452,N_24330,N_22653);
or UO_453 (O_453,N_23627,N_23018);
and UO_454 (O_454,N_22499,N_22990);
nor UO_455 (O_455,N_24013,N_23553);
xnor UO_456 (O_456,N_23801,N_22467);
nor UO_457 (O_457,N_23194,N_23913);
and UO_458 (O_458,N_24823,N_24056);
nor UO_459 (O_459,N_23032,N_24727);
or UO_460 (O_460,N_21884,N_24401);
nand UO_461 (O_461,N_22638,N_24428);
nor UO_462 (O_462,N_23113,N_24370);
or UO_463 (O_463,N_23830,N_23934);
nand UO_464 (O_464,N_22367,N_22704);
or UO_465 (O_465,N_22068,N_24934);
nor UO_466 (O_466,N_24910,N_22193);
nor UO_467 (O_467,N_22481,N_23952);
nor UO_468 (O_468,N_22207,N_23726);
xor UO_469 (O_469,N_24469,N_23634);
xor UO_470 (O_470,N_22402,N_23596);
nor UO_471 (O_471,N_23377,N_23275);
and UO_472 (O_472,N_24164,N_23430);
nand UO_473 (O_473,N_24651,N_24902);
xnor UO_474 (O_474,N_22120,N_22171);
or UO_475 (O_475,N_24528,N_23195);
xor UO_476 (O_476,N_23208,N_22932);
nand UO_477 (O_477,N_23820,N_23705);
nor UO_478 (O_478,N_23237,N_23487);
xor UO_479 (O_479,N_23706,N_22370);
and UO_480 (O_480,N_22414,N_24898);
or UO_481 (O_481,N_22684,N_22213);
xnor UO_482 (O_482,N_22649,N_22231);
nor UO_483 (O_483,N_24772,N_23427);
or UO_484 (O_484,N_23424,N_23360);
nor UO_485 (O_485,N_23321,N_23298);
and UO_486 (O_486,N_24777,N_24175);
nand UO_487 (O_487,N_22373,N_22740);
and UO_488 (O_488,N_23873,N_24470);
and UO_489 (O_489,N_22630,N_24923);
xnor UO_490 (O_490,N_23061,N_23000);
nor UO_491 (O_491,N_23439,N_23920);
nor UO_492 (O_492,N_24545,N_24444);
and UO_493 (O_493,N_23267,N_24109);
and UO_494 (O_494,N_23568,N_24193);
or UO_495 (O_495,N_24129,N_24999);
or UO_496 (O_496,N_22848,N_23347);
nand UO_497 (O_497,N_22240,N_24773);
and UO_498 (O_498,N_21923,N_23684);
or UO_499 (O_499,N_23980,N_21896);
xor UO_500 (O_500,N_23301,N_24108);
or UO_501 (O_501,N_24327,N_24524);
and UO_502 (O_502,N_23921,N_22554);
and UO_503 (O_503,N_23074,N_23915);
xor UO_504 (O_504,N_24415,N_23707);
nand UO_505 (O_505,N_22857,N_22869);
nand UO_506 (O_506,N_24931,N_24570);
xnor UO_507 (O_507,N_22989,N_22864);
or UO_508 (O_508,N_22678,N_22037);
or UO_509 (O_509,N_23549,N_22797);
and UO_510 (O_510,N_23907,N_24811);
xor UO_511 (O_511,N_24683,N_23115);
nor UO_512 (O_512,N_23961,N_22003);
nand UO_513 (O_513,N_23278,N_23520);
or UO_514 (O_514,N_23695,N_23155);
nand UO_515 (O_515,N_23223,N_24069);
nor UO_516 (O_516,N_24270,N_22327);
nand UO_517 (O_517,N_22300,N_24424);
or UO_518 (O_518,N_23701,N_24546);
and UO_519 (O_519,N_22510,N_24080);
or UO_520 (O_520,N_22919,N_22781);
xnor UO_521 (O_521,N_22807,N_24488);
nor UO_522 (O_522,N_21982,N_24413);
xnor UO_523 (O_523,N_23247,N_23316);
nor UO_524 (O_524,N_24394,N_24335);
and UO_525 (O_525,N_21927,N_24497);
nor UO_526 (O_526,N_23575,N_22255);
nand UO_527 (O_527,N_23927,N_22155);
nand UO_528 (O_528,N_23161,N_21909);
xor UO_529 (O_529,N_24659,N_23489);
xor UO_530 (O_530,N_24427,N_24277);
or UO_531 (O_531,N_24347,N_22865);
and UO_532 (O_532,N_23405,N_22893);
xnor UO_533 (O_533,N_23295,N_23309);
nand UO_534 (O_534,N_23722,N_24705);
nor UO_535 (O_535,N_23765,N_24133);
and UO_536 (O_536,N_22161,N_22838);
xnor UO_537 (O_537,N_24144,N_24519);
xor UO_538 (O_538,N_24632,N_22812);
and UO_539 (O_539,N_22820,N_24768);
nor UO_540 (O_540,N_22821,N_22451);
and UO_541 (O_541,N_24271,N_24526);
xor UO_542 (O_542,N_23974,N_22180);
and UO_543 (O_543,N_24051,N_24590);
nor UO_544 (O_544,N_22316,N_22129);
nor UO_545 (O_545,N_23929,N_22014);
or UO_546 (O_546,N_24603,N_23184);
and UO_547 (O_547,N_23767,N_22237);
and UO_548 (O_548,N_24459,N_24060);
and UO_549 (O_549,N_22230,N_24495);
and UO_550 (O_550,N_24406,N_23523);
nor UO_551 (O_551,N_22020,N_24767);
nor UO_552 (O_552,N_24536,N_24911);
nor UO_553 (O_553,N_22707,N_24083);
nand UO_554 (O_554,N_22744,N_24593);
nand UO_555 (O_555,N_24156,N_24691);
nor UO_556 (O_556,N_22108,N_24711);
and UO_557 (O_557,N_24505,N_23292);
nor UO_558 (O_558,N_24245,N_24140);
nor UO_559 (O_559,N_23131,N_24625);
nor UO_560 (O_560,N_22002,N_22553);
nor UO_561 (O_561,N_22153,N_22642);
nor UO_562 (O_562,N_23632,N_23768);
and UO_563 (O_563,N_24411,N_23334);
nand UO_564 (O_564,N_23033,N_22700);
nor UO_565 (O_565,N_24757,N_22943);
or UO_566 (O_566,N_23717,N_24666);
xor UO_567 (O_567,N_24007,N_24043);
and UO_568 (O_568,N_24684,N_23755);
or UO_569 (O_569,N_23604,N_21890);
and UO_570 (O_570,N_22917,N_21941);
and UO_571 (O_571,N_24103,N_23012);
nor UO_572 (O_572,N_22565,N_21913);
xor UO_573 (O_573,N_24714,N_22617);
and UO_574 (O_574,N_24552,N_24455);
nor UO_575 (O_575,N_23446,N_22074);
or UO_576 (O_576,N_22754,N_24674);
nand UO_577 (O_577,N_23599,N_22450);
nor UO_578 (O_578,N_22055,N_23466);
nor UO_579 (O_579,N_22764,N_23916);
xor UO_580 (O_580,N_24722,N_23282);
and UO_581 (O_581,N_24240,N_23290);
nand UO_582 (O_582,N_24653,N_23546);
and UO_583 (O_583,N_23610,N_23176);
and UO_584 (O_584,N_22346,N_24258);
xnor UO_585 (O_585,N_23024,N_24273);
and UO_586 (O_586,N_22566,N_24785);
xor UO_587 (O_587,N_24391,N_22520);
nor UO_588 (O_588,N_24837,N_23132);
xor UO_589 (O_589,N_22355,N_22281);
xnor UO_590 (O_590,N_23864,N_23025);
or UO_591 (O_591,N_23363,N_22045);
nand UO_592 (O_592,N_23390,N_24181);
nand UO_593 (O_593,N_23342,N_22456);
or UO_594 (O_594,N_21999,N_22033);
or UO_595 (O_595,N_23664,N_23620);
xnor UO_596 (O_596,N_22863,N_24450);
nor UO_597 (O_597,N_22053,N_24747);
or UO_598 (O_598,N_23169,N_22877);
nand UO_599 (O_599,N_23783,N_22656);
or UO_600 (O_600,N_22799,N_22154);
xnor UO_601 (O_601,N_24014,N_23887);
and UO_602 (O_602,N_23635,N_23597);
nor UO_603 (O_603,N_22063,N_23151);
nor UO_604 (O_604,N_21972,N_24160);
xor UO_605 (O_605,N_22515,N_24036);
xor UO_606 (O_606,N_24940,N_24436);
xnor UO_607 (O_607,N_24030,N_24344);
nand UO_608 (O_608,N_22392,N_22938);
nor UO_609 (O_609,N_23659,N_23595);
or UO_610 (O_610,N_22910,N_22745);
nor UO_611 (O_611,N_23589,N_23855);
nor UO_612 (O_612,N_23166,N_23449);
and UO_613 (O_613,N_23240,N_24019);
and UO_614 (O_614,N_24204,N_22541);
xnor UO_615 (O_615,N_23841,N_23953);
or UO_616 (O_616,N_22218,N_24792);
nand UO_617 (O_617,N_24012,N_22905);
nand UO_618 (O_618,N_22732,N_24487);
and UO_619 (O_619,N_23419,N_24267);
xnor UO_620 (O_620,N_23518,N_21984);
or UO_621 (O_621,N_22331,N_24588);
or UO_622 (O_622,N_22315,N_24627);
nor UO_623 (O_623,N_24709,N_24813);
or UO_624 (O_624,N_23527,N_23771);
nand UO_625 (O_625,N_22805,N_22752);
and UO_626 (O_626,N_22317,N_24584);
xnor UO_627 (O_627,N_24856,N_24143);
xor UO_628 (O_628,N_22297,N_24749);
nor UO_629 (O_629,N_23450,N_24319);
xnor UO_630 (O_630,N_22151,N_24294);
and UO_631 (O_631,N_22798,N_24098);
nand UO_632 (O_632,N_24735,N_22181);
xor UO_633 (O_633,N_24756,N_23073);
or UO_634 (O_634,N_22596,N_24815);
nor UO_635 (O_635,N_24052,N_23530);
and UO_636 (O_636,N_22039,N_22397);
and UO_637 (O_637,N_22241,N_24035);
and UO_638 (O_638,N_24827,N_24533);
and UO_639 (O_639,N_22387,N_24942);
nand UO_640 (O_640,N_22690,N_24894);
nand UO_641 (O_641,N_22374,N_22247);
or UO_642 (O_642,N_23857,N_22939);
nor UO_643 (O_643,N_23177,N_24431);
and UO_644 (O_644,N_22341,N_22751);
nor UO_645 (O_645,N_22665,N_24621);
and UO_646 (O_646,N_24006,N_23392);
xor UO_647 (O_647,N_23234,N_23432);
and UO_648 (O_648,N_22766,N_24725);
nor UO_649 (O_649,N_23805,N_23447);
and UO_650 (O_650,N_22576,N_23227);
and UO_651 (O_651,N_22861,N_22095);
and UO_652 (O_652,N_24645,N_22883);
nor UO_653 (O_653,N_22289,N_23548);
nor UO_654 (O_654,N_23833,N_24135);
nor UO_655 (O_655,N_22898,N_22895);
xnor UO_656 (O_656,N_24265,N_22444);
nor UO_657 (O_657,N_22493,N_22721);
or UO_658 (O_658,N_23323,N_22878);
or UO_659 (O_659,N_24959,N_22081);
and UO_660 (O_660,N_24483,N_22925);
nand UO_661 (O_661,N_23957,N_24724);
nor UO_662 (O_662,N_23834,N_24514);
nand UO_663 (O_663,N_22076,N_23474);
and UO_664 (O_664,N_22996,N_23912);
and UO_665 (O_665,N_22363,N_23577);
or UO_666 (O_666,N_24623,N_22720);
nand UO_667 (O_667,N_24378,N_23029);
nor UO_668 (O_668,N_24285,N_24176);
and UO_669 (O_669,N_22762,N_24950);
nor UO_670 (O_670,N_24841,N_22334);
nor UO_671 (O_671,N_23822,N_24598);
xnor UO_672 (O_672,N_23322,N_23067);
and UO_673 (O_673,N_22253,N_22605);
nand UO_674 (O_674,N_23668,N_24595);
nand UO_675 (O_675,N_23116,N_23335);
and UO_676 (O_676,N_22609,N_22888);
nor UO_677 (O_677,N_24972,N_23657);
nand UO_678 (O_678,N_24489,N_22731);
xnor UO_679 (O_679,N_23004,N_22209);
nand UO_680 (O_680,N_22141,N_22667);
nand UO_681 (O_681,N_23856,N_23534);
xnor UO_682 (O_682,N_24020,N_23507);
nor UO_683 (O_683,N_21880,N_22742);
nand UO_684 (O_684,N_24805,N_24348);
or UO_685 (O_685,N_23608,N_22960);
nand UO_686 (O_686,N_23485,N_24416);
xor UO_687 (O_687,N_22945,N_23429);
nand UO_688 (O_688,N_23319,N_24071);
nand UO_689 (O_689,N_23035,N_23995);
nor UO_690 (O_690,N_22608,N_24106);
xor UO_691 (O_691,N_22911,N_23694);
nor UO_692 (O_692,N_22041,N_24445);
xnor UO_693 (O_693,N_24739,N_22850);
and UO_694 (O_694,N_23337,N_21919);
or UO_695 (O_695,N_24092,N_22635);
or UO_696 (O_696,N_22793,N_23103);
or UO_697 (O_697,N_23796,N_24601);
nor UO_698 (O_698,N_21959,N_24988);
nand UO_699 (O_699,N_22514,N_22405);
and UO_700 (O_700,N_23385,N_24081);
and UO_701 (O_701,N_22542,N_24656);
and UO_702 (O_702,N_24186,N_22149);
or UO_703 (O_703,N_24703,N_22951);
xor UO_704 (O_704,N_24466,N_24113);
nand UO_705 (O_705,N_23117,N_22527);
and UO_706 (O_706,N_23785,N_24121);
xor UO_707 (O_707,N_22946,N_22204);
and UO_708 (O_708,N_24943,N_23327);
xnor UO_709 (O_709,N_22396,N_24438);
nand UO_710 (O_710,N_22051,N_22836);
and UO_711 (O_711,N_22658,N_24892);
nor UO_712 (O_712,N_24927,N_22529);
xnor UO_713 (O_713,N_24115,N_22394);
or UO_714 (O_714,N_23715,N_23779);
nand UO_715 (O_715,N_24861,N_23248);
or UO_716 (O_716,N_24802,N_24952);
and UO_717 (O_717,N_24197,N_23603);
nor UO_718 (O_718,N_22425,N_24622);
nand UO_719 (O_719,N_24358,N_24061);
and UO_720 (O_720,N_24266,N_22739);
nand UO_721 (O_721,N_23138,N_22735);
nor UO_722 (O_722,N_22319,N_24780);
nand UO_723 (O_723,N_24503,N_23006);
nand UO_724 (O_724,N_22718,N_23792);
and UO_725 (O_725,N_23199,N_24990);
and UO_726 (O_726,N_23666,N_23017);
xor UO_727 (O_727,N_24743,N_23624);
and UO_728 (O_728,N_24843,N_21978);
and UO_729 (O_729,N_24618,N_22162);
and UO_730 (O_730,N_24356,N_24696);
xnor UO_731 (O_731,N_24681,N_24376);
or UO_732 (O_732,N_24769,N_24888);
and UO_733 (O_733,N_24096,N_24075);
xnor UO_734 (O_734,N_23536,N_22621);
nor UO_735 (O_735,N_23683,N_24166);
xor UO_736 (O_736,N_24236,N_22886);
nand UO_737 (O_737,N_23457,N_24937);
or UO_738 (O_738,N_22974,N_24298);
or UO_739 (O_739,N_24230,N_22685);
or UO_740 (O_740,N_22916,N_22663);
nand UO_741 (O_741,N_22085,N_22337);
and UO_742 (O_742,N_22083,N_22845);
and UO_743 (O_743,N_24038,N_24840);
nand UO_744 (O_744,N_24257,N_23425);
nand UO_745 (O_745,N_22269,N_22029);
nor UO_746 (O_746,N_24690,N_24594);
nand UO_747 (O_747,N_23576,N_23013);
nand UO_748 (O_748,N_24511,N_24755);
or UO_749 (O_749,N_22562,N_21895);
xor UO_750 (O_750,N_23050,N_23364);
nand UO_751 (O_751,N_24219,N_24198);
nand UO_752 (O_752,N_23555,N_22266);
and UO_753 (O_753,N_24572,N_22777);
nand UO_754 (O_754,N_23299,N_23781);
and UO_755 (O_755,N_24912,N_21939);
nor UO_756 (O_756,N_24672,N_24024);
nand UO_757 (O_757,N_22817,N_24867);
and UO_758 (O_758,N_22243,N_24915);
nand UO_759 (O_759,N_24093,N_23886);
nor UO_760 (O_760,N_24985,N_22399);
xnor UO_761 (O_761,N_23414,N_22087);
or UO_762 (O_762,N_23403,N_24786);
xor UO_763 (O_763,N_22078,N_23212);
nor UO_764 (O_764,N_24216,N_22361);
nor UO_765 (O_765,N_22539,N_23101);
or UO_766 (O_766,N_22271,N_24563);
nand UO_767 (O_767,N_23896,N_24116);
and UO_768 (O_768,N_23700,N_24323);
nand UO_769 (O_769,N_22602,N_24788);
or UO_770 (O_770,N_24775,N_24456);
nand UO_771 (O_771,N_24685,N_22323);
nor UO_772 (O_772,N_22597,N_24571);
nor UO_773 (O_773,N_24033,N_24305);
or UO_774 (O_774,N_22174,N_23526);
nand UO_775 (O_775,N_22328,N_23633);
or UO_776 (O_776,N_22214,N_23506);
or UO_777 (O_777,N_23730,N_22498);
or UO_778 (O_778,N_24643,N_23167);
nand UO_779 (O_779,N_24362,N_22371);
or UO_780 (O_780,N_24660,N_24909);
nor UO_781 (O_781,N_23438,N_22177);
or UO_782 (O_782,N_22702,N_22887);
xor UO_783 (O_783,N_23808,N_24791);
xnor UO_784 (O_784,N_22988,N_23494);
nand UO_785 (O_785,N_24869,N_22543);
nand UO_786 (O_786,N_23109,N_24547);
xor UO_787 (O_787,N_22522,N_22118);
xor UO_788 (O_788,N_22235,N_24086);
and UO_789 (O_789,N_24425,N_23291);
xnor UO_790 (O_790,N_24479,N_22203);
or UO_791 (O_791,N_22296,N_22458);
xnor UO_792 (O_792,N_24941,N_21910);
xnor UO_793 (O_793,N_22802,N_23571);
nand UO_794 (O_794,N_24303,N_24619);
xor UO_795 (O_795,N_24199,N_22906);
nor UO_796 (O_796,N_24321,N_23198);
or UO_797 (O_797,N_23501,N_22672);
or UO_798 (O_798,N_23754,N_22254);
or UO_799 (O_799,N_23906,N_24515);
nor UO_800 (O_800,N_24010,N_23349);
nand UO_801 (O_801,N_24573,N_24090);
nand UO_802 (O_802,N_23196,N_21954);
xnor UO_803 (O_803,N_22278,N_22629);
or UO_804 (O_804,N_24975,N_21943);
nand UO_805 (O_805,N_22001,N_23988);
or UO_806 (O_806,N_23387,N_24040);
or UO_807 (O_807,N_24873,N_23525);
nand UO_808 (O_808,N_23402,N_22559);
or UO_809 (O_809,N_24393,N_21966);
nand UO_810 (O_810,N_22615,N_24301);
nand UO_811 (O_811,N_23747,N_24730);
or UO_812 (O_812,N_24539,N_21889);
nor UO_813 (O_813,N_22918,N_23607);
and UO_814 (O_814,N_23735,N_22066);
xnor UO_815 (O_815,N_23849,N_22894);
xor UO_816 (O_816,N_24693,N_23579);
or UO_817 (O_817,N_24082,N_22511);
nand UO_818 (O_818,N_22590,N_23122);
or UO_819 (O_819,N_22288,N_23296);
nor UO_820 (O_820,N_23100,N_23945);
nor UO_821 (O_821,N_24150,N_22115);
or UO_822 (O_822,N_22506,N_24716);
nand UO_823 (O_823,N_22476,N_23144);
nor UO_824 (O_824,N_22496,N_22302);
nand UO_825 (O_825,N_24485,N_23040);
xnor UO_826 (O_826,N_23099,N_24256);
and UO_827 (O_827,N_22852,N_24992);
or UO_828 (O_828,N_24649,N_21885);
nand UO_829 (O_829,N_22036,N_22368);
nand UO_830 (O_830,N_24312,N_24222);
xnor UO_831 (O_831,N_22920,N_23736);
nand UO_832 (O_832,N_23241,N_24467);
nand UO_833 (O_833,N_23566,N_22659);
nor UO_834 (O_834,N_24084,N_22011);
or UO_835 (O_835,N_23993,N_23688);
or UO_836 (O_836,N_23181,N_22272);
xnor UO_837 (O_837,N_24964,N_22645);
xor UO_838 (O_838,N_22759,N_22185);
nor UO_839 (O_839,N_24799,N_22265);
or UO_840 (O_840,N_23328,N_24784);
or UO_841 (O_841,N_23897,N_23862);
or UO_842 (O_842,N_24435,N_23271);
or UO_843 (O_843,N_21986,N_23160);
nor UO_844 (O_844,N_22150,N_24125);
xnor UO_845 (O_845,N_22343,N_24338);
nor UO_846 (O_846,N_22062,N_23652);
or UO_847 (O_847,N_24556,N_22881);
or UO_848 (O_848,N_24926,N_24553);
xor UO_849 (O_849,N_22294,N_22308);
nand UO_850 (O_850,N_22624,N_24462);
nand UO_851 (O_851,N_24253,N_22976);
nor UO_852 (O_852,N_24804,N_22157);
nor UO_853 (O_853,N_22275,N_24022);
nand UO_854 (O_854,N_22216,N_23812);
nand UO_855 (O_855,N_24192,N_22725);
or UO_856 (O_856,N_22750,N_22113);
or UO_857 (O_857,N_24663,N_23817);
nand UO_858 (O_858,N_24440,N_24697);
xor UO_859 (O_859,N_22061,N_23543);
nand UO_860 (O_860,N_24689,N_24059);
and UO_861 (O_861,N_22784,N_22604);
and UO_862 (O_862,N_22892,N_23725);
xnor UO_863 (O_863,N_22096,N_21973);
or UO_864 (O_864,N_24770,N_22484);
and UO_865 (O_865,N_22248,N_24908);
nor UO_866 (O_866,N_22344,N_21914);
or UO_867 (O_867,N_24345,N_21912);
xor UO_868 (O_868,N_24016,N_22680);
and UO_869 (O_869,N_24293,N_23370);
or UO_870 (O_870,N_23312,N_22708);
nand UO_871 (O_871,N_22794,N_22738);
and UO_872 (O_872,N_24446,N_24371);
or UO_873 (O_873,N_24901,N_22378);
or UO_874 (O_874,N_22873,N_22310);
xnor UO_875 (O_875,N_23861,N_23353);
and UO_876 (O_876,N_24354,N_23661);
or UO_877 (O_877,N_24408,N_22699);
xor UO_878 (O_878,N_24123,N_24662);
nand UO_879 (O_879,N_23376,N_22380);
nand UO_880 (O_880,N_22084,N_24903);
xnor UO_881 (O_881,N_23815,N_22075);
or UO_882 (O_882,N_22844,N_24254);
nand UO_883 (O_883,N_23210,N_23023);
xor UO_884 (O_884,N_22126,N_22398);
nand UO_885 (O_885,N_24630,N_22422);
nor UO_886 (O_886,N_24372,N_23648);
xor UO_887 (O_887,N_23538,N_24458);
or UO_888 (O_888,N_23052,N_24578);
nor UO_889 (O_889,N_22652,N_23946);
nand UO_890 (O_890,N_23367,N_24790);
and UO_891 (O_891,N_22073,N_23180);
or UO_892 (O_892,N_23235,N_23955);
or UO_893 (O_893,N_23773,N_24202);
xor UO_894 (O_894,N_24011,N_24939);
and UO_895 (O_895,N_24616,N_24464);
nand UO_896 (O_896,N_24833,N_24916);
nand UO_897 (O_897,N_23691,N_23728);
and UO_898 (O_898,N_24906,N_24717);
and UO_899 (O_899,N_22926,N_22353);
xnor UO_900 (O_900,N_22067,N_22987);
xor UO_901 (O_901,N_23791,N_22668);
nand UO_902 (O_902,N_23411,N_22274);
xor UO_903 (O_903,N_22489,N_23225);
or UO_904 (O_904,N_23274,N_24742);
or UO_905 (O_905,N_23910,N_24982);
nand UO_906 (O_906,N_22479,N_24948);
nor UO_907 (O_907,N_24597,N_22591);
nor UO_908 (O_908,N_24169,N_23066);
xor UO_909 (O_909,N_23853,N_23752);
or UO_910 (O_910,N_23098,N_23326);
xnor UO_911 (O_911,N_24386,N_21998);
xor UO_912 (O_912,N_23178,N_22221);
nand UO_913 (O_913,N_21888,N_22572);
nand UO_914 (O_914,N_22226,N_23043);
or UO_915 (O_915,N_22273,N_24357);
and UO_916 (O_916,N_21936,N_24538);
nand UO_917 (O_917,N_21932,N_21907);
or UO_918 (O_918,N_22632,N_21946);
nor UO_919 (O_919,N_24576,N_22048);
nand UO_920 (O_920,N_24921,N_23584);
nand UO_921 (O_921,N_24676,N_23382);
or UO_922 (O_922,N_23724,N_22089);
and UO_923 (O_923,N_22461,N_24712);
nand UO_924 (O_924,N_22313,N_22421);
nor UO_925 (O_925,N_22102,N_22436);
nor UO_926 (O_926,N_24173,N_24064);
nor UO_927 (O_927,N_22486,N_23134);
or UO_928 (O_928,N_21997,N_23087);
and UO_929 (O_929,N_22092,N_23776);
nand UO_930 (O_930,N_24279,N_23991);
and UO_931 (O_931,N_24820,N_22179);
nor UO_932 (O_932,N_23996,N_24648);
xor UO_933 (O_933,N_24879,N_24951);
nand UO_934 (O_934,N_22715,N_22860);
nor UO_935 (O_935,N_23111,N_22059);
and UO_936 (O_936,N_22464,N_24871);
or UO_937 (O_937,N_22469,N_22428);
nor UO_938 (O_938,N_23371,N_21892);
nand UO_939 (O_939,N_22761,N_22567);
or UO_940 (O_940,N_23479,N_24548);
xor UO_941 (O_941,N_22299,N_23690);
nor UO_942 (O_942,N_23002,N_22224);
xnor UO_943 (O_943,N_21916,N_24498);
or UO_944 (O_944,N_23260,N_24532);
nor UO_945 (O_945,N_24816,N_24094);
nor UO_946 (O_946,N_24322,N_24110);
xnor UO_947 (O_947,N_22128,N_23774);
nor UO_948 (O_948,N_23756,N_24581);
and UO_949 (O_949,N_23669,N_24617);
and UO_950 (O_950,N_24737,N_23997);
xor UO_951 (O_951,N_24374,N_23190);
nand UO_952 (O_952,N_22452,N_22874);
nor UO_953 (O_953,N_23734,N_23761);
or UO_954 (O_954,N_22336,N_23977);
nor UO_955 (O_955,N_23202,N_23393);
or UO_956 (O_956,N_22524,N_23539);
and UO_957 (O_957,N_24046,N_23175);
or UO_958 (O_958,N_23831,N_23505);
and UO_959 (O_959,N_22199,N_23136);
nand UO_960 (O_960,N_21937,N_22352);
or UO_961 (O_961,N_21958,N_23016);
or UO_962 (O_962,N_24778,N_23444);
xnor UO_963 (O_963,N_24453,N_22119);
and UO_964 (O_964,N_24611,N_23215);
nor UO_965 (O_965,N_23204,N_23351);
nand UO_966 (O_966,N_22427,N_24241);
and UO_967 (O_967,N_23081,N_24471);
xor UO_968 (O_968,N_23254,N_24938);
nand UO_969 (O_969,N_24658,N_22017);
or UO_970 (O_970,N_24628,N_23203);
or UO_971 (O_971,N_23626,N_24899);
or UO_972 (O_972,N_24053,N_24073);
nor UO_973 (O_973,N_23854,N_22756);
xnor UO_974 (O_974,N_23284,N_24045);
xor UO_975 (O_975,N_24205,N_24218);
nand UO_976 (O_976,N_22104,N_24602);
or UO_977 (O_977,N_23994,N_22079);
and UO_978 (O_978,N_24860,N_24120);
xor UO_979 (O_979,N_23142,N_22485);
nor UO_980 (O_980,N_22618,N_24932);
nor UO_981 (O_981,N_22369,N_22242);
or UO_982 (O_982,N_22028,N_22250);
nor UO_983 (O_983,N_24541,N_23885);
nand UO_984 (O_984,N_23384,N_22424);
or UO_985 (O_985,N_22914,N_24634);
xnor UO_986 (O_986,N_23088,N_24996);
nand UO_987 (O_987,N_24591,N_22737);
xnor UO_988 (O_988,N_24187,N_24260);
xnor UO_989 (O_989,N_23638,N_24300);
or UO_990 (O_990,N_21994,N_23935);
and UO_991 (O_991,N_22696,N_24283);
nor UO_992 (O_992,N_22110,N_22347);
and UO_993 (O_993,N_23036,N_22016);
or UO_994 (O_994,N_22525,N_24812);
xor UO_995 (O_995,N_24977,N_24779);
or UO_996 (O_996,N_23651,N_23172);
nand UO_997 (O_997,N_24842,N_24925);
or UO_998 (O_998,N_24246,N_22947);
xor UO_999 (O_999,N_24607,N_22223);
and UO_1000 (O_1000,N_24555,N_23096);
nand UO_1001 (O_1001,N_23365,N_24206);
or UO_1002 (O_1002,N_22622,N_23598);
xor UO_1003 (O_1003,N_24299,N_22978);
xnor UO_1004 (O_1004,N_24644,N_22245);
or UO_1005 (O_1005,N_22165,N_24665);
xnor UO_1006 (O_1006,N_22849,N_24295);
nor UO_1007 (O_1007,N_24704,N_24810);
nor UO_1008 (O_1008,N_22823,N_23636);
nand UO_1009 (O_1009,N_22277,N_22595);
and UO_1010 (O_1010,N_22263,N_23650);
xor UO_1011 (O_1011,N_22695,N_22901);
nand UO_1012 (O_1012,N_23211,N_24264);
and UO_1013 (O_1013,N_23336,N_23496);
xnor UO_1014 (O_1014,N_24965,N_23628);
nand UO_1015 (O_1015,N_22239,N_22259);
xor UO_1016 (O_1016,N_24849,N_22376);
nor UO_1017 (O_1017,N_22795,N_23079);
nor UO_1018 (O_1018,N_24465,N_24800);
xor UO_1019 (O_1019,N_22748,N_24981);
nor UO_1020 (O_1020,N_21985,N_23014);
and UO_1021 (O_1021,N_23368,N_22921);
nand UO_1022 (O_1022,N_23437,N_22413);
nand UO_1023 (O_1023,N_22880,N_22516);
or UO_1024 (O_1024,N_24227,N_22640);
or UO_1025 (O_1025,N_24317,N_22982);
nand UO_1026 (O_1026,N_24486,N_22669);
and UO_1027 (O_1027,N_22528,N_23616);
and UO_1028 (O_1028,N_22625,N_22012);
nand UO_1029 (O_1029,N_23086,N_21904);
or UO_1030 (O_1030,N_24278,N_22183);
nand UO_1031 (O_1031,N_23751,N_22189);
nor UO_1032 (O_1032,N_23108,N_21929);
xor UO_1033 (O_1033,N_22561,N_22891);
and UO_1034 (O_1034,N_23969,N_21962);
and UO_1035 (O_1035,N_24478,N_23972);
xnor UO_1036 (O_1036,N_23397,N_24978);
and UO_1037 (O_1037,N_22796,N_22488);
or UO_1038 (O_1038,N_23795,N_21930);
and UO_1039 (O_1039,N_23905,N_22019);
xor UO_1040 (O_1040,N_23803,N_23026);
xor UO_1041 (O_1041,N_24893,N_23775);
xnor UO_1042 (O_1042,N_23482,N_22689);
or UO_1043 (O_1043,N_23532,N_23277);
nand UO_1044 (O_1044,N_24961,N_24366);
xor UO_1045 (O_1045,N_24177,N_23629);
nand UO_1046 (O_1046,N_24005,N_23076);
and UO_1047 (O_1047,N_23308,N_23879);
and UO_1048 (O_1048,N_23612,N_21935);
or UO_1049 (O_1049,N_23229,N_22280);
or UO_1050 (O_1050,N_23860,N_23990);
nor UO_1051 (O_1051,N_23590,N_22205);
nand UO_1052 (O_1052,N_22332,N_22131);
and UO_1053 (O_1053,N_23200,N_24333);
nor UO_1054 (O_1054,N_22767,N_23580);
or UO_1055 (O_1055,N_22819,N_22651);
or UO_1056 (O_1056,N_22492,N_22403);
nor UO_1057 (O_1057,N_23984,N_22583);
nand UO_1058 (O_1058,N_23135,N_22311);
xnor UO_1059 (O_1059,N_24957,N_22858);
and UO_1060 (O_1060,N_24207,N_23739);
xnor UO_1061 (O_1061,N_23662,N_22423);
nand UO_1062 (O_1062,N_23509,N_21947);
and UO_1063 (O_1063,N_23838,N_24054);
and UO_1064 (O_1064,N_23793,N_23845);
xor UO_1065 (O_1065,N_21964,N_23173);
and UO_1066 (O_1066,N_23914,N_24326);
and UO_1067 (O_1067,N_24384,N_23760);
and UO_1068 (O_1068,N_23019,N_22435);
xnor UO_1069 (O_1069,N_22448,N_23844);
nand UO_1070 (O_1070,N_22470,N_24284);
and UO_1071 (O_1071,N_23009,N_24209);
and UO_1072 (O_1072,N_24074,N_22478);
xnor UO_1073 (O_1073,N_24525,N_23383);
nor UO_1074 (O_1074,N_22909,N_23021);
xor UO_1075 (O_1075,N_22046,N_24953);
nor UO_1076 (O_1076,N_24491,N_22958);
nor UO_1077 (O_1077,N_23852,N_23925);
nor UO_1078 (O_1078,N_23591,N_24223);
or UO_1079 (O_1079,N_24157,N_24846);
nand UO_1080 (O_1080,N_24194,N_23840);
or UO_1081 (O_1081,N_24868,N_24161);
nand UO_1082 (O_1082,N_22534,N_22351);
and UO_1083 (O_1083,N_21899,N_22746);
nand UO_1084 (O_1084,N_24710,N_24582);
xor UO_1085 (O_1085,N_24613,N_24026);
or UO_1086 (O_1086,N_22571,N_23338);
or UO_1087 (O_1087,N_23719,N_24141);
nand UO_1088 (O_1088,N_24473,N_23110);
or UO_1089 (O_1089,N_23288,N_24447);
and UO_1090 (O_1090,N_24781,N_23529);
xor UO_1091 (O_1091,N_24484,N_22445);
or UO_1092 (O_1092,N_22304,N_22070);
xor UO_1093 (O_1093,N_24829,N_22446);
xnor UO_1094 (O_1094,N_24397,N_23558);
nor UO_1095 (O_1095,N_23689,N_24147);
nor UO_1096 (O_1096,N_23542,N_23452);
nand UO_1097 (O_1097,N_24448,N_24373);
nor UO_1098 (O_1098,N_22438,N_24171);
xor UO_1099 (O_1099,N_22359,N_23975);
xnor UO_1100 (O_1100,N_23508,N_24304);
nand UO_1101 (O_1101,N_23352,N_23692);
nor UO_1102 (O_1102,N_24385,N_23071);
and UO_1103 (O_1103,N_23698,N_22117);
nand UO_1104 (O_1104,N_22188,N_22258);
or UO_1105 (O_1105,N_22497,N_24551);
nor UO_1106 (O_1106,N_22809,N_22674);
nor UO_1107 (O_1107,N_24234,N_24702);
xor UO_1108 (O_1108,N_22345,N_22957);
or UO_1109 (O_1109,N_23149,N_24468);
nand UO_1110 (O_1110,N_23020,N_23307);
and UO_1111 (O_1111,N_24184,N_24874);
and UO_1112 (O_1112,N_24715,N_24070);
nand UO_1113 (O_1113,N_23743,N_22611);
nand UO_1114 (O_1114,N_22806,N_24989);
nand UO_1115 (O_1115,N_24518,N_22600);
nand UO_1116 (O_1116,N_22509,N_22701);
or UO_1117 (O_1117,N_22601,N_23107);
nor UO_1118 (O_1118,N_23656,N_23475);
or UO_1119 (O_1119,N_22992,N_22307);
nor UO_1120 (O_1120,N_22641,N_23317);
nor UO_1121 (O_1121,N_22164,N_21945);
nand UO_1122 (O_1122,N_24008,N_24001);
xnor UO_1123 (O_1123,N_22285,N_22144);
nand UO_1124 (O_1124,N_24152,N_24225);
nand UO_1125 (O_1125,N_22907,N_22090);
xnor UO_1126 (O_1126,N_23524,N_24564);
or UO_1127 (O_1127,N_24762,N_24288);
or UO_1128 (O_1128,N_21975,N_23233);
and UO_1129 (O_1129,N_23152,N_24275);
nand UO_1130 (O_1130,N_23333,N_24698);
or UO_1131 (O_1131,N_24887,N_24158);
nor UO_1132 (O_1132,N_23909,N_23346);
or UO_1133 (O_1133,N_22194,N_22026);
and UO_1134 (O_1134,N_22788,N_22833);
or UO_1135 (O_1135,N_24311,N_23930);
nor UO_1136 (O_1136,N_23703,N_23667);
xor UO_1137 (O_1137,N_24365,N_23948);
and UO_1138 (O_1138,N_22586,N_24806);
nor UO_1139 (O_1139,N_24542,N_24297);
xor UO_1140 (O_1140,N_23226,N_21993);
nor UO_1141 (O_1141,N_23276,N_22801);
and UO_1142 (O_1142,N_23056,N_24566);
nor UO_1143 (O_1143,N_23547,N_24881);
nor UO_1144 (O_1144,N_24400,N_23010);
nand UO_1145 (O_1145,N_23263,N_24599);
nor UO_1146 (O_1146,N_24828,N_22814);
and UO_1147 (O_1147,N_22847,N_22356);
nand UO_1148 (O_1148,N_23217,N_22537);
xnor UO_1149 (O_1149,N_23973,N_23473);
or UO_1150 (O_1150,N_23250,N_23102);
xnor UO_1151 (O_1151,N_24139,N_24896);
nand UO_1152 (O_1152,N_23045,N_23034);
xor UO_1153 (O_1153,N_24801,N_22042);
and UO_1154 (O_1154,N_22437,N_22581);
nand UO_1155 (O_1155,N_24029,N_24771);
nor UO_1156 (O_1156,N_24114,N_22526);
xnor UO_1157 (O_1157,N_23391,N_22099);
and UO_1158 (O_1158,N_22004,N_24633);
nor UO_1159 (O_1159,N_22904,N_22000);
xnor UO_1160 (O_1160,N_22703,N_22264);
or UO_1161 (O_1161,N_22675,N_23372);
nand UO_1162 (O_1162,N_22329,N_23942);
nand UO_1163 (O_1163,N_22791,N_23315);
xnor UO_1164 (O_1164,N_23865,N_23077);
and UO_1165 (O_1165,N_21918,N_23121);
and UO_1166 (O_1166,N_23828,N_22999);
xor UO_1167 (O_1167,N_23746,N_24850);
nor UO_1168 (O_1168,N_24891,N_22786);
and UO_1169 (O_1169,N_21928,N_23564);
or UO_1170 (O_1170,N_24740,N_22071);
or UO_1171 (O_1171,N_22956,N_23007);
or UO_1172 (O_1172,N_22598,N_22453);
and UO_1173 (O_1173,N_23369,N_22375);
xor UO_1174 (O_1174,N_22549,N_22138);
and UO_1175 (O_1175,N_24569,N_23059);
nor UO_1176 (O_1176,N_22049,N_23908);
xnor UO_1177 (O_1177,N_23924,N_23655);
and UO_1178 (O_1178,N_23895,N_22015);
xor UO_1179 (O_1179,N_24248,N_22025);
nor UO_1180 (O_1180,N_24417,N_22546);
nor UO_1181 (O_1181,N_24015,N_23147);
nor UO_1182 (O_1182,N_22159,N_24274);
or UO_1183 (O_1183,N_23516,N_22440);
nor UO_1184 (O_1184,N_21917,N_22813);
xnor UO_1185 (O_1185,N_21877,N_23255);
nand UO_1186 (O_1186,N_23428,N_24579);
and UO_1187 (O_1187,N_23647,N_21952);
nor UO_1188 (O_1188,N_23517,N_24744);
nand UO_1189 (O_1189,N_22899,N_22827);
and UO_1190 (O_1190,N_23574,N_24502);
xnor UO_1191 (O_1191,N_24049,N_22217);
xnor UO_1192 (O_1192,N_22758,N_22643);
xnor UO_1193 (O_1193,N_22580,N_23486);
nand UO_1194 (O_1194,N_23932,N_24315);
and UO_1195 (O_1195,N_22889,N_21971);
and UO_1196 (O_1196,N_22993,N_22145);
or UO_1197 (O_1197,N_23112,N_24517);
or UO_1198 (O_1198,N_22854,N_24838);
xnor UO_1199 (O_1199,N_23105,N_23480);
nor UO_1200 (O_1200,N_22710,N_22309);
xnor UO_1201 (O_1201,N_24130,N_24844);
nor UO_1202 (O_1202,N_22491,N_22198);
and UO_1203 (O_1203,N_24568,N_24381);
nand UO_1204 (O_1204,N_23639,N_21944);
nand UO_1205 (O_1205,N_23049,N_22256);
xnor UO_1206 (O_1206,N_23741,N_22508);
or UO_1207 (O_1207,N_22800,N_22531);
or UO_1208 (O_1208,N_22480,N_23232);
and UO_1209 (O_1209,N_21976,N_24382);
nor UO_1210 (O_1210,N_22228,N_22306);
xor UO_1211 (O_1211,N_24289,N_22686);
nor UO_1212 (O_1212,N_22366,N_22111);
and UO_1213 (O_1213,N_21893,N_23537);
and UO_1214 (O_1214,N_23757,N_24055);
or UO_1215 (O_1215,N_24655,N_24314);
nand UO_1216 (O_1216,N_23443,N_24905);
nor UO_1217 (O_1217,N_24107,N_22882);
xor UO_1218 (O_1218,N_24224,N_22395);
xor UO_1219 (O_1219,N_23559,N_22206);
and UO_1220 (O_1220,N_24574,N_22954);
and UO_1221 (O_1221,N_24339,N_21977);
nand UO_1222 (O_1222,N_24650,N_23228);
nand UO_1223 (O_1223,N_23060,N_21903);
or UO_1224 (O_1224,N_23051,N_24736);
and UO_1225 (O_1225,N_23078,N_23493);
or UO_1226 (O_1226,N_23738,N_24018);
nor UO_1227 (O_1227,N_23522,N_24575);
or UO_1228 (O_1228,N_24308,N_23630);
and UO_1229 (O_1229,N_23037,N_23269);
or UO_1230 (O_1230,N_22122,N_21915);
nor UO_1231 (O_1231,N_24159,N_24287);
and UO_1232 (O_1232,N_23064,N_24037);
xor UO_1233 (O_1233,N_24741,N_22970);
nand UO_1234 (O_1234,N_22192,N_22776);
or UO_1235 (O_1235,N_24091,N_22056);
nand UO_1236 (O_1236,N_22975,N_23476);
or UO_1237 (O_1237,N_23740,N_22324);
nand UO_1238 (O_1238,N_24522,N_22585);
nor UO_1239 (O_1239,N_24983,N_24290);
xor UO_1240 (O_1240,N_22829,N_23408);
nor UO_1241 (O_1241,N_22775,N_24474);
or UO_1242 (O_1242,N_22709,N_22610);
nor UO_1243 (O_1243,N_23264,N_24027);
and UO_1244 (O_1244,N_23435,N_22923);
or UO_1245 (O_1245,N_23983,N_24764);
or UO_1246 (O_1246,N_22502,N_23445);
xor UO_1247 (O_1247,N_22210,N_24922);
xor UO_1248 (O_1248,N_23441,N_23763);
nand UO_1249 (O_1249,N_24437,N_22466);
xnor UO_1250 (O_1250,N_22890,N_23859);
nand UO_1251 (O_1251,N_24501,N_24647);
nand UO_1252 (O_1252,N_24527,N_22401);
or UO_1253 (O_1253,N_23868,N_23285);
xnor UO_1254 (O_1254,N_24798,N_22261);
and UO_1255 (O_1255,N_23047,N_22778);
nand UO_1256 (O_1256,N_23723,N_23600);
nor UO_1257 (O_1257,N_24196,N_23985);
or UO_1258 (O_1258,N_22657,N_23287);
or UO_1259 (O_1259,N_23556,N_24928);
xor UO_1260 (O_1260,N_21948,N_23145);
or UO_1261 (O_1261,N_23710,N_24331);
or UO_1262 (O_1262,N_22415,N_22855);
xor UO_1263 (O_1263,N_23987,N_24752);
nor UO_1264 (O_1264,N_23455,N_22803);
and UO_1265 (O_1265,N_24268,N_24399);
nand UO_1266 (O_1266,N_22949,N_23193);
or UO_1267 (O_1267,N_22010,N_24671);
and UO_1268 (O_1268,N_24041,N_22389);
nor UO_1269 (O_1269,N_23528,N_24839);
or UO_1270 (O_1270,N_24604,N_22166);
xor UO_1271 (O_1271,N_23325,N_23956);
or UO_1272 (O_1272,N_23784,N_22871);
nand UO_1273 (O_1273,N_23030,N_22023);
nand UO_1274 (O_1274,N_24753,N_22134);
nand UO_1275 (O_1275,N_22661,N_23693);
xnor UO_1276 (O_1276,N_24549,N_24670);
nand UO_1277 (O_1277,N_23967,N_22587);
nor UO_1278 (O_1278,N_22749,N_24535);
nand UO_1279 (O_1279,N_22872,N_24731);
nand UO_1280 (O_1280,N_22538,N_24047);
or UO_1281 (O_1281,N_23123,N_23388);
or UO_1282 (O_1282,N_23057,N_24244);
nor UO_1283 (O_1283,N_23311,N_24441);
and UO_1284 (O_1284,N_24247,N_21951);
and UO_1285 (O_1285,N_23357,N_22790);
xor UO_1286 (O_1286,N_22137,N_22612);
xor UO_1287 (O_1287,N_22050,N_23880);
nor UO_1288 (O_1288,N_24492,N_22291);
nor UO_1289 (O_1289,N_21956,N_24682);
and UO_1290 (O_1290,N_23742,N_24520);
or UO_1291 (O_1291,N_22190,N_22143);
or UO_1292 (O_1292,N_24419,N_24870);
nor UO_1293 (O_1293,N_22922,N_23790);
or UO_1294 (O_1294,N_23794,N_22442);
xnor UO_1295 (O_1295,N_24847,N_22839);
nor UO_1296 (O_1296,N_24281,N_24694);
and UO_1297 (O_1297,N_24878,N_22384);
nand UO_1298 (O_1298,N_24155,N_23829);
and UO_1299 (O_1299,N_24134,N_22603);
nor UO_1300 (O_1300,N_24328,N_23119);
nand UO_1301 (O_1301,N_23685,N_24097);
nand UO_1302 (O_1302,N_21898,N_24004);
nand UO_1303 (O_1303,N_22132,N_23065);
or UO_1304 (O_1304,N_24857,N_23259);
nand UO_1305 (O_1305,N_23573,N_23453);
and UO_1306 (O_1306,N_22030,N_23911);
nand UO_1307 (O_1307,N_23048,N_23182);
nand UO_1308 (O_1308,N_22040,N_23606);
nor UO_1309 (O_1309,N_24017,N_23305);
or UO_1310 (O_1310,N_22763,N_24128);
or UO_1311 (O_1311,N_24640,N_23681);
or UO_1312 (O_1312,N_22160,N_22197);
or UO_1313 (O_1313,N_24162,N_23279);
xor UO_1314 (O_1314,N_23581,N_23960);
xnor UO_1315 (O_1315,N_22057,N_23332);
xnor UO_1316 (O_1316,N_22454,N_22482);
and UO_1317 (O_1317,N_22457,N_22503);
and UO_1318 (O_1318,N_23823,N_22364);
xor UO_1319 (O_1319,N_23875,N_24420);
and UO_1320 (O_1320,N_24042,N_23270);
nor UO_1321 (O_1321,N_24142,N_24076);
or UO_1322 (O_1322,N_22969,N_22463);
or UO_1323 (O_1323,N_22140,N_23355);
xor UO_1324 (O_1324,N_23380,N_22681);
xor UO_1325 (O_1325,N_24235,N_22540);
or UO_1326 (O_1326,N_24795,N_24226);
xnor UO_1327 (O_1327,N_23583,N_24387);
nor UO_1328 (O_1328,N_23943,N_22350);
xor UO_1329 (O_1329,N_22202,N_22372);
xor UO_1330 (O_1330,N_22808,N_22133);
xor UO_1331 (O_1331,N_22407,N_23818);
and UO_1332 (O_1332,N_22382,N_22979);
xnor UO_1333 (O_1333,N_23231,N_22569);
and UO_1334 (O_1334,N_21961,N_23302);
and UO_1335 (O_1335,N_24048,N_22260);
or UO_1336 (O_1336,N_23206,N_22728);
nor UO_1337 (O_1337,N_23179,N_24359);
xor UO_1338 (O_1338,N_24119,N_24398);
nor UO_1339 (O_1339,N_24421,N_23251);
xnor UO_1340 (O_1340,N_22191,N_22550);
nor UO_1341 (O_1341,N_22322,N_23483);
and UO_1342 (O_1342,N_24822,N_24543);
or UO_1343 (O_1343,N_24034,N_22842);
nand UO_1344 (O_1344,N_23778,N_24044);
nand UO_1345 (O_1345,N_24292,N_23090);
nor UO_1346 (O_1346,N_24819,N_23137);
xor UO_1347 (O_1347,N_24343,N_23679);
nand UO_1348 (O_1348,N_23622,N_24646);
and UO_1349 (O_1349,N_24853,N_22517);
xor UO_1350 (O_1350,N_23468,N_23070);
and UO_1351 (O_1351,N_24654,N_24699);
nand UO_1352 (O_1352,N_24172,N_22377);
nor UO_1353 (O_1353,N_22439,N_21921);
or UO_1354 (O_1354,N_22032,N_22676);
nand UO_1355 (O_1355,N_23788,N_23968);
xnor UO_1356 (O_1356,N_24980,N_23665);
and UO_1357 (O_1357,N_21980,N_22178);
or UO_1358 (O_1358,N_23440,N_22348);
xnor UO_1359 (O_1359,N_22490,N_24635);
and UO_1360 (O_1360,N_22691,N_23491);
xor UO_1361 (O_1361,N_24313,N_23339);
nand UO_1362 (O_1362,N_23519,N_22853);
nor UO_1363 (O_1363,N_24396,N_23082);
or UO_1364 (O_1364,N_24077,N_24976);
nor UO_1365 (O_1365,N_22065,N_23889);
nor UO_1366 (O_1366,N_22027,N_24679);
nor UO_1367 (O_1367,N_23986,N_23400);
nor UO_1368 (O_1368,N_22995,N_22673);
nor UO_1369 (O_1369,N_22521,N_23646);
and UO_1370 (O_1370,N_24050,N_22942);
and UO_1371 (O_1371,N_22662,N_23869);
nor UO_1372 (O_1372,N_23557,N_22628);
or UO_1373 (O_1373,N_22082,N_23758);
xnor UO_1374 (O_1374,N_24994,N_24180);
and UO_1375 (O_1375,N_23872,N_21965);
nand UO_1376 (O_1376,N_23892,N_22034);
nand UO_1377 (O_1377,N_23870,N_24405);
nand UO_1378 (O_1378,N_23396,N_22314);
and UO_1379 (O_1379,N_24589,N_23129);
nor UO_1380 (O_1380,N_22494,N_24065);
nand UO_1381 (O_1381,N_24960,N_22773);
nand UO_1382 (O_1382,N_24138,N_24987);
nor UO_1383 (O_1383,N_23502,N_24490);
xor UO_1384 (O_1384,N_23811,N_24765);
xor UO_1385 (O_1385,N_24612,N_23404);
xor UO_1386 (O_1386,N_23737,N_24430);
nor UO_1387 (O_1387,N_24540,N_22170);
and UO_1388 (O_1388,N_24914,N_22573);
xor UO_1389 (O_1389,N_22980,N_22060);
xor UO_1390 (O_1390,N_24383,N_23091);
xor UO_1391 (O_1391,N_23979,N_24363);
xor UO_1392 (O_1392,N_23156,N_22955);
nor UO_1393 (O_1393,N_21967,N_22563);
or UO_1394 (O_1394,N_24746,N_23562);
xnor UO_1395 (O_1395,N_23641,N_22831);
or UO_1396 (O_1396,N_24272,N_22136);
nor UO_1397 (O_1397,N_22109,N_23399);
xnor UO_1398 (O_1398,N_24117,N_22613);
nor UO_1399 (O_1399,N_22594,N_23514);
xor UO_1400 (O_1400,N_23762,N_24826);
xor UO_1401 (O_1401,N_24817,N_24148);
nand UO_1402 (O_1402,N_23366,N_22935);
nand UO_1403 (O_1403,N_22755,N_22655);
nor UO_1404 (O_1404,N_23097,N_24250);
and UO_1405 (O_1405,N_24661,N_22098);
or UO_1406 (O_1406,N_24818,N_22393);
nand UO_1407 (O_1407,N_24355,N_24039);
nor UO_1408 (O_1408,N_23931,N_22862);
nand UO_1409 (O_1409,N_23898,N_23787);
or UO_1410 (O_1410,N_22222,N_24499);
xnor UO_1411 (O_1411,N_22693,N_23605);
xor UO_1412 (O_1412,N_22505,N_24087);
and UO_1413 (O_1413,N_23745,N_24340);
nand UO_1414 (O_1414,N_22354,N_22986);
nand UO_1415 (O_1415,N_22647,N_22286);
nor UO_1416 (O_1416,N_23106,N_24808);
and UO_1417 (O_1417,N_22646,N_22639);
nor UO_1418 (O_1418,N_24677,N_22568);
nor UO_1419 (O_1419,N_22431,N_24111);
and UO_1420 (O_1420,N_21970,N_23658);
nor UO_1421 (O_1421,N_24100,N_24422);
nor UO_1422 (O_1422,N_24089,N_24890);
nor UO_1423 (O_1423,N_23197,N_24410);
nor UO_1424 (O_1424,N_22495,N_24239);
nand UO_1425 (O_1425,N_24369,N_24954);
xnor UO_1426 (O_1426,N_22913,N_24754);
and UO_1427 (O_1427,N_22599,N_24751);
nand UO_1428 (O_1428,N_22156,N_24700);
nand UO_1429 (O_1429,N_24876,N_24629);
nor UO_1430 (O_1430,N_24886,N_21901);
nor UO_1431 (O_1431,N_23850,N_23406);
or UO_1432 (O_1432,N_23904,N_24758);
nand UO_1433 (O_1433,N_23964,N_22716);
nand UO_1434 (O_1434,N_23772,N_21878);
nand UO_1435 (O_1435,N_22811,N_23937);
nor UO_1436 (O_1436,N_24404,N_22320);
or UO_1437 (O_1437,N_24918,N_24423);
xnor UO_1438 (O_1438,N_22152,N_22644);
xnor UO_1439 (O_1439,N_22342,N_24920);
nand UO_1440 (O_1440,N_24099,N_23062);
or UO_1441 (O_1441,N_24170,N_24610);
and UO_1442 (O_1442,N_23293,N_22616);
nand UO_1443 (O_1443,N_23422,N_23304);
nor UO_1444 (O_1444,N_22994,N_22365);
nor UO_1445 (O_1445,N_22121,N_23258);
and UO_1446 (O_1446,N_22441,N_22633);
or UO_1447 (O_1447,N_24774,N_24761);
or UO_1448 (O_1448,N_24935,N_24507);
or UO_1449 (O_1449,N_24153,N_23883);
nand UO_1450 (O_1450,N_23863,N_22727);
nor UO_1451 (O_1451,N_23802,N_23675);
or UO_1452 (O_1452,N_24105,N_24668);
or UO_1453 (O_1453,N_24763,N_23313);
and UO_1454 (O_1454,N_23028,N_22186);
nor UO_1455 (O_1455,N_24124,N_23001);
nand UO_1456 (O_1456,N_23836,N_24262);
or UO_1457 (O_1457,N_22009,N_21879);
nor UO_1458 (O_1458,N_24388,N_23825);
nand UO_1459 (O_1459,N_22200,N_23252);
nand UO_1460 (O_1460,N_23188,N_23488);
xnor UO_1461 (O_1461,N_22706,N_23621);
and UO_1462 (O_1462,N_23759,N_22851);
and UO_1463 (O_1463,N_23586,N_24154);
and UO_1464 (O_1464,N_24631,N_23092);
and UO_1465 (O_1465,N_24936,N_24332);
and UO_1466 (O_1466,N_21911,N_24759);
xnor UO_1467 (O_1467,N_24962,N_24687);
and UO_1468 (O_1468,N_23331,N_22411);
and UO_1469 (O_1469,N_22472,N_24057);
xor UO_1470 (O_1470,N_22859,N_21902);
or UO_1471 (O_1471,N_22830,N_23027);
nor UO_1472 (O_1472,N_23713,N_22834);
nand UO_1473 (O_1473,N_24031,N_23789);
or UO_1474 (O_1474,N_24851,N_24733);
nor UO_1475 (O_1475,N_23702,N_23168);
nor UO_1476 (O_1476,N_22998,N_22449);
or UO_1477 (O_1477,N_22234,N_23551);
nor UO_1478 (O_1478,N_23998,N_23578);
nand UO_1479 (O_1479,N_23565,N_23407);
and UO_1480 (O_1480,N_21989,N_23949);
xnor UO_1481 (O_1481,N_23089,N_23128);
nand UO_1482 (O_1482,N_23827,N_22477);
and UO_1483 (O_1483,N_23572,N_24748);
or UO_1484 (O_1484,N_22966,N_23554);
and UO_1485 (O_1485,N_23515,N_22952);
nor UO_1486 (O_1486,N_24432,N_24210);
nand UO_1487 (O_1487,N_23837,N_23839);
and UO_1488 (O_1488,N_23219,N_23375);
nand UO_1489 (O_1489,N_24673,N_24426);
and UO_1490 (O_1490,N_23780,N_23625);
xnor UO_1491 (O_1491,N_24221,N_24062);
nor UO_1492 (O_1492,N_23832,N_23672);
nand UO_1493 (O_1493,N_22391,N_23769);
and UO_1494 (O_1494,N_22504,N_23570);
xor UO_1495 (O_1495,N_21920,N_24686);
or UO_1496 (O_1496,N_22295,N_23126);
nor UO_1497 (O_1497,N_22771,N_22168);
xor UO_1498 (O_1498,N_21894,N_21987);
nor UO_1499 (O_1499,N_23072,N_22357);
nor UO_1500 (O_1500,N_23671,N_24201);
nand UO_1501 (O_1501,N_23923,N_23944);
nand UO_1502 (O_1502,N_24392,N_23660);
xor UO_1503 (O_1503,N_24924,N_22637);
or UO_1504 (O_1504,N_24895,N_23239);
xor UO_1505 (O_1505,N_23878,N_24707);
and UO_1506 (O_1506,N_23958,N_24395);
xnor UO_1507 (O_1507,N_22968,N_23454);
or UO_1508 (O_1508,N_22900,N_24360);
nor UO_1509 (O_1509,N_24477,N_24252);
nand UO_1510 (O_1510,N_23764,N_23164);
xor UO_1511 (O_1511,N_24482,N_24032);
xor UO_1512 (O_1512,N_23417,N_22875);
xor UO_1513 (O_1513,N_23456,N_22101);
nand UO_1514 (O_1514,N_23902,N_23678);
xor UO_1515 (O_1515,N_23777,N_23867);
and UO_1516 (O_1516,N_23499,N_23213);
xnor UO_1517 (O_1517,N_24183,N_22614);
nor UO_1518 (O_1518,N_22930,N_24168);
nand UO_1519 (O_1519,N_24276,N_22885);
or UO_1520 (O_1520,N_24136,N_22512);
xnor UO_1521 (O_1521,N_23966,N_23806);
nor UO_1522 (O_1522,N_22215,N_22634);
nor UO_1523 (O_1523,N_22388,N_22705);
nor UO_1524 (O_1524,N_23613,N_24562);
or UO_1525 (O_1525,N_21933,N_24875);
and UO_1526 (O_1526,N_24606,N_24457);
xnor UO_1527 (O_1527,N_23644,N_23894);
xor UO_1528 (O_1528,N_24997,N_24836);
nand UO_1529 (O_1529,N_24072,N_23901);
nor UO_1530 (O_1530,N_23858,N_23804);
and UO_1531 (O_1531,N_23807,N_22607);
or UO_1532 (O_1532,N_23699,N_24504);
or UO_1533 (O_1533,N_23289,N_24390);
nand UO_1534 (O_1534,N_21925,N_24165);
xor UO_1535 (O_1535,N_21876,N_23294);
nand UO_1536 (O_1536,N_23256,N_24904);
nand UO_1537 (O_1537,N_22293,N_22283);
nor UO_1538 (O_1538,N_24664,N_24554);
and UO_1539 (O_1539,N_21974,N_23552);
and UO_1540 (O_1540,N_23243,N_23146);
xnor UO_1541 (O_1541,N_22582,N_23174);
or UO_1542 (O_1542,N_24877,N_22184);
xnor UO_1543 (O_1543,N_24718,N_22483);
or UO_1544 (O_1544,N_22828,N_23594);
or UO_1545 (O_1545,N_24361,N_22933);
and UO_1546 (O_1546,N_22212,N_23022);
or UO_1547 (O_1547,N_23330,N_23095);
nor UO_1548 (O_1548,N_23314,N_22879);
and UO_1549 (O_1549,N_24088,N_24228);
xor UO_1550 (O_1550,N_22233,N_24973);
and UO_1551 (O_1551,N_24307,N_23345);
and UO_1552 (O_1552,N_23356,N_21990);
nand UO_1553 (O_1553,N_23950,N_23283);
nand UO_1554 (O_1554,N_24167,N_22816);
nor UO_1555 (O_1555,N_22560,N_24085);
xnor UO_1556 (O_1556,N_23874,N_23130);
or UO_1557 (O_1557,N_24229,N_23192);
nand UO_1558 (O_1558,N_23389,N_22409);
or UO_1559 (O_1559,N_22069,N_24451);
nor UO_1560 (O_1560,N_23165,N_24734);
and UO_1561 (O_1561,N_22112,N_23329);
xnor UO_1562 (O_1562,N_23503,N_24197);
and UO_1563 (O_1563,N_22744,N_22517);
xor UO_1564 (O_1564,N_23097,N_23217);
xor UO_1565 (O_1565,N_23577,N_24208);
and UO_1566 (O_1566,N_24007,N_23764);
xnor UO_1567 (O_1567,N_23927,N_24911);
and UO_1568 (O_1568,N_24177,N_24922);
nand UO_1569 (O_1569,N_22420,N_24000);
nand UO_1570 (O_1570,N_23825,N_24203);
nand UO_1571 (O_1571,N_22736,N_22939);
nand UO_1572 (O_1572,N_22892,N_24329);
and UO_1573 (O_1573,N_23869,N_24530);
nor UO_1574 (O_1574,N_22175,N_23782);
or UO_1575 (O_1575,N_22488,N_24583);
nand UO_1576 (O_1576,N_22661,N_23186);
nor UO_1577 (O_1577,N_21939,N_22551);
or UO_1578 (O_1578,N_22286,N_23472);
xnor UO_1579 (O_1579,N_24048,N_22842);
nand UO_1580 (O_1580,N_23534,N_23584);
xnor UO_1581 (O_1581,N_22972,N_23553);
and UO_1582 (O_1582,N_22884,N_23007);
nor UO_1583 (O_1583,N_22794,N_24959);
nand UO_1584 (O_1584,N_22929,N_22640);
xor UO_1585 (O_1585,N_22871,N_23434);
and UO_1586 (O_1586,N_22684,N_22443);
nor UO_1587 (O_1587,N_23749,N_22820);
nand UO_1588 (O_1588,N_24313,N_23522);
xnor UO_1589 (O_1589,N_24594,N_24635);
or UO_1590 (O_1590,N_24615,N_22677);
xor UO_1591 (O_1591,N_23109,N_24619);
nand UO_1592 (O_1592,N_21926,N_22470);
and UO_1593 (O_1593,N_22903,N_24081);
nand UO_1594 (O_1594,N_23592,N_24123);
xnor UO_1595 (O_1595,N_22369,N_23793);
or UO_1596 (O_1596,N_23421,N_24659);
and UO_1597 (O_1597,N_22411,N_23383);
and UO_1598 (O_1598,N_22663,N_24612);
and UO_1599 (O_1599,N_24377,N_23738);
or UO_1600 (O_1600,N_24182,N_24301);
xnor UO_1601 (O_1601,N_23504,N_24822);
or UO_1602 (O_1602,N_24525,N_23070);
xor UO_1603 (O_1603,N_23165,N_23955);
or UO_1604 (O_1604,N_24148,N_24325);
nor UO_1605 (O_1605,N_23363,N_24794);
nor UO_1606 (O_1606,N_23226,N_24376);
or UO_1607 (O_1607,N_22575,N_24605);
nor UO_1608 (O_1608,N_23310,N_23467);
and UO_1609 (O_1609,N_22613,N_23187);
xor UO_1610 (O_1610,N_23084,N_23621);
xor UO_1611 (O_1611,N_24606,N_22000);
and UO_1612 (O_1612,N_22085,N_24117);
nor UO_1613 (O_1613,N_23681,N_22412);
and UO_1614 (O_1614,N_23287,N_23040);
nor UO_1615 (O_1615,N_22004,N_22534);
or UO_1616 (O_1616,N_24302,N_23330);
or UO_1617 (O_1617,N_22730,N_24059);
and UO_1618 (O_1618,N_23312,N_23297);
nand UO_1619 (O_1619,N_21987,N_23622);
nand UO_1620 (O_1620,N_24031,N_23307);
and UO_1621 (O_1621,N_22860,N_23997);
and UO_1622 (O_1622,N_23054,N_22902);
or UO_1623 (O_1623,N_24851,N_22130);
and UO_1624 (O_1624,N_24518,N_23149);
nor UO_1625 (O_1625,N_23173,N_23677);
or UO_1626 (O_1626,N_23288,N_24636);
nand UO_1627 (O_1627,N_23986,N_23817);
nand UO_1628 (O_1628,N_24674,N_24576);
xor UO_1629 (O_1629,N_24965,N_23168);
nor UO_1630 (O_1630,N_22512,N_22675);
nand UO_1631 (O_1631,N_23431,N_22823);
nor UO_1632 (O_1632,N_24393,N_24608);
and UO_1633 (O_1633,N_24184,N_22620);
or UO_1634 (O_1634,N_22755,N_23272);
nand UO_1635 (O_1635,N_22736,N_23980);
nand UO_1636 (O_1636,N_22005,N_23584);
and UO_1637 (O_1637,N_22127,N_22460);
and UO_1638 (O_1638,N_22035,N_24389);
or UO_1639 (O_1639,N_22192,N_24418);
or UO_1640 (O_1640,N_24124,N_22010);
or UO_1641 (O_1641,N_23101,N_23702);
nor UO_1642 (O_1642,N_23302,N_24453);
and UO_1643 (O_1643,N_23981,N_24577);
and UO_1644 (O_1644,N_23603,N_24171);
nor UO_1645 (O_1645,N_23705,N_24764);
and UO_1646 (O_1646,N_23774,N_22765);
and UO_1647 (O_1647,N_22378,N_24045);
xor UO_1648 (O_1648,N_24866,N_22628);
nand UO_1649 (O_1649,N_24103,N_21884);
or UO_1650 (O_1650,N_24785,N_23635);
or UO_1651 (O_1651,N_24840,N_24277);
and UO_1652 (O_1652,N_24831,N_22021);
nor UO_1653 (O_1653,N_24075,N_24307);
xor UO_1654 (O_1654,N_22445,N_24435);
xnor UO_1655 (O_1655,N_24921,N_23727);
or UO_1656 (O_1656,N_24074,N_24049);
nor UO_1657 (O_1657,N_23764,N_23002);
nor UO_1658 (O_1658,N_24060,N_23377);
nand UO_1659 (O_1659,N_24097,N_23932);
nor UO_1660 (O_1660,N_21956,N_23185);
xor UO_1661 (O_1661,N_23304,N_22208);
xnor UO_1662 (O_1662,N_23716,N_23937);
nand UO_1663 (O_1663,N_23817,N_24639);
or UO_1664 (O_1664,N_22908,N_24564);
xor UO_1665 (O_1665,N_24496,N_24473);
and UO_1666 (O_1666,N_23680,N_22699);
or UO_1667 (O_1667,N_24797,N_24800);
nor UO_1668 (O_1668,N_22110,N_23571);
nor UO_1669 (O_1669,N_24643,N_24938);
nor UO_1670 (O_1670,N_24259,N_23857);
and UO_1671 (O_1671,N_24936,N_23513);
nand UO_1672 (O_1672,N_22669,N_24783);
xor UO_1673 (O_1673,N_23092,N_23313);
nor UO_1674 (O_1674,N_24130,N_24252);
nand UO_1675 (O_1675,N_22010,N_22489);
xnor UO_1676 (O_1676,N_23335,N_23407);
or UO_1677 (O_1677,N_23860,N_23430);
and UO_1678 (O_1678,N_23529,N_22820);
or UO_1679 (O_1679,N_22336,N_24380);
xor UO_1680 (O_1680,N_21901,N_24337);
nor UO_1681 (O_1681,N_23897,N_22322);
or UO_1682 (O_1682,N_23162,N_24729);
nand UO_1683 (O_1683,N_22584,N_24833);
or UO_1684 (O_1684,N_24123,N_24619);
xnor UO_1685 (O_1685,N_22152,N_24466);
xnor UO_1686 (O_1686,N_24551,N_24495);
xnor UO_1687 (O_1687,N_24733,N_24277);
xor UO_1688 (O_1688,N_24685,N_22778);
or UO_1689 (O_1689,N_22790,N_23497);
nand UO_1690 (O_1690,N_24509,N_22615);
xnor UO_1691 (O_1691,N_21891,N_23241);
and UO_1692 (O_1692,N_22095,N_23075);
or UO_1693 (O_1693,N_23131,N_22100);
and UO_1694 (O_1694,N_24937,N_22771);
and UO_1695 (O_1695,N_23065,N_21924);
or UO_1696 (O_1696,N_24795,N_23411);
xor UO_1697 (O_1697,N_22941,N_24306);
nor UO_1698 (O_1698,N_23173,N_24219);
and UO_1699 (O_1699,N_21939,N_22612);
nand UO_1700 (O_1700,N_24927,N_22681);
nand UO_1701 (O_1701,N_24566,N_22290);
nand UO_1702 (O_1702,N_22183,N_24365);
or UO_1703 (O_1703,N_24929,N_22924);
nand UO_1704 (O_1704,N_23371,N_23957);
and UO_1705 (O_1705,N_23342,N_23522);
xnor UO_1706 (O_1706,N_23683,N_24747);
or UO_1707 (O_1707,N_24641,N_22705);
nand UO_1708 (O_1708,N_22727,N_22693);
or UO_1709 (O_1709,N_24361,N_22987);
or UO_1710 (O_1710,N_23131,N_22905);
nand UO_1711 (O_1711,N_23056,N_23958);
nand UO_1712 (O_1712,N_24536,N_23431);
and UO_1713 (O_1713,N_22021,N_23151);
nor UO_1714 (O_1714,N_24474,N_22528);
nor UO_1715 (O_1715,N_23914,N_23430);
xor UO_1716 (O_1716,N_23260,N_23473);
xnor UO_1717 (O_1717,N_23438,N_24512);
nor UO_1718 (O_1718,N_23778,N_24917);
nor UO_1719 (O_1719,N_23885,N_23470);
xor UO_1720 (O_1720,N_23216,N_23109);
nor UO_1721 (O_1721,N_22678,N_23059);
and UO_1722 (O_1722,N_23441,N_24050);
nor UO_1723 (O_1723,N_24959,N_23857);
nor UO_1724 (O_1724,N_22601,N_23759);
nor UO_1725 (O_1725,N_23636,N_24683);
and UO_1726 (O_1726,N_22657,N_22513);
or UO_1727 (O_1727,N_23361,N_22051);
nand UO_1728 (O_1728,N_22263,N_23171);
nand UO_1729 (O_1729,N_23271,N_23108);
xnor UO_1730 (O_1730,N_24127,N_24771);
and UO_1731 (O_1731,N_23491,N_24382);
xnor UO_1732 (O_1732,N_23171,N_24023);
nand UO_1733 (O_1733,N_24233,N_22114);
nor UO_1734 (O_1734,N_24126,N_23683);
nand UO_1735 (O_1735,N_24664,N_24458);
and UO_1736 (O_1736,N_24103,N_22310);
or UO_1737 (O_1737,N_22584,N_23001);
and UO_1738 (O_1738,N_24457,N_24195);
nand UO_1739 (O_1739,N_24095,N_22110);
nor UO_1740 (O_1740,N_24378,N_22021);
or UO_1741 (O_1741,N_24888,N_23976);
and UO_1742 (O_1742,N_24736,N_22194);
xnor UO_1743 (O_1743,N_24323,N_23513);
xor UO_1744 (O_1744,N_21975,N_22878);
and UO_1745 (O_1745,N_22953,N_24295);
or UO_1746 (O_1746,N_24407,N_23226);
nor UO_1747 (O_1747,N_24332,N_22511);
and UO_1748 (O_1748,N_24815,N_24198);
and UO_1749 (O_1749,N_23772,N_24560);
or UO_1750 (O_1750,N_23325,N_24413);
and UO_1751 (O_1751,N_23724,N_23329);
and UO_1752 (O_1752,N_22701,N_22206);
nor UO_1753 (O_1753,N_24598,N_24996);
xor UO_1754 (O_1754,N_23295,N_22273);
nand UO_1755 (O_1755,N_24625,N_24218);
and UO_1756 (O_1756,N_22247,N_23463);
xor UO_1757 (O_1757,N_23987,N_24808);
or UO_1758 (O_1758,N_22852,N_24898);
nor UO_1759 (O_1759,N_24733,N_24883);
nor UO_1760 (O_1760,N_22067,N_22314);
or UO_1761 (O_1761,N_23373,N_24937);
and UO_1762 (O_1762,N_22383,N_24603);
xor UO_1763 (O_1763,N_23112,N_22555);
nand UO_1764 (O_1764,N_23303,N_23236);
and UO_1765 (O_1765,N_22843,N_23837);
and UO_1766 (O_1766,N_24879,N_21936);
nand UO_1767 (O_1767,N_24000,N_22592);
or UO_1768 (O_1768,N_24461,N_22670);
nor UO_1769 (O_1769,N_23890,N_22942);
nor UO_1770 (O_1770,N_23281,N_23765);
xor UO_1771 (O_1771,N_21918,N_22692);
and UO_1772 (O_1772,N_22885,N_24503);
nand UO_1773 (O_1773,N_24502,N_23316);
xor UO_1774 (O_1774,N_23392,N_24706);
nand UO_1775 (O_1775,N_23088,N_22343);
nand UO_1776 (O_1776,N_22612,N_22545);
or UO_1777 (O_1777,N_22274,N_23796);
and UO_1778 (O_1778,N_21940,N_23230);
and UO_1779 (O_1779,N_22916,N_21938);
xnor UO_1780 (O_1780,N_23601,N_21917);
and UO_1781 (O_1781,N_23909,N_23921);
and UO_1782 (O_1782,N_23225,N_23940);
nand UO_1783 (O_1783,N_24702,N_22530);
xnor UO_1784 (O_1784,N_23944,N_23951);
or UO_1785 (O_1785,N_23049,N_24665);
nand UO_1786 (O_1786,N_24589,N_24777);
nand UO_1787 (O_1787,N_24717,N_23160);
or UO_1788 (O_1788,N_23180,N_23861);
or UO_1789 (O_1789,N_23171,N_24589);
or UO_1790 (O_1790,N_22611,N_22933);
nand UO_1791 (O_1791,N_22353,N_22572);
xor UO_1792 (O_1792,N_24851,N_24651);
and UO_1793 (O_1793,N_24255,N_22652);
and UO_1794 (O_1794,N_24844,N_22107);
nor UO_1795 (O_1795,N_23873,N_23619);
or UO_1796 (O_1796,N_21899,N_22197);
or UO_1797 (O_1797,N_22211,N_24785);
xnor UO_1798 (O_1798,N_23672,N_23771);
xnor UO_1799 (O_1799,N_22762,N_22488);
or UO_1800 (O_1800,N_22096,N_24413);
xnor UO_1801 (O_1801,N_24330,N_21924);
nor UO_1802 (O_1802,N_22366,N_22439);
xnor UO_1803 (O_1803,N_24327,N_22104);
and UO_1804 (O_1804,N_22068,N_22557);
or UO_1805 (O_1805,N_23939,N_23370);
xnor UO_1806 (O_1806,N_22210,N_24447);
nor UO_1807 (O_1807,N_24959,N_22545);
xnor UO_1808 (O_1808,N_24970,N_24987);
and UO_1809 (O_1809,N_22430,N_24898);
and UO_1810 (O_1810,N_24754,N_24688);
xor UO_1811 (O_1811,N_22608,N_22816);
nand UO_1812 (O_1812,N_24346,N_22597);
or UO_1813 (O_1813,N_22614,N_23719);
xor UO_1814 (O_1814,N_22335,N_22433);
xor UO_1815 (O_1815,N_22996,N_22753);
nand UO_1816 (O_1816,N_24481,N_23378);
and UO_1817 (O_1817,N_24177,N_24781);
nand UO_1818 (O_1818,N_22553,N_24222);
xor UO_1819 (O_1819,N_22235,N_23396);
or UO_1820 (O_1820,N_22368,N_24432);
nor UO_1821 (O_1821,N_24216,N_22160);
nand UO_1822 (O_1822,N_23693,N_22996);
xor UO_1823 (O_1823,N_22795,N_23153);
nor UO_1824 (O_1824,N_23489,N_22816);
nor UO_1825 (O_1825,N_22208,N_24998);
xor UO_1826 (O_1826,N_23088,N_23229);
or UO_1827 (O_1827,N_23755,N_24667);
and UO_1828 (O_1828,N_22330,N_23301);
nor UO_1829 (O_1829,N_22188,N_22493);
xnor UO_1830 (O_1830,N_24953,N_23757);
or UO_1831 (O_1831,N_23087,N_23475);
xor UO_1832 (O_1832,N_24519,N_24282);
or UO_1833 (O_1833,N_23612,N_24451);
and UO_1834 (O_1834,N_23209,N_23731);
xnor UO_1835 (O_1835,N_22100,N_22002);
and UO_1836 (O_1836,N_24539,N_24926);
or UO_1837 (O_1837,N_23953,N_23276);
xor UO_1838 (O_1838,N_23197,N_22864);
xor UO_1839 (O_1839,N_23288,N_23950);
or UO_1840 (O_1840,N_23978,N_24948);
nor UO_1841 (O_1841,N_24798,N_22947);
xor UO_1842 (O_1842,N_24141,N_22917);
or UO_1843 (O_1843,N_23375,N_24859);
and UO_1844 (O_1844,N_24047,N_22524);
nand UO_1845 (O_1845,N_22480,N_23451);
xnor UO_1846 (O_1846,N_23562,N_23383);
nand UO_1847 (O_1847,N_23424,N_21951);
nor UO_1848 (O_1848,N_23935,N_23096);
nand UO_1849 (O_1849,N_24225,N_24304);
nand UO_1850 (O_1850,N_22339,N_22903);
xor UO_1851 (O_1851,N_24158,N_24583);
xnor UO_1852 (O_1852,N_24232,N_23514);
xor UO_1853 (O_1853,N_22976,N_22368);
and UO_1854 (O_1854,N_24768,N_24985);
nor UO_1855 (O_1855,N_23049,N_23340);
xnor UO_1856 (O_1856,N_23646,N_22940);
or UO_1857 (O_1857,N_22267,N_23964);
nand UO_1858 (O_1858,N_23847,N_23856);
or UO_1859 (O_1859,N_24379,N_24621);
xnor UO_1860 (O_1860,N_24896,N_22857);
or UO_1861 (O_1861,N_23212,N_24226);
or UO_1862 (O_1862,N_23060,N_22730);
xnor UO_1863 (O_1863,N_24357,N_23023);
xnor UO_1864 (O_1864,N_24744,N_23958);
xor UO_1865 (O_1865,N_22039,N_24572);
nand UO_1866 (O_1866,N_24817,N_23459);
and UO_1867 (O_1867,N_22725,N_24637);
nand UO_1868 (O_1868,N_22778,N_22142);
nor UO_1869 (O_1869,N_21893,N_24600);
or UO_1870 (O_1870,N_24044,N_22044);
nand UO_1871 (O_1871,N_23759,N_22493);
or UO_1872 (O_1872,N_22117,N_21941);
nor UO_1873 (O_1873,N_22796,N_22063);
or UO_1874 (O_1874,N_23156,N_22755);
or UO_1875 (O_1875,N_22099,N_22045);
nor UO_1876 (O_1876,N_22826,N_22893);
xnor UO_1877 (O_1877,N_24228,N_22310);
or UO_1878 (O_1878,N_22004,N_24024);
or UO_1879 (O_1879,N_22202,N_22063);
xor UO_1880 (O_1880,N_24714,N_23659);
xor UO_1881 (O_1881,N_23732,N_23883);
or UO_1882 (O_1882,N_22895,N_22675);
or UO_1883 (O_1883,N_23454,N_24260);
xnor UO_1884 (O_1884,N_23804,N_24618);
xor UO_1885 (O_1885,N_22837,N_23473);
xnor UO_1886 (O_1886,N_23212,N_24668);
and UO_1887 (O_1887,N_24766,N_23507);
xor UO_1888 (O_1888,N_22792,N_24264);
or UO_1889 (O_1889,N_24573,N_23009);
and UO_1890 (O_1890,N_24101,N_23224);
and UO_1891 (O_1891,N_23741,N_22794);
nand UO_1892 (O_1892,N_23241,N_24564);
xnor UO_1893 (O_1893,N_22470,N_24469);
and UO_1894 (O_1894,N_24151,N_23907);
nor UO_1895 (O_1895,N_24429,N_22206);
or UO_1896 (O_1896,N_23774,N_23078);
nand UO_1897 (O_1897,N_22598,N_23749);
xor UO_1898 (O_1898,N_24392,N_24518);
nor UO_1899 (O_1899,N_22301,N_22039);
nor UO_1900 (O_1900,N_24580,N_23697);
or UO_1901 (O_1901,N_22662,N_23179);
nor UO_1902 (O_1902,N_22886,N_23304);
and UO_1903 (O_1903,N_23673,N_23568);
or UO_1904 (O_1904,N_23483,N_24840);
xnor UO_1905 (O_1905,N_23066,N_22862);
and UO_1906 (O_1906,N_23337,N_22302);
nor UO_1907 (O_1907,N_22620,N_24417);
or UO_1908 (O_1908,N_23630,N_23567);
xor UO_1909 (O_1909,N_22987,N_23159);
or UO_1910 (O_1910,N_23218,N_23166);
and UO_1911 (O_1911,N_23273,N_22342);
and UO_1912 (O_1912,N_22521,N_23104);
nand UO_1913 (O_1913,N_24334,N_23449);
nand UO_1914 (O_1914,N_24354,N_23200);
nand UO_1915 (O_1915,N_22150,N_22088);
nand UO_1916 (O_1916,N_23705,N_23961);
nand UO_1917 (O_1917,N_24970,N_22268);
nor UO_1918 (O_1918,N_22979,N_22327);
xor UO_1919 (O_1919,N_22026,N_23477);
xor UO_1920 (O_1920,N_23088,N_24840);
xnor UO_1921 (O_1921,N_24413,N_24956);
nand UO_1922 (O_1922,N_24308,N_24741);
nand UO_1923 (O_1923,N_23549,N_24403);
nand UO_1924 (O_1924,N_24635,N_24571);
and UO_1925 (O_1925,N_22455,N_24175);
xnor UO_1926 (O_1926,N_24004,N_22457);
xor UO_1927 (O_1927,N_24112,N_22513);
and UO_1928 (O_1928,N_23209,N_23166);
or UO_1929 (O_1929,N_24947,N_22928);
and UO_1930 (O_1930,N_24964,N_23664);
xnor UO_1931 (O_1931,N_24805,N_23513);
and UO_1932 (O_1932,N_22101,N_24344);
xnor UO_1933 (O_1933,N_22382,N_22747);
and UO_1934 (O_1934,N_24289,N_23636);
and UO_1935 (O_1935,N_22528,N_21938);
and UO_1936 (O_1936,N_24659,N_23411);
nor UO_1937 (O_1937,N_23293,N_22938);
nor UO_1938 (O_1938,N_23598,N_23265);
or UO_1939 (O_1939,N_24299,N_24762);
and UO_1940 (O_1940,N_23332,N_22870);
and UO_1941 (O_1941,N_22944,N_23452);
nand UO_1942 (O_1942,N_22885,N_24315);
and UO_1943 (O_1943,N_24357,N_24358);
xor UO_1944 (O_1944,N_24382,N_23964);
xnor UO_1945 (O_1945,N_23917,N_24233);
and UO_1946 (O_1946,N_24785,N_23852);
nor UO_1947 (O_1947,N_24337,N_24868);
xnor UO_1948 (O_1948,N_22903,N_22119);
xor UO_1949 (O_1949,N_23792,N_24796);
nor UO_1950 (O_1950,N_24929,N_24150);
or UO_1951 (O_1951,N_24754,N_24877);
nand UO_1952 (O_1952,N_22181,N_24271);
nor UO_1953 (O_1953,N_23514,N_22302);
and UO_1954 (O_1954,N_24020,N_22550);
xnor UO_1955 (O_1955,N_24667,N_22896);
and UO_1956 (O_1956,N_24039,N_22009);
nand UO_1957 (O_1957,N_24215,N_24078);
or UO_1958 (O_1958,N_23279,N_23507);
nor UO_1959 (O_1959,N_22674,N_22089);
and UO_1960 (O_1960,N_24305,N_22455);
xnor UO_1961 (O_1961,N_22357,N_24786);
nand UO_1962 (O_1962,N_22829,N_22477);
or UO_1963 (O_1963,N_22528,N_24518);
or UO_1964 (O_1964,N_22849,N_24335);
nor UO_1965 (O_1965,N_22609,N_22211);
nor UO_1966 (O_1966,N_22642,N_22492);
nor UO_1967 (O_1967,N_23756,N_24862);
or UO_1968 (O_1968,N_24606,N_23780);
nor UO_1969 (O_1969,N_24826,N_22774);
nor UO_1970 (O_1970,N_24422,N_23248);
nand UO_1971 (O_1971,N_23315,N_24332);
xor UO_1972 (O_1972,N_22457,N_24007);
nor UO_1973 (O_1973,N_22293,N_22163);
or UO_1974 (O_1974,N_23703,N_24416);
and UO_1975 (O_1975,N_24657,N_23007);
nor UO_1976 (O_1976,N_24245,N_22546);
and UO_1977 (O_1977,N_22148,N_24987);
nand UO_1978 (O_1978,N_23506,N_24285);
nand UO_1979 (O_1979,N_24994,N_23374);
xor UO_1980 (O_1980,N_23094,N_22165);
and UO_1981 (O_1981,N_24642,N_22660);
or UO_1982 (O_1982,N_24596,N_22270);
and UO_1983 (O_1983,N_22854,N_22005);
xnor UO_1984 (O_1984,N_24920,N_23686);
nor UO_1985 (O_1985,N_24126,N_23425);
or UO_1986 (O_1986,N_24641,N_24490);
nand UO_1987 (O_1987,N_23917,N_23473);
and UO_1988 (O_1988,N_24499,N_23843);
and UO_1989 (O_1989,N_22814,N_22070);
nor UO_1990 (O_1990,N_23543,N_22380);
and UO_1991 (O_1991,N_22189,N_22939);
and UO_1992 (O_1992,N_22706,N_22547);
or UO_1993 (O_1993,N_23179,N_21962);
and UO_1994 (O_1994,N_22308,N_21979);
xor UO_1995 (O_1995,N_22239,N_23256);
nor UO_1996 (O_1996,N_22053,N_24036);
nand UO_1997 (O_1997,N_23399,N_24769);
xor UO_1998 (O_1998,N_22684,N_23101);
and UO_1999 (O_1999,N_23687,N_24241);
nand UO_2000 (O_2000,N_21986,N_23863);
nand UO_2001 (O_2001,N_22336,N_24126);
nor UO_2002 (O_2002,N_24531,N_22177);
and UO_2003 (O_2003,N_23195,N_24102);
and UO_2004 (O_2004,N_23539,N_23147);
nand UO_2005 (O_2005,N_24644,N_24295);
and UO_2006 (O_2006,N_23437,N_24980);
or UO_2007 (O_2007,N_21981,N_24795);
xnor UO_2008 (O_2008,N_23631,N_24150);
or UO_2009 (O_2009,N_23072,N_23574);
nand UO_2010 (O_2010,N_22882,N_22161);
and UO_2011 (O_2011,N_24987,N_22243);
or UO_2012 (O_2012,N_23904,N_22852);
nand UO_2013 (O_2013,N_21910,N_24887);
nand UO_2014 (O_2014,N_24160,N_22372);
nand UO_2015 (O_2015,N_22625,N_22285);
or UO_2016 (O_2016,N_22854,N_23768);
xnor UO_2017 (O_2017,N_22448,N_23236);
xnor UO_2018 (O_2018,N_24293,N_24163);
nand UO_2019 (O_2019,N_24795,N_23802);
xnor UO_2020 (O_2020,N_23640,N_21915);
and UO_2021 (O_2021,N_23342,N_22215);
xor UO_2022 (O_2022,N_22740,N_22494);
nor UO_2023 (O_2023,N_23233,N_24357);
xnor UO_2024 (O_2024,N_23215,N_22951);
or UO_2025 (O_2025,N_24793,N_24810);
nor UO_2026 (O_2026,N_24376,N_22858);
nand UO_2027 (O_2027,N_23377,N_23255);
xor UO_2028 (O_2028,N_23263,N_24933);
or UO_2029 (O_2029,N_24918,N_24673);
nor UO_2030 (O_2030,N_22692,N_23961);
nand UO_2031 (O_2031,N_24463,N_21952);
or UO_2032 (O_2032,N_24712,N_22409);
or UO_2033 (O_2033,N_22731,N_23727);
xor UO_2034 (O_2034,N_21888,N_22896);
nand UO_2035 (O_2035,N_24378,N_24980);
nand UO_2036 (O_2036,N_23376,N_24912);
xnor UO_2037 (O_2037,N_23649,N_23578);
xnor UO_2038 (O_2038,N_23297,N_22241);
and UO_2039 (O_2039,N_24681,N_23461);
xnor UO_2040 (O_2040,N_22624,N_22410);
or UO_2041 (O_2041,N_23534,N_24929);
nand UO_2042 (O_2042,N_24488,N_22278);
xnor UO_2043 (O_2043,N_24981,N_24872);
nand UO_2044 (O_2044,N_22935,N_22184);
xnor UO_2045 (O_2045,N_24690,N_23238);
nor UO_2046 (O_2046,N_23770,N_22515);
xor UO_2047 (O_2047,N_24057,N_23971);
nor UO_2048 (O_2048,N_24161,N_22185);
nand UO_2049 (O_2049,N_22185,N_23985);
and UO_2050 (O_2050,N_23381,N_22603);
nor UO_2051 (O_2051,N_22277,N_23215);
xor UO_2052 (O_2052,N_22218,N_23326);
xor UO_2053 (O_2053,N_24606,N_23139);
xnor UO_2054 (O_2054,N_22920,N_23619);
or UO_2055 (O_2055,N_23705,N_24539);
xor UO_2056 (O_2056,N_22259,N_24711);
nor UO_2057 (O_2057,N_23542,N_22807);
or UO_2058 (O_2058,N_22762,N_23855);
or UO_2059 (O_2059,N_22982,N_23030);
nand UO_2060 (O_2060,N_23389,N_24647);
or UO_2061 (O_2061,N_21978,N_23316);
xnor UO_2062 (O_2062,N_24103,N_23960);
nor UO_2063 (O_2063,N_22793,N_22493);
or UO_2064 (O_2064,N_22368,N_24970);
or UO_2065 (O_2065,N_23884,N_22094);
xnor UO_2066 (O_2066,N_24575,N_22283);
nor UO_2067 (O_2067,N_22433,N_22684);
or UO_2068 (O_2068,N_24636,N_22803);
and UO_2069 (O_2069,N_23794,N_23487);
xor UO_2070 (O_2070,N_22417,N_24647);
nand UO_2071 (O_2071,N_23302,N_24228);
or UO_2072 (O_2072,N_23795,N_23279);
nor UO_2073 (O_2073,N_23548,N_24130);
xnor UO_2074 (O_2074,N_24240,N_23849);
and UO_2075 (O_2075,N_24157,N_23654);
nand UO_2076 (O_2076,N_23165,N_24236);
or UO_2077 (O_2077,N_22458,N_22535);
nand UO_2078 (O_2078,N_23481,N_23230);
nor UO_2079 (O_2079,N_22959,N_24475);
and UO_2080 (O_2080,N_24105,N_22631);
or UO_2081 (O_2081,N_22923,N_23152);
xnor UO_2082 (O_2082,N_22143,N_24278);
nor UO_2083 (O_2083,N_22758,N_24032);
xor UO_2084 (O_2084,N_22433,N_22704);
nand UO_2085 (O_2085,N_24653,N_22440);
nand UO_2086 (O_2086,N_22288,N_22371);
nor UO_2087 (O_2087,N_24100,N_23666);
or UO_2088 (O_2088,N_22471,N_23324);
xnor UO_2089 (O_2089,N_24223,N_22246);
nor UO_2090 (O_2090,N_22383,N_24817);
nor UO_2091 (O_2091,N_22234,N_24334);
and UO_2092 (O_2092,N_24268,N_24754);
nor UO_2093 (O_2093,N_22306,N_24807);
nor UO_2094 (O_2094,N_23630,N_22305);
nor UO_2095 (O_2095,N_22617,N_22854);
xnor UO_2096 (O_2096,N_22254,N_23624);
or UO_2097 (O_2097,N_24438,N_24888);
nand UO_2098 (O_2098,N_23316,N_24069);
and UO_2099 (O_2099,N_22989,N_22119);
nor UO_2100 (O_2100,N_24442,N_22693);
and UO_2101 (O_2101,N_24291,N_23719);
nand UO_2102 (O_2102,N_24095,N_24886);
nand UO_2103 (O_2103,N_24041,N_22867);
nand UO_2104 (O_2104,N_22200,N_22510);
nor UO_2105 (O_2105,N_23448,N_22990);
nand UO_2106 (O_2106,N_23409,N_22635);
and UO_2107 (O_2107,N_23603,N_22616);
nand UO_2108 (O_2108,N_22661,N_24494);
xnor UO_2109 (O_2109,N_22387,N_23543);
or UO_2110 (O_2110,N_23384,N_24941);
or UO_2111 (O_2111,N_24516,N_24939);
or UO_2112 (O_2112,N_22797,N_24769);
nand UO_2113 (O_2113,N_22720,N_22846);
nor UO_2114 (O_2114,N_22892,N_22494);
xnor UO_2115 (O_2115,N_22275,N_22524);
and UO_2116 (O_2116,N_22913,N_22692);
and UO_2117 (O_2117,N_24429,N_23080);
xor UO_2118 (O_2118,N_23848,N_23995);
xor UO_2119 (O_2119,N_24476,N_23343);
nor UO_2120 (O_2120,N_23097,N_24862);
nor UO_2121 (O_2121,N_23151,N_24058);
or UO_2122 (O_2122,N_24160,N_22805);
nor UO_2123 (O_2123,N_23237,N_23186);
nand UO_2124 (O_2124,N_24382,N_22751);
and UO_2125 (O_2125,N_23103,N_22716);
nor UO_2126 (O_2126,N_23916,N_22100);
xnor UO_2127 (O_2127,N_23374,N_24243);
nand UO_2128 (O_2128,N_21942,N_21878);
xnor UO_2129 (O_2129,N_24647,N_23354);
nor UO_2130 (O_2130,N_24197,N_24878);
or UO_2131 (O_2131,N_23344,N_22062);
xor UO_2132 (O_2132,N_22356,N_24985);
and UO_2133 (O_2133,N_22247,N_24066);
nand UO_2134 (O_2134,N_24746,N_23741);
or UO_2135 (O_2135,N_24347,N_24114);
xnor UO_2136 (O_2136,N_22366,N_23950);
and UO_2137 (O_2137,N_21950,N_23565);
or UO_2138 (O_2138,N_21980,N_23163);
xnor UO_2139 (O_2139,N_23638,N_21914);
and UO_2140 (O_2140,N_23515,N_23510);
nor UO_2141 (O_2141,N_23432,N_24718);
or UO_2142 (O_2142,N_22928,N_24477);
and UO_2143 (O_2143,N_23801,N_22618);
and UO_2144 (O_2144,N_22390,N_24167);
or UO_2145 (O_2145,N_24442,N_23186);
xor UO_2146 (O_2146,N_24450,N_23217);
xor UO_2147 (O_2147,N_24866,N_24214);
and UO_2148 (O_2148,N_22866,N_23910);
and UO_2149 (O_2149,N_23602,N_24813);
nand UO_2150 (O_2150,N_24357,N_22252);
xor UO_2151 (O_2151,N_24154,N_22406);
and UO_2152 (O_2152,N_23823,N_22467);
xnor UO_2153 (O_2153,N_24098,N_21889);
and UO_2154 (O_2154,N_24017,N_24048);
nor UO_2155 (O_2155,N_24215,N_24664);
or UO_2156 (O_2156,N_24883,N_24050);
or UO_2157 (O_2157,N_23404,N_24755);
nor UO_2158 (O_2158,N_23616,N_24373);
nor UO_2159 (O_2159,N_23955,N_22130);
nor UO_2160 (O_2160,N_23217,N_23012);
xor UO_2161 (O_2161,N_22915,N_22706);
or UO_2162 (O_2162,N_23178,N_24834);
nand UO_2163 (O_2163,N_22602,N_24588);
xor UO_2164 (O_2164,N_24412,N_23130);
nor UO_2165 (O_2165,N_22171,N_24570);
and UO_2166 (O_2166,N_22283,N_21952);
xnor UO_2167 (O_2167,N_23850,N_22345);
or UO_2168 (O_2168,N_24411,N_23729);
nor UO_2169 (O_2169,N_24056,N_22389);
or UO_2170 (O_2170,N_23164,N_22165);
xor UO_2171 (O_2171,N_22894,N_24725);
nand UO_2172 (O_2172,N_22856,N_24317);
or UO_2173 (O_2173,N_24622,N_24516);
nand UO_2174 (O_2174,N_23530,N_22588);
nor UO_2175 (O_2175,N_22063,N_23395);
and UO_2176 (O_2176,N_22836,N_24630);
nor UO_2177 (O_2177,N_22504,N_22343);
nor UO_2178 (O_2178,N_24823,N_23449);
or UO_2179 (O_2179,N_24065,N_24921);
and UO_2180 (O_2180,N_24022,N_24053);
xnor UO_2181 (O_2181,N_23326,N_22614);
or UO_2182 (O_2182,N_22971,N_24879);
nor UO_2183 (O_2183,N_24429,N_22862);
xor UO_2184 (O_2184,N_22722,N_22272);
nand UO_2185 (O_2185,N_23791,N_23872);
or UO_2186 (O_2186,N_22493,N_23256);
nand UO_2187 (O_2187,N_22705,N_23895);
nor UO_2188 (O_2188,N_23633,N_23100);
and UO_2189 (O_2189,N_24135,N_22534);
and UO_2190 (O_2190,N_22542,N_24504);
and UO_2191 (O_2191,N_23291,N_22244);
nor UO_2192 (O_2192,N_21885,N_22353);
xor UO_2193 (O_2193,N_23446,N_22374);
xnor UO_2194 (O_2194,N_22663,N_22825);
nand UO_2195 (O_2195,N_24919,N_22137);
nand UO_2196 (O_2196,N_24686,N_22053);
and UO_2197 (O_2197,N_22503,N_22356);
and UO_2198 (O_2198,N_22263,N_23802);
xor UO_2199 (O_2199,N_23306,N_24497);
nor UO_2200 (O_2200,N_22796,N_22813);
nand UO_2201 (O_2201,N_22522,N_24132);
or UO_2202 (O_2202,N_23025,N_24980);
or UO_2203 (O_2203,N_24665,N_22505);
nand UO_2204 (O_2204,N_24131,N_24271);
xnor UO_2205 (O_2205,N_23530,N_24612);
or UO_2206 (O_2206,N_22497,N_24713);
or UO_2207 (O_2207,N_24164,N_21945);
and UO_2208 (O_2208,N_22901,N_24190);
nand UO_2209 (O_2209,N_23351,N_22855);
and UO_2210 (O_2210,N_23836,N_22512);
xor UO_2211 (O_2211,N_22951,N_22119);
and UO_2212 (O_2212,N_22832,N_22508);
nor UO_2213 (O_2213,N_23985,N_24890);
nand UO_2214 (O_2214,N_24862,N_24068);
nand UO_2215 (O_2215,N_23351,N_22734);
or UO_2216 (O_2216,N_23294,N_23218);
and UO_2217 (O_2217,N_24393,N_23582);
and UO_2218 (O_2218,N_22860,N_23004);
nor UO_2219 (O_2219,N_22922,N_22860);
and UO_2220 (O_2220,N_24345,N_24599);
and UO_2221 (O_2221,N_22272,N_22755);
xnor UO_2222 (O_2222,N_24232,N_24824);
xor UO_2223 (O_2223,N_24228,N_24083);
nor UO_2224 (O_2224,N_24822,N_23856);
nor UO_2225 (O_2225,N_21886,N_24669);
nand UO_2226 (O_2226,N_23576,N_23423);
or UO_2227 (O_2227,N_21996,N_23803);
xnor UO_2228 (O_2228,N_23867,N_23555);
and UO_2229 (O_2229,N_22237,N_22894);
and UO_2230 (O_2230,N_23629,N_22370);
nor UO_2231 (O_2231,N_23696,N_23233);
nand UO_2232 (O_2232,N_24058,N_22543);
nand UO_2233 (O_2233,N_24429,N_23541);
xor UO_2234 (O_2234,N_22357,N_22343);
and UO_2235 (O_2235,N_24064,N_21935);
and UO_2236 (O_2236,N_22971,N_24165);
xor UO_2237 (O_2237,N_23425,N_23906);
nand UO_2238 (O_2238,N_22849,N_23932);
and UO_2239 (O_2239,N_23534,N_22433);
xor UO_2240 (O_2240,N_23722,N_22683);
and UO_2241 (O_2241,N_22736,N_23407);
nand UO_2242 (O_2242,N_22327,N_22243);
nor UO_2243 (O_2243,N_22918,N_23377);
xnor UO_2244 (O_2244,N_24874,N_22440);
nand UO_2245 (O_2245,N_24143,N_24837);
nor UO_2246 (O_2246,N_24136,N_24273);
nand UO_2247 (O_2247,N_22248,N_22527);
xor UO_2248 (O_2248,N_23577,N_24910);
nand UO_2249 (O_2249,N_22267,N_24224);
xor UO_2250 (O_2250,N_23198,N_24515);
nand UO_2251 (O_2251,N_23110,N_23652);
nand UO_2252 (O_2252,N_24104,N_23193);
xor UO_2253 (O_2253,N_22595,N_22115);
and UO_2254 (O_2254,N_23595,N_22234);
or UO_2255 (O_2255,N_22553,N_23114);
xnor UO_2256 (O_2256,N_24860,N_24227);
nand UO_2257 (O_2257,N_24368,N_24181);
xor UO_2258 (O_2258,N_23723,N_22942);
or UO_2259 (O_2259,N_21904,N_23993);
xnor UO_2260 (O_2260,N_23755,N_23167);
xnor UO_2261 (O_2261,N_23060,N_22990);
xor UO_2262 (O_2262,N_23721,N_24540);
xnor UO_2263 (O_2263,N_24952,N_23088);
and UO_2264 (O_2264,N_22433,N_23101);
xor UO_2265 (O_2265,N_24686,N_24997);
nand UO_2266 (O_2266,N_24809,N_24464);
or UO_2267 (O_2267,N_24303,N_23156);
and UO_2268 (O_2268,N_22866,N_24529);
or UO_2269 (O_2269,N_23433,N_23701);
nor UO_2270 (O_2270,N_22221,N_23958);
or UO_2271 (O_2271,N_24933,N_24311);
xnor UO_2272 (O_2272,N_23501,N_23977);
xnor UO_2273 (O_2273,N_22425,N_22684);
and UO_2274 (O_2274,N_23690,N_22881);
or UO_2275 (O_2275,N_24534,N_23613);
nor UO_2276 (O_2276,N_23540,N_23774);
xor UO_2277 (O_2277,N_24946,N_23119);
or UO_2278 (O_2278,N_23423,N_23842);
nor UO_2279 (O_2279,N_23857,N_24193);
xnor UO_2280 (O_2280,N_22616,N_22301);
nor UO_2281 (O_2281,N_22395,N_24877);
nor UO_2282 (O_2282,N_23528,N_22644);
or UO_2283 (O_2283,N_24194,N_23794);
nor UO_2284 (O_2284,N_23458,N_24097);
and UO_2285 (O_2285,N_24314,N_24457);
xnor UO_2286 (O_2286,N_22592,N_24719);
or UO_2287 (O_2287,N_22254,N_22728);
xnor UO_2288 (O_2288,N_23554,N_23698);
nor UO_2289 (O_2289,N_22780,N_24159);
xnor UO_2290 (O_2290,N_24999,N_22769);
xor UO_2291 (O_2291,N_22631,N_22325);
xnor UO_2292 (O_2292,N_23740,N_23340);
or UO_2293 (O_2293,N_22956,N_23889);
or UO_2294 (O_2294,N_24342,N_24142);
and UO_2295 (O_2295,N_24655,N_24011);
xor UO_2296 (O_2296,N_24585,N_21945);
xor UO_2297 (O_2297,N_24188,N_23306);
xnor UO_2298 (O_2298,N_22218,N_23279);
nand UO_2299 (O_2299,N_21971,N_24138);
xnor UO_2300 (O_2300,N_22237,N_23313);
nand UO_2301 (O_2301,N_24711,N_21906);
nand UO_2302 (O_2302,N_22578,N_23078);
xor UO_2303 (O_2303,N_22822,N_22133);
xor UO_2304 (O_2304,N_23541,N_22736);
nand UO_2305 (O_2305,N_22391,N_22291);
nand UO_2306 (O_2306,N_22132,N_24165);
xor UO_2307 (O_2307,N_24498,N_22297);
or UO_2308 (O_2308,N_23037,N_24874);
xor UO_2309 (O_2309,N_23842,N_22696);
xnor UO_2310 (O_2310,N_24071,N_23491);
nand UO_2311 (O_2311,N_22873,N_24045);
xnor UO_2312 (O_2312,N_23873,N_24275);
nor UO_2313 (O_2313,N_22434,N_23593);
nand UO_2314 (O_2314,N_22807,N_23448);
xor UO_2315 (O_2315,N_24690,N_22899);
nand UO_2316 (O_2316,N_24053,N_24361);
and UO_2317 (O_2317,N_23051,N_24860);
and UO_2318 (O_2318,N_23677,N_23515);
nand UO_2319 (O_2319,N_23310,N_22843);
xor UO_2320 (O_2320,N_22357,N_22022);
or UO_2321 (O_2321,N_23935,N_24426);
nor UO_2322 (O_2322,N_24557,N_22471);
and UO_2323 (O_2323,N_23507,N_24125);
or UO_2324 (O_2324,N_23799,N_22920);
nand UO_2325 (O_2325,N_24310,N_24458);
nand UO_2326 (O_2326,N_24590,N_23580);
nand UO_2327 (O_2327,N_23236,N_23234);
and UO_2328 (O_2328,N_22807,N_24660);
nor UO_2329 (O_2329,N_24305,N_22378);
nand UO_2330 (O_2330,N_22958,N_22715);
and UO_2331 (O_2331,N_24806,N_23620);
and UO_2332 (O_2332,N_24142,N_22841);
or UO_2333 (O_2333,N_23257,N_22691);
nand UO_2334 (O_2334,N_23420,N_22967);
nor UO_2335 (O_2335,N_24758,N_22180);
or UO_2336 (O_2336,N_21890,N_23871);
nor UO_2337 (O_2337,N_23649,N_23391);
or UO_2338 (O_2338,N_22458,N_23828);
xnor UO_2339 (O_2339,N_24873,N_24156);
or UO_2340 (O_2340,N_24161,N_24572);
and UO_2341 (O_2341,N_22226,N_23490);
nor UO_2342 (O_2342,N_23598,N_24946);
xor UO_2343 (O_2343,N_22275,N_23909);
and UO_2344 (O_2344,N_22524,N_23043);
or UO_2345 (O_2345,N_22750,N_22627);
or UO_2346 (O_2346,N_23590,N_22193);
nand UO_2347 (O_2347,N_23748,N_23905);
xnor UO_2348 (O_2348,N_23552,N_22030);
nand UO_2349 (O_2349,N_23997,N_24470);
or UO_2350 (O_2350,N_23025,N_22298);
xnor UO_2351 (O_2351,N_22811,N_24228);
nand UO_2352 (O_2352,N_23369,N_22823);
and UO_2353 (O_2353,N_23805,N_23970);
or UO_2354 (O_2354,N_24821,N_22322);
nand UO_2355 (O_2355,N_23652,N_22701);
nor UO_2356 (O_2356,N_23327,N_24754);
nor UO_2357 (O_2357,N_22255,N_23949);
and UO_2358 (O_2358,N_23705,N_22997);
xnor UO_2359 (O_2359,N_24555,N_22331);
or UO_2360 (O_2360,N_23415,N_24158);
or UO_2361 (O_2361,N_22405,N_23041);
xor UO_2362 (O_2362,N_22467,N_24041);
nor UO_2363 (O_2363,N_22117,N_24014);
or UO_2364 (O_2364,N_24627,N_22713);
nand UO_2365 (O_2365,N_24534,N_24115);
or UO_2366 (O_2366,N_24045,N_24647);
or UO_2367 (O_2367,N_24597,N_22041);
or UO_2368 (O_2368,N_24851,N_24751);
and UO_2369 (O_2369,N_22505,N_24202);
xor UO_2370 (O_2370,N_22966,N_23049);
and UO_2371 (O_2371,N_22983,N_23930);
and UO_2372 (O_2372,N_23583,N_24571);
or UO_2373 (O_2373,N_23074,N_22038);
nor UO_2374 (O_2374,N_24825,N_24735);
and UO_2375 (O_2375,N_24308,N_24974);
nand UO_2376 (O_2376,N_24474,N_22430);
nand UO_2377 (O_2377,N_22017,N_23222);
or UO_2378 (O_2378,N_24691,N_23901);
xor UO_2379 (O_2379,N_24990,N_24931);
or UO_2380 (O_2380,N_24259,N_23622);
or UO_2381 (O_2381,N_22185,N_23857);
nor UO_2382 (O_2382,N_24364,N_21981);
or UO_2383 (O_2383,N_23914,N_21914);
nand UO_2384 (O_2384,N_23545,N_22501);
or UO_2385 (O_2385,N_23220,N_23223);
xnor UO_2386 (O_2386,N_22562,N_23445);
and UO_2387 (O_2387,N_23588,N_24743);
and UO_2388 (O_2388,N_23892,N_24370);
nor UO_2389 (O_2389,N_22424,N_23086);
nand UO_2390 (O_2390,N_22055,N_24256);
xor UO_2391 (O_2391,N_24278,N_23576);
xor UO_2392 (O_2392,N_23946,N_22564);
and UO_2393 (O_2393,N_24794,N_22971);
nand UO_2394 (O_2394,N_24236,N_23297);
xor UO_2395 (O_2395,N_24175,N_23190);
nand UO_2396 (O_2396,N_24953,N_24643);
nand UO_2397 (O_2397,N_23382,N_22556);
or UO_2398 (O_2398,N_22420,N_22895);
and UO_2399 (O_2399,N_22550,N_24879);
nand UO_2400 (O_2400,N_23550,N_22837);
and UO_2401 (O_2401,N_22504,N_24286);
nand UO_2402 (O_2402,N_23156,N_22534);
or UO_2403 (O_2403,N_23044,N_22996);
or UO_2404 (O_2404,N_23660,N_22793);
or UO_2405 (O_2405,N_24679,N_21890);
or UO_2406 (O_2406,N_22729,N_23934);
nor UO_2407 (O_2407,N_22069,N_23667);
nor UO_2408 (O_2408,N_24479,N_22146);
and UO_2409 (O_2409,N_24982,N_23754);
nor UO_2410 (O_2410,N_23886,N_22563);
nand UO_2411 (O_2411,N_22423,N_24012);
nand UO_2412 (O_2412,N_22710,N_24117);
and UO_2413 (O_2413,N_22631,N_23027);
nor UO_2414 (O_2414,N_21972,N_24457);
and UO_2415 (O_2415,N_22600,N_22606);
and UO_2416 (O_2416,N_24933,N_22820);
and UO_2417 (O_2417,N_22822,N_24329);
and UO_2418 (O_2418,N_24277,N_23027);
xnor UO_2419 (O_2419,N_22727,N_22718);
nor UO_2420 (O_2420,N_24009,N_23522);
nor UO_2421 (O_2421,N_24550,N_22325);
nor UO_2422 (O_2422,N_22443,N_23660);
and UO_2423 (O_2423,N_22394,N_22850);
nor UO_2424 (O_2424,N_23514,N_24804);
nor UO_2425 (O_2425,N_21993,N_24424);
xor UO_2426 (O_2426,N_23106,N_24054);
or UO_2427 (O_2427,N_24149,N_23601);
nor UO_2428 (O_2428,N_23588,N_24873);
or UO_2429 (O_2429,N_24455,N_24304);
and UO_2430 (O_2430,N_24759,N_22050);
nand UO_2431 (O_2431,N_23782,N_23819);
xor UO_2432 (O_2432,N_23180,N_24460);
xor UO_2433 (O_2433,N_23703,N_24628);
nand UO_2434 (O_2434,N_21981,N_24625);
or UO_2435 (O_2435,N_24156,N_24788);
or UO_2436 (O_2436,N_22185,N_24272);
or UO_2437 (O_2437,N_24055,N_21988);
nand UO_2438 (O_2438,N_24713,N_22478);
or UO_2439 (O_2439,N_23972,N_24544);
xnor UO_2440 (O_2440,N_24022,N_22445);
xor UO_2441 (O_2441,N_24000,N_24223);
or UO_2442 (O_2442,N_24071,N_22044);
xor UO_2443 (O_2443,N_21961,N_24007);
nor UO_2444 (O_2444,N_24830,N_24059);
and UO_2445 (O_2445,N_24781,N_22504);
nand UO_2446 (O_2446,N_23525,N_23862);
or UO_2447 (O_2447,N_24620,N_24441);
and UO_2448 (O_2448,N_24472,N_24540);
nor UO_2449 (O_2449,N_22877,N_22285);
and UO_2450 (O_2450,N_24132,N_21948);
and UO_2451 (O_2451,N_22668,N_24324);
xnor UO_2452 (O_2452,N_24986,N_22965);
or UO_2453 (O_2453,N_24655,N_23029);
xnor UO_2454 (O_2454,N_22604,N_24045);
nand UO_2455 (O_2455,N_24023,N_22228);
or UO_2456 (O_2456,N_24713,N_21922);
or UO_2457 (O_2457,N_22777,N_23073);
nor UO_2458 (O_2458,N_22526,N_23901);
nand UO_2459 (O_2459,N_23541,N_22701);
and UO_2460 (O_2460,N_23479,N_24747);
or UO_2461 (O_2461,N_22267,N_24191);
nand UO_2462 (O_2462,N_24101,N_23536);
or UO_2463 (O_2463,N_23409,N_22610);
nor UO_2464 (O_2464,N_22618,N_23231);
xor UO_2465 (O_2465,N_23695,N_24850);
or UO_2466 (O_2466,N_22710,N_24709);
xnor UO_2467 (O_2467,N_24247,N_23257);
nand UO_2468 (O_2468,N_23636,N_23847);
xnor UO_2469 (O_2469,N_22169,N_24366);
nor UO_2470 (O_2470,N_23195,N_23916);
nand UO_2471 (O_2471,N_23391,N_23906);
xnor UO_2472 (O_2472,N_23405,N_23036);
xnor UO_2473 (O_2473,N_21878,N_24105);
or UO_2474 (O_2474,N_24801,N_24011);
or UO_2475 (O_2475,N_22666,N_22574);
xor UO_2476 (O_2476,N_23805,N_24984);
nor UO_2477 (O_2477,N_23585,N_24064);
and UO_2478 (O_2478,N_21960,N_23288);
xor UO_2479 (O_2479,N_23194,N_24155);
and UO_2480 (O_2480,N_23015,N_22709);
xnor UO_2481 (O_2481,N_22415,N_23326);
xnor UO_2482 (O_2482,N_22769,N_22474);
and UO_2483 (O_2483,N_24387,N_23352);
nor UO_2484 (O_2484,N_24077,N_24912);
xnor UO_2485 (O_2485,N_21903,N_24702);
nor UO_2486 (O_2486,N_24727,N_24811);
nand UO_2487 (O_2487,N_24422,N_24836);
xor UO_2488 (O_2488,N_24078,N_22006);
and UO_2489 (O_2489,N_22705,N_23772);
xnor UO_2490 (O_2490,N_21909,N_23899);
nor UO_2491 (O_2491,N_23244,N_22279);
xor UO_2492 (O_2492,N_22016,N_24566);
and UO_2493 (O_2493,N_22735,N_24482);
or UO_2494 (O_2494,N_24574,N_24708);
or UO_2495 (O_2495,N_23812,N_23182);
or UO_2496 (O_2496,N_24364,N_23111);
xnor UO_2497 (O_2497,N_22708,N_22764);
xnor UO_2498 (O_2498,N_23218,N_21942);
nor UO_2499 (O_2499,N_23692,N_23277);
and UO_2500 (O_2500,N_23764,N_23295);
xor UO_2501 (O_2501,N_22865,N_24735);
xnor UO_2502 (O_2502,N_24446,N_21923);
nand UO_2503 (O_2503,N_22148,N_24580);
and UO_2504 (O_2504,N_22113,N_23501);
and UO_2505 (O_2505,N_22929,N_24123);
or UO_2506 (O_2506,N_22000,N_23120);
and UO_2507 (O_2507,N_22550,N_24055);
nor UO_2508 (O_2508,N_24010,N_23438);
nand UO_2509 (O_2509,N_24846,N_22183);
and UO_2510 (O_2510,N_23100,N_22247);
xor UO_2511 (O_2511,N_22800,N_23480);
nor UO_2512 (O_2512,N_23056,N_24432);
and UO_2513 (O_2513,N_22732,N_24457);
and UO_2514 (O_2514,N_23206,N_24448);
xnor UO_2515 (O_2515,N_22173,N_23664);
and UO_2516 (O_2516,N_22177,N_22406);
and UO_2517 (O_2517,N_22361,N_24300);
and UO_2518 (O_2518,N_21906,N_23990);
or UO_2519 (O_2519,N_24127,N_23602);
nand UO_2520 (O_2520,N_22964,N_24685);
nor UO_2521 (O_2521,N_23094,N_23471);
and UO_2522 (O_2522,N_22549,N_24434);
nand UO_2523 (O_2523,N_24609,N_22440);
nor UO_2524 (O_2524,N_22186,N_23796);
xnor UO_2525 (O_2525,N_22663,N_22874);
nand UO_2526 (O_2526,N_22700,N_22235);
nand UO_2527 (O_2527,N_24020,N_24729);
or UO_2528 (O_2528,N_23155,N_24400);
or UO_2529 (O_2529,N_22614,N_22348);
or UO_2530 (O_2530,N_23572,N_24275);
or UO_2531 (O_2531,N_22846,N_22181);
and UO_2532 (O_2532,N_24751,N_23242);
nand UO_2533 (O_2533,N_23375,N_23783);
nor UO_2534 (O_2534,N_22114,N_23618);
or UO_2535 (O_2535,N_23585,N_23080);
xnor UO_2536 (O_2536,N_22043,N_23428);
nor UO_2537 (O_2537,N_23701,N_22905);
xor UO_2538 (O_2538,N_23874,N_23340);
or UO_2539 (O_2539,N_23909,N_21941);
nor UO_2540 (O_2540,N_22321,N_22025);
nand UO_2541 (O_2541,N_23443,N_24187);
or UO_2542 (O_2542,N_23649,N_24301);
xnor UO_2543 (O_2543,N_22044,N_21916);
xor UO_2544 (O_2544,N_24217,N_23255);
xnor UO_2545 (O_2545,N_24292,N_22813);
and UO_2546 (O_2546,N_22975,N_22762);
xor UO_2547 (O_2547,N_24902,N_23482);
xor UO_2548 (O_2548,N_23986,N_24706);
xnor UO_2549 (O_2549,N_23383,N_24788);
xor UO_2550 (O_2550,N_24255,N_24946);
nor UO_2551 (O_2551,N_23282,N_24969);
or UO_2552 (O_2552,N_24400,N_23861);
nand UO_2553 (O_2553,N_22434,N_24377);
nand UO_2554 (O_2554,N_23295,N_23965);
xor UO_2555 (O_2555,N_22745,N_22467);
and UO_2556 (O_2556,N_23935,N_24415);
xnor UO_2557 (O_2557,N_23549,N_23750);
nand UO_2558 (O_2558,N_23037,N_24897);
or UO_2559 (O_2559,N_24467,N_22944);
nand UO_2560 (O_2560,N_22769,N_23092);
and UO_2561 (O_2561,N_22460,N_22238);
xnor UO_2562 (O_2562,N_23300,N_24060);
nand UO_2563 (O_2563,N_22464,N_23797);
and UO_2564 (O_2564,N_22664,N_23262);
and UO_2565 (O_2565,N_23899,N_22532);
nand UO_2566 (O_2566,N_24700,N_24029);
nor UO_2567 (O_2567,N_22817,N_23646);
and UO_2568 (O_2568,N_23102,N_24737);
nor UO_2569 (O_2569,N_21960,N_22577);
and UO_2570 (O_2570,N_24430,N_24738);
and UO_2571 (O_2571,N_22953,N_22805);
and UO_2572 (O_2572,N_24299,N_24014);
xor UO_2573 (O_2573,N_22855,N_23347);
xor UO_2574 (O_2574,N_23384,N_23293);
xor UO_2575 (O_2575,N_24588,N_23971);
and UO_2576 (O_2576,N_24170,N_22139);
nor UO_2577 (O_2577,N_23974,N_23893);
or UO_2578 (O_2578,N_23675,N_23580);
nand UO_2579 (O_2579,N_24194,N_24905);
and UO_2580 (O_2580,N_22834,N_24586);
or UO_2581 (O_2581,N_22595,N_23525);
nand UO_2582 (O_2582,N_23557,N_22978);
xor UO_2583 (O_2583,N_22061,N_23622);
nand UO_2584 (O_2584,N_24559,N_23316);
or UO_2585 (O_2585,N_23806,N_23066);
nor UO_2586 (O_2586,N_23813,N_24994);
xnor UO_2587 (O_2587,N_24239,N_24694);
or UO_2588 (O_2588,N_23725,N_23295);
nor UO_2589 (O_2589,N_22663,N_24580);
or UO_2590 (O_2590,N_24943,N_22031);
or UO_2591 (O_2591,N_22643,N_24539);
nand UO_2592 (O_2592,N_23326,N_22826);
xnor UO_2593 (O_2593,N_23585,N_24994);
and UO_2594 (O_2594,N_23912,N_22680);
nand UO_2595 (O_2595,N_22036,N_22653);
or UO_2596 (O_2596,N_22126,N_24363);
xor UO_2597 (O_2597,N_22124,N_21954);
nand UO_2598 (O_2598,N_24932,N_23233);
nand UO_2599 (O_2599,N_23878,N_22343);
or UO_2600 (O_2600,N_23712,N_23056);
nor UO_2601 (O_2601,N_24331,N_24861);
xnor UO_2602 (O_2602,N_24535,N_24466);
and UO_2603 (O_2603,N_23977,N_23290);
nor UO_2604 (O_2604,N_22858,N_24167);
or UO_2605 (O_2605,N_21930,N_24949);
and UO_2606 (O_2606,N_23956,N_23667);
or UO_2607 (O_2607,N_23671,N_21938);
and UO_2608 (O_2608,N_22768,N_23169);
nor UO_2609 (O_2609,N_21950,N_24117);
and UO_2610 (O_2610,N_22453,N_23933);
nor UO_2611 (O_2611,N_24769,N_23794);
xor UO_2612 (O_2612,N_23519,N_24858);
xor UO_2613 (O_2613,N_21978,N_24580);
or UO_2614 (O_2614,N_23309,N_23968);
xor UO_2615 (O_2615,N_21956,N_24195);
xnor UO_2616 (O_2616,N_22540,N_23299);
nor UO_2617 (O_2617,N_23654,N_22851);
or UO_2618 (O_2618,N_22276,N_21876);
and UO_2619 (O_2619,N_24102,N_24407);
nor UO_2620 (O_2620,N_22297,N_23215);
nor UO_2621 (O_2621,N_23135,N_24185);
or UO_2622 (O_2622,N_24562,N_24580);
nor UO_2623 (O_2623,N_22911,N_24416);
and UO_2624 (O_2624,N_23953,N_23175);
and UO_2625 (O_2625,N_23972,N_24099);
and UO_2626 (O_2626,N_22828,N_22765);
and UO_2627 (O_2627,N_23841,N_22036);
or UO_2628 (O_2628,N_23105,N_23923);
xnor UO_2629 (O_2629,N_22820,N_22198);
xor UO_2630 (O_2630,N_24748,N_23645);
and UO_2631 (O_2631,N_23319,N_22836);
or UO_2632 (O_2632,N_23085,N_22521);
xnor UO_2633 (O_2633,N_22590,N_23445);
nand UO_2634 (O_2634,N_24544,N_24198);
nor UO_2635 (O_2635,N_23381,N_22878);
and UO_2636 (O_2636,N_24426,N_23942);
nor UO_2637 (O_2637,N_23719,N_23506);
nand UO_2638 (O_2638,N_24964,N_23517);
nor UO_2639 (O_2639,N_24781,N_24952);
or UO_2640 (O_2640,N_23926,N_24309);
or UO_2641 (O_2641,N_24221,N_23004);
and UO_2642 (O_2642,N_23154,N_24317);
xor UO_2643 (O_2643,N_22552,N_24759);
or UO_2644 (O_2644,N_23383,N_23296);
xnor UO_2645 (O_2645,N_24467,N_23821);
nand UO_2646 (O_2646,N_23199,N_24171);
or UO_2647 (O_2647,N_24098,N_21991);
or UO_2648 (O_2648,N_22289,N_22294);
xnor UO_2649 (O_2649,N_23990,N_24910);
nor UO_2650 (O_2650,N_23938,N_21913);
and UO_2651 (O_2651,N_23561,N_22375);
or UO_2652 (O_2652,N_22737,N_22861);
or UO_2653 (O_2653,N_23622,N_23111);
xnor UO_2654 (O_2654,N_23438,N_21956);
nand UO_2655 (O_2655,N_24797,N_24891);
and UO_2656 (O_2656,N_23905,N_23707);
nor UO_2657 (O_2657,N_24619,N_24391);
nand UO_2658 (O_2658,N_22936,N_23039);
and UO_2659 (O_2659,N_23598,N_24979);
nor UO_2660 (O_2660,N_23312,N_24581);
xnor UO_2661 (O_2661,N_24395,N_24783);
or UO_2662 (O_2662,N_24382,N_23117);
nand UO_2663 (O_2663,N_22576,N_22407);
nor UO_2664 (O_2664,N_24111,N_23560);
nand UO_2665 (O_2665,N_24776,N_23621);
and UO_2666 (O_2666,N_22778,N_24001);
nor UO_2667 (O_2667,N_23641,N_23740);
or UO_2668 (O_2668,N_24283,N_22613);
nand UO_2669 (O_2669,N_22653,N_22069);
nand UO_2670 (O_2670,N_22741,N_24016);
and UO_2671 (O_2671,N_24942,N_22850);
nand UO_2672 (O_2672,N_22824,N_23830);
xnor UO_2673 (O_2673,N_24159,N_22764);
xor UO_2674 (O_2674,N_22314,N_24692);
xnor UO_2675 (O_2675,N_23877,N_24164);
xnor UO_2676 (O_2676,N_21880,N_22766);
nor UO_2677 (O_2677,N_22115,N_24699);
xnor UO_2678 (O_2678,N_23895,N_24558);
and UO_2679 (O_2679,N_23465,N_22385);
xor UO_2680 (O_2680,N_23287,N_24679);
or UO_2681 (O_2681,N_24279,N_24528);
xnor UO_2682 (O_2682,N_24256,N_24347);
nand UO_2683 (O_2683,N_23235,N_22970);
xnor UO_2684 (O_2684,N_23687,N_23690);
nor UO_2685 (O_2685,N_22971,N_23448);
xnor UO_2686 (O_2686,N_22457,N_22419);
nand UO_2687 (O_2687,N_23497,N_22908);
xor UO_2688 (O_2688,N_24960,N_23635);
nor UO_2689 (O_2689,N_23292,N_24483);
nand UO_2690 (O_2690,N_22014,N_23911);
and UO_2691 (O_2691,N_24250,N_22228);
xor UO_2692 (O_2692,N_24230,N_24711);
or UO_2693 (O_2693,N_23790,N_24631);
and UO_2694 (O_2694,N_22892,N_24123);
nand UO_2695 (O_2695,N_22899,N_24462);
or UO_2696 (O_2696,N_22439,N_24074);
nand UO_2697 (O_2697,N_24425,N_24496);
and UO_2698 (O_2698,N_24028,N_21965);
nand UO_2699 (O_2699,N_23213,N_24564);
or UO_2700 (O_2700,N_23507,N_24685);
nand UO_2701 (O_2701,N_22026,N_23151);
xor UO_2702 (O_2702,N_24311,N_24628);
or UO_2703 (O_2703,N_23614,N_23272);
and UO_2704 (O_2704,N_22011,N_24971);
nand UO_2705 (O_2705,N_23103,N_24076);
xor UO_2706 (O_2706,N_22656,N_22013);
xnor UO_2707 (O_2707,N_22312,N_22714);
nand UO_2708 (O_2708,N_22075,N_23271);
xor UO_2709 (O_2709,N_23559,N_23821);
or UO_2710 (O_2710,N_24966,N_22979);
xor UO_2711 (O_2711,N_22106,N_22595);
and UO_2712 (O_2712,N_23818,N_22200);
or UO_2713 (O_2713,N_24026,N_23683);
nand UO_2714 (O_2714,N_23734,N_24549);
and UO_2715 (O_2715,N_21934,N_22745);
nor UO_2716 (O_2716,N_22609,N_23434);
nor UO_2717 (O_2717,N_22465,N_23859);
nand UO_2718 (O_2718,N_24268,N_24756);
nand UO_2719 (O_2719,N_24498,N_23770);
xor UO_2720 (O_2720,N_24892,N_22748);
and UO_2721 (O_2721,N_24678,N_24401);
nand UO_2722 (O_2722,N_24929,N_22221);
nor UO_2723 (O_2723,N_23967,N_22635);
xnor UO_2724 (O_2724,N_23138,N_23194);
or UO_2725 (O_2725,N_24132,N_23681);
and UO_2726 (O_2726,N_22880,N_23504);
and UO_2727 (O_2727,N_22268,N_21933);
xnor UO_2728 (O_2728,N_22420,N_22344);
nor UO_2729 (O_2729,N_22540,N_23974);
or UO_2730 (O_2730,N_24055,N_23594);
nor UO_2731 (O_2731,N_23193,N_22427);
or UO_2732 (O_2732,N_21995,N_24328);
xnor UO_2733 (O_2733,N_24680,N_22701);
xnor UO_2734 (O_2734,N_21913,N_23890);
or UO_2735 (O_2735,N_22889,N_22138);
and UO_2736 (O_2736,N_23971,N_23353);
nand UO_2737 (O_2737,N_24684,N_24259);
nor UO_2738 (O_2738,N_22580,N_22875);
nor UO_2739 (O_2739,N_24253,N_23344);
nand UO_2740 (O_2740,N_22490,N_24284);
or UO_2741 (O_2741,N_24275,N_24720);
nor UO_2742 (O_2742,N_24761,N_22056);
xnor UO_2743 (O_2743,N_22841,N_24479);
nand UO_2744 (O_2744,N_22251,N_23918);
and UO_2745 (O_2745,N_21894,N_23190);
nor UO_2746 (O_2746,N_24804,N_24829);
nor UO_2747 (O_2747,N_22883,N_24762);
or UO_2748 (O_2748,N_24765,N_23807);
nor UO_2749 (O_2749,N_24183,N_24534);
nor UO_2750 (O_2750,N_24764,N_22232);
nor UO_2751 (O_2751,N_23186,N_24064);
or UO_2752 (O_2752,N_23929,N_24422);
nor UO_2753 (O_2753,N_24451,N_22057);
nand UO_2754 (O_2754,N_23133,N_24033);
xnor UO_2755 (O_2755,N_24771,N_22367);
or UO_2756 (O_2756,N_24885,N_24365);
nor UO_2757 (O_2757,N_24184,N_23205);
nor UO_2758 (O_2758,N_24615,N_21999);
or UO_2759 (O_2759,N_23961,N_23235);
and UO_2760 (O_2760,N_22918,N_22653);
nor UO_2761 (O_2761,N_24540,N_22975);
xor UO_2762 (O_2762,N_24893,N_24243);
nor UO_2763 (O_2763,N_23582,N_22407);
xor UO_2764 (O_2764,N_22339,N_24191);
nand UO_2765 (O_2765,N_24471,N_24846);
and UO_2766 (O_2766,N_23499,N_24064);
nor UO_2767 (O_2767,N_23336,N_22799);
or UO_2768 (O_2768,N_24175,N_23973);
nand UO_2769 (O_2769,N_23347,N_22429);
or UO_2770 (O_2770,N_23752,N_22007);
nor UO_2771 (O_2771,N_23777,N_23850);
xor UO_2772 (O_2772,N_22052,N_22123);
and UO_2773 (O_2773,N_22347,N_23443);
xor UO_2774 (O_2774,N_23224,N_24124);
nor UO_2775 (O_2775,N_21970,N_23497);
xor UO_2776 (O_2776,N_24469,N_23586);
nor UO_2777 (O_2777,N_23796,N_22855);
or UO_2778 (O_2778,N_24301,N_24439);
and UO_2779 (O_2779,N_22977,N_23186);
nor UO_2780 (O_2780,N_22953,N_23122);
or UO_2781 (O_2781,N_22322,N_24188);
and UO_2782 (O_2782,N_23976,N_24115);
nand UO_2783 (O_2783,N_24955,N_24682);
nor UO_2784 (O_2784,N_22868,N_24526);
nor UO_2785 (O_2785,N_23129,N_23145);
or UO_2786 (O_2786,N_23547,N_22009);
nand UO_2787 (O_2787,N_23642,N_24991);
nand UO_2788 (O_2788,N_22568,N_23044);
or UO_2789 (O_2789,N_24292,N_24833);
or UO_2790 (O_2790,N_24828,N_22242);
and UO_2791 (O_2791,N_22978,N_24857);
or UO_2792 (O_2792,N_23506,N_22150);
and UO_2793 (O_2793,N_23627,N_24203);
nand UO_2794 (O_2794,N_21951,N_23173);
or UO_2795 (O_2795,N_22521,N_23211);
and UO_2796 (O_2796,N_23074,N_22392);
and UO_2797 (O_2797,N_22312,N_22056);
or UO_2798 (O_2798,N_22469,N_22709);
and UO_2799 (O_2799,N_24025,N_24417);
or UO_2800 (O_2800,N_23867,N_23554);
or UO_2801 (O_2801,N_23150,N_21904);
or UO_2802 (O_2802,N_23945,N_24367);
xnor UO_2803 (O_2803,N_22485,N_23746);
nor UO_2804 (O_2804,N_22515,N_23561);
xor UO_2805 (O_2805,N_23888,N_22215);
nor UO_2806 (O_2806,N_24409,N_24512);
nor UO_2807 (O_2807,N_23554,N_22793);
and UO_2808 (O_2808,N_24917,N_24674);
or UO_2809 (O_2809,N_24951,N_24937);
and UO_2810 (O_2810,N_23456,N_21997);
and UO_2811 (O_2811,N_24260,N_24912);
or UO_2812 (O_2812,N_23592,N_24875);
nor UO_2813 (O_2813,N_23898,N_22627);
nor UO_2814 (O_2814,N_22755,N_23313);
or UO_2815 (O_2815,N_23270,N_24284);
or UO_2816 (O_2816,N_24351,N_22275);
or UO_2817 (O_2817,N_22805,N_23635);
xor UO_2818 (O_2818,N_22574,N_24949);
xnor UO_2819 (O_2819,N_22831,N_22233);
nor UO_2820 (O_2820,N_23554,N_24796);
xor UO_2821 (O_2821,N_22464,N_24835);
nand UO_2822 (O_2822,N_22352,N_23790);
and UO_2823 (O_2823,N_24872,N_24192);
and UO_2824 (O_2824,N_23824,N_23591);
nor UO_2825 (O_2825,N_24579,N_24588);
xor UO_2826 (O_2826,N_22024,N_22399);
nand UO_2827 (O_2827,N_23348,N_22480);
xnor UO_2828 (O_2828,N_22237,N_22608);
xor UO_2829 (O_2829,N_23706,N_22089);
nand UO_2830 (O_2830,N_22271,N_23481);
nand UO_2831 (O_2831,N_23282,N_23360);
xnor UO_2832 (O_2832,N_24357,N_24100);
nor UO_2833 (O_2833,N_23037,N_22771);
or UO_2834 (O_2834,N_22039,N_22411);
nor UO_2835 (O_2835,N_22177,N_24456);
and UO_2836 (O_2836,N_23271,N_24892);
nor UO_2837 (O_2837,N_22343,N_21971);
or UO_2838 (O_2838,N_22430,N_21878);
xnor UO_2839 (O_2839,N_23648,N_23500);
nand UO_2840 (O_2840,N_23224,N_24085);
nand UO_2841 (O_2841,N_24433,N_23855);
and UO_2842 (O_2842,N_24930,N_23347);
xnor UO_2843 (O_2843,N_24393,N_22267);
nor UO_2844 (O_2844,N_22939,N_22846);
xnor UO_2845 (O_2845,N_24678,N_22610);
or UO_2846 (O_2846,N_21927,N_24159);
nor UO_2847 (O_2847,N_21876,N_23729);
nor UO_2848 (O_2848,N_22522,N_22893);
or UO_2849 (O_2849,N_23249,N_21985);
nor UO_2850 (O_2850,N_23358,N_24329);
nand UO_2851 (O_2851,N_24380,N_22509);
or UO_2852 (O_2852,N_22520,N_23770);
or UO_2853 (O_2853,N_23233,N_22940);
xor UO_2854 (O_2854,N_21929,N_24793);
or UO_2855 (O_2855,N_22571,N_22951);
or UO_2856 (O_2856,N_23010,N_22546);
xor UO_2857 (O_2857,N_23159,N_22421);
nand UO_2858 (O_2858,N_23534,N_23614);
or UO_2859 (O_2859,N_23860,N_23106);
nand UO_2860 (O_2860,N_23942,N_24413);
xor UO_2861 (O_2861,N_21924,N_22500);
nor UO_2862 (O_2862,N_24163,N_23413);
and UO_2863 (O_2863,N_24625,N_24529);
or UO_2864 (O_2864,N_23191,N_23026);
and UO_2865 (O_2865,N_23002,N_24970);
nand UO_2866 (O_2866,N_23983,N_22794);
and UO_2867 (O_2867,N_22743,N_23025);
nand UO_2868 (O_2868,N_23503,N_24756);
xnor UO_2869 (O_2869,N_24364,N_23919);
nand UO_2870 (O_2870,N_22982,N_24894);
or UO_2871 (O_2871,N_22462,N_23782);
xnor UO_2872 (O_2872,N_22878,N_23196);
nand UO_2873 (O_2873,N_24018,N_22610);
and UO_2874 (O_2874,N_22126,N_23954);
xor UO_2875 (O_2875,N_22887,N_22211);
and UO_2876 (O_2876,N_24447,N_23095);
nor UO_2877 (O_2877,N_23776,N_23975);
xor UO_2878 (O_2878,N_23772,N_24302);
or UO_2879 (O_2879,N_22663,N_22070);
xor UO_2880 (O_2880,N_24549,N_23455);
nand UO_2881 (O_2881,N_22257,N_22137);
nand UO_2882 (O_2882,N_24959,N_22951);
nand UO_2883 (O_2883,N_23593,N_24905);
nand UO_2884 (O_2884,N_23911,N_24806);
xor UO_2885 (O_2885,N_22545,N_21994);
nor UO_2886 (O_2886,N_22984,N_23958);
or UO_2887 (O_2887,N_22308,N_24033);
and UO_2888 (O_2888,N_24780,N_24624);
nand UO_2889 (O_2889,N_24274,N_22736);
xor UO_2890 (O_2890,N_23581,N_22420);
xnor UO_2891 (O_2891,N_23171,N_23690);
nand UO_2892 (O_2892,N_24803,N_23960);
xnor UO_2893 (O_2893,N_24525,N_24743);
xnor UO_2894 (O_2894,N_23585,N_23051);
or UO_2895 (O_2895,N_21986,N_24636);
or UO_2896 (O_2896,N_23782,N_23432);
nand UO_2897 (O_2897,N_23243,N_22006);
nand UO_2898 (O_2898,N_22884,N_23700);
nand UO_2899 (O_2899,N_22368,N_24872);
nand UO_2900 (O_2900,N_22201,N_22558);
nor UO_2901 (O_2901,N_23664,N_24295);
and UO_2902 (O_2902,N_22608,N_23443);
or UO_2903 (O_2903,N_21914,N_23666);
or UO_2904 (O_2904,N_23833,N_23399);
and UO_2905 (O_2905,N_22407,N_22393);
and UO_2906 (O_2906,N_23267,N_22650);
xnor UO_2907 (O_2907,N_23235,N_23675);
and UO_2908 (O_2908,N_24781,N_24602);
xor UO_2909 (O_2909,N_23350,N_22544);
nand UO_2910 (O_2910,N_22095,N_24076);
nor UO_2911 (O_2911,N_24266,N_23684);
and UO_2912 (O_2912,N_22601,N_22045);
xor UO_2913 (O_2913,N_22763,N_24463);
or UO_2914 (O_2914,N_23886,N_24090);
nor UO_2915 (O_2915,N_24996,N_22793);
nand UO_2916 (O_2916,N_22249,N_23925);
and UO_2917 (O_2917,N_22479,N_22206);
xnor UO_2918 (O_2918,N_22194,N_24373);
xnor UO_2919 (O_2919,N_23689,N_24381);
nand UO_2920 (O_2920,N_22627,N_22012);
nand UO_2921 (O_2921,N_24212,N_22710);
or UO_2922 (O_2922,N_22029,N_22290);
nor UO_2923 (O_2923,N_24061,N_24663);
xnor UO_2924 (O_2924,N_22571,N_24713);
xnor UO_2925 (O_2925,N_23552,N_24370);
or UO_2926 (O_2926,N_21923,N_23163);
xor UO_2927 (O_2927,N_22332,N_24899);
and UO_2928 (O_2928,N_22176,N_22759);
xnor UO_2929 (O_2929,N_24701,N_23293);
and UO_2930 (O_2930,N_23823,N_24995);
and UO_2931 (O_2931,N_21897,N_21913);
nand UO_2932 (O_2932,N_22744,N_22276);
xnor UO_2933 (O_2933,N_24346,N_23037);
or UO_2934 (O_2934,N_24132,N_21983);
or UO_2935 (O_2935,N_23638,N_24995);
or UO_2936 (O_2936,N_23905,N_23445);
nor UO_2937 (O_2937,N_24220,N_23562);
or UO_2938 (O_2938,N_23419,N_22819);
or UO_2939 (O_2939,N_24511,N_24757);
or UO_2940 (O_2940,N_24836,N_22993);
xnor UO_2941 (O_2941,N_23801,N_21905);
xor UO_2942 (O_2942,N_24726,N_23204);
and UO_2943 (O_2943,N_24041,N_22743);
nor UO_2944 (O_2944,N_24484,N_22985);
nor UO_2945 (O_2945,N_24454,N_22131);
nor UO_2946 (O_2946,N_22066,N_23284);
and UO_2947 (O_2947,N_23062,N_22860);
and UO_2948 (O_2948,N_22575,N_22637);
or UO_2949 (O_2949,N_22120,N_23169);
and UO_2950 (O_2950,N_22287,N_24938);
nor UO_2951 (O_2951,N_23439,N_23753);
nand UO_2952 (O_2952,N_22509,N_24262);
xnor UO_2953 (O_2953,N_22678,N_22024);
nor UO_2954 (O_2954,N_23089,N_24350);
nor UO_2955 (O_2955,N_23597,N_24850);
or UO_2956 (O_2956,N_22316,N_23036);
nor UO_2957 (O_2957,N_24278,N_22319);
nor UO_2958 (O_2958,N_22093,N_24934);
nand UO_2959 (O_2959,N_23741,N_22012);
xnor UO_2960 (O_2960,N_23041,N_24456);
nand UO_2961 (O_2961,N_24935,N_24408);
and UO_2962 (O_2962,N_24917,N_23302);
nor UO_2963 (O_2963,N_23270,N_24647);
or UO_2964 (O_2964,N_22159,N_24104);
or UO_2965 (O_2965,N_24879,N_23400);
or UO_2966 (O_2966,N_23155,N_24145);
xnor UO_2967 (O_2967,N_23272,N_22667);
nor UO_2968 (O_2968,N_24744,N_24155);
nand UO_2969 (O_2969,N_23145,N_22112);
xor UO_2970 (O_2970,N_23431,N_22180);
nand UO_2971 (O_2971,N_24441,N_24516);
or UO_2972 (O_2972,N_24583,N_23923);
or UO_2973 (O_2973,N_24790,N_23162);
nand UO_2974 (O_2974,N_23778,N_24884);
xnor UO_2975 (O_2975,N_24136,N_24117);
nor UO_2976 (O_2976,N_24456,N_24914);
and UO_2977 (O_2977,N_22056,N_24472);
nor UO_2978 (O_2978,N_22686,N_22705);
nand UO_2979 (O_2979,N_24689,N_22571);
nand UO_2980 (O_2980,N_23798,N_24523);
or UO_2981 (O_2981,N_24219,N_23006);
or UO_2982 (O_2982,N_23648,N_24493);
nor UO_2983 (O_2983,N_24880,N_21962);
or UO_2984 (O_2984,N_23638,N_23917);
or UO_2985 (O_2985,N_22885,N_22025);
nor UO_2986 (O_2986,N_23307,N_22305);
xnor UO_2987 (O_2987,N_22571,N_24617);
and UO_2988 (O_2988,N_23195,N_22391);
or UO_2989 (O_2989,N_23712,N_22317);
and UO_2990 (O_2990,N_24689,N_22618);
or UO_2991 (O_2991,N_22286,N_22166);
and UO_2992 (O_2992,N_23072,N_23817);
xor UO_2993 (O_2993,N_22072,N_24929);
nor UO_2994 (O_2994,N_23538,N_22688);
xor UO_2995 (O_2995,N_23674,N_24023);
nor UO_2996 (O_2996,N_24044,N_22450);
and UO_2997 (O_2997,N_23320,N_23659);
nor UO_2998 (O_2998,N_23123,N_24203);
or UO_2999 (O_2999,N_22713,N_24161);
endmodule