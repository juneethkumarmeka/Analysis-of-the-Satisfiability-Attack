module basic_2000_20000_2500_40_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nor U0 (N_0,In_999,In_745);
and U1 (N_1,In_210,In_1352);
or U2 (N_2,In_326,In_1627);
nand U3 (N_3,In_1771,In_311);
nand U4 (N_4,In_297,In_212);
or U5 (N_5,In_353,In_338);
nor U6 (N_6,In_1468,In_215);
nand U7 (N_7,In_77,In_1952);
or U8 (N_8,In_114,In_1529);
nand U9 (N_9,In_273,In_1014);
or U10 (N_10,In_1870,In_1991);
or U11 (N_11,In_381,In_1411);
and U12 (N_12,In_1886,In_61);
or U13 (N_13,In_719,In_1437);
or U14 (N_14,In_433,In_705);
and U15 (N_15,In_1406,In_594);
or U16 (N_16,In_328,In_55);
and U17 (N_17,In_530,In_31);
nand U18 (N_18,In_1005,In_1148);
nor U19 (N_19,In_1994,In_1665);
or U20 (N_20,In_1710,In_331);
or U21 (N_21,In_1938,In_93);
or U22 (N_22,In_111,In_1085);
and U23 (N_23,In_711,In_395);
or U24 (N_24,In_1976,In_1067);
and U25 (N_25,In_193,In_1155);
or U26 (N_26,In_242,In_978);
or U27 (N_27,In_1922,In_302);
xor U28 (N_28,In_109,In_888);
or U29 (N_29,In_583,In_942);
and U30 (N_30,In_1013,In_1720);
or U31 (N_31,In_169,In_883);
or U32 (N_32,In_1091,In_305);
or U33 (N_33,In_57,In_1499);
and U34 (N_34,In_890,In_1254);
nor U35 (N_35,In_576,In_1302);
nand U36 (N_36,In_313,In_68);
nand U37 (N_37,In_1220,In_646);
xor U38 (N_38,In_1989,In_1859);
nor U39 (N_39,In_1436,In_1258);
or U40 (N_40,In_1951,In_1193);
xnor U41 (N_41,In_1472,In_157);
nand U42 (N_42,In_943,In_1312);
nor U43 (N_43,In_799,In_1253);
or U44 (N_44,In_622,In_1849);
nand U45 (N_45,In_636,In_416);
and U46 (N_46,In_428,In_334);
nand U47 (N_47,In_1142,In_1611);
or U48 (N_48,In_534,In_391);
or U49 (N_49,In_1019,In_285);
nor U50 (N_50,In_22,In_648);
nand U51 (N_51,In_1684,In_1761);
or U52 (N_52,In_269,In_1425);
xnor U53 (N_53,In_1433,In_1049);
or U54 (N_54,In_213,In_1281);
xor U55 (N_55,In_744,In_436);
and U56 (N_56,In_1794,In_1896);
or U57 (N_57,In_753,In_1390);
xor U58 (N_58,In_29,In_1486);
or U59 (N_59,In_1179,In_791);
xor U60 (N_60,In_587,In_610);
and U61 (N_61,In_1104,In_1857);
nand U62 (N_62,In_7,In_1249);
nand U63 (N_63,In_1519,In_941);
xor U64 (N_64,In_256,In_1512);
or U65 (N_65,In_567,In_532);
nor U66 (N_66,In_503,In_776);
and U67 (N_67,In_1518,In_1757);
and U68 (N_68,In_1060,In_642);
nand U69 (N_69,In_663,In_143);
or U70 (N_70,In_489,In_1292);
and U71 (N_71,In_1063,In_232);
nor U72 (N_72,In_480,In_1548);
or U73 (N_73,In_747,In_1537);
nor U74 (N_74,In_1076,In_312);
nand U75 (N_75,In_987,In_358);
or U76 (N_76,In_1335,In_1834);
or U77 (N_77,In_1784,In_886);
nor U78 (N_78,In_1031,In_687);
nor U79 (N_79,In_240,In_807);
nand U80 (N_80,In_1588,In_1133);
or U81 (N_81,In_588,In_18);
or U82 (N_82,In_1051,In_97);
or U83 (N_83,In_380,In_1327);
nor U84 (N_84,In_1651,In_1039);
nor U85 (N_85,In_184,In_134);
and U86 (N_86,In_1349,In_118);
nor U87 (N_87,In_1556,In_1384);
nand U88 (N_88,In_609,In_786);
nand U89 (N_89,In_1464,In_1850);
nand U90 (N_90,In_1586,In_488);
and U91 (N_91,In_1610,In_1978);
or U92 (N_92,In_1541,In_1678);
nand U93 (N_93,In_1137,In_102);
or U94 (N_94,In_595,In_1491);
nor U95 (N_95,In_303,In_1904);
or U96 (N_96,In_1176,In_562);
or U97 (N_97,In_1059,In_1191);
nor U98 (N_98,In_710,In_557);
nor U99 (N_99,In_479,In_1073);
xnor U100 (N_100,In_1631,In_657);
nor U101 (N_101,In_1832,In_292);
xnor U102 (N_102,In_348,In_891);
and U103 (N_103,In_905,In_91);
nand U104 (N_104,In_1008,In_1355);
nand U105 (N_105,In_1341,In_1791);
xor U106 (N_106,In_1926,In_493);
nand U107 (N_107,In_1385,In_201);
or U108 (N_108,In_52,In_1065);
nor U109 (N_109,In_108,In_1027);
xor U110 (N_110,In_1102,In_1205);
nand U111 (N_111,In_956,In_1135);
or U112 (N_112,In_1876,In_995);
or U113 (N_113,In_1743,In_1942);
and U114 (N_114,In_33,In_345);
nand U115 (N_115,In_569,In_1026);
and U116 (N_116,In_757,In_873);
xor U117 (N_117,In_1525,In_241);
nor U118 (N_118,In_607,In_767);
and U119 (N_119,In_1195,In_1925);
nor U120 (N_120,In_695,In_1147);
nor U121 (N_121,In_87,In_1021);
and U122 (N_122,In_1774,In_1868);
and U123 (N_123,In_1821,In_809);
and U124 (N_124,In_1666,In_1600);
nor U125 (N_125,In_621,In_803);
nand U126 (N_126,In_746,In_676);
and U127 (N_127,In_680,In_1100);
nand U128 (N_128,In_270,In_290);
or U129 (N_129,In_1323,In_863);
xor U130 (N_130,In_589,In_1722);
or U131 (N_131,In_396,In_885);
nor U132 (N_132,In_1015,In_815);
or U133 (N_133,In_237,In_92);
and U134 (N_134,In_829,In_579);
nor U135 (N_135,In_546,In_1538);
nor U136 (N_136,In_1508,In_1326);
xnor U137 (N_137,In_133,In_1792);
xor U138 (N_138,In_495,In_889);
nand U139 (N_139,In_1605,In_1316);
and U140 (N_140,In_484,In_414);
or U141 (N_141,In_1576,In_513);
or U142 (N_142,In_160,In_743);
nand U143 (N_143,In_1427,In_505);
xor U144 (N_144,In_1010,In_1636);
nand U145 (N_145,In_1511,In_1682);
nand U146 (N_146,In_1816,In_1558);
xnor U147 (N_147,In_497,In_83);
and U148 (N_148,In_1351,In_1932);
nand U149 (N_149,In_633,In_1136);
xnor U150 (N_150,In_1036,In_1339);
xnor U151 (N_151,In_1933,In_1533);
nand U152 (N_152,In_25,In_526);
or U153 (N_153,In_1712,In_1776);
nor U154 (N_154,In_81,In_1278);
and U155 (N_155,In_1843,In_606);
or U156 (N_156,In_1409,In_1838);
nor U157 (N_157,In_822,In_1668);
nor U158 (N_158,In_765,In_867);
xor U159 (N_159,In_1671,In_795);
nand U160 (N_160,In_1413,In_1293);
xnor U161 (N_161,In_1649,In_1095);
and U162 (N_162,In_1345,In_704);
xnor U163 (N_163,In_1828,In_1052);
nor U164 (N_164,In_485,In_733);
or U165 (N_165,In_1419,In_1023);
xor U166 (N_166,In_289,In_1082);
nor U167 (N_167,In_191,In_1454);
and U168 (N_168,In_1704,In_355);
nand U169 (N_169,In_39,In_1184);
nor U170 (N_170,In_399,In_821);
nor U171 (N_171,In_1983,In_792);
xor U172 (N_172,In_1729,In_690);
nand U173 (N_173,In_228,In_573);
or U174 (N_174,In_700,In_1679);
xor U175 (N_175,In_1673,In_117);
nor U176 (N_176,In_1563,In_1961);
nand U177 (N_177,In_1721,In_1144);
nand U178 (N_178,In_234,In_1730);
nand U179 (N_179,In_903,In_946);
or U180 (N_180,In_628,In_726);
xor U181 (N_181,In_1998,In_100);
nor U182 (N_182,In_1751,In_1368);
nor U183 (N_183,In_418,In_623);
nand U184 (N_184,In_349,In_625);
or U185 (N_185,In_1196,In_1947);
xnor U186 (N_186,In_833,In_1417);
or U187 (N_187,In_644,In_1084);
xor U188 (N_188,In_1950,In_1192);
nand U189 (N_189,In_1889,In_1837);
nand U190 (N_190,In_914,In_73);
nand U191 (N_191,In_2,In_1306);
nor U192 (N_192,In_763,In_1820);
or U193 (N_193,In_1798,In_1484);
or U194 (N_194,In_383,In_1995);
or U195 (N_195,In_63,In_1696);
or U196 (N_196,In_80,In_1362);
xnor U197 (N_197,In_1676,In_1455);
or U198 (N_198,In_110,In_1582);
nor U199 (N_199,In_174,In_1140);
nor U200 (N_200,In_966,In_820);
or U201 (N_201,In_1697,In_85);
or U202 (N_202,In_239,In_1752);
and U203 (N_203,In_1270,In_547);
or U204 (N_204,In_1641,In_286);
nor U205 (N_205,In_1002,In_1210);
nand U206 (N_206,In_518,In_857);
nand U207 (N_207,In_1364,In_1233);
nand U208 (N_208,In_361,In_148);
nand U209 (N_209,In_1325,In_1766);
and U210 (N_210,In_564,In_163);
nor U211 (N_211,In_1806,In_951);
xor U212 (N_212,In_948,In_709);
and U213 (N_213,In_751,In_1962);
nor U214 (N_214,In_550,In_1045);
xnor U215 (N_215,In_870,In_1132);
and U216 (N_216,In_1595,In_510);
nand U217 (N_217,In_132,In_1120);
xnor U218 (N_218,In_459,In_40);
or U219 (N_219,In_1447,In_1106);
nor U220 (N_220,In_1307,In_360);
and U221 (N_221,In_684,In_1158);
nand U222 (N_222,In_811,In_1382);
or U223 (N_223,In_973,In_929);
nor U224 (N_224,In_1506,In_899);
and U225 (N_225,In_202,In_1955);
nand U226 (N_226,In_1880,In_861);
nand U227 (N_227,In_1492,In_260);
and U228 (N_228,In_991,In_1501);
and U229 (N_229,In_46,In_912);
or U230 (N_230,In_1675,In_171);
xnor U231 (N_231,In_137,In_410);
and U232 (N_232,In_1072,In_1157);
nand U233 (N_233,In_136,In_363);
and U234 (N_234,In_385,In_483);
nor U235 (N_235,In_1815,In_1161);
xnor U236 (N_236,In_1892,In_961);
nor U237 (N_237,In_298,In_263);
nand U238 (N_238,In_10,In_1698);
nand U239 (N_239,In_1423,In_618);
or U240 (N_240,In_1319,In_1357);
nor U241 (N_241,In_571,In_968);
nand U242 (N_242,In_1213,In_1907);
nor U243 (N_243,In_1753,In_643);
nor U244 (N_244,In_1295,In_1913);
nor U245 (N_245,In_1905,In_565);
nor U246 (N_246,In_1657,In_1223);
nor U247 (N_247,In_1949,In_42);
xnor U248 (N_248,In_11,In_194);
nor U249 (N_249,In_1615,In_832);
or U250 (N_250,In_1536,In_14);
or U251 (N_251,In_1915,In_1872);
nand U252 (N_252,In_1043,In_910);
nor U253 (N_253,In_487,In_1356);
nand U254 (N_254,In_1603,In_960);
nor U255 (N_255,In_1497,In_1153);
and U256 (N_256,In_1963,In_1465);
nor U257 (N_257,In_640,In_279);
and U258 (N_258,In_1788,In_1282);
nor U259 (N_259,In_1453,In_72);
nor U260 (N_260,In_838,In_1953);
nor U261 (N_261,In_317,In_182);
or U262 (N_262,In_1234,In_1207);
nand U263 (N_263,In_1970,In_1919);
or U264 (N_264,In_1139,In_1175);
nand U265 (N_265,In_1030,In_682);
or U266 (N_266,In_918,In_445);
nor U267 (N_267,In_454,In_1024);
or U268 (N_268,In_602,In_1554);
or U269 (N_269,In_438,In_1129);
nor U270 (N_270,In_35,In_220);
xnor U271 (N_271,In_153,In_1804);
or U272 (N_272,In_151,In_959);
and U273 (N_273,In_56,In_390);
nor U274 (N_274,In_1782,In_1958);
and U275 (N_275,In_1037,In_299);
xnor U276 (N_276,In_1927,In_1528);
nand U277 (N_277,In_147,In_983);
nor U278 (N_278,In_359,In_1064);
or U279 (N_279,In_989,In_1112);
nand U280 (N_280,In_1320,In_116);
and U281 (N_281,In_641,In_976);
or U282 (N_282,In_1523,In_904);
or U283 (N_283,In_1865,In_612);
and U284 (N_284,In_1629,In_794);
and U285 (N_285,In_1122,In_1040);
or U286 (N_286,In_1860,In_284);
nor U287 (N_287,In_121,In_1906);
nor U288 (N_288,In_221,In_437);
nor U289 (N_289,In_1899,In_540);
nor U290 (N_290,In_1758,In_253);
and U291 (N_291,In_1909,In_1029);
nand U292 (N_292,In_631,In_674);
nand U293 (N_293,In_536,In_1127);
nor U294 (N_294,In_222,In_1420);
or U295 (N_295,In_1377,In_1910);
nor U296 (N_296,In_928,In_280);
and U297 (N_297,In_766,In_1304);
or U298 (N_298,In_1923,In_1399);
or U299 (N_299,In_817,In_1498);
nor U300 (N_300,In_1831,In_1802);
and U301 (N_301,In_1099,In_1471);
nor U302 (N_302,In_994,In_1439);
nor U303 (N_303,In_231,In_504);
nor U304 (N_304,In_377,In_1050);
or U305 (N_305,In_902,In_535);
nand U306 (N_306,In_1079,In_1248);
or U307 (N_307,In_476,In_668);
nor U308 (N_308,In_601,In_626);
nor U309 (N_309,In_1388,In_1888);
or U310 (N_310,In_1150,In_931);
xor U311 (N_311,In_558,In_1460);
nor U312 (N_312,In_1338,In_1152);
xnor U313 (N_313,In_1931,In_958);
nand U314 (N_314,In_1173,In_1353);
nand U315 (N_315,In_48,In_200);
nor U316 (N_316,In_352,In_1286);
and U317 (N_317,In_458,In_166);
or U318 (N_318,In_1068,In_135);
nand U319 (N_319,In_649,In_1485);
nor U320 (N_320,In_378,In_1103);
nor U321 (N_321,In_407,In_662);
xor U322 (N_322,In_1568,In_1182);
xnor U323 (N_323,In_1186,In_1917);
or U324 (N_324,In_945,In_675);
or U325 (N_325,In_1597,In_1443);
nand U326 (N_326,In_203,In_1984);
and U327 (N_327,In_1006,In_1000);
nor U328 (N_328,In_937,In_1754);
or U329 (N_329,In_1590,In_26);
nand U330 (N_330,In_1354,In_880);
xor U331 (N_331,In_1809,In_1749);
nand U332 (N_332,In_130,In_94);
xor U333 (N_333,In_164,In_551);
or U334 (N_334,In_831,In_1262);
or U335 (N_335,In_1707,In_34);
nand U336 (N_336,In_1584,In_475);
nor U337 (N_337,In_683,In_159);
nor U338 (N_338,In_908,In_638);
and U339 (N_339,In_1674,In_835);
nor U340 (N_340,In_384,In_1208);
nand U341 (N_341,In_217,In_1372);
nor U342 (N_342,In_692,In_1488);
or U343 (N_343,In_1602,In_1882);
nand U344 (N_344,In_1803,In_1392);
xor U345 (N_345,In_271,In_655);
xnor U346 (N_346,In_230,In_1863);
nor U347 (N_347,In_1500,In_16);
nand U348 (N_348,In_1643,In_1549);
or U349 (N_349,In_729,In_150);
or U350 (N_350,In_70,In_1796);
xor U351 (N_351,In_1732,In_499);
nand U352 (N_352,In_1003,In_342);
nor U353 (N_353,In_775,In_1343);
and U354 (N_354,In_825,In_1383);
and U355 (N_355,In_1800,In_382);
and U356 (N_356,In_761,In_1839);
nand U357 (N_357,In_782,In_762);
or U358 (N_358,In_985,In_1482);
xnor U359 (N_359,In_502,In_851);
or U360 (N_360,In_769,In_442);
and U361 (N_361,In_993,In_1061);
nand U362 (N_362,In_1218,In_1146);
nand U363 (N_363,In_759,In_1438);
or U364 (N_364,In_1289,In_412);
nor U365 (N_365,In_369,In_447);
nor U366 (N_366,In_1624,In_1314);
and U367 (N_367,In_1480,In_340);
or U368 (N_368,In_1980,In_477);
and U369 (N_369,In_927,In_661);
nand U370 (N_370,In_736,In_446);
or U371 (N_371,In_611,In_1154);
or U372 (N_372,In_1956,In_106);
nor U373 (N_373,In_79,In_774);
nor U374 (N_374,In_922,In_1038);
or U375 (N_375,In_1539,In_1055);
or U376 (N_376,In_1116,In_560);
xnor U377 (N_377,In_350,In_650);
and U378 (N_378,In_440,In_1378);
nand U379 (N_379,In_176,In_1185);
nand U380 (N_380,In_691,In_1188);
nor U381 (N_381,In_1813,In_1737);
nor U382 (N_382,In_1334,In_1322);
nand U383 (N_383,In_1793,In_1891);
or U384 (N_384,In_1769,In_190);
nor U385 (N_385,In_1448,In_1921);
and U386 (N_386,In_27,In_634);
nand U387 (N_387,In_697,In_1974);
nand U388 (N_388,In_1685,In_1020);
nand U389 (N_389,In_1755,In_366);
xnor U390 (N_390,In_1667,In_1071);
or U391 (N_391,In_876,In_1151);
nand U392 (N_392,In_1594,In_310);
nand U393 (N_393,In_1937,In_406);
nand U394 (N_394,In_327,In_281);
xnor U395 (N_395,In_1244,In_1505);
nand U396 (N_396,In_95,In_1833);
or U397 (N_397,In_371,In_846);
and U398 (N_398,In_1466,In_1789);
nor U399 (N_399,In_1128,In_1424);
xor U400 (N_400,In_251,In_919);
xnor U401 (N_401,In_1180,In_1283);
nand U402 (N_402,In_1194,In_935);
nand U403 (N_403,In_43,In_1768);
and U404 (N_404,In_1756,In_120);
or U405 (N_405,In_575,In_1902);
or U406 (N_406,In_764,In_481);
nor U407 (N_407,In_1267,In_432);
nand U408 (N_408,In_853,In_1521);
and U409 (N_409,In_963,In_88);
or U410 (N_410,In_351,In_1542);
nor U411 (N_411,In_1944,In_466);
and U412 (N_412,In_1878,In_787);
and U413 (N_413,In_1035,In_703);
nor U414 (N_414,In_330,In_843);
xnor U415 (N_415,In_430,In_1404);
and U416 (N_416,In_740,In_915);
and U417 (N_417,In_319,In_104);
xnor U418 (N_418,In_1054,In_1329);
xnor U419 (N_419,In_162,In_1111);
or U420 (N_420,In_972,In_1232);
nand U421 (N_421,In_521,In_1174);
nand U422 (N_422,In_1412,In_852);
or U423 (N_423,In_276,In_879);
or U424 (N_424,In_1559,In_522);
nand U425 (N_425,In_1695,In_1058);
or U426 (N_426,In_431,In_173);
or U427 (N_427,In_146,In_1308);
or U428 (N_428,In_178,In_778);
nand U429 (N_429,In_724,In_1261);
nand U430 (N_430,In_868,In_1125);
nor U431 (N_431,In_1405,In_1869);
or U432 (N_432,In_41,In_1108);
or U433 (N_433,In_347,In_1380);
and U434 (N_434,In_425,In_375);
and U435 (N_435,In_1461,In_1219);
nand U436 (N_436,In_1982,In_858);
and U437 (N_437,In_537,In_1625);
nor U438 (N_438,In_568,In_1226);
or U439 (N_439,In_839,In_1396);
and U440 (N_440,In_13,In_665);
nand U441 (N_441,In_689,In_1187);
nor U442 (N_442,In_596,In_409);
nand U443 (N_443,In_1587,In_1846);
or U444 (N_444,In_1476,In_1459);
nand U445 (N_445,In_460,In_671);
nor U446 (N_446,In_1344,In_258);
and U447 (N_447,In_1545,In_1664);
nor U448 (N_448,In_1993,In_617);
nor U449 (N_449,In_1808,In_1530);
nor U450 (N_450,In_282,In_1216);
nand U451 (N_451,In_300,In_156);
xor U452 (N_452,In_1573,In_894);
and U453 (N_453,In_316,In_1981);
nor U454 (N_454,In_812,In_1171);
and U455 (N_455,In_1034,In_293);
nor U456 (N_456,In_1881,In_1246);
xor U457 (N_457,In_107,In_124);
nor U458 (N_458,In_1092,In_287);
nor U459 (N_459,In_1297,In_706);
and U460 (N_460,In_1048,In_615);
or U461 (N_461,In_600,In_1211);
nor U462 (N_462,In_1109,In_1435);
or U463 (N_463,In_1273,In_1726);
and U464 (N_464,In_364,In_1686);
xnor U465 (N_465,In_60,In_1094);
nor U466 (N_466,In_511,In_1241);
or U467 (N_467,In_967,In_849);
or U468 (N_468,In_509,In_620);
xnor U469 (N_469,In_608,In_1575);
nand U470 (N_470,In_1612,In_936);
nand U471 (N_471,In_1330,In_1514);
xnor U472 (N_472,In_1516,In_1660);
and U473 (N_473,In_1303,In_1767);
nor U474 (N_474,In_913,In_1418);
xor U475 (N_475,In_472,In_1916);
and U476 (N_476,In_785,In_1296);
and U477 (N_477,In_1988,In_1259);
and U478 (N_478,In_1583,In_1557);
xor U479 (N_479,In_582,In_1973);
or U480 (N_480,In_1608,In_1221);
nor U481 (N_481,In_209,In_6);
nor U482 (N_482,In_1748,In_341);
and U483 (N_483,In_1256,In_20);
nand U484 (N_484,In_1337,In_1567);
or U485 (N_485,In_592,In_1535);
or U486 (N_486,In_940,In_871);
or U487 (N_487,In_977,In_1898);
nand U488 (N_488,In_1564,In_186);
and U489 (N_489,In_1366,In_1069);
or U490 (N_490,In_1824,In_129);
or U491 (N_491,In_1251,In_401);
nor U492 (N_492,In_1901,In_1634);
nand U493 (N_493,In_1301,In_605);
and U494 (N_494,In_1941,In_1098);
or U495 (N_495,In_185,In_507);
nand U496 (N_496,In_911,In_955);
nor U497 (N_497,In_336,In_738);
or U498 (N_498,In_1487,In_1017);
xnor U499 (N_499,In_314,In_1126);
or U500 (N_500,N_481,In_179);
nor U501 (N_501,In_758,N_138);
xor U502 (N_502,N_186,In_1170);
nand U503 (N_503,In_494,N_368);
and U504 (N_504,N_320,In_1347);
nor U505 (N_505,In_451,In_616);
nor U506 (N_506,In_172,In_1765);
nor U507 (N_507,In_679,N_196);
nor U508 (N_508,N_98,In_23);
nand U509 (N_509,In_323,In_856);
nor U510 (N_510,In_1149,N_52);
nor U511 (N_511,In_906,N_222);
xor U512 (N_512,In_556,N_273);
nor U513 (N_513,In_688,In_1986);
nor U514 (N_514,In_1169,In_491);
nand U515 (N_515,In_604,In_1740);
nor U516 (N_516,In_1604,In_1799);
or U517 (N_517,In_708,N_231);
and U518 (N_518,In_1745,N_218);
and U519 (N_519,N_499,N_346);
or U520 (N_520,N_289,N_397);
and U521 (N_521,In_544,In_1633);
xnor U522 (N_522,In_500,In_1853);
or U523 (N_523,In_198,In_1400);
nor U524 (N_524,In_1935,In_1893);
nor U525 (N_525,N_295,N_479);
or U526 (N_526,N_369,In_508);
or U527 (N_527,In_1742,In_452);
nor U528 (N_528,In_1997,In_1449);
nand U529 (N_529,In_199,In_990);
and U530 (N_530,In_670,N_469);
nand U531 (N_531,In_468,N_460);
nand U532 (N_532,In_730,In_1566);
or U533 (N_533,In_1416,In_1398);
or U534 (N_534,In_722,In_552);
nor U535 (N_535,In_1847,In_1733);
nor U536 (N_536,N_272,In_715);
and U537 (N_537,In_339,In_1022);
and U538 (N_538,In_800,In_325);
and U539 (N_539,N_213,In_1617);
nand U540 (N_540,In_243,In_128);
or U541 (N_541,In_848,In_555);
nand U542 (N_542,N_8,In_1178);
and U543 (N_543,In_686,In_404);
xor U544 (N_544,In_119,N_489);
and U545 (N_545,N_184,In_854);
nor U546 (N_546,N_119,In_1110);
nor U547 (N_547,In_739,In_1428);
and U548 (N_548,In_970,In_125);
or U549 (N_549,In_737,In_790);
or U550 (N_550,N_71,In_362);
nor U551 (N_551,In_698,N_109);
and U552 (N_552,N_454,In_1515);
xor U553 (N_553,In_1513,In_1840);
and U554 (N_554,N_359,N_327);
and U555 (N_555,In_1546,N_166);
or U556 (N_556,N_363,In_211);
nor U557 (N_557,N_194,In_1894);
and U558 (N_558,In_1096,In_845);
and U559 (N_559,In_1360,N_170);
nor U560 (N_560,N_490,N_461);
and U561 (N_561,In_645,N_115);
or U562 (N_562,In_1272,In_236);
or U563 (N_563,In_149,In_1783);
nor U564 (N_564,N_10,N_235);
nand U565 (N_565,In_779,N_107);
and U566 (N_566,N_313,In_506);
and U567 (N_567,In_1331,In_1948);
and U568 (N_568,In_667,In_872);
nand U569 (N_569,N_134,N_216);
nand U570 (N_570,N_195,N_446);
and U571 (N_571,N_40,N_258);
nand U572 (N_572,In_1924,In_1741);
or U573 (N_573,In_12,In_233);
and U574 (N_574,N_355,In_1862);
nor U575 (N_575,In_554,In_357);
or U576 (N_576,N_285,In_471);
or U577 (N_577,In_827,In_1421);
nor U578 (N_578,In_796,In_75);
or U579 (N_579,N_161,In_818);
and U580 (N_580,In_1805,N_314);
or U581 (N_581,N_457,In_1959);
or U582 (N_582,N_243,In_1348);
or U583 (N_583,N_212,In_1591);
and U584 (N_584,N_20,In_36);
nand U585 (N_585,In_962,In_1252);
nand U586 (N_586,In_1841,N_299);
nor U587 (N_587,In_1265,In_1121);
nor U588 (N_588,N_117,In_1276);
or U589 (N_589,In_1431,N_277);
nor U590 (N_590,N_31,N_56);
or U591 (N_591,N_249,In_881);
nor U592 (N_592,N_447,N_151);
nor U593 (N_593,In_1105,In_1202);
nor U594 (N_594,In_814,N_191);
nand U595 (N_595,N_79,In_321);
or U596 (N_596,In_1452,In_1138);
nor U597 (N_597,N_264,In_1456);
nor U598 (N_598,In_158,In_677);
or U599 (N_599,In_826,In_1217);
or U600 (N_600,N_392,In_714);
xnor U601 (N_601,In_74,In_900);
nand U602 (N_602,In_1628,N_496);
nand U603 (N_603,In_1203,In_520);
nor U604 (N_604,N_57,In_630);
nor U605 (N_605,N_373,In_461);
xnor U606 (N_606,N_303,In_1572);
nor U607 (N_607,In_1277,N_497);
xnor U608 (N_608,N_174,In_647);
and U609 (N_609,N_211,In_1143);
and U610 (N_610,In_1473,In_780);
nand U611 (N_611,In_783,In_467);
or U612 (N_612,In_244,In_701);
nand U613 (N_613,N_436,In_1911);
xor U614 (N_614,In_1908,N_217);
xor U615 (N_615,In_992,In_1845);
and U616 (N_616,N_63,In_1580);
and U617 (N_617,N_493,In_218);
and U618 (N_618,In_197,In_1410);
xor U619 (N_619,N_88,In_823);
nor U620 (N_620,N_55,N_414);
nor U621 (N_621,N_492,In_1728);
nand U622 (N_622,In_1747,In_1550);
nand U623 (N_623,In_541,In_238);
nor U624 (N_624,In_71,N_43);
nand U625 (N_625,In_322,In_96);
or U626 (N_626,N_49,N_472);
nor U627 (N_627,In_1386,N_390);
or U628 (N_628,In_32,N_404);
nor U629 (N_629,In_1522,N_293);
nand U630 (N_630,In_1090,In_1708);
and U631 (N_631,In_816,In_374);
or U632 (N_632,In_664,N_155);
or U633 (N_633,In_1713,N_330);
or U634 (N_634,N_485,In_713);
nor U635 (N_635,N_387,In_748);
nand U636 (N_636,In_548,N_141);
and U637 (N_637,In_367,In_1653);
or U638 (N_638,N_411,N_477);
xnor U639 (N_639,N_149,In_1619);
or U640 (N_640,In_337,In_262);
nand U641 (N_641,In_1985,In_723);
or U642 (N_642,In_947,N_225);
nand U643 (N_643,In_1315,N_97);
or U644 (N_644,In_1943,In_1764);
and U645 (N_645,In_65,N_331);
nor U646 (N_646,In_1999,In_1285);
or U647 (N_647,In_984,N_431);
nor U648 (N_648,In_441,N_190);
and U649 (N_649,In_329,In_632);
nor U650 (N_650,In_1613,In_1781);
nor U651 (N_651,N_172,N_33);
nor U652 (N_652,N_100,In_1763);
nand U653 (N_653,In_1807,In_1407);
or U654 (N_654,In_161,N_257);
nand U655 (N_655,In_252,In_389);
nand U656 (N_656,In_1457,In_265);
and U657 (N_657,N_61,In_226);
nand U658 (N_658,In_1358,N_202);
nor U659 (N_659,N_266,In_1790);
nor U660 (N_660,N_144,In_1242);
nor U661 (N_661,In_1946,In_1688);
nand U662 (N_662,In_673,In_181);
nor U663 (N_663,In_1450,N_72);
nand U664 (N_664,In_402,N_173);
or U665 (N_665,In_397,In_1113);
nand U666 (N_666,In_69,N_104);
nand U667 (N_667,In_1163,In_356);
nand U668 (N_668,N_127,In_1346);
or U669 (N_669,N_23,In_1397);
nand U670 (N_670,In_1543,N_69);
nor U671 (N_671,In_1960,In_1166);
nor U672 (N_672,In_291,N_304);
nand U673 (N_673,N_405,In_1877);
nand U674 (N_674,In_1818,In_1123);
xor U675 (N_675,In_1033,N_244);
nor U676 (N_676,In_860,In_1394);
nor U677 (N_677,In_1700,In_67);
nand U678 (N_678,N_241,In_773);
and U679 (N_679,N_451,In_1992);
or U680 (N_680,In_1810,N_77);
nand U681 (N_681,In_386,In_516);
xnor U682 (N_682,In_435,In_1481);
nand U683 (N_683,N_182,In_1693);
and U684 (N_684,In_1097,In_335);
or U685 (N_685,In_490,In_1694);
nand U686 (N_686,N_408,In_969);
nor U687 (N_687,In_1197,N_311);
or U688 (N_688,In_1716,In_76);
or U689 (N_689,N_70,In_1025);
nor U690 (N_690,In_1592,N_486);
nand U691 (N_691,In_1222,In_926);
nand U692 (N_692,N_201,In_566);
and U693 (N_693,In_1235,N_366);
nor U694 (N_694,In_496,N_324);
and U695 (N_695,In_1614,In_1389);
nand U696 (N_696,In_1240,In_1371);
nor U697 (N_697,In_1574,In_760);
or U698 (N_698,In_444,In_1577);
and U699 (N_699,N_340,In_333);
and U700 (N_700,In_1835,In_1826);
and U701 (N_701,In_1374,In_862);
nor U702 (N_702,N_158,In_570);
and U703 (N_703,In_449,N_78);
nor U704 (N_704,In_1680,N_412);
nor U705 (N_705,N_262,N_465);
xnor U706 (N_706,In_45,In_1229);
or U707 (N_707,In_1047,N_13);
and U708 (N_708,In_1526,In_1585);
nand U709 (N_709,In_702,In_1446);
nor U710 (N_710,N_329,In_1773);
nor U711 (N_711,N_146,N_424);
nor U712 (N_712,In_1160,N_418);
or U713 (N_713,In_195,In_1616);
nor U714 (N_714,N_38,In_804);
and U715 (N_715,N_251,N_448);
or U716 (N_716,N_86,N_323);
xnor U717 (N_717,In_1168,In_343);
and U718 (N_718,In_1662,In_413);
xnor U719 (N_719,N_28,In_1239);
or U720 (N_720,N_420,In_306);
and U721 (N_721,In_866,In_1691);
or U722 (N_722,N_374,In_1328);
or U723 (N_723,In_1403,In_1779);
nand U724 (N_724,In_155,N_47);
and U725 (N_725,N_254,In_1477);
and U726 (N_726,N_268,N_364);
nor U727 (N_727,N_341,In_419);
nand U728 (N_728,In_82,In_875);
nor U729 (N_729,In_1401,In_1164);
nor U730 (N_730,N_230,In_1470);
or U731 (N_731,N_358,In_1760);
nor U732 (N_732,In_519,In_145);
and U733 (N_733,N_3,N_95);
nor U734 (N_734,In_808,In_295);
nor U735 (N_735,N_371,N_16);
nand U736 (N_736,N_440,In_907);
nand U737 (N_737,In_1507,In_1703);
nor U738 (N_738,In_1483,In_175);
and U739 (N_739,In_1134,In_840);
xnor U740 (N_740,N_96,In_1724);
and U741 (N_741,N_206,In_798);
nand U742 (N_742,N_287,In_86);
and U743 (N_743,N_322,N_379);
nor U744 (N_744,N_99,In_1524);
and U745 (N_745,In_1996,In_1502);
and U746 (N_746,N_396,In_1544);
nor U747 (N_747,N_62,N_162);
xor U748 (N_748,In_1209,In_986);
nand U749 (N_749,In_1920,N_430);
or U750 (N_750,In_1672,In_581);
nor U751 (N_751,In_1206,In_268);
xnor U752 (N_752,In_187,In_998);
nand U753 (N_753,N_315,N_383);
and U754 (N_754,In_1622,N_487);
or U755 (N_755,In_266,In_1827);
nand U756 (N_756,In_152,In_586);
nor U757 (N_757,In_214,In_0);
nor U758 (N_758,In_1718,In_464);
nand U759 (N_759,N_80,In_563);
or U760 (N_760,In_1552,In_1451);
nor U761 (N_761,N_349,N_260);
and U762 (N_762,In_887,In_1547);
and U763 (N_763,N_197,In_1369);
or U764 (N_764,In_1639,In_1145);
or U765 (N_765,N_402,N_375);
and U766 (N_766,In_699,In_524);
and U767 (N_767,In_30,In_1663);
nand U768 (N_768,In_421,N_399);
or U769 (N_769,In_1669,N_85);
and U770 (N_770,In_1056,In_113);
nor U771 (N_771,In_712,In_1214);
nor U772 (N_772,N_459,In_1442);
nand U773 (N_773,In_828,In_975);
or U774 (N_774,In_1979,In_1864);
nand U775 (N_775,In_1028,In_1510);
and U776 (N_776,In_1441,In_1569);
nand U777 (N_777,N_473,N_238);
and U778 (N_778,In_770,N_132);
xnor U779 (N_779,In_741,In_627);
nor U780 (N_780,In_453,In_1719);
nor U781 (N_781,In_66,N_35);
or U782 (N_782,In_1842,N_288);
nand U783 (N_783,In_1509,N_438);
and U784 (N_784,In_422,N_279);
or U785 (N_785,N_270,In_1075);
nand U786 (N_786,N_193,In_1532);
nand U787 (N_787,In_659,In_1181);
xnor U788 (N_788,In_405,In_1141);
or U789 (N_789,In_996,In_1009);
nand U790 (N_790,In_917,N_22);
and U791 (N_791,In_574,N_68);
or U792 (N_792,N_164,N_471);
or U793 (N_793,N_7,N_284);
nor U794 (N_794,In_354,In_1640);
nor U795 (N_795,In_1570,N_250);
nor U796 (N_796,In_1971,In_1635);
nor U797 (N_797,N_415,In_1342);
or U798 (N_798,In_275,In_415);
or U799 (N_799,In_1527,In_1081);
nor U800 (N_800,N_318,N_419);
or U801 (N_801,In_577,In_1332);
nor U802 (N_802,In_223,In_1787);
or U803 (N_803,In_971,N_200);
or U804 (N_804,N_9,N_105);
nor U805 (N_805,In_1156,In_277);
nand U806 (N_806,N_307,In_1858);
nor U807 (N_807,In_307,In_1887);
or U808 (N_808,In_981,N_370);
and U809 (N_809,In_1884,In_1263);
and U810 (N_810,In_1900,N_333);
and U811 (N_811,N_253,In_1190);
xor U812 (N_812,N_495,In_553);
nand U813 (N_813,N_208,In_1599);
and U814 (N_814,In_1725,N_305);
nand U815 (N_815,In_140,In_1825);
or U816 (N_816,In_1266,N_136);
and U817 (N_817,In_90,In_308);
nor U818 (N_818,In_1681,N_417);
nor U819 (N_819,In_1236,N_357);
and U820 (N_820,N_456,In_1422);
and U821 (N_821,In_855,N_348);
or U822 (N_822,N_25,In_1734);
and U823 (N_823,N_381,In_1702);
or U824 (N_824,In_1555,N_34);
or U825 (N_825,In_1237,N_367);
nand U826 (N_826,In_1812,In_585);
or U827 (N_827,In_1670,N_214);
nor U828 (N_828,In_1848,In_1965);
nor U829 (N_829,In_561,In_1644);
and U830 (N_830,N_75,N_463);
or U831 (N_831,In_806,In_768);
or U832 (N_832,In_1469,In_965);
nor U833 (N_833,N_179,N_433);
nor U834 (N_834,N_67,N_177);
nor U835 (N_835,N_17,N_306);
nor U836 (N_836,In_580,In_346);
nand U837 (N_837,N_29,N_388);
or U838 (N_838,N_156,In_1746);
nand U839 (N_839,In_789,N_178);
nor U840 (N_840,N_92,In_1086);
nor U841 (N_841,In_1647,In_1291);
or U842 (N_842,In_1593,In_1723);
or U843 (N_843,In_1046,In_545);
nor U844 (N_844,N_292,N_432);
nand U845 (N_845,N_278,N_83);
nand U846 (N_846,In_1093,In_1199);
and U847 (N_847,In_1434,N_345);
nand U848 (N_848,In_1250,N_227);
nor U849 (N_849,In_1299,In_1642);
or U850 (N_850,In_1632,In_474);
nor U851 (N_851,In_1778,In_1245);
or U852 (N_852,N_215,N_312);
or U853 (N_853,N_131,N_393);
nand U854 (N_854,N_452,In_1198);
xor U855 (N_855,In_1124,N_188);
or U856 (N_856,In_974,N_110);
nand U857 (N_857,In_170,In_1630);
or U858 (N_858,N_114,In_376);
or U859 (N_859,In_572,In_469);
and U860 (N_860,N_93,In_1874);
and U861 (N_861,N_353,In_725);
and U862 (N_862,In_259,In_1830);
nor U863 (N_863,In_1990,N_143);
or U864 (N_864,N_439,In_952);
and U865 (N_865,In_315,N_391);
or U866 (N_866,In_728,In_934);
nand U867 (N_867,N_89,N_219);
or U868 (N_868,N_37,In_462);
nand U869 (N_869,In_1011,In_296);
or U870 (N_870,In_653,In_921);
xnor U871 (N_871,N_468,N_30);
nor U872 (N_872,In_115,N_476);
nand U873 (N_873,In_257,In_1);
or U874 (N_874,N_269,In_954);
nand U875 (N_875,In_1626,N_122);
nor U876 (N_876,In_864,In_1689);
nor U877 (N_877,N_297,N_167);
xor U878 (N_878,In_1311,N_263);
nor U879 (N_879,N_44,N_239);
and U880 (N_880,N_450,N_106);
and U881 (N_881,In_1777,N_32);
or U882 (N_882,In_982,In_1890);
nand U883 (N_883,In_720,In_1606);
nor U884 (N_884,In_1032,In_24);
and U885 (N_885,N_221,In_1967);
or U886 (N_886,N_39,In_1772);
nand U887 (N_887,In_1852,N_470);
or U888 (N_888,In_1829,In_1607);
nor U889 (N_889,In_98,In_742);
nand U890 (N_890,N_220,In_1977);
nand U891 (N_891,N_475,In_639);
nor U892 (N_892,N_422,In_1652);
nand U893 (N_893,In_332,N_398);
or U894 (N_894,In_1215,N_224);
nor U895 (N_895,N_280,In_492);
nand U896 (N_896,In_1062,In_127);
nor U897 (N_897,N_232,In_274);
nor U898 (N_898,In_1957,N_81);
nor U899 (N_899,In_1578,In_1936);
and U900 (N_900,In_997,In_1861);
nand U901 (N_901,In_1479,In_771);
nand U902 (N_902,N_434,In_250);
and U903 (N_903,In_1350,N_176);
and U904 (N_904,N_484,N_181);
or U905 (N_905,N_240,In_1376);
and U906 (N_906,In_1114,N_228);
nor U907 (N_907,In_1637,N_283);
nor U908 (N_908,In_1432,In_1310);
and U909 (N_909,In_372,In_448);
xor U910 (N_910,N_118,In_1458);
and U911 (N_911,In_824,In_672);
xor U912 (N_912,In_755,In_1089);
nand U913 (N_913,N_296,In_1930);
nor U914 (N_914,N_441,N_189);
nand U915 (N_915,N_261,In_427);
and U916 (N_916,In_1875,N_108);
nand U917 (N_917,In_1001,N_54);
xnor U918 (N_918,In_1601,In_732);
nor U919 (N_919,In_924,N_223);
or U920 (N_920,In_247,N_103);
or U921 (N_921,N_474,In_1677);
or U922 (N_922,In_538,In_261);
and U923 (N_923,In_1118,In_666);
nor U924 (N_924,N_123,In_142);
or U925 (N_925,N_425,In_457);
nor U926 (N_926,In_707,N_300);
nor U927 (N_927,In_1227,In_1440);
nor U928 (N_928,N_60,N_163);
or U929 (N_929,In_1288,In_1183);
or U930 (N_930,N_207,In_1478);
or U931 (N_931,N_187,In_1393);
or U932 (N_932,In_301,In_896);
and U933 (N_933,In_549,In_1705);
and U934 (N_934,In_901,In_324);
nor U935 (N_935,In_1131,In_1204);
and U936 (N_936,In_17,N_462);
and U937 (N_937,In_1589,In_1867);
and U938 (N_938,N_365,In_1041);
and U939 (N_939,N_302,In_1018);
nor U940 (N_940,In_1621,N_410);
nor U941 (N_941,In_138,In_44);
nand U942 (N_942,In_1279,In_473);
or U943 (N_943,In_1077,In_1618);
nand U944 (N_944,N_413,N_265);
xnor U945 (N_945,In_598,In_533);
nand U946 (N_946,In_141,In_1274);
nand U947 (N_947,In_930,In_944);
xnor U948 (N_948,In_283,In_897);
nand U949 (N_949,In_1224,In_1715);
xnor U950 (N_950,N_157,In_624);
and U951 (N_951,In_916,N_234);
or U952 (N_952,In_1814,In_1711);
nor U953 (N_953,In_272,N_328);
or U954 (N_954,In_320,N_360);
or U955 (N_955,In_1305,N_301);
nand U956 (N_956,In_189,N_111);
xor U957 (N_957,In_1053,N_5);
and U958 (N_958,In_1596,In_264);
xor U959 (N_959,In_1463,In_584);
nor U960 (N_960,In_246,In_1797);
xor U961 (N_961,In_813,In_196);
xnor U962 (N_962,In_456,N_427);
xor U963 (N_963,N_19,In_802);
or U964 (N_964,N_229,In_933);
nand U965 (N_965,In_207,In_1966);
xnor U966 (N_966,In_1495,In_1490);
nand U967 (N_967,In_1856,N_12);
and U968 (N_968,N_325,In_1731);
or U969 (N_969,N_210,In_144);
nor U970 (N_970,In_1964,In_235);
nand U971 (N_971,In_1692,In_1646);
and U972 (N_972,In_388,In_1661);
xor U973 (N_973,In_750,In_1162);
nor U974 (N_974,N_84,In_1871);
nor U975 (N_975,In_681,N_1);
nand U976 (N_976,In_1727,In_834);
nand U977 (N_977,N_247,N_147);
and U978 (N_978,In_1690,N_209);
and U979 (N_979,In_717,N_154);
nor U980 (N_980,N_137,In_635);
and U981 (N_981,In_716,N_233);
nor U982 (N_982,In_1770,In_781);
xor U983 (N_983,In_517,In_1264);
nor U984 (N_984,In_38,In_1088);
xnor U985 (N_985,In_734,In_131);
or U986 (N_986,In_559,N_429);
or U987 (N_987,In_1414,In_224);
nor U988 (N_988,N_421,In_801);
nand U989 (N_989,In_1817,N_2);
nand U990 (N_990,In_370,N_455);
and U991 (N_991,N_126,In_1701);
and U992 (N_992,In_450,In_837);
nor U993 (N_993,In_1503,In_78);
nand U994 (N_994,N_0,In_1786);
or U995 (N_995,In_1294,In_1645);
and U996 (N_996,In_1177,N_11);
nor U997 (N_997,In_1903,In_245);
or U998 (N_998,In_387,In_1811);
or U999 (N_999,In_1321,N_347);
or U1000 (N_1000,N_684,In_498);
nand U1001 (N_1001,In_1238,N_906);
nor U1002 (N_1002,N_946,In_1659);
or U1003 (N_1003,N_663,N_532);
or U1004 (N_1004,N_237,N_896);
nand U1005 (N_1005,N_437,N_308);
or U1006 (N_1006,N_753,N_316);
or U1007 (N_1007,N_389,N_929);
or U1008 (N_1008,N_674,N_483);
nor U1009 (N_1009,N_651,N_394);
nor U1010 (N_1010,In_590,In_398);
and U1011 (N_1011,In_1200,N_872);
or U1012 (N_1012,In_523,N_913);
and U1013 (N_1013,In_1918,N_534);
or U1014 (N_1014,N_925,N_918);
or U1015 (N_1015,N_782,N_698);
and U1016 (N_1016,N_967,N_509);
nand U1017 (N_1017,In_9,N_537);
and U1018 (N_1018,In_1654,N_153);
nand U1019 (N_1019,In_939,In_847);
and U1020 (N_1020,N_423,N_290);
nand U1021 (N_1021,N_703,N_664);
or U1022 (N_1022,N_638,In_842);
and U1023 (N_1023,N_622,N_763);
nand U1024 (N_1024,In_1873,In_1656);
or U1025 (N_1025,In_403,N_678);
nor U1026 (N_1026,N_344,N_994);
nand U1027 (N_1027,In_294,N_718);
and U1028 (N_1028,N_943,N_640);
or U1029 (N_1029,N_591,In_1844);
xor U1030 (N_1030,N_354,N_708);
and U1031 (N_1031,N_866,N_581);
nor U1032 (N_1032,N_593,In_1759);
or U1033 (N_1033,In_658,In_784);
xnor U1034 (N_1034,N_855,In_1370);
nand U1035 (N_1035,N_652,In_1284);
nand U1036 (N_1036,N_931,In_514);
and U1037 (N_1037,In_950,In_613);
and U1038 (N_1038,N_342,N_771);
nand U1039 (N_1039,N_554,N_934);
or U1040 (N_1040,N_976,In_1699);
nand U1041 (N_1041,N_491,N_999);
nand U1042 (N_1042,In_1945,In_216);
nand U1043 (N_1043,In_1940,In_1581);
nor U1044 (N_1044,N_814,N_58);
and U1045 (N_1045,N_794,N_121);
and U1046 (N_1046,N_755,N_849);
nand U1047 (N_1047,N_53,N_565);
or U1048 (N_1048,In_205,N_867);
nand U1049 (N_1049,N_91,N_873);
and U1050 (N_1050,In_865,In_426);
and U1051 (N_1051,N_901,In_1379);
nor U1052 (N_1052,N_401,In_1268);
nand U1053 (N_1053,In_1066,N_274);
or U1054 (N_1054,N_750,N_605);
or U1055 (N_1055,N_525,N_989);
and U1056 (N_1056,N_395,N_799);
and U1057 (N_1057,In_1785,In_1070);
xnor U1058 (N_1058,N_426,N_518);
and U1059 (N_1059,N_572,N_988);
nor U1060 (N_1060,N_571,N_821);
nor U1061 (N_1061,N_893,N_942);
or U1062 (N_1062,N_993,In_515);
and U1063 (N_1063,N_898,N_919);
or U1064 (N_1064,N_905,N_510);
and U1065 (N_1065,N_130,N_842);
or U1066 (N_1066,In_463,In_844);
xnor U1067 (N_1067,N_948,N_908);
and U1068 (N_1068,N_317,In_893);
nand U1069 (N_1069,N_608,In_859);
or U1070 (N_1070,In_1415,In_603);
nand U1071 (N_1071,N_14,N_668);
and U1072 (N_1072,N_659,N_563);
xnor U1073 (N_1073,In_180,N_959);
xor U1074 (N_1074,In_47,In_1167);
nor U1075 (N_1075,N_886,N_998);
nand U1076 (N_1076,N_734,In_735);
nand U1077 (N_1077,In_895,N_667);
and U1078 (N_1078,In_1359,N_791);
nand U1079 (N_1079,N_825,N_310);
or U1080 (N_1080,N_751,In_1257);
nand U1081 (N_1081,In_1489,N_520);
and U1082 (N_1082,N_498,N_850);
and U1083 (N_1083,N_639,In_1402);
nor U1084 (N_1084,N_735,In_614);
nor U1085 (N_1085,In_1287,N_528);
and U1086 (N_1086,N_533,N_4);
or U1087 (N_1087,In_669,N_624);
or U1088 (N_1088,N_592,N_183);
xor U1089 (N_1089,N_599,In_1571);
nand U1090 (N_1090,N_797,N_530);
nand U1091 (N_1091,N_949,N_772);
nor U1092 (N_1092,In_439,N_938);
and U1093 (N_1093,N_321,In_420);
xor U1094 (N_1094,In_344,N_647);
nand U1095 (N_1095,N_150,In_793);
nor U1096 (N_1096,N_578,N_672);
xnor U1097 (N_1097,N_76,N_291);
nand U1098 (N_1098,In_288,In_424);
nor U1099 (N_1099,N_676,N_618);
nor U1100 (N_1100,In_400,In_1298);
or U1101 (N_1101,N_553,In_1300);
and U1102 (N_1102,N_890,N_94);
xor U1103 (N_1103,N_606,N_728);
and U1104 (N_1104,N_981,N_386);
and U1105 (N_1105,In_167,N_248);
nor U1106 (N_1106,In_528,N_653);
xor U1107 (N_1107,In_122,In_1540);
or U1108 (N_1108,In_154,In_1975);
xor U1109 (N_1109,In_920,In_1333);
nor U1110 (N_1110,N_745,N_406);
and U1111 (N_1111,In_654,In_1365);
or U1112 (N_1112,In_1044,In_1243);
nor U1113 (N_1113,N_900,N_936);
nor U1114 (N_1114,N_756,N_644);
and U1115 (N_1115,N_677,In_1225);
and U1116 (N_1116,N_853,In_248);
nand U1117 (N_1117,N_769,In_1119);
nand U1118 (N_1118,N_969,N_688);
or U1119 (N_1119,N_875,N_566);
xnor U1120 (N_1120,N_958,In_1375);
or U1121 (N_1121,N_654,N_48);
nand U1122 (N_1122,N_540,N_953);
nand U1123 (N_1123,In_1275,N_350);
or U1124 (N_1124,N_634,In_1340);
and U1125 (N_1125,N_726,N_727);
or U1126 (N_1126,N_552,N_569);
nor U1127 (N_1127,N_6,In_841);
nor U1128 (N_1128,N_560,N_813);
and U1129 (N_1129,N_990,In_278);
nor U1130 (N_1130,In_1706,N_570);
nand U1131 (N_1131,N_236,N_276);
or U1132 (N_1132,N_812,N_478);
nor U1133 (N_1133,N_620,In_772);
and U1134 (N_1134,N_705,N_862);
nand U1135 (N_1135,In_1373,N_561);
nand U1136 (N_1136,N_818,N_847);
nor U1137 (N_1137,N_830,N_309);
xor U1138 (N_1138,N_376,N_861);
or U1139 (N_1139,N_632,N_579);
and U1140 (N_1140,N_736,In_1387);
and U1141 (N_1141,In_1309,N_74);
xor U1142 (N_1142,N_90,In_1280);
nand U1143 (N_1143,N_687,N_722);
or U1144 (N_1144,N_549,N_758);
nand U1145 (N_1145,N_116,N_543);
nor U1146 (N_1146,N_159,N_779);
nand U1147 (N_1147,N_294,N_603);
or U1148 (N_1148,In_1336,In_754);
nor U1149 (N_1149,In_909,N_914);
and U1150 (N_1150,In_1324,N_500);
and U1151 (N_1151,N_453,In_597);
xnor U1152 (N_1152,N_878,N_980);
xnor U1153 (N_1153,N_643,In_629);
nand U1154 (N_1154,N_256,N_378);
nand U1155 (N_1155,N_595,N_766);
and U1156 (N_1156,N_774,N_319);
nand U1157 (N_1157,N_613,N_140);
and U1158 (N_1158,N_752,In_1007);
nand U1159 (N_1159,N_562,In_225);
or U1160 (N_1160,N_556,N_584);
or U1161 (N_1161,N_858,In_1201);
nor U1162 (N_1162,In_443,In_177);
nor U1163 (N_1163,N_259,N_573);
and U1164 (N_1164,In_1493,N_171);
nand U1165 (N_1165,N_361,N_916);
nand U1166 (N_1166,In_501,In_1709);
and U1167 (N_1167,N_702,N_675);
or U1168 (N_1168,N_860,In_1683);
nor U1169 (N_1169,N_741,N_686);
nor U1170 (N_1170,N_695,In_543);
and U1171 (N_1171,N_596,N_882);
or U1172 (N_1172,In_718,In_756);
nor U1173 (N_1173,N_623,In_1687);
or U1174 (N_1174,In_749,N_586);
nand U1175 (N_1175,N_826,In_304);
or U1176 (N_1176,N_910,In_49);
nand U1177 (N_1177,In_923,N_742);
or U1178 (N_1178,In_1561,In_21);
or U1179 (N_1179,N_641,N_604);
nand U1180 (N_1180,N_614,In_830);
nor U1181 (N_1181,N_912,N_619);
nor U1182 (N_1182,In_309,N_899);
and U1183 (N_1183,In_721,In_1650);
nand U1184 (N_1184,N_600,N_845);
or U1185 (N_1185,N_955,N_458);
nor U1186 (N_1186,N_356,N_793);
nand U1187 (N_1187,In_727,In_417);
nor U1188 (N_1188,N_746,N_715);
xor U1189 (N_1189,N_185,In_1231);
or U1190 (N_1190,In_4,In_660);
xor U1191 (N_1191,N_538,N_242);
and U1192 (N_1192,In_1474,N_598);
or U1193 (N_1193,N_656,In_819);
nand U1194 (N_1194,In_656,In_54);
nand U1195 (N_1195,N_822,N_337);
and U1196 (N_1196,N_710,In_531);
or U1197 (N_1197,N_385,N_977);
and U1198 (N_1198,In_1885,In_486);
or U1199 (N_1199,In_1074,N_550);
or U1200 (N_1200,In_1520,N_635);
or U1201 (N_1201,N_515,N_986);
xor U1202 (N_1202,N_773,N_887);
nand U1203 (N_1203,In_1462,N_521);
nor U1204 (N_1204,N_165,In_267);
or U1205 (N_1205,N_507,In_15);
xor U1206 (N_1206,In_28,N_951);
or U1207 (N_1207,N_42,In_593);
xor U1208 (N_1208,N_494,N_739);
nand U1209 (N_1209,In_1429,N_545);
or U1210 (N_1210,N_542,N_780);
nor U1211 (N_1211,In_1494,N_82);
and U1212 (N_1212,N_978,N_636);
nor U1213 (N_1213,In_1115,N_711);
nor U1214 (N_1214,N_941,N_807);
nor U1215 (N_1215,In_318,N_41);
xor U1216 (N_1216,N_926,N_546);
and U1217 (N_1217,In_392,N_947);
nand U1218 (N_1218,N_940,In_836);
and U1219 (N_1219,N_798,N_963);
nor U1220 (N_1220,N_120,N_135);
and U1221 (N_1221,N_874,N_876);
and U1222 (N_1222,N_516,In_619);
xor U1223 (N_1223,N_51,N_838);
and U1224 (N_1224,N_610,In_255);
nor U1225 (N_1225,N_637,N_693);
xor U1226 (N_1226,N_985,N_881);
nor U1227 (N_1227,N_602,In_1212);
and U1228 (N_1228,In_1823,N_911);
or U1229 (N_1229,N_823,In_470);
nand U1230 (N_1230,In_1795,N_298);
nor U1231 (N_1231,In_1939,N_588);
xnor U1232 (N_1232,N_894,In_1159);
nor U1233 (N_1233,N_840,N_956);
nor U1234 (N_1234,In_652,N_879);
nand U1235 (N_1235,In_1744,In_979);
xor U1236 (N_1236,N_633,In_1954);
nor U1237 (N_1237,In_1317,In_932);
and U1238 (N_1238,N_738,N_199);
nor U1239 (N_1239,In_805,N_657);
nand U1240 (N_1240,N_760,In_1638);
nand U1241 (N_1241,N_351,N_336);
and U1242 (N_1242,N_601,In_59);
and U1243 (N_1243,In_1083,In_1609);
nand U1244 (N_1244,In_694,In_1648);
nand U1245 (N_1245,In_1444,N_551);
xnor U1246 (N_1246,In_434,In_89);
and U1247 (N_1247,N_145,N_897);
nand U1248 (N_1248,In_139,N_964);
and U1249 (N_1249,N_286,In_3);
and U1250 (N_1250,N_282,N_863);
nor U1251 (N_1251,N_721,In_105);
xor U1252 (N_1252,In_1426,N_820);
nand U1253 (N_1253,In_1883,N_271);
nor U1254 (N_1254,N_973,N_714);
nor U1255 (N_1255,N_576,N_903);
or U1256 (N_1256,In_408,N_809);
nand U1257 (N_1257,N_526,N_723);
nand U1258 (N_1258,In_599,N_281);
and U1259 (N_1259,N_706,N_267);
and U1260 (N_1260,In_949,N_856);
nand U1261 (N_1261,N_555,In_1969);
and U1262 (N_1262,In_878,N_700);
nand U1263 (N_1263,In_1560,In_1016);
nand U1264 (N_1264,In_1620,N_859);
nand U1265 (N_1265,In_101,N_529);
nand U1266 (N_1266,N_811,N_865);
nand U1267 (N_1267,N_933,N_255);
or U1268 (N_1268,N_442,N_697);
and U1269 (N_1269,In_5,In_1914);
nor U1270 (N_1270,N_169,N_148);
nand U1271 (N_1271,N_102,N_343);
and U1272 (N_1272,N_558,In_379);
xor U1273 (N_1273,N_466,N_732);
nand U1274 (N_1274,N_974,N_523);
and U1275 (N_1275,In_1087,N_36);
nor U1276 (N_1276,N_991,In_777);
or U1277 (N_1277,In_1255,N_655);
or U1278 (N_1278,N_559,In_1738);
nand U1279 (N_1279,In_731,In_1565);
nor U1280 (N_1280,N_817,N_792);
nand U1281 (N_1281,N_24,In_1517);
or U1282 (N_1282,N_671,N_770);
or U1283 (N_1283,N_45,In_1551);
xnor U1284 (N_1284,N_626,In_394);
or U1285 (N_1285,In_1531,In_1318);
nor U1286 (N_1286,In_1801,In_1897);
nor U1287 (N_1287,N_800,N_939);
or U1288 (N_1288,N_597,N_709);
and U1289 (N_1289,N_101,N_125);
nand U1290 (N_1290,In_1247,N_18);
nor U1291 (N_1291,N_776,In_1762);
nor U1292 (N_1292,In_37,N_204);
and U1293 (N_1293,In_964,N_175);
nand U1294 (N_1294,In_1855,N_679);
nand U1295 (N_1295,N_621,N_508);
and U1296 (N_1296,In_1658,N_759);
nand U1297 (N_1297,N_730,In_578);
nand U1298 (N_1298,N_73,N_683);
nand U1299 (N_1299,N_743,N_972);
and U1300 (N_1300,N_982,N_922);
or U1301 (N_1301,In_64,In_651);
and U1302 (N_1302,N_789,N_984);
nor U1303 (N_1303,In_525,N_962);
or U1304 (N_1304,N_50,N_690);
xor U1305 (N_1305,In_1553,N_372);
or U1306 (N_1306,N_642,N_547);
nor U1307 (N_1307,In_1172,In_1775);
xnor U1308 (N_1308,In_1230,N_806);
or U1309 (N_1309,N_835,N_839);
nand U1310 (N_1310,N_966,N_511);
and U1311 (N_1311,In_1714,In_103);
or U1312 (N_1312,N_767,N_335);
xnor U1313 (N_1313,In_249,N_539);
and U1314 (N_1314,N_907,N_713);
nor U1315 (N_1315,In_874,N_648);
or U1316 (N_1316,N_594,In_365);
nand U1317 (N_1317,N_577,N_616);
nand U1318 (N_1318,In_423,In_898);
or U1319 (N_1319,N_801,In_1735);
and U1320 (N_1320,N_707,N_680);
or U1321 (N_1321,In_1445,In_206);
nor U1322 (N_1322,N_761,In_542);
and U1323 (N_1323,N_660,N_382);
xnor U1324 (N_1324,N_128,In_892);
nor U1325 (N_1325,N_112,N_802);
and U1326 (N_1326,N_609,N_970);
nor U1327 (N_1327,N_630,In_1012);
and U1328 (N_1328,N_864,N_950);
or U1329 (N_1329,N_892,N_27);
nand U1330 (N_1330,In_797,N_548);
or U1331 (N_1331,In_99,N_205);
xor U1332 (N_1332,N_512,N_785);
or U1333 (N_1333,N_694,N_979);
or U1334 (N_1334,N_445,N_954);
or U1335 (N_1335,In_877,In_1972);
or U1336 (N_1336,N_836,In_53);
and U1337 (N_1337,In_165,N_575);
or U1338 (N_1338,In_227,In_1042);
nor U1339 (N_1339,In_58,In_1363);
or U1340 (N_1340,In_1269,N_531);
or U1341 (N_1341,N_891,In_1057);
or U1342 (N_1342,In_1290,In_1467);
nand U1343 (N_1343,N_332,In_50);
nand U1344 (N_1344,In_1822,N_673);
nand U1345 (N_1345,N_403,N_712);
nand U1346 (N_1346,In_957,In_192);
nor U1347 (N_1347,N_902,N_717);
nor U1348 (N_1348,In_1475,N_505);
nand U1349 (N_1349,N_924,In_1080);
xor U1350 (N_1350,N_992,N_580);
or U1351 (N_1351,In_1496,N_790);
and U1352 (N_1352,In_1107,N_670);
xor U1353 (N_1353,N_352,N_944);
nor U1354 (N_1354,N_467,N_384);
xnor U1355 (N_1355,N_245,N_788);
nand U1356 (N_1356,N_699,N_65);
or U1357 (N_1357,In_455,N_681);
nor U1358 (N_1358,N_764,N_564);
or U1359 (N_1359,In_429,In_1912);
or U1360 (N_1360,N_719,N_326);
and U1361 (N_1361,N_889,N_832);
nand U1362 (N_1362,N_920,In_411);
and U1363 (N_1363,In_1367,N_841);
and U1364 (N_1364,In_678,N_557);
and U1365 (N_1365,In_1101,N_409);
and U1366 (N_1366,N_535,N_997);
nor U1367 (N_1367,N_113,In_112);
nand U1368 (N_1368,In_1928,N_203);
and U1369 (N_1369,N_482,N_928);
nand U1370 (N_1370,In_884,In_693);
nor U1371 (N_1371,N_831,N_513);
and U1372 (N_1372,N_139,In_188);
or U1373 (N_1373,N_754,In_1391);
or U1374 (N_1374,N_744,N_904);
and U1375 (N_1375,In_1750,N_781);
nor U1376 (N_1376,N_757,In_1579);
nand U1377 (N_1377,N_589,N_583);
or U1378 (N_1378,N_133,N_628);
nand U1379 (N_1379,In_8,N_834);
nand U1380 (N_1380,In_882,N_803);
nor U1381 (N_1381,N_857,In_1819);
and U1382 (N_1382,N_815,N_26);
nor U1383 (N_1383,In_465,N_816);
nor U1384 (N_1384,In_373,In_126);
nor U1385 (N_1385,N_983,N_15);
nor U1386 (N_1386,N_334,N_996);
and U1387 (N_1387,N_877,N_827);
nand U1388 (N_1388,N_615,N_685);
nor U1389 (N_1389,N_851,N_645);
nor U1390 (N_1390,N_724,N_682);
nor U1391 (N_1391,In_752,N_795);
nand U1392 (N_1392,N_777,N_567);
nor U1393 (N_1393,In_1260,In_1736);
and U1394 (N_1394,N_661,N_160);
nand U1395 (N_1395,N_784,N_884);
and U1396 (N_1396,N_64,N_443);
or U1397 (N_1397,In_1598,N_923);
and U1398 (N_1398,N_650,N_611);
nor U1399 (N_1399,N_504,In_512);
and U1400 (N_1400,N_612,N_960);
nand U1401 (N_1401,In_1430,N_59);
xor U1402 (N_1402,In_478,In_219);
nor U1403 (N_1403,N_464,N_975);
or U1404 (N_1404,N_168,N_968);
nor U1405 (N_1405,N_957,N_880);
and U1406 (N_1406,In_1739,N_658);
nand U1407 (N_1407,In_1228,N_765);
xor U1408 (N_1408,In_168,N_696);
and U1409 (N_1409,N_883,N_885);
or U1410 (N_1410,N_480,N_129);
and U1411 (N_1411,In_1117,N_783);
xnor U1412 (N_1412,N_748,N_400);
nor U1413 (N_1413,N_720,N_871);
and U1414 (N_1414,N_927,N_519);
and U1415 (N_1415,N_852,N_246);
nor U1416 (N_1416,N_501,N_844);
xnor U1417 (N_1417,N_829,N_275);
nand U1418 (N_1418,In_1655,In_1780);
nand U1419 (N_1419,N_775,N_731);
and U1420 (N_1420,In_1381,N_805);
nor U1421 (N_1421,In_1130,In_123);
nand U1422 (N_1422,In_980,N_669);
nand U1423 (N_1423,In_1165,N_909);
xnor U1424 (N_1424,N_808,In_1879);
nand U1425 (N_1425,N_198,N_810);
nor U1426 (N_1426,In_1968,N_804);
and U1427 (N_1427,N_987,N_514);
and U1428 (N_1428,N_937,In_183);
nand U1429 (N_1429,N_87,In_1934);
nand U1430 (N_1430,N_522,N_142);
nand U1431 (N_1431,In_529,In_229);
nor U1432 (N_1432,N_582,In_19);
nor U1433 (N_1433,In_482,N_747);
nand U1434 (N_1434,N_46,N_541);
or U1435 (N_1435,In_1271,N_338);
nor U1436 (N_1436,N_704,N_837);
and U1437 (N_1437,In_1836,In_810);
nand U1438 (N_1438,N_965,In_51);
xor U1439 (N_1439,N_627,N_666);
xnor U1440 (N_1440,N_607,N_935);
nor U1441 (N_1441,N_868,N_665);
or U1442 (N_1442,N_786,In_1717);
or U1443 (N_1443,In_938,In_1534);
or U1444 (N_1444,N_226,N_524);
nor U1445 (N_1445,N_995,N_895);
nand U1446 (N_1446,In_953,In_925);
or U1447 (N_1447,N_869,N_729);
nand U1448 (N_1448,N_625,In_1866);
and U1449 (N_1449,In_850,N_449);
nor U1450 (N_1450,In_591,N_921);
or U1451 (N_1451,N_192,N_819);
nor U1452 (N_1452,N_930,N_716);
and U1453 (N_1453,In_204,N_824);
or U1454 (N_1454,In_1078,N_407);
and U1455 (N_1455,In_539,N_21);
xor U1456 (N_1456,N_339,In_1504);
and U1457 (N_1457,N_536,In_988);
nor U1458 (N_1458,N_961,N_971);
nor U1459 (N_1459,N_762,In_527);
xor U1460 (N_1460,N_733,N_725);
or U1461 (N_1461,N_585,N_796);
and U1462 (N_1462,N_502,N_778);
or U1463 (N_1463,N_587,N_662);
nand U1464 (N_1464,N_870,N_848);
or U1465 (N_1465,In_685,N_503);
nand U1466 (N_1466,N_590,N_527);
and U1467 (N_1467,N_377,In_1987);
and U1468 (N_1468,N_416,N_917);
nand U1469 (N_1469,In_393,N_737);
and U1470 (N_1470,N_517,N_544);
and U1471 (N_1471,In_208,In_696);
nand U1472 (N_1472,N_689,N_701);
or U1473 (N_1473,N_180,In_368);
or U1474 (N_1474,In_637,In_1313);
nand U1475 (N_1475,N_568,N_768);
or U1476 (N_1476,N_915,N_749);
and U1477 (N_1477,In_1854,In_84);
nor U1478 (N_1478,N_629,In_1929);
nand U1479 (N_1479,N_646,N_631);
or U1480 (N_1480,In_1189,In_1623);
and U1481 (N_1481,N_787,N_252);
nor U1482 (N_1482,N_649,N_152);
nand U1483 (N_1483,N_124,N_888);
nor U1484 (N_1484,In_1004,In_1408);
nor U1485 (N_1485,N_952,In_1361);
xor U1486 (N_1486,N_854,In_1851);
or U1487 (N_1487,N_740,N_846);
nand U1488 (N_1488,N_506,N_843);
nor U1489 (N_1489,N_833,In_1562);
nand U1490 (N_1490,N_945,N_574);
xnor U1491 (N_1491,N_435,N_428);
nor U1492 (N_1492,N_828,N_380);
or U1493 (N_1493,N_66,N_617);
nor U1494 (N_1494,N_932,N_488);
nand U1495 (N_1495,In_788,In_1395);
xor U1496 (N_1496,In_869,In_254);
or U1497 (N_1497,N_362,N_691);
and U1498 (N_1498,In_62,N_692);
nand U1499 (N_1499,In_1895,N_444);
and U1500 (N_1500,N_1358,N_1224);
nor U1501 (N_1501,N_1302,N_1321);
xnor U1502 (N_1502,N_1202,N_1460);
or U1503 (N_1503,N_1424,N_1118);
or U1504 (N_1504,N_1024,N_1493);
xnor U1505 (N_1505,N_1407,N_1351);
or U1506 (N_1506,N_1313,N_1296);
nor U1507 (N_1507,N_1100,N_1331);
nor U1508 (N_1508,N_1199,N_1242);
and U1509 (N_1509,N_1219,N_1171);
and U1510 (N_1510,N_1239,N_1338);
or U1511 (N_1511,N_1377,N_1444);
nor U1512 (N_1512,N_1379,N_1099);
or U1513 (N_1513,N_1165,N_1029);
nor U1514 (N_1514,N_1131,N_1163);
nor U1515 (N_1515,N_1426,N_1300);
and U1516 (N_1516,N_1402,N_1413);
and U1517 (N_1517,N_1474,N_1448);
nand U1518 (N_1518,N_1181,N_1012);
and U1519 (N_1519,N_1164,N_1457);
or U1520 (N_1520,N_1294,N_1280);
nand U1521 (N_1521,N_1340,N_1422);
or U1522 (N_1522,N_1499,N_1039);
nand U1523 (N_1523,N_1014,N_1274);
nand U1524 (N_1524,N_1049,N_1222);
nand U1525 (N_1525,N_1465,N_1106);
or U1526 (N_1526,N_1263,N_1365);
and U1527 (N_1527,N_1206,N_1341);
nand U1528 (N_1528,N_1094,N_1185);
nor U1529 (N_1529,N_1030,N_1478);
nor U1530 (N_1530,N_1277,N_1088);
or U1531 (N_1531,N_1031,N_1308);
nor U1532 (N_1532,N_1125,N_1211);
nand U1533 (N_1533,N_1393,N_1168);
nand U1534 (N_1534,N_1028,N_1266);
or U1535 (N_1535,N_1287,N_1160);
or U1536 (N_1536,N_1273,N_1364);
nor U1537 (N_1537,N_1354,N_1489);
or U1538 (N_1538,N_1084,N_1495);
or U1539 (N_1539,N_1447,N_1285);
nor U1540 (N_1540,N_1357,N_1490);
nand U1541 (N_1541,N_1371,N_1486);
and U1542 (N_1542,N_1262,N_1021);
xor U1543 (N_1543,N_1240,N_1394);
and U1544 (N_1544,N_1214,N_1392);
or U1545 (N_1545,N_1268,N_1190);
or U1546 (N_1546,N_1347,N_1055);
or U1547 (N_1547,N_1337,N_1419);
and U1548 (N_1548,N_1256,N_1400);
nand U1549 (N_1549,N_1389,N_1405);
and U1550 (N_1550,N_1417,N_1150);
or U1551 (N_1551,N_1298,N_1162);
xor U1552 (N_1552,N_1312,N_1013);
and U1553 (N_1553,N_1025,N_1428);
or U1554 (N_1554,N_1090,N_1497);
nor U1555 (N_1555,N_1235,N_1065);
xnor U1556 (N_1556,N_1144,N_1310);
or U1557 (N_1557,N_1323,N_1397);
or U1558 (N_1558,N_1140,N_1368);
nand U1559 (N_1559,N_1427,N_1480);
nand U1560 (N_1560,N_1068,N_1335);
and U1561 (N_1561,N_1059,N_1184);
nor U1562 (N_1562,N_1261,N_1492);
xor U1563 (N_1563,N_1311,N_1267);
xnor U1564 (N_1564,N_1126,N_1195);
nor U1565 (N_1565,N_1324,N_1454);
nor U1566 (N_1566,N_1384,N_1320);
nand U1567 (N_1567,N_1194,N_1343);
nor U1568 (N_1568,N_1336,N_1141);
nor U1569 (N_1569,N_1241,N_1291);
xnor U1570 (N_1570,N_1498,N_1443);
nor U1571 (N_1571,N_1197,N_1083);
and U1572 (N_1572,N_1119,N_1103);
nor U1573 (N_1573,N_1155,N_1440);
and U1574 (N_1574,N_1390,N_1376);
nand U1575 (N_1575,N_1076,N_1123);
nor U1576 (N_1576,N_1200,N_1381);
nor U1577 (N_1577,N_1309,N_1130);
nor U1578 (N_1578,N_1000,N_1369);
or U1579 (N_1579,N_1432,N_1189);
and U1580 (N_1580,N_1134,N_1361);
and U1581 (N_1581,N_1048,N_1359);
nor U1582 (N_1582,N_1270,N_1468);
nand U1583 (N_1583,N_1382,N_1481);
nor U1584 (N_1584,N_1105,N_1036);
and U1585 (N_1585,N_1091,N_1179);
nand U1586 (N_1586,N_1386,N_1108);
nand U1587 (N_1587,N_1362,N_1040);
xor U1588 (N_1588,N_1353,N_1412);
nand U1589 (N_1589,N_1207,N_1257);
nor U1590 (N_1590,N_1018,N_1439);
nor U1591 (N_1591,N_1002,N_1325);
nand U1592 (N_1592,N_1205,N_1079);
nand U1593 (N_1593,N_1062,N_1295);
xor U1594 (N_1594,N_1398,N_1132);
nand U1595 (N_1595,N_1374,N_1104);
or U1596 (N_1596,N_1322,N_1438);
nand U1597 (N_1597,N_1366,N_1097);
nand U1598 (N_1598,N_1290,N_1360);
nand U1599 (N_1599,N_1033,N_1234);
or U1600 (N_1600,N_1057,N_1107);
or U1601 (N_1601,N_1434,N_1334);
or U1602 (N_1602,N_1067,N_1078);
and U1603 (N_1603,N_1225,N_1327);
and U1604 (N_1604,N_1201,N_1149);
and U1605 (N_1605,N_1232,N_1293);
or U1606 (N_1606,N_1198,N_1248);
nor U1607 (N_1607,N_1192,N_1053);
and U1608 (N_1608,N_1373,N_1026);
xnor U1609 (N_1609,N_1109,N_1175);
nor U1610 (N_1610,N_1349,N_1350);
nor U1611 (N_1611,N_1469,N_1128);
xnor U1612 (N_1612,N_1072,N_1186);
and U1613 (N_1613,N_1082,N_1156);
nor U1614 (N_1614,N_1410,N_1370);
and U1615 (N_1615,N_1339,N_1281);
nor U1616 (N_1616,N_1375,N_1102);
and U1617 (N_1617,N_1135,N_1254);
nand U1618 (N_1618,N_1395,N_1085);
or U1619 (N_1619,N_1152,N_1001);
or U1620 (N_1620,N_1045,N_1080);
or U1621 (N_1621,N_1101,N_1196);
or U1622 (N_1622,N_1050,N_1210);
and U1623 (N_1623,N_1473,N_1114);
or U1624 (N_1624,N_1077,N_1292);
and U1625 (N_1625,N_1213,N_1462);
or U1626 (N_1626,N_1483,N_1110);
nor U1627 (N_1627,N_1143,N_1208);
nand U1628 (N_1628,N_1064,N_1403);
or U1629 (N_1629,N_1271,N_1008);
or U1630 (N_1630,N_1463,N_1459);
xor U1631 (N_1631,N_1147,N_1329);
nor U1632 (N_1632,N_1431,N_1051);
or U1633 (N_1633,N_1496,N_1279);
and U1634 (N_1634,N_1276,N_1414);
and U1635 (N_1635,N_1148,N_1346);
nand U1636 (N_1636,N_1236,N_1467);
xnor U1637 (N_1637,N_1316,N_1095);
nor U1638 (N_1638,N_1058,N_1301);
nand U1639 (N_1639,N_1066,N_1124);
nand U1640 (N_1640,N_1054,N_1151);
nor U1641 (N_1641,N_1265,N_1117);
and U1642 (N_1642,N_1133,N_1178);
and U1643 (N_1643,N_1042,N_1482);
nand U1644 (N_1644,N_1437,N_1435);
or U1645 (N_1645,N_1433,N_1145);
nand U1646 (N_1646,N_1015,N_1278);
nand U1647 (N_1647,N_1352,N_1034);
or U1648 (N_1648,N_1476,N_1245);
nor U1649 (N_1649,N_1446,N_1136);
and U1650 (N_1650,N_1157,N_1415);
xor U1651 (N_1651,N_1250,N_1429);
and U1652 (N_1652,N_1430,N_1212);
and U1653 (N_1653,N_1345,N_1093);
xnor U1654 (N_1654,N_1069,N_1247);
nand U1655 (N_1655,N_1442,N_1063);
or U1656 (N_1656,N_1170,N_1282);
or U1657 (N_1657,N_1022,N_1218);
and U1658 (N_1658,N_1319,N_1041);
or U1659 (N_1659,N_1075,N_1204);
xnor U1660 (N_1660,N_1342,N_1356);
and U1661 (N_1661,N_1061,N_1203);
or U1662 (N_1662,N_1477,N_1056);
xnor U1663 (N_1663,N_1304,N_1318);
nand U1664 (N_1664,N_1191,N_1209);
or U1665 (N_1665,N_1344,N_1307);
or U1666 (N_1666,N_1387,N_1260);
xnor U1667 (N_1667,N_1215,N_1264);
nor U1668 (N_1668,N_1193,N_1038);
nand U1669 (N_1669,N_1120,N_1073);
or U1670 (N_1670,N_1449,N_1409);
or U1671 (N_1671,N_1005,N_1253);
xnor U1672 (N_1672,N_1116,N_1009);
and U1673 (N_1673,N_1081,N_1315);
nor U1674 (N_1674,N_1399,N_1037);
or U1675 (N_1675,N_1139,N_1098);
and U1676 (N_1676,N_1173,N_1086);
and U1677 (N_1677,N_1408,N_1305);
xnor U1678 (N_1678,N_1418,N_1158);
or U1679 (N_1679,N_1188,N_1217);
nor U1680 (N_1680,N_1472,N_1159);
or U1681 (N_1681,N_1047,N_1003);
or U1682 (N_1682,N_1032,N_1092);
and U1683 (N_1683,N_1259,N_1111);
or U1684 (N_1684,N_1220,N_1404);
xnor U1685 (N_1685,N_1044,N_1421);
nor U1686 (N_1686,N_1233,N_1378);
nand U1687 (N_1687,N_1436,N_1046);
and U1688 (N_1688,N_1238,N_1016);
or U1689 (N_1689,N_1471,N_1406);
xor U1690 (N_1690,N_1450,N_1174);
or U1691 (N_1691,N_1231,N_1401);
nand U1692 (N_1692,N_1416,N_1303);
xor U1693 (N_1693,N_1187,N_1491);
nand U1694 (N_1694,N_1183,N_1020);
nand U1695 (N_1695,N_1228,N_1035);
and U1696 (N_1696,N_1122,N_1355);
or U1697 (N_1697,N_1461,N_1367);
nand U1698 (N_1698,N_1146,N_1494);
or U1699 (N_1699,N_1441,N_1153);
nor U1700 (N_1700,N_1297,N_1385);
nand U1701 (N_1701,N_1328,N_1363);
or U1702 (N_1702,N_1172,N_1138);
xnor U1703 (N_1703,N_1475,N_1216);
nand U1704 (N_1704,N_1167,N_1019);
and U1705 (N_1705,N_1288,N_1246);
nor U1706 (N_1706,N_1388,N_1142);
nand U1707 (N_1707,N_1348,N_1176);
nor U1708 (N_1708,N_1177,N_1221);
nor U1709 (N_1709,N_1237,N_1284);
nor U1710 (N_1710,N_1226,N_1479);
nand U1711 (N_1711,N_1017,N_1330);
xnor U1712 (N_1712,N_1314,N_1027);
and U1713 (N_1713,N_1485,N_1007);
xor U1714 (N_1714,N_1396,N_1023);
nand U1715 (N_1715,N_1372,N_1089);
xor U1716 (N_1716,N_1010,N_1252);
or U1717 (N_1717,N_1458,N_1052);
xor U1718 (N_1718,N_1333,N_1243);
or U1719 (N_1719,N_1169,N_1466);
nor U1720 (N_1720,N_1425,N_1289);
or U1721 (N_1721,N_1182,N_1154);
or U1722 (N_1722,N_1113,N_1451);
nand U1723 (N_1723,N_1456,N_1258);
nor U1724 (N_1724,N_1223,N_1137);
nor U1725 (N_1725,N_1380,N_1011);
nand U1726 (N_1726,N_1251,N_1121);
nor U1727 (N_1727,N_1161,N_1071);
nand U1728 (N_1728,N_1249,N_1269);
or U1729 (N_1729,N_1074,N_1115);
or U1730 (N_1730,N_1455,N_1487);
xor U1731 (N_1731,N_1420,N_1229);
or U1732 (N_1732,N_1230,N_1332);
nor U1733 (N_1733,N_1070,N_1383);
nor U1734 (N_1734,N_1423,N_1283);
nor U1735 (N_1735,N_1112,N_1453);
nor U1736 (N_1736,N_1306,N_1470);
xnor U1737 (N_1737,N_1180,N_1166);
and U1738 (N_1738,N_1488,N_1129);
nor U1739 (N_1739,N_1272,N_1060);
or U1740 (N_1740,N_1275,N_1484);
and U1741 (N_1741,N_1244,N_1286);
nor U1742 (N_1742,N_1096,N_1004);
and U1743 (N_1743,N_1255,N_1043);
nand U1744 (N_1744,N_1006,N_1445);
nand U1745 (N_1745,N_1299,N_1464);
or U1746 (N_1746,N_1391,N_1411);
nand U1747 (N_1747,N_1317,N_1087);
nor U1748 (N_1748,N_1127,N_1452);
or U1749 (N_1749,N_1227,N_1326);
nand U1750 (N_1750,N_1471,N_1343);
or U1751 (N_1751,N_1425,N_1178);
nand U1752 (N_1752,N_1443,N_1279);
or U1753 (N_1753,N_1472,N_1084);
and U1754 (N_1754,N_1483,N_1357);
and U1755 (N_1755,N_1282,N_1381);
nor U1756 (N_1756,N_1499,N_1395);
nor U1757 (N_1757,N_1135,N_1430);
nor U1758 (N_1758,N_1239,N_1108);
and U1759 (N_1759,N_1179,N_1137);
or U1760 (N_1760,N_1021,N_1325);
nand U1761 (N_1761,N_1431,N_1377);
nor U1762 (N_1762,N_1469,N_1313);
nand U1763 (N_1763,N_1085,N_1422);
nor U1764 (N_1764,N_1440,N_1148);
nor U1765 (N_1765,N_1073,N_1227);
nand U1766 (N_1766,N_1478,N_1222);
and U1767 (N_1767,N_1317,N_1150);
nand U1768 (N_1768,N_1234,N_1271);
or U1769 (N_1769,N_1166,N_1099);
xor U1770 (N_1770,N_1465,N_1363);
nor U1771 (N_1771,N_1458,N_1492);
nor U1772 (N_1772,N_1201,N_1380);
nand U1773 (N_1773,N_1019,N_1023);
and U1774 (N_1774,N_1483,N_1045);
nor U1775 (N_1775,N_1278,N_1002);
or U1776 (N_1776,N_1154,N_1103);
nand U1777 (N_1777,N_1096,N_1116);
or U1778 (N_1778,N_1439,N_1020);
or U1779 (N_1779,N_1038,N_1080);
or U1780 (N_1780,N_1012,N_1268);
nand U1781 (N_1781,N_1023,N_1445);
and U1782 (N_1782,N_1217,N_1030);
nand U1783 (N_1783,N_1107,N_1489);
or U1784 (N_1784,N_1101,N_1217);
or U1785 (N_1785,N_1303,N_1107);
nand U1786 (N_1786,N_1183,N_1215);
xnor U1787 (N_1787,N_1439,N_1075);
or U1788 (N_1788,N_1159,N_1264);
nor U1789 (N_1789,N_1182,N_1424);
and U1790 (N_1790,N_1424,N_1098);
and U1791 (N_1791,N_1480,N_1241);
and U1792 (N_1792,N_1153,N_1077);
and U1793 (N_1793,N_1482,N_1280);
xnor U1794 (N_1794,N_1466,N_1473);
nor U1795 (N_1795,N_1271,N_1031);
nor U1796 (N_1796,N_1178,N_1063);
or U1797 (N_1797,N_1175,N_1124);
nor U1798 (N_1798,N_1052,N_1017);
and U1799 (N_1799,N_1025,N_1078);
nand U1800 (N_1800,N_1158,N_1479);
and U1801 (N_1801,N_1205,N_1130);
or U1802 (N_1802,N_1488,N_1457);
or U1803 (N_1803,N_1378,N_1422);
nand U1804 (N_1804,N_1284,N_1179);
and U1805 (N_1805,N_1353,N_1354);
nand U1806 (N_1806,N_1262,N_1089);
or U1807 (N_1807,N_1464,N_1011);
nand U1808 (N_1808,N_1463,N_1430);
or U1809 (N_1809,N_1430,N_1194);
nor U1810 (N_1810,N_1082,N_1110);
or U1811 (N_1811,N_1317,N_1421);
nor U1812 (N_1812,N_1042,N_1316);
or U1813 (N_1813,N_1090,N_1324);
nand U1814 (N_1814,N_1105,N_1035);
and U1815 (N_1815,N_1223,N_1316);
xnor U1816 (N_1816,N_1331,N_1284);
and U1817 (N_1817,N_1420,N_1456);
nor U1818 (N_1818,N_1371,N_1268);
and U1819 (N_1819,N_1499,N_1016);
and U1820 (N_1820,N_1297,N_1259);
and U1821 (N_1821,N_1417,N_1180);
or U1822 (N_1822,N_1236,N_1310);
xor U1823 (N_1823,N_1026,N_1378);
xnor U1824 (N_1824,N_1315,N_1291);
nor U1825 (N_1825,N_1378,N_1358);
or U1826 (N_1826,N_1419,N_1486);
nand U1827 (N_1827,N_1252,N_1277);
xnor U1828 (N_1828,N_1228,N_1347);
nor U1829 (N_1829,N_1015,N_1018);
xnor U1830 (N_1830,N_1333,N_1011);
nor U1831 (N_1831,N_1278,N_1321);
xor U1832 (N_1832,N_1093,N_1354);
nand U1833 (N_1833,N_1143,N_1431);
nand U1834 (N_1834,N_1199,N_1297);
nand U1835 (N_1835,N_1212,N_1392);
or U1836 (N_1836,N_1296,N_1366);
xnor U1837 (N_1837,N_1205,N_1486);
or U1838 (N_1838,N_1220,N_1411);
xor U1839 (N_1839,N_1457,N_1235);
xnor U1840 (N_1840,N_1334,N_1357);
nor U1841 (N_1841,N_1171,N_1410);
or U1842 (N_1842,N_1172,N_1170);
xor U1843 (N_1843,N_1123,N_1374);
xor U1844 (N_1844,N_1009,N_1344);
nand U1845 (N_1845,N_1460,N_1010);
or U1846 (N_1846,N_1391,N_1379);
nor U1847 (N_1847,N_1167,N_1452);
and U1848 (N_1848,N_1221,N_1017);
nand U1849 (N_1849,N_1475,N_1250);
and U1850 (N_1850,N_1414,N_1309);
or U1851 (N_1851,N_1467,N_1312);
or U1852 (N_1852,N_1080,N_1026);
nand U1853 (N_1853,N_1357,N_1105);
and U1854 (N_1854,N_1361,N_1383);
and U1855 (N_1855,N_1196,N_1225);
nand U1856 (N_1856,N_1177,N_1383);
nor U1857 (N_1857,N_1439,N_1281);
or U1858 (N_1858,N_1019,N_1498);
nand U1859 (N_1859,N_1001,N_1000);
or U1860 (N_1860,N_1029,N_1175);
and U1861 (N_1861,N_1217,N_1296);
nor U1862 (N_1862,N_1461,N_1097);
nor U1863 (N_1863,N_1048,N_1446);
and U1864 (N_1864,N_1292,N_1113);
and U1865 (N_1865,N_1269,N_1001);
and U1866 (N_1866,N_1001,N_1242);
nand U1867 (N_1867,N_1016,N_1284);
and U1868 (N_1868,N_1265,N_1338);
nand U1869 (N_1869,N_1355,N_1437);
or U1870 (N_1870,N_1284,N_1400);
nand U1871 (N_1871,N_1144,N_1040);
nor U1872 (N_1872,N_1096,N_1140);
nor U1873 (N_1873,N_1207,N_1234);
nand U1874 (N_1874,N_1326,N_1060);
nand U1875 (N_1875,N_1164,N_1265);
nand U1876 (N_1876,N_1049,N_1180);
xnor U1877 (N_1877,N_1439,N_1151);
and U1878 (N_1878,N_1474,N_1334);
and U1879 (N_1879,N_1238,N_1173);
nor U1880 (N_1880,N_1300,N_1203);
nand U1881 (N_1881,N_1199,N_1266);
nand U1882 (N_1882,N_1315,N_1244);
or U1883 (N_1883,N_1024,N_1283);
nand U1884 (N_1884,N_1293,N_1111);
nand U1885 (N_1885,N_1387,N_1218);
or U1886 (N_1886,N_1082,N_1095);
nor U1887 (N_1887,N_1215,N_1477);
nor U1888 (N_1888,N_1081,N_1017);
and U1889 (N_1889,N_1121,N_1473);
nand U1890 (N_1890,N_1287,N_1342);
and U1891 (N_1891,N_1220,N_1259);
and U1892 (N_1892,N_1015,N_1098);
nand U1893 (N_1893,N_1231,N_1233);
or U1894 (N_1894,N_1100,N_1364);
and U1895 (N_1895,N_1434,N_1065);
or U1896 (N_1896,N_1247,N_1287);
or U1897 (N_1897,N_1297,N_1150);
and U1898 (N_1898,N_1191,N_1001);
nor U1899 (N_1899,N_1174,N_1421);
nand U1900 (N_1900,N_1469,N_1247);
or U1901 (N_1901,N_1189,N_1470);
nor U1902 (N_1902,N_1000,N_1169);
nor U1903 (N_1903,N_1121,N_1031);
and U1904 (N_1904,N_1477,N_1172);
nor U1905 (N_1905,N_1444,N_1226);
nand U1906 (N_1906,N_1089,N_1303);
and U1907 (N_1907,N_1263,N_1069);
or U1908 (N_1908,N_1269,N_1152);
nand U1909 (N_1909,N_1249,N_1069);
and U1910 (N_1910,N_1076,N_1115);
nand U1911 (N_1911,N_1117,N_1350);
and U1912 (N_1912,N_1158,N_1276);
nand U1913 (N_1913,N_1223,N_1098);
nand U1914 (N_1914,N_1262,N_1020);
and U1915 (N_1915,N_1378,N_1304);
nor U1916 (N_1916,N_1089,N_1020);
nand U1917 (N_1917,N_1441,N_1132);
nor U1918 (N_1918,N_1286,N_1453);
or U1919 (N_1919,N_1384,N_1100);
nand U1920 (N_1920,N_1243,N_1377);
and U1921 (N_1921,N_1269,N_1317);
nor U1922 (N_1922,N_1426,N_1393);
nor U1923 (N_1923,N_1110,N_1175);
and U1924 (N_1924,N_1012,N_1204);
or U1925 (N_1925,N_1454,N_1108);
nor U1926 (N_1926,N_1426,N_1476);
nand U1927 (N_1927,N_1331,N_1406);
xor U1928 (N_1928,N_1366,N_1412);
nor U1929 (N_1929,N_1484,N_1025);
xnor U1930 (N_1930,N_1418,N_1424);
nand U1931 (N_1931,N_1418,N_1145);
or U1932 (N_1932,N_1280,N_1249);
and U1933 (N_1933,N_1061,N_1498);
or U1934 (N_1934,N_1444,N_1374);
or U1935 (N_1935,N_1316,N_1436);
nor U1936 (N_1936,N_1203,N_1181);
nand U1937 (N_1937,N_1428,N_1061);
xnor U1938 (N_1938,N_1484,N_1016);
or U1939 (N_1939,N_1470,N_1280);
nand U1940 (N_1940,N_1018,N_1250);
and U1941 (N_1941,N_1093,N_1411);
or U1942 (N_1942,N_1190,N_1242);
xnor U1943 (N_1943,N_1120,N_1026);
nor U1944 (N_1944,N_1449,N_1313);
or U1945 (N_1945,N_1144,N_1439);
and U1946 (N_1946,N_1454,N_1457);
nand U1947 (N_1947,N_1229,N_1093);
xnor U1948 (N_1948,N_1055,N_1126);
or U1949 (N_1949,N_1020,N_1152);
and U1950 (N_1950,N_1325,N_1034);
or U1951 (N_1951,N_1407,N_1339);
or U1952 (N_1952,N_1107,N_1462);
or U1953 (N_1953,N_1105,N_1084);
xor U1954 (N_1954,N_1413,N_1483);
nor U1955 (N_1955,N_1067,N_1364);
xnor U1956 (N_1956,N_1280,N_1237);
and U1957 (N_1957,N_1033,N_1093);
or U1958 (N_1958,N_1420,N_1166);
nand U1959 (N_1959,N_1204,N_1230);
nor U1960 (N_1960,N_1201,N_1437);
nand U1961 (N_1961,N_1295,N_1234);
nand U1962 (N_1962,N_1089,N_1404);
xor U1963 (N_1963,N_1412,N_1380);
or U1964 (N_1964,N_1222,N_1437);
nand U1965 (N_1965,N_1378,N_1398);
nor U1966 (N_1966,N_1322,N_1084);
nor U1967 (N_1967,N_1053,N_1448);
or U1968 (N_1968,N_1023,N_1479);
or U1969 (N_1969,N_1392,N_1383);
and U1970 (N_1970,N_1214,N_1470);
and U1971 (N_1971,N_1146,N_1359);
and U1972 (N_1972,N_1032,N_1360);
and U1973 (N_1973,N_1434,N_1148);
xor U1974 (N_1974,N_1194,N_1182);
nand U1975 (N_1975,N_1315,N_1111);
nor U1976 (N_1976,N_1071,N_1468);
or U1977 (N_1977,N_1177,N_1345);
and U1978 (N_1978,N_1339,N_1132);
nand U1979 (N_1979,N_1028,N_1000);
nand U1980 (N_1980,N_1424,N_1089);
and U1981 (N_1981,N_1040,N_1323);
nor U1982 (N_1982,N_1142,N_1170);
and U1983 (N_1983,N_1152,N_1431);
nor U1984 (N_1984,N_1436,N_1411);
nor U1985 (N_1985,N_1056,N_1356);
nor U1986 (N_1986,N_1494,N_1334);
nand U1987 (N_1987,N_1389,N_1237);
or U1988 (N_1988,N_1441,N_1238);
nor U1989 (N_1989,N_1368,N_1132);
or U1990 (N_1990,N_1062,N_1436);
or U1991 (N_1991,N_1129,N_1320);
nand U1992 (N_1992,N_1248,N_1225);
nor U1993 (N_1993,N_1146,N_1214);
xor U1994 (N_1994,N_1115,N_1428);
or U1995 (N_1995,N_1403,N_1184);
nor U1996 (N_1996,N_1184,N_1387);
and U1997 (N_1997,N_1319,N_1282);
nor U1998 (N_1998,N_1260,N_1466);
and U1999 (N_1999,N_1218,N_1312);
and U2000 (N_2000,N_1543,N_1777);
nor U2001 (N_2001,N_1998,N_1875);
nor U2002 (N_2002,N_1989,N_1546);
nor U2003 (N_2003,N_1613,N_1534);
or U2004 (N_2004,N_1908,N_1902);
nand U2005 (N_2005,N_1725,N_1655);
and U2006 (N_2006,N_1944,N_1909);
or U2007 (N_2007,N_1624,N_1775);
or U2008 (N_2008,N_1743,N_1644);
nor U2009 (N_2009,N_1979,N_1574);
nand U2010 (N_2010,N_1922,N_1951);
and U2011 (N_2011,N_1924,N_1699);
and U2012 (N_2012,N_1698,N_1940);
and U2013 (N_2013,N_1550,N_1763);
nand U2014 (N_2014,N_1586,N_1936);
and U2015 (N_2015,N_1567,N_1905);
or U2016 (N_2016,N_1693,N_1745);
nor U2017 (N_2017,N_1508,N_1617);
nor U2018 (N_2018,N_1893,N_1570);
nand U2019 (N_2019,N_1649,N_1781);
xor U2020 (N_2020,N_1672,N_1657);
nor U2021 (N_2021,N_1977,N_1600);
or U2022 (N_2022,N_1798,N_1929);
nor U2023 (N_2023,N_1872,N_1547);
and U2024 (N_2024,N_1500,N_1688);
and U2025 (N_2025,N_1641,N_1604);
or U2026 (N_2026,N_1642,N_1766);
or U2027 (N_2027,N_1884,N_1939);
nor U2028 (N_2028,N_1796,N_1726);
nor U2029 (N_2029,N_1588,N_1737);
or U2030 (N_2030,N_1591,N_1563);
nor U2031 (N_2031,N_1987,N_1815);
or U2032 (N_2032,N_1595,N_1530);
or U2033 (N_2033,N_1890,N_1622);
or U2034 (N_2034,N_1851,N_1732);
nor U2035 (N_2035,N_1943,N_1941);
and U2036 (N_2036,N_1728,N_1901);
or U2037 (N_2037,N_1632,N_1945);
or U2038 (N_2038,N_1599,N_1621);
nand U2039 (N_2039,N_1501,N_1637);
or U2040 (N_2040,N_1878,N_1587);
xor U2041 (N_2041,N_1866,N_1718);
nand U2042 (N_2042,N_1910,N_1799);
and U2043 (N_2043,N_1949,N_1981);
or U2044 (N_2044,N_1665,N_1895);
nor U2045 (N_2045,N_1551,N_1610);
and U2046 (N_2046,N_1876,N_1807);
and U2047 (N_2047,N_1727,N_1572);
nor U2048 (N_2048,N_1994,N_1933);
or U2049 (N_2049,N_1723,N_1707);
or U2050 (N_2050,N_1535,N_1660);
or U2051 (N_2051,N_1537,N_1602);
nand U2052 (N_2052,N_1605,N_1514);
nor U2053 (N_2053,N_1680,N_1823);
or U2054 (N_2054,N_1806,N_1555);
nor U2055 (N_2055,N_1831,N_1695);
nor U2056 (N_2056,N_1970,N_1957);
nand U2057 (N_2057,N_1790,N_1955);
xnor U2058 (N_2058,N_1579,N_1669);
nor U2059 (N_2059,N_1703,N_1717);
or U2060 (N_2060,N_1874,N_1923);
or U2061 (N_2061,N_1756,N_1846);
and U2062 (N_2062,N_1673,N_1962);
or U2063 (N_2063,N_1653,N_1540);
or U2064 (N_2064,N_1668,N_1697);
or U2065 (N_2065,N_1797,N_1837);
or U2066 (N_2066,N_1536,N_1864);
or U2067 (N_2067,N_1542,N_1930);
or U2068 (N_2068,N_1868,N_1964);
or U2069 (N_2069,N_1674,N_1640);
xnor U2070 (N_2070,N_1650,N_1681);
nand U2071 (N_2071,N_1808,N_1947);
nor U2072 (N_2072,N_1889,N_1504);
or U2073 (N_2073,N_1869,N_1883);
or U2074 (N_2074,N_1925,N_1912);
nor U2075 (N_2075,N_1871,N_1829);
and U2076 (N_2076,N_1577,N_1916);
or U2077 (N_2077,N_1854,N_1608);
nor U2078 (N_2078,N_1990,N_1708);
nand U2079 (N_2079,N_1956,N_1556);
and U2080 (N_2080,N_1541,N_1735);
nor U2081 (N_2081,N_1946,N_1772);
nand U2082 (N_2082,N_1842,N_1841);
nor U2083 (N_2083,N_1965,N_1954);
or U2084 (N_2084,N_1862,N_1667);
xnor U2085 (N_2085,N_1803,N_1716);
nand U2086 (N_2086,N_1670,N_1897);
xnor U2087 (N_2087,N_1611,N_1646);
or U2088 (N_2088,N_1553,N_1592);
or U2089 (N_2089,N_1704,N_1568);
and U2090 (N_2090,N_1515,N_1952);
nand U2091 (N_2091,N_1522,N_1830);
and U2092 (N_2092,N_1817,N_1742);
or U2093 (N_2093,N_1700,N_1762);
or U2094 (N_2094,N_1526,N_1926);
nand U2095 (N_2095,N_1792,N_1776);
nor U2096 (N_2096,N_1887,N_1788);
nand U2097 (N_2097,N_1532,N_1692);
and U2098 (N_2098,N_1658,N_1654);
and U2099 (N_2099,N_1919,N_1791);
xor U2100 (N_2100,N_1683,N_1983);
and U2101 (N_2101,N_1898,N_1696);
nor U2102 (N_2102,N_1710,N_1740);
xnor U2103 (N_2103,N_1517,N_1664);
and U2104 (N_2104,N_1639,N_1507);
nor U2105 (N_2105,N_1516,N_1715);
nand U2106 (N_2106,N_1519,N_1769);
or U2107 (N_2107,N_1991,N_1980);
nand U2108 (N_2108,N_1794,N_1523);
or U2109 (N_2109,N_1774,N_1531);
and U2110 (N_2110,N_1958,N_1731);
nand U2111 (N_2111,N_1953,N_1764);
or U2112 (N_2112,N_1719,N_1671);
xor U2113 (N_2113,N_1734,N_1684);
xor U2114 (N_2114,N_1961,N_1721);
nand U2115 (N_2115,N_1593,N_1963);
xnor U2116 (N_2116,N_1513,N_1984);
nor U2117 (N_2117,N_1896,N_1565);
xnor U2118 (N_2118,N_1720,N_1822);
or U2119 (N_2119,N_1971,N_1659);
nand U2120 (N_2120,N_1583,N_1818);
xor U2121 (N_2121,N_1966,N_1877);
nor U2122 (N_2122,N_1638,N_1629);
nand U2123 (N_2123,N_1913,N_1960);
nand U2124 (N_2124,N_1510,N_1575);
nand U2125 (N_2125,N_1741,N_1627);
nor U2126 (N_2126,N_1571,N_1856);
and U2127 (N_2127,N_1948,N_1882);
or U2128 (N_2128,N_1757,N_1739);
or U2129 (N_2129,N_1607,N_1789);
nor U2130 (N_2130,N_1663,N_1705);
nor U2131 (N_2131,N_1675,N_1503);
and U2132 (N_2132,N_1904,N_1761);
and U2133 (N_2133,N_1906,N_1937);
nand U2134 (N_2134,N_1770,N_1651);
and U2135 (N_2135,N_1618,N_1678);
nand U2136 (N_2136,N_1524,N_1558);
or U2137 (N_2137,N_1580,N_1623);
nand U2138 (N_2138,N_1748,N_1528);
and U2139 (N_2139,N_1722,N_1691);
and U2140 (N_2140,N_1746,N_1560);
nor U2141 (N_2141,N_1753,N_1578);
or U2142 (N_2142,N_1601,N_1802);
nand U2143 (N_2143,N_1589,N_1879);
or U2144 (N_2144,N_1927,N_1931);
and U2145 (N_2145,N_1685,N_1816);
and U2146 (N_2146,N_1917,N_1934);
nor U2147 (N_2147,N_1986,N_1648);
or U2148 (N_2148,N_1950,N_1942);
nand U2149 (N_2149,N_1967,N_1714);
xnor U2150 (N_2150,N_1838,N_1525);
nor U2151 (N_2151,N_1811,N_1747);
and U2152 (N_2152,N_1502,N_1972);
nand U2153 (N_2153,N_1585,N_1850);
nand U2154 (N_2154,N_1938,N_1784);
and U2155 (N_2155,N_1900,N_1767);
nand U2156 (N_2156,N_1820,N_1544);
nand U2157 (N_2157,N_1828,N_1554);
nor U2158 (N_2158,N_1630,N_1582);
or U2159 (N_2159,N_1750,N_1885);
xor U2160 (N_2160,N_1867,N_1738);
and U2161 (N_2161,N_1545,N_1821);
and U2162 (N_2162,N_1518,N_1911);
nor U2163 (N_2163,N_1694,N_1992);
xnor U2164 (N_2164,N_1921,N_1612);
and U2165 (N_2165,N_1676,N_1628);
xnor U2166 (N_2166,N_1888,N_1539);
and U2167 (N_2167,N_1855,N_1566);
nor U2168 (N_2168,N_1881,N_1538);
nor U2169 (N_2169,N_1616,N_1614);
nor U2170 (N_2170,N_1701,N_1813);
nand U2171 (N_2171,N_1596,N_1928);
nand U2172 (N_2172,N_1857,N_1765);
or U2173 (N_2173,N_1509,N_1982);
xnor U2174 (N_2174,N_1873,N_1999);
nor U2175 (N_2175,N_1755,N_1935);
nor U2176 (N_2176,N_1549,N_1810);
and U2177 (N_2177,N_1891,N_1758);
or U2178 (N_2178,N_1870,N_1853);
or U2179 (N_2179,N_1760,N_1836);
and U2180 (N_2180,N_1619,N_1969);
and U2181 (N_2181,N_1787,N_1843);
or U2182 (N_2182,N_1557,N_1749);
and U2183 (N_2183,N_1780,N_1724);
nand U2184 (N_2184,N_1915,N_1859);
nand U2185 (N_2185,N_1863,N_1903);
or U2186 (N_2186,N_1712,N_1552);
nand U2187 (N_2187,N_1975,N_1752);
nor U2188 (N_2188,N_1733,N_1751);
or U2189 (N_2189,N_1584,N_1625);
nand U2190 (N_2190,N_1886,N_1597);
or U2191 (N_2191,N_1744,N_1844);
nand U2192 (N_2192,N_1609,N_1677);
nand U2193 (N_2193,N_1690,N_1832);
nor U2194 (N_2194,N_1559,N_1711);
or U2195 (N_2195,N_1506,N_1603);
nand U2196 (N_2196,N_1768,N_1564);
nor U2197 (N_2197,N_1505,N_1835);
nor U2198 (N_2198,N_1615,N_1899);
nand U2199 (N_2199,N_1894,N_1804);
nand U2200 (N_2200,N_1824,N_1631);
nor U2201 (N_2201,N_1996,N_1976);
or U2202 (N_2202,N_1666,N_1907);
or U2203 (N_2203,N_1988,N_1848);
nand U2204 (N_2204,N_1581,N_1521);
nor U2205 (N_2205,N_1713,N_1573);
xnor U2206 (N_2206,N_1968,N_1702);
or U2207 (N_2207,N_1634,N_1834);
xor U2208 (N_2208,N_1995,N_1771);
nor U2209 (N_2209,N_1635,N_1974);
and U2210 (N_2210,N_1754,N_1801);
nor U2211 (N_2211,N_1569,N_1918);
or U2212 (N_2212,N_1778,N_1795);
nand U2213 (N_2213,N_1997,N_1729);
or U2214 (N_2214,N_1840,N_1865);
and U2215 (N_2215,N_1914,N_1773);
and U2216 (N_2216,N_1860,N_1783);
and U2217 (N_2217,N_1689,N_1520);
nor U2218 (N_2218,N_1800,N_1827);
or U2219 (N_2219,N_1686,N_1656);
nand U2220 (N_2220,N_1529,N_1759);
nand U2221 (N_2221,N_1819,N_1661);
nand U2222 (N_2222,N_1812,N_1643);
xor U2223 (N_2223,N_1647,N_1576);
nand U2224 (N_2224,N_1786,N_1993);
nor U2225 (N_2225,N_1932,N_1920);
nand U2226 (N_2226,N_1626,N_1849);
nor U2227 (N_2227,N_1662,N_1861);
and U2228 (N_2228,N_1633,N_1814);
or U2229 (N_2229,N_1785,N_1533);
and U2230 (N_2230,N_1892,N_1706);
nor U2231 (N_2231,N_1782,N_1512);
nand U2232 (N_2232,N_1736,N_1598);
or U2233 (N_2233,N_1959,N_1793);
nand U2234 (N_2234,N_1825,N_1645);
nor U2235 (N_2235,N_1594,N_1858);
nor U2236 (N_2236,N_1973,N_1880);
or U2237 (N_2237,N_1590,N_1682);
nand U2238 (N_2238,N_1687,N_1511);
nor U2239 (N_2239,N_1852,N_1826);
and U2240 (N_2240,N_1652,N_1833);
and U2241 (N_2241,N_1548,N_1805);
nand U2242 (N_2242,N_1636,N_1562);
or U2243 (N_2243,N_1839,N_1809);
or U2244 (N_2244,N_1779,N_1978);
nor U2245 (N_2245,N_1620,N_1985);
nand U2246 (N_2246,N_1561,N_1709);
xor U2247 (N_2247,N_1606,N_1527);
nor U2248 (N_2248,N_1847,N_1679);
nand U2249 (N_2249,N_1730,N_1845);
nand U2250 (N_2250,N_1513,N_1935);
xor U2251 (N_2251,N_1537,N_1556);
nand U2252 (N_2252,N_1955,N_1578);
and U2253 (N_2253,N_1949,N_1848);
xor U2254 (N_2254,N_1544,N_1843);
and U2255 (N_2255,N_1876,N_1740);
nand U2256 (N_2256,N_1586,N_1690);
nand U2257 (N_2257,N_1672,N_1720);
nand U2258 (N_2258,N_1513,N_1992);
xnor U2259 (N_2259,N_1964,N_1785);
and U2260 (N_2260,N_1562,N_1772);
nor U2261 (N_2261,N_1891,N_1549);
or U2262 (N_2262,N_1683,N_1846);
nor U2263 (N_2263,N_1894,N_1527);
and U2264 (N_2264,N_1778,N_1966);
nand U2265 (N_2265,N_1974,N_1820);
nor U2266 (N_2266,N_1760,N_1744);
nor U2267 (N_2267,N_1921,N_1707);
nand U2268 (N_2268,N_1581,N_1725);
or U2269 (N_2269,N_1700,N_1893);
and U2270 (N_2270,N_1928,N_1745);
nor U2271 (N_2271,N_1862,N_1869);
xor U2272 (N_2272,N_1648,N_1852);
xor U2273 (N_2273,N_1737,N_1898);
nand U2274 (N_2274,N_1764,N_1567);
nand U2275 (N_2275,N_1812,N_1600);
or U2276 (N_2276,N_1583,N_1504);
nor U2277 (N_2277,N_1927,N_1851);
nor U2278 (N_2278,N_1504,N_1915);
nand U2279 (N_2279,N_1733,N_1670);
or U2280 (N_2280,N_1950,N_1753);
nor U2281 (N_2281,N_1555,N_1796);
or U2282 (N_2282,N_1699,N_1913);
nand U2283 (N_2283,N_1734,N_1801);
xnor U2284 (N_2284,N_1781,N_1625);
and U2285 (N_2285,N_1781,N_1835);
nor U2286 (N_2286,N_1518,N_1558);
and U2287 (N_2287,N_1834,N_1934);
xnor U2288 (N_2288,N_1683,N_1688);
and U2289 (N_2289,N_1685,N_1752);
and U2290 (N_2290,N_1709,N_1678);
and U2291 (N_2291,N_1524,N_1885);
nand U2292 (N_2292,N_1579,N_1851);
and U2293 (N_2293,N_1965,N_1533);
nor U2294 (N_2294,N_1772,N_1935);
nand U2295 (N_2295,N_1779,N_1953);
nor U2296 (N_2296,N_1862,N_1665);
nor U2297 (N_2297,N_1963,N_1635);
nand U2298 (N_2298,N_1952,N_1850);
and U2299 (N_2299,N_1661,N_1510);
or U2300 (N_2300,N_1612,N_1898);
and U2301 (N_2301,N_1761,N_1705);
and U2302 (N_2302,N_1542,N_1560);
or U2303 (N_2303,N_1663,N_1741);
or U2304 (N_2304,N_1791,N_1652);
or U2305 (N_2305,N_1622,N_1985);
or U2306 (N_2306,N_1964,N_1530);
and U2307 (N_2307,N_1830,N_1986);
and U2308 (N_2308,N_1862,N_1780);
and U2309 (N_2309,N_1556,N_1605);
or U2310 (N_2310,N_1714,N_1565);
nand U2311 (N_2311,N_1580,N_1957);
and U2312 (N_2312,N_1605,N_1654);
nand U2313 (N_2313,N_1605,N_1982);
nor U2314 (N_2314,N_1546,N_1662);
nand U2315 (N_2315,N_1520,N_1949);
nor U2316 (N_2316,N_1922,N_1626);
nor U2317 (N_2317,N_1822,N_1570);
nor U2318 (N_2318,N_1723,N_1895);
nand U2319 (N_2319,N_1535,N_1882);
nor U2320 (N_2320,N_1934,N_1671);
and U2321 (N_2321,N_1529,N_1536);
and U2322 (N_2322,N_1649,N_1811);
and U2323 (N_2323,N_1525,N_1831);
or U2324 (N_2324,N_1683,N_1778);
xnor U2325 (N_2325,N_1824,N_1798);
nand U2326 (N_2326,N_1968,N_1533);
or U2327 (N_2327,N_1697,N_1928);
nand U2328 (N_2328,N_1846,N_1636);
nor U2329 (N_2329,N_1956,N_1783);
xnor U2330 (N_2330,N_1601,N_1989);
nor U2331 (N_2331,N_1874,N_1902);
nand U2332 (N_2332,N_1711,N_1988);
nand U2333 (N_2333,N_1871,N_1752);
nand U2334 (N_2334,N_1663,N_1649);
or U2335 (N_2335,N_1677,N_1550);
or U2336 (N_2336,N_1819,N_1738);
or U2337 (N_2337,N_1850,N_1853);
nor U2338 (N_2338,N_1701,N_1738);
nor U2339 (N_2339,N_1752,N_1705);
xnor U2340 (N_2340,N_1906,N_1968);
nand U2341 (N_2341,N_1916,N_1564);
and U2342 (N_2342,N_1672,N_1634);
or U2343 (N_2343,N_1764,N_1630);
xnor U2344 (N_2344,N_1866,N_1794);
nand U2345 (N_2345,N_1583,N_1800);
and U2346 (N_2346,N_1853,N_1839);
nor U2347 (N_2347,N_1755,N_1689);
or U2348 (N_2348,N_1983,N_1934);
or U2349 (N_2349,N_1798,N_1871);
nand U2350 (N_2350,N_1666,N_1890);
nand U2351 (N_2351,N_1808,N_1661);
or U2352 (N_2352,N_1655,N_1519);
nand U2353 (N_2353,N_1832,N_1853);
xnor U2354 (N_2354,N_1756,N_1750);
nor U2355 (N_2355,N_1631,N_1595);
nor U2356 (N_2356,N_1660,N_1792);
nand U2357 (N_2357,N_1697,N_1564);
nand U2358 (N_2358,N_1925,N_1712);
nand U2359 (N_2359,N_1943,N_1605);
or U2360 (N_2360,N_1563,N_1508);
and U2361 (N_2361,N_1928,N_1723);
and U2362 (N_2362,N_1839,N_1731);
or U2363 (N_2363,N_1913,N_1524);
or U2364 (N_2364,N_1794,N_1612);
nand U2365 (N_2365,N_1792,N_1994);
nand U2366 (N_2366,N_1604,N_1870);
nand U2367 (N_2367,N_1889,N_1614);
nor U2368 (N_2368,N_1564,N_1925);
nand U2369 (N_2369,N_1899,N_1601);
and U2370 (N_2370,N_1702,N_1841);
and U2371 (N_2371,N_1648,N_1552);
or U2372 (N_2372,N_1848,N_1829);
nand U2373 (N_2373,N_1543,N_1569);
and U2374 (N_2374,N_1614,N_1923);
or U2375 (N_2375,N_1668,N_1736);
and U2376 (N_2376,N_1701,N_1623);
or U2377 (N_2377,N_1932,N_1854);
xor U2378 (N_2378,N_1847,N_1677);
or U2379 (N_2379,N_1938,N_1806);
nand U2380 (N_2380,N_1989,N_1753);
and U2381 (N_2381,N_1869,N_1842);
xor U2382 (N_2382,N_1811,N_1784);
nor U2383 (N_2383,N_1726,N_1756);
nor U2384 (N_2384,N_1576,N_1875);
nand U2385 (N_2385,N_1650,N_1917);
nor U2386 (N_2386,N_1580,N_1925);
or U2387 (N_2387,N_1878,N_1752);
nand U2388 (N_2388,N_1748,N_1859);
nor U2389 (N_2389,N_1503,N_1663);
nor U2390 (N_2390,N_1636,N_1780);
or U2391 (N_2391,N_1959,N_1982);
or U2392 (N_2392,N_1763,N_1724);
and U2393 (N_2393,N_1858,N_1703);
and U2394 (N_2394,N_1953,N_1997);
xor U2395 (N_2395,N_1690,N_1599);
nand U2396 (N_2396,N_1669,N_1565);
nor U2397 (N_2397,N_1650,N_1733);
nand U2398 (N_2398,N_1980,N_1813);
and U2399 (N_2399,N_1796,N_1785);
xnor U2400 (N_2400,N_1820,N_1946);
nor U2401 (N_2401,N_1947,N_1983);
nand U2402 (N_2402,N_1884,N_1992);
nand U2403 (N_2403,N_1606,N_1801);
or U2404 (N_2404,N_1530,N_1853);
or U2405 (N_2405,N_1873,N_1871);
nor U2406 (N_2406,N_1529,N_1719);
or U2407 (N_2407,N_1716,N_1968);
and U2408 (N_2408,N_1795,N_1637);
nor U2409 (N_2409,N_1541,N_1658);
and U2410 (N_2410,N_1824,N_1836);
or U2411 (N_2411,N_1522,N_1773);
and U2412 (N_2412,N_1781,N_1762);
nor U2413 (N_2413,N_1721,N_1892);
or U2414 (N_2414,N_1626,N_1641);
xnor U2415 (N_2415,N_1788,N_1527);
or U2416 (N_2416,N_1634,N_1712);
nor U2417 (N_2417,N_1628,N_1917);
and U2418 (N_2418,N_1516,N_1600);
or U2419 (N_2419,N_1971,N_1874);
nor U2420 (N_2420,N_1708,N_1687);
or U2421 (N_2421,N_1914,N_1952);
nor U2422 (N_2422,N_1645,N_1695);
nand U2423 (N_2423,N_1968,N_1827);
or U2424 (N_2424,N_1849,N_1848);
xor U2425 (N_2425,N_1611,N_1975);
nand U2426 (N_2426,N_1704,N_1777);
or U2427 (N_2427,N_1559,N_1848);
or U2428 (N_2428,N_1814,N_1974);
or U2429 (N_2429,N_1615,N_1769);
and U2430 (N_2430,N_1666,N_1557);
nand U2431 (N_2431,N_1583,N_1670);
or U2432 (N_2432,N_1714,N_1665);
nand U2433 (N_2433,N_1978,N_1511);
and U2434 (N_2434,N_1607,N_1979);
and U2435 (N_2435,N_1721,N_1801);
nor U2436 (N_2436,N_1652,N_1773);
or U2437 (N_2437,N_1938,N_1888);
nor U2438 (N_2438,N_1643,N_1743);
nor U2439 (N_2439,N_1502,N_1677);
or U2440 (N_2440,N_1843,N_1829);
or U2441 (N_2441,N_1859,N_1615);
nor U2442 (N_2442,N_1965,N_1762);
or U2443 (N_2443,N_1837,N_1900);
or U2444 (N_2444,N_1970,N_1714);
and U2445 (N_2445,N_1591,N_1521);
nor U2446 (N_2446,N_1748,N_1787);
and U2447 (N_2447,N_1845,N_1631);
or U2448 (N_2448,N_1686,N_1659);
nor U2449 (N_2449,N_1559,N_1685);
xor U2450 (N_2450,N_1605,N_1607);
nor U2451 (N_2451,N_1773,N_1809);
or U2452 (N_2452,N_1703,N_1794);
and U2453 (N_2453,N_1950,N_1825);
nand U2454 (N_2454,N_1818,N_1783);
or U2455 (N_2455,N_1648,N_1578);
or U2456 (N_2456,N_1563,N_1891);
nand U2457 (N_2457,N_1685,N_1897);
and U2458 (N_2458,N_1926,N_1535);
xnor U2459 (N_2459,N_1762,N_1544);
and U2460 (N_2460,N_1970,N_1877);
or U2461 (N_2461,N_1862,N_1685);
nand U2462 (N_2462,N_1616,N_1760);
and U2463 (N_2463,N_1704,N_1598);
and U2464 (N_2464,N_1863,N_1841);
nor U2465 (N_2465,N_1947,N_1719);
nor U2466 (N_2466,N_1942,N_1822);
or U2467 (N_2467,N_1635,N_1688);
or U2468 (N_2468,N_1804,N_1622);
nor U2469 (N_2469,N_1936,N_1735);
or U2470 (N_2470,N_1586,N_1509);
xor U2471 (N_2471,N_1725,N_1598);
and U2472 (N_2472,N_1568,N_1971);
and U2473 (N_2473,N_1582,N_1959);
nand U2474 (N_2474,N_1559,N_1846);
nor U2475 (N_2475,N_1950,N_1542);
nor U2476 (N_2476,N_1834,N_1916);
and U2477 (N_2477,N_1935,N_1643);
xor U2478 (N_2478,N_1611,N_1706);
and U2479 (N_2479,N_1898,N_1742);
xor U2480 (N_2480,N_1630,N_1650);
nand U2481 (N_2481,N_1581,N_1579);
nand U2482 (N_2482,N_1769,N_1770);
nor U2483 (N_2483,N_1581,N_1655);
nand U2484 (N_2484,N_1595,N_1689);
and U2485 (N_2485,N_1868,N_1995);
nor U2486 (N_2486,N_1897,N_1501);
or U2487 (N_2487,N_1740,N_1968);
or U2488 (N_2488,N_1952,N_1901);
nor U2489 (N_2489,N_1863,N_1681);
or U2490 (N_2490,N_1651,N_1782);
and U2491 (N_2491,N_1554,N_1817);
and U2492 (N_2492,N_1609,N_1604);
or U2493 (N_2493,N_1577,N_1729);
nand U2494 (N_2494,N_1958,N_1781);
xnor U2495 (N_2495,N_1683,N_1920);
or U2496 (N_2496,N_1666,N_1608);
nor U2497 (N_2497,N_1986,N_1759);
or U2498 (N_2498,N_1881,N_1537);
and U2499 (N_2499,N_1990,N_1745);
xnor U2500 (N_2500,N_2354,N_2128);
nor U2501 (N_2501,N_2203,N_2178);
and U2502 (N_2502,N_2239,N_2171);
and U2503 (N_2503,N_2197,N_2134);
nor U2504 (N_2504,N_2157,N_2492);
or U2505 (N_2505,N_2450,N_2117);
and U2506 (N_2506,N_2436,N_2408);
nand U2507 (N_2507,N_2221,N_2010);
nor U2508 (N_2508,N_2074,N_2388);
nor U2509 (N_2509,N_2270,N_2481);
nor U2510 (N_2510,N_2497,N_2030);
or U2511 (N_2511,N_2173,N_2261);
nand U2512 (N_2512,N_2195,N_2381);
nand U2513 (N_2513,N_2147,N_2183);
nor U2514 (N_2514,N_2319,N_2426);
or U2515 (N_2515,N_2027,N_2371);
and U2516 (N_2516,N_2475,N_2015);
nand U2517 (N_2517,N_2046,N_2367);
nand U2518 (N_2518,N_2004,N_2212);
nor U2519 (N_2519,N_2132,N_2440);
nor U2520 (N_2520,N_2277,N_2357);
nor U2521 (N_2521,N_2441,N_2324);
and U2522 (N_2522,N_2122,N_2405);
or U2523 (N_2523,N_2269,N_2148);
xor U2524 (N_2524,N_2067,N_2322);
xnor U2525 (N_2525,N_2411,N_2244);
or U2526 (N_2526,N_2320,N_2126);
and U2527 (N_2527,N_2169,N_2361);
or U2528 (N_2528,N_2020,N_2356);
and U2529 (N_2529,N_2069,N_2394);
or U2530 (N_2530,N_2419,N_2323);
or U2531 (N_2531,N_2168,N_2434);
or U2532 (N_2532,N_2136,N_2124);
nor U2533 (N_2533,N_2120,N_2187);
and U2534 (N_2534,N_2123,N_2284);
nor U2535 (N_2535,N_2303,N_2457);
or U2536 (N_2536,N_2039,N_2421);
or U2537 (N_2537,N_2036,N_2154);
and U2538 (N_2538,N_2080,N_2352);
nor U2539 (N_2539,N_2174,N_2179);
nand U2540 (N_2540,N_2002,N_2022);
and U2541 (N_2541,N_2012,N_2344);
or U2542 (N_2542,N_2470,N_2077);
and U2543 (N_2543,N_2149,N_2225);
nand U2544 (N_2544,N_2376,N_2140);
nor U2545 (N_2545,N_2137,N_2101);
nand U2546 (N_2546,N_2307,N_2448);
xor U2547 (N_2547,N_2274,N_2446);
or U2548 (N_2548,N_2218,N_2034);
and U2549 (N_2549,N_2198,N_2420);
or U2550 (N_2550,N_2283,N_2143);
nor U2551 (N_2551,N_2483,N_2110);
nand U2552 (N_2552,N_2162,N_2360);
and U2553 (N_2553,N_2488,N_2359);
nor U2554 (N_2554,N_2484,N_2460);
or U2555 (N_2555,N_2445,N_2275);
or U2556 (N_2556,N_2098,N_2097);
nand U2557 (N_2557,N_2316,N_2469);
xor U2558 (N_2558,N_2427,N_2145);
and U2559 (N_2559,N_2202,N_2008);
nand U2560 (N_2560,N_2175,N_2247);
nor U2561 (N_2561,N_2415,N_2289);
or U2562 (N_2562,N_2418,N_2035);
nand U2563 (N_2563,N_2048,N_2076);
and U2564 (N_2564,N_2262,N_2482);
nor U2565 (N_2565,N_2089,N_2437);
nor U2566 (N_2566,N_2465,N_2379);
and U2567 (N_2567,N_2204,N_2127);
and U2568 (N_2568,N_2406,N_2314);
and U2569 (N_2569,N_2310,N_2332);
or U2570 (N_2570,N_2208,N_2150);
or U2571 (N_2571,N_2409,N_2064);
xor U2572 (N_2572,N_2164,N_2188);
or U2573 (N_2573,N_2373,N_2059);
or U2574 (N_2574,N_2321,N_2290);
and U2575 (N_2575,N_2205,N_2199);
or U2576 (N_2576,N_2263,N_2298);
nand U2577 (N_2577,N_2103,N_2302);
or U2578 (N_2578,N_2196,N_2153);
nand U2579 (N_2579,N_2336,N_2297);
or U2580 (N_2580,N_2313,N_2000);
and U2581 (N_2581,N_2232,N_2037);
and U2582 (N_2582,N_2100,N_2119);
nand U2583 (N_2583,N_2057,N_2021);
nor U2584 (N_2584,N_2439,N_2180);
nand U2585 (N_2585,N_2355,N_2487);
or U2586 (N_2586,N_2172,N_2102);
nand U2587 (N_2587,N_2209,N_2493);
nor U2588 (N_2588,N_2392,N_2294);
or U2589 (N_2589,N_2315,N_2082);
nor U2590 (N_2590,N_2312,N_2073);
nor U2591 (N_2591,N_2366,N_2351);
nor U2592 (N_2592,N_2045,N_2139);
and U2593 (N_2593,N_2333,N_2473);
nor U2594 (N_2594,N_2248,N_2402);
nor U2595 (N_2595,N_2112,N_2087);
or U2596 (N_2596,N_2255,N_2217);
xnor U2597 (N_2597,N_2412,N_2184);
nand U2598 (N_2598,N_2335,N_2466);
nand U2599 (N_2599,N_2456,N_2029);
and U2600 (N_2600,N_2464,N_2194);
nor U2601 (N_2601,N_2115,N_2243);
xnor U2602 (N_2602,N_2461,N_2489);
or U2603 (N_2603,N_2267,N_2328);
or U2604 (N_2604,N_2084,N_2014);
and U2605 (N_2605,N_2295,N_2342);
nand U2606 (N_2606,N_2214,N_2276);
nand U2607 (N_2607,N_2410,N_2395);
or U2608 (N_2608,N_2404,N_2398);
and U2609 (N_2609,N_2341,N_2279);
or U2610 (N_2610,N_2038,N_2495);
nand U2611 (N_2611,N_2401,N_2040);
nand U2612 (N_2612,N_2161,N_2216);
and U2613 (N_2613,N_2167,N_2451);
and U2614 (N_2614,N_2477,N_2429);
xnor U2615 (N_2615,N_2215,N_2416);
nand U2616 (N_2616,N_2058,N_2236);
and U2617 (N_2617,N_2424,N_2479);
xor U2618 (N_2618,N_2056,N_2079);
nand U2619 (N_2619,N_2235,N_2054);
or U2620 (N_2620,N_2330,N_2345);
and U2621 (N_2621,N_2085,N_2386);
and U2622 (N_2622,N_2285,N_2287);
nand U2623 (N_2623,N_2304,N_2467);
and U2624 (N_2624,N_2348,N_2016);
nand U2625 (N_2625,N_2389,N_2340);
nor U2626 (N_2626,N_2374,N_2141);
or U2627 (N_2627,N_2219,N_2350);
nand U2628 (N_2628,N_2189,N_2220);
or U2629 (N_2629,N_2156,N_2454);
nand U2630 (N_2630,N_2393,N_2023);
or U2631 (N_2631,N_2111,N_2490);
or U2632 (N_2632,N_2377,N_2009);
and U2633 (N_2633,N_2363,N_2498);
nand U2634 (N_2634,N_2170,N_2055);
or U2635 (N_2635,N_2397,N_2468);
or U2636 (N_2636,N_2472,N_2017);
nor U2637 (N_2637,N_2181,N_2301);
nand U2638 (N_2638,N_2364,N_2449);
nor U2639 (N_2639,N_2288,N_2400);
nand U2640 (N_2640,N_2268,N_2391);
nand U2641 (N_2641,N_2086,N_2072);
or U2642 (N_2642,N_2240,N_2191);
or U2643 (N_2643,N_2083,N_2491);
nor U2644 (N_2644,N_2192,N_2380);
and U2645 (N_2645,N_2200,N_2226);
nand U2646 (N_2646,N_2423,N_2003);
nor U2647 (N_2647,N_2052,N_2019);
nand U2648 (N_2648,N_2211,N_2384);
nand U2649 (N_2649,N_2358,N_2455);
and U2650 (N_2650,N_2264,N_2249);
nor U2651 (N_2651,N_2349,N_2442);
nor U2652 (N_2652,N_2485,N_2066);
and U2653 (N_2653,N_2337,N_2458);
and U2654 (N_2654,N_2210,N_2193);
nor U2655 (N_2655,N_2043,N_2362);
nor U2656 (N_2656,N_2387,N_2265);
nor U2657 (N_2657,N_2282,N_2432);
nand U2658 (N_2658,N_2163,N_2113);
or U2659 (N_2659,N_2447,N_2453);
or U2660 (N_2660,N_2329,N_2166);
xor U2661 (N_2661,N_2372,N_2254);
or U2662 (N_2662,N_2185,N_2257);
or U2663 (N_2663,N_2144,N_2496);
nand U2664 (N_2664,N_2026,N_2025);
and U2665 (N_2665,N_2096,N_2234);
or U2666 (N_2666,N_2223,N_2383);
or U2667 (N_2667,N_2070,N_2047);
or U2668 (N_2668,N_2382,N_2186);
nand U2669 (N_2669,N_2272,N_2031);
nor U2670 (N_2670,N_2499,N_2001);
xor U2671 (N_2671,N_2114,N_2463);
and U2672 (N_2672,N_2281,N_2241);
and U2673 (N_2673,N_2414,N_2266);
nand U2674 (N_2674,N_2133,N_2271);
or U2675 (N_2675,N_2011,N_2245);
nor U2676 (N_2676,N_2152,N_2233);
nand U2677 (N_2677,N_2155,N_2273);
nor U2678 (N_2678,N_2078,N_2190);
and U2679 (N_2679,N_2251,N_2396);
or U2680 (N_2680,N_2105,N_2293);
nor U2681 (N_2681,N_2231,N_2109);
nand U2682 (N_2682,N_2068,N_2378);
or U2683 (N_2683,N_2435,N_2088);
nand U2684 (N_2684,N_2028,N_2075);
and U2685 (N_2685,N_2158,N_2253);
nand U2686 (N_2686,N_2032,N_2474);
or U2687 (N_2687,N_2159,N_2121);
nor U2688 (N_2688,N_2090,N_2252);
or U2689 (N_2689,N_2176,N_2042);
or U2690 (N_2690,N_2227,N_2331);
or U2691 (N_2691,N_2049,N_2033);
xnor U2692 (N_2692,N_2428,N_2370);
nor U2693 (N_2693,N_2369,N_2146);
xnor U2694 (N_2694,N_2177,N_2403);
xnor U2695 (N_2695,N_2041,N_2259);
nor U2696 (N_2696,N_2125,N_2480);
or U2697 (N_2697,N_2308,N_2325);
nor U2698 (N_2698,N_2433,N_2305);
nor U2699 (N_2699,N_2237,N_2095);
nand U2700 (N_2700,N_2151,N_2062);
and U2701 (N_2701,N_2007,N_2365);
nor U2702 (N_2702,N_2334,N_2182);
nand U2703 (N_2703,N_2063,N_2207);
or U2704 (N_2704,N_2104,N_2343);
and U2705 (N_2705,N_2051,N_2230);
nand U2706 (N_2706,N_2224,N_2246);
and U2707 (N_2707,N_2107,N_2385);
nor U2708 (N_2708,N_2462,N_2353);
xnor U2709 (N_2709,N_2229,N_2425);
or U2710 (N_2710,N_2339,N_2430);
nand U2711 (N_2711,N_2222,N_2013);
nand U2712 (N_2712,N_2443,N_2160);
or U2713 (N_2713,N_2138,N_2309);
nor U2714 (N_2714,N_2306,N_2093);
nand U2715 (N_2715,N_2478,N_2044);
xnor U2716 (N_2716,N_2201,N_2286);
nor U2717 (N_2717,N_2053,N_2071);
nand U2718 (N_2718,N_2135,N_2399);
and U2719 (N_2719,N_2118,N_2296);
and U2720 (N_2720,N_2486,N_2311);
nor U2721 (N_2721,N_2317,N_2094);
and U2722 (N_2722,N_2061,N_2347);
or U2723 (N_2723,N_2129,N_2116);
nand U2724 (N_2724,N_2250,N_2368);
and U2725 (N_2725,N_2142,N_2131);
nor U2726 (N_2726,N_2476,N_2299);
or U2727 (N_2727,N_2228,N_2108);
nand U2728 (N_2728,N_2238,N_2318);
nand U2729 (N_2729,N_2291,N_2431);
xnor U2730 (N_2730,N_2407,N_2422);
nor U2731 (N_2731,N_2390,N_2438);
or U2732 (N_2732,N_2459,N_2256);
nand U2733 (N_2733,N_2258,N_2081);
or U2734 (N_2734,N_2006,N_2024);
nor U2735 (N_2735,N_2280,N_2060);
and U2736 (N_2736,N_2018,N_2413);
xor U2737 (N_2737,N_2292,N_2091);
nor U2738 (N_2738,N_2494,N_2346);
nand U2739 (N_2739,N_2452,N_2375);
or U2740 (N_2740,N_2213,N_2444);
and U2741 (N_2741,N_2165,N_2326);
nor U2742 (N_2742,N_2260,N_2417);
and U2743 (N_2743,N_2471,N_2338);
and U2744 (N_2744,N_2278,N_2206);
and U2745 (N_2745,N_2005,N_2106);
xnor U2746 (N_2746,N_2050,N_2065);
nand U2747 (N_2747,N_2092,N_2099);
or U2748 (N_2748,N_2242,N_2130);
or U2749 (N_2749,N_2300,N_2327);
or U2750 (N_2750,N_2263,N_2187);
and U2751 (N_2751,N_2015,N_2433);
or U2752 (N_2752,N_2174,N_2315);
nor U2753 (N_2753,N_2094,N_2467);
nand U2754 (N_2754,N_2470,N_2440);
and U2755 (N_2755,N_2265,N_2328);
and U2756 (N_2756,N_2015,N_2219);
nand U2757 (N_2757,N_2453,N_2461);
and U2758 (N_2758,N_2090,N_2026);
or U2759 (N_2759,N_2257,N_2245);
or U2760 (N_2760,N_2015,N_2499);
xor U2761 (N_2761,N_2026,N_2203);
xnor U2762 (N_2762,N_2443,N_2023);
nand U2763 (N_2763,N_2191,N_2342);
nor U2764 (N_2764,N_2354,N_2161);
nand U2765 (N_2765,N_2145,N_2008);
nand U2766 (N_2766,N_2378,N_2012);
nand U2767 (N_2767,N_2473,N_2438);
nor U2768 (N_2768,N_2369,N_2178);
or U2769 (N_2769,N_2398,N_2177);
nor U2770 (N_2770,N_2378,N_2186);
and U2771 (N_2771,N_2353,N_2467);
nand U2772 (N_2772,N_2161,N_2111);
nor U2773 (N_2773,N_2360,N_2335);
nand U2774 (N_2774,N_2352,N_2252);
or U2775 (N_2775,N_2351,N_2339);
or U2776 (N_2776,N_2354,N_2010);
and U2777 (N_2777,N_2242,N_2019);
nor U2778 (N_2778,N_2108,N_2103);
nand U2779 (N_2779,N_2079,N_2082);
nand U2780 (N_2780,N_2010,N_2282);
and U2781 (N_2781,N_2485,N_2011);
and U2782 (N_2782,N_2221,N_2250);
nor U2783 (N_2783,N_2038,N_2006);
and U2784 (N_2784,N_2387,N_2211);
and U2785 (N_2785,N_2186,N_2080);
xnor U2786 (N_2786,N_2314,N_2045);
nor U2787 (N_2787,N_2154,N_2239);
or U2788 (N_2788,N_2455,N_2335);
nand U2789 (N_2789,N_2139,N_2163);
nand U2790 (N_2790,N_2407,N_2240);
or U2791 (N_2791,N_2158,N_2218);
nor U2792 (N_2792,N_2484,N_2214);
nand U2793 (N_2793,N_2282,N_2216);
and U2794 (N_2794,N_2488,N_2001);
nand U2795 (N_2795,N_2375,N_2496);
or U2796 (N_2796,N_2070,N_2406);
nor U2797 (N_2797,N_2371,N_2357);
and U2798 (N_2798,N_2188,N_2436);
nor U2799 (N_2799,N_2141,N_2498);
or U2800 (N_2800,N_2198,N_2460);
nor U2801 (N_2801,N_2213,N_2434);
nand U2802 (N_2802,N_2484,N_2376);
nor U2803 (N_2803,N_2178,N_2101);
and U2804 (N_2804,N_2464,N_2356);
or U2805 (N_2805,N_2175,N_2339);
xor U2806 (N_2806,N_2308,N_2370);
or U2807 (N_2807,N_2167,N_2046);
nor U2808 (N_2808,N_2284,N_2198);
nand U2809 (N_2809,N_2430,N_2452);
or U2810 (N_2810,N_2036,N_2168);
or U2811 (N_2811,N_2233,N_2160);
or U2812 (N_2812,N_2340,N_2077);
or U2813 (N_2813,N_2234,N_2468);
and U2814 (N_2814,N_2040,N_2087);
nand U2815 (N_2815,N_2044,N_2489);
xnor U2816 (N_2816,N_2327,N_2317);
xor U2817 (N_2817,N_2138,N_2319);
and U2818 (N_2818,N_2005,N_2049);
and U2819 (N_2819,N_2071,N_2162);
or U2820 (N_2820,N_2285,N_2262);
nor U2821 (N_2821,N_2055,N_2496);
nand U2822 (N_2822,N_2073,N_2322);
nor U2823 (N_2823,N_2498,N_2399);
and U2824 (N_2824,N_2348,N_2424);
xnor U2825 (N_2825,N_2465,N_2155);
nor U2826 (N_2826,N_2303,N_2151);
or U2827 (N_2827,N_2138,N_2235);
and U2828 (N_2828,N_2475,N_2461);
nand U2829 (N_2829,N_2402,N_2102);
and U2830 (N_2830,N_2190,N_2185);
nor U2831 (N_2831,N_2467,N_2212);
and U2832 (N_2832,N_2257,N_2467);
and U2833 (N_2833,N_2403,N_2107);
or U2834 (N_2834,N_2465,N_2170);
xor U2835 (N_2835,N_2068,N_2344);
nor U2836 (N_2836,N_2162,N_2474);
or U2837 (N_2837,N_2491,N_2328);
nor U2838 (N_2838,N_2211,N_2118);
nand U2839 (N_2839,N_2179,N_2397);
nand U2840 (N_2840,N_2352,N_2159);
xor U2841 (N_2841,N_2235,N_2233);
xor U2842 (N_2842,N_2125,N_2360);
xnor U2843 (N_2843,N_2438,N_2244);
nand U2844 (N_2844,N_2361,N_2350);
nor U2845 (N_2845,N_2050,N_2110);
nor U2846 (N_2846,N_2280,N_2421);
nor U2847 (N_2847,N_2306,N_2132);
xnor U2848 (N_2848,N_2120,N_2015);
xnor U2849 (N_2849,N_2023,N_2204);
xor U2850 (N_2850,N_2049,N_2465);
and U2851 (N_2851,N_2039,N_2377);
or U2852 (N_2852,N_2285,N_2468);
nand U2853 (N_2853,N_2080,N_2313);
or U2854 (N_2854,N_2404,N_2422);
and U2855 (N_2855,N_2313,N_2388);
xnor U2856 (N_2856,N_2000,N_2228);
or U2857 (N_2857,N_2266,N_2281);
nand U2858 (N_2858,N_2404,N_2409);
nand U2859 (N_2859,N_2007,N_2290);
nor U2860 (N_2860,N_2027,N_2171);
nor U2861 (N_2861,N_2227,N_2462);
nor U2862 (N_2862,N_2408,N_2213);
or U2863 (N_2863,N_2274,N_2412);
or U2864 (N_2864,N_2492,N_2377);
nor U2865 (N_2865,N_2441,N_2252);
and U2866 (N_2866,N_2118,N_2129);
nor U2867 (N_2867,N_2393,N_2312);
nor U2868 (N_2868,N_2090,N_2112);
or U2869 (N_2869,N_2132,N_2488);
or U2870 (N_2870,N_2407,N_2390);
or U2871 (N_2871,N_2002,N_2042);
nand U2872 (N_2872,N_2191,N_2343);
nor U2873 (N_2873,N_2002,N_2006);
nor U2874 (N_2874,N_2134,N_2431);
or U2875 (N_2875,N_2120,N_2190);
or U2876 (N_2876,N_2490,N_2416);
nor U2877 (N_2877,N_2131,N_2180);
nor U2878 (N_2878,N_2060,N_2115);
xnor U2879 (N_2879,N_2140,N_2485);
nand U2880 (N_2880,N_2417,N_2423);
xnor U2881 (N_2881,N_2468,N_2250);
or U2882 (N_2882,N_2380,N_2410);
or U2883 (N_2883,N_2123,N_2430);
and U2884 (N_2884,N_2076,N_2071);
nand U2885 (N_2885,N_2353,N_2407);
nor U2886 (N_2886,N_2119,N_2087);
and U2887 (N_2887,N_2312,N_2035);
and U2888 (N_2888,N_2016,N_2438);
nand U2889 (N_2889,N_2210,N_2127);
nand U2890 (N_2890,N_2109,N_2235);
or U2891 (N_2891,N_2341,N_2259);
nor U2892 (N_2892,N_2114,N_2269);
or U2893 (N_2893,N_2452,N_2112);
or U2894 (N_2894,N_2380,N_2286);
nand U2895 (N_2895,N_2333,N_2039);
nand U2896 (N_2896,N_2066,N_2070);
and U2897 (N_2897,N_2403,N_2176);
nand U2898 (N_2898,N_2169,N_2307);
or U2899 (N_2899,N_2064,N_2350);
nand U2900 (N_2900,N_2070,N_2456);
nor U2901 (N_2901,N_2059,N_2409);
and U2902 (N_2902,N_2468,N_2142);
and U2903 (N_2903,N_2248,N_2304);
nand U2904 (N_2904,N_2415,N_2237);
or U2905 (N_2905,N_2236,N_2474);
nand U2906 (N_2906,N_2076,N_2233);
nor U2907 (N_2907,N_2186,N_2157);
and U2908 (N_2908,N_2011,N_2007);
and U2909 (N_2909,N_2121,N_2259);
or U2910 (N_2910,N_2210,N_2170);
xnor U2911 (N_2911,N_2356,N_2078);
or U2912 (N_2912,N_2281,N_2396);
and U2913 (N_2913,N_2087,N_2110);
and U2914 (N_2914,N_2358,N_2032);
xnor U2915 (N_2915,N_2127,N_2004);
nor U2916 (N_2916,N_2117,N_2237);
nand U2917 (N_2917,N_2453,N_2030);
nand U2918 (N_2918,N_2268,N_2081);
and U2919 (N_2919,N_2163,N_2119);
nand U2920 (N_2920,N_2497,N_2389);
or U2921 (N_2921,N_2457,N_2130);
nand U2922 (N_2922,N_2205,N_2299);
nor U2923 (N_2923,N_2377,N_2339);
and U2924 (N_2924,N_2283,N_2128);
and U2925 (N_2925,N_2370,N_2472);
nor U2926 (N_2926,N_2005,N_2186);
or U2927 (N_2927,N_2104,N_2008);
nand U2928 (N_2928,N_2308,N_2265);
xnor U2929 (N_2929,N_2390,N_2258);
nand U2930 (N_2930,N_2139,N_2237);
or U2931 (N_2931,N_2079,N_2048);
nor U2932 (N_2932,N_2466,N_2086);
or U2933 (N_2933,N_2438,N_2132);
and U2934 (N_2934,N_2029,N_2414);
xor U2935 (N_2935,N_2421,N_2305);
nand U2936 (N_2936,N_2092,N_2141);
nor U2937 (N_2937,N_2083,N_2433);
or U2938 (N_2938,N_2300,N_2121);
or U2939 (N_2939,N_2112,N_2091);
or U2940 (N_2940,N_2039,N_2078);
nor U2941 (N_2941,N_2483,N_2263);
nand U2942 (N_2942,N_2356,N_2442);
nand U2943 (N_2943,N_2197,N_2030);
nor U2944 (N_2944,N_2276,N_2138);
or U2945 (N_2945,N_2244,N_2314);
and U2946 (N_2946,N_2381,N_2371);
xor U2947 (N_2947,N_2005,N_2336);
nand U2948 (N_2948,N_2154,N_2398);
nand U2949 (N_2949,N_2499,N_2080);
and U2950 (N_2950,N_2201,N_2413);
or U2951 (N_2951,N_2253,N_2411);
and U2952 (N_2952,N_2498,N_2135);
and U2953 (N_2953,N_2474,N_2329);
and U2954 (N_2954,N_2428,N_2065);
nor U2955 (N_2955,N_2430,N_2336);
or U2956 (N_2956,N_2110,N_2467);
or U2957 (N_2957,N_2195,N_2052);
nor U2958 (N_2958,N_2175,N_2487);
or U2959 (N_2959,N_2225,N_2374);
xnor U2960 (N_2960,N_2048,N_2400);
nand U2961 (N_2961,N_2276,N_2414);
or U2962 (N_2962,N_2468,N_2258);
and U2963 (N_2963,N_2119,N_2285);
and U2964 (N_2964,N_2102,N_2214);
nand U2965 (N_2965,N_2024,N_2484);
nor U2966 (N_2966,N_2071,N_2368);
nand U2967 (N_2967,N_2498,N_2440);
or U2968 (N_2968,N_2198,N_2204);
and U2969 (N_2969,N_2226,N_2131);
or U2970 (N_2970,N_2169,N_2048);
or U2971 (N_2971,N_2253,N_2210);
nor U2972 (N_2972,N_2324,N_2325);
and U2973 (N_2973,N_2438,N_2314);
and U2974 (N_2974,N_2405,N_2088);
or U2975 (N_2975,N_2229,N_2432);
xnor U2976 (N_2976,N_2470,N_2318);
and U2977 (N_2977,N_2320,N_2137);
nor U2978 (N_2978,N_2331,N_2446);
nor U2979 (N_2979,N_2141,N_2178);
nand U2980 (N_2980,N_2087,N_2106);
nor U2981 (N_2981,N_2211,N_2180);
and U2982 (N_2982,N_2307,N_2111);
xnor U2983 (N_2983,N_2474,N_2231);
xnor U2984 (N_2984,N_2143,N_2019);
or U2985 (N_2985,N_2217,N_2393);
or U2986 (N_2986,N_2472,N_2050);
nor U2987 (N_2987,N_2422,N_2231);
or U2988 (N_2988,N_2386,N_2184);
or U2989 (N_2989,N_2335,N_2037);
and U2990 (N_2990,N_2259,N_2268);
nand U2991 (N_2991,N_2126,N_2177);
nor U2992 (N_2992,N_2142,N_2465);
xor U2993 (N_2993,N_2474,N_2212);
nand U2994 (N_2994,N_2193,N_2396);
and U2995 (N_2995,N_2114,N_2295);
nor U2996 (N_2996,N_2107,N_2056);
nor U2997 (N_2997,N_2385,N_2191);
and U2998 (N_2998,N_2317,N_2057);
xor U2999 (N_2999,N_2359,N_2066);
and U3000 (N_3000,N_2841,N_2911);
and U3001 (N_3001,N_2940,N_2877);
and U3002 (N_3002,N_2776,N_2824);
xnor U3003 (N_3003,N_2893,N_2927);
and U3004 (N_3004,N_2848,N_2992);
nor U3005 (N_3005,N_2552,N_2757);
nand U3006 (N_3006,N_2980,N_2801);
and U3007 (N_3007,N_2574,N_2862);
nand U3008 (N_3008,N_2813,N_2668);
nand U3009 (N_3009,N_2703,N_2968);
nand U3010 (N_3010,N_2545,N_2570);
and U3011 (N_3011,N_2993,N_2736);
or U3012 (N_3012,N_2505,N_2669);
nand U3013 (N_3013,N_2963,N_2845);
and U3014 (N_3014,N_2662,N_2796);
and U3015 (N_3015,N_2831,N_2956);
nand U3016 (N_3016,N_2648,N_2800);
or U3017 (N_3017,N_2684,N_2603);
nand U3018 (N_3018,N_2667,N_2925);
nor U3019 (N_3019,N_2853,N_2926);
nor U3020 (N_3020,N_2503,N_2528);
nand U3021 (N_3021,N_2971,N_2683);
xor U3022 (N_3022,N_2642,N_2794);
or U3023 (N_3023,N_2581,N_2799);
or U3024 (N_3024,N_2594,N_2534);
xor U3025 (N_3025,N_2596,N_2816);
nor U3026 (N_3026,N_2663,N_2515);
xnor U3027 (N_3027,N_2611,N_2692);
nor U3028 (N_3028,N_2922,N_2543);
nand U3029 (N_3029,N_2510,N_2532);
xnor U3030 (N_3030,N_2826,N_2641);
nand U3031 (N_3031,N_2944,N_2818);
or U3032 (N_3032,N_2599,N_2654);
nand U3033 (N_3033,N_2855,N_2598);
or U3034 (N_3034,N_2814,N_2961);
nand U3035 (N_3035,N_2907,N_2681);
nor U3036 (N_3036,N_2604,N_2873);
and U3037 (N_3037,N_2633,N_2730);
and U3038 (N_3038,N_2538,N_2626);
and U3039 (N_3039,N_2728,N_2595);
xnor U3040 (N_3040,N_2660,N_2951);
nand U3041 (N_3041,N_2618,N_2714);
nand U3042 (N_3042,N_2664,N_2973);
nand U3043 (N_3043,N_2665,N_2750);
nand U3044 (N_3044,N_2895,N_2868);
nor U3045 (N_3045,N_2754,N_2830);
nand U3046 (N_3046,N_2921,N_2740);
nand U3047 (N_3047,N_2960,N_2582);
xnor U3048 (N_3048,N_2704,N_2939);
xnor U3049 (N_3049,N_2717,N_2601);
nand U3050 (N_3050,N_2808,N_2896);
or U3051 (N_3051,N_2820,N_2978);
and U3052 (N_3052,N_2825,N_2766);
nor U3053 (N_3053,N_2865,N_2742);
nand U3054 (N_3054,N_2988,N_2624);
nor U3055 (N_3055,N_2914,N_2749);
xor U3056 (N_3056,N_2527,N_2649);
xnor U3057 (N_3057,N_2763,N_2919);
nand U3058 (N_3058,N_2844,N_2874);
or U3059 (N_3059,N_2615,N_2881);
nand U3060 (N_3060,N_2937,N_2608);
nor U3061 (N_3061,N_2835,N_2652);
and U3062 (N_3062,N_2561,N_2802);
or U3063 (N_3063,N_2872,N_2863);
or U3064 (N_3064,N_2936,N_2834);
nor U3065 (N_3065,N_2588,N_2774);
nor U3066 (N_3066,N_2780,N_2555);
nor U3067 (N_3067,N_2621,N_2902);
xnor U3068 (N_3068,N_2729,N_2924);
and U3069 (N_3069,N_2784,N_2905);
or U3070 (N_3070,N_2879,N_2509);
nor U3071 (N_3071,N_2628,N_2635);
and U3072 (N_3072,N_2962,N_2560);
xor U3073 (N_3073,N_2612,N_2568);
and U3074 (N_3074,N_2995,N_2644);
nor U3075 (N_3075,N_2760,N_2948);
and U3076 (N_3076,N_2823,N_2975);
nand U3077 (N_3077,N_2672,N_2932);
nand U3078 (N_3078,N_2526,N_2519);
nor U3079 (N_3079,N_2691,N_2753);
or U3080 (N_3080,N_2787,N_2622);
or U3081 (N_3081,N_2548,N_2550);
nor U3082 (N_3082,N_2501,N_2585);
nor U3083 (N_3083,N_2707,N_2954);
or U3084 (N_3084,N_2678,N_2958);
or U3085 (N_3085,N_2609,N_2945);
nor U3086 (N_3086,N_2976,N_2777);
nor U3087 (N_3087,N_2508,N_2812);
nand U3088 (N_3088,N_2647,N_2843);
or U3089 (N_3089,N_2955,N_2803);
nand U3090 (N_3090,N_2629,N_2688);
or U3091 (N_3091,N_2762,N_2979);
xor U3092 (N_3092,N_2748,N_2770);
and U3093 (N_3093,N_2689,N_2655);
and U3094 (N_3094,N_2864,N_2785);
xor U3095 (N_3095,N_2989,N_2910);
and U3096 (N_3096,N_2786,N_2553);
or U3097 (N_3097,N_2999,N_2767);
nor U3098 (N_3098,N_2852,N_2579);
nor U3099 (N_3099,N_2788,N_2677);
xor U3100 (N_3100,N_2875,N_2711);
xnor U3101 (N_3101,N_2790,N_2733);
or U3102 (N_3102,N_2698,N_2952);
and U3103 (N_3103,N_2638,N_2970);
nor U3104 (N_3104,N_2985,N_2653);
xor U3105 (N_3105,N_2791,N_2871);
or U3106 (N_3106,N_2718,N_2904);
and U3107 (N_3107,N_2577,N_2616);
nand U3108 (N_3108,N_2511,N_2929);
or U3109 (N_3109,N_2755,N_2732);
or U3110 (N_3110,N_2706,N_2583);
xnor U3111 (N_3111,N_2751,N_2889);
and U3112 (N_3112,N_2696,N_2589);
nor U3113 (N_3113,N_2513,N_2783);
or U3114 (N_3114,N_2815,N_2725);
nor U3115 (N_3115,N_2811,N_2798);
or U3116 (N_3116,N_2572,N_2938);
nand U3117 (N_3117,N_2942,N_2977);
or U3118 (N_3118,N_2747,N_2634);
nand U3119 (N_3119,N_2849,N_2759);
or U3120 (N_3120,N_2984,N_2933);
and U3121 (N_3121,N_2632,N_2602);
nor U3122 (N_3122,N_2656,N_2500);
and U3123 (N_3123,N_2556,N_2861);
or U3124 (N_3124,N_2745,N_2716);
nor U3125 (N_3125,N_2891,N_2590);
xor U3126 (N_3126,N_2946,N_2885);
and U3127 (N_3127,N_2769,N_2947);
or U3128 (N_3128,N_2643,N_2521);
or U3129 (N_3129,N_2743,N_2883);
nor U3130 (N_3130,N_2744,N_2886);
or U3131 (N_3131,N_2580,N_2700);
and U3132 (N_3132,N_2837,N_2539);
and U3133 (N_3133,N_2876,N_2900);
xor U3134 (N_3134,N_2957,N_2607);
or U3135 (N_3135,N_2913,N_2727);
nor U3136 (N_3136,N_2890,N_2569);
xnor U3137 (N_3137,N_2878,N_2705);
nor U3138 (N_3138,N_2636,N_2827);
nor U3139 (N_3139,N_2771,N_2565);
or U3140 (N_3140,N_2866,N_2828);
or U3141 (N_3141,N_2722,N_2752);
or U3142 (N_3142,N_2779,N_2906);
nor U3143 (N_3143,N_2912,N_2666);
nand U3144 (N_3144,N_2593,N_2950);
and U3145 (N_3145,N_2614,N_2559);
nand U3146 (N_3146,N_2854,N_2639);
or U3147 (N_3147,N_2546,N_2531);
nand U3148 (N_3148,N_2573,N_2567);
nand U3149 (N_3149,N_2838,N_2516);
or U3150 (N_3150,N_2512,N_2514);
and U3151 (N_3151,N_2880,N_2797);
nor U3152 (N_3152,N_2529,N_2735);
xnor U3153 (N_3153,N_2650,N_2726);
nand U3154 (N_3154,N_2564,N_2923);
and U3155 (N_3155,N_2737,N_2734);
or U3156 (N_3156,N_2631,N_2541);
and U3157 (N_3157,N_2600,N_2524);
and U3158 (N_3158,N_2807,N_2829);
nand U3159 (N_3159,N_2536,N_2899);
nor U3160 (N_3160,N_2934,N_2520);
nand U3161 (N_3161,N_2699,N_2540);
or U3162 (N_3162,N_2773,N_2804);
or U3163 (N_3163,N_2964,N_2920);
or U3164 (N_3164,N_2544,N_2627);
and U3165 (N_3165,N_2659,N_2709);
nor U3166 (N_3166,N_2897,N_2967);
nand U3167 (N_3167,N_2789,N_2741);
or U3168 (N_3168,N_2675,N_2965);
or U3169 (N_3169,N_2554,N_2658);
and U3170 (N_3170,N_2930,N_2915);
and U3171 (N_3171,N_2935,N_2620);
nand U3172 (N_3172,N_2679,N_2859);
nand U3173 (N_3173,N_2990,N_2821);
xnor U3174 (N_3174,N_2533,N_2746);
nand U3175 (N_3175,N_2623,N_2858);
nand U3176 (N_3176,N_2617,N_2587);
nand U3177 (N_3177,N_2606,N_2504);
xnor U3178 (N_3178,N_2535,N_2972);
xnor U3179 (N_3179,N_2645,N_2557);
nand U3180 (N_3180,N_2781,N_2613);
nand U3181 (N_3181,N_2867,N_2630);
nand U3182 (N_3182,N_2860,N_2576);
or U3183 (N_3183,N_2793,N_2685);
nand U3184 (N_3184,N_2840,N_2888);
or U3185 (N_3185,N_2832,N_2953);
nand U3186 (N_3186,N_2822,N_2597);
nand U3187 (N_3187,N_2870,N_2959);
and U3188 (N_3188,N_2836,N_2670);
nor U3189 (N_3189,N_2943,N_2674);
nor U3190 (N_3190,N_2928,N_2758);
nand U3191 (N_3191,N_2918,N_2856);
or U3192 (N_3192,N_2549,N_2537);
and U3193 (N_3193,N_2562,N_2850);
nor U3194 (N_3194,N_2584,N_2949);
and U3195 (N_3195,N_2833,N_2673);
nor U3196 (N_3196,N_2592,N_2806);
nor U3197 (N_3197,N_2739,N_2903);
xor U3198 (N_3198,N_2941,N_2701);
nor U3199 (N_3199,N_2817,N_2782);
or U3200 (N_3200,N_2894,N_2682);
nand U3201 (N_3201,N_2917,N_2676);
nand U3202 (N_3202,N_2558,N_2724);
nand U3203 (N_3203,N_2610,N_2712);
xor U3204 (N_3204,N_2916,N_2710);
and U3205 (N_3205,N_2671,N_2982);
or U3206 (N_3206,N_2931,N_2761);
and U3207 (N_3207,N_2996,N_2731);
and U3208 (N_3208,N_2723,N_2756);
nand U3209 (N_3209,N_2846,N_2908);
xnor U3210 (N_3210,N_2694,N_2551);
and U3211 (N_3211,N_2695,N_2591);
nor U3212 (N_3212,N_2687,N_2715);
or U3213 (N_3213,N_2571,N_2839);
nand U3214 (N_3214,N_2775,N_2765);
nand U3215 (N_3215,N_2680,N_2566);
nand U3216 (N_3216,N_2713,N_2778);
xnor U3217 (N_3217,N_2884,N_2869);
and U3218 (N_3218,N_2809,N_2901);
and U3219 (N_3219,N_2518,N_2819);
and U3220 (N_3220,N_2795,N_2974);
nand U3221 (N_3221,N_2575,N_2686);
nand U3222 (N_3222,N_2997,N_2892);
and U3223 (N_3223,N_2764,N_2983);
nand U3224 (N_3224,N_2810,N_2586);
nor U3225 (N_3225,N_2842,N_2547);
xor U3226 (N_3226,N_2563,N_2805);
or U3227 (N_3227,N_2651,N_2502);
nor U3228 (N_3228,N_2693,N_2851);
nor U3229 (N_3229,N_2605,N_2994);
and U3230 (N_3230,N_2966,N_2986);
and U3231 (N_3231,N_2991,N_2719);
nor U3232 (N_3232,N_2507,N_2772);
nor U3233 (N_3233,N_2987,N_2882);
nand U3234 (N_3234,N_2998,N_2857);
nand U3235 (N_3235,N_2720,N_2697);
and U3236 (N_3236,N_2517,N_2522);
and U3237 (N_3237,N_2661,N_2637);
nand U3238 (N_3238,N_2530,N_2898);
or U3239 (N_3239,N_2506,N_2792);
or U3240 (N_3240,N_2847,N_2909);
xor U3241 (N_3241,N_2646,N_2525);
or U3242 (N_3242,N_2578,N_2969);
nor U3243 (N_3243,N_2619,N_2708);
xnor U3244 (N_3244,N_2523,N_2738);
and U3245 (N_3245,N_2657,N_2981);
nor U3246 (N_3246,N_2768,N_2542);
nand U3247 (N_3247,N_2887,N_2625);
nor U3248 (N_3248,N_2640,N_2702);
xnor U3249 (N_3249,N_2721,N_2690);
and U3250 (N_3250,N_2609,N_2991);
nand U3251 (N_3251,N_2759,N_2917);
nand U3252 (N_3252,N_2944,N_2660);
xnor U3253 (N_3253,N_2690,N_2649);
and U3254 (N_3254,N_2610,N_2599);
and U3255 (N_3255,N_2942,N_2983);
nand U3256 (N_3256,N_2771,N_2998);
nand U3257 (N_3257,N_2834,N_2681);
nand U3258 (N_3258,N_2895,N_2964);
and U3259 (N_3259,N_2790,N_2597);
nor U3260 (N_3260,N_2919,N_2841);
nor U3261 (N_3261,N_2835,N_2893);
nor U3262 (N_3262,N_2586,N_2982);
and U3263 (N_3263,N_2914,N_2978);
nor U3264 (N_3264,N_2687,N_2754);
and U3265 (N_3265,N_2922,N_2511);
and U3266 (N_3266,N_2670,N_2840);
xor U3267 (N_3267,N_2800,N_2827);
and U3268 (N_3268,N_2788,N_2569);
nor U3269 (N_3269,N_2924,N_2701);
nand U3270 (N_3270,N_2644,N_2960);
nand U3271 (N_3271,N_2530,N_2891);
nor U3272 (N_3272,N_2793,N_2785);
and U3273 (N_3273,N_2827,N_2860);
and U3274 (N_3274,N_2518,N_2931);
nor U3275 (N_3275,N_2918,N_2910);
nor U3276 (N_3276,N_2730,N_2745);
nand U3277 (N_3277,N_2739,N_2993);
or U3278 (N_3278,N_2581,N_2658);
nor U3279 (N_3279,N_2848,N_2768);
nor U3280 (N_3280,N_2592,N_2793);
nor U3281 (N_3281,N_2658,N_2910);
nand U3282 (N_3282,N_2734,N_2679);
nand U3283 (N_3283,N_2509,N_2773);
and U3284 (N_3284,N_2873,N_2811);
or U3285 (N_3285,N_2938,N_2668);
nor U3286 (N_3286,N_2538,N_2660);
nand U3287 (N_3287,N_2708,N_2958);
or U3288 (N_3288,N_2700,N_2815);
nand U3289 (N_3289,N_2857,N_2696);
xnor U3290 (N_3290,N_2881,N_2629);
and U3291 (N_3291,N_2851,N_2977);
or U3292 (N_3292,N_2765,N_2939);
and U3293 (N_3293,N_2760,N_2649);
and U3294 (N_3294,N_2781,N_2933);
nand U3295 (N_3295,N_2641,N_2952);
nand U3296 (N_3296,N_2691,N_2730);
nand U3297 (N_3297,N_2520,N_2993);
nor U3298 (N_3298,N_2699,N_2653);
and U3299 (N_3299,N_2984,N_2520);
xnor U3300 (N_3300,N_2511,N_2947);
xor U3301 (N_3301,N_2688,N_2512);
or U3302 (N_3302,N_2759,N_2590);
nor U3303 (N_3303,N_2742,N_2599);
nor U3304 (N_3304,N_2677,N_2828);
or U3305 (N_3305,N_2829,N_2689);
nor U3306 (N_3306,N_2982,N_2597);
nand U3307 (N_3307,N_2783,N_2570);
nor U3308 (N_3308,N_2670,N_2729);
or U3309 (N_3309,N_2548,N_2825);
or U3310 (N_3310,N_2678,N_2766);
and U3311 (N_3311,N_2618,N_2997);
nand U3312 (N_3312,N_2882,N_2738);
xnor U3313 (N_3313,N_2547,N_2559);
and U3314 (N_3314,N_2688,N_2866);
nor U3315 (N_3315,N_2715,N_2776);
nand U3316 (N_3316,N_2808,N_2878);
or U3317 (N_3317,N_2677,N_2617);
nor U3318 (N_3318,N_2890,N_2789);
and U3319 (N_3319,N_2931,N_2798);
or U3320 (N_3320,N_2847,N_2697);
nand U3321 (N_3321,N_2582,N_2557);
and U3322 (N_3322,N_2989,N_2868);
and U3323 (N_3323,N_2986,N_2953);
nand U3324 (N_3324,N_2879,N_2521);
and U3325 (N_3325,N_2516,N_2981);
or U3326 (N_3326,N_2629,N_2545);
xor U3327 (N_3327,N_2791,N_2731);
and U3328 (N_3328,N_2783,N_2622);
nor U3329 (N_3329,N_2984,N_2949);
nor U3330 (N_3330,N_2535,N_2668);
nor U3331 (N_3331,N_2763,N_2963);
nor U3332 (N_3332,N_2793,N_2643);
nand U3333 (N_3333,N_2565,N_2718);
nand U3334 (N_3334,N_2570,N_2753);
and U3335 (N_3335,N_2694,N_2814);
and U3336 (N_3336,N_2827,N_2779);
and U3337 (N_3337,N_2900,N_2909);
nor U3338 (N_3338,N_2766,N_2949);
or U3339 (N_3339,N_2964,N_2998);
and U3340 (N_3340,N_2816,N_2507);
nand U3341 (N_3341,N_2789,N_2672);
and U3342 (N_3342,N_2506,N_2870);
and U3343 (N_3343,N_2771,N_2900);
nand U3344 (N_3344,N_2930,N_2829);
nor U3345 (N_3345,N_2953,N_2862);
and U3346 (N_3346,N_2806,N_2932);
nand U3347 (N_3347,N_2726,N_2944);
nor U3348 (N_3348,N_2844,N_2593);
and U3349 (N_3349,N_2949,N_2777);
or U3350 (N_3350,N_2881,N_2645);
or U3351 (N_3351,N_2711,N_2988);
nor U3352 (N_3352,N_2860,N_2552);
and U3353 (N_3353,N_2644,N_2553);
nor U3354 (N_3354,N_2837,N_2508);
or U3355 (N_3355,N_2637,N_2957);
nor U3356 (N_3356,N_2770,N_2615);
and U3357 (N_3357,N_2840,N_2716);
or U3358 (N_3358,N_2678,N_2596);
xnor U3359 (N_3359,N_2658,N_2764);
nand U3360 (N_3360,N_2964,N_2893);
and U3361 (N_3361,N_2687,N_2850);
nor U3362 (N_3362,N_2900,N_2626);
and U3363 (N_3363,N_2776,N_2851);
and U3364 (N_3364,N_2770,N_2773);
nand U3365 (N_3365,N_2715,N_2666);
nand U3366 (N_3366,N_2530,N_2696);
and U3367 (N_3367,N_2781,N_2963);
nand U3368 (N_3368,N_2928,N_2600);
or U3369 (N_3369,N_2911,N_2685);
nand U3370 (N_3370,N_2755,N_2679);
nand U3371 (N_3371,N_2784,N_2972);
or U3372 (N_3372,N_2858,N_2822);
and U3373 (N_3373,N_2864,N_2830);
and U3374 (N_3374,N_2851,N_2579);
and U3375 (N_3375,N_2972,N_2984);
nor U3376 (N_3376,N_2816,N_2619);
nor U3377 (N_3377,N_2946,N_2974);
nand U3378 (N_3378,N_2653,N_2630);
nand U3379 (N_3379,N_2939,N_2822);
nor U3380 (N_3380,N_2896,N_2693);
nor U3381 (N_3381,N_2719,N_2590);
nor U3382 (N_3382,N_2957,N_2923);
nor U3383 (N_3383,N_2903,N_2755);
nand U3384 (N_3384,N_2871,N_2945);
and U3385 (N_3385,N_2925,N_2506);
nand U3386 (N_3386,N_2782,N_2883);
nor U3387 (N_3387,N_2873,N_2601);
nand U3388 (N_3388,N_2797,N_2796);
nor U3389 (N_3389,N_2948,N_2577);
nand U3390 (N_3390,N_2640,N_2884);
xnor U3391 (N_3391,N_2744,N_2870);
or U3392 (N_3392,N_2937,N_2893);
nand U3393 (N_3393,N_2959,N_2982);
or U3394 (N_3394,N_2666,N_2748);
and U3395 (N_3395,N_2842,N_2839);
nor U3396 (N_3396,N_2786,N_2950);
nor U3397 (N_3397,N_2796,N_2906);
and U3398 (N_3398,N_2955,N_2951);
or U3399 (N_3399,N_2689,N_2719);
nand U3400 (N_3400,N_2948,N_2865);
nor U3401 (N_3401,N_2576,N_2623);
and U3402 (N_3402,N_2656,N_2604);
nor U3403 (N_3403,N_2982,N_2546);
or U3404 (N_3404,N_2967,N_2829);
and U3405 (N_3405,N_2819,N_2800);
nand U3406 (N_3406,N_2963,N_2578);
or U3407 (N_3407,N_2565,N_2647);
nand U3408 (N_3408,N_2841,N_2559);
nand U3409 (N_3409,N_2890,N_2810);
nand U3410 (N_3410,N_2834,N_2532);
xnor U3411 (N_3411,N_2979,N_2517);
nor U3412 (N_3412,N_2998,N_2517);
and U3413 (N_3413,N_2622,N_2943);
nor U3414 (N_3414,N_2910,N_2941);
and U3415 (N_3415,N_2693,N_2874);
or U3416 (N_3416,N_2531,N_2836);
nand U3417 (N_3417,N_2946,N_2882);
nor U3418 (N_3418,N_2593,N_2583);
nand U3419 (N_3419,N_2636,N_2756);
nor U3420 (N_3420,N_2517,N_2866);
nand U3421 (N_3421,N_2610,N_2877);
or U3422 (N_3422,N_2939,N_2909);
nor U3423 (N_3423,N_2599,N_2538);
xnor U3424 (N_3424,N_2844,N_2616);
or U3425 (N_3425,N_2721,N_2787);
nand U3426 (N_3426,N_2772,N_2850);
or U3427 (N_3427,N_2618,N_2752);
and U3428 (N_3428,N_2832,N_2544);
or U3429 (N_3429,N_2861,N_2881);
nor U3430 (N_3430,N_2706,N_2986);
xnor U3431 (N_3431,N_2858,N_2719);
or U3432 (N_3432,N_2627,N_2504);
and U3433 (N_3433,N_2774,N_2941);
nor U3434 (N_3434,N_2759,N_2852);
and U3435 (N_3435,N_2678,N_2897);
or U3436 (N_3436,N_2922,N_2549);
nand U3437 (N_3437,N_2522,N_2584);
and U3438 (N_3438,N_2741,N_2505);
nor U3439 (N_3439,N_2622,N_2895);
and U3440 (N_3440,N_2717,N_2566);
nand U3441 (N_3441,N_2977,N_2645);
xor U3442 (N_3442,N_2766,N_2750);
nand U3443 (N_3443,N_2693,N_2950);
nor U3444 (N_3444,N_2644,N_2892);
or U3445 (N_3445,N_2931,N_2552);
nand U3446 (N_3446,N_2887,N_2780);
or U3447 (N_3447,N_2599,N_2835);
xor U3448 (N_3448,N_2549,N_2604);
nand U3449 (N_3449,N_2914,N_2869);
nor U3450 (N_3450,N_2833,N_2630);
or U3451 (N_3451,N_2987,N_2846);
or U3452 (N_3452,N_2983,N_2797);
nor U3453 (N_3453,N_2700,N_2907);
or U3454 (N_3454,N_2959,N_2986);
and U3455 (N_3455,N_2667,N_2681);
or U3456 (N_3456,N_2579,N_2793);
xnor U3457 (N_3457,N_2651,N_2590);
nand U3458 (N_3458,N_2826,N_2865);
or U3459 (N_3459,N_2831,N_2749);
or U3460 (N_3460,N_2872,N_2718);
xor U3461 (N_3461,N_2583,N_2753);
and U3462 (N_3462,N_2558,N_2943);
nor U3463 (N_3463,N_2812,N_2917);
nand U3464 (N_3464,N_2545,N_2774);
nand U3465 (N_3465,N_2604,N_2820);
nand U3466 (N_3466,N_2522,N_2579);
and U3467 (N_3467,N_2711,N_2574);
nor U3468 (N_3468,N_2904,N_2734);
nand U3469 (N_3469,N_2713,N_2945);
xnor U3470 (N_3470,N_2816,N_2879);
xnor U3471 (N_3471,N_2573,N_2796);
nand U3472 (N_3472,N_2690,N_2688);
and U3473 (N_3473,N_2602,N_2972);
nand U3474 (N_3474,N_2785,N_2972);
nor U3475 (N_3475,N_2615,N_2833);
xor U3476 (N_3476,N_2590,N_2781);
nand U3477 (N_3477,N_2538,N_2602);
nand U3478 (N_3478,N_2985,N_2826);
nand U3479 (N_3479,N_2695,N_2946);
nand U3480 (N_3480,N_2667,N_2649);
nor U3481 (N_3481,N_2613,N_2557);
and U3482 (N_3482,N_2804,N_2780);
nor U3483 (N_3483,N_2523,N_2839);
nor U3484 (N_3484,N_2597,N_2857);
nor U3485 (N_3485,N_2670,N_2563);
or U3486 (N_3486,N_2514,N_2797);
xor U3487 (N_3487,N_2788,N_2737);
or U3488 (N_3488,N_2680,N_2650);
or U3489 (N_3489,N_2712,N_2593);
or U3490 (N_3490,N_2872,N_2816);
or U3491 (N_3491,N_2672,N_2683);
nand U3492 (N_3492,N_2759,N_2967);
and U3493 (N_3493,N_2601,N_2737);
or U3494 (N_3494,N_2566,N_2543);
nand U3495 (N_3495,N_2925,N_2891);
or U3496 (N_3496,N_2609,N_2807);
and U3497 (N_3497,N_2980,N_2977);
nand U3498 (N_3498,N_2838,N_2758);
or U3499 (N_3499,N_2655,N_2869);
or U3500 (N_3500,N_3095,N_3372);
and U3501 (N_3501,N_3349,N_3240);
xor U3502 (N_3502,N_3261,N_3435);
nor U3503 (N_3503,N_3439,N_3178);
nand U3504 (N_3504,N_3212,N_3491);
nor U3505 (N_3505,N_3450,N_3025);
and U3506 (N_3506,N_3346,N_3341);
nor U3507 (N_3507,N_3065,N_3404);
or U3508 (N_3508,N_3074,N_3276);
nor U3509 (N_3509,N_3168,N_3344);
xor U3510 (N_3510,N_3174,N_3166);
nand U3511 (N_3511,N_3198,N_3296);
or U3512 (N_3512,N_3078,N_3157);
nor U3513 (N_3513,N_3177,N_3447);
or U3514 (N_3514,N_3154,N_3081);
nor U3515 (N_3515,N_3457,N_3170);
and U3516 (N_3516,N_3121,N_3102);
nand U3517 (N_3517,N_3335,N_3472);
and U3518 (N_3518,N_3229,N_3355);
nor U3519 (N_3519,N_3233,N_3018);
nor U3520 (N_3520,N_3329,N_3131);
xnor U3521 (N_3521,N_3122,N_3399);
and U3522 (N_3522,N_3071,N_3080);
and U3523 (N_3523,N_3182,N_3140);
nor U3524 (N_3524,N_3101,N_3141);
and U3525 (N_3525,N_3211,N_3258);
or U3526 (N_3526,N_3187,N_3361);
and U3527 (N_3527,N_3072,N_3339);
nand U3528 (N_3528,N_3064,N_3208);
nand U3529 (N_3529,N_3228,N_3094);
and U3530 (N_3530,N_3282,N_3167);
nor U3531 (N_3531,N_3186,N_3386);
or U3532 (N_3532,N_3196,N_3285);
nor U3533 (N_3533,N_3482,N_3234);
xnor U3534 (N_3534,N_3437,N_3035);
or U3535 (N_3535,N_3044,N_3043);
nor U3536 (N_3536,N_3469,N_3200);
nand U3537 (N_3537,N_3175,N_3345);
or U3538 (N_3538,N_3327,N_3325);
and U3539 (N_3539,N_3269,N_3366);
xnor U3540 (N_3540,N_3380,N_3295);
nor U3541 (N_3541,N_3231,N_3181);
nor U3542 (N_3542,N_3085,N_3495);
or U3543 (N_3543,N_3287,N_3456);
and U3544 (N_3544,N_3298,N_3426);
nand U3545 (N_3545,N_3489,N_3013);
and U3546 (N_3546,N_3383,N_3308);
nor U3547 (N_3547,N_3148,N_3446);
or U3548 (N_3548,N_3427,N_3352);
xnor U3549 (N_3549,N_3220,N_3125);
or U3550 (N_3550,N_3496,N_3486);
xnor U3551 (N_3551,N_3313,N_3000);
and U3552 (N_3552,N_3307,N_3063);
nand U3553 (N_3553,N_3089,N_3049);
nor U3554 (N_3554,N_3470,N_3090);
and U3555 (N_3555,N_3487,N_3146);
or U3556 (N_3556,N_3418,N_3445);
nor U3557 (N_3557,N_3252,N_3423);
or U3558 (N_3558,N_3387,N_3483);
nor U3559 (N_3559,N_3406,N_3143);
nand U3560 (N_3560,N_3051,N_3218);
and U3561 (N_3561,N_3442,N_3056);
or U3562 (N_3562,N_3020,N_3407);
or U3563 (N_3563,N_3488,N_3398);
or U3564 (N_3564,N_3392,N_3015);
or U3565 (N_3565,N_3249,N_3040);
xnor U3566 (N_3566,N_3328,N_3251);
nor U3567 (N_3567,N_3219,N_3052);
or U3568 (N_3568,N_3476,N_3153);
and U3569 (N_3569,N_3395,N_3410);
or U3570 (N_3570,N_3024,N_3203);
or U3571 (N_3571,N_3343,N_3274);
and U3572 (N_3572,N_3272,N_3379);
and U3573 (N_3573,N_3227,N_3223);
nand U3574 (N_3574,N_3058,N_3191);
nand U3575 (N_3575,N_3422,N_3238);
xor U3576 (N_3576,N_3008,N_3312);
nand U3577 (N_3577,N_3232,N_3265);
and U3578 (N_3578,N_3097,N_3088);
and U3579 (N_3579,N_3351,N_3120);
and U3580 (N_3580,N_3403,N_3443);
nor U3581 (N_3581,N_3452,N_3286);
nand U3582 (N_3582,N_3291,N_3067);
nand U3583 (N_3583,N_3358,N_3019);
or U3584 (N_3584,N_3086,N_3139);
nand U3585 (N_3585,N_3293,N_3050);
nand U3586 (N_3586,N_3250,N_3244);
or U3587 (N_3587,N_3350,N_3388);
nor U3588 (N_3588,N_3205,N_3468);
nor U3589 (N_3589,N_3164,N_3353);
or U3590 (N_3590,N_3448,N_3356);
and U3591 (N_3591,N_3245,N_3033);
or U3592 (N_3592,N_3451,N_3160);
xor U3593 (N_3593,N_3390,N_3192);
xor U3594 (N_3594,N_3173,N_3159);
and U3595 (N_3595,N_3270,N_3068);
and U3596 (N_3596,N_3384,N_3107);
nor U3597 (N_3597,N_3389,N_3059);
nor U3598 (N_3598,N_3204,N_3412);
nor U3599 (N_3599,N_3053,N_3332);
nor U3600 (N_3600,N_3179,N_3303);
nor U3601 (N_3601,N_3340,N_3299);
and U3602 (N_3602,N_3414,N_3010);
or U3603 (N_3603,N_3333,N_3479);
nor U3604 (N_3604,N_3155,N_3188);
or U3605 (N_3605,N_3111,N_3458);
nand U3606 (N_3606,N_3374,N_3243);
nor U3607 (N_3607,N_3171,N_3461);
nor U3608 (N_3608,N_3169,N_3185);
nor U3609 (N_3609,N_3117,N_3342);
or U3610 (N_3610,N_3375,N_3241);
or U3611 (N_3611,N_3042,N_3417);
or U3612 (N_3612,N_3357,N_3324);
nor U3613 (N_3613,N_3454,N_3069);
and U3614 (N_3614,N_3096,N_3256);
or U3615 (N_3615,N_3359,N_3289);
or U3616 (N_3616,N_3093,N_3364);
nand U3617 (N_3617,N_3315,N_3077);
nor U3618 (N_3618,N_3378,N_3278);
and U3619 (N_3619,N_3430,N_3322);
or U3620 (N_3620,N_3263,N_3266);
nor U3621 (N_3621,N_3225,N_3055);
nand U3622 (N_3622,N_3323,N_3429);
xor U3623 (N_3623,N_3401,N_3360);
and U3624 (N_3624,N_3310,N_3376);
and U3625 (N_3625,N_3206,N_3199);
nor U3626 (N_3626,N_3134,N_3076);
or U3627 (N_3627,N_3235,N_3112);
nor U3628 (N_3628,N_3441,N_3129);
nor U3629 (N_3629,N_3029,N_3433);
and U3630 (N_3630,N_3354,N_3115);
and U3631 (N_3631,N_3014,N_3114);
and U3632 (N_3632,N_3498,N_3138);
or U3633 (N_3633,N_3151,N_3474);
nor U3634 (N_3634,N_3124,N_3130);
or U3635 (N_3635,N_3082,N_3041);
nor U3636 (N_3636,N_3434,N_3330);
nor U3637 (N_3637,N_3411,N_3224);
and U3638 (N_3638,N_3247,N_3497);
or U3639 (N_3639,N_3083,N_3464);
nand U3640 (N_3640,N_3316,N_3193);
nor U3641 (N_3641,N_3079,N_3408);
or U3642 (N_3642,N_3126,N_3004);
nand U3643 (N_3643,N_3023,N_3216);
nand U3644 (N_3644,N_3294,N_3163);
nand U3645 (N_3645,N_3254,N_3432);
nand U3646 (N_3646,N_3003,N_3002);
nand U3647 (N_3647,N_3116,N_3336);
nor U3648 (N_3648,N_3222,N_3419);
nor U3649 (N_3649,N_3321,N_3046);
and U3650 (N_3650,N_3136,N_3373);
or U3651 (N_3651,N_3109,N_3475);
nand U3652 (N_3652,N_3363,N_3039);
and U3653 (N_3653,N_3215,N_3156);
nor U3654 (N_3654,N_3075,N_3070);
nand U3655 (N_3655,N_3425,N_3467);
nor U3656 (N_3656,N_3396,N_3260);
and U3657 (N_3657,N_3444,N_3368);
nor U3658 (N_3658,N_3123,N_3133);
or U3659 (N_3659,N_3119,N_3060);
or U3660 (N_3660,N_3214,N_3180);
nand U3661 (N_3661,N_3463,N_3268);
nor U3662 (N_3662,N_3462,N_3239);
and U3663 (N_3663,N_3031,N_3201);
and U3664 (N_3664,N_3012,N_3026);
xor U3665 (N_3665,N_3132,N_3028);
nand U3666 (N_3666,N_3290,N_3326);
and U3667 (N_3667,N_3037,N_3271);
nand U3668 (N_3668,N_3259,N_3370);
nor U3669 (N_3669,N_3103,N_3183);
nand U3670 (N_3670,N_3001,N_3347);
and U3671 (N_3671,N_3011,N_3034);
nand U3672 (N_3672,N_3084,N_3300);
nand U3673 (N_3673,N_3217,N_3455);
nand U3674 (N_3674,N_3453,N_3431);
and U3675 (N_3675,N_3184,N_3213);
or U3676 (N_3676,N_3100,N_3027);
or U3677 (N_3677,N_3098,N_3428);
or U3678 (N_3678,N_3334,N_3253);
or U3679 (N_3679,N_3165,N_3314);
nand U3680 (N_3680,N_3311,N_3402);
or U3681 (N_3681,N_3473,N_3030);
and U3682 (N_3682,N_3409,N_3032);
or U3683 (N_3683,N_3158,N_3162);
xor U3684 (N_3684,N_3485,N_3045);
and U3685 (N_3685,N_3494,N_3391);
nand U3686 (N_3686,N_3304,N_3207);
or U3687 (N_3687,N_3394,N_3492);
and U3688 (N_3688,N_3062,N_3262);
nor U3689 (N_3689,N_3288,N_3194);
nor U3690 (N_3690,N_3365,N_3255);
and U3691 (N_3691,N_3038,N_3318);
xor U3692 (N_3692,N_3230,N_3257);
nor U3693 (N_3693,N_3499,N_3017);
xnor U3694 (N_3694,N_3248,N_3436);
and U3695 (N_3695,N_3277,N_3273);
xor U3696 (N_3696,N_3319,N_3210);
xnor U3697 (N_3697,N_3301,N_3369);
nor U3698 (N_3698,N_3091,N_3061);
xnor U3699 (N_3699,N_3149,N_3221);
nor U3700 (N_3700,N_3275,N_3400);
nor U3701 (N_3701,N_3066,N_3302);
and U3702 (N_3702,N_3281,N_3338);
nand U3703 (N_3703,N_3264,N_3292);
nor U3704 (N_3704,N_3087,N_3137);
xor U3705 (N_3705,N_3128,N_3237);
nand U3706 (N_3706,N_3477,N_3176);
or U3707 (N_3707,N_3110,N_3306);
nand U3708 (N_3708,N_3415,N_3416);
and U3709 (N_3709,N_3144,N_3305);
nor U3710 (N_3710,N_3147,N_3459);
nor U3711 (N_3711,N_3465,N_3279);
and U3712 (N_3712,N_3104,N_3135);
nand U3713 (N_3713,N_3466,N_3284);
nor U3714 (N_3714,N_3007,N_3348);
xor U3715 (N_3715,N_3283,N_3242);
and U3716 (N_3716,N_3421,N_3009);
nor U3717 (N_3717,N_3073,N_3016);
and U3718 (N_3718,N_3118,N_3021);
xnor U3719 (N_3719,N_3189,N_3317);
or U3720 (N_3720,N_3190,N_3484);
and U3721 (N_3721,N_3377,N_3152);
nand U3722 (N_3722,N_3367,N_3054);
nor U3723 (N_3723,N_3106,N_3142);
nor U3724 (N_3724,N_3320,N_3460);
nor U3725 (N_3725,N_3280,N_3385);
nor U3726 (N_3726,N_3362,N_3022);
nand U3727 (N_3727,N_3478,N_3005);
xor U3728 (N_3728,N_3209,N_3297);
or U3729 (N_3729,N_3331,N_3405);
nand U3730 (N_3730,N_3420,N_3337);
and U3731 (N_3731,N_3267,N_3057);
xor U3732 (N_3732,N_3202,N_3197);
nand U3733 (N_3733,N_3449,N_3172);
or U3734 (N_3734,N_3413,N_3490);
nor U3735 (N_3735,N_3006,N_3493);
or U3736 (N_3736,N_3099,N_3161);
or U3737 (N_3737,N_3105,N_3393);
or U3738 (N_3738,N_3150,N_3309);
xnor U3739 (N_3739,N_3424,N_3226);
nand U3740 (N_3740,N_3036,N_3371);
nand U3741 (N_3741,N_3246,N_3236);
nand U3742 (N_3742,N_3047,N_3048);
or U3743 (N_3743,N_3440,N_3438);
and U3744 (N_3744,N_3480,N_3127);
and U3745 (N_3745,N_3113,N_3145);
nor U3746 (N_3746,N_3381,N_3108);
xor U3747 (N_3747,N_3092,N_3481);
nand U3748 (N_3748,N_3471,N_3397);
nand U3749 (N_3749,N_3382,N_3195);
nor U3750 (N_3750,N_3038,N_3158);
nor U3751 (N_3751,N_3055,N_3057);
or U3752 (N_3752,N_3202,N_3237);
or U3753 (N_3753,N_3284,N_3062);
nor U3754 (N_3754,N_3257,N_3446);
or U3755 (N_3755,N_3454,N_3129);
or U3756 (N_3756,N_3104,N_3244);
nor U3757 (N_3757,N_3230,N_3454);
and U3758 (N_3758,N_3244,N_3377);
and U3759 (N_3759,N_3037,N_3371);
nor U3760 (N_3760,N_3225,N_3438);
nand U3761 (N_3761,N_3093,N_3060);
and U3762 (N_3762,N_3307,N_3200);
or U3763 (N_3763,N_3053,N_3136);
nand U3764 (N_3764,N_3470,N_3216);
xor U3765 (N_3765,N_3071,N_3048);
xnor U3766 (N_3766,N_3099,N_3306);
nand U3767 (N_3767,N_3316,N_3074);
xor U3768 (N_3768,N_3044,N_3372);
or U3769 (N_3769,N_3002,N_3347);
or U3770 (N_3770,N_3293,N_3395);
nand U3771 (N_3771,N_3348,N_3222);
xor U3772 (N_3772,N_3422,N_3270);
nand U3773 (N_3773,N_3068,N_3353);
and U3774 (N_3774,N_3254,N_3298);
nand U3775 (N_3775,N_3494,N_3113);
nand U3776 (N_3776,N_3371,N_3281);
or U3777 (N_3777,N_3201,N_3080);
or U3778 (N_3778,N_3312,N_3241);
xnor U3779 (N_3779,N_3099,N_3481);
and U3780 (N_3780,N_3245,N_3340);
and U3781 (N_3781,N_3232,N_3258);
nor U3782 (N_3782,N_3168,N_3395);
nand U3783 (N_3783,N_3299,N_3147);
and U3784 (N_3784,N_3148,N_3423);
nand U3785 (N_3785,N_3193,N_3036);
or U3786 (N_3786,N_3214,N_3081);
or U3787 (N_3787,N_3063,N_3253);
xnor U3788 (N_3788,N_3241,N_3411);
or U3789 (N_3789,N_3081,N_3271);
nand U3790 (N_3790,N_3370,N_3426);
xnor U3791 (N_3791,N_3114,N_3492);
nor U3792 (N_3792,N_3116,N_3488);
nand U3793 (N_3793,N_3252,N_3068);
nor U3794 (N_3794,N_3350,N_3192);
xor U3795 (N_3795,N_3207,N_3341);
and U3796 (N_3796,N_3342,N_3092);
nor U3797 (N_3797,N_3390,N_3480);
or U3798 (N_3798,N_3373,N_3057);
nand U3799 (N_3799,N_3470,N_3237);
nor U3800 (N_3800,N_3193,N_3215);
and U3801 (N_3801,N_3411,N_3110);
and U3802 (N_3802,N_3014,N_3008);
nor U3803 (N_3803,N_3029,N_3470);
and U3804 (N_3804,N_3180,N_3194);
xnor U3805 (N_3805,N_3257,N_3350);
nand U3806 (N_3806,N_3290,N_3129);
xnor U3807 (N_3807,N_3221,N_3477);
and U3808 (N_3808,N_3378,N_3469);
xor U3809 (N_3809,N_3433,N_3038);
or U3810 (N_3810,N_3289,N_3352);
nor U3811 (N_3811,N_3441,N_3432);
and U3812 (N_3812,N_3155,N_3045);
xnor U3813 (N_3813,N_3492,N_3433);
nor U3814 (N_3814,N_3123,N_3157);
or U3815 (N_3815,N_3262,N_3073);
nand U3816 (N_3816,N_3331,N_3321);
nor U3817 (N_3817,N_3205,N_3358);
nand U3818 (N_3818,N_3181,N_3263);
nor U3819 (N_3819,N_3319,N_3395);
nand U3820 (N_3820,N_3008,N_3329);
and U3821 (N_3821,N_3470,N_3211);
nand U3822 (N_3822,N_3091,N_3356);
or U3823 (N_3823,N_3279,N_3071);
xnor U3824 (N_3824,N_3477,N_3154);
xor U3825 (N_3825,N_3227,N_3466);
or U3826 (N_3826,N_3339,N_3488);
or U3827 (N_3827,N_3152,N_3200);
or U3828 (N_3828,N_3155,N_3058);
nor U3829 (N_3829,N_3300,N_3368);
or U3830 (N_3830,N_3428,N_3047);
or U3831 (N_3831,N_3051,N_3415);
nor U3832 (N_3832,N_3235,N_3063);
or U3833 (N_3833,N_3253,N_3266);
nor U3834 (N_3834,N_3397,N_3060);
xnor U3835 (N_3835,N_3363,N_3442);
and U3836 (N_3836,N_3498,N_3238);
nand U3837 (N_3837,N_3228,N_3058);
nor U3838 (N_3838,N_3102,N_3067);
nor U3839 (N_3839,N_3169,N_3494);
nand U3840 (N_3840,N_3392,N_3264);
xor U3841 (N_3841,N_3095,N_3415);
and U3842 (N_3842,N_3169,N_3382);
nor U3843 (N_3843,N_3014,N_3002);
nor U3844 (N_3844,N_3131,N_3465);
nor U3845 (N_3845,N_3061,N_3343);
nor U3846 (N_3846,N_3411,N_3275);
nor U3847 (N_3847,N_3071,N_3146);
or U3848 (N_3848,N_3458,N_3370);
and U3849 (N_3849,N_3281,N_3243);
nor U3850 (N_3850,N_3238,N_3293);
nand U3851 (N_3851,N_3424,N_3361);
nand U3852 (N_3852,N_3367,N_3302);
and U3853 (N_3853,N_3170,N_3000);
and U3854 (N_3854,N_3154,N_3091);
nand U3855 (N_3855,N_3367,N_3487);
and U3856 (N_3856,N_3472,N_3309);
and U3857 (N_3857,N_3193,N_3248);
nand U3858 (N_3858,N_3068,N_3236);
and U3859 (N_3859,N_3235,N_3127);
or U3860 (N_3860,N_3062,N_3116);
or U3861 (N_3861,N_3037,N_3169);
or U3862 (N_3862,N_3401,N_3396);
or U3863 (N_3863,N_3058,N_3156);
or U3864 (N_3864,N_3303,N_3322);
nor U3865 (N_3865,N_3115,N_3160);
nand U3866 (N_3866,N_3251,N_3197);
or U3867 (N_3867,N_3093,N_3463);
and U3868 (N_3868,N_3121,N_3238);
or U3869 (N_3869,N_3149,N_3208);
nor U3870 (N_3870,N_3117,N_3390);
or U3871 (N_3871,N_3128,N_3025);
or U3872 (N_3872,N_3201,N_3194);
nand U3873 (N_3873,N_3434,N_3360);
nand U3874 (N_3874,N_3451,N_3320);
or U3875 (N_3875,N_3305,N_3291);
and U3876 (N_3876,N_3462,N_3335);
nand U3877 (N_3877,N_3029,N_3234);
and U3878 (N_3878,N_3113,N_3337);
nand U3879 (N_3879,N_3049,N_3024);
nand U3880 (N_3880,N_3124,N_3031);
nor U3881 (N_3881,N_3152,N_3084);
xor U3882 (N_3882,N_3282,N_3371);
nor U3883 (N_3883,N_3240,N_3272);
and U3884 (N_3884,N_3046,N_3414);
nor U3885 (N_3885,N_3432,N_3001);
and U3886 (N_3886,N_3363,N_3412);
nand U3887 (N_3887,N_3005,N_3495);
nand U3888 (N_3888,N_3333,N_3278);
nand U3889 (N_3889,N_3419,N_3024);
nor U3890 (N_3890,N_3320,N_3008);
or U3891 (N_3891,N_3269,N_3423);
nand U3892 (N_3892,N_3138,N_3343);
nor U3893 (N_3893,N_3298,N_3189);
nor U3894 (N_3894,N_3419,N_3376);
and U3895 (N_3895,N_3072,N_3314);
nand U3896 (N_3896,N_3476,N_3167);
and U3897 (N_3897,N_3247,N_3441);
and U3898 (N_3898,N_3199,N_3434);
or U3899 (N_3899,N_3028,N_3417);
or U3900 (N_3900,N_3453,N_3233);
nor U3901 (N_3901,N_3451,N_3328);
nand U3902 (N_3902,N_3411,N_3474);
and U3903 (N_3903,N_3362,N_3161);
xnor U3904 (N_3904,N_3012,N_3187);
xor U3905 (N_3905,N_3033,N_3352);
or U3906 (N_3906,N_3390,N_3246);
nor U3907 (N_3907,N_3377,N_3021);
nand U3908 (N_3908,N_3498,N_3124);
or U3909 (N_3909,N_3415,N_3230);
or U3910 (N_3910,N_3076,N_3003);
nor U3911 (N_3911,N_3391,N_3118);
or U3912 (N_3912,N_3206,N_3010);
xnor U3913 (N_3913,N_3399,N_3001);
nand U3914 (N_3914,N_3355,N_3056);
nand U3915 (N_3915,N_3479,N_3290);
nand U3916 (N_3916,N_3066,N_3351);
nand U3917 (N_3917,N_3264,N_3312);
and U3918 (N_3918,N_3048,N_3312);
and U3919 (N_3919,N_3391,N_3178);
nor U3920 (N_3920,N_3488,N_3480);
nor U3921 (N_3921,N_3034,N_3265);
nor U3922 (N_3922,N_3483,N_3437);
nor U3923 (N_3923,N_3179,N_3446);
or U3924 (N_3924,N_3080,N_3209);
nor U3925 (N_3925,N_3498,N_3331);
nand U3926 (N_3926,N_3016,N_3142);
or U3927 (N_3927,N_3146,N_3023);
xnor U3928 (N_3928,N_3304,N_3132);
or U3929 (N_3929,N_3135,N_3172);
nor U3930 (N_3930,N_3093,N_3385);
nand U3931 (N_3931,N_3008,N_3110);
and U3932 (N_3932,N_3086,N_3352);
xnor U3933 (N_3933,N_3408,N_3061);
and U3934 (N_3934,N_3340,N_3119);
and U3935 (N_3935,N_3401,N_3423);
nand U3936 (N_3936,N_3027,N_3486);
nor U3937 (N_3937,N_3028,N_3297);
or U3938 (N_3938,N_3406,N_3418);
and U3939 (N_3939,N_3318,N_3035);
nand U3940 (N_3940,N_3492,N_3072);
nor U3941 (N_3941,N_3012,N_3455);
nor U3942 (N_3942,N_3119,N_3280);
or U3943 (N_3943,N_3221,N_3231);
and U3944 (N_3944,N_3176,N_3072);
or U3945 (N_3945,N_3464,N_3297);
nor U3946 (N_3946,N_3399,N_3087);
and U3947 (N_3947,N_3429,N_3484);
and U3948 (N_3948,N_3478,N_3370);
nor U3949 (N_3949,N_3127,N_3229);
nor U3950 (N_3950,N_3467,N_3358);
and U3951 (N_3951,N_3054,N_3044);
nor U3952 (N_3952,N_3331,N_3210);
nand U3953 (N_3953,N_3370,N_3424);
and U3954 (N_3954,N_3047,N_3320);
and U3955 (N_3955,N_3258,N_3293);
nor U3956 (N_3956,N_3368,N_3468);
or U3957 (N_3957,N_3248,N_3498);
nand U3958 (N_3958,N_3058,N_3174);
or U3959 (N_3959,N_3344,N_3137);
and U3960 (N_3960,N_3031,N_3303);
xor U3961 (N_3961,N_3216,N_3291);
nor U3962 (N_3962,N_3445,N_3043);
xnor U3963 (N_3963,N_3065,N_3136);
and U3964 (N_3964,N_3216,N_3138);
and U3965 (N_3965,N_3287,N_3051);
nand U3966 (N_3966,N_3361,N_3126);
and U3967 (N_3967,N_3381,N_3458);
or U3968 (N_3968,N_3146,N_3155);
nor U3969 (N_3969,N_3392,N_3008);
nor U3970 (N_3970,N_3207,N_3127);
and U3971 (N_3971,N_3332,N_3433);
nand U3972 (N_3972,N_3425,N_3033);
and U3973 (N_3973,N_3453,N_3438);
nand U3974 (N_3974,N_3133,N_3005);
and U3975 (N_3975,N_3366,N_3347);
nor U3976 (N_3976,N_3309,N_3017);
nand U3977 (N_3977,N_3419,N_3385);
and U3978 (N_3978,N_3167,N_3361);
nor U3979 (N_3979,N_3358,N_3473);
or U3980 (N_3980,N_3255,N_3446);
and U3981 (N_3981,N_3202,N_3271);
nand U3982 (N_3982,N_3007,N_3202);
and U3983 (N_3983,N_3459,N_3277);
or U3984 (N_3984,N_3283,N_3289);
nand U3985 (N_3985,N_3470,N_3453);
or U3986 (N_3986,N_3384,N_3469);
nand U3987 (N_3987,N_3283,N_3290);
nor U3988 (N_3988,N_3421,N_3112);
and U3989 (N_3989,N_3367,N_3403);
or U3990 (N_3990,N_3121,N_3096);
and U3991 (N_3991,N_3457,N_3223);
or U3992 (N_3992,N_3012,N_3310);
and U3993 (N_3993,N_3196,N_3022);
nand U3994 (N_3994,N_3267,N_3293);
nor U3995 (N_3995,N_3100,N_3243);
and U3996 (N_3996,N_3234,N_3143);
or U3997 (N_3997,N_3261,N_3438);
nor U3998 (N_3998,N_3102,N_3468);
or U3999 (N_3999,N_3095,N_3098);
nand U4000 (N_4000,N_3937,N_3554);
or U4001 (N_4001,N_3650,N_3998);
xnor U4002 (N_4002,N_3673,N_3785);
nand U4003 (N_4003,N_3832,N_3806);
or U4004 (N_4004,N_3798,N_3863);
and U4005 (N_4005,N_3507,N_3997);
xnor U4006 (N_4006,N_3957,N_3787);
nand U4007 (N_4007,N_3663,N_3769);
or U4008 (N_4008,N_3774,N_3909);
nor U4009 (N_4009,N_3784,N_3600);
nand U4010 (N_4010,N_3963,N_3604);
nor U4011 (N_4011,N_3585,N_3760);
and U4012 (N_4012,N_3599,N_3685);
nor U4013 (N_4013,N_3880,N_3964);
xnor U4014 (N_4014,N_3775,N_3879);
nor U4015 (N_4015,N_3830,N_3906);
or U4016 (N_4016,N_3613,N_3645);
nor U4017 (N_4017,N_3624,N_3897);
nor U4018 (N_4018,N_3522,N_3958);
and U4019 (N_4019,N_3719,N_3690);
xnor U4020 (N_4020,N_3709,N_3623);
or U4021 (N_4021,N_3628,N_3900);
nor U4022 (N_4022,N_3710,N_3676);
nand U4023 (N_4023,N_3705,N_3500);
and U4024 (N_4024,N_3682,N_3873);
nor U4025 (N_4025,N_3751,N_3727);
nand U4026 (N_4026,N_3702,N_3947);
nor U4027 (N_4027,N_3892,N_3874);
and U4028 (N_4028,N_3872,N_3923);
xor U4029 (N_4029,N_3890,N_3514);
nor U4030 (N_4030,N_3856,N_3807);
and U4031 (N_4031,N_3548,N_3840);
or U4032 (N_4032,N_3951,N_3869);
xor U4033 (N_4033,N_3992,N_3936);
nor U4034 (N_4034,N_3694,N_3731);
and U4035 (N_4035,N_3979,N_3509);
or U4036 (N_4036,N_3805,N_3552);
nand U4037 (N_4037,N_3648,N_3859);
nor U4038 (N_4038,N_3758,N_3582);
nand U4039 (N_4039,N_3962,N_3686);
nand U4040 (N_4040,N_3955,N_3542);
or U4041 (N_4041,N_3596,N_3788);
and U4042 (N_4042,N_3521,N_3938);
or U4043 (N_4043,N_3864,N_3952);
nand U4044 (N_4044,N_3529,N_3825);
or U4045 (N_4045,N_3671,N_3611);
nor U4046 (N_4046,N_3954,N_3925);
or U4047 (N_4047,N_3844,N_3752);
nand U4048 (N_4048,N_3738,N_3630);
and U4049 (N_4049,N_3818,N_3723);
nand U4050 (N_4050,N_3586,N_3767);
and U4051 (N_4051,N_3689,N_3516);
nor U4052 (N_4052,N_3991,N_3770);
nand U4053 (N_4053,N_3989,N_3993);
nor U4054 (N_4054,N_3720,N_3640);
nand U4055 (N_4055,N_3974,N_3776);
xor U4056 (N_4056,N_3627,N_3933);
nand U4057 (N_4057,N_3766,N_3660);
xnor U4058 (N_4058,N_3916,N_3817);
or U4059 (N_4059,N_3948,N_3986);
or U4060 (N_4060,N_3753,N_3826);
xnor U4061 (N_4061,N_3644,N_3846);
or U4062 (N_4062,N_3754,N_3943);
xor U4063 (N_4063,N_3764,N_3677);
nand U4064 (N_4064,N_3625,N_3654);
nor U4065 (N_4065,N_3917,N_3949);
nand U4066 (N_4066,N_3990,N_3519);
nand U4067 (N_4067,N_3961,N_3575);
or U4068 (N_4068,N_3960,N_3935);
nor U4069 (N_4069,N_3852,N_3994);
and U4070 (N_4070,N_3574,N_3668);
xnor U4071 (N_4071,N_3884,N_3814);
and U4072 (N_4072,N_3584,N_3978);
nand U4073 (N_4073,N_3816,N_3861);
and U4074 (N_4074,N_3571,N_3740);
xor U4075 (N_4075,N_3793,N_3576);
nand U4076 (N_4076,N_3748,N_3970);
nand U4077 (N_4077,N_3794,N_3587);
and U4078 (N_4078,N_3837,N_3609);
xnor U4079 (N_4079,N_3711,N_3842);
or U4080 (N_4080,N_3946,N_3866);
xnor U4081 (N_4081,N_3715,N_3637);
and U4082 (N_4082,N_3579,N_3749);
and U4083 (N_4083,N_3792,N_3786);
nand U4084 (N_4084,N_3534,N_3595);
and U4085 (N_4085,N_3667,N_3821);
nor U4086 (N_4086,N_3583,N_3718);
and U4087 (N_4087,N_3911,N_3893);
or U4088 (N_4088,N_3691,N_3982);
xnor U4089 (N_4089,N_3539,N_3606);
nor U4090 (N_4090,N_3607,N_3578);
and U4091 (N_4091,N_3891,N_3959);
xnor U4092 (N_4092,N_3932,N_3547);
and U4093 (N_4093,N_3987,N_3950);
or U4094 (N_4094,N_3590,N_3795);
and U4095 (N_4095,N_3887,N_3546);
and U4096 (N_4096,N_3977,N_3618);
nand U4097 (N_4097,N_3538,N_3940);
and U4098 (N_4098,N_3915,N_3652);
nor U4099 (N_4099,N_3898,N_3918);
nor U4100 (N_4100,N_3980,N_3706);
nand U4101 (N_4101,N_3803,N_3865);
nor U4102 (N_4102,N_3850,N_3531);
nand U4103 (N_4103,N_3843,N_3616);
nand U4104 (N_4104,N_3881,N_3501);
nor U4105 (N_4105,N_3800,N_3867);
or U4106 (N_4106,N_3526,N_3908);
nand U4107 (N_4107,N_3765,N_3988);
nor U4108 (N_4108,N_3976,N_3510);
and U4109 (N_4109,N_3780,N_3502);
or U4110 (N_4110,N_3756,N_3612);
and U4111 (N_4111,N_3561,N_3833);
nand U4112 (N_4112,N_3828,N_3601);
nor U4113 (N_4113,N_3617,N_3907);
nand U4114 (N_4114,N_3801,N_3506);
nand U4115 (N_4115,N_3570,N_3781);
and U4116 (N_4116,N_3675,N_3921);
and U4117 (N_4117,N_3762,N_3944);
nor U4118 (N_4118,N_3820,N_3678);
nand U4119 (N_4119,N_3920,N_3855);
and U4120 (N_4120,N_3562,N_3773);
xnor U4121 (N_4121,N_3995,N_3631);
or U4122 (N_4122,N_3537,N_3975);
nor U4123 (N_4123,N_3520,N_3504);
and U4124 (N_4124,N_3905,N_3602);
nor U4125 (N_4125,N_3622,N_3722);
nand U4126 (N_4126,N_3877,N_3741);
and U4127 (N_4127,N_3849,N_3638);
nor U4128 (N_4128,N_3589,N_3730);
or U4129 (N_4129,N_3704,N_3896);
xnor U4130 (N_4130,N_3902,N_3608);
or U4131 (N_4131,N_3953,N_3544);
and U4132 (N_4132,N_3512,N_3680);
or U4133 (N_4133,N_3610,N_3941);
xor U4134 (N_4134,N_3838,N_3692);
or U4135 (N_4135,N_3559,N_3634);
nor U4136 (N_4136,N_3672,N_3647);
and U4137 (N_4137,N_3513,N_3746);
nor U4138 (N_4138,N_3808,N_3942);
nor U4139 (N_4139,N_3854,N_3687);
and U4140 (N_4140,N_3525,N_3824);
or U4141 (N_4141,N_3603,N_3588);
or U4142 (N_4142,N_3656,N_3569);
xor U4143 (N_4143,N_3763,N_3666);
nand U4144 (N_4144,N_3708,N_3904);
or U4145 (N_4145,N_3858,N_3665);
nand U4146 (N_4146,N_3528,N_3910);
nor U4147 (N_4147,N_3733,N_3927);
or U4148 (N_4148,N_3836,N_3819);
nor U4149 (N_4149,N_3553,N_3919);
or U4150 (N_4150,N_3924,N_3659);
nand U4151 (N_4151,N_3939,N_3649);
and U4152 (N_4152,N_3655,N_3593);
and U4153 (N_4153,N_3984,N_3533);
and U4154 (N_4154,N_3750,N_3619);
nor U4155 (N_4155,N_3956,N_3688);
nand U4156 (N_4156,N_3577,N_3851);
or U4157 (N_4157,N_3965,N_3875);
nand U4158 (N_4158,N_3620,N_3658);
nand U4159 (N_4159,N_3834,N_3888);
and U4160 (N_4160,N_3983,N_3564);
or U4161 (N_4161,N_3563,N_3968);
nor U4162 (N_4162,N_3703,N_3789);
and U4163 (N_4163,N_3515,N_3532);
nor U4164 (N_4164,N_3772,N_3653);
nand U4165 (N_4165,N_3717,N_3527);
nand U4166 (N_4166,N_3996,N_3549);
or U4167 (N_4167,N_3973,N_3699);
and U4168 (N_4168,N_3629,N_3848);
nand U4169 (N_4169,N_3886,N_3860);
nor U4170 (N_4170,N_3934,N_3580);
nand U4171 (N_4171,N_3812,N_3729);
and U4172 (N_4172,N_3728,N_3759);
or U4173 (N_4173,N_3573,N_3822);
nor U4174 (N_4174,N_3734,N_3868);
nand U4175 (N_4175,N_3566,N_3966);
nor U4176 (N_4176,N_3701,N_3945);
nand U4177 (N_4177,N_3598,N_3591);
xor U4178 (N_4178,N_3739,N_3661);
xor U4179 (N_4179,N_3930,N_3985);
nor U4180 (N_4180,N_3804,N_3810);
nor U4181 (N_4181,N_3929,N_3724);
nor U4182 (N_4182,N_3894,N_3845);
or U4183 (N_4183,N_3732,N_3736);
nand U4184 (N_4184,N_3827,N_3523);
or U4185 (N_4185,N_3568,N_3922);
nor U4186 (N_4186,N_3878,N_3565);
xor U4187 (N_4187,N_3857,N_3913);
or U4188 (N_4188,N_3742,N_3597);
xnor U4189 (N_4189,N_3777,N_3518);
or U4190 (N_4190,N_3714,N_3581);
and U4191 (N_4191,N_3768,N_3883);
nand U4192 (N_4192,N_3725,N_3664);
nand U4193 (N_4193,N_3971,N_3651);
or U4194 (N_4194,N_3572,N_3707);
and U4195 (N_4195,N_3761,N_3882);
or U4196 (N_4196,N_3558,N_3981);
or U4197 (N_4197,N_3632,N_3684);
or U4198 (N_4198,N_3614,N_3605);
and U4199 (N_4199,N_3639,N_3551);
or U4200 (N_4200,N_3594,N_3726);
and U4201 (N_4201,N_3835,N_3779);
and U4202 (N_4202,N_3670,N_3643);
and U4203 (N_4203,N_3969,N_3626);
nor U4204 (N_4204,N_3926,N_3536);
nor U4205 (N_4205,N_3791,N_3592);
nand U4206 (N_4206,N_3555,N_3782);
and U4207 (N_4207,N_3799,N_3901);
nor U4208 (N_4208,N_3889,N_3674);
or U4209 (N_4209,N_3876,N_3839);
and U4210 (N_4210,N_3811,N_3560);
or U4211 (N_4211,N_3831,N_3641);
or U4212 (N_4212,N_3735,N_3517);
nand U4213 (N_4213,N_3669,N_3737);
or U4214 (N_4214,N_3870,N_3567);
or U4215 (N_4215,N_3899,N_3615);
or U4216 (N_4216,N_3545,N_3895);
nand U4217 (N_4217,N_3871,N_3796);
nand U4218 (N_4218,N_3928,N_3642);
or U4219 (N_4219,N_3550,N_3695);
or U4220 (N_4220,N_3681,N_3530);
nor U4221 (N_4221,N_3967,N_3679);
xor U4222 (N_4222,N_3716,N_3797);
or U4223 (N_4223,N_3743,N_3721);
and U4224 (N_4224,N_3541,N_3621);
and U4225 (N_4225,N_3757,N_3885);
and U4226 (N_4226,N_3557,N_3696);
nor U4227 (N_4227,N_3503,N_3698);
nand U4228 (N_4228,N_3809,N_3511);
nand U4229 (N_4229,N_3931,N_3771);
nor U4230 (N_4230,N_3853,N_3744);
nand U4231 (N_4231,N_3829,N_3543);
xor U4232 (N_4232,N_3633,N_3662);
and U4233 (N_4233,N_3700,N_3813);
or U4234 (N_4234,N_3841,N_3999);
or U4235 (N_4235,N_3505,N_3508);
nand U4236 (N_4236,N_3657,N_3745);
xnor U4237 (N_4237,N_3697,N_3683);
and U4238 (N_4238,N_3862,N_3636);
and U4239 (N_4239,N_3747,N_3903);
nor U4240 (N_4240,N_3972,N_3524);
and U4241 (N_4241,N_3693,N_3646);
nand U4242 (N_4242,N_3635,N_3783);
xor U4243 (N_4243,N_3540,N_3914);
xnor U4244 (N_4244,N_3755,N_3815);
and U4245 (N_4245,N_3912,N_3713);
nand U4246 (N_4246,N_3802,N_3556);
xor U4247 (N_4247,N_3535,N_3790);
and U4248 (N_4248,N_3778,N_3847);
xor U4249 (N_4249,N_3823,N_3712);
and U4250 (N_4250,N_3928,N_3616);
or U4251 (N_4251,N_3613,N_3971);
nand U4252 (N_4252,N_3531,N_3628);
and U4253 (N_4253,N_3934,N_3902);
nor U4254 (N_4254,N_3709,N_3586);
and U4255 (N_4255,N_3842,N_3791);
and U4256 (N_4256,N_3661,N_3727);
nor U4257 (N_4257,N_3848,N_3705);
nand U4258 (N_4258,N_3582,N_3599);
nand U4259 (N_4259,N_3705,N_3658);
nand U4260 (N_4260,N_3571,N_3710);
and U4261 (N_4261,N_3906,N_3614);
and U4262 (N_4262,N_3850,N_3854);
or U4263 (N_4263,N_3967,N_3924);
xnor U4264 (N_4264,N_3657,N_3637);
nand U4265 (N_4265,N_3838,N_3904);
or U4266 (N_4266,N_3551,N_3788);
nor U4267 (N_4267,N_3946,N_3947);
xnor U4268 (N_4268,N_3924,N_3926);
nor U4269 (N_4269,N_3906,N_3665);
or U4270 (N_4270,N_3796,N_3625);
nand U4271 (N_4271,N_3527,N_3568);
nand U4272 (N_4272,N_3547,N_3971);
nand U4273 (N_4273,N_3768,N_3830);
and U4274 (N_4274,N_3865,N_3561);
nor U4275 (N_4275,N_3961,N_3972);
and U4276 (N_4276,N_3742,N_3805);
nor U4277 (N_4277,N_3563,N_3823);
nor U4278 (N_4278,N_3594,N_3792);
xor U4279 (N_4279,N_3964,N_3532);
nand U4280 (N_4280,N_3948,N_3526);
nor U4281 (N_4281,N_3698,N_3924);
nand U4282 (N_4282,N_3968,N_3599);
nand U4283 (N_4283,N_3632,N_3668);
nand U4284 (N_4284,N_3685,N_3738);
or U4285 (N_4285,N_3636,N_3631);
nand U4286 (N_4286,N_3902,N_3730);
and U4287 (N_4287,N_3606,N_3868);
nor U4288 (N_4288,N_3804,N_3559);
nand U4289 (N_4289,N_3620,N_3524);
and U4290 (N_4290,N_3514,N_3889);
and U4291 (N_4291,N_3775,N_3568);
nor U4292 (N_4292,N_3533,N_3510);
or U4293 (N_4293,N_3945,N_3912);
nand U4294 (N_4294,N_3720,N_3991);
nor U4295 (N_4295,N_3646,N_3546);
and U4296 (N_4296,N_3917,N_3698);
or U4297 (N_4297,N_3615,N_3779);
xor U4298 (N_4298,N_3710,N_3947);
or U4299 (N_4299,N_3877,N_3798);
and U4300 (N_4300,N_3795,N_3909);
nor U4301 (N_4301,N_3935,N_3809);
xnor U4302 (N_4302,N_3830,N_3684);
and U4303 (N_4303,N_3788,N_3872);
nand U4304 (N_4304,N_3734,N_3599);
and U4305 (N_4305,N_3950,N_3967);
xor U4306 (N_4306,N_3988,N_3922);
or U4307 (N_4307,N_3639,N_3772);
and U4308 (N_4308,N_3502,N_3651);
and U4309 (N_4309,N_3912,N_3582);
xor U4310 (N_4310,N_3932,N_3701);
or U4311 (N_4311,N_3577,N_3876);
or U4312 (N_4312,N_3506,N_3527);
nor U4313 (N_4313,N_3903,N_3720);
xor U4314 (N_4314,N_3852,N_3678);
nor U4315 (N_4315,N_3704,N_3508);
nand U4316 (N_4316,N_3884,N_3837);
or U4317 (N_4317,N_3588,N_3880);
xnor U4318 (N_4318,N_3877,N_3774);
and U4319 (N_4319,N_3517,N_3786);
or U4320 (N_4320,N_3666,N_3768);
nand U4321 (N_4321,N_3543,N_3572);
nor U4322 (N_4322,N_3810,N_3901);
and U4323 (N_4323,N_3557,N_3888);
nand U4324 (N_4324,N_3942,N_3835);
nor U4325 (N_4325,N_3567,N_3882);
nor U4326 (N_4326,N_3897,N_3620);
xor U4327 (N_4327,N_3969,N_3654);
nand U4328 (N_4328,N_3835,N_3510);
nand U4329 (N_4329,N_3761,N_3560);
nand U4330 (N_4330,N_3706,N_3943);
or U4331 (N_4331,N_3672,N_3870);
and U4332 (N_4332,N_3696,N_3566);
and U4333 (N_4333,N_3810,N_3982);
nand U4334 (N_4334,N_3821,N_3968);
nor U4335 (N_4335,N_3883,N_3857);
and U4336 (N_4336,N_3926,N_3662);
nor U4337 (N_4337,N_3754,N_3831);
nor U4338 (N_4338,N_3595,N_3845);
and U4339 (N_4339,N_3825,N_3573);
nor U4340 (N_4340,N_3587,N_3834);
xnor U4341 (N_4341,N_3887,N_3924);
nor U4342 (N_4342,N_3531,N_3664);
nor U4343 (N_4343,N_3955,N_3726);
nor U4344 (N_4344,N_3744,N_3835);
or U4345 (N_4345,N_3563,N_3961);
xnor U4346 (N_4346,N_3864,N_3795);
and U4347 (N_4347,N_3665,N_3840);
nand U4348 (N_4348,N_3545,N_3800);
and U4349 (N_4349,N_3580,N_3548);
nor U4350 (N_4350,N_3602,N_3962);
nand U4351 (N_4351,N_3684,N_3658);
nand U4352 (N_4352,N_3682,N_3985);
or U4353 (N_4353,N_3921,N_3661);
nand U4354 (N_4354,N_3507,N_3639);
nor U4355 (N_4355,N_3643,N_3960);
or U4356 (N_4356,N_3591,N_3800);
or U4357 (N_4357,N_3933,N_3636);
nand U4358 (N_4358,N_3954,N_3661);
and U4359 (N_4359,N_3942,N_3794);
nor U4360 (N_4360,N_3571,N_3654);
and U4361 (N_4361,N_3533,N_3874);
and U4362 (N_4362,N_3991,N_3865);
or U4363 (N_4363,N_3977,N_3837);
or U4364 (N_4364,N_3960,N_3986);
and U4365 (N_4365,N_3598,N_3695);
xor U4366 (N_4366,N_3582,N_3553);
or U4367 (N_4367,N_3656,N_3954);
and U4368 (N_4368,N_3690,N_3663);
xnor U4369 (N_4369,N_3914,N_3547);
nor U4370 (N_4370,N_3516,N_3752);
or U4371 (N_4371,N_3899,N_3656);
nor U4372 (N_4372,N_3588,N_3971);
or U4373 (N_4373,N_3959,N_3510);
or U4374 (N_4374,N_3566,N_3699);
nand U4375 (N_4375,N_3535,N_3636);
and U4376 (N_4376,N_3757,N_3830);
nand U4377 (N_4377,N_3895,N_3743);
nand U4378 (N_4378,N_3987,N_3526);
nor U4379 (N_4379,N_3942,N_3960);
and U4380 (N_4380,N_3526,N_3761);
nor U4381 (N_4381,N_3816,N_3959);
xor U4382 (N_4382,N_3673,N_3712);
and U4383 (N_4383,N_3590,N_3905);
or U4384 (N_4384,N_3812,N_3559);
or U4385 (N_4385,N_3705,N_3739);
nor U4386 (N_4386,N_3524,N_3970);
or U4387 (N_4387,N_3842,N_3885);
and U4388 (N_4388,N_3897,N_3832);
or U4389 (N_4389,N_3582,N_3940);
nor U4390 (N_4390,N_3870,N_3613);
nand U4391 (N_4391,N_3696,N_3861);
nor U4392 (N_4392,N_3806,N_3650);
and U4393 (N_4393,N_3761,N_3710);
xnor U4394 (N_4394,N_3877,N_3949);
nand U4395 (N_4395,N_3580,N_3918);
nor U4396 (N_4396,N_3830,N_3836);
or U4397 (N_4397,N_3770,N_3743);
nor U4398 (N_4398,N_3693,N_3618);
or U4399 (N_4399,N_3724,N_3676);
or U4400 (N_4400,N_3544,N_3894);
and U4401 (N_4401,N_3925,N_3842);
and U4402 (N_4402,N_3737,N_3820);
and U4403 (N_4403,N_3817,N_3733);
or U4404 (N_4404,N_3762,N_3812);
or U4405 (N_4405,N_3679,N_3917);
or U4406 (N_4406,N_3745,N_3715);
nand U4407 (N_4407,N_3646,N_3865);
nand U4408 (N_4408,N_3783,N_3845);
nand U4409 (N_4409,N_3978,N_3755);
nand U4410 (N_4410,N_3624,N_3918);
or U4411 (N_4411,N_3502,N_3686);
or U4412 (N_4412,N_3771,N_3909);
nand U4413 (N_4413,N_3888,N_3501);
and U4414 (N_4414,N_3752,N_3724);
nand U4415 (N_4415,N_3638,N_3725);
nand U4416 (N_4416,N_3660,N_3829);
and U4417 (N_4417,N_3669,N_3846);
and U4418 (N_4418,N_3785,N_3928);
or U4419 (N_4419,N_3618,N_3513);
or U4420 (N_4420,N_3953,N_3552);
or U4421 (N_4421,N_3771,N_3594);
nand U4422 (N_4422,N_3672,N_3969);
nand U4423 (N_4423,N_3846,N_3724);
nand U4424 (N_4424,N_3537,N_3719);
nand U4425 (N_4425,N_3954,N_3975);
or U4426 (N_4426,N_3714,N_3944);
nand U4427 (N_4427,N_3996,N_3674);
nand U4428 (N_4428,N_3706,N_3553);
and U4429 (N_4429,N_3673,N_3566);
nand U4430 (N_4430,N_3707,N_3556);
or U4431 (N_4431,N_3585,N_3658);
nand U4432 (N_4432,N_3602,N_3875);
nor U4433 (N_4433,N_3608,N_3732);
and U4434 (N_4434,N_3693,N_3629);
nor U4435 (N_4435,N_3689,N_3782);
xor U4436 (N_4436,N_3795,N_3509);
or U4437 (N_4437,N_3553,N_3849);
nand U4438 (N_4438,N_3683,N_3749);
and U4439 (N_4439,N_3520,N_3963);
and U4440 (N_4440,N_3910,N_3787);
nor U4441 (N_4441,N_3724,N_3961);
and U4442 (N_4442,N_3914,N_3517);
and U4443 (N_4443,N_3632,N_3945);
nor U4444 (N_4444,N_3503,N_3733);
nand U4445 (N_4445,N_3564,N_3923);
or U4446 (N_4446,N_3693,N_3663);
nand U4447 (N_4447,N_3696,N_3606);
or U4448 (N_4448,N_3878,N_3943);
xor U4449 (N_4449,N_3510,N_3871);
nor U4450 (N_4450,N_3793,N_3932);
xnor U4451 (N_4451,N_3574,N_3661);
and U4452 (N_4452,N_3737,N_3678);
nor U4453 (N_4453,N_3534,N_3801);
nor U4454 (N_4454,N_3655,N_3801);
xnor U4455 (N_4455,N_3867,N_3604);
nand U4456 (N_4456,N_3884,N_3941);
nand U4457 (N_4457,N_3692,N_3954);
nor U4458 (N_4458,N_3831,N_3867);
nand U4459 (N_4459,N_3809,N_3701);
nand U4460 (N_4460,N_3708,N_3617);
and U4461 (N_4461,N_3533,N_3937);
nor U4462 (N_4462,N_3909,N_3856);
nor U4463 (N_4463,N_3885,N_3658);
and U4464 (N_4464,N_3637,N_3690);
nand U4465 (N_4465,N_3531,N_3837);
and U4466 (N_4466,N_3718,N_3952);
or U4467 (N_4467,N_3582,N_3768);
or U4468 (N_4468,N_3962,N_3863);
nand U4469 (N_4469,N_3868,N_3532);
nand U4470 (N_4470,N_3575,N_3594);
xor U4471 (N_4471,N_3892,N_3727);
and U4472 (N_4472,N_3985,N_3573);
or U4473 (N_4473,N_3857,N_3965);
nand U4474 (N_4474,N_3677,N_3755);
nand U4475 (N_4475,N_3870,N_3822);
xor U4476 (N_4476,N_3824,N_3760);
and U4477 (N_4477,N_3890,N_3920);
and U4478 (N_4478,N_3817,N_3598);
xnor U4479 (N_4479,N_3780,N_3874);
and U4480 (N_4480,N_3531,N_3824);
or U4481 (N_4481,N_3534,N_3719);
xnor U4482 (N_4482,N_3717,N_3833);
nand U4483 (N_4483,N_3864,N_3676);
and U4484 (N_4484,N_3850,N_3673);
xor U4485 (N_4485,N_3928,N_3843);
nand U4486 (N_4486,N_3590,N_3745);
or U4487 (N_4487,N_3995,N_3959);
xor U4488 (N_4488,N_3668,N_3757);
or U4489 (N_4489,N_3806,N_3667);
or U4490 (N_4490,N_3831,N_3608);
nand U4491 (N_4491,N_3666,N_3936);
or U4492 (N_4492,N_3600,N_3914);
nor U4493 (N_4493,N_3830,N_3558);
and U4494 (N_4494,N_3919,N_3722);
nor U4495 (N_4495,N_3936,N_3676);
nand U4496 (N_4496,N_3852,N_3855);
or U4497 (N_4497,N_3672,N_3686);
or U4498 (N_4498,N_3600,N_3707);
and U4499 (N_4499,N_3881,N_3926);
or U4500 (N_4500,N_4326,N_4283);
or U4501 (N_4501,N_4376,N_4112);
xnor U4502 (N_4502,N_4397,N_4205);
nor U4503 (N_4503,N_4477,N_4480);
and U4504 (N_4504,N_4104,N_4476);
and U4505 (N_4505,N_4304,N_4448);
or U4506 (N_4506,N_4415,N_4273);
nor U4507 (N_4507,N_4022,N_4206);
xnor U4508 (N_4508,N_4243,N_4497);
or U4509 (N_4509,N_4481,N_4096);
or U4510 (N_4510,N_4435,N_4229);
nor U4511 (N_4511,N_4340,N_4043);
and U4512 (N_4512,N_4218,N_4475);
nand U4513 (N_4513,N_4157,N_4212);
nand U4514 (N_4514,N_4001,N_4027);
or U4515 (N_4515,N_4299,N_4482);
or U4516 (N_4516,N_4225,N_4441);
nor U4517 (N_4517,N_4343,N_4199);
or U4518 (N_4518,N_4172,N_4436);
nor U4519 (N_4519,N_4169,N_4339);
and U4520 (N_4520,N_4242,N_4453);
nor U4521 (N_4521,N_4041,N_4018);
nor U4522 (N_4522,N_4325,N_4191);
or U4523 (N_4523,N_4222,N_4474);
and U4524 (N_4524,N_4345,N_4364);
nor U4525 (N_4525,N_4236,N_4454);
or U4526 (N_4526,N_4073,N_4368);
and U4527 (N_4527,N_4449,N_4267);
or U4528 (N_4528,N_4126,N_4342);
or U4529 (N_4529,N_4045,N_4127);
or U4530 (N_4530,N_4058,N_4496);
and U4531 (N_4531,N_4113,N_4327);
nand U4532 (N_4532,N_4274,N_4303);
or U4533 (N_4533,N_4386,N_4285);
or U4534 (N_4534,N_4166,N_4296);
or U4535 (N_4535,N_4445,N_4450);
and U4536 (N_4536,N_4403,N_4138);
xnor U4537 (N_4537,N_4300,N_4451);
and U4538 (N_4538,N_4470,N_4056);
nand U4539 (N_4539,N_4133,N_4163);
and U4540 (N_4540,N_4484,N_4239);
or U4541 (N_4541,N_4069,N_4434);
and U4542 (N_4542,N_4038,N_4311);
nor U4543 (N_4543,N_4263,N_4430);
nand U4544 (N_4544,N_4298,N_4004);
xnor U4545 (N_4545,N_4100,N_4356);
or U4546 (N_4546,N_4357,N_4131);
nor U4547 (N_4547,N_4396,N_4091);
xnor U4548 (N_4548,N_4193,N_4071);
nor U4549 (N_4549,N_4125,N_4361);
or U4550 (N_4550,N_4329,N_4366);
or U4551 (N_4551,N_4249,N_4068);
nand U4552 (N_4552,N_4044,N_4110);
and U4553 (N_4553,N_4008,N_4197);
nand U4554 (N_4554,N_4287,N_4078);
xnor U4555 (N_4555,N_4432,N_4232);
nand U4556 (N_4556,N_4036,N_4035);
and U4557 (N_4557,N_4101,N_4455);
and U4558 (N_4558,N_4049,N_4135);
nor U4559 (N_4559,N_4377,N_4442);
nor U4560 (N_4560,N_4016,N_4116);
and U4561 (N_4561,N_4148,N_4405);
xor U4562 (N_4562,N_4334,N_4065);
nor U4563 (N_4563,N_4379,N_4279);
and U4564 (N_4564,N_4362,N_4266);
and U4565 (N_4565,N_4227,N_4170);
nand U4566 (N_4566,N_4105,N_4438);
nand U4567 (N_4567,N_4444,N_4021);
nand U4568 (N_4568,N_4276,N_4050);
nand U4569 (N_4569,N_4416,N_4107);
or U4570 (N_4570,N_4427,N_4067);
or U4571 (N_4571,N_4037,N_4318);
xor U4572 (N_4572,N_4490,N_4042);
and U4573 (N_4573,N_4289,N_4161);
and U4574 (N_4574,N_4374,N_4070);
and U4575 (N_4575,N_4143,N_4241);
or U4576 (N_4576,N_4047,N_4423);
and U4577 (N_4577,N_4137,N_4499);
and U4578 (N_4578,N_4057,N_4132);
xnor U4579 (N_4579,N_4254,N_4262);
or U4580 (N_4580,N_4238,N_4309);
nor U4581 (N_4581,N_4082,N_4014);
xor U4582 (N_4582,N_4282,N_4176);
or U4583 (N_4583,N_4433,N_4024);
xor U4584 (N_4584,N_4194,N_4284);
nor U4585 (N_4585,N_4278,N_4235);
and U4586 (N_4586,N_4203,N_4198);
and U4587 (N_4587,N_4372,N_4246);
nand U4588 (N_4588,N_4346,N_4080);
and U4589 (N_4589,N_4458,N_4465);
and U4590 (N_4590,N_4040,N_4466);
or U4591 (N_4591,N_4154,N_4352);
nor U4592 (N_4592,N_4258,N_4461);
nor U4593 (N_4593,N_4139,N_4420);
and U4594 (N_4594,N_4272,N_4085);
nor U4595 (N_4595,N_4464,N_4215);
and U4596 (N_4596,N_4000,N_4265);
and U4597 (N_4597,N_4214,N_4237);
nor U4598 (N_4598,N_4180,N_4090);
xnor U4599 (N_4599,N_4039,N_4079);
xor U4600 (N_4600,N_4297,N_4425);
or U4601 (N_4601,N_4373,N_4392);
or U4602 (N_4602,N_4393,N_4378);
or U4603 (N_4603,N_4335,N_4494);
or U4604 (N_4604,N_4145,N_4315);
xnor U4605 (N_4605,N_4251,N_4492);
nor U4606 (N_4606,N_4463,N_4367);
and U4607 (N_4607,N_4398,N_4115);
and U4608 (N_4608,N_4333,N_4390);
nor U4609 (N_4609,N_4223,N_4472);
or U4610 (N_4610,N_4487,N_4006);
nand U4611 (N_4611,N_4338,N_4207);
or U4612 (N_4612,N_4310,N_4128);
nor U4613 (N_4613,N_4248,N_4409);
or U4614 (N_4614,N_4122,N_4414);
nor U4615 (N_4615,N_4189,N_4025);
xnor U4616 (N_4616,N_4389,N_4328);
nor U4617 (N_4617,N_4077,N_4064);
nor U4618 (N_4618,N_4341,N_4033);
or U4619 (N_4619,N_4271,N_4181);
and U4620 (N_4620,N_4011,N_4256);
or U4621 (N_4621,N_4129,N_4075);
nor U4622 (N_4622,N_4410,N_4192);
nor U4623 (N_4623,N_4220,N_4358);
nor U4624 (N_4624,N_4365,N_4401);
or U4625 (N_4625,N_4422,N_4097);
nand U4626 (N_4626,N_4007,N_4005);
or U4627 (N_4627,N_4030,N_4179);
or U4628 (N_4628,N_4412,N_4388);
nor U4629 (N_4629,N_4404,N_4066);
nand U4630 (N_4630,N_4061,N_4209);
nand U4631 (N_4631,N_4228,N_4158);
nand U4632 (N_4632,N_4439,N_4233);
and U4633 (N_4633,N_4332,N_4098);
nand U4634 (N_4634,N_4291,N_4336);
nand U4635 (N_4635,N_4424,N_4247);
nor U4636 (N_4636,N_4184,N_4408);
or U4637 (N_4637,N_4290,N_4010);
or U4638 (N_4638,N_4305,N_4146);
nor U4639 (N_4639,N_4120,N_4469);
or U4640 (N_4640,N_4350,N_4468);
and U4641 (N_4641,N_4400,N_4103);
or U4642 (N_4642,N_4063,N_4034);
nor U4643 (N_4643,N_4003,N_4084);
or U4644 (N_4644,N_4117,N_4029);
xnor U4645 (N_4645,N_4182,N_4440);
xnor U4646 (N_4646,N_4407,N_4413);
nor U4647 (N_4647,N_4224,N_4156);
and U4648 (N_4648,N_4221,N_4149);
or U4649 (N_4649,N_4160,N_4230);
xnor U4650 (N_4650,N_4086,N_4402);
or U4651 (N_4651,N_4351,N_4312);
xor U4652 (N_4652,N_4421,N_4320);
nand U4653 (N_4653,N_4015,N_4316);
or U4654 (N_4654,N_4190,N_4260);
nand U4655 (N_4655,N_4281,N_4399);
and U4656 (N_4656,N_4359,N_4406);
nor U4657 (N_4657,N_4292,N_4046);
and U4658 (N_4658,N_4380,N_4252);
or U4659 (N_4659,N_4462,N_4394);
nand U4660 (N_4660,N_4074,N_4028);
or U4661 (N_4661,N_4369,N_4321);
and U4662 (N_4662,N_4013,N_4319);
and U4663 (N_4663,N_4355,N_4240);
or U4664 (N_4664,N_4196,N_4459);
nand U4665 (N_4665,N_4293,N_4418);
nand U4666 (N_4666,N_4183,N_4323);
and U4667 (N_4667,N_4211,N_4486);
and U4668 (N_4668,N_4250,N_4411);
and U4669 (N_4669,N_4147,N_4452);
or U4670 (N_4670,N_4088,N_4200);
and U4671 (N_4671,N_4457,N_4142);
or U4672 (N_4672,N_4141,N_4419);
and U4673 (N_4673,N_4185,N_4443);
nor U4674 (N_4674,N_4210,N_4174);
nor U4675 (N_4675,N_4032,N_4280);
xnor U4676 (N_4676,N_4017,N_4330);
or U4677 (N_4677,N_4375,N_4155);
nor U4678 (N_4678,N_4168,N_4178);
nand U4679 (N_4679,N_4314,N_4313);
nor U4680 (N_4680,N_4264,N_4216);
nand U4681 (N_4681,N_4483,N_4479);
nand U4682 (N_4682,N_4099,N_4089);
nand U4683 (N_4683,N_4217,N_4245);
and U4684 (N_4684,N_4052,N_4055);
nor U4685 (N_4685,N_4151,N_4226);
nand U4686 (N_4686,N_4093,N_4109);
nand U4687 (N_4687,N_4322,N_4124);
xnor U4688 (N_4688,N_4307,N_4130);
and U4689 (N_4689,N_4188,N_4261);
and U4690 (N_4690,N_4485,N_4121);
or U4691 (N_4691,N_4437,N_4153);
nand U4692 (N_4692,N_4026,N_4171);
and U4693 (N_4693,N_4277,N_4446);
nand U4694 (N_4694,N_4165,N_4294);
nand U4695 (N_4695,N_4456,N_4354);
nor U4696 (N_4696,N_4162,N_4471);
nand U4697 (N_4697,N_4255,N_4159);
nand U4698 (N_4698,N_4144,N_4253);
nor U4699 (N_4699,N_4383,N_4152);
and U4700 (N_4700,N_4337,N_4387);
or U4701 (N_4701,N_4053,N_4134);
and U4702 (N_4702,N_4363,N_4349);
xnor U4703 (N_4703,N_4391,N_4173);
or U4704 (N_4704,N_4308,N_4083);
nand U4705 (N_4705,N_4167,N_4295);
nor U4706 (N_4706,N_4429,N_4094);
nand U4707 (N_4707,N_4259,N_4488);
nand U4708 (N_4708,N_4114,N_4136);
nand U4709 (N_4709,N_4395,N_4219);
nor U4710 (N_4710,N_4385,N_4020);
nor U4711 (N_4711,N_4062,N_4270);
nand U4712 (N_4712,N_4467,N_4382);
nand U4713 (N_4713,N_4498,N_4324);
and U4714 (N_4714,N_4119,N_4473);
and U4715 (N_4715,N_4353,N_4087);
nand U4716 (N_4716,N_4360,N_4431);
xor U4717 (N_4717,N_4051,N_4201);
nand U4718 (N_4718,N_4111,N_4381);
and U4719 (N_4719,N_4306,N_4371);
xnor U4720 (N_4720,N_4208,N_4428);
and U4721 (N_4721,N_4317,N_4108);
nand U4722 (N_4722,N_4031,N_4202);
and U4723 (N_4723,N_4102,N_4460);
nand U4724 (N_4724,N_4268,N_4489);
nand U4725 (N_4725,N_4257,N_4076);
and U4726 (N_4726,N_4447,N_4417);
xor U4727 (N_4727,N_4301,N_4302);
and U4728 (N_4728,N_4495,N_4213);
and U4729 (N_4729,N_4072,N_4140);
or U4730 (N_4730,N_4331,N_4177);
and U4731 (N_4731,N_4426,N_4009);
and U4732 (N_4732,N_4344,N_4092);
nor U4733 (N_4733,N_4095,N_4118);
xnor U4734 (N_4734,N_4060,N_4186);
or U4735 (N_4735,N_4150,N_4019);
or U4736 (N_4736,N_4123,N_4286);
nor U4737 (N_4737,N_4244,N_4269);
nand U4738 (N_4738,N_4231,N_4275);
nor U4739 (N_4739,N_4048,N_4175);
nor U4740 (N_4740,N_4288,N_4002);
nor U4741 (N_4741,N_4195,N_4081);
xnor U4742 (N_4742,N_4384,N_4204);
or U4743 (N_4743,N_4493,N_4059);
xnor U4744 (N_4744,N_4478,N_4234);
and U4745 (N_4745,N_4187,N_4023);
nor U4746 (N_4746,N_4348,N_4012);
and U4747 (N_4747,N_4491,N_4054);
and U4748 (N_4748,N_4106,N_4164);
nand U4749 (N_4749,N_4370,N_4347);
and U4750 (N_4750,N_4330,N_4386);
nand U4751 (N_4751,N_4194,N_4105);
and U4752 (N_4752,N_4082,N_4366);
xor U4753 (N_4753,N_4095,N_4396);
nand U4754 (N_4754,N_4170,N_4173);
nand U4755 (N_4755,N_4125,N_4271);
xnor U4756 (N_4756,N_4076,N_4485);
or U4757 (N_4757,N_4458,N_4212);
nor U4758 (N_4758,N_4340,N_4117);
nor U4759 (N_4759,N_4140,N_4020);
nor U4760 (N_4760,N_4122,N_4319);
and U4761 (N_4761,N_4180,N_4300);
and U4762 (N_4762,N_4272,N_4087);
and U4763 (N_4763,N_4200,N_4203);
or U4764 (N_4764,N_4482,N_4019);
nand U4765 (N_4765,N_4172,N_4315);
or U4766 (N_4766,N_4022,N_4299);
and U4767 (N_4767,N_4147,N_4210);
nor U4768 (N_4768,N_4399,N_4432);
xnor U4769 (N_4769,N_4325,N_4073);
or U4770 (N_4770,N_4045,N_4128);
or U4771 (N_4771,N_4308,N_4048);
nand U4772 (N_4772,N_4105,N_4217);
or U4773 (N_4773,N_4267,N_4189);
nor U4774 (N_4774,N_4453,N_4084);
and U4775 (N_4775,N_4075,N_4366);
nand U4776 (N_4776,N_4000,N_4013);
xor U4777 (N_4777,N_4385,N_4459);
and U4778 (N_4778,N_4484,N_4040);
xor U4779 (N_4779,N_4429,N_4173);
and U4780 (N_4780,N_4369,N_4404);
or U4781 (N_4781,N_4025,N_4140);
xor U4782 (N_4782,N_4118,N_4345);
nand U4783 (N_4783,N_4385,N_4305);
or U4784 (N_4784,N_4335,N_4109);
nand U4785 (N_4785,N_4350,N_4291);
nand U4786 (N_4786,N_4433,N_4109);
or U4787 (N_4787,N_4268,N_4458);
and U4788 (N_4788,N_4464,N_4456);
nor U4789 (N_4789,N_4069,N_4000);
and U4790 (N_4790,N_4231,N_4165);
nor U4791 (N_4791,N_4093,N_4041);
nor U4792 (N_4792,N_4175,N_4449);
nand U4793 (N_4793,N_4157,N_4124);
or U4794 (N_4794,N_4466,N_4147);
and U4795 (N_4795,N_4443,N_4036);
or U4796 (N_4796,N_4053,N_4059);
or U4797 (N_4797,N_4362,N_4195);
nor U4798 (N_4798,N_4291,N_4081);
xor U4799 (N_4799,N_4048,N_4160);
nor U4800 (N_4800,N_4241,N_4029);
and U4801 (N_4801,N_4427,N_4180);
and U4802 (N_4802,N_4163,N_4029);
or U4803 (N_4803,N_4438,N_4116);
or U4804 (N_4804,N_4219,N_4182);
xnor U4805 (N_4805,N_4331,N_4432);
nand U4806 (N_4806,N_4449,N_4365);
nor U4807 (N_4807,N_4217,N_4303);
nor U4808 (N_4808,N_4122,N_4392);
nand U4809 (N_4809,N_4107,N_4147);
nor U4810 (N_4810,N_4207,N_4461);
nor U4811 (N_4811,N_4127,N_4343);
nor U4812 (N_4812,N_4116,N_4173);
and U4813 (N_4813,N_4126,N_4299);
nand U4814 (N_4814,N_4299,N_4458);
or U4815 (N_4815,N_4282,N_4364);
or U4816 (N_4816,N_4488,N_4172);
nor U4817 (N_4817,N_4464,N_4361);
nor U4818 (N_4818,N_4423,N_4451);
or U4819 (N_4819,N_4240,N_4035);
xnor U4820 (N_4820,N_4160,N_4062);
nor U4821 (N_4821,N_4036,N_4388);
nand U4822 (N_4822,N_4097,N_4016);
and U4823 (N_4823,N_4020,N_4494);
nor U4824 (N_4824,N_4331,N_4191);
nand U4825 (N_4825,N_4310,N_4169);
nor U4826 (N_4826,N_4416,N_4378);
nor U4827 (N_4827,N_4383,N_4452);
or U4828 (N_4828,N_4220,N_4314);
nor U4829 (N_4829,N_4023,N_4270);
and U4830 (N_4830,N_4385,N_4088);
nor U4831 (N_4831,N_4245,N_4014);
or U4832 (N_4832,N_4304,N_4454);
or U4833 (N_4833,N_4321,N_4117);
nand U4834 (N_4834,N_4293,N_4010);
and U4835 (N_4835,N_4465,N_4004);
xnor U4836 (N_4836,N_4073,N_4333);
or U4837 (N_4837,N_4473,N_4136);
xor U4838 (N_4838,N_4244,N_4290);
and U4839 (N_4839,N_4160,N_4312);
nor U4840 (N_4840,N_4240,N_4056);
xor U4841 (N_4841,N_4008,N_4038);
and U4842 (N_4842,N_4482,N_4294);
nand U4843 (N_4843,N_4303,N_4096);
nor U4844 (N_4844,N_4496,N_4314);
nand U4845 (N_4845,N_4332,N_4019);
nor U4846 (N_4846,N_4210,N_4077);
nand U4847 (N_4847,N_4491,N_4335);
nor U4848 (N_4848,N_4294,N_4490);
nand U4849 (N_4849,N_4259,N_4489);
and U4850 (N_4850,N_4206,N_4225);
xnor U4851 (N_4851,N_4045,N_4081);
nand U4852 (N_4852,N_4303,N_4120);
nand U4853 (N_4853,N_4441,N_4018);
nand U4854 (N_4854,N_4473,N_4340);
or U4855 (N_4855,N_4318,N_4422);
or U4856 (N_4856,N_4077,N_4387);
or U4857 (N_4857,N_4006,N_4202);
or U4858 (N_4858,N_4327,N_4313);
nand U4859 (N_4859,N_4088,N_4465);
and U4860 (N_4860,N_4328,N_4348);
or U4861 (N_4861,N_4220,N_4299);
or U4862 (N_4862,N_4010,N_4313);
and U4863 (N_4863,N_4322,N_4155);
and U4864 (N_4864,N_4138,N_4464);
nand U4865 (N_4865,N_4181,N_4133);
or U4866 (N_4866,N_4027,N_4420);
and U4867 (N_4867,N_4186,N_4286);
nor U4868 (N_4868,N_4171,N_4415);
nand U4869 (N_4869,N_4091,N_4314);
nor U4870 (N_4870,N_4299,N_4273);
or U4871 (N_4871,N_4148,N_4147);
or U4872 (N_4872,N_4371,N_4034);
or U4873 (N_4873,N_4310,N_4033);
xnor U4874 (N_4874,N_4499,N_4321);
or U4875 (N_4875,N_4077,N_4148);
or U4876 (N_4876,N_4101,N_4056);
and U4877 (N_4877,N_4155,N_4128);
or U4878 (N_4878,N_4251,N_4203);
nor U4879 (N_4879,N_4257,N_4198);
and U4880 (N_4880,N_4146,N_4094);
or U4881 (N_4881,N_4458,N_4153);
nand U4882 (N_4882,N_4493,N_4255);
nand U4883 (N_4883,N_4477,N_4060);
nor U4884 (N_4884,N_4392,N_4403);
nor U4885 (N_4885,N_4186,N_4250);
or U4886 (N_4886,N_4175,N_4002);
and U4887 (N_4887,N_4374,N_4174);
or U4888 (N_4888,N_4235,N_4338);
xor U4889 (N_4889,N_4052,N_4273);
and U4890 (N_4890,N_4276,N_4302);
nor U4891 (N_4891,N_4205,N_4007);
and U4892 (N_4892,N_4183,N_4115);
nand U4893 (N_4893,N_4391,N_4421);
or U4894 (N_4894,N_4493,N_4495);
nand U4895 (N_4895,N_4108,N_4155);
xnor U4896 (N_4896,N_4245,N_4357);
nor U4897 (N_4897,N_4434,N_4162);
nor U4898 (N_4898,N_4298,N_4442);
or U4899 (N_4899,N_4234,N_4002);
and U4900 (N_4900,N_4345,N_4204);
nand U4901 (N_4901,N_4429,N_4101);
xnor U4902 (N_4902,N_4418,N_4361);
or U4903 (N_4903,N_4300,N_4052);
nand U4904 (N_4904,N_4299,N_4162);
nor U4905 (N_4905,N_4410,N_4179);
xnor U4906 (N_4906,N_4389,N_4255);
nor U4907 (N_4907,N_4456,N_4116);
and U4908 (N_4908,N_4475,N_4262);
nand U4909 (N_4909,N_4195,N_4015);
nor U4910 (N_4910,N_4208,N_4343);
nor U4911 (N_4911,N_4331,N_4473);
and U4912 (N_4912,N_4076,N_4158);
and U4913 (N_4913,N_4431,N_4299);
or U4914 (N_4914,N_4435,N_4196);
nor U4915 (N_4915,N_4478,N_4244);
nand U4916 (N_4916,N_4118,N_4066);
nand U4917 (N_4917,N_4161,N_4017);
nand U4918 (N_4918,N_4370,N_4186);
or U4919 (N_4919,N_4223,N_4270);
or U4920 (N_4920,N_4011,N_4429);
and U4921 (N_4921,N_4485,N_4027);
and U4922 (N_4922,N_4024,N_4441);
nor U4923 (N_4923,N_4026,N_4010);
or U4924 (N_4924,N_4498,N_4088);
and U4925 (N_4925,N_4386,N_4117);
or U4926 (N_4926,N_4222,N_4438);
and U4927 (N_4927,N_4481,N_4492);
and U4928 (N_4928,N_4462,N_4282);
and U4929 (N_4929,N_4293,N_4021);
and U4930 (N_4930,N_4434,N_4422);
nor U4931 (N_4931,N_4335,N_4437);
and U4932 (N_4932,N_4271,N_4089);
and U4933 (N_4933,N_4310,N_4411);
nand U4934 (N_4934,N_4022,N_4488);
nand U4935 (N_4935,N_4247,N_4158);
nor U4936 (N_4936,N_4060,N_4162);
and U4937 (N_4937,N_4008,N_4425);
or U4938 (N_4938,N_4211,N_4489);
nor U4939 (N_4939,N_4023,N_4436);
or U4940 (N_4940,N_4268,N_4492);
or U4941 (N_4941,N_4049,N_4067);
xor U4942 (N_4942,N_4448,N_4144);
nand U4943 (N_4943,N_4397,N_4202);
or U4944 (N_4944,N_4372,N_4105);
nand U4945 (N_4945,N_4292,N_4342);
xor U4946 (N_4946,N_4091,N_4417);
or U4947 (N_4947,N_4060,N_4330);
nor U4948 (N_4948,N_4347,N_4459);
or U4949 (N_4949,N_4197,N_4335);
nand U4950 (N_4950,N_4071,N_4413);
or U4951 (N_4951,N_4419,N_4181);
or U4952 (N_4952,N_4471,N_4451);
and U4953 (N_4953,N_4217,N_4124);
and U4954 (N_4954,N_4450,N_4075);
xor U4955 (N_4955,N_4164,N_4473);
or U4956 (N_4956,N_4258,N_4257);
or U4957 (N_4957,N_4484,N_4367);
and U4958 (N_4958,N_4424,N_4490);
nand U4959 (N_4959,N_4193,N_4209);
nor U4960 (N_4960,N_4401,N_4412);
xnor U4961 (N_4961,N_4101,N_4163);
nand U4962 (N_4962,N_4015,N_4330);
and U4963 (N_4963,N_4427,N_4205);
or U4964 (N_4964,N_4382,N_4259);
and U4965 (N_4965,N_4220,N_4344);
and U4966 (N_4966,N_4180,N_4329);
nor U4967 (N_4967,N_4145,N_4092);
xnor U4968 (N_4968,N_4332,N_4433);
and U4969 (N_4969,N_4282,N_4144);
xor U4970 (N_4970,N_4329,N_4370);
nor U4971 (N_4971,N_4397,N_4463);
or U4972 (N_4972,N_4487,N_4199);
nand U4973 (N_4973,N_4160,N_4331);
and U4974 (N_4974,N_4404,N_4056);
nand U4975 (N_4975,N_4442,N_4234);
nor U4976 (N_4976,N_4472,N_4354);
or U4977 (N_4977,N_4056,N_4298);
nand U4978 (N_4978,N_4340,N_4397);
xor U4979 (N_4979,N_4438,N_4198);
nor U4980 (N_4980,N_4036,N_4137);
or U4981 (N_4981,N_4115,N_4082);
nand U4982 (N_4982,N_4328,N_4400);
nand U4983 (N_4983,N_4193,N_4045);
or U4984 (N_4984,N_4334,N_4108);
and U4985 (N_4985,N_4327,N_4400);
nor U4986 (N_4986,N_4093,N_4430);
nor U4987 (N_4987,N_4472,N_4203);
or U4988 (N_4988,N_4030,N_4107);
or U4989 (N_4989,N_4305,N_4365);
xnor U4990 (N_4990,N_4318,N_4327);
nor U4991 (N_4991,N_4317,N_4445);
nor U4992 (N_4992,N_4231,N_4011);
or U4993 (N_4993,N_4300,N_4288);
nand U4994 (N_4994,N_4274,N_4476);
and U4995 (N_4995,N_4177,N_4483);
or U4996 (N_4996,N_4020,N_4175);
xnor U4997 (N_4997,N_4483,N_4105);
nor U4998 (N_4998,N_4028,N_4213);
nor U4999 (N_4999,N_4325,N_4447);
and U5000 (N_5000,N_4680,N_4918);
or U5001 (N_5001,N_4517,N_4778);
nor U5002 (N_5002,N_4622,N_4961);
or U5003 (N_5003,N_4915,N_4828);
and U5004 (N_5004,N_4742,N_4962);
and U5005 (N_5005,N_4757,N_4790);
nand U5006 (N_5006,N_4955,N_4522);
and U5007 (N_5007,N_4638,N_4510);
nor U5008 (N_5008,N_4660,N_4545);
and U5009 (N_5009,N_4605,N_4741);
and U5010 (N_5010,N_4960,N_4966);
or U5011 (N_5011,N_4783,N_4969);
nand U5012 (N_5012,N_4667,N_4930);
and U5013 (N_5013,N_4939,N_4873);
and U5014 (N_5014,N_4890,N_4670);
xnor U5015 (N_5015,N_4713,N_4781);
and U5016 (N_5016,N_4506,N_4722);
or U5017 (N_5017,N_4989,N_4976);
or U5018 (N_5018,N_4829,N_4628);
and U5019 (N_5019,N_4661,N_4631);
nand U5020 (N_5020,N_4685,N_4926);
or U5021 (N_5021,N_4769,N_4771);
nor U5022 (N_5022,N_4991,N_4659);
nand U5023 (N_5023,N_4501,N_4699);
or U5024 (N_5024,N_4744,N_4750);
nand U5025 (N_5025,N_4526,N_4603);
xor U5026 (N_5026,N_4999,N_4726);
nor U5027 (N_5027,N_4747,N_4513);
and U5028 (N_5028,N_4723,N_4898);
and U5029 (N_5029,N_4871,N_4932);
xor U5030 (N_5030,N_4693,N_4564);
nor U5031 (N_5031,N_4646,N_4888);
or U5032 (N_5032,N_4911,N_4563);
nand U5033 (N_5033,N_4627,N_4602);
nor U5034 (N_5034,N_4633,N_4562);
nor U5035 (N_5035,N_4889,N_4706);
xor U5036 (N_5036,N_4597,N_4585);
xor U5037 (N_5037,N_4756,N_4511);
nor U5038 (N_5038,N_4805,N_4814);
nor U5039 (N_5039,N_4674,N_4573);
xnor U5040 (N_5040,N_4864,N_4752);
nand U5041 (N_5041,N_4621,N_4934);
and U5042 (N_5042,N_4555,N_4874);
nand U5043 (N_5043,N_4524,N_4780);
and U5044 (N_5044,N_4859,N_4914);
or U5045 (N_5045,N_4763,N_4698);
and U5046 (N_5046,N_4664,N_4635);
xnor U5047 (N_5047,N_4988,N_4529);
xor U5048 (N_5048,N_4532,N_4839);
nand U5049 (N_5049,N_4979,N_4982);
or U5050 (N_5050,N_4779,N_4578);
xor U5051 (N_5051,N_4834,N_4904);
xor U5052 (N_5052,N_4694,N_4589);
nand U5053 (N_5053,N_4948,N_4662);
and U5054 (N_5054,N_4987,N_4596);
xnor U5055 (N_5055,N_4590,N_4758);
or U5056 (N_5056,N_4668,N_4574);
nand U5057 (N_5057,N_4802,N_4725);
xor U5058 (N_5058,N_4575,N_4868);
and U5059 (N_5059,N_4774,N_4531);
nor U5060 (N_5060,N_4942,N_4576);
or U5061 (N_5061,N_4831,N_4559);
or U5062 (N_5062,N_4552,N_4708);
and U5063 (N_5063,N_4536,N_4965);
and U5064 (N_5064,N_4862,N_4765);
nand U5065 (N_5065,N_4908,N_4666);
and U5066 (N_5066,N_4619,N_4714);
and U5067 (N_5067,N_4586,N_4587);
nor U5068 (N_5068,N_4858,N_4967);
nor U5069 (N_5069,N_4544,N_4500);
and U5070 (N_5070,N_4632,N_4951);
nor U5071 (N_5071,N_4823,N_4557);
or U5072 (N_5072,N_4877,N_4815);
and U5073 (N_5073,N_4560,N_4715);
nor U5074 (N_5074,N_4849,N_4737);
or U5075 (N_5075,N_4792,N_4755);
nand U5076 (N_5076,N_4860,N_4830);
or U5077 (N_5077,N_4535,N_4920);
or U5078 (N_5078,N_4882,N_4600);
nor U5079 (N_5079,N_4804,N_4593);
or U5080 (N_5080,N_4682,N_4712);
or U5081 (N_5081,N_4970,N_4952);
or U5082 (N_5082,N_4998,N_4703);
or U5083 (N_5083,N_4912,N_4876);
and U5084 (N_5084,N_4630,N_4727);
nand U5085 (N_5085,N_4690,N_4863);
or U5086 (N_5086,N_4766,N_4992);
nor U5087 (N_5087,N_4683,N_4577);
nand U5088 (N_5088,N_4520,N_4537);
and U5089 (N_5089,N_4672,N_4571);
nand U5090 (N_5090,N_4826,N_4624);
nand U5091 (N_5091,N_4907,N_4673);
nand U5092 (N_5092,N_4964,N_4717);
or U5093 (N_5093,N_4940,N_4933);
xor U5094 (N_5094,N_4611,N_4957);
or U5095 (N_5095,N_4827,N_4917);
or U5096 (N_5096,N_4903,N_4588);
xor U5097 (N_5097,N_4840,N_4656);
or U5098 (N_5098,N_4985,N_4865);
or U5099 (N_5099,N_4867,N_4938);
or U5100 (N_5100,N_4734,N_4515);
nor U5101 (N_5101,N_4767,N_4636);
or U5102 (N_5102,N_4838,N_4910);
xor U5103 (N_5103,N_4639,N_4824);
and U5104 (N_5104,N_4533,N_4579);
and U5105 (N_5105,N_4762,N_4978);
nand U5106 (N_5106,N_4740,N_4990);
nand U5107 (N_5107,N_4665,N_4836);
and U5108 (N_5108,N_4896,N_4794);
nor U5109 (N_5109,N_4566,N_4754);
or U5110 (N_5110,N_4642,N_4810);
and U5111 (N_5111,N_4900,N_4539);
nand U5112 (N_5112,N_4542,N_4658);
and U5113 (N_5113,N_4953,N_4791);
or U5114 (N_5114,N_4947,N_4720);
or U5115 (N_5115,N_4972,N_4521);
nor U5116 (N_5116,N_4637,N_4850);
and U5117 (N_5117,N_4817,N_4993);
nand U5118 (N_5118,N_4844,N_4565);
or U5119 (N_5119,N_4608,N_4806);
nand U5120 (N_5120,N_4676,N_4893);
nand U5121 (N_5121,N_4950,N_4880);
or U5122 (N_5122,N_4663,N_4869);
nor U5123 (N_5123,N_4975,N_4853);
and U5124 (N_5124,N_4581,N_4540);
nor U5125 (N_5125,N_4785,N_4886);
or U5126 (N_5126,N_4921,N_4944);
and U5127 (N_5127,N_4803,N_4701);
nor U5128 (N_5128,N_4746,N_4580);
nor U5129 (N_5129,N_4971,N_4695);
and U5130 (N_5130,N_4935,N_4984);
nor U5131 (N_5131,N_4775,N_4753);
xor U5132 (N_5132,N_4881,N_4786);
nor U5133 (N_5133,N_4652,N_4797);
or U5134 (N_5134,N_4813,N_4568);
or U5135 (N_5135,N_4875,N_4538);
or U5136 (N_5136,N_4937,N_4556);
xor U5137 (N_5137,N_4980,N_4997);
nor U5138 (N_5138,N_4894,N_4929);
or U5139 (N_5139,N_4892,N_4609);
or U5140 (N_5140,N_4719,N_4825);
nand U5141 (N_5141,N_4731,N_4958);
nor U5142 (N_5142,N_4856,N_4678);
or U5143 (N_5143,N_4807,N_4547);
nor U5144 (N_5144,N_4629,N_4800);
nor U5145 (N_5145,N_4710,N_4927);
and U5146 (N_5146,N_4743,N_4648);
nor U5147 (N_5147,N_4749,N_4567);
and U5148 (N_5148,N_4595,N_4759);
nand U5149 (N_5149,N_4525,N_4702);
or U5150 (N_5150,N_4822,N_4634);
nor U5151 (N_5151,N_4709,N_4891);
nor U5152 (N_5152,N_4773,N_4931);
nand U5153 (N_5153,N_4919,N_4909);
nor U5154 (N_5154,N_4924,N_4508);
nand U5155 (N_5155,N_4543,N_4684);
nor U5156 (N_5156,N_4598,N_4643);
nor U5157 (N_5157,N_4738,N_4902);
or U5158 (N_5158,N_4857,N_4729);
and U5159 (N_5159,N_4623,N_4973);
or U5160 (N_5160,N_4691,N_4721);
xnor U5161 (N_5161,N_4732,N_4570);
and U5162 (N_5162,N_4735,N_4761);
nor U5163 (N_5163,N_4554,N_4872);
or U5164 (N_5164,N_4616,N_4977);
xor U5165 (N_5165,N_4705,N_4620);
or U5166 (N_5166,N_4878,N_4884);
nand U5167 (N_5167,N_4841,N_4610);
nor U5168 (N_5168,N_4808,N_4916);
nand U5169 (N_5169,N_4711,N_4716);
nand U5170 (N_5170,N_4941,N_4764);
nor U5171 (N_5171,N_4870,N_4730);
nand U5172 (N_5172,N_4528,N_4718);
or U5173 (N_5173,N_4561,N_4640);
xor U5174 (N_5174,N_4550,N_4548);
nor U5175 (N_5175,N_4549,N_4645);
xor U5176 (N_5176,N_4745,N_4594);
and U5177 (N_5177,N_4922,N_4760);
nand U5178 (N_5178,N_4599,N_4959);
nand U5179 (N_5179,N_4897,N_4866);
nand U5180 (N_5180,N_4943,N_4677);
nor U5181 (N_5181,N_4887,N_4818);
and U5182 (N_5182,N_4696,N_4899);
xnor U5183 (N_5183,N_4504,N_4649);
or U5184 (N_5184,N_4795,N_4861);
or U5185 (N_5185,N_4527,N_4883);
nor U5186 (N_5186,N_4626,N_4518);
and U5187 (N_5187,N_4788,N_4514);
and U5188 (N_5188,N_4607,N_4821);
nand U5189 (N_5189,N_4687,N_4816);
and U5190 (N_5190,N_4995,N_4854);
nor U5191 (N_5191,N_4986,N_4669);
and U5192 (N_5192,N_4697,N_4534);
or U5193 (N_5193,N_4801,N_4644);
or U5194 (N_5194,N_4613,N_4601);
or U5195 (N_5195,N_4583,N_4798);
xnor U5196 (N_5196,N_4905,N_4612);
nor U5197 (N_5197,N_4768,N_4519);
or U5198 (N_5198,N_4782,N_4592);
nor U5199 (N_5199,N_4777,N_4641);
or U5200 (N_5200,N_4983,N_4657);
or U5201 (N_5201,N_4647,N_4946);
nor U5202 (N_5202,N_4895,N_4704);
nor U5203 (N_5203,N_4879,N_4981);
and U5204 (N_5204,N_4654,N_4772);
nand U5205 (N_5205,N_4688,N_4546);
nand U5206 (N_5206,N_4655,N_4848);
nor U5207 (N_5207,N_4625,N_4681);
nor U5208 (N_5208,N_4728,N_4776);
or U5209 (N_5209,N_4724,N_4617);
nand U5210 (N_5210,N_4820,N_4949);
nor U5211 (N_5211,N_4692,N_4507);
or U5212 (N_5212,N_4516,N_4503);
and U5213 (N_5213,N_4901,N_4923);
nor U5214 (N_5214,N_4842,N_4653);
nand U5215 (N_5215,N_4906,N_4591);
and U5216 (N_5216,N_4584,N_4835);
nor U5217 (N_5217,N_4799,N_4523);
xor U5218 (N_5218,N_4847,N_4582);
and U5219 (N_5219,N_4679,N_4700);
nor U5220 (N_5220,N_4819,N_4651);
nand U5221 (N_5221,N_4925,N_4811);
nor U5222 (N_5222,N_4968,N_4650);
nand U5223 (N_5223,N_4748,N_4945);
nor U5224 (N_5224,N_4996,N_4604);
nor U5225 (N_5225,N_4541,N_4796);
xor U5226 (N_5226,N_4689,N_4793);
or U5227 (N_5227,N_4509,N_4936);
xor U5228 (N_5228,N_4787,N_4733);
and U5229 (N_5229,N_4675,N_4809);
or U5230 (N_5230,N_4974,N_4671);
nand U5231 (N_5231,N_4707,N_4551);
or U5232 (N_5232,N_4852,N_4770);
or U5233 (N_5233,N_4994,N_4812);
or U5234 (N_5234,N_4928,N_4851);
or U5235 (N_5235,N_4956,N_4569);
or U5236 (N_5236,N_4614,N_4739);
or U5237 (N_5237,N_4963,N_4736);
xor U5238 (N_5238,N_4789,N_4530);
and U5239 (N_5239,N_4837,N_4505);
xor U5240 (N_5240,N_4606,N_4833);
or U5241 (N_5241,N_4751,N_4855);
nor U5242 (N_5242,N_4615,N_4553);
nand U5243 (N_5243,N_4784,N_4572);
nand U5244 (N_5244,N_4846,N_4913);
nand U5245 (N_5245,N_4845,N_4885);
and U5246 (N_5246,N_4832,N_4618);
nor U5247 (N_5247,N_4558,N_4686);
nand U5248 (N_5248,N_4512,N_4954);
or U5249 (N_5249,N_4843,N_4502);
nor U5250 (N_5250,N_4959,N_4933);
nor U5251 (N_5251,N_4520,N_4928);
nand U5252 (N_5252,N_4822,N_4905);
and U5253 (N_5253,N_4594,N_4716);
nor U5254 (N_5254,N_4748,N_4779);
or U5255 (N_5255,N_4686,N_4819);
and U5256 (N_5256,N_4762,N_4988);
nor U5257 (N_5257,N_4544,N_4542);
nand U5258 (N_5258,N_4540,N_4606);
nand U5259 (N_5259,N_4800,N_4949);
nand U5260 (N_5260,N_4613,N_4615);
and U5261 (N_5261,N_4795,N_4960);
and U5262 (N_5262,N_4704,N_4625);
nor U5263 (N_5263,N_4587,N_4794);
and U5264 (N_5264,N_4752,N_4891);
or U5265 (N_5265,N_4509,N_4776);
or U5266 (N_5266,N_4556,N_4636);
or U5267 (N_5267,N_4618,N_4723);
and U5268 (N_5268,N_4710,N_4547);
nor U5269 (N_5269,N_4810,N_4645);
nor U5270 (N_5270,N_4762,N_4586);
nor U5271 (N_5271,N_4802,N_4787);
nor U5272 (N_5272,N_4930,N_4973);
nand U5273 (N_5273,N_4535,N_4940);
nand U5274 (N_5274,N_4910,N_4519);
nor U5275 (N_5275,N_4546,N_4930);
or U5276 (N_5276,N_4698,N_4987);
nor U5277 (N_5277,N_4545,N_4910);
and U5278 (N_5278,N_4569,N_4580);
and U5279 (N_5279,N_4574,N_4858);
nand U5280 (N_5280,N_4583,N_4557);
or U5281 (N_5281,N_4800,N_4925);
nor U5282 (N_5282,N_4842,N_4595);
nor U5283 (N_5283,N_4946,N_4597);
or U5284 (N_5284,N_4780,N_4875);
and U5285 (N_5285,N_4706,N_4712);
xnor U5286 (N_5286,N_4799,N_4548);
nor U5287 (N_5287,N_4823,N_4566);
and U5288 (N_5288,N_4592,N_4954);
nand U5289 (N_5289,N_4616,N_4907);
or U5290 (N_5290,N_4549,N_4919);
nand U5291 (N_5291,N_4839,N_4761);
or U5292 (N_5292,N_4575,N_4677);
nand U5293 (N_5293,N_4524,N_4567);
nor U5294 (N_5294,N_4766,N_4677);
nand U5295 (N_5295,N_4790,N_4509);
nor U5296 (N_5296,N_4858,N_4890);
nor U5297 (N_5297,N_4818,N_4848);
and U5298 (N_5298,N_4716,N_4526);
xnor U5299 (N_5299,N_4515,N_4908);
nand U5300 (N_5300,N_4537,N_4655);
and U5301 (N_5301,N_4652,N_4620);
and U5302 (N_5302,N_4886,N_4568);
nor U5303 (N_5303,N_4606,N_4745);
nand U5304 (N_5304,N_4775,N_4641);
nor U5305 (N_5305,N_4855,N_4551);
or U5306 (N_5306,N_4902,N_4943);
nand U5307 (N_5307,N_4797,N_4915);
or U5308 (N_5308,N_4848,N_4747);
and U5309 (N_5309,N_4983,N_4706);
and U5310 (N_5310,N_4855,N_4836);
and U5311 (N_5311,N_4995,N_4838);
nand U5312 (N_5312,N_4576,N_4878);
and U5313 (N_5313,N_4733,N_4554);
nand U5314 (N_5314,N_4829,N_4569);
nor U5315 (N_5315,N_4725,N_4807);
nand U5316 (N_5316,N_4696,N_4600);
nor U5317 (N_5317,N_4760,N_4586);
and U5318 (N_5318,N_4714,N_4765);
and U5319 (N_5319,N_4990,N_4714);
xor U5320 (N_5320,N_4964,N_4980);
nand U5321 (N_5321,N_4936,N_4944);
nor U5322 (N_5322,N_4903,N_4936);
or U5323 (N_5323,N_4803,N_4597);
or U5324 (N_5324,N_4804,N_4608);
and U5325 (N_5325,N_4951,N_4893);
nor U5326 (N_5326,N_4851,N_4538);
nor U5327 (N_5327,N_4591,N_4750);
or U5328 (N_5328,N_4614,N_4965);
nor U5329 (N_5329,N_4748,N_4535);
and U5330 (N_5330,N_4810,N_4964);
nand U5331 (N_5331,N_4944,N_4615);
and U5332 (N_5332,N_4782,N_4733);
nor U5333 (N_5333,N_4730,N_4667);
or U5334 (N_5334,N_4793,N_4939);
and U5335 (N_5335,N_4771,N_4722);
or U5336 (N_5336,N_4562,N_4952);
xnor U5337 (N_5337,N_4792,N_4647);
and U5338 (N_5338,N_4859,N_4674);
and U5339 (N_5339,N_4783,N_4743);
and U5340 (N_5340,N_4776,N_4827);
nor U5341 (N_5341,N_4520,N_4777);
and U5342 (N_5342,N_4998,N_4881);
and U5343 (N_5343,N_4643,N_4565);
nor U5344 (N_5344,N_4996,N_4946);
nor U5345 (N_5345,N_4538,N_4745);
or U5346 (N_5346,N_4567,N_4799);
xnor U5347 (N_5347,N_4860,N_4511);
xor U5348 (N_5348,N_4930,N_4698);
nand U5349 (N_5349,N_4827,N_4547);
or U5350 (N_5350,N_4583,N_4746);
nand U5351 (N_5351,N_4835,N_4883);
or U5352 (N_5352,N_4978,N_4810);
nor U5353 (N_5353,N_4511,N_4609);
nor U5354 (N_5354,N_4625,N_4725);
nand U5355 (N_5355,N_4661,N_4732);
nor U5356 (N_5356,N_4505,N_4904);
and U5357 (N_5357,N_4638,N_4541);
and U5358 (N_5358,N_4803,N_4854);
nor U5359 (N_5359,N_4831,N_4869);
and U5360 (N_5360,N_4978,N_4796);
or U5361 (N_5361,N_4641,N_4959);
and U5362 (N_5362,N_4601,N_4618);
or U5363 (N_5363,N_4882,N_4678);
and U5364 (N_5364,N_4863,N_4634);
and U5365 (N_5365,N_4934,N_4611);
or U5366 (N_5366,N_4834,N_4823);
nor U5367 (N_5367,N_4733,N_4809);
nand U5368 (N_5368,N_4772,N_4800);
nor U5369 (N_5369,N_4819,N_4976);
or U5370 (N_5370,N_4656,N_4737);
nand U5371 (N_5371,N_4686,N_4954);
nor U5372 (N_5372,N_4774,N_4831);
nand U5373 (N_5373,N_4622,N_4672);
nor U5374 (N_5374,N_4851,N_4937);
nand U5375 (N_5375,N_4534,N_4877);
xnor U5376 (N_5376,N_4931,N_4825);
or U5377 (N_5377,N_4867,N_4970);
or U5378 (N_5378,N_4702,N_4736);
and U5379 (N_5379,N_4971,N_4962);
or U5380 (N_5380,N_4648,N_4974);
or U5381 (N_5381,N_4867,N_4694);
and U5382 (N_5382,N_4673,N_4816);
and U5383 (N_5383,N_4624,N_4766);
nor U5384 (N_5384,N_4560,N_4957);
and U5385 (N_5385,N_4726,N_4831);
or U5386 (N_5386,N_4879,N_4663);
or U5387 (N_5387,N_4736,N_4957);
and U5388 (N_5388,N_4801,N_4824);
nand U5389 (N_5389,N_4514,N_4511);
xor U5390 (N_5390,N_4520,N_4636);
nand U5391 (N_5391,N_4774,N_4867);
and U5392 (N_5392,N_4666,N_4811);
xor U5393 (N_5393,N_4876,N_4530);
nor U5394 (N_5394,N_4975,N_4905);
nor U5395 (N_5395,N_4759,N_4545);
nand U5396 (N_5396,N_4937,N_4551);
or U5397 (N_5397,N_4695,N_4922);
nand U5398 (N_5398,N_4848,N_4555);
and U5399 (N_5399,N_4650,N_4635);
nand U5400 (N_5400,N_4803,N_4692);
xnor U5401 (N_5401,N_4779,N_4633);
nand U5402 (N_5402,N_4754,N_4930);
xnor U5403 (N_5403,N_4549,N_4665);
and U5404 (N_5404,N_4581,N_4664);
or U5405 (N_5405,N_4984,N_4617);
or U5406 (N_5406,N_4969,N_4904);
and U5407 (N_5407,N_4894,N_4852);
nor U5408 (N_5408,N_4983,N_4674);
nor U5409 (N_5409,N_4917,N_4895);
nand U5410 (N_5410,N_4640,N_4828);
nand U5411 (N_5411,N_4956,N_4763);
nand U5412 (N_5412,N_4968,N_4823);
and U5413 (N_5413,N_4929,N_4761);
nand U5414 (N_5414,N_4903,N_4830);
and U5415 (N_5415,N_4540,N_4580);
xnor U5416 (N_5416,N_4645,N_4529);
or U5417 (N_5417,N_4512,N_4897);
or U5418 (N_5418,N_4891,N_4576);
nand U5419 (N_5419,N_4519,N_4515);
or U5420 (N_5420,N_4977,N_4755);
nor U5421 (N_5421,N_4841,N_4871);
nand U5422 (N_5422,N_4788,N_4608);
nand U5423 (N_5423,N_4674,N_4546);
or U5424 (N_5424,N_4835,N_4708);
and U5425 (N_5425,N_4835,N_4864);
nor U5426 (N_5426,N_4750,N_4565);
xor U5427 (N_5427,N_4968,N_4994);
nor U5428 (N_5428,N_4764,N_4675);
nor U5429 (N_5429,N_4748,N_4742);
and U5430 (N_5430,N_4656,N_4524);
or U5431 (N_5431,N_4948,N_4955);
nand U5432 (N_5432,N_4805,N_4748);
or U5433 (N_5433,N_4784,N_4864);
nand U5434 (N_5434,N_4678,N_4628);
nand U5435 (N_5435,N_4640,N_4833);
or U5436 (N_5436,N_4967,N_4954);
or U5437 (N_5437,N_4837,N_4695);
xnor U5438 (N_5438,N_4659,N_4844);
xnor U5439 (N_5439,N_4709,N_4517);
or U5440 (N_5440,N_4675,N_4667);
nand U5441 (N_5441,N_4781,N_4587);
and U5442 (N_5442,N_4979,N_4995);
nand U5443 (N_5443,N_4842,N_4897);
nand U5444 (N_5444,N_4533,N_4624);
nand U5445 (N_5445,N_4544,N_4625);
nor U5446 (N_5446,N_4630,N_4853);
and U5447 (N_5447,N_4665,N_4652);
xor U5448 (N_5448,N_4515,N_4593);
nor U5449 (N_5449,N_4804,N_4644);
and U5450 (N_5450,N_4813,N_4782);
nor U5451 (N_5451,N_4677,N_4805);
nor U5452 (N_5452,N_4893,N_4541);
and U5453 (N_5453,N_4870,N_4610);
or U5454 (N_5454,N_4980,N_4634);
nand U5455 (N_5455,N_4878,N_4868);
and U5456 (N_5456,N_4677,N_4908);
xor U5457 (N_5457,N_4943,N_4774);
nor U5458 (N_5458,N_4854,N_4653);
or U5459 (N_5459,N_4925,N_4859);
and U5460 (N_5460,N_4864,N_4677);
and U5461 (N_5461,N_4843,N_4774);
nor U5462 (N_5462,N_4632,N_4547);
nand U5463 (N_5463,N_4540,N_4564);
or U5464 (N_5464,N_4976,N_4668);
xnor U5465 (N_5465,N_4816,N_4639);
and U5466 (N_5466,N_4868,N_4518);
nand U5467 (N_5467,N_4839,N_4553);
xnor U5468 (N_5468,N_4544,N_4618);
nor U5469 (N_5469,N_4580,N_4586);
and U5470 (N_5470,N_4682,N_4590);
or U5471 (N_5471,N_4876,N_4880);
and U5472 (N_5472,N_4535,N_4589);
nor U5473 (N_5473,N_4995,N_4878);
xnor U5474 (N_5474,N_4995,N_4829);
and U5475 (N_5475,N_4723,N_4749);
nor U5476 (N_5476,N_4963,N_4716);
nand U5477 (N_5477,N_4866,N_4596);
nor U5478 (N_5478,N_4900,N_4876);
nor U5479 (N_5479,N_4823,N_4517);
or U5480 (N_5480,N_4511,N_4863);
xnor U5481 (N_5481,N_4758,N_4576);
xnor U5482 (N_5482,N_4882,N_4704);
nor U5483 (N_5483,N_4530,N_4825);
nor U5484 (N_5484,N_4852,N_4872);
and U5485 (N_5485,N_4800,N_4513);
or U5486 (N_5486,N_4740,N_4591);
xnor U5487 (N_5487,N_4804,N_4701);
and U5488 (N_5488,N_4701,N_4645);
xnor U5489 (N_5489,N_4555,N_4880);
and U5490 (N_5490,N_4943,N_4524);
nand U5491 (N_5491,N_4724,N_4983);
and U5492 (N_5492,N_4743,N_4737);
nand U5493 (N_5493,N_4772,N_4535);
and U5494 (N_5494,N_4749,N_4857);
xnor U5495 (N_5495,N_4756,N_4683);
nor U5496 (N_5496,N_4572,N_4610);
nand U5497 (N_5497,N_4772,N_4880);
and U5498 (N_5498,N_4713,N_4631);
and U5499 (N_5499,N_4613,N_4763);
or U5500 (N_5500,N_5294,N_5188);
nor U5501 (N_5501,N_5228,N_5110);
nor U5502 (N_5502,N_5205,N_5279);
or U5503 (N_5503,N_5030,N_5135);
nand U5504 (N_5504,N_5160,N_5190);
nor U5505 (N_5505,N_5398,N_5231);
xnor U5506 (N_5506,N_5291,N_5462);
nor U5507 (N_5507,N_5070,N_5498);
nand U5508 (N_5508,N_5393,N_5060);
xnor U5509 (N_5509,N_5109,N_5375);
and U5510 (N_5510,N_5112,N_5009);
or U5511 (N_5511,N_5316,N_5148);
xor U5512 (N_5512,N_5366,N_5194);
and U5513 (N_5513,N_5330,N_5132);
nand U5514 (N_5514,N_5390,N_5441);
and U5515 (N_5515,N_5453,N_5467);
or U5516 (N_5516,N_5254,N_5180);
and U5517 (N_5517,N_5040,N_5173);
nand U5518 (N_5518,N_5384,N_5359);
and U5519 (N_5519,N_5172,N_5195);
or U5520 (N_5520,N_5347,N_5058);
nand U5521 (N_5521,N_5078,N_5167);
or U5522 (N_5522,N_5007,N_5349);
xnor U5523 (N_5523,N_5481,N_5090);
nand U5524 (N_5524,N_5120,N_5168);
nor U5525 (N_5525,N_5171,N_5389);
and U5526 (N_5526,N_5494,N_5333);
and U5527 (N_5527,N_5037,N_5255);
or U5528 (N_5528,N_5154,N_5065);
nand U5529 (N_5529,N_5401,N_5286);
nand U5530 (N_5530,N_5408,N_5406);
nand U5531 (N_5531,N_5162,N_5410);
nor U5532 (N_5532,N_5118,N_5287);
nand U5533 (N_5533,N_5310,N_5015);
nand U5534 (N_5534,N_5385,N_5034);
and U5535 (N_5535,N_5274,N_5036);
nand U5536 (N_5536,N_5415,N_5491);
and U5537 (N_5537,N_5456,N_5331);
nand U5538 (N_5538,N_5003,N_5478);
and U5539 (N_5539,N_5332,N_5016);
nor U5540 (N_5540,N_5069,N_5426);
nand U5541 (N_5541,N_5062,N_5271);
or U5542 (N_5542,N_5409,N_5305);
or U5543 (N_5543,N_5068,N_5425);
nor U5544 (N_5544,N_5073,N_5327);
and U5545 (N_5545,N_5430,N_5324);
xor U5546 (N_5546,N_5296,N_5391);
and U5547 (N_5547,N_5397,N_5284);
or U5548 (N_5548,N_5292,N_5353);
and U5549 (N_5549,N_5202,N_5434);
nand U5550 (N_5550,N_5107,N_5270);
and U5551 (N_5551,N_5224,N_5127);
nand U5552 (N_5552,N_5479,N_5043);
nor U5553 (N_5553,N_5265,N_5155);
and U5554 (N_5554,N_5304,N_5309);
or U5555 (N_5555,N_5227,N_5241);
nor U5556 (N_5556,N_5178,N_5496);
or U5557 (N_5557,N_5087,N_5288);
and U5558 (N_5558,N_5215,N_5192);
nand U5559 (N_5559,N_5350,N_5329);
nand U5560 (N_5560,N_5437,N_5031);
or U5561 (N_5561,N_5485,N_5454);
and U5562 (N_5562,N_5337,N_5232);
nand U5563 (N_5563,N_5199,N_5374);
or U5564 (N_5564,N_5251,N_5080);
and U5565 (N_5565,N_5487,N_5318);
or U5566 (N_5566,N_5448,N_5138);
and U5567 (N_5567,N_5463,N_5365);
nand U5568 (N_5568,N_5189,N_5362);
and U5569 (N_5569,N_5412,N_5308);
or U5570 (N_5570,N_5339,N_5466);
or U5571 (N_5571,N_5064,N_5085);
nor U5572 (N_5572,N_5414,N_5367);
nand U5573 (N_5573,N_5262,N_5044);
nand U5574 (N_5574,N_5038,N_5157);
or U5575 (N_5575,N_5095,N_5026);
nor U5576 (N_5576,N_5144,N_5495);
nor U5577 (N_5577,N_5045,N_5360);
or U5578 (N_5578,N_5092,N_5295);
or U5579 (N_5579,N_5442,N_5435);
nor U5580 (N_5580,N_5021,N_5388);
nor U5581 (N_5581,N_5394,N_5220);
nor U5582 (N_5582,N_5383,N_5222);
or U5583 (N_5583,N_5404,N_5125);
nand U5584 (N_5584,N_5378,N_5020);
nand U5585 (N_5585,N_5124,N_5055);
xnor U5586 (N_5586,N_5186,N_5142);
or U5587 (N_5587,N_5381,N_5019);
and U5588 (N_5588,N_5100,N_5297);
nor U5589 (N_5589,N_5281,N_5244);
nand U5590 (N_5590,N_5084,N_5344);
or U5591 (N_5591,N_5252,N_5351);
nor U5592 (N_5592,N_5032,N_5126);
or U5593 (N_5593,N_5290,N_5341);
nand U5594 (N_5594,N_5129,N_5438);
or U5595 (N_5595,N_5276,N_5358);
xnor U5596 (N_5596,N_5348,N_5153);
and U5597 (N_5597,N_5312,N_5427);
nor U5598 (N_5598,N_5470,N_5493);
or U5599 (N_5599,N_5422,N_5443);
xnor U5600 (N_5600,N_5203,N_5147);
nand U5601 (N_5601,N_5176,N_5379);
nand U5602 (N_5602,N_5008,N_5041);
or U5603 (N_5603,N_5460,N_5216);
nor U5604 (N_5604,N_5074,N_5079);
or U5605 (N_5605,N_5277,N_5407);
nor U5606 (N_5606,N_5417,N_5091);
nor U5607 (N_5607,N_5424,N_5400);
and U5608 (N_5608,N_5285,N_5429);
xnor U5609 (N_5609,N_5187,N_5421);
nand U5610 (N_5610,N_5206,N_5177);
and U5611 (N_5611,N_5063,N_5071);
nand U5612 (N_5612,N_5455,N_5081);
and U5613 (N_5613,N_5150,N_5159);
nand U5614 (N_5614,N_5257,N_5418);
and U5615 (N_5615,N_5102,N_5137);
or U5616 (N_5616,N_5122,N_5136);
or U5617 (N_5617,N_5240,N_5233);
xnor U5618 (N_5618,N_5245,N_5230);
or U5619 (N_5619,N_5130,N_5354);
or U5620 (N_5620,N_5372,N_5301);
nor U5621 (N_5621,N_5208,N_5121);
or U5622 (N_5622,N_5183,N_5447);
or U5623 (N_5623,N_5403,N_5311);
nand U5624 (N_5624,N_5017,N_5077);
or U5625 (N_5625,N_5143,N_5345);
and U5626 (N_5626,N_5432,N_5209);
xnor U5627 (N_5627,N_5317,N_5005);
or U5628 (N_5628,N_5185,N_5486);
xor U5629 (N_5629,N_5174,N_5335);
and U5630 (N_5630,N_5357,N_5000);
nand U5631 (N_5631,N_5169,N_5196);
nor U5632 (N_5632,N_5247,N_5175);
nor U5633 (N_5633,N_5035,N_5246);
nand U5634 (N_5634,N_5259,N_5483);
nor U5635 (N_5635,N_5033,N_5269);
or U5636 (N_5636,N_5303,N_5342);
and U5637 (N_5637,N_5067,N_5096);
or U5638 (N_5638,N_5219,N_5115);
xor U5639 (N_5639,N_5086,N_5113);
nand U5640 (N_5640,N_5472,N_5218);
nor U5641 (N_5641,N_5264,N_5278);
nand U5642 (N_5642,N_5371,N_5315);
nor U5643 (N_5643,N_5382,N_5306);
and U5644 (N_5644,N_5061,N_5198);
nand U5645 (N_5645,N_5399,N_5461);
nand U5646 (N_5646,N_5156,N_5238);
nor U5647 (N_5647,N_5013,N_5165);
nand U5648 (N_5648,N_5321,N_5346);
nor U5649 (N_5649,N_5475,N_5322);
or U5650 (N_5650,N_5313,N_5014);
or U5651 (N_5651,N_5088,N_5166);
and U5652 (N_5652,N_5179,N_5093);
and U5653 (N_5653,N_5201,N_5082);
or U5654 (N_5654,N_5370,N_5225);
nor U5655 (N_5655,N_5488,N_5193);
nor U5656 (N_5656,N_5207,N_5001);
and U5657 (N_5657,N_5145,N_5465);
nand U5658 (N_5658,N_5151,N_5268);
and U5659 (N_5659,N_5048,N_5140);
nand U5660 (N_5660,N_5146,N_5103);
or U5661 (N_5661,N_5056,N_5094);
nand U5662 (N_5662,N_5029,N_5413);
and U5663 (N_5663,N_5267,N_5027);
and U5664 (N_5664,N_5307,N_5200);
nand U5665 (N_5665,N_5119,N_5053);
nand U5666 (N_5666,N_5158,N_5051);
xnor U5667 (N_5667,N_5428,N_5010);
and U5668 (N_5668,N_5490,N_5273);
nor U5669 (N_5669,N_5433,N_5239);
or U5670 (N_5670,N_5226,N_5364);
nor U5671 (N_5671,N_5477,N_5237);
and U5672 (N_5672,N_5340,N_5046);
nor U5673 (N_5673,N_5387,N_5235);
nor U5674 (N_5674,N_5012,N_5212);
nor U5675 (N_5675,N_5280,N_5163);
and U5676 (N_5676,N_5057,N_5320);
xnor U5677 (N_5677,N_5473,N_5242);
and U5678 (N_5678,N_5452,N_5319);
nand U5679 (N_5679,N_5039,N_5289);
nand U5680 (N_5680,N_5386,N_5023);
or U5681 (N_5681,N_5223,N_5117);
nor U5682 (N_5682,N_5217,N_5499);
nand U5683 (N_5683,N_5028,N_5256);
xor U5684 (N_5684,N_5170,N_5469);
nor U5685 (N_5685,N_5105,N_5396);
nand U5686 (N_5686,N_5373,N_5152);
and U5687 (N_5687,N_5369,N_5336);
nor U5688 (N_5688,N_5101,N_5423);
nand U5689 (N_5689,N_5464,N_5139);
nor U5690 (N_5690,N_5492,N_5002);
nand U5691 (N_5691,N_5263,N_5444);
nor U5692 (N_5692,N_5323,N_5293);
or U5693 (N_5693,N_5299,N_5368);
nand U5694 (N_5694,N_5474,N_5141);
xor U5695 (N_5695,N_5076,N_5440);
nor U5696 (N_5696,N_5468,N_5376);
xor U5697 (N_5697,N_5116,N_5405);
nand U5698 (N_5698,N_5451,N_5022);
and U5699 (N_5699,N_5004,N_5355);
or U5700 (N_5700,N_5213,N_5131);
and U5701 (N_5701,N_5184,N_5449);
xnor U5702 (N_5702,N_5352,N_5210);
and U5703 (N_5703,N_5392,N_5204);
nor U5704 (N_5704,N_5300,N_5108);
and U5705 (N_5705,N_5497,N_5250);
or U5706 (N_5706,N_5052,N_5458);
xnor U5707 (N_5707,N_5083,N_5164);
or U5708 (N_5708,N_5211,N_5361);
and U5709 (N_5709,N_5134,N_5197);
or U5710 (N_5710,N_5334,N_5042);
nand U5711 (N_5711,N_5283,N_5325);
or U5712 (N_5712,N_5221,N_5482);
xor U5713 (N_5713,N_5050,N_5298);
or U5714 (N_5714,N_5018,N_5395);
nor U5715 (N_5715,N_5272,N_5236);
xnor U5716 (N_5716,N_5099,N_5450);
xnor U5717 (N_5717,N_5161,N_5114);
nor U5718 (N_5718,N_5420,N_5006);
and U5719 (N_5719,N_5266,N_5459);
and U5720 (N_5720,N_5181,N_5243);
or U5721 (N_5721,N_5123,N_5229);
and U5722 (N_5722,N_5098,N_5234);
nor U5723 (N_5723,N_5054,N_5457);
nand U5724 (N_5724,N_5302,N_5328);
nand U5725 (N_5725,N_5377,N_5326);
xnor U5726 (N_5726,N_5275,N_5416);
xor U5727 (N_5727,N_5439,N_5431);
or U5728 (N_5728,N_5260,N_5066);
nand U5729 (N_5729,N_5261,N_5191);
nor U5730 (N_5730,N_5446,N_5097);
nand U5731 (N_5731,N_5104,N_5106);
and U5732 (N_5732,N_5248,N_5476);
nor U5733 (N_5733,N_5363,N_5149);
nand U5734 (N_5734,N_5356,N_5489);
or U5735 (N_5735,N_5258,N_5182);
or U5736 (N_5736,N_5419,N_5445);
nand U5737 (N_5737,N_5480,N_5047);
or U5738 (N_5738,N_5075,N_5471);
xor U5739 (N_5739,N_5049,N_5214);
xnor U5740 (N_5740,N_5025,N_5072);
nand U5741 (N_5741,N_5282,N_5133);
nor U5742 (N_5742,N_5402,N_5059);
or U5743 (N_5743,N_5024,N_5253);
and U5744 (N_5744,N_5011,N_5111);
nor U5745 (N_5745,N_5314,N_5128);
and U5746 (N_5746,N_5343,N_5089);
nand U5747 (N_5747,N_5411,N_5380);
or U5748 (N_5748,N_5338,N_5436);
and U5749 (N_5749,N_5249,N_5484);
nor U5750 (N_5750,N_5469,N_5491);
or U5751 (N_5751,N_5412,N_5102);
and U5752 (N_5752,N_5216,N_5160);
or U5753 (N_5753,N_5013,N_5494);
nor U5754 (N_5754,N_5470,N_5027);
nor U5755 (N_5755,N_5265,N_5254);
xor U5756 (N_5756,N_5290,N_5005);
xnor U5757 (N_5757,N_5359,N_5403);
nand U5758 (N_5758,N_5438,N_5377);
xnor U5759 (N_5759,N_5287,N_5340);
or U5760 (N_5760,N_5057,N_5084);
or U5761 (N_5761,N_5170,N_5322);
nand U5762 (N_5762,N_5384,N_5370);
xnor U5763 (N_5763,N_5461,N_5380);
or U5764 (N_5764,N_5372,N_5113);
nor U5765 (N_5765,N_5299,N_5278);
nand U5766 (N_5766,N_5107,N_5374);
and U5767 (N_5767,N_5062,N_5457);
and U5768 (N_5768,N_5338,N_5485);
and U5769 (N_5769,N_5240,N_5004);
nor U5770 (N_5770,N_5184,N_5388);
nand U5771 (N_5771,N_5140,N_5200);
and U5772 (N_5772,N_5377,N_5003);
and U5773 (N_5773,N_5479,N_5340);
nand U5774 (N_5774,N_5165,N_5133);
xnor U5775 (N_5775,N_5424,N_5394);
nor U5776 (N_5776,N_5245,N_5432);
and U5777 (N_5777,N_5499,N_5311);
nor U5778 (N_5778,N_5185,N_5349);
nor U5779 (N_5779,N_5370,N_5345);
nor U5780 (N_5780,N_5080,N_5254);
nand U5781 (N_5781,N_5408,N_5052);
nand U5782 (N_5782,N_5403,N_5065);
xor U5783 (N_5783,N_5450,N_5000);
nor U5784 (N_5784,N_5278,N_5391);
and U5785 (N_5785,N_5007,N_5131);
nand U5786 (N_5786,N_5143,N_5228);
or U5787 (N_5787,N_5119,N_5098);
or U5788 (N_5788,N_5049,N_5430);
xor U5789 (N_5789,N_5387,N_5324);
nor U5790 (N_5790,N_5298,N_5466);
and U5791 (N_5791,N_5239,N_5242);
or U5792 (N_5792,N_5235,N_5072);
nand U5793 (N_5793,N_5090,N_5173);
or U5794 (N_5794,N_5083,N_5469);
and U5795 (N_5795,N_5435,N_5071);
and U5796 (N_5796,N_5010,N_5142);
nor U5797 (N_5797,N_5175,N_5318);
or U5798 (N_5798,N_5481,N_5086);
or U5799 (N_5799,N_5450,N_5091);
nor U5800 (N_5800,N_5283,N_5437);
and U5801 (N_5801,N_5486,N_5391);
nor U5802 (N_5802,N_5303,N_5458);
and U5803 (N_5803,N_5457,N_5367);
nand U5804 (N_5804,N_5466,N_5263);
or U5805 (N_5805,N_5039,N_5312);
xnor U5806 (N_5806,N_5438,N_5136);
nand U5807 (N_5807,N_5294,N_5471);
and U5808 (N_5808,N_5204,N_5166);
nand U5809 (N_5809,N_5320,N_5153);
and U5810 (N_5810,N_5344,N_5413);
and U5811 (N_5811,N_5466,N_5398);
and U5812 (N_5812,N_5398,N_5080);
or U5813 (N_5813,N_5393,N_5139);
nor U5814 (N_5814,N_5203,N_5217);
xnor U5815 (N_5815,N_5170,N_5244);
and U5816 (N_5816,N_5451,N_5334);
nand U5817 (N_5817,N_5410,N_5138);
nand U5818 (N_5818,N_5209,N_5126);
and U5819 (N_5819,N_5469,N_5196);
nor U5820 (N_5820,N_5017,N_5021);
nand U5821 (N_5821,N_5291,N_5385);
and U5822 (N_5822,N_5408,N_5026);
nor U5823 (N_5823,N_5279,N_5339);
nand U5824 (N_5824,N_5147,N_5278);
nor U5825 (N_5825,N_5180,N_5419);
or U5826 (N_5826,N_5467,N_5148);
nand U5827 (N_5827,N_5289,N_5317);
nand U5828 (N_5828,N_5111,N_5389);
nor U5829 (N_5829,N_5086,N_5065);
xnor U5830 (N_5830,N_5497,N_5268);
nand U5831 (N_5831,N_5048,N_5255);
nand U5832 (N_5832,N_5142,N_5220);
xnor U5833 (N_5833,N_5158,N_5148);
or U5834 (N_5834,N_5298,N_5446);
and U5835 (N_5835,N_5407,N_5207);
nand U5836 (N_5836,N_5259,N_5040);
nor U5837 (N_5837,N_5425,N_5375);
nor U5838 (N_5838,N_5294,N_5321);
or U5839 (N_5839,N_5425,N_5484);
or U5840 (N_5840,N_5060,N_5048);
nand U5841 (N_5841,N_5208,N_5357);
nor U5842 (N_5842,N_5192,N_5086);
nor U5843 (N_5843,N_5105,N_5008);
xor U5844 (N_5844,N_5088,N_5049);
or U5845 (N_5845,N_5458,N_5207);
nand U5846 (N_5846,N_5301,N_5414);
or U5847 (N_5847,N_5245,N_5478);
nand U5848 (N_5848,N_5088,N_5035);
nand U5849 (N_5849,N_5458,N_5205);
or U5850 (N_5850,N_5453,N_5491);
nor U5851 (N_5851,N_5163,N_5485);
and U5852 (N_5852,N_5259,N_5482);
xor U5853 (N_5853,N_5399,N_5438);
or U5854 (N_5854,N_5299,N_5114);
or U5855 (N_5855,N_5485,N_5150);
and U5856 (N_5856,N_5352,N_5491);
nand U5857 (N_5857,N_5289,N_5227);
nor U5858 (N_5858,N_5211,N_5256);
or U5859 (N_5859,N_5388,N_5451);
nand U5860 (N_5860,N_5367,N_5386);
nor U5861 (N_5861,N_5144,N_5370);
xnor U5862 (N_5862,N_5367,N_5116);
and U5863 (N_5863,N_5251,N_5141);
nor U5864 (N_5864,N_5263,N_5216);
or U5865 (N_5865,N_5264,N_5473);
and U5866 (N_5866,N_5416,N_5307);
nand U5867 (N_5867,N_5421,N_5418);
or U5868 (N_5868,N_5481,N_5107);
or U5869 (N_5869,N_5010,N_5106);
nor U5870 (N_5870,N_5470,N_5309);
and U5871 (N_5871,N_5074,N_5102);
nand U5872 (N_5872,N_5094,N_5483);
nor U5873 (N_5873,N_5165,N_5487);
xnor U5874 (N_5874,N_5189,N_5091);
or U5875 (N_5875,N_5102,N_5157);
and U5876 (N_5876,N_5041,N_5185);
nand U5877 (N_5877,N_5399,N_5394);
nand U5878 (N_5878,N_5017,N_5327);
or U5879 (N_5879,N_5466,N_5109);
nor U5880 (N_5880,N_5458,N_5457);
nor U5881 (N_5881,N_5213,N_5490);
or U5882 (N_5882,N_5009,N_5301);
nor U5883 (N_5883,N_5496,N_5324);
or U5884 (N_5884,N_5011,N_5224);
nor U5885 (N_5885,N_5068,N_5469);
xor U5886 (N_5886,N_5037,N_5212);
or U5887 (N_5887,N_5300,N_5466);
xor U5888 (N_5888,N_5407,N_5050);
nand U5889 (N_5889,N_5336,N_5381);
nor U5890 (N_5890,N_5177,N_5060);
nand U5891 (N_5891,N_5398,N_5168);
and U5892 (N_5892,N_5326,N_5460);
and U5893 (N_5893,N_5063,N_5407);
and U5894 (N_5894,N_5173,N_5137);
or U5895 (N_5895,N_5112,N_5460);
nand U5896 (N_5896,N_5222,N_5036);
nor U5897 (N_5897,N_5491,N_5356);
or U5898 (N_5898,N_5071,N_5430);
nand U5899 (N_5899,N_5178,N_5357);
and U5900 (N_5900,N_5402,N_5015);
or U5901 (N_5901,N_5475,N_5065);
nor U5902 (N_5902,N_5050,N_5281);
xnor U5903 (N_5903,N_5404,N_5093);
nand U5904 (N_5904,N_5239,N_5345);
and U5905 (N_5905,N_5111,N_5308);
nor U5906 (N_5906,N_5466,N_5304);
xor U5907 (N_5907,N_5162,N_5486);
nor U5908 (N_5908,N_5239,N_5498);
or U5909 (N_5909,N_5251,N_5451);
or U5910 (N_5910,N_5380,N_5276);
or U5911 (N_5911,N_5043,N_5220);
nand U5912 (N_5912,N_5496,N_5417);
xor U5913 (N_5913,N_5361,N_5394);
and U5914 (N_5914,N_5458,N_5137);
nand U5915 (N_5915,N_5084,N_5374);
xor U5916 (N_5916,N_5497,N_5159);
nand U5917 (N_5917,N_5431,N_5373);
and U5918 (N_5918,N_5391,N_5242);
xnor U5919 (N_5919,N_5487,N_5418);
nand U5920 (N_5920,N_5241,N_5390);
nand U5921 (N_5921,N_5086,N_5132);
and U5922 (N_5922,N_5125,N_5329);
nor U5923 (N_5923,N_5347,N_5141);
nor U5924 (N_5924,N_5145,N_5071);
nor U5925 (N_5925,N_5403,N_5110);
and U5926 (N_5926,N_5447,N_5060);
xnor U5927 (N_5927,N_5334,N_5344);
nor U5928 (N_5928,N_5326,N_5451);
or U5929 (N_5929,N_5169,N_5025);
or U5930 (N_5930,N_5108,N_5462);
and U5931 (N_5931,N_5027,N_5074);
or U5932 (N_5932,N_5128,N_5182);
nand U5933 (N_5933,N_5155,N_5404);
xor U5934 (N_5934,N_5075,N_5254);
or U5935 (N_5935,N_5148,N_5135);
nor U5936 (N_5936,N_5329,N_5223);
and U5937 (N_5937,N_5172,N_5058);
nor U5938 (N_5938,N_5279,N_5012);
or U5939 (N_5939,N_5223,N_5064);
and U5940 (N_5940,N_5357,N_5308);
nand U5941 (N_5941,N_5078,N_5137);
nand U5942 (N_5942,N_5038,N_5342);
or U5943 (N_5943,N_5385,N_5197);
or U5944 (N_5944,N_5400,N_5196);
xor U5945 (N_5945,N_5469,N_5487);
nor U5946 (N_5946,N_5252,N_5310);
or U5947 (N_5947,N_5057,N_5383);
or U5948 (N_5948,N_5260,N_5317);
or U5949 (N_5949,N_5197,N_5046);
or U5950 (N_5950,N_5256,N_5218);
or U5951 (N_5951,N_5481,N_5306);
nor U5952 (N_5952,N_5443,N_5434);
nand U5953 (N_5953,N_5250,N_5304);
and U5954 (N_5954,N_5440,N_5311);
nor U5955 (N_5955,N_5292,N_5248);
or U5956 (N_5956,N_5027,N_5356);
or U5957 (N_5957,N_5200,N_5384);
or U5958 (N_5958,N_5498,N_5275);
and U5959 (N_5959,N_5170,N_5203);
nor U5960 (N_5960,N_5135,N_5401);
nor U5961 (N_5961,N_5151,N_5292);
nor U5962 (N_5962,N_5239,N_5400);
and U5963 (N_5963,N_5099,N_5277);
or U5964 (N_5964,N_5317,N_5316);
nor U5965 (N_5965,N_5145,N_5376);
nand U5966 (N_5966,N_5387,N_5315);
or U5967 (N_5967,N_5295,N_5149);
xnor U5968 (N_5968,N_5317,N_5032);
xnor U5969 (N_5969,N_5074,N_5119);
or U5970 (N_5970,N_5103,N_5399);
nand U5971 (N_5971,N_5050,N_5415);
or U5972 (N_5972,N_5240,N_5153);
nor U5973 (N_5973,N_5433,N_5219);
or U5974 (N_5974,N_5275,N_5055);
nor U5975 (N_5975,N_5186,N_5219);
or U5976 (N_5976,N_5252,N_5302);
xnor U5977 (N_5977,N_5134,N_5385);
nor U5978 (N_5978,N_5448,N_5002);
nor U5979 (N_5979,N_5351,N_5331);
or U5980 (N_5980,N_5117,N_5206);
and U5981 (N_5981,N_5065,N_5456);
and U5982 (N_5982,N_5237,N_5198);
and U5983 (N_5983,N_5127,N_5440);
and U5984 (N_5984,N_5289,N_5003);
nor U5985 (N_5985,N_5009,N_5024);
nand U5986 (N_5986,N_5390,N_5024);
nand U5987 (N_5987,N_5206,N_5271);
nor U5988 (N_5988,N_5137,N_5017);
nor U5989 (N_5989,N_5147,N_5196);
or U5990 (N_5990,N_5397,N_5377);
and U5991 (N_5991,N_5430,N_5254);
or U5992 (N_5992,N_5177,N_5127);
nand U5993 (N_5993,N_5444,N_5092);
and U5994 (N_5994,N_5226,N_5195);
and U5995 (N_5995,N_5031,N_5156);
nor U5996 (N_5996,N_5097,N_5075);
or U5997 (N_5997,N_5478,N_5054);
and U5998 (N_5998,N_5241,N_5357);
nor U5999 (N_5999,N_5063,N_5479);
and U6000 (N_6000,N_5654,N_5616);
nor U6001 (N_6001,N_5737,N_5523);
xor U6002 (N_6002,N_5912,N_5543);
and U6003 (N_6003,N_5745,N_5636);
nand U6004 (N_6004,N_5645,N_5607);
and U6005 (N_6005,N_5811,N_5780);
nor U6006 (N_6006,N_5991,N_5520);
xnor U6007 (N_6007,N_5787,N_5741);
nand U6008 (N_6008,N_5539,N_5877);
and U6009 (N_6009,N_5593,N_5582);
and U6010 (N_6010,N_5566,N_5519);
nand U6011 (N_6011,N_5958,N_5812);
nand U6012 (N_6012,N_5989,N_5659);
and U6013 (N_6013,N_5799,N_5555);
or U6014 (N_6014,N_5669,N_5621);
nor U6015 (N_6015,N_5854,N_5584);
nor U6016 (N_6016,N_5571,N_5511);
nor U6017 (N_6017,N_5966,N_5867);
or U6018 (N_6018,N_5541,N_5765);
nand U6019 (N_6019,N_5500,N_5890);
nand U6020 (N_6020,N_5944,N_5853);
or U6021 (N_6021,N_5866,N_5802);
and U6022 (N_6022,N_5684,N_5777);
nand U6023 (N_6023,N_5702,N_5893);
or U6024 (N_6024,N_5878,N_5590);
nor U6025 (N_6025,N_5530,N_5885);
and U6026 (N_6026,N_5528,N_5762);
or U6027 (N_6027,N_5864,N_5722);
or U6028 (N_6028,N_5831,N_5552);
nor U6029 (N_6029,N_5772,N_5790);
nand U6030 (N_6030,N_5792,N_5779);
nand U6031 (N_6031,N_5943,N_5588);
and U6032 (N_6032,N_5980,N_5677);
nor U6033 (N_6033,N_5691,N_5585);
nand U6034 (N_6034,N_5613,N_5969);
nor U6035 (N_6035,N_5568,N_5857);
or U6036 (N_6036,N_5567,N_5904);
or U6037 (N_6037,N_5559,N_5679);
nor U6038 (N_6038,N_5846,N_5707);
nand U6039 (N_6039,N_5518,N_5955);
or U6040 (N_6040,N_5914,N_5711);
nor U6041 (N_6041,N_5922,N_5531);
or U6042 (N_6042,N_5696,N_5766);
and U6043 (N_6043,N_5673,N_5791);
xor U6044 (N_6044,N_5892,N_5532);
nand U6045 (N_6045,N_5693,N_5968);
nand U6046 (N_6046,N_5870,N_5981);
nor U6047 (N_6047,N_5656,N_5917);
xor U6048 (N_6048,N_5538,N_5573);
and U6049 (N_6049,N_5907,N_5628);
or U6050 (N_6050,N_5658,N_5774);
and U6051 (N_6051,N_5550,N_5743);
or U6052 (N_6052,N_5839,N_5876);
or U6053 (N_6053,N_5860,N_5920);
and U6054 (N_6054,N_5634,N_5576);
and U6055 (N_6055,N_5648,N_5849);
or U6056 (N_6056,N_5661,N_5807);
nand U6057 (N_6057,N_5855,N_5882);
nor U6058 (N_6058,N_5845,N_5942);
nor U6059 (N_6059,N_5763,N_5984);
nor U6060 (N_6060,N_5606,N_5574);
nor U6061 (N_6061,N_5514,N_5879);
or U6062 (N_6062,N_5668,N_5672);
nor U6063 (N_6063,N_5665,N_5803);
and U6064 (N_6064,N_5887,N_5675);
nor U6065 (N_6065,N_5965,N_5516);
nor U6066 (N_6066,N_5861,N_5889);
nand U6067 (N_6067,N_5517,N_5577);
and U6068 (N_6068,N_5683,N_5848);
nand U6069 (N_6069,N_5947,N_5830);
or U6070 (N_6070,N_5556,N_5758);
nor U6071 (N_6071,N_5983,N_5542);
xor U6072 (N_6072,N_5662,N_5896);
nor U6073 (N_6073,N_5915,N_5631);
nand U6074 (N_6074,N_5975,N_5721);
xor U6075 (N_6075,N_5717,N_5587);
or U6076 (N_6076,N_5701,N_5624);
and U6077 (N_6077,N_5581,N_5823);
and U6078 (N_6078,N_5547,N_5757);
and U6079 (N_6079,N_5862,N_5940);
nand U6080 (N_6080,N_5881,N_5740);
xnor U6081 (N_6081,N_5509,N_5936);
nor U6082 (N_6082,N_5610,N_5923);
nand U6083 (N_6083,N_5639,N_5753);
and U6084 (N_6084,N_5689,N_5805);
nor U6085 (N_6085,N_5682,N_5789);
nand U6086 (N_6086,N_5713,N_5771);
or U6087 (N_6087,N_5651,N_5818);
xnor U6088 (N_6088,N_5733,N_5680);
and U6089 (N_6089,N_5562,N_5793);
and U6090 (N_6090,N_5918,N_5996);
nor U6091 (N_6091,N_5794,N_5508);
and U6092 (N_6092,N_5714,N_5700);
or U6093 (N_6093,N_5640,N_5545);
or U6094 (N_6094,N_5501,N_5863);
nand U6095 (N_6095,N_5769,N_5951);
and U6096 (N_6096,N_5838,N_5897);
xnor U6097 (N_6097,N_5869,N_5649);
or U6098 (N_6098,N_5934,N_5524);
nor U6099 (N_6099,N_5596,N_5629);
and U6100 (N_6100,N_5919,N_5536);
nor U6101 (N_6101,N_5956,N_5671);
nand U6102 (N_6102,N_5973,N_5641);
and U6103 (N_6103,N_5952,N_5681);
nand U6104 (N_6104,N_5899,N_5828);
and U6105 (N_6105,N_5935,N_5938);
and U6106 (N_6106,N_5505,N_5695);
and U6107 (N_6107,N_5954,N_5603);
nand U6108 (N_6108,N_5822,N_5929);
and U6109 (N_6109,N_5832,N_5716);
nand U6110 (N_6110,N_5525,N_5623);
nand U6111 (N_6111,N_5515,N_5962);
nor U6112 (N_6112,N_5865,N_5950);
nand U6113 (N_6113,N_5835,N_5997);
nor U6114 (N_6114,N_5974,N_5821);
or U6115 (N_6115,N_5959,N_5589);
nand U6116 (N_6116,N_5638,N_5670);
or U6117 (N_6117,N_5776,N_5916);
or U6118 (N_6118,N_5507,N_5548);
nor U6119 (N_6119,N_5945,N_5580);
nor U6120 (N_6120,N_5808,N_5768);
nor U6121 (N_6121,N_5786,N_5874);
or U6122 (N_6122,N_5946,N_5715);
nor U6123 (N_6123,N_5926,N_5512);
or U6124 (N_6124,N_5815,N_5971);
nor U6125 (N_6125,N_5572,N_5688);
nand U6126 (N_6126,N_5674,N_5643);
or U6127 (N_6127,N_5647,N_5570);
nor U6128 (N_6128,N_5527,N_5522);
or U6129 (N_6129,N_5637,N_5905);
nor U6130 (N_6130,N_5801,N_5728);
nand U6131 (N_6131,N_5970,N_5948);
nor U6132 (N_6132,N_5698,N_5901);
nor U6133 (N_6133,N_5978,N_5837);
and U6134 (N_6134,N_5960,N_5685);
and U6135 (N_6135,N_5502,N_5746);
or U6136 (N_6136,N_5709,N_5544);
and U6137 (N_6137,N_5626,N_5883);
nand U6138 (N_6138,N_5602,N_5827);
nor U6139 (N_6139,N_5504,N_5964);
and U6140 (N_6140,N_5609,N_5739);
nand U6141 (N_6141,N_5908,N_5903);
and U6142 (N_6142,N_5842,N_5732);
nand U6143 (N_6143,N_5731,N_5751);
and U6144 (N_6144,N_5872,N_5650);
and U6145 (N_6145,N_5804,N_5900);
nor U6146 (N_6146,N_5927,N_5612);
nand U6147 (N_6147,N_5906,N_5994);
nand U6148 (N_6148,N_5836,N_5655);
nand U6149 (N_6149,N_5859,N_5708);
nor U6150 (N_6150,N_5727,N_5937);
or U6151 (N_6151,N_5736,N_5730);
or U6152 (N_6152,N_5692,N_5586);
nor U6153 (N_6153,N_5521,N_5747);
and U6154 (N_6154,N_5987,N_5744);
and U6155 (N_6155,N_5814,N_5657);
nand U6156 (N_6156,N_5884,N_5749);
xnor U6157 (N_6157,N_5642,N_5785);
or U6158 (N_6158,N_5933,N_5597);
nor U6159 (N_6159,N_5844,N_5773);
or U6160 (N_6160,N_5699,N_5660);
nand U6161 (N_6161,N_5537,N_5601);
xnor U6162 (N_6162,N_5760,N_5949);
nand U6163 (N_6163,N_5748,N_5710);
or U6164 (N_6164,N_5913,N_5513);
or U6165 (N_6165,N_5961,N_5625);
xor U6166 (N_6166,N_5888,N_5678);
or U6167 (N_6167,N_5619,N_5506);
nand U6168 (N_6168,N_5594,N_5579);
nor U6169 (N_6169,N_5535,N_5843);
nand U6170 (N_6170,N_5614,N_5930);
or U6171 (N_6171,N_5569,N_5604);
nand U6172 (N_6172,N_5620,N_5534);
and U6173 (N_6173,N_5825,N_5939);
and U6174 (N_6174,N_5967,N_5895);
nor U6175 (N_6175,N_5925,N_5979);
or U6176 (N_6176,N_5719,N_5540);
xnor U6177 (N_6177,N_5554,N_5560);
or U6178 (N_6178,N_5990,N_5781);
and U6179 (N_6179,N_5533,N_5510);
or U6180 (N_6180,N_5756,N_5813);
and U6181 (N_6181,N_5563,N_5810);
and U6182 (N_6182,N_5826,N_5750);
or U6183 (N_6183,N_5795,N_5738);
nor U6184 (N_6184,N_5663,N_5558);
or U6185 (N_6185,N_5561,N_5622);
or U6186 (N_6186,N_5856,N_5858);
nor U6187 (N_6187,N_5608,N_5788);
nand U6188 (N_6188,N_5591,N_5986);
or U6189 (N_6189,N_5529,N_5754);
and U6190 (N_6190,N_5578,N_5690);
xor U6191 (N_6191,N_5605,N_5592);
nand U6192 (N_6192,N_5988,N_5886);
nand U6193 (N_6193,N_5898,N_5632);
or U6194 (N_6194,N_5667,N_5976);
and U6195 (N_6195,N_5551,N_5503);
nor U6196 (N_6196,N_5599,N_5783);
nor U6197 (N_6197,N_5953,N_5553);
or U6198 (N_6198,N_5932,N_5871);
nor U6199 (N_6199,N_5615,N_5850);
xor U6200 (N_6200,N_5729,N_5921);
xor U6201 (N_6201,N_5704,N_5635);
and U6202 (N_6202,N_5797,N_5646);
xor U6203 (N_6203,N_5924,N_5611);
nor U6204 (N_6204,N_5633,N_5734);
nor U6205 (N_6205,N_5820,N_5928);
nor U6206 (N_6206,N_5666,N_5720);
or U6207 (N_6207,N_5800,N_5841);
xnor U6208 (N_6208,N_5575,N_5875);
and U6209 (N_6209,N_5706,N_5724);
nand U6210 (N_6210,N_5782,N_5546);
nor U6211 (N_6211,N_5767,N_5617);
or U6212 (N_6212,N_5694,N_5873);
or U6213 (N_6213,N_5796,N_5764);
and U6214 (N_6214,N_5557,N_5653);
nor U6215 (N_6215,N_5784,N_5806);
nor U6216 (N_6216,N_5565,N_5600);
nand U6217 (N_6217,N_5992,N_5957);
or U6218 (N_6218,N_5676,N_5995);
nor U6219 (N_6219,N_5998,N_5759);
nand U6220 (N_6220,N_5618,N_5726);
and U6221 (N_6221,N_5770,N_5816);
nor U6222 (N_6222,N_5705,N_5735);
nand U6223 (N_6223,N_5829,N_5902);
or U6224 (N_6224,N_5868,N_5798);
or U6225 (N_6225,N_5644,N_5595);
or U6226 (N_6226,N_5999,N_5834);
nand U6227 (N_6227,N_5909,N_5712);
nand U6228 (N_6228,N_5977,N_5809);
or U6229 (N_6229,N_5664,N_5775);
nand U6230 (N_6230,N_5564,N_5652);
nor U6231 (N_6231,N_5833,N_5819);
or U6232 (N_6232,N_5526,N_5941);
and U6233 (N_6233,N_5824,N_5851);
nand U6234 (N_6234,N_5549,N_5985);
and U6235 (N_6235,N_5963,N_5891);
and U6236 (N_6236,N_5778,N_5982);
nand U6237 (N_6237,N_5627,N_5761);
nand U6238 (N_6238,N_5817,N_5583);
nor U6239 (N_6239,N_5755,N_5993);
nor U6240 (N_6240,N_5742,N_5972);
or U6241 (N_6241,N_5752,N_5840);
and U6242 (N_6242,N_5894,N_5725);
and U6243 (N_6243,N_5852,N_5687);
nor U6244 (N_6244,N_5686,N_5911);
or U6245 (N_6245,N_5910,N_5598);
or U6246 (N_6246,N_5703,N_5697);
nand U6247 (N_6247,N_5723,N_5880);
and U6248 (N_6248,N_5718,N_5931);
nor U6249 (N_6249,N_5847,N_5630);
xnor U6250 (N_6250,N_5903,N_5965);
and U6251 (N_6251,N_5991,N_5818);
nor U6252 (N_6252,N_5627,N_5646);
and U6253 (N_6253,N_5943,N_5945);
xnor U6254 (N_6254,N_5732,N_5730);
nor U6255 (N_6255,N_5729,N_5671);
nor U6256 (N_6256,N_5952,N_5884);
nand U6257 (N_6257,N_5708,N_5670);
nand U6258 (N_6258,N_5808,N_5631);
and U6259 (N_6259,N_5562,N_5544);
xnor U6260 (N_6260,N_5533,N_5580);
or U6261 (N_6261,N_5500,N_5968);
or U6262 (N_6262,N_5557,N_5856);
or U6263 (N_6263,N_5547,N_5768);
nor U6264 (N_6264,N_5557,N_5914);
nand U6265 (N_6265,N_5578,N_5732);
and U6266 (N_6266,N_5690,N_5946);
xor U6267 (N_6267,N_5934,N_5848);
and U6268 (N_6268,N_5727,N_5604);
or U6269 (N_6269,N_5937,N_5608);
nand U6270 (N_6270,N_5622,N_5563);
nor U6271 (N_6271,N_5757,N_5946);
and U6272 (N_6272,N_5611,N_5739);
nor U6273 (N_6273,N_5976,N_5572);
nand U6274 (N_6274,N_5728,N_5755);
nand U6275 (N_6275,N_5763,N_5975);
nand U6276 (N_6276,N_5964,N_5522);
and U6277 (N_6277,N_5908,N_5538);
nor U6278 (N_6278,N_5719,N_5746);
xor U6279 (N_6279,N_5950,N_5559);
xnor U6280 (N_6280,N_5631,N_5855);
xor U6281 (N_6281,N_5620,N_5916);
or U6282 (N_6282,N_5855,N_5690);
and U6283 (N_6283,N_5548,N_5588);
nor U6284 (N_6284,N_5647,N_5770);
or U6285 (N_6285,N_5961,N_5903);
and U6286 (N_6286,N_5990,N_5716);
xnor U6287 (N_6287,N_5690,N_5715);
nand U6288 (N_6288,N_5502,N_5799);
or U6289 (N_6289,N_5784,N_5909);
nor U6290 (N_6290,N_5517,N_5942);
or U6291 (N_6291,N_5596,N_5991);
and U6292 (N_6292,N_5942,N_5921);
or U6293 (N_6293,N_5698,N_5919);
nand U6294 (N_6294,N_5893,N_5906);
nand U6295 (N_6295,N_5875,N_5754);
nand U6296 (N_6296,N_5716,N_5846);
xor U6297 (N_6297,N_5967,N_5613);
nor U6298 (N_6298,N_5561,N_5502);
or U6299 (N_6299,N_5570,N_5532);
nor U6300 (N_6300,N_5574,N_5525);
xnor U6301 (N_6301,N_5822,N_5631);
or U6302 (N_6302,N_5896,N_5516);
and U6303 (N_6303,N_5741,N_5770);
nand U6304 (N_6304,N_5526,N_5696);
nand U6305 (N_6305,N_5996,N_5892);
nor U6306 (N_6306,N_5943,N_5638);
nor U6307 (N_6307,N_5724,N_5650);
xnor U6308 (N_6308,N_5759,N_5815);
nand U6309 (N_6309,N_5601,N_5583);
xnor U6310 (N_6310,N_5843,N_5853);
and U6311 (N_6311,N_5928,N_5513);
nand U6312 (N_6312,N_5764,N_5826);
nand U6313 (N_6313,N_5760,N_5653);
xnor U6314 (N_6314,N_5946,N_5543);
nand U6315 (N_6315,N_5906,N_5896);
nand U6316 (N_6316,N_5542,N_5562);
xnor U6317 (N_6317,N_5856,N_5711);
or U6318 (N_6318,N_5705,N_5516);
xnor U6319 (N_6319,N_5834,N_5846);
or U6320 (N_6320,N_5759,N_5653);
and U6321 (N_6321,N_5690,N_5983);
and U6322 (N_6322,N_5612,N_5564);
nor U6323 (N_6323,N_5949,N_5792);
nand U6324 (N_6324,N_5725,N_5695);
nand U6325 (N_6325,N_5919,N_5947);
xnor U6326 (N_6326,N_5665,N_5727);
nor U6327 (N_6327,N_5828,N_5608);
or U6328 (N_6328,N_5996,N_5847);
and U6329 (N_6329,N_5886,N_5822);
nor U6330 (N_6330,N_5759,N_5664);
nand U6331 (N_6331,N_5905,N_5514);
nor U6332 (N_6332,N_5751,N_5754);
nor U6333 (N_6333,N_5962,N_5504);
nor U6334 (N_6334,N_5651,N_5922);
nand U6335 (N_6335,N_5520,N_5631);
and U6336 (N_6336,N_5559,N_5850);
and U6337 (N_6337,N_5598,N_5905);
and U6338 (N_6338,N_5864,N_5784);
nor U6339 (N_6339,N_5973,N_5707);
and U6340 (N_6340,N_5554,N_5746);
nor U6341 (N_6341,N_5869,N_5860);
nor U6342 (N_6342,N_5872,N_5816);
and U6343 (N_6343,N_5542,N_5729);
and U6344 (N_6344,N_5948,N_5719);
or U6345 (N_6345,N_5713,N_5846);
nand U6346 (N_6346,N_5746,N_5834);
nand U6347 (N_6347,N_5644,N_5942);
or U6348 (N_6348,N_5539,N_5582);
or U6349 (N_6349,N_5773,N_5591);
nand U6350 (N_6350,N_5776,N_5995);
or U6351 (N_6351,N_5852,N_5816);
nor U6352 (N_6352,N_5699,N_5923);
nand U6353 (N_6353,N_5854,N_5571);
xnor U6354 (N_6354,N_5883,N_5959);
and U6355 (N_6355,N_5905,N_5866);
nand U6356 (N_6356,N_5651,N_5787);
nor U6357 (N_6357,N_5842,N_5690);
nand U6358 (N_6358,N_5631,N_5812);
nand U6359 (N_6359,N_5652,N_5839);
or U6360 (N_6360,N_5718,N_5984);
nor U6361 (N_6361,N_5507,N_5586);
nand U6362 (N_6362,N_5964,N_5646);
nand U6363 (N_6363,N_5850,N_5587);
nor U6364 (N_6364,N_5513,N_5999);
nand U6365 (N_6365,N_5969,N_5946);
xnor U6366 (N_6366,N_5808,N_5585);
nor U6367 (N_6367,N_5695,N_5919);
nand U6368 (N_6368,N_5861,N_5762);
nand U6369 (N_6369,N_5828,N_5772);
or U6370 (N_6370,N_5870,N_5735);
nor U6371 (N_6371,N_5863,N_5712);
and U6372 (N_6372,N_5785,N_5848);
nor U6373 (N_6373,N_5568,N_5759);
xor U6374 (N_6374,N_5568,N_5564);
nand U6375 (N_6375,N_5752,N_5820);
or U6376 (N_6376,N_5773,N_5870);
nor U6377 (N_6377,N_5532,N_5995);
nand U6378 (N_6378,N_5945,N_5835);
and U6379 (N_6379,N_5729,N_5694);
and U6380 (N_6380,N_5970,N_5641);
and U6381 (N_6381,N_5979,N_5661);
xnor U6382 (N_6382,N_5512,N_5964);
or U6383 (N_6383,N_5696,N_5553);
and U6384 (N_6384,N_5863,N_5885);
and U6385 (N_6385,N_5807,N_5755);
nand U6386 (N_6386,N_5749,N_5893);
nand U6387 (N_6387,N_5691,N_5636);
and U6388 (N_6388,N_5897,N_5638);
or U6389 (N_6389,N_5877,N_5607);
xor U6390 (N_6390,N_5633,N_5804);
nor U6391 (N_6391,N_5746,N_5929);
and U6392 (N_6392,N_5568,N_5796);
and U6393 (N_6393,N_5982,N_5810);
nand U6394 (N_6394,N_5998,N_5792);
nand U6395 (N_6395,N_5602,N_5954);
xnor U6396 (N_6396,N_5846,N_5689);
nor U6397 (N_6397,N_5633,N_5624);
or U6398 (N_6398,N_5816,N_5801);
nand U6399 (N_6399,N_5869,N_5573);
nand U6400 (N_6400,N_5671,N_5990);
or U6401 (N_6401,N_5968,N_5790);
or U6402 (N_6402,N_5814,N_5640);
nor U6403 (N_6403,N_5805,N_5627);
or U6404 (N_6404,N_5855,N_5511);
or U6405 (N_6405,N_5525,N_5515);
or U6406 (N_6406,N_5986,N_5566);
nand U6407 (N_6407,N_5916,N_5875);
nor U6408 (N_6408,N_5783,N_5972);
nor U6409 (N_6409,N_5847,N_5579);
xnor U6410 (N_6410,N_5758,N_5854);
or U6411 (N_6411,N_5870,N_5914);
nand U6412 (N_6412,N_5581,N_5668);
nor U6413 (N_6413,N_5658,N_5561);
nor U6414 (N_6414,N_5904,N_5671);
xnor U6415 (N_6415,N_5900,N_5997);
and U6416 (N_6416,N_5931,N_5579);
and U6417 (N_6417,N_5560,N_5901);
xnor U6418 (N_6418,N_5867,N_5876);
nand U6419 (N_6419,N_5522,N_5566);
xor U6420 (N_6420,N_5676,N_5576);
and U6421 (N_6421,N_5846,N_5619);
nand U6422 (N_6422,N_5571,N_5523);
nand U6423 (N_6423,N_5808,N_5885);
nor U6424 (N_6424,N_5539,N_5832);
nor U6425 (N_6425,N_5504,N_5590);
nand U6426 (N_6426,N_5737,N_5869);
or U6427 (N_6427,N_5812,N_5758);
xnor U6428 (N_6428,N_5535,N_5894);
or U6429 (N_6429,N_5999,N_5709);
nor U6430 (N_6430,N_5670,N_5847);
or U6431 (N_6431,N_5732,N_5984);
nor U6432 (N_6432,N_5875,N_5889);
and U6433 (N_6433,N_5734,N_5807);
nand U6434 (N_6434,N_5541,N_5556);
xor U6435 (N_6435,N_5701,N_5825);
xnor U6436 (N_6436,N_5606,N_5848);
nand U6437 (N_6437,N_5595,N_5717);
or U6438 (N_6438,N_5988,N_5810);
nand U6439 (N_6439,N_5832,N_5709);
and U6440 (N_6440,N_5707,N_5944);
xor U6441 (N_6441,N_5785,N_5596);
and U6442 (N_6442,N_5639,N_5546);
nor U6443 (N_6443,N_5836,N_5948);
nand U6444 (N_6444,N_5851,N_5513);
or U6445 (N_6445,N_5851,N_5755);
and U6446 (N_6446,N_5955,N_5563);
nand U6447 (N_6447,N_5672,N_5763);
or U6448 (N_6448,N_5754,N_5685);
and U6449 (N_6449,N_5857,N_5821);
or U6450 (N_6450,N_5885,N_5759);
nand U6451 (N_6451,N_5899,N_5982);
or U6452 (N_6452,N_5580,N_5812);
and U6453 (N_6453,N_5640,N_5657);
nand U6454 (N_6454,N_5707,N_5856);
and U6455 (N_6455,N_5944,N_5951);
nand U6456 (N_6456,N_5660,N_5861);
nand U6457 (N_6457,N_5545,N_5841);
nor U6458 (N_6458,N_5628,N_5607);
and U6459 (N_6459,N_5869,N_5644);
xor U6460 (N_6460,N_5960,N_5734);
and U6461 (N_6461,N_5745,N_5855);
or U6462 (N_6462,N_5828,N_5709);
or U6463 (N_6463,N_5881,N_5966);
nor U6464 (N_6464,N_5661,N_5683);
and U6465 (N_6465,N_5528,N_5976);
nor U6466 (N_6466,N_5823,N_5670);
nor U6467 (N_6467,N_5944,N_5564);
and U6468 (N_6468,N_5504,N_5893);
nand U6469 (N_6469,N_5855,N_5709);
or U6470 (N_6470,N_5843,N_5561);
and U6471 (N_6471,N_5617,N_5706);
and U6472 (N_6472,N_5962,N_5986);
or U6473 (N_6473,N_5919,N_5596);
and U6474 (N_6474,N_5504,N_5897);
or U6475 (N_6475,N_5994,N_5793);
nor U6476 (N_6476,N_5795,N_5881);
nor U6477 (N_6477,N_5947,N_5982);
and U6478 (N_6478,N_5635,N_5794);
or U6479 (N_6479,N_5839,N_5825);
and U6480 (N_6480,N_5945,N_5940);
and U6481 (N_6481,N_5651,N_5722);
nand U6482 (N_6482,N_5943,N_5755);
nand U6483 (N_6483,N_5886,N_5663);
xor U6484 (N_6484,N_5829,N_5694);
nand U6485 (N_6485,N_5713,N_5847);
nand U6486 (N_6486,N_5633,N_5701);
nor U6487 (N_6487,N_5961,N_5603);
nand U6488 (N_6488,N_5743,N_5727);
and U6489 (N_6489,N_5607,N_5980);
xor U6490 (N_6490,N_5847,N_5614);
or U6491 (N_6491,N_5910,N_5713);
nand U6492 (N_6492,N_5571,N_5934);
or U6493 (N_6493,N_5834,N_5907);
nor U6494 (N_6494,N_5968,N_5751);
or U6495 (N_6495,N_5763,N_5684);
nor U6496 (N_6496,N_5735,N_5570);
nor U6497 (N_6497,N_5763,N_5964);
nor U6498 (N_6498,N_5787,N_5977);
nor U6499 (N_6499,N_5500,N_5670);
nand U6500 (N_6500,N_6310,N_6420);
nand U6501 (N_6501,N_6052,N_6419);
and U6502 (N_6502,N_6188,N_6351);
or U6503 (N_6503,N_6013,N_6426);
xor U6504 (N_6504,N_6380,N_6169);
xor U6505 (N_6505,N_6308,N_6312);
nor U6506 (N_6506,N_6099,N_6112);
and U6507 (N_6507,N_6360,N_6243);
nand U6508 (N_6508,N_6039,N_6444);
and U6509 (N_6509,N_6495,N_6359);
nand U6510 (N_6510,N_6323,N_6059);
xnor U6511 (N_6511,N_6375,N_6027);
or U6512 (N_6512,N_6441,N_6081);
or U6513 (N_6513,N_6305,N_6407);
nand U6514 (N_6514,N_6125,N_6181);
nand U6515 (N_6515,N_6050,N_6185);
or U6516 (N_6516,N_6452,N_6488);
or U6517 (N_6517,N_6491,N_6131);
and U6518 (N_6518,N_6272,N_6124);
nand U6519 (N_6519,N_6378,N_6071);
nand U6520 (N_6520,N_6172,N_6321);
nand U6521 (N_6521,N_6240,N_6073);
or U6522 (N_6522,N_6034,N_6428);
nor U6523 (N_6523,N_6347,N_6306);
and U6524 (N_6524,N_6342,N_6412);
or U6525 (N_6525,N_6033,N_6108);
xnor U6526 (N_6526,N_6416,N_6037);
xor U6527 (N_6527,N_6403,N_6228);
and U6528 (N_6528,N_6004,N_6182);
nand U6529 (N_6529,N_6277,N_6390);
nor U6530 (N_6530,N_6090,N_6411);
nor U6531 (N_6531,N_6436,N_6496);
nor U6532 (N_6532,N_6450,N_6137);
and U6533 (N_6533,N_6054,N_6348);
xor U6534 (N_6534,N_6022,N_6468);
nor U6535 (N_6535,N_6386,N_6106);
xor U6536 (N_6536,N_6116,N_6275);
and U6537 (N_6537,N_6232,N_6060);
or U6538 (N_6538,N_6366,N_6269);
or U6539 (N_6539,N_6025,N_6015);
nor U6540 (N_6540,N_6330,N_6104);
xor U6541 (N_6541,N_6457,N_6126);
or U6542 (N_6542,N_6211,N_6461);
nor U6543 (N_6543,N_6417,N_6362);
nor U6544 (N_6544,N_6118,N_6455);
nor U6545 (N_6545,N_6463,N_6156);
nand U6546 (N_6546,N_6371,N_6418);
or U6547 (N_6547,N_6353,N_6437);
nor U6548 (N_6548,N_6247,N_6499);
nor U6549 (N_6549,N_6194,N_6467);
nor U6550 (N_6550,N_6460,N_6497);
and U6551 (N_6551,N_6421,N_6476);
and U6552 (N_6552,N_6024,N_6392);
or U6553 (N_6553,N_6307,N_6096);
and U6554 (N_6554,N_6264,N_6120);
nor U6555 (N_6555,N_6408,N_6248);
nor U6556 (N_6556,N_6079,N_6021);
nor U6557 (N_6557,N_6216,N_6260);
nor U6558 (N_6558,N_6374,N_6334);
xor U6559 (N_6559,N_6414,N_6433);
nor U6560 (N_6560,N_6242,N_6173);
xor U6561 (N_6561,N_6494,N_6431);
xnor U6562 (N_6562,N_6128,N_6335);
and U6563 (N_6563,N_6014,N_6432);
nand U6564 (N_6564,N_6162,N_6427);
or U6565 (N_6565,N_6202,N_6447);
nor U6566 (N_6566,N_6332,N_6008);
or U6567 (N_6567,N_6413,N_6017);
or U6568 (N_6568,N_6175,N_6029);
nand U6569 (N_6569,N_6152,N_6134);
nor U6570 (N_6570,N_6195,N_6398);
and U6571 (N_6571,N_6477,N_6296);
nor U6572 (N_6572,N_6214,N_6006);
or U6573 (N_6573,N_6459,N_6192);
or U6574 (N_6574,N_6235,N_6102);
and U6575 (N_6575,N_6114,N_6258);
nand U6576 (N_6576,N_6231,N_6227);
nand U6577 (N_6577,N_6075,N_6254);
xnor U6578 (N_6578,N_6011,N_6067);
nand U6579 (N_6579,N_6047,N_6139);
or U6580 (N_6580,N_6395,N_6357);
nand U6581 (N_6581,N_6005,N_6379);
nor U6582 (N_6582,N_6087,N_6474);
nor U6583 (N_6583,N_6291,N_6063);
or U6584 (N_6584,N_6123,N_6145);
nand U6585 (N_6585,N_6391,N_6262);
xnor U6586 (N_6586,N_6072,N_6385);
nor U6587 (N_6587,N_6387,N_6184);
nor U6588 (N_6588,N_6141,N_6191);
or U6589 (N_6589,N_6328,N_6485);
nor U6590 (N_6590,N_6065,N_6148);
and U6591 (N_6591,N_6209,N_6201);
nand U6592 (N_6592,N_6253,N_6121);
xor U6593 (N_6593,N_6239,N_6055);
nor U6594 (N_6594,N_6405,N_6249);
and U6595 (N_6595,N_6035,N_6278);
or U6596 (N_6596,N_6367,N_6281);
and U6597 (N_6597,N_6113,N_6489);
and U6598 (N_6598,N_6032,N_6294);
nand U6599 (N_6599,N_6160,N_6225);
nor U6600 (N_6600,N_6205,N_6293);
nand U6601 (N_6601,N_6446,N_6265);
or U6602 (N_6602,N_6333,N_6095);
or U6603 (N_6603,N_6337,N_6180);
nor U6604 (N_6604,N_6373,N_6163);
or U6605 (N_6605,N_6479,N_6422);
nor U6606 (N_6606,N_6161,N_6402);
xnor U6607 (N_6607,N_6498,N_6028);
xnor U6608 (N_6608,N_6316,N_6224);
or U6609 (N_6609,N_6443,N_6016);
nand U6610 (N_6610,N_6368,N_6273);
nor U6611 (N_6611,N_6044,N_6127);
nand U6612 (N_6612,N_6010,N_6056);
xnor U6613 (N_6613,N_6001,N_6199);
nor U6614 (N_6614,N_6100,N_6434);
xor U6615 (N_6615,N_6178,N_6279);
nor U6616 (N_6616,N_6057,N_6300);
nor U6617 (N_6617,N_6136,N_6492);
or U6618 (N_6618,N_6110,N_6345);
and U6619 (N_6619,N_6343,N_6089);
nand U6620 (N_6620,N_6149,N_6266);
and U6621 (N_6621,N_6062,N_6023);
or U6622 (N_6622,N_6221,N_6361);
nor U6623 (N_6623,N_6097,N_6190);
nand U6624 (N_6624,N_6170,N_6174);
and U6625 (N_6625,N_6066,N_6338);
nor U6626 (N_6626,N_6233,N_6241);
nand U6627 (N_6627,N_6246,N_6210);
and U6628 (N_6628,N_6256,N_6440);
and U6629 (N_6629,N_6215,N_6168);
and U6630 (N_6630,N_6255,N_6030);
and U6631 (N_6631,N_6200,N_6103);
nor U6632 (N_6632,N_6471,N_6206);
and U6633 (N_6633,N_6478,N_6142);
xor U6634 (N_6634,N_6197,N_6171);
nand U6635 (N_6635,N_6074,N_6179);
and U6636 (N_6636,N_6287,N_6208);
or U6637 (N_6637,N_6276,N_6372);
nor U6638 (N_6638,N_6166,N_6115);
nor U6639 (N_6639,N_6456,N_6198);
and U6640 (N_6640,N_6158,N_6018);
xor U6641 (N_6641,N_6263,N_6245);
or U6642 (N_6642,N_6451,N_6311);
or U6643 (N_6643,N_6290,N_6314);
nand U6644 (N_6644,N_6250,N_6389);
xor U6645 (N_6645,N_6061,N_6122);
nand U6646 (N_6646,N_6085,N_6448);
or U6647 (N_6647,N_6458,N_6352);
and U6648 (N_6648,N_6473,N_6077);
and U6649 (N_6649,N_6346,N_6219);
and U6650 (N_6650,N_6318,N_6466);
and U6651 (N_6651,N_6322,N_6155);
nand U6652 (N_6652,N_6292,N_6482);
or U6653 (N_6653,N_6415,N_6226);
xor U6654 (N_6654,N_6327,N_6020);
or U6655 (N_6655,N_6135,N_6252);
xnor U6656 (N_6656,N_6370,N_6355);
nor U6657 (N_6657,N_6177,N_6289);
and U6658 (N_6658,N_6117,N_6094);
or U6659 (N_6659,N_6339,N_6220);
or U6660 (N_6660,N_6012,N_6237);
xor U6661 (N_6661,N_6109,N_6381);
xnor U6662 (N_6662,N_6302,N_6167);
nor U6663 (N_6663,N_6383,N_6404);
and U6664 (N_6664,N_6165,N_6406);
and U6665 (N_6665,N_6146,N_6119);
and U6666 (N_6666,N_6157,N_6377);
nor U6667 (N_6667,N_6423,N_6326);
nand U6668 (N_6668,N_6299,N_6341);
nand U6669 (N_6669,N_6007,N_6144);
nor U6670 (N_6670,N_6396,N_6217);
xor U6671 (N_6671,N_6331,N_6189);
nor U6672 (N_6672,N_6401,N_6078);
nand U6673 (N_6673,N_6435,N_6356);
xnor U6674 (N_6674,N_6193,N_6251);
and U6675 (N_6675,N_6069,N_6212);
nor U6676 (N_6676,N_6105,N_6349);
xor U6677 (N_6677,N_6301,N_6397);
or U6678 (N_6678,N_6439,N_6230);
nor U6679 (N_6679,N_6469,N_6133);
and U6680 (N_6680,N_6438,N_6288);
xor U6681 (N_6681,N_6150,N_6064);
nand U6682 (N_6682,N_6138,N_6453);
nor U6683 (N_6683,N_6303,N_6049);
and U6684 (N_6684,N_6130,N_6388);
nand U6685 (N_6685,N_6143,N_6261);
nor U6686 (N_6686,N_6462,N_6369);
xor U6687 (N_6687,N_6045,N_6358);
nand U6688 (N_6688,N_6487,N_6223);
and U6689 (N_6689,N_6207,N_6019);
and U6690 (N_6690,N_6259,N_6236);
nor U6691 (N_6691,N_6042,N_6297);
nand U6692 (N_6692,N_6465,N_6229);
and U6693 (N_6693,N_6298,N_6445);
nor U6694 (N_6694,N_6313,N_6365);
and U6695 (N_6695,N_6329,N_6410);
nand U6696 (N_6696,N_6304,N_6084);
nor U6697 (N_6697,N_6394,N_6176);
nand U6698 (N_6698,N_6058,N_6092);
and U6699 (N_6699,N_6282,N_6043);
and U6700 (N_6700,N_6083,N_6430);
nor U6701 (N_6701,N_6480,N_6009);
nand U6702 (N_6702,N_6336,N_6164);
nand U6703 (N_6703,N_6257,N_6154);
or U6704 (N_6704,N_6222,N_6040);
or U6705 (N_6705,N_6093,N_6484);
nand U6706 (N_6706,N_6268,N_6442);
and U6707 (N_6707,N_6384,N_6036);
nor U6708 (N_6708,N_6286,N_6325);
nor U6709 (N_6709,N_6283,N_6376);
and U6710 (N_6710,N_6000,N_6234);
xnor U6711 (N_6711,N_6159,N_6213);
nor U6712 (N_6712,N_6101,N_6354);
xnor U6713 (N_6713,N_6424,N_6086);
nand U6714 (N_6714,N_6151,N_6107);
and U6715 (N_6715,N_6284,N_6393);
nand U6716 (N_6716,N_6350,N_6409);
xnor U6717 (N_6717,N_6132,N_6280);
nand U6718 (N_6718,N_6051,N_6319);
or U6719 (N_6719,N_6481,N_6046);
nand U6720 (N_6720,N_6003,N_6204);
and U6721 (N_6721,N_6475,N_6098);
and U6722 (N_6722,N_6324,N_6068);
xnor U6723 (N_6723,N_6203,N_6076);
nand U6724 (N_6724,N_6267,N_6271);
or U6725 (N_6725,N_6002,N_6317);
and U6726 (N_6726,N_6186,N_6238);
nor U6727 (N_6727,N_6295,N_6340);
and U6728 (N_6728,N_6309,N_6449);
and U6729 (N_6729,N_6270,N_6041);
nor U6730 (N_6730,N_6274,N_6082);
xnor U6731 (N_6731,N_6031,N_6454);
xor U6732 (N_6732,N_6364,N_6425);
or U6733 (N_6733,N_6490,N_6111);
xnor U6734 (N_6734,N_6429,N_6218);
nand U6735 (N_6735,N_6196,N_6285);
or U6736 (N_6736,N_6183,N_6187);
and U6737 (N_6737,N_6363,N_6244);
and U6738 (N_6738,N_6400,N_6038);
or U6739 (N_6739,N_6320,N_6026);
nand U6740 (N_6740,N_6382,N_6088);
or U6741 (N_6741,N_6147,N_6493);
xnor U6742 (N_6742,N_6344,N_6140);
or U6743 (N_6743,N_6053,N_6129);
nand U6744 (N_6744,N_6470,N_6464);
or U6745 (N_6745,N_6091,N_6315);
nor U6746 (N_6746,N_6080,N_6153);
nor U6747 (N_6747,N_6399,N_6483);
or U6748 (N_6748,N_6486,N_6472);
and U6749 (N_6749,N_6048,N_6070);
nand U6750 (N_6750,N_6248,N_6324);
nor U6751 (N_6751,N_6261,N_6387);
and U6752 (N_6752,N_6339,N_6369);
xnor U6753 (N_6753,N_6437,N_6179);
nand U6754 (N_6754,N_6280,N_6282);
and U6755 (N_6755,N_6130,N_6359);
or U6756 (N_6756,N_6453,N_6028);
and U6757 (N_6757,N_6354,N_6173);
nor U6758 (N_6758,N_6477,N_6367);
or U6759 (N_6759,N_6412,N_6270);
xnor U6760 (N_6760,N_6303,N_6244);
nand U6761 (N_6761,N_6350,N_6005);
nand U6762 (N_6762,N_6234,N_6156);
or U6763 (N_6763,N_6419,N_6107);
nand U6764 (N_6764,N_6209,N_6361);
and U6765 (N_6765,N_6222,N_6158);
and U6766 (N_6766,N_6228,N_6104);
nor U6767 (N_6767,N_6002,N_6117);
and U6768 (N_6768,N_6368,N_6010);
and U6769 (N_6769,N_6252,N_6123);
or U6770 (N_6770,N_6289,N_6235);
or U6771 (N_6771,N_6038,N_6116);
xnor U6772 (N_6772,N_6090,N_6214);
xor U6773 (N_6773,N_6007,N_6263);
nand U6774 (N_6774,N_6084,N_6178);
nor U6775 (N_6775,N_6186,N_6032);
nor U6776 (N_6776,N_6354,N_6274);
nand U6777 (N_6777,N_6356,N_6436);
nor U6778 (N_6778,N_6076,N_6180);
xor U6779 (N_6779,N_6018,N_6464);
nand U6780 (N_6780,N_6182,N_6433);
and U6781 (N_6781,N_6147,N_6475);
or U6782 (N_6782,N_6223,N_6443);
nand U6783 (N_6783,N_6310,N_6362);
or U6784 (N_6784,N_6017,N_6363);
or U6785 (N_6785,N_6441,N_6157);
or U6786 (N_6786,N_6373,N_6391);
and U6787 (N_6787,N_6320,N_6144);
or U6788 (N_6788,N_6094,N_6025);
and U6789 (N_6789,N_6374,N_6109);
or U6790 (N_6790,N_6262,N_6078);
and U6791 (N_6791,N_6467,N_6034);
and U6792 (N_6792,N_6197,N_6175);
nand U6793 (N_6793,N_6277,N_6430);
and U6794 (N_6794,N_6292,N_6092);
nand U6795 (N_6795,N_6117,N_6324);
and U6796 (N_6796,N_6431,N_6165);
and U6797 (N_6797,N_6203,N_6347);
and U6798 (N_6798,N_6149,N_6444);
and U6799 (N_6799,N_6024,N_6043);
and U6800 (N_6800,N_6045,N_6377);
nor U6801 (N_6801,N_6051,N_6244);
xnor U6802 (N_6802,N_6483,N_6159);
nor U6803 (N_6803,N_6433,N_6028);
or U6804 (N_6804,N_6146,N_6294);
and U6805 (N_6805,N_6084,N_6414);
nand U6806 (N_6806,N_6302,N_6368);
or U6807 (N_6807,N_6093,N_6193);
and U6808 (N_6808,N_6475,N_6262);
nor U6809 (N_6809,N_6123,N_6455);
nand U6810 (N_6810,N_6161,N_6065);
or U6811 (N_6811,N_6095,N_6317);
xor U6812 (N_6812,N_6213,N_6271);
and U6813 (N_6813,N_6085,N_6277);
and U6814 (N_6814,N_6375,N_6385);
xor U6815 (N_6815,N_6092,N_6328);
nand U6816 (N_6816,N_6303,N_6334);
or U6817 (N_6817,N_6164,N_6435);
or U6818 (N_6818,N_6222,N_6096);
nor U6819 (N_6819,N_6056,N_6489);
nand U6820 (N_6820,N_6328,N_6300);
and U6821 (N_6821,N_6322,N_6368);
xnor U6822 (N_6822,N_6076,N_6021);
nor U6823 (N_6823,N_6004,N_6492);
nor U6824 (N_6824,N_6370,N_6365);
and U6825 (N_6825,N_6078,N_6219);
nor U6826 (N_6826,N_6300,N_6473);
nor U6827 (N_6827,N_6044,N_6400);
nand U6828 (N_6828,N_6381,N_6362);
and U6829 (N_6829,N_6013,N_6212);
or U6830 (N_6830,N_6128,N_6420);
or U6831 (N_6831,N_6102,N_6021);
or U6832 (N_6832,N_6335,N_6109);
xnor U6833 (N_6833,N_6112,N_6421);
xor U6834 (N_6834,N_6043,N_6298);
or U6835 (N_6835,N_6409,N_6010);
xor U6836 (N_6836,N_6183,N_6461);
xnor U6837 (N_6837,N_6232,N_6021);
nand U6838 (N_6838,N_6442,N_6337);
nor U6839 (N_6839,N_6229,N_6008);
and U6840 (N_6840,N_6252,N_6416);
nand U6841 (N_6841,N_6186,N_6163);
and U6842 (N_6842,N_6467,N_6446);
and U6843 (N_6843,N_6024,N_6415);
nor U6844 (N_6844,N_6253,N_6158);
nand U6845 (N_6845,N_6138,N_6388);
and U6846 (N_6846,N_6260,N_6297);
and U6847 (N_6847,N_6166,N_6290);
nand U6848 (N_6848,N_6394,N_6357);
nand U6849 (N_6849,N_6477,N_6122);
or U6850 (N_6850,N_6296,N_6028);
or U6851 (N_6851,N_6079,N_6405);
or U6852 (N_6852,N_6117,N_6168);
nand U6853 (N_6853,N_6454,N_6499);
nor U6854 (N_6854,N_6231,N_6308);
nor U6855 (N_6855,N_6221,N_6239);
and U6856 (N_6856,N_6386,N_6394);
xnor U6857 (N_6857,N_6275,N_6304);
nor U6858 (N_6858,N_6424,N_6376);
xnor U6859 (N_6859,N_6004,N_6369);
xor U6860 (N_6860,N_6482,N_6101);
nor U6861 (N_6861,N_6122,N_6010);
nor U6862 (N_6862,N_6401,N_6187);
and U6863 (N_6863,N_6103,N_6047);
or U6864 (N_6864,N_6011,N_6029);
nor U6865 (N_6865,N_6105,N_6111);
xnor U6866 (N_6866,N_6247,N_6152);
nand U6867 (N_6867,N_6130,N_6416);
or U6868 (N_6868,N_6420,N_6314);
and U6869 (N_6869,N_6185,N_6270);
and U6870 (N_6870,N_6323,N_6345);
nand U6871 (N_6871,N_6181,N_6217);
and U6872 (N_6872,N_6262,N_6299);
or U6873 (N_6873,N_6108,N_6188);
and U6874 (N_6874,N_6463,N_6389);
nand U6875 (N_6875,N_6452,N_6086);
and U6876 (N_6876,N_6281,N_6053);
and U6877 (N_6877,N_6365,N_6350);
or U6878 (N_6878,N_6048,N_6247);
xnor U6879 (N_6879,N_6036,N_6249);
xor U6880 (N_6880,N_6399,N_6197);
and U6881 (N_6881,N_6216,N_6058);
or U6882 (N_6882,N_6455,N_6461);
and U6883 (N_6883,N_6408,N_6456);
xor U6884 (N_6884,N_6371,N_6399);
nor U6885 (N_6885,N_6245,N_6261);
or U6886 (N_6886,N_6394,N_6481);
nor U6887 (N_6887,N_6221,N_6030);
or U6888 (N_6888,N_6441,N_6380);
nor U6889 (N_6889,N_6288,N_6277);
nand U6890 (N_6890,N_6055,N_6451);
and U6891 (N_6891,N_6456,N_6187);
nor U6892 (N_6892,N_6200,N_6301);
xnor U6893 (N_6893,N_6122,N_6428);
nand U6894 (N_6894,N_6123,N_6325);
and U6895 (N_6895,N_6367,N_6125);
and U6896 (N_6896,N_6147,N_6311);
nor U6897 (N_6897,N_6272,N_6367);
nand U6898 (N_6898,N_6126,N_6130);
nand U6899 (N_6899,N_6203,N_6176);
nand U6900 (N_6900,N_6069,N_6420);
and U6901 (N_6901,N_6436,N_6101);
nand U6902 (N_6902,N_6237,N_6097);
nand U6903 (N_6903,N_6154,N_6080);
nand U6904 (N_6904,N_6429,N_6302);
and U6905 (N_6905,N_6493,N_6087);
xnor U6906 (N_6906,N_6470,N_6298);
xnor U6907 (N_6907,N_6288,N_6120);
nand U6908 (N_6908,N_6327,N_6199);
nor U6909 (N_6909,N_6390,N_6062);
and U6910 (N_6910,N_6467,N_6089);
nand U6911 (N_6911,N_6362,N_6359);
xnor U6912 (N_6912,N_6001,N_6332);
xor U6913 (N_6913,N_6171,N_6014);
xor U6914 (N_6914,N_6014,N_6225);
nand U6915 (N_6915,N_6442,N_6063);
or U6916 (N_6916,N_6026,N_6213);
xor U6917 (N_6917,N_6297,N_6492);
and U6918 (N_6918,N_6252,N_6383);
xnor U6919 (N_6919,N_6392,N_6425);
nor U6920 (N_6920,N_6036,N_6147);
and U6921 (N_6921,N_6451,N_6133);
or U6922 (N_6922,N_6041,N_6346);
and U6923 (N_6923,N_6133,N_6492);
and U6924 (N_6924,N_6430,N_6225);
nor U6925 (N_6925,N_6248,N_6195);
and U6926 (N_6926,N_6014,N_6297);
or U6927 (N_6927,N_6444,N_6353);
xor U6928 (N_6928,N_6390,N_6294);
and U6929 (N_6929,N_6050,N_6236);
or U6930 (N_6930,N_6323,N_6196);
nand U6931 (N_6931,N_6124,N_6294);
nor U6932 (N_6932,N_6478,N_6451);
and U6933 (N_6933,N_6059,N_6309);
nand U6934 (N_6934,N_6074,N_6095);
nand U6935 (N_6935,N_6076,N_6360);
nor U6936 (N_6936,N_6384,N_6105);
or U6937 (N_6937,N_6076,N_6393);
and U6938 (N_6938,N_6011,N_6095);
and U6939 (N_6939,N_6415,N_6313);
nand U6940 (N_6940,N_6255,N_6293);
or U6941 (N_6941,N_6022,N_6439);
xor U6942 (N_6942,N_6407,N_6166);
nand U6943 (N_6943,N_6012,N_6375);
nand U6944 (N_6944,N_6410,N_6337);
xnor U6945 (N_6945,N_6108,N_6124);
and U6946 (N_6946,N_6104,N_6089);
or U6947 (N_6947,N_6472,N_6044);
nand U6948 (N_6948,N_6012,N_6191);
nor U6949 (N_6949,N_6012,N_6355);
or U6950 (N_6950,N_6209,N_6453);
or U6951 (N_6951,N_6271,N_6070);
nand U6952 (N_6952,N_6468,N_6067);
nor U6953 (N_6953,N_6109,N_6378);
nand U6954 (N_6954,N_6419,N_6464);
and U6955 (N_6955,N_6228,N_6318);
nor U6956 (N_6956,N_6479,N_6344);
nor U6957 (N_6957,N_6474,N_6244);
and U6958 (N_6958,N_6120,N_6103);
and U6959 (N_6959,N_6407,N_6148);
nor U6960 (N_6960,N_6301,N_6120);
nor U6961 (N_6961,N_6059,N_6404);
and U6962 (N_6962,N_6184,N_6032);
nor U6963 (N_6963,N_6110,N_6007);
or U6964 (N_6964,N_6275,N_6235);
or U6965 (N_6965,N_6038,N_6182);
nand U6966 (N_6966,N_6082,N_6375);
xor U6967 (N_6967,N_6139,N_6039);
nor U6968 (N_6968,N_6018,N_6433);
nor U6969 (N_6969,N_6276,N_6345);
nand U6970 (N_6970,N_6032,N_6130);
nor U6971 (N_6971,N_6380,N_6144);
nor U6972 (N_6972,N_6010,N_6228);
nand U6973 (N_6973,N_6107,N_6223);
nor U6974 (N_6974,N_6217,N_6453);
nand U6975 (N_6975,N_6312,N_6302);
nor U6976 (N_6976,N_6028,N_6111);
and U6977 (N_6977,N_6008,N_6378);
nor U6978 (N_6978,N_6229,N_6110);
or U6979 (N_6979,N_6499,N_6498);
and U6980 (N_6980,N_6455,N_6381);
xnor U6981 (N_6981,N_6442,N_6208);
nand U6982 (N_6982,N_6348,N_6424);
and U6983 (N_6983,N_6051,N_6427);
nor U6984 (N_6984,N_6267,N_6416);
and U6985 (N_6985,N_6401,N_6020);
and U6986 (N_6986,N_6132,N_6480);
and U6987 (N_6987,N_6384,N_6053);
or U6988 (N_6988,N_6426,N_6165);
nor U6989 (N_6989,N_6286,N_6305);
and U6990 (N_6990,N_6446,N_6077);
and U6991 (N_6991,N_6183,N_6394);
or U6992 (N_6992,N_6115,N_6197);
or U6993 (N_6993,N_6379,N_6157);
xor U6994 (N_6994,N_6378,N_6020);
nand U6995 (N_6995,N_6363,N_6178);
nor U6996 (N_6996,N_6211,N_6350);
xor U6997 (N_6997,N_6094,N_6148);
or U6998 (N_6998,N_6025,N_6135);
or U6999 (N_6999,N_6322,N_6345);
and U7000 (N_7000,N_6934,N_6910);
nor U7001 (N_7001,N_6595,N_6665);
nor U7002 (N_7002,N_6800,N_6796);
nand U7003 (N_7003,N_6885,N_6827);
xor U7004 (N_7004,N_6502,N_6893);
or U7005 (N_7005,N_6658,N_6830);
or U7006 (N_7006,N_6767,N_6669);
and U7007 (N_7007,N_6702,N_6552);
xnor U7008 (N_7008,N_6585,N_6906);
or U7009 (N_7009,N_6788,N_6829);
nor U7010 (N_7010,N_6613,N_6543);
xnor U7011 (N_7011,N_6940,N_6873);
and U7012 (N_7012,N_6807,N_6919);
and U7013 (N_7013,N_6510,N_6735);
xnor U7014 (N_7014,N_6652,N_6857);
nor U7015 (N_7015,N_6986,N_6842);
or U7016 (N_7016,N_6773,N_6549);
nor U7017 (N_7017,N_6805,N_6538);
or U7018 (N_7018,N_6603,N_6594);
and U7019 (N_7019,N_6834,N_6911);
or U7020 (N_7020,N_6928,N_6582);
and U7021 (N_7021,N_6943,N_6682);
and U7022 (N_7022,N_6612,N_6650);
or U7023 (N_7023,N_6960,N_6721);
nor U7024 (N_7024,N_6540,N_6964);
or U7025 (N_7025,N_6792,N_6671);
or U7026 (N_7026,N_6741,N_6775);
nor U7027 (N_7027,N_6769,N_6719);
nor U7028 (N_7028,N_6664,N_6624);
nand U7029 (N_7029,N_6533,N_6812);
nand U7030 (N_7030,N_6779,N_6674);
and U7031 (N_7031,N_6746,N_6634);
nand U7032 (N_7032,N_6705,N_6630);
nand U7033 (N_7033,N_6751,N_6899);
and U7034 (N_7034,N_6967,N_6615);
and U7035 (N_7035,N_6713,N_6924);
or U7036 (N_7036,N_6505,N_6852);
xor U7037 (N_7037,N_6878,N_6791);
and U7038 (N_7038,N_6628,N_6635);
nand U7039 (N_7039,N_6514,N_6680);
nor U7040 (N_7040,N_6740,N_6776);
xnor U7041 (N_7041,N_6806,N_6987);
nor U7042 (N_7042,N_6872,N_6737);
nand U7043 (N_7043,N_6564,N_6932);
and U7044 (N_7044,N_6927,N_6575);
or U7045 (N_7045,N_6882,N_6606);
nand U7046 (N_7046,N_6780,N_6536);
nor U7047 (N_7047,N_6747,N_6637);
and U7048 (N_7048,N_6766,N_6983);
and U7049 (N_7049,N_6617,N_6811);
nand U7050 (N_7050,N_6693,N_6743);
or U7051 (N_7051,N_6631,N_6869);
xor U7052 (N_7052,N_6826,N_6849);
and U7053 (N_7053,N_6823,N_6557);
nor U7054 (N_7054,N_6600,N_6633);
nand U7055 (N_7055,N_6706,N_6623);
nor U7056 (N_7056,N_6565,N_6627);
nor U7057 (N_7057,N_6678,N_6738);
xnor U7058 (N_7058,N_6709,N_6944);
and U7059 (N_7059,N_6941,N_6534);
or U7060 (N_7060,N_6523,N_6781);
or U7061 (N_7061,N_6537,N_6856);
xor U7062 (N_7062,N_6722,N_6607);
nor U7063 (N_7063,N_6880,N_6618);
xor U7064 (N_7064,N_6808,N_6690);
nor U7065 (N_7065,N_6714,N_6556);
or U7066 (N_7066,N_6889,N_6995);
or U7067 (N_7067,N_6949,N_6951);
and U7068 (N_7068,N_6904,N_6670);
nand U7069 (N_7069,N_6844,N_6982);
nand U7070 (N_7070,N_6660,N_6578);
or U7071 (N_7071,N_6922,N_6599);
xor U7072 (N_7072,N_6583,N_6527);
nor U7073 (N_7073,N_6590,N_6587);
and U7074 (N_7074,N_6589,N_6711);
or U7075 (N_7075,N_6994,N_6501);
and U7076 (N_7076,N_6626,N_6588);
nand U7077 (N_7077,N_6659,N_6621);
xnor U7078 (N_7078,N_6522,N_6655);
or U7079 (N_7079,N_6916,N_6636);
nor U7080 (N_7080,N_6526,N_6610);
xnor U7081 (N_7081,N_6959,N_6981);
xnor U7082 (N_7082,N_6803,N_6619);
xor U7083 (N_7083,N_6917,N_6864);
nand U7084 (N_7084,N_6815,N_6768);
and U7085 (N_7085,N_6684,N_6931);
and U7086 (N_7086,N_6831,N_6528);
xnor U7087 (N_7087,N_6957,N_6611);
or U7088 (N_7088,N_6962,N_6760);
nand U7089 (N_7089,N_6790,N_6687);
and U7090 (N_7090,N_6953,N_6572);
nor U7091 (N_7091,N_6997,N_6896);
nand U7092 (N_7092,N_6942,N_6666);
and U7093 (N_7093,N_6581,N_6672);
and U7094 (N_7094,N_6989,N_6677);
xnor U7095 (N_7095,N_6914,N_6545);
nor U7096 (N_7096,N_6716,N_6692);
nand U7097 (N_7097,N_6563,N_6854);
and U7098 (N_7098,N_6833,N_6836);
nand U7099 (N_7099,N_6755,N_6947);
or U7100 (N_7100,N_6511,N_6647);
nand U7101 (N_7101,N_6886,N_6728);
and U7102 (N_7102,N_6723,N_6784);
and U7103 (N_7103,N_6871,N_6879);
nand U7104 (N_7104,N_6912,N_6843);
nor U7105 (N_7105,N_6697,N_6846);
nor U7106 (N_7106,N_6966,N_6688);
and U7107 (N_7107,N_6888,N_6818);
nor U7108 (N_7108,N_6535,N_6555);
nor U7109 (N_7109,N_6971,N_6657);
xnor U7110 (N_7110,N_6504,N_6945);
or U7111 (N_7111,N_6601,N_6804);
and U7112 (N_7112,N_6980,N_6883);
nor U7113 (N_7113,N_6956,N_6898);
nor U7114 (N_7114,N_6785,N_6976);
nand U7115 (N_7115,N_6681,N_6820);
and U7116 (N_7116,N_6707,N_6759);
nor U7117 (N_7117,N_6783,N_6978);
xnor U7118 (N_7118,N_6559,N_6547);
nor U7119 (N_7119,N_6999,N_6965);
nand U7120 (N_7120,N_6734,N_6661);
nor U7121 (N_7121,N_6770,N_6763);
nand U7122 (N_7122,N_6905,N_6866);
or U7123 (N_7123,N_6524,N_6546);
and U7124 (N_7124,N_6689,N_6969);
nor U7125 (N_7125,N_6616,N_6525);
or U7126 (N_7126,N_6608,N_6638);
nand U7127 (N_7127,N_6518,N_6668);
or U7128 (N_7128,N_6758,N_6925);
nor U7129 (N_7129,N_6541,N_6908);
and U7130 (N_7130,N_6907,N_6691);
nor U7131 (N_7131,N_6570,N_6667);
or U7132 (N_7132,N_6900,N_6991);
and U7133 (N_7133,N_6596,N_6732);
and U7134 (N_7134,N_6929,N_6996);
or U7135 (N_7135,N_6649,N_6926);
and U7136 (N_7136,N_6673,N_6712);
and U7137 (N_7137,N_6903,N_6729);
nand U7138 (N_7138,N_6993,N_6998);
or U7139 (N_7139,N_6500,N_6662);
xor U7140 (N_7140,N_6742,N_6822);
and U7141 (N_7141,N_6895,N_6860);
nor U7142 (N_7142,N_6726,N_6724);
nand U7143 (N_7143,N_6985,N_6816);
xor U7144 (N_7144,N_6569,N_6855);
and U7145 (N_7145,N_6554,N_6739);
or U7146 (N_7146,N_6890,N_6937);
nand U7147 (N_7147,N_6909,N_6946);
and U7148 (N_7148,N_6863,N_6507);
xor U7149 (N_7149,N_6799,N_6850);
or U7150 (N_7150,N_6861,N_6977);
nor U7151 (N_7151,N_6694,N_6774);
or U7152 (N_7152,N_6891,N_6913);
and U7153 (N_7153,N_6961,N_6837);
and U7154 (N_7154,N_6625,N_6643);
nor U7155 (N_7155,N_6529,N_6935);
or U7156 (N_7156,N_6853,N_6897);
and U7157 (N_7157,N_6765,N_6756);
xor U7158 (N_7158,N_6579,N_6530);
nor U7159 (N_7159,N_6506,N_6952);
and U7160 (N_7160,N_6571,N_6519);
nor U7161 (N_7161,N_6839,N_6787);
or U7162 (N_7162,N_6870,N_6715);
nor U7163 (N_7163,N_6503,N_6851);
or U7164 (N_7164,N_6686,N_6512);
and U7165 (N_7165,N_6620,N_6685);
xnor U7166 (N_7166,N_6642,N_6761);
and U7167 (N_7167,N_6797,N_6824);
and U7168 (N_7168,N_6972,N_6553);
nor U7169 (N_7169,N_6639,N_6605);
nor U7170 (N_7170,N_6876,N_6884);
and U7171 (N_7171,N_6520,N_6574);
and U7172 (N_7172,N_6825,N_6532);
and U7173 (N_7173,N_6892,N_6558);
nand U7174 (N_7174,N_6704,N_6641);
or U7175 (N_7175,N_6561,N_6745);
nor U7176 (N_7176,N_6592,N_6874);
nor U7177 (N_7177,N_6531,N_6591);
and U7178 (N_7178,N_6580,N_6542);
and U7179 (N_7179,N_6764,N_6720);
nor U7180 (N_7180,N_6923,N_6699);
and U7181 (N_7181,N_6567,N_6789);
and U7182 (N_7182,N_6614,N_6819);
nand U7183 (N_7183,N_6809,N_6835);
xnor U7184 (N_7184,N_6752,N_6508);
nor U7185 (N_7185,N_6821,N_6597);
nor U7186 (N_7186,N_6696,N_6566);
nor U7187 (N_7187,N_6539,N_6648);
or U7188 (N_7188,N_6653,N_6921);
or U7189 (N_7189,N_6663,N_6782);
xor U7190 (N_7190,N_6598,N_6901);
and U7191 (N_7191,N_6798,N_6845);
and U7192 (N_7192,N_6609,N_6568);
or U7193 (N_7193,N_6701,N_6710);
or U7194 (N_7194,N_6725,N_6772);
nand U7195 (N_7195,N_6560,N_6700);
nor U7196 (N_7196,N_6936,N_6676);
nand U7197 (N_7197,N_6984,N_6840);
xor U7198 (N_7198,N_6604,N_6915);
and U7199 (N_7199,N_6974,N_6675);
and U7200 (N_7200,N_6794,N_6573);
xnor U7201 (N_7201,N_6736,N_6813);
nand U7202 (N_7202,N_6562,N_6733);
nor U7203 (N_7203,N_6646,N_6730);
or U7204 (N_7204,N_6717,N_6754);
nand U7205 (N_7205,N_6778,N_6881);
and U7206 (N_7206,N_6753,N_6862);
xnor U7207 (N_7207,N_6838,N_6990);
and U7208 (N_7208,N_6644,N_6795);
xor U7209 (N_7209,N_6801,N_6859);
nor U7210 (N_7210,N_6586,N_6938);
and U7211 (N_7211,N_6731,N_6515);
or U7212 (N_7212,N_6877,N_6920);
nor U7213 (N_7213,N_6679,N_6656);
and U7214 (N_7214,N_6894,N_6875);
and U7215 (N_7215,N_6577,N_6548);
nand U7216 (N_7216,N_6576,N_6748);
or U7217 (N_7217,N_6744,N_6973);
nand U7218 (N_7218,N_6516,N_6550);
or U7219 (N_7219,N_6654,N_6698);
or U7220 (N_7220,N_6930,N_6727);
nand U7221 (N_7221,N_6970,N_6867);
and U7222 (N_7222,N_6793,N_6988);
nand U7223 (N_7223,N_6683,N_6513);
and U7224 (N_7224,N_6887,N_6718);
and U7225 (N_7225,N_6521,N_6629);
and U7226 (N_7226,N_6848,N_6954);
xor U7227 (N_7227,N_6975,N_6828);
nand U7228 (N_7228,N_6645,N_6749);
nand U7229 (N_7229,N_6865,N_6777);
nand U7230 (N_7230,N_6802,N_6979);
and U7231 (N_7231,N_6602,N_6858);
or U7232 (N_7232,N_6786,N_6708);
nand U7233 (N_7233,N_6517,N_6832);
nand U7234 (N_7234,N_6593,N_6814);
nor U7235 (N_7235,N_6918,N_6817);
and U7236 (N_7236,N_6544,N_6771);
and U7237 (N_7237,N_6868,N_6622);
and U7238 (N_7238,N_6902,N_6968);
nor U7239 (N_7239,N_6651,N_6757);
or U7240 (N_7240,N_6810,N_6703);
nand U7241 (N_7241,N_6632,N_6584);
nand U7242 (N_7242,N_6939,N_6847);
and U7243 (N_7243,N_6992,N_6948);
xnor U7244 (N_7244,N_6841,N_6640);
or U7245 (N_7245,N_6509,N_6762);
or U7246 (N_7246,N_6955,N_6963);
or U7247 (N_7247,N_6750,N_6695);
or U7248 (N_7248,N_6958,N_6933);
and U7249 (N_7249,N_6950,N_6551);
and U7250 (N_7250,N_6912,N_6617);
nand U7251 (N_7251,N_6886,N_6560);
or U7252 (N_7252,N_6730,N_6757);
nand U7253 (N_7253,N_6767,N_6586);
or U7254 (N_7254,N_6885,N_6864);
nor U7255 (N_7255,N_6623,N_6799);
nand U7256 (N_7256,N_6788,N_6978);
and U7257 (N_7257,N_6620,N_6961);
nand U7258 (N_7258,N_6705,N_6957);
and U7259 (N_7259,N_6939,N_6702);
and U7260 (N_7260,N_6942,N_6675);
nand U7261 (N_7261,N_6904,N_6753);
nand U7262 (N_7262,N_6577,N_6621);
nor U7263 (N_7263,N_6555,N_6701);
and U7264 (N_7264,N_6549,N_6954);
nand U7265 (N_7265,N_6764,N_6762);
nor U7266 (N_7266,N_6872,N_6962);
or U7267 (N_7267,N_6788,N_6750);
nor U7268 (N_7268,N_6913,N_6935);
nand U7269 (N_7269,N_6900,N_6980);
and U7270 (N_7270,N_6556,N_6817);
or U7271 (N_7271,N_6807,N_6603);
nand U7272 (N_7272,N_6957,N_6542);
nand U7273 (N_7273,N_6801,N_6739);
nor U7274 (N_7274,N_6836,N_6589);
or U7275 (N_7275,N_6872,N_6881);
nor U7276 (N_7276,N_6657,N_6771);
nand U7277 (N_7277,N_6927,N_6871);
or U7278 (N_7278,N_6526,N_6605);
or U7279 (N_7279,N_6729,N_6848);
nand U7280 (N_7280,N_6917,N_6985);
or U7281 (N_7281,N_6784,N_6686);
nor U7282 (N_7282,N_6727,N_6622);
xor U7283 (N_7283,N_6578,N_6506);
nor U7284 (N_7284,N_6960,N_6686);
nand U7285 (N_7285,N_6742,N_6727);
or U7286 (N_7286,N_6985,N_6870);
nand U7287 (N_7287,N_6845,N_6683);
nor U7288 (N_7288,N_6932,N_6744);
or U7289 (N_7289,N_6895,N_6940);
and U7290 (N_7290,N_6871,N_6706);
nor U7291 (N_7291,N_6664,N_6958);
and U7292 (N_7292,N_6694,N_6510);
xnor U7293 (N_7293,N_6800,N_6864);
nor U7294 (N_7294,N_6860,N_6891);
or U7295 (N_7295,N_6501,N_6772);
and U7296 (N_7296,N_6665,N_6995);
or U7297 (N_7297,N_6832,N_6546);
or U7298 (N_7298,N_6822,N_6973);
and U7299 (N_7299,N_6589,N_6692);
and U7300 (N_7300,N_6595,N_6505);
or U7301 (N_7301,N_6606,N_6506);
nand U7302 (N_7302,N_6637,N_6604);
and U7303 (N_7303,N_6976,N_6565);
and U7304 (N_7304,N_6528,N_6519);
or U7305 (N_7305,N_6901,N_6936);
or U7306 (N_7306,N_6802,N_6852);
or U7307 (N_7307,N_6578,N_6744);
nand U7308 (N_7308,N_6574,N_6903);
nand U7309 (N_7309,N_6745,N_6589);
nand U7310 (N_7310,N_6963,N_6713);
nor U7311 (N_7311,N_6640,N_6751);
or U7312 (N_7312,N_6941,N_6980);
or U7313 (N_7313,N_6624,N_6892);
and U7314 (N_7314,N_6715,N_6856);
and U7315 (N_7315,N_6758,N_6842);
and U7316 (N_7316,N_6654,N_6541);
xnor U7317 (N_7317,N_6952,N_6837);
and U7318 (N_7318,N_6567,N_6607);
and U7319 (N_7319,N_6881,N_6756);
and U7320 (N_7320,N_6884,N_6744);
or U7321 (N_7321,N_6970,N_6648);
xnor U7322 (N_7322,N_6543,N_6969);
and U7323 (N_7323,N_6584,N_6533);
xnor U7324 (N_7324,N_6631,N_6870);
or U7325 (N_7325,N_6860,N_6731);
and U7326 (N_7326,N_6553,N_6742);
and U7327 (N_7327,N_6570,N_6548);
or U7328 (N_7328,N_6994,N_6641);
nor U7329 (N_7329,N_6508,N_6571);
nand U7330 (N_7330,N_6943,N_6869);
nor U7331 (N_7331,N_6604,N_6652);
or U7332 (N_7332,N_6988,N_6547);
xnor U7333 (N_7333,N_6815,N_6742);
nand U7334 (N_7334,N_6521,N_6805);
and U7335 (N_7335,N_6593,N_6668);
nor U7336 (N_7336,N_6844,N_6651);
and U7337 (N_7337,N_6796,N_6905);
or U7338 (N_7338,N_6803,N_6953);
nand U7339 (N_7339,N_6707,N_6594);
nand U7340 (N_7340,N_6809,N_6871);
nor U7341 (N_7341,N_6835,N_6855);
or U7342 (N_7342,N_6927,N_6793);
nor U7343 (N_7343,N_6924,N_6925);
nor U7344 (N_7344,N_6836,N_6754);
nand U7345 (N_7345,N_6639,N_6835);
nand U7346 (N_7346,N_6585,N_6820);
or U7347 (N_7347,N_6752,N_6958);
nor U7348 (N_7348,N_6915,N_6646);
or U7349 (N_7349,N_6526,N_6545);
and U7350 (N_7350,N_6831,N_6572);
or U7351 (N_7351,N_6855,N_6925);
xor U7352 (N_7352,N_6986,N_6551);
nor U7353 (N_7353,N_6636,N_6678);
or U7354 (N_7354,N_6642,N_6844);
nor U7355 (N_7355,N_6947,N_6859);
or U7356 (N_7356,N_6638,N_6530);
nor U7357 (N_7357,N_6931,N_6633);
or U7358 (N_7358,N_6838,N_6758);
or U7359 (N_7359,N_6742,N_6944);
xor U7360 (N_7360,N_6651,N_6542);
nand U7361 (N_7361,N_6577,N_6897);
and U7362 (N_7362,N_6938,N_6969);
nor U7363 (N_7363,N_6668,N_6887);
nor U7364 (N_7364,N_6972,N_6708);
and U7365 (N_7365,N_6623,N_6755);
and U7366 (N_7366,N_6583,N_6737);
nor U7367 (N_7367,N_6811,N_6608);
or U7368 (N_7368,N_6766,N_6619);
or U7369 (N_7369,N_6848,N_6873);
xor U7370 (N_7370,N_6589,N_6538);
nor U7371 (N_7371,N_6954,N_6528);
or U7372 (N_7372,N_6613,N_6558);
xor U7373 (N_7373,N_6832,N_6863);
nand U7374 (N_7374,N_6618,N_6602);
nand U7375 (N_7375,N_6715,N_6910);
and U7376 (N_7376,N_6856,N_6605);
nor U7377 (N_7377,N_6611,N_6821);
nor U7378 (N_7378,N_6979,N_6815);
and U7379 (N_7379,N_6790,N_6604);
and U7380 (N_7380,N_6836,N_6591);
and U7381 (N_7381,N_6823,N_6874);
or U7382 (N_7382,N_6649,N_6592);
or U7383 (N_7383,N_6694,N_6652);
nand U7384 (N_7384,N_6707,N_6750);
nor U7385 (N_7385,N_6810,N_6786);
nand U7386 (N_7386,N_6829,N_6521);
nor U7387 (N_7387,N_6643,N_6615);
or U7388 (N_7388,N_6553,N_6783);
and U7389 (N_7389,N_6873,N_6800);
and U7390 (N_7390,N_6890,N_6866);
and U7391 (N_7391,N_6630,N_6914);
xnor U7392 (N_7392,N_6744,N_6849);
or U7393 (N_7393,N_6678,N_6671);
or U7394 (N_7394,N_6997,N_6764);
xnor U7395 (N_7395,N_6548,N_6868);
nor U7396 (N_7396,N_6715,N_6792);
nand U7397 (N_7397,N_6552,N_6949);
and U7398 (N_7398,N_6559,N_6896);
nor U7399 (N_7399,N_6759,N_6703);
and U7400 (N_7400,N_6832,N_6926);
nand U7401 (N_7401,N_6526,N_6951);
nand U7402 (N_7402,N_6692,N_6843);
xnor U7403 (N_7403,N_6559,N_6730);
or U7404 (N_7404,N_6630,N_6739);
xnor U7405 (N_7405,N_6942,N_6653);
nand U7406 (N_7406,N_6954,N_6554);
or U7407 (N_7407,N_6723,N_6513);
or U7408 (N_7408,N_6661,N_6884);
xnor U7409 (N_7409,N_6788,N_6758);
and U7410 (N_7410,N_6907,N_6628);
nand U7411 (N_7411,N_6923,N_6679);
and U7412 (N_7412,N_6551,N_6603);
or U7413 (N_7413,N_6786,N_6724);
nor U7414 (N_7414,N_6582,N_6979);
nor U7415 (N_7415,N_6557,N_6993);
and U7416 (N_7416,N_6633,N_6729);
nor U7417 (N_7417,N_6926,N_6747);
nand U7418 (N_7418,N_6788,N_6859);
nor U7419 (N_7419,N_6617,N_6924);
nand U7420 (N_7420,N_6645,N_6686);
nor U7421 (N_7421,N_6776,N_6877);
nand U7422 (N_7422,N_6851,N_6985);
xor U7423 (N_7423,N_6797,N_6668);
nor U7424 (N_7424,N_6748,N_6638);
nor U7425 (N_7425,N_6999,N_6551);
nand U7426 (N_7426,N_6528,N_6969);
nor U7427 (N_7427,N_6957,N_6968);
or U7428 (N_7428,N_6525,N_6967);
nand U7429 (N_7429,N_6952,N_6935);
nor U7430 (N_7430,N_6563,N_6805);
nand U7431 (N_7431,N_6542,N_6635);
and U7432 (N_7432,N_6659,N_6866);
or U7433 (N_7433,N_6961,N_6944);
nor U7434 (N_7434,N_6733,N_6619);
or U7435 (N_7435,N_6725,N_6829);
and U7436 (N_7436,N_6582,N_6657);
nor U7437 (N_7437,N_6859,N_6677);
nor U7438 (N_7438,N_6937,N_6744);
nand U7439 (N_7439,N_6633,N_6901);
nor U7440 (N_7440,N_6529,N_6572);
nand U7441 (N_7441,N_6653,N_6986);
nor U7442 (N_7442,N_6889,N_6708);
nor U7443 (N_7443,N_6798,N_6644);
xnor U7444 (N_7444,N_6850,N_6809);
nor U7445 (N_7445,N_6983,N_6749);
or U7446 (N_7446,N_6993,N_6716);
and U7447 (N_7447,N_6892,N_6840);
and U7448 (N_7448,N_6966,N_6793);
nand U7449 (N_7449,N_6925,N_6668);
or U7450 (N_7450,N_6716,N_6543);
and U7451 (N_7451,N_6755,N_6576);
or U7452 (N_7452,N_6835,N_6783);
or U7453 (N_7453,N_6768,N_6998);
and U7454 (N_7454,N_6719,N_6908);
and U7455 (N_7455,N_6969,N_6822);
nor U7456 (N_7456,N_6912,N_6939);
or U7457 (N_7457,N_6960,N_6572);
or U7458 (N_7458,N_6673,N_6856);
and U7459 (N_7459,N_6942,N_6618);
nand U7460 (N_7460,N_6646,N_6799);
and U7461 (N_7461,N_6755,N_6831);
nand U7462 (N_7462,N_6743,N_6505);
xnor U7463 (N_7463,N_6930,N_6858);
or U7464 (N_7464,N_6539,N_6662);
and U7465 (N_7465,N_6878,N_6871);
nor U7466 (N_7466,N_6900,N_6982);
and U7467 (N_7467,N_6563,N_6686);
nand U7468 (N_7468,N_6699,N_6884);
nand U7469 (N_7469,N_6859,N_6684);
xnor U7470 (N_7470,N_6578,N_6697);
or U7471 (N_7471,N_6911,N_6614);
nor U7472 (N_7472,N_6701,N_6876);
nor U7473 (N_7473,N_6552,N_6781);
or U7474 (N_7474,N_6872,N_6649);
and U7475 (N_7475,N_6834,N_6824);
nor U7476 (N_7476,N_6679,N_6991);
and U7477 (N_7477,N_6753,N_6919);
or U7478 (N_7478,N_6558,N_6753);
nor U7479 (N_7479,N_6801,N_6964);
and U7480 (N_7480,N_6823,N_6793);
and U7481 (N_7481,N_6783,N_6559);
nand U7482 (N_7482,N_6996,N_6721);
and U7483 (N_7483,N_6952,N_6944);
nand U7484 (N_7484,N_6709,N_6910);
or U7485 (N_7485,N_6793,N_6637);
nor U7486 (N_7486,N_6731,N_6759);
and U7487 (N_7487,N_6560,N_6608);
or U7488 (N_7488,N_6632,N_6682);
and U7489 (N_7489,N_6564,N_6588);
and U7490 (N_7490,N_6544,N_6829);
or U7491 (N_7491,N_6667,N_6942);
nor U7492 (N_7492,N_6865,N_6932);
nor U7493 (N_7493,N_6548,N_6757);
nor U7494 (N_7494,N_6860,N_6649);
and U7495 (N_7495,N_6999,N_6832);
nand U7496 (N_7496,N_6647,N_6532);
nor U7497 (N_7497,N_6853,N_6950);
or U7498 (N_7498,N_6524,N_6565);
xnor U7499 (N_7499,N_6690,N_6742);
or U7500 (N_7500,N_7150,N_7110);
and U7501 (N_7501,N_7214,N_7469);
nand U7502 (N_7502,N_7377,N_7248);
or U7503 (N_7503,N_7168,N_7277);
nor U7504 (N_7504,N_7448,N_7157);
or U7505 (N_7505,N_7333,N_7477);
and U7506 (N_7506,N_7271,N_7149);
or U7507 (N_7507,N_7370,N_7140);
nand U7508 (N_7508,N_7031,N_7159);
nand U7509 (N_7509,N_7101,N_7267);
xnor U7510 (N_7510,N_7073,N_7083);
or U7511 (N_7511,N_7230,N_7053);
nor U7512 (N_7512,N_7126,N_7480);
or U7513 (N_7513,N_7385,N_7086);
nor U7514 (N_7514,N_7438,N_7146);
and U7515 (N_7515,N_7381,N_7300);
or U7516 (N_7516,N_7362,N_7250);
and U7517 (N_7517,N_7346,N_7118);
xnor U7518 (N_7518,N_7051,N_7495);
and U7519 (N_7519,N_7039,N_7494);
nand U7520 (N_7520,N_7177,N_7044);
nor U7521 (N_7521,N_7211,N_7336);
and U7522 (N_7522,N_7270,N_7142);
nand U7523 (N_7523,N_7202,N_7123);
or U7524 (N_7524,N_7069,N_7249);
nor U7525 (N_7525,N_7190,N_7310);
nand U7526 (N_7526,N_7196,N_7290);
nor U7527 (N_7527,N_7392,N_7225);
xnor U7528 (N_7528,N_7371,N_7025);
nand U7529 (N_7529,N_7062,N_7203);
xor U7530 (N_7530,N_7332,N_7032);
nand U7531 (N_7531,N_7339,N_7048);
nand U7532 (N_7532,N_7008,N_7218);
or U7533 (N_7533,N_7487,N_7374);
nand U7534 (N_7534,N_7012,N_7348);
and U7535 (N_7535,N_7158,N_7263);
nand U7536 (N_7536,N_7397,N_7176);
and U7537 (N_7537,N_7119,N_7446);
nor U7538 (N_7538,N_7458,N_7052);
nand U7539 (N_7539,N_7360,N_7317);
nand U7540 (N_7540,N_7319,N_7496);
or U7541 (N_7541,N_7375,N_7217);
or U7542 (N_7542,N_7476,N_7365);
and U7543 (N_7543,N_7350,N_7246);
or U7544 (N_7544,N_7213,N_7103);
nor U7545 (N_7545,N_7296,N_7399);
and U7546 (N_7546,N_7005,N_7037);
and U7547 (N_7547,N_7147,N_7148);
nor U7548 (N_7548,N_7413,N_7390);
and U7549 (N_7549,N_7046,N_7467);
and U7550 (N_7550,N_7459,N_7231);
nor U7551 (N_7551,N_7207,N_7324);
and U7552 (N_7552,N_7015,N_7412);
nor U7553 (N_7553,N_7279,N_7283);
nor U7554 (N_7554,N_7445,N_7185);
nor U7555 (N_7555,N_7182,N_7482);
nor U7556 (N_7556,N_7474,N_7255);
xor U7557 (N_7557,N_7261,N_7434);
xor U7558 (N_7558,N_7206,N_7063);
nand U7559 (N_7559,N_7120,N_7268);
nand U7560 (N_7560,N_7491,N_7338);
nor U7561 (N_7561,N_7368,N_7428);
or U7562 (N_7562,N_7030,N_7334);
nand U7563 (N_7563,N_7287,N_7414);
nor U7564 (N_7564,N_7096,N_7275);
or U7565 (N_7565,N_7179,N_7163);
and U7566 (N_7566,N_7306,N_7386);
and U7567 (N_7567,N_7369,N_7138);
and U7568 (N_7568,N_7026,N_7498);
nor U7569 (N_7569,N_7416,N_7393);
or U7570 (N_7570,N_7418,N_7252);
nand U7571 (N_7571,N_7235,N_7254);
xor U7572 (N_7572,N_7253,N_7098);
and U7573 (N_7573,N_7167,N_7401);
or U7574 (N_7574,N_7180,N_7437);
nor U7575 (N_7575,N_7162,N_7092);
or U7576 (N_7576,N_7499,N_7439);
xor U7577 (N_7577,N_7132,N_7361);
nor U7578 (N_7578,N_7088,N_7014);
nor U7579 (N_7579,N_7197,N_7041);
xnor U7580 (N_7580,N_7427,N_7233);
and U7581 (N_7581,N_7156,N_7049);
or U7582 (N_7582,N_7372,N_7405);
or U7583 (N_7583,N_7085,N_7077);
or U7584 (N_7584,N_7042,N_7109);
nand U7585 (N_7585,N_7050,N_7059);
and U7586 (N_7586,N_7121,N_7061);
nor U7587 (N_7587,N_7170,N_7128);
or U7588 (N_7588,N_7466,N_7314);
nor U7589 (N_7589,N_7321,N_7341);
or U7590 (N_7590,N_7293,N_7429);
xnor U7591 (N_7591,N_7442,N_7236);
and U7592 (N_7592,N_7072,N_7492);
nor U7593 (N_7593,N_7289,N_7278);
nor U7594 (N_7594,N_7407,N_7454);
or U7595 (N_7595,N_7302,N_7355);
and U7596 (N_7596,N_7431,N_7432);
nand U7597 (N_7597,N_7464,N_7342);
xor U7598 (N_7598,N_7485,N_7097);
nor U7599 (N_7599,N_7227,N_7137);
and U7600 (N_7600,N_7286,N_7394);
or U7601 (N_7601,N_7111,N_7007);
nor U7602 (N_7602,N_7001,N_7335);
nand U7603 (N_7603,N_7018,N_7478);
nand U7604 (N_7604,N_7391,N_7175);
nand U7605 (N_7605,N_7160,N_7065);
or U7606 (N_7606,N_7345,N_7356);
nand U7607 (N_7607,N_7130,N_7328);
nor U7608 (N_7608,N_7387,N_7057);
and U7609 (N_7609,N_7316,N_7288);
and U7610 (N_7610,N_7460,N_7192);
or U7611 (N_7611,N_7272,N_7105);
nor U7612 (N_7612,N_7367,N_7090);
and U7613 (N_7613,N_7465,N_7173);
or U7614 (N_7614,N_7463,N_7004);
or U7615 (N_7615,N_7228,N_7078);
or U7616 (N_7616,N_7450,N_7043);
or U7617 (N_7617,N_7166,N_7080);
nand U7618 (N_7618,N_7280,N_7011);
or U7619 (N_7619,N_7276,N_7262);
or U7620 (N_7620,N_7234,N_7444);
nand U7621 (N_7621,N_7389,N_7481);
nand U7622 (N_7622,N_7396,N_7323);
or U7623 (N_7623,N_7074,N_7423);
and U7624 (N_7624,N_7411,N_7003);
xor U7625 (N_7625,N_7269,N_7219);
and U7626 (N_7626,N_7419,N_7484);
nand U7627 (N_7627,N_7112,N_7409);
and U7628 (N_7628,N_7127,N_7164);
nand U7629 (N_7629,N_7388,N_7285);
nor U7630 (N_7630,N_7415,N_7410);
or U7631 (N_7631,N_7304,N_7084);
nand U7632 (N_7632,N_7373,N_7452);
nand U7633 (N_7633,N_7376,N_7135);
nor U7634 (N_7634,N_7244,N_7010);
or U7635 (N_7635,N_7307,N_7479);
or U7636 (N_7636,N_7047,N_7161);
nand U7637 (N_7637,N_7295,N_7238);
or U7638 (N_7638,N_7215,N_7068);
nand U7639 (N_7639,N_7038,N_7058);
nor U7640 (N_7640,N_7151,N_7171);
nand U7641 (N_7641,N_7122,N_7184);
or U7642 (N_7642,N_7357,N_7461);
nand U7643 (N_7643,N_7404,N_7449);
nor U7644 (N_7644,N_7199,N_7406);
nor U7645 (N_7645,N_7353,N_7113);
or U7646 (N_7646,N_7091,N_7124);
nor U7647 (N_7647,N_7033,N_7089);
nor U7648 (N_7648,N_7027,N_7294);
or U7649 (N_7649,N_7311,N_7129);
nand U7650 (N_7650,N_7237,N_7241);
nor U7651 (N_7651,N_7006,N_7054);
nor U7652 (N_7652,N_7331,N_7079);
nor U7653 (N_7653,N_7106,N_7284);
nand U7654 (N_7654,N_7155,N_7395);
or U7655 (N_7655,N_7071,N_7384);
or U7656 (N_7656,N_7036,N_7318);
and U7657 (N_7657,N_7139,N_7322);
or U7658 (N_7658,N_7125,N_7327);
xnor U7659 (N_7659,N_7013,N_7240);
nand U7660 (N_7660,N_7301,N_7497);
and U7661 (N_7661,N_7028,N_7174);
xor U7662 (N_7662,N_7273,N_7108);
xnor U7663 (N_7663,N_7222,N_7299);
nor U7664 (N_7664,N_7420,N_7178);
nor U7665 (N_7665,N_7486,N_7076);
or U7666 (N_7666,N_7440,N_7475);
nand U7667 (N_7667,N_7380,N_7358);
nand U7668 (N_7668,N_7201,N_7379);
or U7669 (N_7669,N_7408,N_7344);
nand U7670 (N_7670,N_7035,N_7451);
xnor U7671 (N_7671,N_7191,N_7210);
or U7672 (N_7672,N_7455,N_7100);
nand U7673 (N_7673,N_7422,N_7169);
xor U7674 (N_7674,N_7326,N_7424);
nand U7675 (N_7675,N_7195,N_7000);
and U7676 (N_7676,N_7297,N_7021);
nor U7677 (N_7677,N_7264,N_7243);
or U7678 (N_7678,N_7141,N_7453);
nor U7679 (N_7679,N_7020,N_7183);
nand U7680 (N_7680,N_7468,N_7205);
xor U7681 (N_7681,N_7274,N_7425);
or U7682 (N_7682,N_7070,N_7343);
nor U7683 (N_7683,N_7352,N_7116);
or U7684 (N_7684,N_7320,N_7347);
nand U7685 (N_7685,N_7378,N_7009);
nor U7686 (N_7686,N_7447,N_7329);
xnor U7687 (N_7687,N_7292,N_7383);
and U7688 (N_7688,N_7117,N_7133);
nand U7689 (N_7689,N_7312,N_7060);
nand U7690 (N_7690,N_7441,N_7443);
and U7691 (N_7691,N_7456,N_7154);
and U7692 (N_7692,N_7056,N_7403);
nor U7693 (N_7693,N_7024,N_7398);
nor U7694 (N_7694,N_7212,N_7239);
and U7695 (N_7695,N_7082,N_7200);
and U7696 (N_7696,N_7066,N_7359);
xor U7697 (N_7697,N_7426,N_7349);
and U7698 (N_7698,N_7457,N_7114);
and U7699 (N_7699,N_7232,N_7220);
nand U7700 (N_7700,N_7136,N_7143);
nand U7701 (N_7701,N_7305,N_7016);
and U7702 (N_7702,N_7291,N_7019);
or U7703 (N_7703,N_7165,N_7226);
or U7704 (N_7704,N_7298,N_7189);
nor U7705 (N_7705,N_7430,N_7489);
nor U7706 (N_7706,N_7194,N_7055);
nand U7707 (N_7707,N_7187,N_7340);
nand U7708 (N_7708,N_7266,N_7483);
or U7709 (N_7709,N_7308,N_7134);
and U7710 (N_7710,N_7067,N_7313);
and U7711 (N_7711,N_7436,N_7256);
xor U7712 (N_7712,N_7221,N_7223);
xor U7713 (N_7713,N_7259,N_7198);
and U7714 (N_7714,N_7488,N_7462);
nand U7715 (N_7715,N_7099,N_7186);
xnor U7716 (N_7716,N_7265,N_7172);
nand U7717 (N_7717,N_7064,N_7022);
and U7718 (N_7718,N_7145,N_7257);
nand U7719 (N_7719,N_7382,N_7282);
nor U7720 (N_7720,N_7045,N_7017);
nor U7721 (N_7721,N_7303,N_7029);
or U7722 (N_7722,N_7040,N_7034);
and U7723 (N_7723,N_7400,N_7131);
and U7724 (N_7724,N_7081,N_7087);
or U7725 (N_7725,N_7115,N_7471);
or U7726 (N_7726,N_7258,N_7152);
and U7727 (N_7727,N_7095,N_7229);
and U7728 (N_7728,N_7104,N_7363);
nand U7729 (N_7729,N_7337,N_7075);
nand U7730 (N_7730,N_7493,N_7102);
xnor U7731 (N_7731,N_7281,N_7366);
nand U7732 (N_7732,N_7354,N_7433);
and U7733 (N_7733,N_7204,N_7153);
xor U7734 (N_7734,N_7002,N_7473);
nand U7735 (N_7735,N_7023,N_7093);
or U7736 (N_7736,N_7208,N_7245);
nor U7737 (N_7737,N_7251,N_7325);
nor U7738 (N_7738,N_7364,N_7224);
or U7739 (N_7739,N_7216,N_7315);
and U7740 (N_7740,N_7470,N_7490);
nor U7741 (N_7741,N_7209,N_7193);
nor U7742 (N_7742,N_7260,N_7417);
nor U7743 (N_7743,N_7402,N_7242);
and U7744 (N_7744,N_7107,N_7181);
nor U7745 (N_7745,N_7094,N_7330);
nor U7746 (N_7746,N_7421,N_7472);
and U7747 (N_7747,N_7435,N_7188);
and U7748 (N_7748,N_7247,N_7309);
nand U7749 (N_7749,N_7351,N_7144);
nand U7750 (N_7750,N_7221,N_7075);
or U7751 (N_7751,N_7342,N_7491);
nand U7752 (N_7752,N_7362,N_7446);
and U7753 (N_7753,N_7205,N_7354);
nor U7754 (N_7754,N_7402,N_7083);
nand U7755 (N_7755,N_7462,N_7299);
nor U7756 (N_7756,N_7297,N_7419);
nand U7757 (N_7757,N_7372,N_7193);
or U7758 (N_7758,N_7015,N_7311);
or U7759 (N_7759,N_7044,N_7497);
or U7760 (N_7760,N_7160,N_7347);
or U7761 (N_7761,N_7247,N_7036);
and U7762 (N_7762,N_7345,N_7119);
or U7763 (N_7763,N_7051,N_7292);
nand U7764 (N_7764,N_7209,N_7168);
nand U7765 (N_7765,N_7189,N_7109);
nand U7766 (N_7766,N_7093,N_7352);
nor U7767 (N_7767,N_7104,N_7149);
and U7768 (N_7768,N_7185,N_7322);
or U7769 (N_7769,N_7225,N_7491);
and U7770 (N_7770,N_7342,N_7380);
or U7771 (N_7771,N_7472,N_7001);
xor U7772 (N_7772,N_7345,N_7150);
and U7773 (N_7773,N_7435,N_7390);
nor U7774 (N_7774,N_7388,N_7443);
and U7775 (N_7775,N_7335,N_7093);
nor U7776 (N_7776,N_7200,N_7276);
or U7777 (N_7777,N_7200,N_7081);
or U7778 (N_7778,N_7489,N_7334);
nand U7779 (N_7779,N_7413,N_7067);
or U7780 (N_7780,N_7302,N_7294);
and U7781 (N_7781,N_7328,N_7058);
or U7782 (N_7782,N_7010,N_7193);
xnor U7783 (N_7783,N_7450,N_7145);
nand U7784 (N_7784,N_7169,N_7240);
nand U7785 (N_7785,N_7349,N_7286);
or U7786 (N_7786,N_7185,N_7034);
xnor U7787 (N_7787,N_7495,N_7161);
nor U7788 (N_7788,N_7139,N_7153);
or U7789 (N_7789,N_7031,N_7460);
nand U7790 (N_7790,N_7089,N_7196);
xnor U7791 (N_7791,N_7257,N_7013);
nand U7792 (N_7792,N_7418,N_7169);
nor U7793 (N_7793,N_7062,N_7414);
nor U7794 (N_7794,N_7308,N_7116);
nor U7795 (N_7795,N_7409,N_7375);
nor U7796 (N_7796,N_7225,N_7483);
nor U7797 (N_7797,N_7120,N_7469);
nand U7798 (N_7798,N_7318,N_7173);
nand U7799 (N_7799,N_7380,N_7481);
nor U7800 (N_7800,N_7431,N_7079);
nand U7801 (N_7801,N_7297,N_7313);
nor U7802 (N_7802,N_7467,N_7012);
nand U7803 (N_7803,N_7234,N_7385);
and U7804 (N_7804,N_7225,N_7208);
nand U7805 (N_7805,N_7122,N_7495);
nor U7806 (N_7806,N_7375,N_7181);
nand U7807 (N_7807,N_7162,N_7297);
or U7808 (N_7808,N_7317,N_7124);
nand U7809 (N_7809,N_7003,N_7351);
nor U7810 (N_7810,N_7420,N_7230);
or U7811 (N_7811,N_7053,N_7031);
and U7812 (N_7812,N_7226,N_7204);
nor U7813 (N_7813,N_7075,N_7015);
nor U7814 (N_7814,N_7173,N_7372);
nand U7815 (N_7815,N_7271,N_7185);
nor U7816 (N_7816,N_7026,N_7437);
or U7817 (N_7817,N_7030,N_7115);
nand U7818 (N_7818,N_7326,N_7333);
and U7819 (N_7819,N_7187,N_7325);
nand U7820 (N_7820,N_7045,N_7435);
or U7821 (N_7821,N_7376,N_7268);
nand U7822 (N_7822,N_7419,N_7196);
xnor U7823 (N_7823,N_7005,N_7043);
nor U7824 (N_7824,N_7436,N_7161);
and U7825 (N_7825,N_7167,N_7072);
nand U7826 (N_7826,N_7125,N_7091);
or U7827 (N_7827,N_7162,N_7366);
nor U7828 (N_7828,N_7241,N_7335);
xnor U7829 (N_7829,N_7358,N_7261);
xnor U7830 (N_7830,N_7071,N_7327);
or U7831 (N_7831,N_7468,N_7498);
nor U7832 (N_7832,N_7331,N_7039);
xor U7833 (N_7833,N_7138,N_7146);
or U7834 (N_7834,N_7155,N_7094);
nor U7835 (N_7835,N_7406,N_7462);
nor U7836 (N_7836,N_7034,N_7000);
nand U7837 (N_7837,N_7336,N_7341);
and U7838 (N_7838,N_7380,N_7329);
xor U7839 (N_7839,N_7181,N_7246);
and U7840 (N_7840,N_7028,N_7144);
nand U7841 (N_7841,N_7469,N_7115);
nand U7842 (N_7842,N_7126,N_7323);
nand U7843 (N_7843,N_7105,N_7474);
nor U7844 (N_7844,N_7368,N_7309);
nor U7845 (N_7845,N_7287,N_7271);
nor U7846 (N_7846,N_7113,N_7398);
or U7847 (N_7847,N_7072,N_7401);
and U7848 (N_7848,N_7446,N_7169);
or U7849 (N_7849,N_7283,N_7107);
and U7850 (N_7850,N_7499,N_7273);
or U7851 (N_7851,N_7125,N_7071);
nor U7852 (N_7852,N_7473,N_7444);
nor U7853 (N_7853,N_7267,N_7151);
and U7854 (N_7854,N_7113,N_7042);
nand U7855 (N_7855,N_7320,N_7101);
nand U7856 (N_7856,N_7185,N_7148);
or U7857 (N_7857,N_7221,N_7477);
or U7858 (N_7858,N_7110,N_7332);
nand U7859 (N_7859,N_7011,N_7406);
and U7860 (N_7860,N_7132,N_7068);
nand U7861 (N_7861,N_7025,N_7337);
or U7862 (N_7862,N_7116,N_7107);
nor U7863 (N_7863,N_7371,N_7457);
and U7864 (N_7864,N_7030,N_7090);
nand U7865 (N_7865,N_7222,N_7425);
and U7866 (N_7866,N_7371,N_7108);
nor U7867 (N_7867,N_7159,N_7222);
and U7868 (N_7868,N_7207,N_7235);
nand U7869 (N_7869,N_7138,N_7202);
and U7870 (N_7870,N_7357,N_7415);
and U7871 (N_7871,N_7396,N_7414);
or U7872 (N_7872,N_7259,N_7147);
and U7873 (N_7873,N_7255,N_7199);
xnor U7874 (N_7874,N_7089,N_7100);
nor U7875 (N_7875,N_7278,N_7035);
or U7876 (N_7876,N_7479,N_7251);
or U7877 (N_7877,N_7354,N_7464);
xnor U7878 (N_7878,N_7480,N_7018);
or U7879 (N_7879,N_7286,N_7115);
and U7880 (N_7880,N_7204,N_7417);
nor U7881 (N_7881,N_7335,N_7033);
nand U7882 (N_7882,N_7061,N_7469);
nor U7883 (N_7883,N_7336,N_7265);
or U7884 (N_7884,N_7013,N_7103);
xor U7885 (N_7885,N_7464,N_7356);
or U7886 (N_7886,N_7476,N_7370);
or U7887 (N_7887,N_7293,N_7195);
xor U7888 (N_7888,N_7199,N_7167);
or U7889 (N_7889,N_7009,N_7309);
and U7890 (N_7890,N_7183,N_7099);
or U7891 (N_7891,N_7370,N_7273);
and U7892 (N_7892,N_7342,N_7381);
and U7893 (N_7893,N_7370,N_7017);
or U7894 (N_7894,N_7268,N_7364);
nand U7895 (N_7895,N_7173,N_7078);
and U7896 (N_7896,N_7095,N_7339);
nor U7897 (N_7897,N_7422,N_7317);
or U7898 (N_7898,N_7424,N_7284);
or U7899 (N_7899,N_7479,N_7424);
and U7900 (N_7900,N_7177,N_7161);
and U7901 (N_7901,N_7240,N_7306);
and U7902 (N_7902,N_7109,N_7264);
nor U7903 (N_7903,N_7194,N_7225);
or U7904 (N_7904,N_7096,N_7427);
or U7905 (N_7905,N_7401,N_7423);
and U7906 (N_7906,N_7391,N_7117);
nor U7907 (N_7907,N_7213,N_7469);
nor U7908 (N_7908,N_7482,N_7038);
nand U7909 (N_7909,N_7122,N_7467);
and U7910 (N_7910,N_7179,N_7314);
nor U7911 (N_7911,N_7363,N_7372);
nand U7912 (N_7912,N_7496,N_7249);
nand U7913 (N_7913,N_7336,N_7494);
nand U7914 (N_7914,N_7380,N_7448);
and U7915 (N_7915,N_7108,N_7351);
nand U7916 (N_7916,N_7101,N_7031);
xnor U7917 (N_7917,N_7424,N_7446);
nor U7918 (N_7918,N_7086,N_7234);
nor U7919 (N_7919,N_7454,N_7131);
and U7920 (N_7920,N_7117,N_7227);
and U7921 (N_7921,N_7369,N_7011);
or U7922 (N_7922,N_7042,N_7470);
nor U7923 (N_7923,N_7385,N_7379);
nor U7924 (N_7924,N_7458,N_7228);
xor U7925 (N_7925,N_7406,N_7084);
and U7926 (N_7926,N_7261,N_7465);
nand U7927 (N_7927,N_7098,N_7154);
or U7928 (N_7928,N_7218,N_7027);
and U7929 (N_7929,N_7442,N_7255);
nand U7930 (N_7930,N_7329,N_7277);
and U7931 (N_7931,N_7253,N_7215);
nor U7932 (N_7932,N_7078,N_7140);
and U7933 (N_7933,N_7421,N_7440);
nand U7934 (N_7934,N_7085,N_7248);
and U7935 (N_7935,N_7098,N_7396);
nand U7936 (N_7936,N_7349,N_7174);
nor U7937 (N_7937,N_7404,N_7486);
and U7938 (N_7938,N_7117,N_7374);
xnor U7939 (N_7939,N_7099,N_7438);
and U7940 (N_7940,N_7091,N_7378);
nand U7941 (N_7941,N_7369,N_7148);
and U7942 (N_7942,N_7466,N_7209);
and U7943 (N_7943,N_7481,N_7458);
nor U7944 (N_7944,N_7007,N_7070);
and U7945 (N_7945,N_7245,N_7397);
xor U7946 (N_7946,N_7032,N_7038);
and U7947 (N_7947,N_7232,N_7383);
nand U7948 (N_7948,N_7170,N_7205);
or U7949 (N_7949,N_7200,N_7435);
nor U7950 (N_7950,N_7043,N_7099);
or U7951 (N_7951,N_7312,N_7157);
nand U7952 (N_7952,N_7102,N_7464);
or U7953 (N_7953,N_7456,N_7039);
nor U7954 (N_7954,N_7443,N_7247);
nor U7955 (N_7955,N_7018,N_7230);
xor U7956 (N_7956,N_7261,N_7075);
nor U7957 (N_7957,N_7115,N_7094);
or U7958 (N_7958,N_7230,N_7079);
xor U7959 (N_7959,N_7040,N_7333);
nand U7960 (N_7960,N_7306,N_7268);
nor U7961 (N_7961,N_7013,N_7432);
nand U7962 (N_7962,N_7496,N_7204);
or U7963 (N_7963,N_7128,N_7100);
xnor U7964 (N_7964,N_7231,N_7464);
and U7965 (N_7965,N_7260,N_7349);
xnor U7966 (N_7966,N_7443,N_7048);
nor U7967 (N_7967,N_7002,N_7377);
nand U7968 (N_7968,N_7204,N_7358);
and U7969 (N_7969,N_7312,N_7405);
and U7970 (N_7970,N_7215,N_7204);
nand U7971 (N_7971,N_7272,N_7063);
and U7972 (N_7972,N_7489,N_7434);
nor U7973 (N_7973,N_7462,N_7437);
nand U7974 (N_7974,N_7412,N_7136);
nand U7975 (N_7975,N_7280,N_7166);
nand U7976 (N_7976,N_7149,N_7259);
nand U7977 (N_7977,N_7131,N_7406);
and U7978 (N_7978,N_7336,N_7209);
nor U7979 (N_7979,N_7498,N_7198);
nand U7980 (N_7980,N_7058,N_7057);
or U7981 (N_7981,N_7193,N_7451);
nor U7982 (N_7982,N_7346,N_7232);
nand U7983 (N_7983,N_7097,N_7431);
nand U7984 (N_7984,N_7060,N_7426);
nor U7985 (N_7985,N_7173,N_7274);
and U7986 (N_7986,N_7017,N_7242);
and U7987 (N_7987,N_7217,N_7341);
nand U7988 (N_7988,N_7248,N_7499);
xor U7989 (N_7989,N_7423,N_7179);
nor U7990 (N_7990,N_7348,N_7411);
nand U7991 (N_7991,N_7130,N_7025);
or U7992 (N_7992,N_7242,N_7182);
xnor U7993 (N_7993,N_7074,N_7336);
nor U7994 (N_7994,N_7104,N_7255);
nand U7995 (N_7995,N_7130,N_7298);
nand U7996 (N_7996,N_7026,N_7448);
nand U7997 (N_7997,N_7093,N_7150);
or U7998 (N_7998,N_7340,N_7089);
nand U7999 (N_7999,N_7007,N_7033);
and U8000 (N_8000,N_7544,N_7993);
nor U8001 (N_8001,N_7634,N_7819);
nor U8002 (N_8002,N_7962,N_7813);
and U8003 (N_8003,N_7615,N_7742);
nand U8004 (N_8004,N_7638,N_7933);
and U8005 (N_8005,N_7884,N_7964);
or U8006 (N_8006,N_7881,N_7624);
nor U8007 (N_8007,N_7579,N_7764);
nor U8008 (N_8008,N_7576,N_7865);
or U8009 (N_8009,N_7805,N_7581);
or U8010 (N_8010,N_7732,N_7533);
or U8011 (N_8011,N_7722,N_7556);
nor U8012 (N_8012,N_7654,N_7888);
or U8013 (N_8013,N_7738,N_7977);
xor U8014 (N_8014,N_7734,N_7783);
and U8015 (N_8015,N_7970,N_7617);
nor U8016 (N_8016,N_7514,N_7880);
and U8017 (N_8017,N_7577,N_7875);
or U8018 (N_8018,N_7820,N_7739);
or U8019 (N_8019,N_7906,N_7768);
or U8020 (N_8020,N_7811,N_7668);
nand U8021 (N_8021,N_7748,N_7952);
nor U8022 (N_8022,N_7862,N_7703);
xor U8023 (N_8023,N_7570,N_7817);
or U8024 (N_8024,N_7803,N_7737);
or U8025 (N_8025,N_7950,N_7765);
nor U8026 (N_8026,N_7625,N_7678);
and U8027 (N_8027,N_7789,N_7958);
or U8028 (N_8028,N_7542,N_7599);
and U8029 (N_8029,N_7727,N_7616);
or U8030 (N_8030,N_7868,N_7893);
nor U8031 (N_8031,N_7587,N_7800);
nor U8032 (N_8032,N_7818,N_7930);
nand U8033 (N_8033,N_7746,N_7736);
nor U8034 (N_8034,N_7671,N_7909);
and U8035 (N_8035,N_7706,N_7883);
nand U8036 (N_8036,N_7641,N_7960);
and U8037 (N_8037,N_7698,N_7924);
or U8038 (N_8038,N_7953,N_7597);
and U8039 (N_8039,N_7915,N_7998);
nand U8040 (N_8040,N_7546,N_7506);
or U8041 (N_8041,N_7561,N_7938);
or U8042 (N_8042,N_7630,N_7507);
or U8043 (N_8043,N_7645,N_7785);
nor U8044 (N_8044,N_7954,N_7908);
nand U8045 (N_8045,N_7872,N_7921);
or U8046 (N_8046,N_7999,N_7613);
or U8047 (N_8047,N_7759,N_7740);
and U8048 (N_8048,N_7791,N_7979);
or U8049 (N_8049,N_7699,N_7829);
nand U8050 (N_8050,N_7666,N_7589);
nand U8051 (N_8051,N_7583,N_7601);
nand U8052 (N_8052,N_7588,N_7835);
and U8053 (N_8053,N_7640,N_7989);
or U8054 (N_8054,N_7943,N_7790);
and U8055 (N_8055,N_7503,N_7539);
nor U8056 (N_8056,N_7725,N_7913);
nand U8057 (N_8057,N_7844,N_7766);
and U8058 (N_8058,N_7516,N_7530);
and U8059 (N_8059,N_7508,N_7767);
nand U8060 (N_8060,N_7551,N_7956);
nor U8061 (N_8061,N_7716,N_7802);
and U8062 (N_8062,N_7664,N_7959);
nor U8063 (N_8063,N_7529,N_7787);
nand U8064 (N_8064,N_7709,N_7607);
and U8065 (N_8065,N_7660,N_7717);
and U8066 (N_8066,N_7935,N_7794);
nor U8067 (N_8067,N_7547,N_7704);
nor U8068 (N_8068,N_7842,N_7809);
or U8069 (N_8069,N_7670,N_7578);
or U8070 (N_8070,N_7863,N_7808);
nor U8071 (N_8071,N_7940,N_7598);
and U8072 (N_8072,N_7786,N_7537);
nor U8073 (N_8073,N_7733,N_7629);
nand U8074 (N_8074,N_7584,N_7710);
nand U8075 (N_8075,N_7777,N_7775);
nand U8076 (N_8076,N_7502,N_7713);
nor U8077 (N_8077,N_7782,N_7948);
xor U8078 (N_8078,N_7887,N_7922);
nand U8079 (N_8079,N_7974,N_7894);
or U8080 (N_8080,N_7788,N_7694);
or U8081 (N_8081,N_7804,N_7779);
nor U8082 (N_8082,N_7554,N_7562);
or U8083 (N_8083,N_7504,N_7936);
xor U8084 (N_8084,N_7778,N_7643);
nand U8085 (N_8085,N_7620,N_7712);
or U8086 (N_8086,N_7637,N_7966);
nor U8087 (N_8087,N_7511,N_7895);
nand U8088 (N_8088,N_7968,N_7608);
or U8089 (N_8089,N_7754,N_7832);
and U8090 (N_8090,N_7651,N_7897);
nand U8091 (N_8091,N_7540,N_7867);
nand U8092 (N_8092,N_7510,N_7946);
nor U8093 (N_8093,N_7891,N_7911);
nor U8094 (N_8094,N_7569,N_7916);
or U8095 (N_8095,N_7923,N_7571);
nand U8096 (N_8096,N_7776,N_7991);
nor U8097 (N_8097,N_7855,N_7854);
and U8098 (N_8098,N_7614,N_7934);
and U8099 (N_8099,N_7967,N_7644);
nand U8100 (N_8100,N_7806,N_7830);
nor U8101 (N_8101,N_7944,N_7825);
xnor U8102 (N_8102,N_7873,N_7566);
or U8103 (N_8103,N_7552,N_7689);
or U8104 (N_8104,N_7980,N_7839);
nor U8105 (N_8105,N_7621,N_7847);
nand U8106 (N_8106,N_7892,N_7986);
nand U8107 (N_8107,N_7871,N_7995);
nor U8108 (N_8108,N_7850,N_7902);
and U8109 (N_8109,N_7877,N_7647);
xor U8110 (N_8110,N_7563,N_7889);
nor U8111 (N_8111,N_7941,N_7928);
nor U8112 (N_8112,N_7864,N_7674);
nand U8113 (N_8113,N_7860,N_7816);
nor U8114 (N_8114,N_7659,N_7618);
and U8115 (N_8115,N_7602,N_7550);
nand U8116 (N_8116,N_7683,N_7929);
nor U8117 (N_8117,N_7726,N_7885);
or U8118 (N_8118,N_7823,N_7665);
xor U8119 (N_8119,N_7837,N_7564);
or U8120 (N_8120,N_7965,N_7600);
nand U8121 (N_8121,N_7910,N_7815);
or U8122 (N_8122,N_7627,N_7500);
and U8123 (N_8123,N_7961,N_7807);
and U8124 (N_8124,N_7750,N_7635);
nor U8125 (N_8125,N_7730,N_7982);
xnor U8126 (N_8126,N_7751,N_7701);
or U8127 (N_8127,N_7692,N_7735);
nor U8128 (N_8128,N_7975,N_7515);
and U8129 (N_8129,N_7639,N_7682);
and U8130 (N_8130,N_7708,N_7610);
nor U8131 (N_8131,N_7840,N_7685);
nand U8132 (N_8132,N_7870,N_7905);
nor U8133 (N_8133,N_7762,N_7519);
and U8134 (N_8134,N_7882,N_7797);
nor U8135 (N_8135,N_7796,N_7667);
and U8136 (N_8136,N_7575,N_7719);
and U8137 (N_8137,N_7555,N_7903);
nand U8138 (N_8138,N_7693,N_7912);
or U8139 (N_8139,N_7755,N_7512);
nand U8140 (N_8140,N_7623,N_7646);
or U8141 (N_8141,N_7679,N_7942);
or U8142 (N_8142,N_7925,N_7874);
or U8143 (N_8143,N_7520,N_7846);
and U8144 (N_8144,N_7773,N_7955);
nor U8145 (N_8145,N_7605,N_7549);
nand U8146 (N_8146,N_7586,N_7747);
or U8147 (N_8147,N_7781,N_7609);
or U8148 (N_8148,N_7932,N_7557);
xnor U8149 (N_8149,N_7688,N_7675);
or U8150 (N_8150,N_7987,N_7714);
nand U8151 (N_8151,N_7983,N_7972);
xor U8152 (N_8152,N_7836,N_7758);
and U8153 (N_8153,N_7574,N_7729);
and U8154 (N_8154,N_7947,N_7522);
nand U8155 (N_8155,N_7594,N_7799);
or U8156 (N_8156,N_7743,N_7592);
or U8157 (N_8157,N_7538,N_7760);
or U8158 (N_8158,N_7749,N_7939);
nor U8159 (N_8159,N_7904,N_7501);
nand U8160 (N_8160,N_7591,N_7505);
or U8161 (N_8161,N_7531,N_7509);
nand U8162 (N_8162,N_7628,N_7653);
and U8163 (N_8163,N_7834,N_7696);
and U8164 (N_8164,N_7920,N_7560);
or U8165 (N_8165,N_7559,N_7687);
nand U8166 (N_8166,N_7763,N_7988);
nor U8167 (N_8167,N_7728,N_7851);
and U8168 (N_8168,N_7852,N_7526);
nand U8169 (N_8169,N_7814,N_7593);
nor U8170 (N_8170,N_7590,N_7723);
nor U8171 (N_8171,N_7642,N_7702);
and U8172 (N_8172,N_7572,N_7757);
or U8173 (N_8173,N_7535,N_7858);
and U8174 (N_8174,N_7949,N_7724);
nor U8175 (N_8175,N_7721,N_7826);
nor U8176 (N_8176,N_7876,N_7582);
and U8177 (N_8177,N_7774,N_7937);
or U8178 (N_8178,N_7756,N_7573);
or U8179 (N_8179,N_7784,N_7994);
xnor U8180 (N_8180,N_7833,N_7541);
and U8181 (N_8181,N_7527,N_7532);
nand U8182 (N_8182,N_7899,N_7780);
and U8183 (N_8183,N_7845,N_7798);
or U8184 (N_8184,N_7772,N_7886);
or U8185 (N_8185,N_7669,N_7700);
nand U8186 (N_8186,N_7793,N_7856);
or U8187 (N_8187,N_7684,N_7707);
xnor U8188 (N_8188,N_7673,N_7691);
xor U8189 (N_8189,N_7633,N_7663);
nand U8190 (N_8190,N_7984,N_7553);
nand U8191 (N_8191,N_7525,N_7612);
or U8192 (N_8192,N_7731,N_7718);
or U8193 (N_8193,N_7878,N_7869);
nor U8194 (N_8194,N_7761,N_7849);
or U8195 (N_8195,N_7831,N_7534);
xnor U8196 (N_8196,N_7810,N_7568);
and U8197 (N_8197,N_7859,N_7841);
or U8198 (N_8198,N_7861,N_7711);
nor U8199 (N_8199,N_7655,N_7741);
nor U8200 (N_8200,N_7523,N_7705);
and U8201 (N_8201,N_7611,N_7686);
and U8202 (N_8202,N_7992,N_7567);
and U8203 (N_8203,N_7681,N_7720);
nor U8204 (N_8204,N_7821,N_7857);
nand U8205 (N_8205,N_7548,N_7973);
nand U8206 (N_8206,N_7971,N_7565);
and U8207 (N_8207,N_7838,N_7622);
nand U8208 (N_8208,N_7604,N_7648);
and U8209 (N_8209,N_7680,N_7978);
nor U8210 (N_8210,N_7580,N_7558);
nor U8211 (N_8211,N_7985,N_7896);
nor U8212 (N_8212,N_7907,N_7914);
nor U8213 (N_8213,N_7963,N_7715);
nor U8214 (N_8214,N_7672,N_7596);
and U8215 (N_8215,N_7812,N_7990);
xnor U8216 (N_8216,N_7697,N_7957);
or U8217 (N_8217,N_7848,N_7677);
or U8218 (N_8218,N_7824,N_7976);
xnor U8219 (N_8219,N_7853,N_7662);
and U8220 (N_8220,N_7656,N_7676);
nor U8221 (N_8221,N_7901,N_7931);
and U8222 (N_8222,N_7661,N_7603);
and U8223 (N_8223,N_7513,N_7649);
nand U8224 (N_8224,N_7595,N_7822);
nor U8225 (N_8225,N_7918,N_7585);
nor U8226 (N_8226,N_7969,N_7606);
and U8227 (N_8227,N_7631,N_7951);
nand U8228 (N_8228,N_7636,N_7866);
nor U8229 (N_8229,N_7828,N_7769);
nand U8230 (N_8230,N_7771,N_7545);
nand U8231 (N_8231,N_7827,N_7898);
and U8232 (N_8232,N_7657,N_7652);
and U8233 (N_8233,N_7536,N_7927);
or U8234 (N_8234,N_7981,N_7795);
or U8235 (N_8235,N_7632,N_7801);
nand U8236 (N_8236,N_7919,N_7997);
nor U8237 (N_8237,N_7518,N_7543);
xnor U8238 (N_8238,N_7996,N_7528);
and U8239 (N_8239,N_7745,N_7792);
nor U8240 (N_8240,N_7843,N_7695);
xor U8241 (N_8241,N_7770,N_7752);
xor U8242 (N_8242,N_7917,N_7690);
and U8243 (N_8243,N_7879,N_7619);
nand U8244 (N_8244,N_7626,N_7658);
or U8245 (N_8245,N_7744,N_7900);
nor U8246 (N_8246,N_7524,N_7650);
nand U8247 (N_8247,N_7945,N_7517);
nand U8248 (N_8248,N_7753,N_7926);
nor U8249 (N_8249,N_7890,N_7521);
and U8250 (N_8250,N_7731,N_7817);
or U8251 (N_8251,N_7965,N_7700);
nand U8252 (N_8252,N_7643,N_7542);
nor U8253 (N_8253,N_7605,N_7962);
and U8254 (N_8254,N_7879,N_7858);
xnor U8255 (N_8255,N_7820,N_7717);
and U8256 (N_8256,N_7960,N_7928);
nor U8257 (N_8257,N_7583,N_7826);
nand U8258 (N_8258,N_7714,N_7796);
or U8259 (N_8259,N_7619,N_7540);
or U8260 (N_8260,N_7566,N_7895);
and U8261 (N_8261,N_7961,N_7595);
xor U8262 (N_8262,N_7964,N_7676);
or U8263 (N_8263,N_7890,N_7704);
nand U8264 (N_8264,N_7934,N_7754);
or U8265 (N_8265,N_7996,N_7631);
nand U8266 (N_8266,N_7574,N_7511);
or U8267 (N_8267,N_7684,N_7817);
xnor U8268 (N_8268,N_7898,N_7862);
or U8269 (N_8269,N_7916,N_7664);
nand U8270 (N_8270,N_7584,N_7526);
nand U8271 (N_8271,N_7881,N_7892);
nor U8272 (N_8272,N_7969,N_7999);
and U8273 (N_8273,N_7723,N_7867);
nand U8274 (N_8274,N_7730,N_7567);
xnor U8275 (N_8275,N_7938,N_7538);
nor U8276 (N_8276,N_7538,N_7798);
or U8277 (N_8277,N_7593,N_7718);
and U8278 (N_8278,N_7776,N_7810);
nand U8279 (N_8279,N_7781,N_7651);
and U8280 (N_8280,N_7513,N_7947);
nand U8281 (N_8281,N_7634,N_7820);
or U8282 (N_8282,N_7559,N_7934);
or U8283 (N_8283,N_7636,N_7925);
and U8284 (N_8284,N_7765,N_7629);
nand U8285 (N_8285,N_7643,N_7795);
and U8286 (N_8286,N_7990,N_7808);
or U8287 (N_8287,N_7811,N_7506);
and U8288 (N_8288,N_7890,N_7782);
xor U8289 (N_8289,N_7888,N_7929);
or U8290 (N_8290,N_7503,N_7757);
nand U8291 (N_8291,N_7873,N_7996);
nor U8292 (N_8292,N_7697,N_7574);
nor U8293 (N_8293,N_7539,N_7669);
xor U8294 (N_8294,N_7780,N_7542);
and U8295 (N_8295,N_7854,N_7607);
nor U8296 (N_8296,N_7866,N_7590);
xor U8297 (N_8297,N_7883,N_7746);
nor U8298 (N_8298,N_7879,N_7767);
nor U8299 (N_8299,N_7934,N_7810);
and U8300 (N_8300,N_7883,N_7578);
or U8301 (N_8301,N_7700,N_7900);
xnor U8302 (N_8302,N_7849,N_7854);
nor U8303 (N_8303,N_7527,N_7932);
or U8304 (N_8304,N_7795,N_7646);
or U8305 (N_8305,N_7744,N_7579);
xnor U8306 (N_8306,N_7696,N_7769);
and U8307 (N_8307,N_7919,N_7809);
or U8308 (N_8308,N_7557,N_7878);
nor U8309 (N_8309,N_7633,N_7895);
xor U8310 (N_8310,N_7905,N_7685);
nor U8311 (N_8311,N_7784,N_7589);
nor U8312 (N_8312,N_7552,N_7679);
nor U8313 (N_8313,N_7930,N_7898);
nand U8314 (N_8314,N_7836,N_7830);
and U8315 (N_8315,N_7978,N_7833);
nand U8316 (N_8316,N_7940,N_7664);
nor U8317 (N_8317,N_7860,N_7749);
nor U8318 (N_8318,N_7881,N_7711);
nand U8319 (N_8319,N_7834,N_7531);
xnor U8320 (N_8320,N_7516,N_7961);
or U8321 (N_8321,N_7936,N_7899);
nand U8322 (N_8322,N_7537,N_7931);
nand U8323 (N_8323,N_7788,N_7580);
or U8324 (N_8324,N_7618,N_7938);
and U8325 (N_8325,N_7684,N_7515);
xor U8326 (N_8326,N_7807,N_7653);
and U8327 (N_8327,N_7821,N_7795);
or U8328 (N_8328,N_7763,N_7947);
nor U8329 (N_8329,N_7786,N_7829);
and U8330 (N_8330,N_7743,N_7832);
or U8331 (N_8331,N_7848,N_7565);
or U8332 (N_8332,N_7539,N_7963);
nand U8333 (N_8333,N_7876,N_7500);
nand U8334 (N_8334,N_7744,N_7851);
nand U8335 (N_8335,N_7763,N_7769);
nand U8336 (N_8336,N_7945,N_7629);
and U8337 (N_8337,N_7902,N_7774);
and U8338 (N_8338,N_7963,N_7671);
or U8339 (N_8339,N_7815,N_7500);
or U8340 (N_8340,N_7853,N_7534);
nor U8341 (N_8341,N_7990,N_7739);
nand U8342 (N_8342,N_7501,N_7780);
xnor U8343 (N_8343,N_7692,N_7908);
or U8344 (N_8344,N_7632,N_7858);
xor U8345 (N_8345,N_7962,N_7980);
nand U8346 (N_8346,N_7934,N_7563);
or U8347 (N_8347,N_7540,N_7930);
or U8348 (N_8348,N_7841,N_7544);
nand U8349 (N_8349,N_7711,N_7992);
or U8350 (N_8350,N_7856,N_7852);
or U8351 (N_8351,N_7675,N_7732);
and U8352 (N_8352,N_7919,N_7846);
nand U8353 (N_8353,N_7901,N_7856);
nor U8354 (N_8354,N_7854,N_7696);
nand U8355 (N_8355,N_7894,N_7743);
or U8356 (N_8356,N_7510,N_7637);
and U8357 (N_8357,N_7778,N_7687);
nor U8358 (N_8358,N_7721,N_7586);
nand U8359 (N_8359,N_7832,N_7874);
or U8360 (N_8360,N_7634,N_7883);
nand U8361 (N_8361,N_7656,N_7595);
xnor U8362 (N_8362,N_7826,N_7852);
or U8363 (N_8363,N_7587,N_7556);
nor U8364 (N_8364,N_7719,N_7940);
nor U8365 (N_8365,N_7931,N_7895);
or U8366 (N_8366,N_7721,N_7650);
and U8367 (N_8367,N_7602,N_7502);
nor U8368 (N_8368,N_7579,N_7571);
nand U8369 (N_8369,N_7808,N_7840);
and U8370 (N_8370,N_7583,N_7774);
nand U8371 (N_8371,N_7608,N_7637);
nor U8372 (N_8372,N_7931,N_7532);
or U8373 (N_8373,N_7904,N_7844);
and U8374 (N_8374,N_7767,N_7561);
and U8375 (N_8375,N_7617,N_7709);
or U8376 (N_8376,N_7804,N_7764);
or U8377 (N_8377,N_7776,N_7963);
and U8378 (N_8378,N_7925,N_7633);
or U8379 (N_8379,N_7538,N_7704);
or U8380 (N_8380,N_7592,N_7553);
nor U8381 (N_8381,N_7615,N_7641);
nor U8382 (N_8382,N_7512,N_7848);
nand U8383 (N_8383,N_7530,N_7827);
and U8384 (N_8384,N_7732,N_7589);
nand U8385 (N_8385,N_7906,N_7855);
nand U8386 (N_8386,N_7838,N_7632);
nand U8387 (N_8387,N_7875,N_7970);
or U8388 (N_8388,N_7894,N_7952);
nor U8389 (N_8389,N_7941,N_7561);
or U8390 (N_8390,N_7984,N_7856);
and U8391 (N_8391,N_7622,N_7832);
nor U8392 (N_8392,N_7932,N_7704);
and U8393 (N_8393,N_7650,N_7967);
nand U8394 (N_8394,N_7543,N_7509);
nand U8395 (N_8395,N_7825,N_7696);
nor U8396 (N_8396,N_7637,N_7994);
and U8397 (N_8397,N_7627,N_7907);
xor U8398 (N_8398,N_7519,N_7586);
or U8399 (N_8399,N_7875,N_7589);
nand U8400 (N_8400,N_7889,N_7863);
or U8401 (N_8401,N_7830,N_7505);
nor U8402 (N_8402,N_7554,N_7970);
xnor U8403 (N_8403,N_7846,N_7546);
and U8404 (N_8404,N_7760,N_7658);
and U8405 (N_8405,N_7530,N_7811);
or U8406 (N_8406,N_7650,N_7724);
and U8407 (N_8407,N_7504,N_7800);
or U8408 (N_8408,N_7520,N_7635);
and U8409 (N_8409,N_7630,N_7790);
and U8410 (N_8410,N_7721,N_7926);
nor U8411 (N_8411,N_7525,N_7651);
nand U8412 (N_8412,N_7921,N_7648);
or U8413 (N_8413,N_7551,N_7558);
nand U8414 (N_8414,N_7560,N_7525);
xnor U8415 (N_8415,N_7988,N_7910);
and U8416 (N_8416,N_7667,N_7742);
nor U8417 (N_8417,N_7988,N_7774);
nand U8418 (N_8418,N_7639,N_7857);
xnor U8419 (N_8419,N_7737,N_7889);
and U8420 (N_8420,N_7995,N_7801);
nand U8421 (N_8421,N_7852,N_7564);
and U8422 (N_8422,N_7537,N_7908);
and U8423 (N_8423,N_7528,N_7971);
nand U8424 (N_8424,N_7611,N_7766);
and U8425 (N_8425,N_7965,N_7830);
or U8426 (N_8426,N_7666,N_7717);
nor U8427 (N_8427,N_7636,N_7953);
nor U8428 (N_8428,N_7516,N_7659);
or U8429 (N_8429,N_7666,N_7502);
nor U8430 (N_8430,N_7677,N_7553);
and U8431 (N_8431,N_7857,N_7647);
nand U8432 (N_8432,N_7869,N_7520);
nand U8433 (N_8433,N_7875,N_7780);
and U8434 (N_8434,N_7816,N_7775);
nor U8435 (N_8435,N_7526,N_7962);
or U8436 (N_8436,N_7560,N_7757);
nor U8437 (N_8437,N_7820,N_7645);
nand U8438 (N_8438,N_7963,N_7548);
nor U8439 (N_8439,N_7914,N_7791);
nor U8440 (N_8440,N_7894,N_7844);
and U8441 (N_8441,N_7640,N_7619);
or U8442 (N_8442,N_7716,N_7852);
nand U8443 (N_8443,N_7613,N_7745);
or U8444 (N_8444,N_7985,N_7884);
nand U8445 (N_8445,N_7822,N_7775);
or U8446 (N_8446,N_7581,N_7653);
or U8447 (N_8447,N_7733,N_7681);
xnor U8448 (N_8448,N_7865,N_7961);
nor U8449 (N_8449,N_7522,N_7871);
and U8450 (N_8450,N_7794,N_7511);
and U8451 (N_8451,N_7965,N_7784);
or U8452 (N_8452,N_7798,N_7764);
nand U8453 (N_8453,N_7545,N_7559);
or U8454 (N_8454,N_7605,N_7834);
or U8455 (N_8455,N_7740,N_7881);
and U8456 (N_8456,N_7672,N_7638);
nor U8457 (N_8457,N_7731,N_7599);
or U8458 (N_8458,N_7911,N_7643);
nor U8459 (N_8459,N_7793,N_7740);
and U8460 (N_8460,N_7525,N_7541);
nor U8461 (N_8461,N_7544,N_7835);
nor U8462 (N_8462,N_7762,N_7752);
and U8463 (N_8463,N_7722,N_7998);
and U8464 (N_8464,N_7612,N_7506);
nand U8465 (N_8465,N_7797,N_7510);
nand U8466 (N_8466,N_7970,N_7623);
xnor U8467 (N_8467,N_7790,N_7920);
nand U8468 (N_8468,N_7884,N_7836);
or U8469 (N_8469,N_7527,N_7759);
or U8470 (N_8470,N_7898,N_7942);
xnor U8471 (N_8471,N_7710,N_7960);
nand U8472 (N_8472,N_7754,N_7534);
or U8473 (N_8473,N_7990,N_7679);
or U8474 (N_8474,N_7780,N_7729);
and U8475 (N_8475,N_7887,N_7778);
nand U8476 (N_8476,N_7735,N_7706);
or U8477 (N_8477,N_7523,N_7751);
and U8478 (N_8478,N_7809,N_7665);
nand U8479 (N_8479,N_7931,N_7611);
nor U8480 (N_8480,N_7631,N_7558);
nand U8481 (N_8481,N_7750,N_7633);
and U8482 (N_8482,N_7619,N_7844);
and U8483 (N_8483,N_7890,N_7894);
and U8484 (N_8484,N_7883,N_7769);
or U8485 (N_8485,N_7800,N_7574);
nor U8486 (N_8486,N_7723,N_7779);
nor U8487 (N_8487,N_7560,N_7606);
nor U8488 (N_8488,N_7572,N_7728);
or U8489 (N_8489,N_7708,N_7511);
or U8490 (N_8490,N_7532,N_7735);
nor U8491 (N_8491,N_7626,N_7747);
and U8492 (N_8492,N_7747,N_7647);
nand U8493 (N_8493,N_7926,N_7863);
nand U8494 (N_8494,N_7955,N_7859);
nor U8495 (N_8495,N_7809,N_7973);
nand U8496 (N_8496,N_7972,N_7862);
xor U8497 (N_8497,N_7739,N_7753);
and U8498 (N_8498,N_7762,N_7758);
nor U8499 (N_8499,N_7555,N_7974);
nor U8500 (N_8500,N_8122,N_8436);
or U8501 (N_8501,N_8393,N_8205);
nand U8502 (N_8502,N_8408,N_8375);
xor U8503 (N_8503,N_8415,N_8155);
and U8504 (N_8504,N_8254,N_8282);
xor U8505 (N_8505,N_8230,N_8276);
nand U8506 (N_8506,N_8498,N_8462);
nor U8507 (N_8507,N_8249,N_8487);
nand U8508 (N_8508,N_8416,N_8484);
and U8509 (N_8509,N_8043,N_8466);
nor U8510 (N_8510,N_8026,N_8104);
and U8511 (N_8511,N_8397,N_8123);
nand U8512 (N_8512,N_8495,N_8364);
nand U8513 (N_8513,N_8022,N_8417);
and U8514 (N_8514,N_8346,N_8036);
or U8515 (N_8515,N_8315,N_8423);
nor U8516 (N_8516,N_8051,N_8030);
nand U8517 (N_8517,N_8363,N_8367);
and U8518 (N_8518,N_8180,N_8300);
or U8519 (N_8519,N_8211,N_8110);
nand U8520 (N_8520,N_8455,N_8134);
nor U8521 (N_8521,N_8279,N_8411);
or U8522 (N_8522,N_8214,N_8328);
nand U8523 (N_8523,N_8251,N_8304);
and U8524 (N_8524,N_8437,N_8331);
nor U8525 (N_8525,N_8201,N_8053);
and U8526 (N_8526,N_8366,N_8118);
nor U8527 (N_8527,N_8075,N_8137);
and U8528 (N_8528,N_8133,N_8294);
nand U8529 (N_8529,N_8035,N_8139);
and U8530 (N_8530,N_8243,N_8383);
and U8531 (N_8531,N_8309,N_8336);
or U8532 (N_8532,N_8358,N_8247);
or U8533 (N_8533,N_8096,N_8368);
nor U8534 (N_8534,N_8070,N_8019);
and U8535 (N_8535,N_8492,N_8288);
or U8536 (N_8536,N_8355,N_8089);
nor U8537 (N_8537,N_8079,N_8322);
nand U8538 (N_8538,N_8285,N_8156);
and U8539 (N_8539,N_8373,N_8286);
nor U8540 (N_8540,N_8164,N_8112);
nor U8541 (N_8541,N_8120,N_8460);
nor U8542 (N_8542,N_8266,N_8225);
or U8543 (N_8543,N_8080,N_8493);
nor U8544 (N_8544,N_8277,N_8024);
xnor U8545 (N_8545,N_8206,N_8392);
nand U8546 (N_8546,N_8319,N_8356);
or U8547 (N_8547,N_8153,N_8264);
or U8548 (N_8548,N_8441,N_8342);
nand U8549 (N_8549,N_8138,N_8208);
nor U8550 (N_8550,N_8020,N_8330);
and U8551 (N_8551,N_8385,N_8056);
or U8552 (N_8552,N_8376,N_8023);
nand U8553 (N_8553,N_8052,N_8351);
nand U8554 (N_8554,N_8181,N_8165);
and U8555 (N_8555,N_8060,N_8203);
nor U8556 (N_8556,N_8287,N_8188);
nand U8557 (N_8557,N_8109,N_8433);
nand U8558 (N_8558,N_8413,N_8042);
and U8559 (N_8559,N_8017,N_8140);
nand U8560 (N_8560,N_8103,N_8320);
and U8561 (N_8561,N_8174,N_8175);
nand U8562 (N_8562,N_8260,N_8057);
nor U8563 (N_8563,N_8069,N_8152);
nand U8564 (N_8564,N_8028,N_8115);
and U8565 (N_8565,N_8407,N_8136);
nand U8566 (N_8566,N_8298,N_8268);
nor U8567 (N_8567,N_8278,N_8015);
xor U8568 (N_8568,N_8475,N_8173);
nand U8569 (N_8569,N_8159,N_8077);
xnor U8570 (N_8570,N_8410,N_8442);
and U8571 (N_8571,N_8213,N_8388);
and U8572 (N_8572,N_8100,N_8227);
xor U8573 (N_8573,N_8339,N_8337);
nand U8574 (N_8574,N_8325,N_8202);
nand U8575 (N_8575,N_8114,N_8255);
or U8576 (N_8576,N_8234,N_8222);
and U8577 (N_8577,N_8365,N_8468);
or U8578 (N_8578,N_8360,N_8435);
nand U8579 (N_8579,N_8326,N_8353);
or U8580 (N_8580,N_8029,N_8135);
and U8581 (N_8581,N_8297,N_8160);
xor U8582 (N_8582,N_8169,N_8296);
and U8583 (N_8583,N_8073,N_8163);
and U8584 (N_8584,N_8018,N_8485);
or U8585 (N_8585,N_8039,N_8207);
or U8586 (N_8586,N_8049,N_8313);
xor U8587 (N_8587,N_8419,N_8065);
and U8588 (N_8588,N_8497,N_8426);
nor U8589 (N_8589,N_8293,N_8223);
or U8590 (N_8590,N_8246,N_8295);
nand U8591 (N_8591,N_8305,N_8098);
and U8592 (N_8592,N_8198,N_8094);
xnor U8593 (N_8593,N_8220,N_8302);
nand U8594 (N_8594,N_8312,N_8184);
nand U8595 (N_8595,N_8479,N_8438);
or U8596 (N_8596,N_8146,N_8378);
or U8597 (N_8597,N_8116,N_8344);
nand U8598 (N_8598,N_8352,N_8003);
nor U8599 (N_8599,N_8008,N_8168);
nor U8600 (N_8600,N_8464,N_8387);
nand U8601 (N_8601,N_8093,N_8239);
xnor U8602 (N_8602,N_8161,N_8384);
nand U8603 (N_8603,N_8209,N_8048);
and U8604 (N_8604,N_8306,N_8290);
nor U8605 (N_8605,N_8047,N_8476);
nor U8606 (N_8606,N_8199,N_8228);
xnor U8607 (N_8607,N_8252,N_8263);
and U8608 (N_8608,N_8453,N_8142);
nor U8609 (N_8609,N_8217,N_8004);
or U8610 (N_8610,N_8126,N_8045);
nor U8611 (N_8611,N_8481,N_8350);
nand U8612 (N_8612,N_8055,N_8488);
nor U8613 (N_8613,N_8427,N_8005);
and U8614 (N_8614,N_8265,N_8068);
or U8615 (N_8615,N_8292,N_8391);
and U8616 (N_8616,N_8235,N_8272);
or U8617 (N_8617,N_8379,N_8374);
and U8618 (N_8618,N_8333,N_8002);
nand U8619 (N_8619,N_8483,N_8066);
nand U8620 (N_8620,N_8324,N_8218);
and U8621 (N_8621,N_8021,N_8113);
or U8622 (N_8622,N_8398,N_8219);
nor U8623 (N_8623,N_8414,N_8171);
and U8624 (N_8624,N_8038,N_8480);
and U8625 (N_8625,N_8395,N_8041);
nor U8626 (N_8626,N_8046,N_8095);
nand U8627 (N_8627,N_8000,N_8025);
nor U8628 (N_8628,N_8237,N_8308);
nand U8629 (N_8629,N_8341,N_8486);
or U8630 (N_8630,N_8314,N_8033);
nor U8631 (N_8631,N_8338,N_8343);
nand U8632 (N_8632,N_8177,N_8016);
or U8633 (N_8633,N_8001,N_8143);
and U8634 (N_8634,N_8196,N_8490);
and U8635 (N_8635,N_8489,N_8221);
or U8636 (N_8636,N_8145,N_8244);
or U8637 (N_8637,N_8061,N_8409);
or U8638 (N_8638,N_8245,N_8463);
nand U8639 (N_8639,N_8076,N_8499);
nand U8640 (N_8640,N_8050,N_8081);
xnor U8641 (N_8641,N_8162,N_8191);
nor U8642 (N_8642,N_8248,N_8399);
xor U8643 (N_8643,N_8108,N_8232);
and U8644 (N_8644,N_8386,N_8451);
xnor U8645 (N_8645,N_8179,N_8403);
nand U8646 (N_8646,N_8259,N_8151);
nor U8647 (N_8647,N_8470,N_8348);
nand U8648 (N_8648,N_8370,N_8064);
or U8649 (N_8649,N_8456,N_8054);
nor U8650 (N_8650,N_8258,N_8400);
nand U8651 (N_8651,N_8382,N_8147);
nand U8652 (N_8652,N_8284,N_8472);
xor U8653 (N_8653,N_8271,N_8197);
or U8654 (N_8654,N_8212,N_8347);
or U8655 (N_8655,N_8085,N_8090);
and U8656 (N_8656,N_8121,N_8185);
and U8657 (N_8657,N_8450,N_8394);
or U8658 (N_8658,N_8454,N_8241);
and U8659 (N_8659,N_8253,N_8105);
nor U8660 (N_8660,N_8469,N_8083);
nand U8661 (N_8661,N_8091,N_8187);
or U8662 (N_8662,N_8310,N_8461);
and U8663 (N_8663,N_8011,N_8465);
or U8664 (N_8664,N_8457,N_8210);
and U8665 (N_8665,N_8111,N_8067);
nor U8666 (N_8666,N_8215,N_8086);
nand U8667 (N_8667,N_8131,N_8377);
nand U8668 (N_8668,N_8381,N_8372);
or U8669 (N_8669,N_8327,N_8303);
and U8670 (N_8670,N_8178,N_8194);
or U8671 (N_8671,N_8006,N_8148);
nor U8672 (N_8672,N_8154,N_8291);
or U8673 (N_8673,N_8473,N_8270);
and U8674 (N_8674,N_8170,N_8149);
and U8675 (N_8675,N_8158,N_8236);
nor U8676 (N_8676,N_8396,N_8299);
or U8677 (N_8677,N_8283,N_8329);
nand U8678 (N_8678,N_8013,N_8340);
xor U8679 (N_8679,N_8204,N_8354);
xor U8680 (N_8680,N_8192,N_8256);
nand U8681 (N_8681,N_8032,N_8150);
or U8682 (N_8682,N_8014,N_8183);
and U8683 (N_8683,N_8088,N_8301);
or U8684 (N_8684,N_8405,N_8037);
nor U8685 (N_8685,N_8467,N_8471);
and U8686 (N_8686,N_8072,N_8380);
nor U8687 (N_8687,N_8242,N_8474);
nor U8688 (N_8688,N_8349,N_8157);
or U8689 (N_8689,N_8063,N_8097);
nand U8690 (N_8690,N_8010,N_8269);
nor U8691 (N_8691,N_8362,N_8318);
nand U8692 (N_8692,N_8240,N_8231);
nand U8693 (N_8693,N_8430,N_8311);
nand U8694 (N_8694,N_8317,N_8084);
or U8695 (N_8695,N_8401,N_8267);
nand U8696 (N_8696,N_8273,N_8429);
nand U8697 (N_8697,N_8425,N_8216);
and U8698 (N_8698,N_8321,N_8458);
xnor U8699 (N_8699,N_8117,N_8332);
and U8700 (N_8700,N_8129,N_8390);
nor U8701 (N_8701,N_8224,N_8092);
xnor U8702 (N_8702,N_8238,N_8359);
nor U8703 (N_8703,N_8262,N_8074);
nor U8704 (N_8704,N_8034,N_8130);
and U8705 (N_8705,N_8418,N_8452);
or U8706 (N_8706,N_8007,N_8281);
and U8707 (N_8707,N_8477,N_8428);
or U8708 (N_8708,N_8141,N_8494);
xnor U8709 (N_8709,N_8449,N_8369);
nand U8710 (N_8710,N_8482,N_8044);
nor U8711 (N_8711,N_8058,N_8389);
or U8712 (N_8712,N_8127,N_8186);
nor U8713 (N_8713,N_8446,N_8226);
or U8714 (N_8714,N_8334,N_8439);
and U8715 (N_8715,N_8361,N_8009);
or U8716 (N_8716,N_8193,N_8357);
nor U8717 (N_8717,N_8445,N_8345);
or U8718 (N_8718,N_8106,N_8335);
nand U8719 (N_8719,N_8402,N_8406);
or U8720 (N_8720,N_8099,N_8434);
xor U8721 (N_8721,N_8448,N_8078);
nand U8722 (N_8722,N_8189,N_8459);
nand U8723 (N_8723,N_8440,N_8082);
and U8724 (N_8724,N_8443,N_8424);
xnor U8725 (N_8725,N_8275,N_8059);
and U8726 (N_8726,N_8200,N_8027);
nor U8727 (N_8727,N_8444,N_8229);
nand U8728 (N_8728,N_8166,N_8420);
nand U8729 (N_8729,N_8132,N_8031);
or U8730 (N_8730,N_8280,N_8107);
nor U8731 (N_8731,N_8431,N_8167);
or U8732 (N_8732,N_8087,N_8257);
or U8733 (N_8733,N_8119,N_8233);
or U8734 (N_8734,N_8062,N_8101);
and U8735 (N_8735,N_8478,N_8404);
nor U8736 (N_8736,N_8307,N_8316);
or U8737 (N_8737,N_8172,N_8412);
and U8738 (N_8738,N_8422,N_8182);
and U8739 (N_8739,N_8012,N_8124);
nand U8740 (N_8740,N_8250,N_8274);
and U8741 (N_8741,N_8195,N_8421);
nor U8742 (N_8742,N_8040,N_8261);
nand U8743 (N_8743,N_8190,N_8323);
nor U8744 (N_8744,N_8102,N_8432);
nor U8745 (N_8745,N_8289,N_8371);
or U8746 (N_8746,N_8491,N_8447);
and U8747 (N_8747,N_8071,N_8125);
nand U8748 (N_8748,N_8128,N_8176);
and U8749 (N_8749,N_8496,N_8144);
and U8750 (N_8750,N_8148,N_8286);
xor U8751 (N_8751,N_8420,N_8389);
nand U8752 (N_8752,N_8011,N_8410);
nor U8753 (N_8753,N_8109,N_8175);
nor U8754 (N_8754,N_8232,N_8446);
xor U8755 (N_8755,N_8283,N_8425);
xnor U8756 (N_8756,N_8037,N_8072);
and U8757 (N_8757,N_8026,N_8428);
xnor U8758 (N_8758,N_8283,N_8476);
nand U8759 (N_8759,N_8238,N_8352);
nand U8760 (N_8760,N_8355,N_8337);
nor U8761 (N_8761,N_8224,N_8365);
or U8762 (N_8762,N_8218,N_8335);
nand U8763 (N_8763,N_8479,N_8029);
or U8764 (N_8764,N_8085,N_8010);
and U8765 (N_8765,N_8038,N_8048);
and U8766 (N_8766,N_8346,N_8050);
nor U8767 (N_8767,N_8393,N_8423);
xor U8768 (N_8768,N_8018,N_8330);
nand U8769 (N_8769,N_8482,N_8460);
and U8770 (N_8770,N_8041,N_8147);
and U8771 (N_8771,N_8204,N_8394);
and U8772 (N_8772,N_8118,N_8450);
nand U8773 (N_8773,N_8007,N_8203);
or U8774 (N_8774,N_8305,N_8329);
or U8775 (N_8775,N_8451,N_8461);
or U8776 (N_8776,N_8367,N_8316);
and U8777 (N_8777,N_8427,N_8456);
nor U8778 (N_8778,N_8305,N_8263);
nor U8779 (N_8779,N_8061,N_8457);
or U8780 (N_8780,N_8151,N_8369);
xor U8781 (N_8781,N_8327,N_8026);
or U8782 (N_8782,N_8282,N_8004);
nor U8783 (N_8783,N_8274,N_8049);
or U8784 (N_8784,N_8451,N_8109);
xor U8785 (N_8785,N_8155,N_8085);
and U8786 (N_8786,N_8197,N_8121);
nand U8787 (N_8787,N_8005,N_8050);
and U8788 (N_8788,N_8062,N_8494);
and U8789 (N_8789,N_8123,N_8414);
nor U8790 (N_8790,N_8380,N_8389);
nor U8791 (N_8791,N_8115,N_8162);
nand U8792 (N_8792,N_8243,N_8455);
or U8793 (N_8793,N_8193,N_8049);
or U8794 (N_8794,N_8049,N_8201);
and U8795 (N_8795,N_8181,N_8119);
nor U8796 (N_8796,N_8059,N_8024);
and U8797 (N_8797,N_8047,N_8013);
nor U8798 (N_8798,N_8353,N_8080);
nor U8799 (N_8799,N_8265,N_8278);
nand U8800 (N_8800,N_8320,N_8045);
or U8801 (N_8801,N_8113,N_8180);
nand U8802 (N_8802,N_8230,N_8045);
or U8803 (N_8803,N_8364,N_8108);
and U8804 (N_8804,N_8464,N_8073);
and U8805 (N_8805,N_8176,N_8489);
and U8806 (N_8806,N_8211,N_8056);
xor U8807 (N_8807,N_8183,N_8483);
nand U8808 (N_8808,N_8452,N_8287);
nand U8809 (N_8809,N_8430,N_8152);
and U8810 (N_8810,N_8241,N_8123);
nor U8811 (N_8811,N_8358,N_8315);
or U8812 (N_8812,N_8083,N_8180);
and U8813 (N_8813,N_8197,N_8352);
and U8814 (N_8814,N_8315,N_8416);
nand U8815 (N_8815,N_8143,N_8290);
or U8816 (N_8816,N_8087,N_8466);
nor U8817 (N_8817,N_8279,N_8201);
or U8818 (N_8818,N_8317,N_8235);
nor U8819 (N_8819,N_8114,N_8137);
xnor U8820 (N_8820,N_8082,N_8254);
nand U8821 (N_8821,N_8440,N_8124);
xor U8822 (N_8822,N_8181,N_8184);
nor U8823 (N_8823,N_8423,N_8173);
xor U8824 (N_8824,N_8072,N_8137);
nand U8825 (N_8825,N_8103,N_8180);
nor U8826 (N_8826,N_8431,N_8393);
and U8827 (N_8827,N_8038,N_8475);
or U8828 (N_8828,N_8323,N_8202);
nor U8829 (N_8829,N_8179,N_8351);
nor U8830 (N_8830,N_8300,N_8165);
nand U8831 (N_8831,N_8236,N_8432);
and U8832 (N_8832,N_8067,N_8106);
nand U8833 (N_8833,N_8028,N_8289);
nor U8834 (N_8834,N_8057,N_8085);
nand U8835 (N_8835,N_8184,N_8356);
nor U8836 (N_8836,N_8143,N_8220);
nand U8837 (N_8837,N_8461,N_8061);
nand U8838 (N_8838,N_8308,N_8132);
or U8839 (N_8839,N_8034,N_8013);
nand U8840 (N_8840,N_8167,N_8009);
nor U8841 (N_8841,N_8192,N_8057);
or U8842 (N_8842,N_8279,N_8066);
nand U8843 (N_8843,N_8184,N_8225);
nor U8844 (N_8844,N_8024,N_8010);
nand U8845 (N_8845,N_8349,N_8281);
and U8846 (N_8846,N_8350,N_8169);
nor U8847 (N_8847,N_8243,N_8415);
or U8848 (N_8848,N_8181,N_8487);
xnor U8849 (N_8849,N_8178,N_8173);
nor U8850 (N_8850,N_8164,N_8190);
nand U8851 (N_8851,N_8320,N_8396);
nand U8852 (N_8852,N_8079,N_8096);
or U8853 (N_8853,N_8170,N_8395);
xnor U8854 (N_8854,N_8128,N_8224);
nor U8855 (N_8855,N_8099,N_8042);
nand U8856 (N_8856,N_8365,N_8344);
or U8857 (N_8857,N_8495,N_8119);
nor U8858 (N_8858,N_8079,N_8069);
or U8859 (N_8859,N_8003,N_8063);
nand U8860 (N_8860,N_8170,N_8112);
nand U8861 (N_8861,N_8394,N_8140);
nor U8862 (N_8862,N_8235,N_8321);
nor U8863 (N_8863,N_8130,N_8036);
and U8864 (N_8864,N_8205,N_8168);
and U8865 (N_8865,N_8039,N_8005);
nand U8866 (N_8866,N_8087,N_8242);
nand U8867 (N_8867,N_8400,N_8462);
or U8868 (N_8868,N_8108,N_8351);
nor U8869 (N_8869,N_8034,N_8448);
and U8870 (N_8870,N_8357,N_8278);
or U8871 (N_8871,N_8233,N_8307);
and U8872 (N_8872,N_8319,N_8090);
xor U8873 (N_8873,N_8396,N_8148);
or U8874 (N_8874,N_8443,N_8198);
and U8875 (N_8875,N_8359,N_8074);
or U8876 (N_8876,N_8144,N_8472);
nand U8877 (N_8877,N_8354,N_8105);
and U8878 (N_8878,N_8004,N_8019);
nand U8879 (N_8879,N_8024,N_8156);
nand U8880 (N_8880,N_8114,N_8187);
nand U8881 (N_8881,N_8161,N_8053);
and U8882 (N_8882,N_8129,N_8491);
and U8883 (N_8883,N_8180,N_8037);
nand U8884 (N_8884,N_8386,N_8475);
nand U8885 (N_8885,N_8138,N_8192);
or U8886 (N_8886,N_8345,N_8244);
nor U8887 (N_8887,N_8166,N_8039);
and U8888 (N_8888,N_8202,N_8178);
and U8889 (N_8889,N_8448,N_8411);
and U8890 (N_8890,N_8076,N_8026);
xor U8891 (N_8891,N_8186,N_8083);
nand U8892 (N_8892,N_8192,N_8414);
nor U8893 (N_8893,N_8376,N_8253);
or U8894 (N_8894,N_8300,N_8181);
and U8895 (N_8895,N_8334,N_8420);
or U8896 (N_8896,N_8282,N_8086);
and U8897 (N_8897,N_8431,N_8274);
xnor U8898 (N_8898,N_8082,N_8487);
or U8899 (N_8899,N_8226,N_8335);
and U8900 (N_8900,N_8018,N_8178);
xnor U8901 (N_8901,N_8181,N_8177);
xor U8902 (N_8902,N_8257,N_8146);
or U8903 (N_8903,N_8204,N_8363);
or U8904 (N_8904,N_8297,N_8281);
xor U8905 (N_8905,N_8091,N_8409);
nand U8906 (N_8906,N_8020,N_8496);
nand U8907 (N_8907,N_8137,N_8142);
nand U8908 (N_8908,N_8154,N_8369);
nand U8909 (N_8909,N_8460,N_8414);
nor U8910 (N_8910,N_8083,N_8089);
or U8911 (N_8911,N_8404,N_8239);
nor U8912 (N_8912,N_8190,N_8266);
nor U8913 (N_8913,N_8254,N_8030);
nand U8914 (N_8914,N_8250,N_8434);
and U8915 (N_8915,N_8412,N_8131);
or U8916 (N_8916,N_8063,N_8052);
nand U8917 (N_8917,N_8421,N_8235);
and U8918 (N_8918,N_8002,N_8371);
nor U8919 (N_8919,N_8459,N_8307);
or U8920 (N_8920,N_8471,N_8162);
and U8921 (N_8921,N_8351,N_8413);
or U8922 (N_8922,N_8351,N_8132);
nor U8923 (N_8923,N_8081,N_8389);
and U8924 (N_8924,N_8325,N_8461);
nor U8925 (N_8925,N_8058,N_8438);
nand U8926 (N_8926,N_8034,N_8045);
or U8927 (N_8927,N_8393,N_8168);
xor U8928 (N_8928,N_8470,N_8402);
and U8929 (N_8929,N_8296,N_8129);
xor U8930 (N_8930,N_8332,N_8191);
nand U8931 (N_8931,N_8353,N_8157);
nand U8932 (N_8932,N_8432,N_8131);
nand U8933 (N_8933,N_8116,N_8299);
and U8934 (N_8934,N_8130,N_8161);
or U8935 (N_8935,N_8388,N_8068);
or U8936 (N_8936,N_8448,N_8307);
or U8937 (N_8937,N_8202,N_8362);
and U8938 (N_8938,N_8068,N_8209);
and U8939 (N_8939,N_8307,N_8497);
or U8940 (N_8940,N_8492,N_8092);
or U8941 (N_8941,N_8065,N_8238);
nand U8942 (N_8942,N_8370,N_8389);
and U8943 (N_8943,N_8339,N_8373);
or U8944 (N_8944,N_8135,N_8043);
nand U8945 (N_8945,N_8420,N_8426);
nor U8946 (N_8946,N_8056,N_8256);
nor U8947 (N_8947,N_8426,N_8314);
nand U8948 (N_8948,N_8037,N_8224);
nand U8949 (N_8949,N_8253,N_8121);
nor U8950 (N_8950,N_8497,N_8261);
or U8951 (N_8951,N_8128,N_8197);
nand U8952 (N_8952,N_8394,N_8163);
and U8953 (N_8953,N_8389,N_8325);
or U8954 (N_8954,N_8324,N_8349);
or U8955 (N_8955,N_8083,N_8491);
nand U8956 (N_8956,N_8364,N_8259);
or U8957 (N_8957,N_8130,N_8490);
or U8958 (N_8958,N_8314,N_8116);
and U8959 (N_8959,N_8438,N_8134);
nor U8960 (N_8960,N_8270,N_8430);
or U8961 (N_8961,N_8149,N_8385);
nor U8962 (N_8962,N_8340,N_8191);
nand U8963 (N_8963,N_8498,N_8330);
nand U8964 (N_8964,N_8496,N_8223);
nor U8965 (N_8965,N_8316,N_8319);
xor U8966 (N_8966,N_8183,N_8362);
nand U8967 (N_8967,N_8270,N_8087);
or U8968 (N_8968,N_8393,N_8101);
nor U8969 (N_8969,N_8167,N_8236);
nand U8970 (N_8970,N_8094,N_8230);
and U8971 (N_8971,N_8223,N_8257);
and U8972 (N_8972,N_8000,N_8459);
nand U8973 (N_8973,N_8422,N_8312);
nand U8974 (N_8974,N_8188,N_8381);
or U8975 (N_8975,N_8326,N_8051);
nor U8976 (N_8976,N_8120,N_8134);
nor U8977 (N_8977,N_8052,N_8159);
or U8978 (N_8978,N_8208,N_8084);
and U8979 (N_8979,N_8469,N_8361);
nand U8980 (N_8980,N_8299,N_8229);
nor U8981 (N_8981,N_8296,N_8210);
nor U8982 (N_8982,N_8134,N_8187);
or U8983 (N_8983,N_8207,N_8120);
and U8984 (N_8984,N_8166,N_8350);
or U8985 (N_8985,N_8274,N_8411);
nor U8986 (N_8986,N_8201,N_8108);
or U8987 (N_8987,N_8101,N_8351);
or U8988 (N_8988,N_8439,N_8190);
and U8989 (N_8989,N_8010,N_8050);
nor U8990 (N_8990,N_8335,N_8017);
xor U8991 (N_8991,N_8393,N_8088);
nor U8992 (N_8992,N_8305,N_8487);
xor U8993 (N_8993,N_8219,N_8336);
nor U8994 (N_8994,N_8471,N_8349);
or U8995 (N_8995,N_8073,N_8428);
or U8996 (N_8996,N_8418,N_8117);
nand U8997 (N_8997,N_8000,N_8190);
or U8998 (N_8998,N_8351,N_8010);
or U8999 (N_8999,N_8266,N_8342);
xnor U9000 (N_9000,N_8544,N_8901);
nor U9001 (N_9001,N_8594,N_8591);
and U9002 (N_9002,N_8836,N_8515);
nor U9003 (N_9003,N_8759,N_8932);
nor U9004 (N_9004,N_8774,N_8847);
nor U9005 (N_9005,N_8802,N_8850);
or U9006 (N_9006,N_8589,N_8621);
xor U9007 (N_9007,N_8894,N_8731);
nor U9008 (N_9008,N_8790,N_8839);
nand U9009 (N_9009,N_8912,N_8552);
or U9010 (N_9010,N_8728,N_8587);
xnor U9011 (N_9011,N_8844,N_8871);
nor U9012 (N_9012,N_8739,N_8672);
or U9013 (N_9013,N_8502,N_8596);
nand U9014 (N_9014,N_8954,N_8800);
and U9015 (N_9015,N_8560,N_8978);
or U9016 (N_9016,N_8692,N_8911);
and U9017 (N_9017,N_8971,N_8549);
nand U9018 (N_9018,N_8733,N_8946);
nor U9019 (N_9019,N_8758,N_8631);
and U9020 (N_9020,N_8866,N_8522);
and U9021 (N_9021,N_8547,N_8930);
nor U9022 (N_9022,N_8517,N_8590);
nand U9023 (N_9023,N_8757,N_8961);
nor U9024 (N_9024,N_8712,N_8838);
and U9025 (N_9025,N_8941,N_8753);
or U9026 (N_9026,N_8943,N_8679);
nand U9027 (N_9027,N_8684,N_8663);
and U9028 (N_9028,N_8833,N_8756);
nand U9029 (N_9029,N_8516,N_8632);
or U9030 (N_9030,N_8834,N_8737);
nor U9031 (N_9031,N_8500,N_8769);
and U9032 (N_9032,N_8881,N_8540);
nand U9033 (N_9033,N_8857,N_8593);
or U9034 (N_9034,N_8778,N_8584);
or U9035 (N_9035,N_8695,N_8965);
nor U9036 (N_9036,N_8734,N_8773);
or U9037 (N_9037,N_8597,N_8819);
or U9038 (N_9038,N_8503,N_8822);
nor U9039 (N_9039,N_8874,N_8869);
nand U9040 (N_9040,N_8626,N_8546);
nand U9041 (N_9041,N_8754,N_8750);
nand U9042 (N_9042,N_8524,N_8798);
or U9043 (N_9043,N_8771,N_8969);
and U9044 (N_9044,N_8570,N_8916);
nand U9045 (N_9045,N_8542,N_8519);
nor U9046 (N_9046,N_8891,N_8713);
or U9047 (N_9047,N_8561,N_8801);
nor U9048 (N_9048,N_8666,N_8685);
or U9049 (N_9049,N_8976,N_8554);
nand U9050 (N_9050,N_8831,N_8892);
nor U9051 (N_9051,N_8719,N_8949);
and U9052 (N_9052,N_8856,N_8652);
and U9053 (N_9053,N_8760,N_8691);
and U9054 (N_9054,N_8948,N_8537);
or U9055 (N_9055,N_8812,N_8929);
or U9056 (N_9056,N_8556,N_8922);
nand U9057 (N_9057,N_8867,N_8607);
and U9058 (N_9058,N_8848,N_8842);
xor U9059 (N_9059,N_8803,N_8787);
and U9060 (N_9060,N_8781,N_8643);
nand U9061 (N_9061,N_8751,N_8662);
nor U9062 (N_9062,N_8532,N_8824);
nand U9063 (N_9063,N_8637,N_8531);
nand U9064 (N_9064,N_8588,N_8973);
or U9065 (N_9065,N_8818,N_8989);
and U9066 (N_9066,N_8606,N_8854);
or U9067 (N_9067,N_8676,N_8615);
nand U9068 (N_9068,N_8744,N_8799);
and U9069 (N_9069,N_8680,N_8723);
nand U9070 (N_9070,N_8700,N_8997);
nand U9071 (N_9071,N_8683,N_8986);
nand U9072 (N_9072,N_8791,N_8722);
nor U9073 (N_9073,N_8920,N_8964);
nand U9074 (N_9074,N_8648,N_8727);
and U9075 (N_9075,N_8815,N_8709);
and U9076 (N_9076,N_8772,N_8660);
xnor U9077 (N_9077,N_8828,N_8998);
and U9078 (N_9078,N_8826,N_8938);
xor U9079 (N_9079,N_8855,N_8653);
and U9080 (N_9080,N_8947,N_8592);
nor U9081 (N_9081,N_8706,N_8902);
nor U9082 (N_9082,N_8928,N_8914);
nor U9083 (N_9083,N_8512,N_8821);
and U9084 (N_9084,N_8908,N_8991);
xor U9085 (N_9085,N_8764,N_8707);
nand U9086 (N_9086,N_8553,N_8646);
or U9087 (N_9087,N_8649,N_8956);
nor U9088 (N_9088,N_8619,N_8686);
or U9089 (N_9089,N_8761,N_8795);
and U9090 (N_9090,N_8887,N_8658);
nor U9091 (N_9091,N_8578,N_8749);
and U9092 (N_9092,N_8975,N_8535);
and U9093 (N_9093,N_8521,N_8984);
xor U9094 (N_9094,N_8746,N_8677);
xnor U9095 (N_9095,N_8783,N_8840);
nor U9096 (N_9096,N_8678,N_8858);
xnor U9097 (N_9097,N_8843,N_8513);
nor U9098 (N_9098,N_8609,N_8714);
xor U9099 (N_9099,N_8738,N_8918);
and U9100 (N_9100,N_8952,N_8505);
nor U9101 (N_9101,N_8704,N_8568);
nand U9102 (N_9102,N_8715,N_8823);
nor U9103 (N_9103,N_8852,N_8923);
or U9104 (N_9104,N_8899,N_8527);
or U9105 (N_9105,N_8681,N_8782);
nor U9106 (N_9106,N_8698,N_8897);
nand U9107 (N_9107,N_8917,N_8878);
or U9108 (N_9108,N_8879,N_8766);
and U9109 (N_9109,N_8729,N_8794);
nand U9110 (N_9110,N_8972,N_8741);
or U9111 (N_9111,N_8921,N_8639);
and U9112 (N_9112,N_8555,N_8551);
or U9113 (N_9113,N_8699,N_8618);
xnor U9114 (N_9114,N_8694,N_8886);
nor U9115 (N_9115,N_8518,N_8673);
nor U9116 (N_9116,N_8633,N_8569);
nor U9117 (N_9117,N_8665,N_8508);
and U9118 (N_9118,N_8611,N_8720);
nor U9119 (N_9119,N_8612,N_8813);
or U9120 (N_9120,N_8526,N_8933);
nand U9121 (N_9121,N_8820,N_8579);
and U9122 (N_9122,N_8581,N_8752);
nand U9123 (N_9123,N_8654,N_8784);
nand U9124 (N_9124,N_8939,N_8598);
nor U9125 (N_9125,N_8945,N_8955);
xnor U9126 (N_9126,N_8638,N_8870);
nand U9127 (N_9127,N_8688,N_8862);
xor U9128 (N_9128,N_8661,N_8807);
and U9129 (N_9129,N_8536,N_8634);
nand U9130 (N_9130,N_8924,N_8864);
and U9131 (N_9131,N_8564,N_8559);
nand U9132 (N_9132,N_8725,N_8927);
nand U9133 (N_9133,N_8905,N_8966);
nor U9134 (N_9134,N_8613,N_8806);
nor U9135 (N_9135,N_8573,N_8735);
nand U9136 (N_9136,N_8716,N_8583);
nor U9137 (N_9137,N_8835,N_8804);
nor U9138 (N_9138,N_8523,N_8558);
or U9139 (N_9139,N_8763,N_8792);
and U9140 (N_9140,N_8600,N_8747);
nor U9141 (N_9141,N_8796,N_8814);
or U9142 (N_9142,N_8689,N_8877);
or U9143 (N_9143,N_8900,N_8884);
nor U9144 (N_9144,N_8545,N_8793);
nor U9145 (N_9145,N_8510,N_8825);
and U9146 (N_9146,N_8979,N_8690);
nor U9147 (N_9147,N_8736,N_8853);
nand U9148 (N_9148,N_8687,N_8967);
and U9149 (N_9149,N_8827,N_8616);
or U9150 (N_9150,N_8904,N_8987);
nand U9151 (N_9151,N_8868,N_8996);
and U9152 (N_9152,N_8501,N_8888);
xor U9153 (N_9153,N_8797,N_8861);
nand U9154 (N_9154,N_8624,N_8846);
and U9155 (N_9155,N_8710,N_8935);
nand U9156 (N_9156,N_8701,N_8711);
or U9157 (N_9157,N_8898,N_8717);
nor U9158 (N_9158,N_8651,N_8999);
nor U9159 (N_9159,N_8909,N_8557);
nand U9160 (N_9160,N_8656,N_8608);
and U9161 (N_9161,N_8575,N_8730);
and U9162 (N_9162,N_8628,N_8708);
and U9163 (N_9163,N_8504,N_8983);
nand U9164 (N_9164,N_8768,N_8776);
nand U9165 (N_9165,N_8525,N_8913);
nand U9166 (N_9166,N_8883,N_8697);
and U9167 (N_9167,N_8627,N_8896);
or U9168 (N_9168,N_8577,N_8963);
nor U9169 (N_9169,N_8994,N_8880);
and U9170 (N_9170,N_8860,N_8595);
nand U9171 (N_9171,N_8995,N_8674);
nand U9172 (N_9172,N_8548,N_8944);
nand U9173 (N_9173,N_8657,N_8992);
or U9174 (N_9174,N_8571,N_8957);
and U9175 (N_9175,N_8630,N_8970);
nand U9176 (N_9176,N_8926,N_8507);
xnor U9177 (N_9177,N_8693,N_8780);
and U9178 (N_9178,N_8885,N_8603);
or U9179 (N_9179,N_8958,N_8762);
nand U9180 (N_9180,N_8718,N_8845);
and U9181 (N_9181,N_8876,N_8566);
nor U9182 (N_9182,N_8982,N_8614);
and U9183 (N_9183,N_8936,N_8668);
or U9184 (N_9184,N_8629,N_8988);
xnor U9185 (N_9185,N_8740,N_8703);
and U9186 (N_9186,N_8650,N_8808);
and U9187 (N_9187,N_8779,N_8851);
or U9188 (N_9188,N_8937,N_8533);
and U9189 (N_9189,N_8925,N_8642);
nand U9190 (N_9190,N_8765,N_8514);
nand U9191 (N_9191,N_8742,N_8696);
nand U9192 (N_9192,N_8726,N_8873);
and U9193 (N_9193,N_8530,N_8829);
nand U9194 (N_9194,N_8915,N_8859);
or U9195 (N_9195,N_8528,N_8601);
or U9196 (N_9196,N_8671,N_8636);
or U9197 (N_9197,N_8980,N_8562);
nand U9198 (N_9198,N_8617,N_8786);
nand U9199 (N_9199,N_8610,N_8644);
nand U9200 (N_9200,N_8974,N_8968);
or U9201 (N_9201,N_8940,N_8981);
xor U9202 (N_9202,N_8659,N_8942);
xor U9203 (N_9203,N_8865,N_8959);
nor U9204 (N_9204,N_8931,N_8622);
nand U9205 (N_9205,N_8872,N_8705);
nand U9206 (N_9206,N_8906,N_8599);
and U9207 (N_9207,N_8520,N_8785);
xnor U9208 (N_9208,N_8667,N_8574);
nor U9209 (N_9209,N_8721,N_8805);
or U9210 (N_9210,N_8541,N_8664);
and U9211 (N_9211,N_8849,N_8640);
xnor U9212 (N_9212,N_8645,N_8841);
nand U9213 (N_9213,N_8882,N_8810);
and U9214 (N_9214,N_8724,N_8910);
or U9215 (N_9215,N_8550,N_8511);
or U9216 (N_9216,N_8539,N_8602);
xnor U9217 (N_9217,N_8670,N_8582);
nor U9218 (N_9218,N_8837,N_8748);
nor U9219 (N_9219,N_8506,N_8777);
or U9220 (N_9220,N_8572,N_8565);
and U9221 (N_9221,N_8788,N_8953);
and U9222 (N_9222,N_8903,N_8811);
or U9223 (N_9223,N_8647,N_8985);
or U9224 (N_9224,N_8641,N_8755);
nor U9225 (N_9225,N_8534,N_8604);
and U9226 (N_9226,N_8809,N_8990);
and U9227 (N_9227,N_8775,N_8767);
nand U9228 (N_9228,N_8563,N_8893);
nand U9229 (N_9229,N_8950,N_8605);
and U9230 (N_9230,N_8567,N_8585);
nand U9231 (N_9231,N_8580,N_8509);
and U9232 (N_9232,N_8538,N_8830);
or U9233 (N_9233,N_8586,N_8789);
or U9234 (N_9234,N_8817,N_8702);
nand U9235 (N_9235,N_8655,N_8623);
nor U9236 (N_9236,N_8934,N_8832);
nor U9237 (N_9237,N_8919,N_8977);
and U9238 (N_9238,N_8907,N_8743);
nand U9239 (N_9239,N_8890,N_8895);
nor U9240 (N_9240,N_8962,N_8960);
and U9241 (N_9241,N_8745,N_8951);
or U9242 (N_9242,N_8576,N_8889);
nand U9243 (N_9243,N_8770,N_8875);
nor U9244 (N_9244,N_8625,N_8675);
or U9245 (N_9245,N_8635,N_8816);
xnor U9246 (N_9246,N_8669,N_8543);
and U9247 (N_9247,N_8682,N_8732);
nor U9248 (N_9248,N_8529,N_8863);
and U9249 (N_9249,N_8993,N_8620);
and U9250 (N_9250,N_8664,N_8695);
nor U9251 (N_9251,N_8563,N_8969);
xnor U9252 (N_9252,N_8623,N_8718);
nand U9253 (N_9253,N_8596,N_8581);
or U9254 (N_9254,N_8500,N_8943);
nor U9255 (N_9255,N_8542,N_8778);
nand U9256 (N_9256,N_8572,N_8576);
xor U9257 (N_9257,N_8707,N_8812);
nand U9258 (N_9258,N_8905,N_8775);
and U9259 (N_9259,N_8550,N_8901);
or U9260 (N_9260,N_8755,N_8682);
nand U9261 (N_9261,N_8749,N_8655);
or U9262 (N_9262,N_8891,N_8779);
nand U9263 (N_9263,N_8867,N_8899);
xnor U9264 (N_9264,N_8834,N_8530);
nor U9265 (N_9265,N_8521,N_8824);
nand U9266 (N_9266,N_8883,N_8975);
nand U9267 (N_9267,N_8868,N_8867);
and U9268 (N_9268,N_8834,N_8515);
nor U9269 (N_9269,N_8988,N_8502);
and U9270 (N_9270,N_8872,N_8527);
or U9271 (N_9271,N_8561,N_8752);
and U9272 (N_9272,N_8837,N_8515);
or U9273 (N_9273,N_8582,N_8708);
nand U9274 (N_9274,N_8573,N_8534);
nor U9275 (N_9275,N_8560,N_8843);
nand U9276 (N_9276,N_8722,N_8963);
nand U9277 (N_9277,N_8672,N_8723);
nor U9278 (N_9278,N_8991,N_8543);
or U9279 (N_9279,N_8574,N_8547);
or U9280 (N_9280,N_8848,N_8552);
or U9281 (N_9281,N_8565,N_8897);
nor U9282 (N_9282,N_8913,N_8602);
or U9283 (N_9283,N_8906,N_8577);
nand U9284 (N_9284,N_8944,N_8852);
xor U9285 (N_9285,N_8992,N_8521);
and U9286 (N_9286,N_8782,N_8989);
and U9287 (N_9287,N_8705,N_8711);
nand U9288 (N_9288,N_8769,N_8937);
xor U9289 (N_9289,N_8593,N_8976);
nand U9290 (N_9290,N_8767,N_8957);
or U9291 (N_9291,N_8749,N_8524);
nand U9292 (N_9292,N_8884,N_8579);
or U9293 (N_9293,N_8513,N_8621);
nand U9294 (N_9294,N_8767,N_8872);
nor U9295 (N_9295,N_8607,N_8600);
nor U9296 (N_9296,N_8659,N_8925);
nand U9297 (N_9297,N_8516,N_8750);
xnor U9298 (N_9298,N_8642,N_8969);
nand U9299 (N_9299,N_8507,N_8859);
nand U9300 (N_9300,N_8926,N_8867);
and U9301 (N_9301,N_8746,N_8789);
nor U9302 (N_9302,N_8806,N_8855);
and U9303 (N_9303,N_8581,N_8790);
and U9304 (N_9304,N_8791,N_8915);
xor U9305 (N_9305,N_8675,N_8746);
and U9306 (N_9306,N_8676,N_8822);
and U9307 (N_9307,N_8548,N_8621);
and U9308 (N_9308,N_8669,N_8576);
or U9309 (N_9309,N_8746,N_8991);
nand U9310 (N_9310,N_8881,N_8792);
xnor U9311 (N_9311,N_8736,N_8804);
or U9312 (N_9312,N_8670,N_8715);
nand U9313 (N_9313,N_8541,N_8923);
nand U9314 (N_9314,N_8850,N_8528);
nor U9315 (N_9315,N_8903,N_8819);
and U9316 (N_9316,N_8852,N_8639);
and U9317 (N_9317,N_8688,N_8820);
or U9318 (N_9318,N_8766,N_8752);
nor U9319 (N_9319,N_8708,N_8851);
and U9320 (N_9320,N_8708,N_8834);
and U9321 (N_9321,N_8817,N_8938);
nor U9322 (N_9322,N_8725,N_8971);
xor U9323 (N_9323,N_8735,N_8545);
or U9324 (N_9324,N_8763,N_8625);
or U9325 (N_9325,N_8570,N_8885);
xnor U9326 (N_9326,N_8818,N_8769);
xor U9327 (N_9327,N_8971,N_8885);
nor U9328 (N_9328,N_8713,N_8931);
and U9329 (N_9329,N_8712,N_8569);
nor U9330 (N_9330,N_8504,N_8634);
or U9331 (N_9331,N_8594,N_8656);
nand U9332 (N_9332,N_8863,N_8984);
xor U9333 (N_9333,N_8870,N_8794);
nor U9334 (N_9334,N_8541,N_8846);
nor U9335 (N_9335,N_8816,N_8905);
or U9336 (N_9336,N_8754,N_8764);
and U9337 (N_9337,N_8962,N_8869);
xor U9338 (N_9338,N_8565,N_8788);
xor U9339 (N_9339,N_8760,N_8756);
or U9340 (N_9340,N_8626,N_8551);
and U9341 (N_9341,N_8924,N_8513);
and U9342 (N_9342,N_8888,N_8620);
nand U9343 (N_9343,N_8962,N_8947);
nand U9344 (N_9344,N_8896,N_8930);
xor U9345 (N_9345,N_8506,N_8921);
nor U9346 (N_9346,N_8908,N_8818);
xor U9347 (N_9347,N_8503,N_8602);
and U9348 (N_9348,N_8739,N_8766);
or U9349 (N_9349,N_8765,N_8802);
nand U9350 (N_9350,N_8767,N_8709);
or U9351 (N_9351,N_8764,N_8914);
nand U9352 (N_9352,N_8664,N_8739);
nor U9353 (N_9353,N_8709,N_8913);
and U9354 (N_9354,N_8593,N_8594);
nand U9355 (N_9355,N_8855,N_8717);
and U9356 (N_9356,N_8813,N_8851);
or U9357 (N_9357,N_8559,N_8705);
or U9358 (N_9358,N_8838,N_8807);
or U9359 (N_9359,N_8798,N_8938);
or U9360 (N_9360,N_8668,N_8827);
xnor U9361 (N_9361,N_8952,N_8689);
nand U9362 (N_9362,N_8889,N_8675);
xor U9363 (N_9363,N_8845,N_8795);
and U9364 (N_9364,N_8607,N_8771);
nand U9365 (N_9365,N_8546,N_8699);
nor U9366 (N_9366,N_8758,N_8529);
or U9367 (N_9367,N_8539,N_8695);
nand U9368 (N_9368,N_8840,N_8785);
nor U9369 (N_9369,N_8621,N_8777);
nor U9370 (N_9370,N_8751,N_8618);
nor U9371 (N_9371,N_8530,N_8696);
nand U9372 (N_9372,N_8724,N_8812);
nand U9373 (N_9373,N_8756,N_8745);
and U9374 (N_9374,N_8720,N_8895);
nand U9375 (N_9375,N_8946,N_8746);
and U9376 (N_9376,N_8815,N_8895);
xnor U9377 (N_9377,N_8695,N_8923);
nor U9378 (N_9378,N_8518,N_8613);
or U9379 (N_9379,N_8752,N_8606);
xnor U9380 (N_9380,N_8556,N_8713);
and U9381 (N_9381,N_8783,N_8944);
xor U9382 (N_9382,N_8958,N_8502);
or U9383 (N_9383,N_8509,N_8860);
nor U9384 (N_9384,N_8640,N_8870);
and U9385 (N_9385,N_8843,N_8569);
nor U9386 (N_9386,N_8521,N_8529);
and U9387 (N_9387,N_8841,N_8847);
nor U9388 (N_9388,N_8769,N_8870);
nor U9389 (N_9389,N_8565,N_8632);
and U9390 (N_9390,N_8871,N_8721);
xor U9391 (N_9391,N_8754,N_8596);
nor U9392 (N_9392,N_8836,N_8830);
xor U9393 (N_9393,N_8906,N_8892);
and U9394 (N_9394,N_8681,N_8884);
nand U9395 (N_9395,N_8554,N_8773);
nand U9396 (N_9396,N_8822,N_8623);
nor U9397 (N_9397,N_8915,N_8780);
nand U9398 (N_9398,N_8954,N_8709);
or U9399 (N_9399,N_8765,N_8553);
nand U9400 (N_9400,N_8669,N_8662);
and U9401 (N_9401,N_8650,N_8641);
nor U9402 (N_9402,N_8533,N_8808);
xor U9403 (N_9403,N_8572,N_8923);
nor U9404 (N_9404,N_8715,N_8910);
or U9405 (N_9405,N_8890,N_8766);
or U9406 (N_9406,N_8594,N_8953);
nand U9407 (N_9407,N_8772,N_8715);
or U9408 (N_9408,N_8595,N_8554);
and U9409 (N_9409,N_8955,N_8969);
nor U9410 (N_9410,N_8611,N_8779);
nand U9411 (N_9411,N_8741,N_8968);
or U9412 (N_9412,N_8642,N_8615);
xnor U9413 (N_9413,N_8970,N_8760);
or U9414 (N_9414,N_8971,N_8537);
nand U9415 (N_9415,N_8703,N_8581);
xor U9416 (N_9416,N_8845,N_8837);
and U9417 (N_9417,N_8843,N_8594);
xnor U9418 (N_9418,N_8619,N_8530);
or U9419 (N_9419,N_8776,N_8509);
nor U9420 (N_9420,N_8906,N_8788);
or U9421 (N_9421,N_8567,N_8631);
nor U9422 (N_9422,N_8556,N_8589);
nand U9423 (N_9423,N_8759,N_8990);
and U9424 (N_9424,N_8732,N_8870);
nor U9425 (N_9425,N_8851,N_8591);
nor U9426 (N_9426,N_8708,N_8903);
and U9427 (N_9427,N_8523,N_8741);
nor U9428 (N_9428,N_8775,N_8845);
and U9429 (N_9429,N_8915,N_8895);
and U9430 (N_9430,N_8786,N_8843);
or U9431 (N_9431,N_8928,N_8523);
nor U9432 (N_9432,N_8855,N_8638);
xnor U9433 (N_9433,N_8969,N_8570);
nand U9434 (N_9434,N_8887,N_8500);
or U9435 (N_9435,N_8844,N_8512);
or U9436 (N_9436,N_8852,N_8620);
or U9437 (N_9437,N_8966,N_8672);
or U9438 (N_9438,N_8828,N_8825);
nand U9439 (N_9439,N_8758,N_8512);
or U9440 (N_9440,N_8687,N_8864);
and U9441 (N_9441,N_8690,N_8654);
or U9442 (N_9442,N_8689,N_8680);
nor U9443 (N_9443,N_8746,N_8797);
or U9444 (N_9444,N_8560,N_8798);
xnor U9445 (N_9445,N_8816,N_8888);
or U9446 (N_9446,N_8698,N_8935);
or U9447 (N_9447,N_8653,N_8805);
or U9448 (N_9448,N_8840,N_8505);
or U9449 (N_9449,N_8765,N_8650);
and U9450 (N_9450,N_8508,N_8700);
xor U9451 (N_9451,N_8896,N_8656);
nand U9452 (N_9452,N_8560,N_8864);
or U9453 (N_9453,N_8500,N_8715);
or U9454 (N_9454,N_8912,N_8969);
nand U9455 (N_9455,N_8682,N_8821);
xor U9456 (N_9456,N_8545,N_8866);
nor U9457 (N_9457,N_8775,N_8977);
nor U9458 (N_9458,N_8657,N_8928);
xnor U9459 (N_9459,N_8703,N_8682);
nor U9460 (N_9460,N_8686,N_8946);
and U9461 (N_9461,N_8541,N_8523);
xor U9462 (N_9462,N_8618,N_8776);
or U9463 (N_9463,N_8686,N_8632);
or U9464 (N_9464,N_8811,N_8905);
nand U9465 (N_9465,N_8803,N_8874);
nor U9466 (N_9466,N_8644,N_8796);
xor U9467 (N_9467,N_8667,N_8522);
nand U9468 (N_9468,N_8799,N_8662);
nand U9469 (N_9469,N_8729,N_8784);
xnor U9470 (N_9470,N_8577,N_8804);
and U9471 (N_9471,N_8515,N_8810);
nand U9472 (N_9472,N_8887,N_8801);
nand U9473 (N_9473,N_8791,N_8873);
or U9474 (N_9474,N_8892,N_8822);
nand U9475 (N_9475,N_8813,N_8658);
or U9476 (N_9476,N_8700,N_8954);
and U9477 (N_9477,N_8979,N_8995);
nand U9478 (N_9478,N_8907,N_8768);
and U9479 (N_9479,N_8781,N_8658);
and U9480 (N_9480,N_8643,N_8650);
nor U9481 (N_9481,N_8620,N_8847);
nor U9482 (N_9482,N_8769,N_8839);
or U9483 (N_9483,N_8706,N_8860);
nand U9484 (N_9484,N_8851,N_8558);
nand U9485 (N_9485,N_8767,N_8620);
and U9486 (N_9486,N_8907,N_8562);
xnor U9487 (N_9487,N_8658,N_8528);
nor U9488 (N_9488,N_8670,N_8737);
nand U9489 (N_9489,N_8831,N_8928);
nand U9490 (N_9490,N_8547,N_8761);
nor U9491 (N_9491,N_8679,N_8586);
nor U9492 (N_9492,N_8616,N_8961);
and U9493 (N_9493,N_8620,N_8682);
nand U9494 (N_9494,N_8864,N_8941);
nor U9495 (N_9495,N_8976,N_8745);
or U9496 (N_9496,N_8793,N_8558);
nand U9497 (N_9497,N_8703,N_8763);
nand U9498 (N_9498,N_8666,N_8889);
nand U9499 (N_9499,N_8775,N_8619);
nor U9500 (N_9500,N_9424,N_9322);
nor U9501 (N_9501,N_9149,N_9387);
and U9502 (N_9502,N_9276,N_9338);
nand U9503 (N_9503,N_9079,N_9174);
or U9504 (N_9504,N_9358,N_9319);
or U9505 (N_9505,N_9126,N_9313);
and U9506 (N_9506,N_9056,N_9105);
and U9507 (N_9507,N_9172,N_9396);
nor U9508 (N_9508,N_9188,N_9478);
and U9509 (N_9509,N_9164,N_9234);
nor U9510 (N_9510,N_9167,N_9066);
and U9511 (N_9511,N_9236,N_9349);
nor U9512 (N_9512,N_9406,N_9481);
and U9513 (N_9513,N_9493,N_9185);
xor U9514 (N_9514,N_9088,N_9299);
nand U9515 (N_9515,N_9013,N_9046);
and U9516 (N_9516,N_9000,N_9304);
nand U9517 (N_9517,N_9118,N_9180);
nor U9518 (N_9518,N_9353,N_9489);
nor U9519 (N_9519,N_9280,N_9003);
and U9520 (N_9520,N_9421,N_9197);
nand U9521 (N_9521,N_9354,N_9246);
or U9522 (N_9522,N_9433,N_9265);
and U9523 (N_9523,N_9277,N_9183);
or U9524 (N_9524,N_9070,N_9207);
or U9525 (N_9525,N_9272,N_9331);
or U9526 (N_9526,N_9028,N_9286);
xor U9527 (N_9527,N_9098,N_9275);
nand U9528 (N_9528,N_9315,N_9057);
and U9529 (N_9529,N_9374,N_9243);
nand U9530 (N_9530,N_9371,N_9366);
and U9531 (N_9531,N_9259,N_9208);
or U9532 (N_9532,N_9125,N_9404);
nor U9533 (N_9533,N_9038,N_9093);
nor U9534 (N_9534,N_9170,N_9081);
or U9535 (N_9535,N_9018,N_9453);
and U9536 (N_9536,N_9006,N_9309);
nor U9537 (N_9537,N_9449,N_9410);
nor U9538 (N_9538,N_9177,N_9488);
and U9539 (N_9539,N_9251,N_9369);
nor U9540 (N_9540,N_9378,N_9132);
and U9541 (N_9541,N_9184,N_9089);
or U9542 (N_9542,N_9201,N_9362);
or U9543 (N_9543,N_9162,N_9026);
nor U9544 (N_9544,N_9456,N_9323);
nand U9545 (N_9545,N_9150,N_9249);
or U9546 (N_9546,N_9023,N_9037);
nor U9547 (N_9547,N_9182,N_9465);
and U9548 (N_9548,N_9128,N_9096);
nand U9549 (N_9549,N_9082,N_9446);
nor U9550 (N_9550,N_9332,N_9291);
and U9551 (N_9551,N_9289,N_9022);
and U9552 (N_9552,N_9194,N_9255);
and U9553 (N_9553,N_9067,N_9068);
nand U9554 (N_9554,N_9240,N_9448);
nor U9555 (N_9555,N_9241,N_9014);
nand U9556 (N_9556,N_9395,N_9140);
or U9557 (N_9557,N_9175,N_9392);
and U9558 (N_9558,N_9407,N_9209);
nand U9559 (N_9559,N_9334,N_9494);
and U9560 (N_9560,N_9238,N_9035);
nor U9561 (N_9561,N_9095,N_9031);
nor U9562 (N_9562,N_9033,N_9300);
nor U9563 (N_9563,N_9254,N_9024);
or U9564 (N_9564,N_9273,N_9475);
nor U9565 (N_9565,N_9131,N_9482);
and U9566 (N_9566,N_9283,N_9034);
nand U9567 (N_9567,N_9411,N_9141);
nor U9568 (N_9568,N_9110,N_9186);
xnor U9569 (N_9569,N_9080,N_9191);
nor U9570 (N_9570,N_9414,N_9495);
nand U9571 (N_9571,N_9460,N_9069);
nand U9572 (N_9572,N_9491,N_9450);
or U9573 (N_9573,N_9200,N_9156);
or U9574 (N_9574,N_9356,N_9423);
xnor U9575 (N_9575,N_9308,N_9106);
xnor U9576 (N_9576,N_9157,N_9333);
nand U9577 (N_9577,N_9377,N_9152);
or U9578 (N_9578,N_9444,N_9245);
nand U9579 (N_9579,N_9373,N_9107);
nand U9580 (N_9580,N_9094,N_9496);
or U9581 (N_9581,N_9384,N_9393);
xnor U9582 (N_9582,N_9466,N_9270);
or U9583 (N_9583,N_9434,N_9441);
xor U9584 (N_9584,N_9459,N_9016);
or U9585 (N_9585,N_9004,N_9136);
nand U9586 (N_9586,N_9168,N_9085);
and U9587 (N_9587,N_9281,N_9400);
nor U9588 (N_9588,N_9160,N_9363);
or U9589 (N_9589,N_9403,N_9497);
nor U9590 (N_9590,N_9102,N_9399);
or U9591 (N_9591,N_9159,N_9357);
nor U9592 (N_9592,N_9445,N_9019);
and U9593 (N_9593,N_9415,N_9100);
xor U9594 (N_9594,N_9116,N_9282);
nand U9595 (N_9595,N_9134,N_9065);
nand U9596 (N_9596,N_9361,N_9454);
nor U9597 (N_9597,N_9213,N_9228);
or U9598 (N_9598,N_9268,N_9101);
nor U9599 (N_9599,N_9327,N_9347);
and U9600 (N_9600,N_9412,N_9295);
or U9601 (N_9601,N_9340,N_9408);
or U9602 (N_9602,N_9051,N_9321);
nor U9603 (N_9603,N_9360,N_9311);
nand U9604 (N_9604,N_9429,N_9165);
nand U9605 (N_9605,N_9196,N_9122);
or U9606 (N_9606,N_9325,N_9344);
nand U9607 (N_9607,N_9485,N_9279);
and U9608 (N_9608,N_9062,N_9244);
nand U9609 (N_9609,N_9405,N_9350);
or U9610 (N_9610,N_9169,N_9119);
or U9611 (N_9611,N_9090,N_9012);
nand U9612 (N_9612,N_9058,N_9301);
xor U9613 (N_9613,N_9047,N_9452);
xor U9614 (N_9614,N_9135,N_9432);
xnor U9615 (N_9615,N_9237,N_9198);
nand U9616 (N_9616,N_9111,N_9040);
and U9617 (N_9617,N_9455,N_9469);
xnor U9618 (N_9618,N_9148,N_9044);
and U9619 (N_9619,N_9355,N_9231);
nand U9620 (N_9620,N_9263,N_9179);
nand U9621 (N_9621,N_9235,N_9413);
nand U9622 (N_9622,N_9464,N_9375);
and U9623 (N_9623,N_9316,N_9473);
nor U9624 (N_9624,N_9064,N_9389);
and U9625 (N_9625,N_9425,N_9351);
and U9626 (N_9626,N_9206,N_9269);
or U9627 (N_9627,N_9250,N_9345);
nand U9628 (N_9628,N_9042,N_9161);
or U9629 (N_9629,N_9457,N_9226);
or U9630 (N_9630,N_9470,N_9290);
or U9631 (N_9631,N_9383,N_9010);
nor U9632 (N_9632,N_9216,N_9428);
nor U9633 (N_9633,N_9054,N_9123);
xnor U9634 (N_9634,N_9438,N_9391);
nor U9635 (N_9635,N_9242,N_9124);
and U9636 (N_9636,N_9143,N_9002);
nand U9637 (N_9637,N_9144,N_9227);
or U9638 (N_9638,N_9223,N_9121);
nor U9639 (N_9639,N_9097,N_9092);
nor U9640 (N_9640,N_9009,N_9086);
nand U9641 (N_9641,N_9490,N_9352);
xor U9642 (N_9642,N_9139,N_9048);
nor U9643 (N_9643,N_9147,N_9137);
nand U9644 (N_9644,N_9442,N_9229);
nor U9645 (N_9645,N_9380,N_9402);
and U9646 (N_9646,N_9278,N_9176);
or U9647 (N_9647,N_9303,N_9030);
nor U9648 (N_9648,N_9328,N_9181);
and U9649 (N_9649,N_9193,N_9153);
or U9650 (N_9650,N_9341,N_9215);
nand U9651 (N_9651,N_9114,N_9379);
and U9652 (N_9652,N_9027,N_9293);
nand U9653 (N_9653,N_9307,N_9078);
and U9654 (N_9654,N_9133,N_9072);
xnor U9655 (N_9655,N_9113,N_9376);
nor U9656 (N_9656,N_9025,N_9173);
nor U9657 (N_9657,N_9075,N_9049);
nand U9658 (N_9658,N_9032,N_9195);
xor U9659 (N_9659,N_9440,N_9348);
or U9660 (N_9660,N_9084,N_9339);
and U9661 (N_9661,N_9431,N_9330);
or U9662 (N_9662,N_9427,N_9318);
or U9663 (N_9663,N_9008,N_9492);
nand U9664 (N_9664,N_9274,N_9294);
nor U9665 (N_9665,N_9346,N_9073);
nand U9666 (N_9666,N_9011,N_9053);
nand U9667 (N_9667,N_9225,N_9061);
and U9668 (N_9668,N_9288,N_9120);
or U9669 (N_9669,N_9214,N_9480);
nand U9670 (N_9670,N_9007,N_9462);
nand U9671 (N_9671,N_9261,N_9296);
and U9672 (N_9672,N_9484,N_9359);
or U9673 (N_9673,N_9381,N_9262);
nand U9674 (N_9674,N_9409,N_9076);
or U9675 (N_9675,N_9386,N_9258);
nor U9676 (N_9676,N_9217,N_9043);
and U9677 (N_9677,N_9219,N_9397);
nand U9678 (N_9678,N_9052,N_9055);
nand U9679 (N_9679,N_9189,N_9230);
and U9680 (N_9680,N_9474,N_9285);
and U9681 (N_9681,N_9050,N_9302);
or U9682 (N_9682,N_9256,N_9320);
or U9683 (N_9683,N_9416,N_9297);
and U9684 (N_9684,N_9127,N_9142);
or U9685 (N_9685,N_9109,N_9239);
nand U9686 (N_9686,N_9232,N_9021);
or U9687 (N_9687,N_9151,N_9368);
nand U9688 (N_9688,N_9247,N_9264);
or U9689 (N_9689,N_9099,N_9398);
nor U9690 (N_9690,N_9337,N_9103);
and U9691 (N_9691,N_9372,N_9401);
xnor U9692 (N_9692,N_9166,N_9171);
nor U9693 (N_9693,N_9267,N_9390);
or U9694 (N_9694,N_9417,N_9312);
or U9695 (N_9695,N_9483,N_9467);
or U9696 (N_9696,N_9104,N_9146);
nand U9697 (N_9697,N_9222,N_9001);
nor U9698 (N_9698,N_9203,N_9451);
nand U9699 (N_9699,N_9463,N_9310);
and U9700 (N_9700,N_9115,N_9447);
and U9701 (N_9701,N_9045,N_9422);
nor U9702 (N_9702,N_9477,N_9343);
nor U9703 (N_9703,N_9498,N_9336);
nand U9704 (N_9704,N_9471,N_9430);
or U9705 (N_9705,N_9439,N_9419);
nand U9706 (N_9706,N_9029,N_9365);
or U9707 (N_9707,N_9020,N_9117);
nor U9708 (N_9708,N_9314,N_9071);
nor U9709 (N_9709,N_9087,N_9298);
xor U9710 (N_9710,N_9145,N_9252);
nor U9711 (N_9711,N_9017,N_9284);
or U9712 (N_9712,N_9317,N_9248);
or U9713 (N_9713,N_9158,N_9108);
nor U9714 (N_9714,N_9260,N_9305);
or U9715 (N_9715,N_9130,N_9199);
and U9716 (N_9716,N_9155,N_9039);
or U9717 (N_9717,N_9487,N_9212);
nand U9718 (N_9718,N_9205,N_9192);
nand U9719 (N_9719,N_9202,N_9479);
nand U9720 (N_9720,N_9015,N_9426);
nand U9721 (N_9721,N_9435,N_9233);
nor U9722 (N_9722,N_9499,N_9436);
or U9723 (N_9723,N_9370,N_9324);
nand U9724 (N_9724,N_9394,N_9091);
nand U9725 (N_9725,N_9224,N_9129);
or U9726 (N_9726,N_9083,N_9138);
and U9727 (N_9727,N_9163,N_9266);
and U9728 (N_9728,N_9154,N_9178);
nor U9729 (N_9729,N_9437,N_9041);
or U9730 (N_9730,N_9486,N_9077);
nor U9731 (N_9731,N_9221,N_9210);
or U9732 (N_9732,N_9306,N_9220);
and U9733 (N_9733,N_9187,N_9476);
nor U9734 (N_9734,N_9074,N_9257);
nor U9735 (N_9735,N_9063,N_9458);
xor U9736 (N_9736,N_9059,N_9253);
nor U9737 (N_9737,N_9005,N_9385);
nor U9738 (N_9738,N_9461,N_9287);
and U9739 (N_9739,N_9190,N_9060);
or U9740 (N_9740,N_9204,N_9420);
xnor U9741 (N_9741,N_9364,N_9418);
and U9742 (N_9742,N_9292,N_9388);
nor U9743 (N_9743,N_9382,N_9326);
nand U9744 (N_9744,N_9335,N_9271);
or U9745 (N_9745,N_9036,N_9443);
nor U9746 (N_9746,N_9329,N_9367);
nor U9747 (N_9747,N_9342,N_9468);
nor U9748 (N_9748,N_9211,N_9472);
xnor U9749 (N_9749,N_9112,N_9218);
nand U9750 (N_9750,N_9297,N_9043);
nand U9751 (N_9751,N_9344,N_9073);
nand U9752 (N_9752,N_9372,N_9010);
nand U9753 (N_9753,N_9312,N_9437);
nor U9754 (N_9754,N_9429,N_9135);
and U9755 (N_9755,N_9080,N_9290);
nand U9756 (N_9756,N_9186,N_9332);
nand U9757 (N_9757,N_9353,N_9254);
nor U9758 (N_9758,N_9104,N_9026);
nand U9759 (N_9759,N_9296,N_9055);
nor U9760 (N_9760,N_9072,N_9019);
nand U9761 (N_9761,N_9075,N_9320);
or U9762 (N_9762,N_9025,N_9455);
or U9763 (N_9763,N_9466,N_9424);
nand U9764 (N_9764,N_9218,N_9488);
nor U9765 (N_9765,N_9483,N_9052);
nand U9766 (N_9766,N_9398,N_9078);
or U9767 (N_9767,N_9433,N_9228);
nor U9768 (N_9768,N_9256,N_9362);
and U9769 (N_9769,N_9130,N_9261);
and U9770 (N_9770,N_9184,N_9314);
nor U9771 (N_9771,N_9366,N_9368);
or U9772 (N_9772,N_9477,N_9287);
nand U9773 (N_9773,N_9374,N_9018);
xnor U9774 (N_9774,N_9377,N_9064);
nand U9775 (N_9775,N_9159,N_9337);
or U9776 (N_9776,N_9348,N_9096);
or U9777 (N_9777,N_9123,N_9029);
nand U9778 (N_9778,N_9215,N_9163);
xnor U9779 (N_9779,N_9210,N_9218);
nand U9780 (N_9780,N_9300,N_9140);
or U9781 (N_9781,N_9312,N_9457);
nand U9782 (N_9782,N_9399,N_9212);
nand U9783 (N_9783,N_9275,N_9465);
and U9784 (N_9784,N_9317,N_9275);
nor U9785 (N_9785,N_9340,N_9417);
nor U9786 (N_9786,N_9185,N_9478);
and U9787 (N_9787,N_9061,N_9484);
nand U9788 (N_9788,N_9076,N_9419);
nand U9789 (N_9789,N_9429,N_9244);
nor U9790 (N_9790,N_9373,N_9051);
nand U9791 (N_9791,N_9307,N_9090);
xnor U9792 (N_9792,N_9492,N_9305);
and U9793 (N_9793,N_9340,N_9262);
nor U9794 (N_9794,N_9427,N_9479);
nand U9795 (N_9795,N_9224,N_9200);
or U9796 (N_9796,N_9108,N_9498);
or U9797 (N_9797,N_9028,N_9199);
xor U9798 (N_9798,N_9367,N_9120);
nand U9799 (N_9799,N_9466,N_9445);
nand U9800 (N_9800,N_9476,N_9021);
nor U9801 (N_9801,N_9091,N_9336);
or U9802 (N_9802,N_9012,N_9149);
xor U9803 (N_9803,N_9187,N_9207);
nor U9804 (N_9804,N_9289,N_9444);
nand U9805 (N_9805,N_9041,N_9078);
nand U9806 (N_9806,N_9202,N_9048);
and U9807 (N_9807,N_9103,N_9402);
nor U9808 (N_9808,N_9111,N_9062);
or U9809 (N_9809,N_9131,N_9165);
or U9810 (N_9810,N_9111,N_9023);
nand U9811 (N_9811,N_9396,N_9069);
nand U9812 (N_9812,N_9248,N_9138);
nor U9813 (N_9813,N_9003,N_9277);
nand U9814 (N_9814,N_9177,N_9011);
and U9815 (N_9815,N_9261,N_9001);
and U9816 (N_9816,N_9476,N_9036);
nand U9817 (N_9817,N_9163,N_9288);
and U9818 (N_9818,N_9239,N_9310);
or U9819 (N_9819,N_9228,N_9327);
and U9820 (N_9820,N_9036,N_9253);
and U9821 (N_9821,N_9128,N_9064);
nand U9822 (N_9822,N_9351,N_9167);
nand U9823 (N_9823,N_9285,N_9363);
xnor U9824 (N_9824,N_9236,N_9134);
nor U9825 (N_9825,N_9449,N_9232);
or U9826 (N_9826,N_9194,N_9372);
nor U9827 (N_9827,N_9196,N_9247);
nand U9828 (N_9828,N_9322,N_9106);
xnor U9829 (N_9829,N_9358,N_9300);
nor U9830 (N_9830,N_9435,N_9110);
or U9831 (N_9831,N_9274,N_9024);
nand U9832 (N_9832,N_9474,N_9422);
xor U9833 (N_9833,N_9196,N_9069);
or U9834 (N_9834,N_9430,N_9284);
xnor U9835 (N_9835,N_9266,N_9039);
nand U9836 (N_9836,N_9067,N_9234);
xor U9837 (N_9837,N_9496,N_9133);
nor U9838 (N_9838,N_9127,N_9311);
nor U9839 (N_9839,N_9328,N_9241);
xnor U9840 (N_9840,N_9412,N_9235);
and U9841 (N_9841,N_9314,N_9425);
or U9842 (N_9842,N_9109,N_9324);
nand U9843 (N_9843,N_9072,N_9163);
or U9844 (N_9844,N_9439,N_9084);
xor U9845 (N_9845,N_9305,N_9468);
xor U9846 (N_9846,N_9375,N_9196);
and U9847 (N_9847,N_9475,N_9126);
nor U9848 (N_9848,N_9257,N_9174);
xor U9849 (N_9849,N_9369,N_9002);
and U9850 (N_9850,N_9263,N_9065);
nor U9851 (N_9851,N_9079,N_9450);
or U9852 (N_9852,N_9141,N_9039);
and U9853 (N_9853,N_9159,N_9483);
or U9854 (N_9854,N_9270,N_9101);
nor U9855 (N_9855,N_9070,N_9480);
or U9856 (N_9856,N_9064,N_9304);
xor U9857 (N_9857,N_9254,N_9056);
or U9858 (N_9858,N_9254,N_9119);
nand U9859 (N_9859,N_9484,N_9429);
nand U9860 (N_9860,N_9303,N_9184);
nor U9861 (N_9861,N_9217,N_9464);
or U9862 (N_9862,N_9241,N_9194);
nor U9863 (N_9863,N_9393,N_9330);
nor U9864 (N_9864,N_9497,N_9239);
nand U9865 (N_9865,N_9175,N_9322);
or U9866 (N_9866,N_9100,N_9288);
nor U9867 (N_9867,N_9195,N_9303);
and U9868 (N_9868,N_9347,N_9216);
nand U9869 (N_9869,N_9364,N_9053);
and U9870 (N_9870,N_9229,N_9279);
or U9871 (N_9871,N_9406,N_9165);
nor U9872 (N_9872,N_9377,N_9199);
or U9873 (N_9873,N_9405,N_9355);
or U9874 (N_9874,N_9290,N_9196);
nor U9875 (N_9875,N_9244,N_9311);
and U9876 (N_9876,N_9472,N_9131);
xor U9877 (N_9877,N_9127,N_9145);
nor U9878 (N_9878,N_9018,N_9479);
xor U9879 (N_9879,N_9178,N_9276);
or U9880 (N_9880,N_9131,N_9092);
nand U9881 (N_9881,N_9303,N_9226);
nor U9882 (N_9882,N_9091,N_9274);
and U9883 (N_9883,N_9365,N_9448);
nand U9884 (N_9884,N_9498,N_9280);
or U9885 (N_9885,N_9116,N_9334);
nand U9886 (N_9886,N_9453,N_9102);
nand U9887 (N_9887,N_9176,N_9133);
nor U9888 (N_9888,N_9217,N_9099);
xor U9889 (N_9889,N_9348,N_9397);
nand U9890 (N_9890,N_9016,N_9390);
or U9891 (N_9891,N_9423,N_9057);
or U9892 (N_9892,N_9016,N_9406);
nand U9893 (N_9893,N_9298,N_9419);
and U9894 (N_9894,N_9446,N_9333);
nand U9895 (N_9895,N_9251,N_9054);
or U9896 (N_9896,N_9411,N_9294);
or U9897 (N_9897,N_9400,N_9325);
nor U9898 (N_9898,N_9395,N_9447);
nand U9899 (N_9899,N_9185,N_9370);
nor U9900 (N_9900,N_9199,N_9163);
nand U9901 (N_9901,N_9070,N_9201);
or U9902 (N_9902,N_9028,N_9448);
or U9903 (N_9903,N_9250,N_9160);
or U9904 (N_9904,N_9385,N_9127);
nor U9905 (N_9905,N_9085,N_9486);
and U9906 (N_9906,N_9161,N_9476);
nor U9907 (N_9907,N_9439,N_9440);
nor U9908 (N_9908,N_9394,N_9125);
xnor U9909 (N_9909,N_9294,N_9163);
xnor U9910 (N_9910,N_9178,N_9374);
or U9911 (N_9911,N_9474,N_9300);
nand U9912 (N_9912,N_9334,N_9193);
nor U9913 (N_9913,N_9449,N_9377);
nand U9914 (N_9914,N_9037,N_9246);
nor U9915 (N_9915,N_9336,N_9180);
and U9916 (N_9916,N_9285,N_9186);
nor U9917 (N_9917,N_9422,N_9285);
nor U9918 (N_9918,N_9314,N_9010);
or U9919 (N_9919,N_9294,N_9030);
nand U9920 (N_9920,N_9387,N_9378);
nor U9921 (N_9921,N_9326,N_9202);
nor U9922 (N_9922,N_9284,N_9249);
or U9923 (N_9923,N_9467,N_9144);
or U9924 (N_9924,N_9151,N_9445);
nor U9925 (N_9925,N_9193,N_9307);
nor U9926 (N_9926,N_9173,N_9022);
nand U9927 (N_9927,N_9261,N_9377);
or U9928 (N_9928,N_9018,N_9244);
or U9929 (N_9929,N_9347,N_9122);
nand U9930 (N_9930,N_9074,N_9390);
or U9931 (N_9931,N_9476,N_9258);
nor U9932 (N_9932,N_9337,N_9369);
and U9933 (N_9933,N_9442,N_9349);
or U9934 (N_9934,N_9003,N_9276);
nand U9935 (N_9935,N_9449,N_9009);
and U9936 (N_9936,N_9095,N_9154);
nor U9937 (N_9937,N_9132,N_9307);
nor U9938 (N_9938,N_9330,N_9085);
nand U9939 (N_9939,N_9175,N_9070);
nor U9940 (N_9940,N_9159,N_9145);
or U9941 (N_9941,N_9125,N_9399);
nand U9942 (N_9942,N_9029,N_9364);
nor U9943 (N_9943,N_9430,N_9395);
and U9944 (N_9944,N_9394,N_9292);
nor U9945 (N_9945,N_9164,N_9420);
nand U9946 (N_9946,N_9146,N_9076);
nand U9947 (N_9947,N_9455,N_9033);
and U9948 (N_9948,N_9062,N_9326);
nor U9949 (N_9949,N_9392,N_9045);
and U9950 (N_9950,N_9368,N_9339);
and U9951 (N_9951,N_9044,N_9031);
nor U9952 (N_9952,N_9329,N_9354);
nor U9953 (N_9953,N_9270,N_9168);
nand U9954 (N_9954,N_9136,N_9293);
and U9955 (N_9955,N_9027,N_9100);
or U9956 (N_9956,N_9061,N_9380);
and U9957 (N_9957,N_9391,N_9387);
or U9958 (N_9958,N_9253,N_9186);
nand U9959 (N_9959,N_9344,N_9214);
nor U9960 (N_9960,N_9225,N_9334);
nor U9961 (N_9961,N_9097,N_9001);
nor U9962 (N_9962,N_9335,N_9202);
nand U9963 (N_9963,N_9032,N_9232);
xnor U9964 (N_9964,N_9166,N_9326);
nor U9965 (N_9965,N_9046,N_9342);
and U9966 (N_9966,N_9352,N_9364);
xor U9967 (N_9967,N_9072,N_9466);
or U9968 (N_9968,N_9124,N_9207);
nand U9969 (N_9969,N_9054,N_9063);
xor U9970 (N_9970,N_9252,N_9390);
and U9971 (N_9971,N_9202,N_9316);
nor U9972 (N_9972,N_9355,N_9044);
nor U9973 (N_9973,N_9168,N_9379);
nand U9974 (N_9974,N_9231,N_9258);
or U9975 (N_9975,N_9188,N_9454);
nand U9976 (N_9976,N_9361,N_9035);
nor U9977 (N_9977,N_9203,N_9120);
or U9978 (N_9978,N_9020,N_9103);
nor U9979 (N_9979,N_9119,N_9201);
and U9980 (N_9980,N_9049,N_9198);
nor U9981 (N_9981,N_9160,N_9122);
or U9982 (N_9982,N_9460,N_9391);
or U9983 (N_9983,N_9378,N_9278);
or U9984 (N_9984,N_9332,N_9049);
nor U9985 (N_9985,N_9055,N_9348);
nor U9986 (N_9986,N_9226,N_9017);
nand U9987 (N_9987,N_9291,N_9148);
nand U9988 (N_9988,N_9406,N_9391);
nand U9989 (N_9989,N_9225,N_9193);
and U9990 (N_9990,N_9005,N_9135);
nand U9991 (N_9991,N_9476,N_9042);
xnor U9992 (N_9992,N_9100,N_9181);
or U9993 (N_9993,N_9450,N_9270);
nand U9994 (N_9994,N_9058,N_9188);
nor U9995 (N_9995,N_9325,N_9118);
and U9996 (N_9996,N_9443,N_9164);
or U9997 (N_9997,N_9034,N_9152);
nor U9998 (N_9998,N_9179,N_9084);
or U9999 (N_9999,N_9099,N_9025);
or U10000 (N_10000,N_9862,N_9597);
nand U10001 (N_10001,N_9795,N_9755);
xor U10002 (N_10002,N_9901,N_9968);
and U10003 (N_10003,N_9926,N_9943);
nor U10004 (N_10004,N_9650,N_9891);
or U10005 (N_10005,N_9548,N_9687);
nor U10006 (N_10006,N_9974,N_9937);
nor U10007 (N_10007,N_9619,N_9515);
nor U10008 (N_10008,N_9531,N_9574);
xor U10009 (N_10009,N_9736,N_9859);
nand U10010 (N_10010,N_9964,N_9777);
nor U10011 (N_10011,N_9931,N_9723);
or U10012 (N_10012,N_9607,N_9939);
xnor U10013 (N_10013,N_9642,N_9789);
xnor U10014 (N_10014,N_9667,N_9684);
and U10015 (N_10015,N_9646,N_9598);
nand U10016 (N_10016,N_9674,N_9616);
or U10017 (N_10017,N_9893,N_9634);
or U10018 (N_10018,N_9711,N_9912);
and U10019 (N_10019,N_9949,N_9641);
nand U10020 (N_10020,N_9657,N_9779);
nor U10021 (N_10021,N_9975,N_9860);
nor U10022 (N_10022,N_9782,N_9997);
nor U10023 (N_10023,N_9883,N_9742);
or U10024 (N_10024,N_9835,N_9735);
or U10025 (N_10025,N_9524,N_9986);
and U10026 (N_10026,N_9856,N_9694);
nor U10027 (N_10027,N_9849,N_9588);
or U10028 (N_10028,N_9505,N_9567);
or U10029 (N_10029,N_9638,N_9722);
or U10030 (N_10030,N_9831,N_9513);
xnor U10031 (N_10031,N_9727,N_9999);
nand U10032 (N_10032,N_9786,N_9996);
and U10033 (N_10033,N_9960,N_9594);
or U10034 (N_10034,N_9550,N_9698);
nor U10035 (N_10035,N_9544,N_9644);
xnor U10036 (N_10036,N_9927,N_9696);
nand U10037 (N_10037,N_9848,N_9649);
nand U10038 (N_10038,N_9998,N_9867);
and U10039 (N_10039,N_9826,N_9523);
or U10040 (N_10040,N_9655,N_9717);
nor U10041 (N_10041,N_9765,N_9857);
and U10042 (N_10042,N_9551,N_9695);
and U10043 (N_10043,N_9706,N_9784);
or U10044 (N_10044,N_9744,N_9908);
nor U10045 (N_10045,N_9560,N_9572);
xor U10046 (N_10046,N_9580,N_9971);
or U10047 (N_10047,N_9842,N_9953);
nand U10048 (N_10048,N_9764,N_9658);
and U10049 (N_10049,N_9704,N_9525);
nor U10050 (N_10050,N_9627,N_9679);
nand U10051 (N_10051,N_9639,N_9762);
nand U10052 (N_10052,N_9942,N_9577);
nand U10053 (N_10053,N_9756,N_9804);
nor U10054 (N_10054,N_9571,N_9824);
or U10055 (N_10055,N_9903,N_9909);
xor U10056 (N_10056,N_9759,N_9651);
nand U10057 (N_10057,N_9946,N_9589);
or U10058 (N_10058,N_9618,N_9885);
or U10059 (N_10059,N_9892,N_9630);
and U10060 (N_10060,N_9739,N_9967);
nand U10061 (N_10061,N_9512,N_9582);
or U10062 (N_10062,N_9629,N_9771);
xor U10063 (N_10063,N_9747,N_9873);
nand U10064 (N_10064,N_9570,N_9624);
or U10065 (N_10065,N_9569,N_9614);
or U10066 (N_10066,N_9750,N_9621);
nor U10067 (N_10067,N_9994,N_9781);
nand U10068 (N_10068,N_9635,N_9534);
or U10069 (N_10069,N_9836,N_9693);
nor U10070 (N_10070,N_9915,N_9886);
and U10071 (N_10071,N_9626,N_9982);
nand U10072 (N_10072,N_9713,N_9977);
xnor U10073 (N_10073,N_9905,N_9681);
nor U10074 (N_10074,N_9659,N_9884);
nand U10075 (N_10075,N_9729,N_9832);
nand U10076 (N_10076,N_9555,N_9591);
and U10077 (N_10077,N_9530,N_9925);
and U10078 (N_10078,N_9888,N_9951);
and U10079 (N_10079,N_9928,N_9734);
xnor U10080 (N_10080,N_9522,N_9573);
nand U10081 (N_10081,N_9520,N_9583);
and U10082 (N_10082,N_9774,N_9984);
nor U10083 (N_10083,N_9954,N_9558);
nor U10084 (N_10084,N_9894,N_9830);
or U10085 (N_10085,N_9839,N_9890);
and U10086 (N_10086,N_9669,N_9564);
or U10087 (N_10087,N_9853,N_9615);
and U10088 (N_10088,N_9796,N_9748);
or U10089 (N_10089,N_9566,N_9633);
xnor U10090 (N_10090,N_9606,N_9906);
or U10091 (N_10091,N_9604,N_9897);
nor U10092 (N_10092,N_9590,N_9881);
and U10093 (N_10093,N_9872,N_9563);
or U10094 (N_10094,N_9846,N_9691);
nand U10095 (N_10095,N_9837,N_9985);
or U10096 (N_10096,N_9533,N_9780);
and U10097 (N_10097,N_9840,N_9958);
nor U10098 (N_10098,N_9677,N_9625);
or U10099 (N_10099,N_9654,N_9632);
and U10100 (N_10100,N_9851,N_9876);
nand U10101 (N_10101,N_9553,N_9724);
or U10102 (N_10102,N_9913,N_9866);
and U10103 (N_10103,N_9602,N_9965);
nand U10104 (N_10104,N_9895,N_9957);
xor U10105 (N_10105,N_9709,N_9676);
and U10106 (N_10106,N_9559,N_9705);
and U10107 (N_10107,N_9944,N_9834);
nand U10108 (N_10108,N_9617,N_9763);
xor U10109 (N_10109,N_9510,N_9543);
nand U10110 (N_10110,N_9752,N_9686);
and U10111 (N_10111,N_9929,N_9934);
or U10112 (N_10112,N_9767,N_9875);
xnor U10113 (N_10113,N_9869,N_9757);
nor U10114 (N_10114,N_9532,N_9863);
nor U10115 (N_10115,N_9508,N_9562);
or U10116 (N_10116,N_9899,N_9587);
and U10117 (N_10117,N_9637,N_9678);
xor U10118 (N_10118,N_9683,N_9714);
nand U10119 (N_10119,N_9807,N_9575);
nand U10120 (N_10120,N_9993,N_9665);
nand U10121 (N_10121,N_9932,N_9506);
or U10122 (N_10122,N_9648,N_9672);
and U10123 (N_10123,N_9877,N_9671);
nand U10124 (N_10124,N_9896,N_9690);
and U10125 (N_10125,N_9864,N_9822);
nor U10126 (N_10126,N_9502,N_9865);
and U10127 (N_10127,N_9702,N_9666);
and U10128 (N_10128,N_9956,N_9668);
xor U10129 (N_10129,N_9970,N_9940);
and U10130 (N_10130,N_9811,N_9511);
nand U10131 (N_10131,N_9697,N_9976);
nand U10132 (N_10132,N_9791,N_9730);
nor U10133 (N_10133,N_9586,N_9871);
nor U10134 (N_10134,N_9647,N_9808);
xor U10135 (N_10135,N_9947,N_9825);
nand U10136 (N_10136,N_9797,N_9814);
nor U10137 (N_10137,N_9518,N_9992);
nor U10138 (N_10138,N_9879,N_9663);
and U10139 (N_10139,N_9904,N_9978);
or U10140 (N_10140,N_9703,N_9517);
or U10141 (N_10141,N_9770,N_9847);
and U10142 (N_10142,N_9973,N_9787);
or U10143 (N_10143,N_9661,N_9793);
nor U10144 (N_10144,N_9778,N_9546);
nor U10145 (N_10145,N_9898,N_9568);
xor U10146 (N_10146,N_9753,N_9952);
and U10147 (N_10147,N_9631,N_9504);
or U10148 (N_10148,N_9963,N_9838);
or U10149 (N_10149,N_9813,N_9552);
and U10150 (N_10150,N_9707,N_9576);
and U10151 (N_10151,N_9751,N_9861);
nand U10152 (N_10152,N_9745,N_9785);
or U10153 (N_10153,N_9930,N_9989);
nand U10154 (N_10154,N_9538,N_9628);
nand U10155 (N_10155,N_9981,N_9950);
or U10156 (N_10156,N_9802,N_9775);
or U10157 (N_10157,N_9578,N_9673);
nor U10158 (N_10158,N_9556,N_9592);
and U10159 (N_10159,N_9919,N_9819);
or U10160 (N_10160,N_9844,N_9719);
nor U10161 (N_10161,N_9605,N_9741);
nor U10162 (N_10162,N_9725,N_9535);
nand U10163 (N_10163,N_9938,N_9769);
or U10164 (N_10164,N_9593,N_9924);
or U10165 (N_10165,N_9521,N_9547);
or U10166 (N_10166,N_9603,N_9728);
or U10167 (N_10167,N_9699,N_9921);
or U10168 (N_10168,N_9917,N_9500);
nor U10169 (N_10169,N_9596,N_9817);
or U10170 (N_10170,N_9554,N_9988);
nand U10171 (N_10171,N_9746,N_9540);
and U10172 (N_10172,N_9608,N_9829);
or U10173 (N_10173,N_9772,N_9613);
and U10174 (N_10174,N_9688,N_9692);
nand U10175 (N_10175,N_9945,N_9806);
or U10176 (N_10176,N_9955,N_9972);
or U10177 (N_10177,N_9761,N_9527);
xor U10178 (N_10178,N_9889,N_9969);
nand U10179 (N_10179,N_9983,N_9815);
nand U10180 (N_10180,N_9536,N_9620);
and U10181 (N_10181,N_9800,N_9870);
xnor U10182 (N_10182,N_9636,N_9855);
nand U10183 (N_10183,N_9599,N_9907);
nor U10184 (N_10184,N_9935,N_9585);
or U10185 (N_10185,N_9933,N_9816);
nor U10186 (N_10186,N_9812,N_9660);
and U10187 (N_10187,N_9652,N_9941);
and U10188 (N_10188,N_9503,N_9680);
nor U10189 (N_10189,N_9959,N_9990);
nand U10190 (N_10190,N_9731,N_9541);
or U10191 (N_10191,N_9880,N_9737);
and U10192 (N_10192,N_9507,N_9902);
nor U10193 (N_10193,N_9612,N_9987);
and U10194 (N_10194,N_9961,N_9827);
xor U10195 (N_10195,N_9850,N_9766);
or U10196 (N_10196,N_9798,N_9640);
or U10197 (N_10197,N_9716,N_9682);
xor U10198 (N_10198,N_9776,N_9514);
and U10199 (N_10199,N_9519,N_9708);
xor U10200 (N_10200,N_9841,N_9623);
and U10201 (N_10201,N_9738,N_9843);
and U10202 (N_10202,N_9732,N_9528);
xor U10203 (N_10203,N_9557,N_9754);
nand U10204 (N_10204,N_9675,N_9743);
nor U10205 (N_10205,N_9995,N_9792);
nor U10206 (N_10206,N_9720,N_9622);
nand U10207 (N_10207,N_9794,N_9882);
or U10208 (N_10208,N_9565,N_9936);
nand U10209 (N_10209,N_9579,N_9611);
nand U10210 (N_10210,N_9664,N_9733);
and U10211 (N_10211,N_9918,N_9799);
or U10212 (N_10212,N_9874,N_9509);
xor U10213 (N_10213,N_9803,N_9878);
nor U10214 (N_10214,N_9670,N_9581);
xor U10215 (N_10215,N_9833,N_9601);
and U10216 (N_10216,N_9689,N_9962);
nand U10217 (N_10217,N_9828,N_9810);
and U10218 (N_10218,N_9600,N_9783);
or U10219 (N_10219,N_9539,N_9922);
nor U10220 (N_10220,N_9823,N_9920);
or U10221 (N_10221,N_9718,N_9561);
or U10222 (N_10222,N_9662,N_9760);
nand U10223 (N_10223,N_9914,N_9790);
or U10224 (N_10224,N_9609,N_9758);
nand U10225 (N_10225,N_9645,N_9726);
or U10226 (N_10226,N_9820,N_9773);
nand U10227 (N_10227,N_9801,N_9653);
nand U10228 (N_10228,N_9911,N_9549);
nand U10229 (N_10229,N_9916,N_9740);
and U10230 (N_10230,N_9685,N_9845);
nand U10231 (N_10231,N_9818,N_9529);
or U10232 (N_10232,N_9710,N_9542);
or U10233 (N_10233,N_9501,N_9809);
and U10234 (N_10234,N_9656,N_9923);
nor U10235 (N_10235,N_9537,N_9712);
and U10236 (N_10236,N_9910,N_9721);
or U10237 (N_10237,N_9545,N_9854);
nor U10238 (N_10238,N_9526,N_9584);
xor U10239 (N_10239,N_9979,N_9610);
nand U10240 (N_10240,N_9991,N_9948);
and U10241 (N_10241,N_9768,N_9643);
nand U10242 (N_10242,N_9868,N_9805);
or U10243 (N_10243,N_9701,N_9858);
nor U10244 (N_10244,N_9900,N_9700);
or U10245 (N_10245,N_9516,N_9980);
or U10246 (N_10246,N_9715,N_9595);
nor U10247 (N_10247,N_9821,N_9966);
nor U10248 (N_10248,N_9788,N_9887);
nor U10249 (N_10249,N_9852,N_9749);
nand U10250 (N_10250,N_9607,N_9687);
or U10251 (N_10251,N_9787,N_9740);
and U10252 (N_10252,N_9522,N_9882);
and U10253 (N_10253,N_9604,N_9737);
or U10254 (N_10254,N_9809,N_9851);
nor U10255 (N_10255,N_9743,N_9613);
or U10256 (N_10256,N_9573,N_9995);
or U10257 (N_10257,N_9902,N_9832);
and U10258 (N_10258,N_9636,N_9875);
nor U10259 (N_10259,N_9721,N_9600);
or U10260 (N_10260,N_9792,N_9721);
or U10261 (N_10261,N_9635,N_9674);
and U10262 (N_10262,N_9931,N_9825);
or U10263 (N_10263,N_9660,N_9772);
and U10264 (N_10264,N_9993,N_9690);
xnor U10265 (N_10265,N_9997,N_9509);
and U10266 (N_10266,N_9970,N_9744);
and U10267 (N_10267,N_9750,N_9756);
or U10268 (N_10268,N_9599,N_9729);
or U10269 (N_10269,N_9831,N_9789);
nor U10270 (N_10270,N_9866,N_9559);
xor U10271 (N_10271,N_9819,N_9838);
nand U10272 (N_10272,N_9757,N_9906);
and U10273 (N_10273,N_9815,N_9916);
nor U10274 (N_10274,N_9836,N_9812);
nor U10275 (N_10275,N_9923,N_9620);
nand U10276 (N_10276,N_9862,N_9705);
nand U10277 (N_10277,N_9774,N_9861);
nor U10278 (N_10278,N_9506,N_9616);
or U10279 (N_10279,N_9678,N_9990);
nand U10280 (N_10280,N_9590,N_9610);
nor U10281 (N_10281,N_9622,N_9662);
and U10282 (N_10282,N_9923,N_9568);
nor U10283 (N_10283,N_9773,N_9743);
or U10284 (N_10284,N_9545,N_9766);
nor U10285 (N_10285,N_9989,N_9882);
nand U10286 (N_10286,N_9905,N_9871);
nand U10287 (N_10287,N_9955,N_9967);
nor U10288 (N_10288,N_9687,N_9732);
xor U10289 (N_10289,N_9818,N_9637);
nand U10290 (N_10290,N_9867,N_9598);
xor U10291 (N_10291,N_9853,N_9540);
xnor U10292 (N_10292,N_9745,N_9647);
or U10293 (N_10293,N_9642,N_9704);
nor U10294 (N_10294,N_9514,N_9740);
nor U10295 (N_10295,N_9893,N_9698);
and U10296 (N_10296,N_9507,N_9590);
nand U10297 (N_10297,N_9983,N_9826);
nand U10298 (N_10298,N_9653,N_9944);
xnor U10299 (N_10299,N_9595,N_9716);
or U10300 (N_10300,N_9767,N_9534);
xor U10301 (N_10301,N_9845,N_9791);
and U10302 (N_10302,N_9989,N_9668);
nand U10303 (N_10303,N_9821,N_9518);
or U10304 (N_10304,N_9686,N_9619);
or U10305 (N_10305,N_9816,N_9647);
xnor U10306 (N_10306,N_9595,N_9698);
nor U10307 (N_10307,N_9864,N_9624);
and U10308 (N_10308,N_9692,N_9569);
and U10309 (N_10309,N_9522,N_9878);
nor U10310 (N_10310,N_9780,N_9891);
or U10311 (N_10311,N_9778,N_9836);
nand U10312 (N_10312,N_9836,N_9740);
nand U10313 (N_10313,N_9823,N_9896);
or U10314 (N_10314,N_9784,N_9959);
and U10315 (N_10315,N_9954,N_9531);
and U10316 (N_10316,N_9577,N_9637);
or U10317 (N_10317,N_9542,N_9789);
nor U10318 (N_10318,N_9954,N_9958);
nor U10319 (N_10319,N_9772,N_9795);
or U10320 (N_10320,N_9754,N_9704);
or U10321 (N_10321,N_9916,N_9509);
and U10322 (N_10322,N_9903,N_9736);
or U10323 (N_10323,N_9664,N_9776);
and U10324 (N_10324,N_9919,N_9869);
nand U10325 (N_10325,N_9843,N_9621);
and U10326 (N_10326,N_9741,N_9728);
nand U10327 (N_10327,N_9584,N_9751);
xor U10328 (N_10328,N_9871,N_9557);
or U10329 (N_10329,N_9878,N_9663);
or U10330 (N_10330,N_9706,N_9538);
or U10331 (N_10331,N_9788,N_9612);
nand U10332 (N_10332,N_9990,N_9611);
nand U10333 (N_10333,N_9688,N_9860);
or U10334 (N_10334,N_9986,N_9765);
nand U10335 (N_10335,N_9688,N_9750);
nor U10336 (N_10336,N_9977,N_9773);
and U10337 (N_10337,N_9607,N_9873);
nand U10338 (N_10338,N_9796,N_9861);
or U10339 (N_10339,N_9719,N_9634);
nor U10340 (N_10340,N_9978,N_9945);
xor U10341 (N_10341,N_9560,N_9792);
xor U10342 (N_10342,N_9791,N_9907);
nor U10343 (N_10343,N_9748,N_9747);
or U10344 (N_10344,N_9914,N_9500);
nor U10345 (N_10345,N_9903,N_9832);
nand U10346 (N_10346,N_9725,N_9839);
nand U10347 (N_10347,N_9917,N_9695);
xor U10348 (N_10348,N_9700,N_9551);
and U10349 (N_10349,N_9527,N_9531);
or U10350 (N_10350,N_9986,N_9790);
nand U10351 (N_10351,N_9941,N_9834);
nand U10352 (N_10352,N_9615,N_9550);
and U10353 (N_10353,N_9619,N_9800);
and U10354 (N_10354,N_9722,N_9694);
xor U10355 (N_10355,N_9953,N_9803);
nand U10356 (N_10356,N_9608,N_9830);
and U10357 (N_10357,N_9708,N_9684);
xnor U10358 (N_10358,N_9877,N_9726);
or U10359 (N_10359,N_9586,N_9823);
and U10360 (N_10360,N_9558,N_9907);
or U10361 (N_10361,N_9761,N_9658);
nor U10362 (N_10362,N_9969,N_9839);
or U10363 (N_10363,N_9743,N_9975);
and U10364 (N_10364,N_9738,N_9826);
and U10365 (N_10365,N_9745,N_9793);
nor U10366 (N_10366,N_9699,N_9557);
nand U10367 (N_10367,N_9877,N_9981);
nor U10368 (N_10368,N_9746,N_9551);
nor U10369 (N_10369,N_9568,N_9683);
or U10370 (N_10370,N_9520,N_9553);
nand U10371 (N_10371,N_9730,N_9669);
and U10372 (N_10372,N_9502,N_9678);
nand U10373 (N_10373,N_9939,N_9602);
nor U10374 (N_10374,N_9695,N_9733);
or U10375 (N_10375,N_9847,N_9941);
nand U10376 (N_10376,N_9503,N_9701);
and U10377 (N_10377,N_9918,N_9938);
xnor U10378 (N_10378,N_9822,N_9517);
nor U10379 (N_10379,N_9624,N_9577);
nor U10380 (N_10380,N_9649,N_9648);
or U10381 (N_10381,N_9621,N_9972);
nand U10382 (N_10382,N_9509,N_9998);
and U10383 (N_10383,N_9841,N_9566);
or U10384 (N_10384,N_9711,N_9673);
nand U10385 (N_10385,N_9924,N_9959);
xnor U10386 (N_10386,N_9665,N_9981);
or U10387 (N_10387,N_9842,N_9950);
or U10388 (N_10388,N_9788,N_9746);
and U10389 (N_10389,N_9738,N_9705);
nand U10390 (N_10390,N_9763,N_9689);
nand U10391 (N_10391,N_9514,N_9882);
xnor U10392 (N_10392,N_9624,N_9627);
or U10393 (N_10393,N_9769,N_9856);
xor U10394 (N_10394,N_9632,N_9700);
xnor U10395 (N_10395,N_9545,N_9578);
nand U10396 (N_10396,N_9632,N_9578);
nor U10397 (N_10397,N_9863,N_9768);
nor U10398 (N_10398,N_9936,N_9643);
xnor U10399 (N_10399,N_9560,N_9953);
and U10400 (N_10400,N_9635,N_9899);
nor U10401 (N_10401,N_9878,N_9582);
and U10402 (N_10402,N_9847,N_9991);
nor U10403 (N_10403,N_9889,N_9761);
xor U10404 (N_10404,N_9956,N_9882);
nand U10405 (N_10405,N_9747,N_9876);
xnor U10406 (N_10406,N_9532,N_9921);
nor U10407 (N_10407,N_9975,N_9620);
and U10408 (N_10408,N_9750,N_9513);
nor U10409 (N_10409,N_9524,N_9582);
nand U10410 (N_10410,N_9618,N_9610);
or U10411 (N_10411,N_9579,N_9817);
xor U10412 (N_10412,N_9663,N_9785);
or U10413 (N_10413,N_9880,N_9555);
or U10414 (N_10414,N_9956,N_9670);
or U10415 (N_10415,N_9936,N_9571);
and U10416 (N_10416,N_9877,N_9992);
and U10417 (N_10417,N_9688,N_9851);
nor U10418 (N_10418,N_9662,N_9834);
or U10419 (N_10419,N_9992,N_9703);
or U10420 (N_10420,N_9704,N_9970);
or U10421 (N_10421,N_9988,N_9598);
xnor U10422 (N_10422,N_9510,N_9564);
nand U10423 (N_10423,N_9586,N_9761);
or U10424 (N_10424,N_9931,N_9750);
or U10425 (N_10425,N_9711,N_9659);
and U10426 (N_10426,N_9893,N_9633);
nor U10427 (N_10427,N_9916,N_9906);
xnor U10428 (N_10428,N_9756,N_9642);
xor U10429 (N_10429,N_9790,N_9983);
xnor U10430 (N_10430,N_9674,N_9940);
nor U10431 (N_10431,N_9540,N_9781);
and U10432 (N_10432,N_9549,N_9540);
nor U10433 (N_10433,N_9508,N_9633);
xor U10434 (N_10434,N_9759,N_9864);
or U10435 (N_10435,N_9861,N_9712);
nand U10436 (N_10436,N_9712,N_9595);
nand U10437 (N_10437,N_9767,N_9506);
or U10438 (N_10438,N_9544,N_9906);
nand U10439 (N_10439,N_9561,N_9837);
nor U10440 (N_10440,N_9990,N_9644);
nor U10441 (N_10441,N_9971,N_9615);
and U10442 (N_10442,N_9872,N_9816);
and U10443 (N_10443,N_9715,N_9942);
nand U10444 (N_10444,N_9600,N_9887);
or U10445 (N_10445,N_9673,N_9582);
nand U10446 (N_10446,N_9837,N_9743);
nand U10447 (N_10447,N_9793,N_9627);
and U10448 (N_10448,N_9539,N_9904);
nor U10449 (N_10449,N_9630,N_9787);
and U10450 (N_10450,N_9548,N_9725);
and U10451 (N_10451,N_9652,N_9821);
nand U10452 (N_10452,N_9652,N_9642);
and U10453 (N_10453,N_9779,N_9635);
or U10454 (N_10454,N_9747,N_9941);
or U10455 (N_10455,N_9802,N_9739);
and U10456 (N_10456,N_9874,N_9720);
or U10457 (N_10457,N_9915,N_9547);
nand U10458 (N_10458,N_9876,N_9559);
nand U10459 (N_10459,N_9723,N_9829);
nor U10460 (N_10460,N_9564,N_9605);
or U10461 (N_10461,N_9729,N_9665);
xor U10462 (N_10462,N_9619,N_9549);
xor U10463 (N_10463,N_9866,N_9940);
and U10464 (N_10464,N_9893,N_9718);
nand U10465 (N_10465,N_9560,N_9791);
nand U10466 (N_10466,N_9796,N_9879);
nor U10467 (N_10467,N_9784,N_9734);
nand U10468 (N_10468,N_9733,N_9811);
and U10469 (N_10469,N_9510,N_9597);
nor U10470 (N_10470,N_9862,N_9884);
nor U10471 (N_10471,N_9996,N_9703);
nor U10472 (N_10472,N_9669,N_9651);
nand U10473 (N_10473,N_9953,N_9532);
or U10474 (N_10474,N_9869,N_9691);
xor U10475 (N_10475,N_9670,N_9846);
or U10476 (N_10476,N_9694,N_9648);
nor U10477 (N_10477,N_9659,N_9683);
or U10478 (N_10478,N_9627,N_9885);
nand U10479 (N_10479,N_9543,N_9990);
or U10480 (N_10480,N_9708,N_9687);
nand U10481 (N_10481,N_9810,N_9715);
nand U10482 (N_10482,N_9757,N_9622);
nand U10483 (N_10483,N_9527,N_9953);
nand U10484 (N_10484,N_9644,N_9968);
or U10485 (N_10485,N_9555,N_9561);
nor U10486 (N_10486,N_9868,N_9887);
and U10487 (N_10487,N_9821,N_9784);
nand U10488 (N_10488,N_9589,N_9655);
nor U10489 (N_10489,N_9832,N_9761);
nand U10490 (N_10490,N_9870,N_9806);
nand U10491 (N_10491,N_9970,N_9701);
or U10492 (N_10492,N_9855,N_9556);
nand U10493 (N_10493,N_9910,N_9812);
nor U10494 (N_10494,N_9778,N_9766);
nand U10495 (N_10495,N_9919,N_9579);
nor U10496 (N_10496,N_9502,N_9897);
nand U10497 (N_10497,N_9918,N_9758);
nand U10498 (N_10498,N_9637,N_9898);
nand U10499 (N_10499,N_9991,N_9950);
xor U10500 (N_10500,N_10000,N_10346);
and U10501 (N_10501,N_10242,N_10126);
nand U10502 (N_10502,N_10337,N_10127);
xnor U10503 (N_10503,N_10104,N_10143);
nor U10504 (N_10504,N_10198,N_10328);
and U10505 (N_10505,N_10443,N_10116);
or U10506 (N_10506,N_10339,N_10172);
nor U10507 (N_10507,N_10332,N_10473);
xnor U10508 (N_10508,N_10350,N_10268);
nor U10509 (N_10509,N_10037,N_10378);
and U10510 (N_10510,N_10330,N_10239);
xor U10511 (N_10511,N_10015,N_10275);
xnor U10512 (N_10512,N_10438,N_10007);
nand U10513 (N_10513,N_10179,N_10412);
nor U10514 (N_10514,N_10379,N_10449);
or U10515 (N_10515,N_10170,N_10358);
nand U10516 (N_10516,N_10311,N_10025);
nand U10517 (N_10517,N_10314,N_10383);
or U10518 (N_10518,N_10023,N_10221);
nand U10519 (N_10519,N_10130,N_10257);
and U10520 (N_10520,N_10207,N_10128);
nand U10521 (N_10521,N_10133,N_10093);
xnor U10522 (N_10522,N_10353,N_10120);
and U10523 (N_10523,N_10177,N_10114);
nand U10524 (N_10524,N_10453,N_10399);
nand U10525 (N_10525,N_10169,N_10039);
nand U10526 (N_10526,N_10360,N_10220);
nand U10527 (N_10527,N_10495,N_10077);
or U10528 (N_10528,N_10302,N_10209);
nor U10529 (N_10529,N_10151,N_10471);
nor U10530 (N_10530,N_10183,N_10206);
xnor U10531 (N_10531,N_10167,N_10042);
xor U10532 (N_10532,N_10331,N_10058);
and U10533 (N_10533,N_10244,N_10241);
or U10534 (N_10534,N_10131,N_10173);
nand U10535 (N_10535,N_10430,N_10470);
or U10536 (N_10536,N_10057,N_10103);
nor U10537 (N_10537,N_10138,N_10456);
or U10538 (N_10538,N_10124,N_10272);
or U10539 (N_10539,N_10299,N_10301);
nor U10540 (N_10540,N_10361,N_10408);
and U10541 (N_10541,N_10459,N_10026);
nor U10542 (N_10542,N_10341,N_10251);
or U10543 (N_10543,N_10188,N_10118);
nor U10544 (N_10544,N_10297,N_10451);
xor U10545 (N_10545,N_10038,N_10392);
xor U10546 (N_10546,N_10010,N_10098);
or U10547 (N_10547,N_10181,N_10248);
nor U10548 (N_10548,N_10427,N_10310);
and U10549 (N_10549,N_10215,N_10434);
and U10550 (N_10550,N_10067,N_10278);
nand U10551 (N_10551,N_10422,N_10082);
nor U10552 (N_10552,N_10288,N_10006);
xnor U10553 (N_10553,N_10364,N_10236);
and U10554 (N_10554,N_10458,N_10031);
nor U10555 (N_10555,N_10429,N_10185);
nor U10556 (N_10556,N_10426,N_10070);
nand U10557 (N_10557,N_10411,N_10295);
xor U10558 (N_10558,N_10217,N_10385);
and U10559 (N_10559,N_10410,N_10322);
or U10560 (N_10560,N_10400,N_10072);
and U10561 (N_10561,N_10155,N_10159);
or U10562 (N_10562,N_10324,N_10327);
and U10563 (N_10563,N_10457,N_10212);
nand U10564 (N_10564,N_10321,N_10208);
nand U10565 (N_10565,N_10040,N_10441);
and U10566 (N_10566,N_10001,N_10352);
nor U10567 (N_10567,N_10413,N_10111);
nand U10568 (N_10568,N_10276,N_10291);
nor U10569 (N_10569,N_10498,N_10326);
xor U10570 (N_10570,N_10474,N_10191);
or U10571 (N_10571,N_10432,N_10223);
or U10572 (N_10572,N_10329,N_10219);
nor U10573 (N_10573,N_10323,N_10303);
nor U10574 (N_10574,N_10240,N_10439);
nor U10575 (N_10575,N_10189,N_10238);
nor U10576 (N_10576,N_10109,N_10161);
and U10577 (N_10577,N_10149,N_10390);
nor U10578 (N_10578,N_10335,N_10068);
and U10579 (N_10579,N_10256,N_10099);
and U10580 (N_10580,N_10313,N_10416);
xnor U10581 (N_10581,N_10389,N_10482);
nand U10582 (N_10582,N_10370,N_10259);
and U10583 (N_10583,N_10063,N_10483);
or U10584 (N_10584,N_10394,N_10014);
nand U10585 (N_10585,N_10190,N_10154);
and U10586 (N_10586,N_10147,N_10083);
xor U10587 (N_10587,N_10137,N_10445);
nand U10588 (N_10588,N_10407,N_10317);
nor U10589 (N_10589,N_10405,N_10105);
and U10590 (N_10590,N_10139,N_10032);
and U10591 (N_10591,N_10363,N_10140);
nand U10592 (N_10592,N_10296,N_10287);
and U10593 (N_10593,N_10271,N_10371);
nor U10594 (N_10594,N_10395,N_10008);
or U10595 (N_10595,N_10146,N_10141);
nor U10596 (N_10596,N_10267,N_10162);
xnor U10597 (N_10597,N_10334,N_10125);
nor U10598 (N_10598,N_10309,N_10064);
nand U10599 (N_10599,N_10305,N_10112);
and U10600 (N_10600,N_10499,N_10036);
nor U10601 (N_10601,N_10076,N_10002);
nand U10602 (N_10602,N_10092,N_10380);
nor U10603 (N_10603,N_10053,N_10199);
nor U10604 (N_10604,N_10101,N_10466);
nor U10605 (N_10605,N_10168,N_10454);
nor U10606 (N_10606,N_10487,N_10056);
and U10607 (N_10607,N_10234,N_10013);
nand U10608 (N_10608,N_10372,N_10343);
nand U10609 (N_10609,N_10210,N_10280);
or U10610 (N_10610,N_10480,N_10315);
nor U10611 (N_10611,N_10110,N_10373);
nor U10612 (N_10612,N_10387,N_10145);
nor U10613 (N_10613,N_10467,N_10096);
nand U10614 (N_10614,N_10362,N_10277);
or U10615 (N_10615,N_10213,N_10122);
nand U10616 (N_10616,N_10347,N_10193);
and U10617 (N_10617,N_10368,N_10021);
and U10618 (N_10618,N_10074,N_10100);
and U10619 (N_10619,N_10090,N_10293);
or U10620 (N_10620,N_10428,N_10022);
or U10621 (N_10621,N_10142,N_10418);
and U10622 (N_10622,N_10160,N_10084);
or U10623 (N_10623,N_10086,N_10226);
and U10624 (N_10624,N_10034,N_10342);
nand U10625 (N_10625,N_10113,N_10490);
or U10626 (N_10626,N_10369,N_10479);
and U10627 (N_10627,N_10166,N_10175);
and U10628 (N_10628,N_10320,N_10005);
or U10629 (N_10629,N_10018,N_10153);
nand U10630 (N_10630,N_10393,N_10406);
and U10631 (N_10631,N_10115,N_10069);
nor U10632 (N_10632,N_10060,N_10089);
and U10633 (N_10633,N_10150,N_10071);
nor U10634 (N_10634,N_10435,N_10016);
or U10635 (N_10635,N_10455,N_10450);
nand U10636 (N_10636,N_10041,N_10079);
or U10637 (N_10637,N_10349,N_10059);
and U10638 (N_10638,N_10247,N_10357);
and U10639 (N_10639,N_10306,N_10384);
nand U10640 (N_10640,N_10003,N_10237);
and U10641 (N_10641,N_10123,N_10336);
and U10642 (N_10642,N_10431,N_10365);
or U10643 (N_10643,N_10048,N_10318);
and U10644 (N_10644,N_10367,N_10419);
and U10645 (N_10645,N_10216,N_10028);
xnor U10646 (N_10646,N_10469,N_10134);
nand U10647 (N_10647,N_10121,N_10494);
nor U10648 (N_10648,N_10255,N_10496);
and U10649 (N_10649,N_10289,N_10464);
or U10650 (N_10650,N_10078,N_10017);
nor U10651 (N_10651,N_10300,N_10081);
and U10652 (N_10652,N_10231,N_10214);
nor U10653 (N_10653,N_10135,N_10264);
nor U10654 (N_10654,N_10396,N_10061);
nand U10655 (N_10655,N_10417,N_10273);
and U10656 (N_10656,N_10148,N_10436);
xnor U10657 (N_10657,N_10024,N_10187);
nor U10658 (N_10658,N_10117,N_10243);
or U10659 (N_10659,N_10286,N_10265);
and U10660 (N_10660,N_10027,N_10062);
nand U10661 (N_10661,N_10157,N_10262);
xnor U10662 (N_10662,N_10492,N_10233);
nor U10663 (N_10663,N_10433,N_10283);
or U10664 (N_10664,N_10468,N_10182);
and U10665 (N_10665,N_10020,N_10230);
and U10666 (N_10666,N_10075,N_10246);
and U10667 (N_10667,N_10478,N_10088);
nor U10668 (N_10668,N_10398,N_10340);
nand U10669 (N_10669,N_10448,N_10249);
and U10670 (N_10670,N_10282,N_10202);
and U10671 (N_10671,N_10260,N_10054);
nor U10672 (N_10672,N_10366,N_10475);
or U10673 (N_10673,N_10012,N_10356);
nor U10674 (N_10674,N_10106,N_10194);
and U10675 (N_10675,N_10298,N_10333);
or U10676 (N_10676,N_10144,N_10269);
nand U10677 (N_10677,N_10164,N_10107);
nand U10678 (N_10678,N_10044,N_10294);
nand U10679 (N_10679,N_10196,N_10091);
or U10680 (N_10680,N_10055,N_10319);
nand U10681 (N_10681,N_10108,N_10222);
nor U10682 (N_10682,N_10488,N_10472);
nor U10683 (N_10683,N_10258,N_10035);
or U10684 (N_10684,N_10095,N_10484);
nor U10685 (N_10685,N_10355,N_10174);
nand U10686 (N_10686,N_10485,N_10308);
nor U10687 (N_10687,N_10119,N_10442);
nor U10688 (N_10688,N_10029,N_10270);
and U10689 (N_10689,N_10386,N_10489);
nand U10690 (N_10690,N_10486,N_10359);
nand U10691 (N_10691,N_10403,N_10197);
nand U10692 (N_10692,N_10129,N_10052);
and U10693 (N_10693,N_10253,N_10065);
and U10694 (N_10694,N_10254,N_10465);
nand U10695 (N_10695,N_10046,N_10171);
nor U10696 (N_10696,N_10307,N_10178);
or U10697 (N_10697,N_10225,N_10163);
nand U10698 (N_10698,N_10376,N_10304);
or U10699 (N_10699,N_10446,N_10043);
nor U10700 (N_10700,N_10045,N_10437);
xor U10701 (N_10701,N_10476,N_10423);
and U10702 (N_10702,N_10227,N_10094);
and U10703 (N_10703,N_10011,N_10425);
xor U10704 (N_10704,N_10452,N_10477);
and U10705 (N_10705,N_10132,N_10284);
and U10706 (N_10706,N_10158,N_10415);
and U10707 (N_10707,N_10377,N_10201);
nor U10708 (N_10708,N_10374,N_10424);
nor U10709 (N_10709,N_10420,N_10281);
or U10710 (N_10710,N_10338,N_10229);
nand U10711 (N_10711,N_10051,N_10218);
nand U10712 (N_10712,N_10290,N_10312);
nand U10713 (N_10713,N_10261,N_10030);
and U10714 (N_10714,N_10404,N_10049);
nand U10715 (N_10715,N_10156,N_10414);
or U10716 (N_10716,N_10136,N_10224);
nor U10717 (N_10717,N_10354,N_10263);
nor U10718 (N_10718,N_10004,N_10087);
and U10719 (N_10719,N_10345,N_10292);
nor U10720 (N_10720,N_10200,N_10344);
and U10721 (N_10721,N_10388,N_10402);
nor U10722 (N_10722,N_10497,N_10325);
nor U10723 (N_10723,N_10205,N_10176);
nand U10724 (N_10724,N_10409,N_10204);
nand U10725 (N_10725,N_10316,N_10401);
and U10726 (N_10726,N_10444,N_10186);
or U10727 (N_10727,N_10245,N_10252);
nor U10728 (N_10728,N_10381,N_10203);
and U10729 (N_10729,N_10211,N_10235);
nand U10730 (N_10730,N_10180,N_10232);
nor U10731 (N_10731,N_10009,N_10461);
or U10732 (N_10732,N_10080,N_10397);
nand U10733 (N_10733,N_10285,N_10491);
xor U10734 (N_10734,N_10375,N_10279);
xnor U10735 (N_10735,N_10462,N_10066);
or U10736 (N_10736,N_10195,N_10097);
xnor U10737 (N_10737,N_10351,N_10152);
nand U10738 (N_10738,N_10391,N_10050);
nand U10739 (N_10739,N_10274,N_10493);
nor U10740 (N_10740,N_10184,N_10481);
nand U10741 (N_10741,N_10421,N_10073);
nand U10742 (N_10742,N_10192,N_10348);
or U10743 (N_10743,N_10460,N_10447);
nor U10744 (N_10744,N_10382,N_10085);
nor U10745 (N_10745,N_10228,N_10250);
and U10746 (N_10746,N_10165,N_10033);
and U10747 (N_10747,N_10102,N_10440);
nor U10748 (N_10748,N_10019,N_10266);
or U10749 (N_10749,N_10463,N_10047);
nor U10750 (N_10750,N_10414,N_10461);
nor U10751 (N_10751,N_10245,N_10442);
nand U10752 (N_10752,N_10331,N_10399);
xnor U10753 (N_10753,N_10304,N_10188);
nand U10754 (N_10754,N_10035,N_10034);
or U10755 (N_10755,N_10097,N_10306);
xor U10756 (N_10756,N_10158,N_10232);
or U10757 (N_10757,N_10438,N_10378);
nand U10758 (N_10758,N_10050,N_10085);
nor U10759 (N_10759,N_10469,N_10467);
nand U10760 (N_10760,N_10050,N_10186);
and U10761 (N_10761,N_10263,N_10379);
nor U10762 (N_10762,N_10174,N_10417);
or U10763 (N_10763,N_10207,N_10482);
nor U10764 (N_10764,N_10112,N_10191);
or U10765 (N_10765,N_10049,N_10195);
and U10766 (N_10766,N_10039,N_10311);
and U10767 (N_10767,N_10017,N_10118);
xor U10768 (N_10768,N_10292,N_10001);
nor U10769 (N_10769,N_10384,N_10005);
or U10770 (N_10770,N_10061,N_10244);
xor U10771 (N_10771,N_10389,N_10305);
nand U10772 (N_10772,N_10076,N_10222);
or U10773 (N_10773,N_10276,N_10413);
and U10774 (N_10774,N_10118,N_10057);
and U10775 (N_10775,N_10149,N_10133);
or U10776 (N_10776,N_10255,N_10471);
nor U10777 (N_10777,N_10065,N_10494);
and U10778 (N_10778,N_10300,N_10338);
nand U10779 (N_10779,N_10163,N_10271);
or U10780 (N_10780,N_10018,N_10451);
nor U10781 (N_10781,N_10288,N_10370);
or U10782 (N_10782,N_10281,N_10011);
nand U10783 (N_10783,N_10496,N_10034);
or U10784 (N_10784,N_10460,N_10094);
or U10785 (N_10785,N_10346,N_10479);
or U10786 (N_10786,N_10026,N_10348);
nor U10787 (N_10787,N_10225,N_10354);
and U10788 (N_10788,N_10426,N_10425);
xnor U10789 (N_10789,N_10333,N_10284);
nand U10790 (N_10790,N_10396,N_10377);
nand U10791 (N_10791,N_10473,N_10498);
and U10792 (N_10792,N_10378,N_10087);
nand U10793 (N_10793,N_10146,N_10347);
nor U10794 (N_10794,N_10433,N_10373);
nand U10795 (N_10795,N_10152,N_10126);
or U10796 (N_10796,N_10320,N_10069);
or U10797 (N_10797,N_10202,N_10022);
and U10798 (N_10798,N_10235,N_10384);
or U10799 (N_10799,N_10185,N_10419);
xnor U10800 (N_10800,N_10435,N_10171);
and U10801 (N_10801,N_10190,N_10274);
nor U10802 (N_10802,N_10354,N_10188);
xor U10803 (N_10803,N_10407,N_10264);
and U10804 (N_10804,N_10299,N_10410);
nor U10805 (N_10805,N_10313,N_10431);
and U10806 (N_10806,N_10214,N_10272);
xor U10807 (N_10807,N_10377,N_10286);
nor U10808 (N_10808,N_10471,N_10201);
or U10809 (N_10809,N_10093,N_10332);
xnor U10810 (N_10810,N_10085,N_10138);
or U10811 (N_10811,N_10466,N_10204);
and U10812 (N_10812,N_10064,N_10499);
xor U10813 (N_10813,N_10205,N_10499);
or U10814 (N_10814,N_10055,N_10028);
and U10815 (N_10815,N_10160,N_10415);
and U10816 (N_10816,N_10151,N_10136);
nor U10817 (N_10817,N_10194,N_10161);
nand U10818 (N_10818,N_10466,N_10479);
and U10819 (N_10819,N_10479,N_10311);
nor U10820 (N_10820,N_10140,N_10124);
nand U10821 (N_10821,N_10221,N_10115);
or U10822 (N_10822,N_10086,N_10253);
nand U10823 (N_10823,N_10333,N_10189);
nor U10824 (N_10824,N_10243,N_10465);
nor U10825 (N_10825,N_10390,N_10272);
or U10826 (N_10826,N_10228,N_10171);
and U10827 (N_10827,N_10013,N_10243);
nor U10828 (N_10828,N_10117,N_10320);
or U10829 (N_10829,N_10428,N_10385);
nand U10830 (N_10830,N_10251,N_10174);
nand U10831 (N_10831,N_10381,N_10347);
xnor U10832 (N_10832,N_10195,N_10266);
or U10833 (N_10833,N_10013,N_10216);
and U10834 (N_10834,N_10462,N_10094);
nor U10835 (N_10835,N_10119,N_10253);
and U10836 (N_10836,N_10303,N_10247);
nand U10837 (N_10837,N_10032,N_10087);
or U10838 (N_10838,N_10369,N_10016);
nand U10839 (N_10839,N_10085,N_10342);
or U10840 (N_10840,N_10197,N_10391);
nor U10841 (N_10841,N_10283,N_10133);
and U10842 (N_10842,N_10057,N_10023);
xor U10843 (N_10843,N_10087,N_10396);
nor U10844 (N_10844,N_10004,N_10366);
nor U10845 (N_10845,N_10452,N_10214);
and U10846 (N_10846,N_10356,N_10145);
or U10847 (N_10847,N_10353,N_10449);
nand U10848 (N_10848,N_10272,N_10343);
nor U10849 (N_10849,N_10063,N_10193);
or U10850 (N_10850,N_10370,N_10389);
nand U10851 (N_10851,N_10145,N_10316);
or U10852 (N_10852,N_10486,N_10345);
nor U10853 (N_10853,N_10070,N_10486);
nor U10854 (N_10854,N_10158,N_10320);
xnor U10855 (N_10855,N_10101,N_10001);
nand U10856 (N_10856,N_10317,N_10443);
and U10857 (N_10857,N_10101,N_10156);
xor U10858 (N_10858,N_10347,N_10186);
or U10859 (N_10859,N_10416,N_10021);
xor U10860 (N_10860,N_10170,N_10013);
nor U10861 (N_10861,N_10356,N_10336);
nand U10862 (N_10862,N_10480,N_10032);
and U10863 (N_10863,N_10363,N_10055);
nor U10864 (N_10864,N_10171,N_10099);
nand U10865 (N_10865,N_10278,N_10471);
nand U10866 (N_10866,N_10040,N_10015);
or U10867 (N_10867,N_10393,N_10124);
and U10868 (N_10868,N_10254,N_10437);
nor U10869 (N_10869,N_10435,N_10425);
or U10870 (N_10870,N_10230,N_10070);
or U10871 (N_10871,N_10359,N_10287);
or U10872 (N_10872,N_10289,N_10434);
nand U10873 (N_10873,N_10301,N_10371);
xor U10874 (N_10874,N_10372,N_10091);
or U10875 (N_10875,N_10243,N_10251);
and U10876 (N_10876,N_10328,N_10450);
nand U10877 (N_10877,N_10104,N_10478);
nand U10878 (N_10878,N_10174,N_10075);
or U10879 (N_10879,N_10330,N_10201);
nand U10880 (N_10880,N_10172,N_10018);
or U10881 (N_10881,N_10159,N_10156);
and U10882 (N_10882,N_10448,N_10103);
nand U10883 (N_10883,N_10265,N_10143);
or U10884 (N_10884,N_10190,N_10078);
and U10885 (N_10885,N_10011,N_10211);
nand U10886 (N_10886,N_10000,N_10243);
nor U10887 (N_10887,N_10189,N_10022);
xnor U10888 (N_10888,N_10354,N_10387);
or U10889 (N_10889,N_10141,N_10340);
nor U10890 (N_10890,N_10390,N_10264);
nor U10891 (N_10891,N_10146,N_10327);
or U10892 (N_10892,N_10462,N_10033);
or U10893 (N_10893,N_10394,N_10452);
and U10894 (N_10894,N_10491,N_10080);
nand U10895 (N_10895,N_10362,N_10080);
xnor U10896 (N_10896,N_10399,N_10330);
nor U10897 (N_10897,N_10287,N_10026);
nor U10898 (N_10898,N_10240,N_10134);
xor U10899 (N_10899,N_10078,N_10479);
or U10900 (N_10900,N_10484,N_10195);
or U10901 (N_10901,N_10235,N_10190);
and U10902 (N_10902,N_10326,N_10389);
nand U10903 (N_10903,N_10182,N_10364);
nand U10904 (N_10904,N_10491,N_10197);
nor U10905 (N_10905,N_10103,N_10426);
xor U10906 (N_10906,N_10288,N_10277);
nor U10907 (N_10907,N_10120,N_10344);
and U10908 (N_10908,N_10461,N_10201);
nor U10909 (N_10909,N_10174,N_10475);
and U10910 (N_10910,N_10497,N_10354);
and U10911 (N_10911,N_10124,N_10431);
or U10912 (N_10912,N_10256,N_10162);
and U10913 (N_10913,N_10028,N_10220);
or U10914 (N_10914,N_10135,N_10314);
and U10915 (N_10915,N_10460,N_10395);
or U10916 (N_10916,N_10007,N_10201);
xnor U10917 (N_10917,N_10127,N_10024);
nand U10918 (N_10918,N_10286,N_10174);
xnor U10919 (N_10919,N_10305,N_10074);
nand U10920 (N_10920,N_10060,N_10169);
xnor U10921 (N_10921,N_10261,N_10089);
or U10922 (N_10922,N_10370,N_10347);
or U10923 (N_10923,N_10298,N_10451);
nor U10924 (N_10924,N_10129,N_10417);
and U10925 (N_10925,N_10373,N_10268);
nand U10926 (N_10926,N_10043,N_10420);
and U10927 (N_10927,N_10013,N_10186);
or U10928 (N_10928,N_10334,N_10078);
nand U10929 (N_10929,N_10206,N_10156);
xnor U10930 (N_10930,N_10044,N_10014);
nand U10931 (N_10931,N_10221,N_10211);
and U10932 (N_10932,N_10187,N_10129);
or U10933 (N_10933,N_10430,N_10055);
nor U10934 (N_10934,N_10017,N_10437);
nand U10935 (N_10935,N_10463,N_10247);
nor U10936 (N_10936,N_10198,N_10247);
nand U10937 (N_10937,N_10130,N_10485);
nor U10938 (N_10938,N_10038,N_10335);
nand U10939 (N_10939,N_10172,N_10228);
or U10940 (N_10940,N_10060,N_10313);
nand U10941 (N_10941,N_10080,N_10089);
or U10942 (N_10942,N_10208,N_10244);
nor U10943 (N_10943,N_10306,N_10074);
and U10944 (N_10944,N_10084,N_10221);
and U10945 (N_10945,N_10040,N_10342);
nand U10946 (N_10946,N_10145,N_10483);
and U10947 (N_10947,N_10448,N_10233);
or U10948 (N_10948,N_10182,N_10098);
nand U10949 (N_10949,N_10257,N_10446);
and U10950 (N_10950,N_10341,N_10410);
and U10951 (N_10951,N_10251,N_10325);
nand U10952 (N_10952,N_10418,N_10459);
or U10953 (N_10953,N_10431,N_10006);
nand U10954 (N_10954,N_10078,N_10363);
and U10955 (N_10955,N_10438,N_10376);
and U10956 (N_10956,N_10036,N_10246);
nand U10957 (N_10957,N_10296,N_10465);
nor U10958 (N_10958,N_10494,N_10486);
or U10959 (N_10959,N_10067,N_10150);
or U10960 (N_10960,N_10049,N_10451);
nand U10961 (N_10961,N_10110,N_10138);
and U10962 (N_10962,N_10371,N_10356);
nand U10963 (N_10963,N_10169,N_10451);
xnor U10964 (N_10964,N_10323,N_10435);
and U10965 (N_10965,N_10337,N_10308);
or U10966 (N_10966,N_10248,N_10200);
or U10967 (N_10967,N_10249,N_10092);
and U10968 (N_10968,N_10162,N_10186);
and U10969 (N_10969,N_10091,N_10050);
nand U10970 (N_10970,N_10147,N_10317);
or U10971 (N_10971,N_10034,N_10258);
nand U10972 (N_10972,N_10044,N_10408);
nand U10973 (N_10973,N_10225,N_10290);
or U10974 (N_10974,N_10285,N_10404);
and U10975 (N_10975,N_10373,N_10150);
nand U10976 (N_10976,N_10385,N_10235);
or U10977 (N_10977,N_10391,N_10120);
or U10978 (N_10978,N_10201,N_10225);
nand U10979 (N_10979,N_10174,N_10200);
nand U10980 (N_10980,N_10127,N_10341);
nand U10981 (N_10981,N_10453,N_10052);
or U10982 (N_10982,N_10032,N_10293);
and U10983 (N_10983,N_10292,N_10372);
xnor U10984 (N_10984,N_10200,N_10214);
and U10985 (N_10985,N_10256,N_10345);
nor U10986 (N_10986,N_10424,N_10031);
nand U10987 (N_10987,N_10292,N_10057);
nor U10988 (N_10988,N_10285,N_10060);
and U10989 (N_10989,N_10293,N_10088);
nand U10990 (N_10990,N_10327,N_10013);
or U10991 (N_10991,N_10096,N_10345);
xor U10992 (N_10992,N_10110,N_10054);
and U10993 (N_10993,N_10471,N_10024);
and U10994 (N_10994,N_10324,N_10421);
and U10995 (N_10995,N_10164,N_10467);
or U10996 (N_10996,N_10168,N_10150);
nor U10997 (N_10997,N_10129,N_10451);
xor U10998 (N_10998,N_10437,N_10247);
or U10999 (N_10999,N_10480,N_10465);
nor U11000 (N_11000,N_10630,N_10656);
nor U11001 (N_11001,N_10927,N_10524);
and U11002 (N_11002,N_10980,N_10783);
nand U11003 (N_11003,N_10887,N_10610);
or U11004 (N_11004,N_10684,N_10922);
and U11005 (N_11005,N_10811,N_10691);
and U11006 (N_11006,N_10506,N_10869);
or U11007 (N_11007,N_10649,N_10819);
nor U11008 (N_11008,N_10725,N_10778);
and U11009 (N_11009,N_10872,N_10708);
nor U11010 (N_11010,N_10860,N_10667);
or U11011 (N_11011,N_10623,N_10702);
and U11012 (N_11012,N_10902,N_10930);
or U11013 (N_11013,N_10554,N_10719);
or U11014 (N_11014,N_10535,N_10786);
and U11015 (N_11015,N_10877,N_10764);
nor U11016 (N_11016,N_10852,N_10798);
and U11017 (N_11017,N_10886,N_10678);
or U11018 (N_11018,N_10876,N_10611);
nand U11019 (N_11019,N_10654,N_10742);
or U11020 (N_11020,N_10991,N_10963);
or U11021 (N_11021,N_10933,N_10743);
nor U11022 (N_11022,N_10787,N_10788);
or U11023 (N_11023,N_10957,N_10964);
xor U11024 (N_11024,N_10646,N_10879);
nor U11025 (N_11025,N_10587,N_10899);
xnor U11026 (N_11026,N_10936,N_10552);
or U11027 (N_11027,N_10857,N_10500);
nor U11028 (N_11028,N_10975,N_10782);
and U11029 (N_11029,N_10873,N_10961);
and U11030 (N_11030,N_10695,N_10648);
nand U11031 (N_11031,N_10780,N_10501);
or U11032 (N_11032,N_10817,N_10588);
nor U11033 (N_11033,N_10697,N_10514);
nor U11034 (N_11034,N_10973,N_10511);
nand U11035 (N_11035,N_10745,N_10823);
nor U11036 (N_11036,N_10673,N_10521);
nor U11037 (N_11037,N_10659,N_10901);
nor U11038 (N_11038,N_10700,N_10891);
nor U11039 (N_11039,N_10612,N_10502);
and U11040 (N_11040,N_10769,N_10557);
and U11041 (N_11041,N_10631,N_10945);
and U11042 (N_11042,N_10875,N_10781);
nand U11043 (N_11043,N_10520,N_10672);
nor U11044 (N_11044,N_10806,N_10613);
or U11045 (N_11045,N_10878,N_10794);
nand U11046 (N_11046,N_10638,N_10739);
xor U11047 (N_11047,N_10994,N_10581);
nor U11048 (N_11048,N_10950,N_10504);
and U11049 (N_11049,N_10566,N_10944);
nand U11050 (N_11050,N_10932,N_10776);
or U11051 (N_11051,N_10931,N_10664);
xor U11052 (N_11052,N_10698,N_10705);
and U11053 (N_11053,N_10815,N_10563);
and U11054 (N_11054,N_10885,N_10871);
or U11055 (N_11055,N_10578,N_10749);
nor U11056 (N_11056,N_10625,N_10666);
xor U11057 (N_11057,N_10660,N_10734);
and U11058 (N_11058,N_10926,N_10959);
and U11059 (N_11059,N_10593,N_10692);
or U11060 (N_11060,N_10689,N_10534);
nor U11061 (N_11061,N_10997,N_10846);
and U11062 (N_11062,N_10863,N_10981);
nand U11063 (N_11063,N_10632,N_10828);
nor U11064 (N_11064,N_10727,N_10835);
nor U11065 (N_11065,N_10586,N_10602);
nor U11066 (N_11066,N_10917,N_10532);
or U11067 (N_11067,N_10643,N_10791);
or U11068 (N_11068,N_10988,N_10754);
nor U11069 (N_11069,N_10516,N_10544);
nand U11070 (N_11070,N_10919,N_10870);
or U11071 (N_11071,N_10647,N_10948);
nand U11072 (N_11072,N_10847,N_10999);
or U11073 (N_11073,N_10793,N_10717);
or U11074 (N_11074,N_10607,N_10840);
nor U11075 (N_11075,N_10967,N_10571);
or U11076 (N_11076,N_10954,N_10834);
or U11077 (N_11077,N_10699,N_10536);
and U11078 (N_11078,N_10731,N_10539);
or U11079 (N_11079,N_10796,N_10960);
xor U11080 (N_11080,N_10748,N_10547);
nand U11081 (N_11081,N_10512,N_10738);
or U11082 (N_11082,N_10810,N_10867);
and U11083 (N_11083,N_10858,N_10903);
and U11084 (N_11084,N_10851,N_10530);
and U11085 (N_11085,N_10838,N_10909);
nand U11086 (N_11086,N_10803,N_10519);
nor U11087 (N_11087,N_10895,N_10938);
or U11088 (N_11088,N_10998,N_10768);
nor U11089 (N_11089,N_10543,N_10814);
or U11090 (N_11090,N_10579,N_10820);
nor U11091 (N_11091,N_10622,N_10560);
nor U11092 (N_11092,N_10690,N_10693);
nor U11093 (N_11093,N_10608,N_10883);
xnor U11094 (N_11094,N_10681,N_10865);
or U11095 (N_11095,N_10671,N_10812);
nand U11096 (N_11096,N_10939,N_10559);
xnor U11097 (N_11097,N_10929,N_10735);
or U11098 (N_11098,N_10561,N_10669);
xnor U11099 (N_11099,N_10525,N_10528);
xor U11100 (N_11100,N_10844,N_10890);
or U11101 (N_11101,N_10789,N_10985);
and U11102 (N_11102,N_10841,N_10972);
xnor U11103 (N_11103,N_10590,N_10624);
nand U11104 (N_11104,N_10567,N_10913);
nor U11105 (N_11105,N_10549,N_10683);
nand U11106 (N_11106,N_10912,N_10962);
or U11107 (N_11107,N_10992,N_10824);
or U11108 (N_11108,N_10598,N_10657);
nand U11109 (N_11109,N_10505,N_10976);
nand U11110 (N_11110,N_10915,N_10984);
and U11111 (N_11111,N_10759,N_10617);
nor U11112 (N_11112,N_10658,N_10849);
or U11113 (N_11113,N_10510,N_10827);
and U11114 (N_11114,N_10515,N_10644);
nor U11115 (N_11115,N_10527,N_10934);
and U11116 (N_11116,N_10688,N_10861);
nor U11117 (N_11117,N_10522,N_10682);
nor U11118 (N_11118,N_10898,N_10799);
or U11119 (N_11119,N_10836,N_10969);
or U11120 (N_11120,N_10965,N_10637);
or U11121 (N_11121,N_10509,N_10640);
nand U11122 (N_11122,N_10585,N_10952);
and U11123 (N_11123,N_10756,N_10541);
and U11124 (N_11124,N_10596,N_10765);
nor U11125 (N_11125,N_10779,N_10545);
or U11126 (N_11126,N_10795,N_10784);
nor U11127 (N_11127,N_10553,N_10568);
nor U11128 (N_11128,N_10755,N_10573);
nor U11129 (N_11129,N_10940,N_10661);
nor U11130 (N_11130,N_10816,N_10966);
xor U11131 (N_11131,N_10881,N_10642);
nand U11132 (N_11132,N_10508,N_10868);
xor U11133 (N_11133,N_10686,N_10813);
nand U11134 (N_11134,N_10629,N_10709);
nand U11135 (N_11135,N_10805,N_10925);
or U11136 (N_11136,N_10848,N_10874);
and U11137 (N_11137,N_10729,N_10518);
nor U11138 (N_11138,N_10685,N_10721);
and U11139 (N_11139,N_10777,N_10542);
xnor U11140 (N_11140,N_10880,N_10905);
nor U11141 (N_11141,N_10641,N_10946);
or U11142 (N_11142,N_10856,N_10750);
or U11143 (N_11143,N_10604,N_10548);
nand U11144 (N_11144,N_10947,N_10958);
nand U11145 (N_11145,N_10722,N_10723);
nand U11146 (N_11146,N_10970,N_10911);
or U11147 (N_11147,N_10626,N_10983);
and U11148 (N_11148,N_10942,N_10853);
nand U11149 (N_11149,N_10715,N_10996);
xor U11150 (N_11150,N_10503,N_10760);
and U11151 (N_11151,N_10758,N_10540);
nor U11152 (N_11152,N_10845,N_10884);
nor U11153 (N_11153,N_10757,N_10572);
xnor U11154 (N_11154,N_10974,N_10651);
or U11155 (N_11155,N_10740,N_10986);
nand U11156 (N_11156,N_10989,N_10652);
nor U11157 (N_11157,N_10894,N_10565);
nor U11158 (N_11158,N_10943,N_10562);
and U11159 (N_11159,N_10538,N_10804);
xor U11160 (N_11160,N_10928,N_10687);
nand U11161 (N_11161,N_10977,N_10951);
nor U11162 (N_11162,N_10546,N_10599);
nand U11163 (N_11163,N_10718,N_10713);
nor U11164 (N_11164,N_10730,N_10882);
nand U11165 (N_11165,N_10826,N_10897);
nor U11166 (N_11166,N_10821,N_10818);
nor U11167 (N_11167,N_10595,N_10751);
nor U11168 (N_11168,N_10792,N_10843);
nand U11169 (N_11169,N_10703,N_10569);
nand U11170 (N_11170,N_10766,N_10770);
and U11171 (N_11171,N_10771,N_10767);
and U11172 (N_11172,N_10580,N_10955);
and U11173 (N_11173,N_10710,N_10907);
nor U11174 (N_11174,N_10639,N_10918);
and U11175 (N_11175,N_10935,N_10716);
and U11176 (N_11176,N_10971,N_10577);
nor U11177 (N_11177,N_10707,N_10551);
and U11178 (N_11178,N_10908,N_10712);
nor U11179 (N_11179,N_10910,N_10773);
or U11180 (N_11180,N_10862,N_10592);
or U11181 (N_11181,N_10513,N_10696);
nor U11182 (N_11182,N_10825,N_10761);
nand U11183 (N_11183,N_10829,N_10726);
and U11184 (N_11184,N_10753,N_10724);
xor U11185 (N_11185,N_10859,N_10762);
or U11186 (N_11186,N_10990,N_10855);
and U11187 (N_11187,N_10746,N_10822);
or U11188 (N_11188,N_10674,N_10892);
or U11189 (N_11189,N_10645,N_10555);
xnor U11190 (N_11190,N_10529,N_10653);
or U11191 (N_11191,N_10741,N_10614);
nand U11192 (N_11192,N_10634,N_10763);
nand U11193 (N_11193,N_10728,N_10558);
and U11194 (N_11194,N_10982,N_10675);
and U11195 (N_11195,N_10774,N_10635);
nand U11196 (N_11196,N_10866,N_10550);
nor U11197 (N_11197,N_10920,N_10864);
or U11198 (N_11198,N_10680,N_10785);
nand U11199 (N_11199,N_10790,N_10801);
nand U11200 (N_11200,N_10582,N_10616);
nor U11201 (N_11201,N_10854,N_10628);
xor U11202 (N_11202,N_10526,N_10670);
and U11203 (N_11203,N_10995,N_10594);
nand U11204 (N_11204,N_10618,N_10591);
or U11205 (N_11205,N_10677,N_10747);
and U11206 (N_11206,N_10837,N_10663);
or U11207 (N_11207,N_10993,N_10606);
and U11208 (N_11208,N_10619,N_10701);
xnor U11209 (N_11209,N_10956,N_10733);
and U11210 (N_11210,N_10900,N_10775);
xnor U11211 (N_11211,N_10978,N_10711);
and U11212 (N_11212,N_10809,N_10802);
nand U11213 (N_11213,N_10842,N_10523);
or U11214 (N_11214,N_10831,N_10797);
nor U11215 (N_11215,N_10916,N_10807);
and U11216 (N_11216,N_10633,N_10636);
nand U11217 (N_11217,N_10839,N_10714);
nand U11218 (N_11218,N_10665,N_10850);
xor U11219 (N_11219,N_10570,N_10923);
nor U11220 (N_11220,N_10676,N_10583);
or U11221 (N_11221,N_10650,N_10889);
and U11222 (N_11222,N_10906,N_10833);
and U11223 (N_11223,N_10832,N_10600);
and U11224 (N_11224,N_10904,N_10941);
nor U11225 (N_11225,N_10979,N_10517);
and U11226 (N_11226,N_10737,N_10888);
nand U11227 (N_11227,N_10575,N_10830);
and U11228 (N_11228,N_10704,N_10921);
or U11229 (N_11229,N_10937,N_10968);
nand U11230 (N_11230,N_10533,N_10720);
and U11231 (N_11231,N_10736,N_10627);
or U11232 (N_11232,N_10603,N_10507);
or U11233 (N_11233,N_10987,N_10949);
or U11234 (N_11234,N_10589,N_10615);
and U11235 (N_11235,N_10621,N_10609);
or U11236 (N_11236,N_10574,N_10732);
nor U11237 (N_11237,N_10679,N_10655);
xor U11238 (N_11238,N_10601,N_10576);
nand U11239 (N_11239,N_10772,N_10556);
or U11240 (N_11240,N_10668,N_10564);
nor U11241 (N_11241,N_10744,N_10694);
and U11242 (N_11242,N_10620,N_10800);
or U11243 (N_11243,N_10706,N_10896);
nand U11244 (N_11244,N_10584,N_10531);
and U11245 (N_11245,N_10924,N_10597);
nor U11246 (N_11246,N_10605,N_10953);
xnor U11247 (N_11247,N_10893,N_10662);
xor U11248 (N_11248,N_10914,N_10752);
or U11249 (N_11249,N_10537,N_10808);
or U11250 (N_11250,N_10517,N_10789);
or U11251 (N_11251,N_10537,N_10884);
nor U11252 (N_11252,N_10900,N_10599);
xnor U11253 (N_11253,N_10612,N_10884);
and U11254 (N_11254,N_10832,N_10839);
nand U11255 (N_11255,N_10896,N_10569);
or U11256 (N_11256,N_10502,N_10583);
or U11257 (N_11257,N_10816,N_10800);
xor U11258 (N_11258,N_10976,N_10922);
nand U11259 (N_11259,N_10558,N_10612);
nand U11260 (N_11260,N_10650,N_10929);
nand U11261 (N_11261,N_10980,N_10770);
or U11262 (N_11262,N_10884,N_10507);
nor U11263 (N_11263,N_10703,N_10686);
or U11264 (N_11264,N_10993,N_10646);
xnor U11265 (N_11265,N_10752,N_10681);
nand U11266 (N_11266,N_10864,N_10724);
nor U11267 (N_11267,N_10949,N_10980);
nor U11268 (N_11268,N_10542,N_10829);
nand U11269 (N_11269,N_10829,N_10626);
nor U11270 (N_11270,N_10565,N_10649);
and U11271 (N_11271,N_10781,N_10784);
nand U11272 (N_11272,N_10904,N_10715);
and U11273 (N_11273,N_10780,N_10866);
nand U11274 (N_11274,N_10807,N_10957);
nor U11275 (N_11275,N_10540,N_10912);
or U11276 (N_11276,N_10842,N_10964);
or U11277 (N_11277,N_10877,N_10755);
nor U11278 (N_11278,N_10772,N_10935);
or U11279 (N_11279,N_10834,N_10716);
xnor U11280 (N_11280,N_10556,N_10947);
xnor U11281 (N_11281,N_10568,N_10524);
nand U11282 (N_11282,N_10947,N_10783);
nand U11283 (N_11283,N_10730,N_10818);
and U11284 (N_11284,N_10836,N_10881);
and U11285 (N_11285,N_10529,N_10556);
or U11286 (N_11286,N_10947,N_10950);
xnor U11287 (N_11287,N_10657,N_10761);
and U11288 (N_11288,N_10972,N_10667);
and U11289 (N_11289,N_10930,N_10854);
nor U11290 (N_11290,N_10613,N_10909);
or U11291 (N_11291,N_10802,N_10971);
and U11292 (N_11292,N_10677,N_10652);
xnor U11293 (N_11293,N_10847,N_10675);
and U11294 (N_11294,N_10737,N_10573);
or U11295 (N_11295,N_10670,N_10763);
xor U11296 (N_11296,N_10690,N_10826);
and U11297 (N_11297,N_10753,N_10729);
and U11298 (N_11298,N_10584,N_10753);
and U11299 (N_11299,N_10592,N_10952);
nor U11300 (N_11300,N_10508,N_10596);
xnor U11301 (N_11301,N_10751,N_10619);
nor U11302 (N_11302,N_10601,N_10930);
xor U11303 (N_11303,N_10771,N_10885);
and U11304 (N_11304,N_10796,N_10905);
or U11305 (N_11305,N_10800,N_10917);
nand U11306 (N_11306,N_10676,N_10525);
nand U11307 (N_11307,N_10870,N_10512);
or U11308 (N_11308,N_10920,N_10916);
nand U11309 (N_11309,N_10910,N_10785);
or U11310 (N_11310,N_10996,N_10514);
nand U11311 (N_11311,N_10705,N_10693);
and U11312 (N_11312,N_10684,N_10997);
or U11313 (N_11313,N_10810,N_10651);
and U11314 (N_11314,N_10791,N_10817);
nand U11315 (N_11315,N_10589,N_10598);
nor U11316 (N_11316,N_10822,N_10982);
or U11317 (N_11317,N_10643,N_10681);
xor U11318 (N_11318,N_10965,N_10663);
or U11319 (N_11319,N_10658,N_10601);
nand U11320 (N_11320,N_10528,N_10949);
nand U11321 (N_11321,N_10648,N_10786);
and U11322 (N_11322,N_10984,N_10692);
or U11323 (N_11323,N_10514,N_10783);
or U11324 (N_11324,N_10770,N_10791);
nand U11325 (N_11325,N_10687,N_10918);
nor U11326 (N_11326,N_10647,N_10846);
nand U11327 (N_11327,N_10644,N_10656);
xnor U11328 (N_11328,N_10680,N_10860);
nor U11329 (N_11329,N_10764,N_10855);
xor U11330 (N_11330,N_10811,N_10767);
nand U11331 (N_11331,N_10614,N_10623);
nand U11332 (N_11332,N_10748,N_10817);
nand U11333 (N_11333,N_10548,N_10538);
xnor U11334 (N_11334,N_10871,N_10632);
and U11335 (N_11335,N_10802,N_10614);
nor U11336 (N_11336,N_10525,N_10831);
nand U11337 (N_11337,N_10549,N_10932);
and U11338 (N_11338,N_10722,N_10645);
nor U11339 (N_11339,N_10860,N_10947);
xnor U11340 (N_11340,N_10894,N_10577);
and U11341 (N_11341,N_10929,N_10544);
xnor U11342 (N_11342,N_10999,N_10951);
and U11343 (N_11343,N_10828,N_10998);
nor U11344 (N_11344,N_10500,N_10955);
xor U11345 (N_11345,N_10958,N_10989);
or U11346 (N_11346,N_10936,N_10558);
nor U11347 (N_11347,N_10939,N_10879);
and U11348 (N_11348,N_10581,N_10981);
and U11349 (N_11349,N_10552,N_10706);
or U11350 (N_11350,N_10786,N_10608);
and U11351 (N_11351,N_10637,N_10867);
nor U11352 (N_11352,N_10609,N_10667);
nand U11353 (N_11353,N_10906,N_10631);
or U11354 (N_11354,N_10763,N_10631);
or U11355 (N_11355,N_10775,N_10591);
or U11356 (N_11356,N_10668,N_10736);
xnor U11357 (N_11357,N_10638,N_10606);
or U11358 (N_11358,N_10849,N_10897);
xnor U11359 (N_11359,N_10812,N_10879);
or U11360 (N_11360,N_10838,N_10973);
nand U11361 (N_11361,N_10900,N_10823);
nand U11362 (N_11362,N_10851,N_10899);
nand U11363 (N_11363,N_10884,N_10627);
or U11364 (N_11364,N_10917,N_10727);
nand U11365 (N_11365,N_10974,N_10797);
nor U11366 (N_11366,N_10743,N_10846);
or U11367 (N_11367,N_10707,N_10821);
nor U11368 (N_11368,N_10543,N_10808);
and U11369 (N_11369,N_10836,N_10882);
nor U11370 (N_11370,N_10618,N_10734);
nand U11371 (N_11371,N_10813,N_10561);
xor U11372 (N_11372,N_10716,N_10619);
nor U11373 (N_11373,N_10636,N_10856);
nor U11374 (N_11374,N_10741,N_10574);
or U11375 (N_11375,N_10778,N_10715);
nand U11376 (N_11376,N_10628,N_10636);
and U11377 (N_11377,N_10903,N_10861);
and U11378 (N_11378,N_10925,N_10560);
nor U11379 (N_11379,N_10911,N_10700);
or U11380 (N_11380,N_10757,N_10985);
nor U11381 (N_11381,N_10708,N_10565);
and U11382 (N_11382,N_10538,N_10714);
or U11383 (N_11383,N_10992,N_10633);
or U11384 (N_11384,N_10793,N_10597);
nor U11385 (N_11385,N_10542,N_10999);
nand U11386 (N_11386,N_10874,N_10775);
and U11387 (N_11387,N_10607,N_10770);
and U11388 (N_11388,N_10881,N_10524);
nor U11389 (N_11389,N_10714,N_10772);
and U11390 (N_11390,N_10560,N_10950);
or U11391 (N_11391,N_10506,N_10659);
xor U11392 (N_11392,N_10533,N_10755);
nor U11393 (N_11393,N_10806,N_10858);
nand U11394 (N_11394,N_10773,N_10587);
nand U11395 (N_11395,N_10904,N_10731);
and U11396 (N_11396,N_10704,N_10562);
and U11397 (N_11397,N_10992,N_10709);
nand U11398 (N_11398,N_10617,N_10791);
and U11399 (N_11399,N_10698,N_10861);
and U11400 (N_11400,N_10758,N_10728);
xnor U11401 (N_11401,N_10883,N_10683);
and U11402 (N_11402,N_10575,N_10810);
and U11403 (N_11403,N_10986,N_10617);
nand U11404 (N_11404,N_10970,N_10936);
and U11405 (N_11405,N_10515,N_10970);
nor U11406 (N_11406,N_10573,N_10926);
nor U11407 (N_11407,N_10606,N_10933);
nor U11408 (N_11408,N_10866,N_10668);
nand U11409 (N_11409,N_10770,N_10957);
nand U11410 (N_11410,N_10520,N_10714);
xor U11411 (N_11411,N_10516,N_10999);
and U11412 (N_11412,N_10751,N_10794);
nand U11413 (N_11413,N_10790,N_10810);
xnor U11414 (N_11414,N_10654,N_10798);
and U11415 (N_11415,N_10516,N_10912);
and U11416 (N_11416,N_10874,N_10952);
nand U11417 (N_11417,N_10761,N_10930);
nand U11418 (N_11418,N_10692,N_10750);
or U11419 (N_11419,N_10922,N_10797);
xor U11420 (N_11420,N_10679,N_10862);
nor U11421 (N_11421,N_10962,N_10984);
and U11422 (N_11422,N_10586,N_10714);
nor U11423 (N_11423,N_10717,N_10600);
nand U11424 (N_11424,N_10989,N_10826);
nand U11425 (N_11425,N_10726,N_10581);
nand U11426 (N_11426,N_10988,N_10681);
or U11427 (N_11427,N_10517,N_10683);
or U11428 (N_11428,N_10638,N_10756);
xnor U11429 (N_11429,N_10537,N_10724);
or U11430 (N_11430,N_10715,N_10620);
nand U11431 (N_11431,N_10701,N_10939);
nor U11432 (N_11432,N_10869,N_10713);
or U11433 (N_11433,N_10619,N_10547);
nor U11434 (N_11434,N_10615,N_10875);
xor U11435 (N_11435,N_10665,N_10962);
or U11436 (N_11436,N_10988,N_10669);
nor U11437 (N_11437,N_10940,N_10627);
or U11438 (N_11438,N_10797,N_10587);
and U11439 (N_11439,N_10818,N_10755);
xor U11440 (N_11440,N_10959,N_10653);
and U11441 (N_11441,N_10919,N_10820);
xor U11442 (N_11442,N_10664,N_10646);
or U11443 (N_11443,N_10869,N_10750);
nand U11444 (N_11444,N_10828,N_10928);
and U11445 (N_11445,N_10981,N_10817);
xor U11446 (N_11446,N_10906,N_10721);
nor U11447 (N_11447,N_10980,N_10750);
and U11448 (N_11448,N_10617,N_10952);
and U11449 (N_11449,N_10810,N_10525);
or U11450 (N_11450,N_10645,N_10593);
nor U11451 (N_11451,N_10742,N_10523);
or U11452 (N_11452,N_10629,N_10534);
nand U11453 (N_11453,N_10511,N_10581);
or U11454 (N_11454,N_10726,N_10952);
or U11455 (N_11455,N_10976,N_10580);
and U11456 (N_11456,N_10821,N_10572);
nor U11457 (N_11457,N_10915,N_10534);
nor U11458 (N_11458,N_10986,N_10872);
and U11459 (N_11459,N_10713,N_10979);
or U11460 (N_11460,N_10861,N_10765);
or U11461 (N_11461,N_10857,N_10919);
nor U11462 (N_11462,N_10648,N_10801);
nand U11463 (N_11463,N_10672,N_10764);
or U11464 (N_11464,N_10726,N_10590);
and U11465 (N_11465,N_10919,N_10613);
nand U11466 (N_11466,N_10578,N_10646);
or U11467 (N_11467,N_10693,N_10926);
nand U11468 (N_11468,N_10694,N_10503);
xor U11469 (N_11469,N_10883,N_10658);
or U11470 (N_11470,N_10557,N_10668);
or U11471 (N_11471,N_10729,N_10877);
or U11472 (N_11472,N_10989,N_10851);
nor U11473 (N_11473,N_10904,N_10916);
xnor U11474 (N_11474,N_10935,N_10642);
nand U11475 (N_11475,N_10580,N_10541);
nor U11476 (N_11476,N_10780,N_10789);
or U11477 (N_11477,N_10606,N_10946);
and U11478 (N_11478,N_10875,N_10699);
nand U11479 (N_11479,N_10784,N_10581);
or U11480 (N_11480,N_10737,N_10801);
nand U11481 (N_11481,N_10912,N_10966);
and U11482 (N_11482,N_10880,N_10650);
nand U11483 (N_11483,N_10614,N_10548);
and U11484 (N_11484,N_10762,N_10840);
or U11485 (N_11485,N_10778,N_10608);
xnor U11486 (N_11486,N_10837,N_10533);
xor U11487 (N_11487,N_10718,N_10647);
and U11488 (N_11488,N_10792,N_10644);
and U11489 (N_11489,N_10863,N_10792);
nor U11490 (N_11490,N_10653,N_10936);
xor U11491 (N_11491,N_10930,N_10592);
or U11492 (N_11492,N_10799,N_10647);
nor U11493 (N_11493,N_10599,N_10976);
or U11494 (N_11494,N_10832,N_10582);
nand U11495 (N_11495,N_10569,N_10659);
xor U11496 (N_11496,N_10807,N_10599);
xor U11497 (N_11497,N_10547,N_10525);
and U11498 (N_11498,N_10586,N_10980);
nand U11499 (N_11499,N_10618,N_10552);
and U11500 (N_11500,N_11087,N_11245);
xnor U11501 (N_11501,N_11280,N_11478);
nand U11502 (N_11502,N_11160,N_11052);
or U11503 (N_11503,N_11187,N_11413);
or U11504 (N_11504,N_11110,N_11104);
nor U11505 (N_11505,N_11246,N_11290);
nor U11506 (N_11506,N_11143,N_11232);
xor U11507 (N_11507,N_11208,N_11310);
and U11508 (N_11508,N_11020,N_11100);
and U11509 (N_11509,N_11205,N_11119);
and U11510 (N_11510,N_11046,N_11498);
or U11511 (N_11511,N_11499,N_11121);
nor U11512 (N_11512,N_11481,N_11383);
nand U11513 (N_11513,N_11170,N_11157);
nand U11514 (N_11514,N_11353,N_11103);
nand U11515 (N_11515,N_11029,N_11146);
xnor U11516 (N_11516,N_11471,N_11359);
nor U11517 (N_11517,N_11089,N_11321);
nor U11518 (N_11518,N_11124,N_11377);
and U11519 (N_11519,N_11236,N_11319);
nand U11520 (N_11520,N_11128,N_11283);
or U11521 (N_11521,N_11333,N_11425);
and U11522 (N_11522,N_11265,N_11045);
xnor U11523 (N_11523,N_11060,N_11204);
nand U11524 (N_11524,N_11444,N_11196);
nand U11525 (N_11525,N_11426,N_11311);
or U11526 (N_11526,N_11022,N_11497);
and U11527 (N_11527,N_11320,N_11276);
and U11528 (N_11528,N_11023,N_11431);
nand U11529 (N_11529,N_11449,N_11443);
nor U11530 (N_11530,N_11420,N_11317);
nor U11531 (N_11531,N_11194,N_11423);
nand U11532 (N_11532,N_11483,N_11343);
and U11533 (N_11533,N_11244,N_11237);
nor U11534 (N_11534,N_11145,N_11054);
xnor U11535 (N_11535,N_11493,N_11010);
and U11536 (N_11536,N_11374,N_11486);
nor U11537 (N_11537,N_11357,N_11177);
and U11538 (N_11538,N_11451,N_11132);
nand U11539 (N_11539,N_11172,N_11150);
or U11540 (N_11540,N_11301,N_11082);
and U11541 (N_11541,N_11180,N_11432);
or U11542 (N_11542,N_11488,N_11101);
nand U11543 (N_11543,N_11448,N_11238);
or U11544 (N_11544,N_11026,N_11436);
or U11545 (N_11545,N_11464,N_11324);
xor U11546 (N_11546,N_11427,N_11279);
or U11547 (N_11547,N_11171,N_11085);
and U11548 (N_11548,N_11458,N_11215);
nor U11549 (N_11549,N_11140,N_11491);
and U11550 (N_11550,N_11003,N_11252);
and U11551 (N_11551,N_11259,N_11284);
xor U11552 (N_11552,N_11038,N_11162);
nor U11553 (N_11553,N_11064,N_11393);
nor U11554 (N_11554,N_11013,N_11113);
and U11555 (N_11555,N_11401,N_11164);
and U11556 (N_11556,N_11463,N_11175);
nand U11557 (N_11557,N_11335,N_11061);
and U11558 (N_11558,N_11278,N_11330);
nand U11559 (N_11559,N_11461,N_11467);
nor U11560 (N_11560,N_11405,N_11350);
or U11561 (N_11561,N_11342,N_11167);
nand U11562 (N_11562,N_11201,N_11091);
and U11563 (N_11563,N_11056,N_11302);
nor U11564 (N_11564,N_11406,N_11161);
and U11565 (N_11565,N_11385,N_11270);
and U11566 (N_11566,N_11078,N_11037);
nand U11567 (N_11567,N_11351,N_11239);
nand U11568 (N_11568,N_11067,N_11370);
nand U11569 (N_11569,N_11039,N_11105);
and U11570 (N_11570,N_11218,N_11466);
nor U11571 (N_11571,N_11347,N_11084);
xnor U11572 (N_11572,N_11277,N_11072);
xor U11573 (N_11573,N_11378,N_11261);
nand U11574 (N_11574,N_11178,N_11477);
nor U11575 (N_11575,N_11005,N_11266);
nor U11576 (N_11576,N_11095,N_11395);
nor U11577 (N_11577,N_11168,N_11441);
and U11578 (N_11578,N_11040,N_11271);
nor U11579 (N_11579,N_11358,N_11211);
or U11580 (N_11580,N_11484,N_11041);
xor U11581 (N_11581,N_11231,N_11349);
or U11582 (N_11582,N_11249,N_11016);
nand U11583 (N_11583,N_11473,N_11438);
or U11584 (N_11584,N_11248,N_11356);
and U11585 (N_11585,N_11344,N_11086);
and U11586 (N_11586,N_11126,N_11305);
xnor U11587 (N_11587,N_11043,N_11116);
nor U11588 (N_11588,N_11409,N_11313);
and U11589 (N_11589,N_11314,N_11312);
nand U11590 (N_11590,N_11340,N_11053);
nor U11591 (N_11591,N_11185,N_11400);
and U11592 (N_11592,N_11285,N_11366);
nand U11593 (N_11593,N_11228,N_11000);
nor U11594 (N_11594,N_11027,N_11057);
xnor U11595 (N_11595,N_11256,N_11325);
nand U11596 (N_11596,N_11118,N_11114);
or U11597 (N_11597,N_11042,N_11480);
and U11598 (N_11598,N_11223,N_11364);
and U11599 (N_11599,N_11083,N_11068);
nor U11600 (N_11600,N_11058,N_11273);
nand U11601 (N_11601,N_11470,N_11389);
and U11602 (N_11602,N_11482,N_11099);
nand U11603 (N_11603,N_11227,N_11354);
and U11604 (N_11604,N_11345,N_11012);
and U11605 (N_11605,N_11080,N_11474);
nor U11606 (N_11606,N_11050,N_11148);
nand U11607 (N_11607,N_11049,N_11450);
or U11608 (N_11608,N_11291,N_11092);
xnor U11609 (N_11609,N_11308,N_11492);
nor U11610 (N_11610,N_11323,N_11251);
and U11611 (N_11611,N_11074,N_11025);
and U11612 (N_11612,N_11006,N_11334);
xnor U11613 (N_11613,N_11048,N_11288);
nor U11614 (N_11614,N_11066,N_11106);
nand U11615 (N_11615,N_11281,N_11033);
nor U11616 (N_11616,N_11004,N_11202);
or U11617 (N_11617,N_11376,N_11348);
or U11618 (N_11618,N_11390,N_11338);
or U11619 (N_11619,N_11047,N_11260);
nand U11620 (N_11620,N_11123,N_11191);
nor U11621 (N_11621,N_11015,N_11240);
or U11622 (N_11622,N_11254,N_11117);
nand U11623 (N_11623,N_11065,N_11199);
and U11624 (N_11624,N_11156,N_11032);
or U11625 (N_11625,N_11293,N_11217);
nand U11626 (N_11626,N_11138,N_11297);
nor U11627 (N_11627,N_11158,N_11306);
or U11628 (N_11628,N_11460,N_11055);
or U11629 (N_11629,N_11435,N_11115);
and U11630 (N_11630,N_11303,N_11275);
and U11631 (N_11631,N_11404,N_11188);
and U11632 (N_11632,N_11130,N_11415);
and U11633 (N_11633,N_11380,N_11430);
and U11634 (N_11634,N_11402,N_11387);
nand U11635 (N_11635,N_11331,N_11298);
and U11636 (N_11636,N_11332,N_11274);
or U11637 (N_11637,N_11440,N_11372);
nor U11638 (N_11638,N_11184,N_11129);
and U11639 (N_11639,N_11031,N_11394);
nor U11640 (N_11640,N_11447,N_11398);
xor U11641 (N_11641,N_11382,N_11097);
xor U11642 (N_11642,N_11076,N_11469);
nor U11643 (N_11643,N_11397,N_11063);
or U11644 (N_11644,N_11229,N_11001);
nand U11645 (N_11645,N_11221,N_11485);
or U11646 (N_11646,N_11365,N_11336);
nand U11647 (N_11647,N_11011,N_11088);
nand U11648 (N_11648,N_11292,N_11141);
xor U11649 (N_11649,N_11257,N_11139);
nor U11650 (N_11650,N_11422,N_11424);
or U11651 (N_11651,N_11384,N_11135);
or U11652 (N_11652,N_11225,N_11392);
nor U11653 (N_11653,N_11263,N_11341);
or U11654 (N_11654,N_11416,N_11316);
or U11655 (N_11655,N_11154,N_11017);
nor U11656 (N_11656,N_11081,N_11465);
nor U11657 (N_11657,N_11200,N_11127);
nand U11658 (N_11658,N_11073,N_11433);
or U11659 (N_11659,N_11247,N_11445);
nand U11660 (N_11660,N_11371,N_11457);
or U11661 (N_11661,N_11173,N_11136);
or U11662 (N_11662,N_11472,N_11242);
xor U11663 (N_11663,N_11018,N_11019);
or U11664 (N_11664,N_11071,N_11059);
nand U11665 (N_11665,N_11176,N_11077);
nor U11666 (N_11666,N_11355,N_11147);
nand U11667 (N_11667,N_11207,N_11375);
or U11668 (N_11668,N_11429,N_11210);
xnor U11669 (N_11669,N_11093,N_11024);
and U11670 (N_11670,N_11152,N_11109);
nand U11671 (N_11671,N_11407,N_11206);
and U11672 (N_11672,N_11307,N_11434);
and U11673 (N_11673,N_11367,N_11149);
xnor U11674 (N_11674,N_11243,N_11134);
nor U11675 (N_11675,N_11396,N_11189);
nand U11676 (N_11676,N_11021,N_11296);
and U11677 (N_11677,N_11386,N_11002);
nor U11678 (N_11678,N_11107,N_11241);
nand U11679 (N_11679,N_11326,N_11165);
and U11680 (N_11680,N_11159,N_11198);
or U11681 (N_11681,N_11454,N_11090);
or U11682 (N_11682,N_11412,N_11190);
or U11683 (N_11683,N_11036,N_11258);
nand U11684 (N_11684,N_11142,N_11182);
xor U11685 (N_11685,N_11219,N_11111);
nor U11686 (N_11686,N_11169,N_11309);
or U11687 (N_11687,N_11179,N_11192);
nand U11688 (N_11688,N_11337,N_11346);
nand U11689 (N_11689,N_11220,N_11213);
and U11690 (N_11690,N_11414,N_11203);
nor U11691 (N_11691,N_11233,N_11391);
nor U11692 (N_11692,N_11339,N_11030);
nand U11693 (N_11693,N_11442,N_11222);
nor U11694 (N_11694,N_11352,N_11120);
xnor U11695 (N_11695,N_11329,N_11315);
nor U11696 (N_11696,N_11153,N_11098);
nor U11697 (N_11697,N_11009,N_11155);
nand U11698 (N_11698,N_11094,N_11295);
or U11699 (N_11699,N_11379,N_11131);
nand U11700 (N_11700,N_11209,N_11495);
nand U11701 (N_11701,N_11253,N_11403);
nand U11702 (N_11702,N_11456,N_11195);
or U11703 (N_11703,N_11193,N_11363);
nand U11704 (N_11704,N_11008,N_11262);
or U11705 (N_11705,N_11272,N_11070);
xnor U11706 (N_11706,N_11388,N_11490);
and U11707 (N_11707,N_11294,N_11226);
and U11708 (N_11708,N_11328,N_11112);
and U11709 (N_11709,N_11181,N_11028);
and U11710 (N_11710,N_11102,N_11286);
and U11711 (N_11711,N_11418,N_11368);
nand U11712 (N_11712,N_11069,N_11322);
nor U11713 (N_11713,N_11411,N_11327);
or U11714 (N_11714,N_11034,N_11361);
nor U11715 (N_11715,N_11452,N_11264);
or U11716 (N_11716,N_11459,N_11166);
nor U11717 (N_11717,N_11075,N_11318);
nor U11718 (N_11718,N_11035,N_11489);
nand U11719 (N_11719,N_11137,N_11462);
or U11720 (N_11720,N_11269,N_11234);
nand U11721 (N_11721,N_11455,N_11122);
or U11722 (N_11722,N_11373,N_11428);
nand U11723 (N_11723,N_11133,N_11487);
or U11724 (N_11724,N_11062,N_11079);
or U11725 (N_11725,N_11051,N_11282);
or U11726 (N_11726,N_11216,N_11235);
nor U11727 (N_11727,N_11299,N_11439);
or U11728 (N_11728,N_11287,N_11362);
nor U11729 (N_11729,N_11007,N_11214);
or U11730 (N_11730,N_11475,N_11151);
or U11731 (N_11731,N_11419,N_11267);
and U11732 (N_11732,N_11197,N_11186);
xnor U11733 (N_11733,N_11453,N_11212);
or U11734 (N_11734,N_11446,N_11014);
nor U11735 (N_11735,N_11408,N_11468);
or U11736 (N_11736,N_11410,N_11096);
nand U11737 (N_11737,N_11479,N_11496);
nor U11738 (N_11738,N_11224,N_11174);
xor U11739 (N_11739,N_11163,N_11421);
nand U11740 (N_11740,N_11183,N_11250);
xor U11741 (N_11741,N_11289,N_11300);
nor U11742 (N_11742,N_11108,N_11417);
and U11743 (N_11743,N_11369,N_11044);
nor U11744 (N_11744,N_11144,N_11360);
nor U11745 (N_11745,N_11255,N_11381);
or U11746 (N_11746,N_11230,N_11494);
or U11747 (N_11747,N_11268,N_11476);
or U11748 (N_11748,N_11399,N_11125);
nor U11749 (N_11749,N_11437,N_11304);
and U11750 (N_11750,N_11364,N_11051);
and U11751 (N_11751,N_11179,N_11342);
nor U11752 (N_11752,N_11074,N_11033);
nor U11753 (N_11753,N_11413,N_11341);
nand U11754 (N_11754,N_11134,N_11392);
nand U11755 (N_11755,N_11136,N_11050);
nor U11756 (N_11756,N_11366,N_11220);
xnor U11757 (N_11757,N_11334,N_11331);
and U11758 (N_11758,N_11254,N_11229);
nor U11759 (N_11759,N_11097,N_11136);
nand U11760 (N_11760,N_11462,N_11102);
nor U11761 (N_11761,N_11264,N_11313);
nor U11762 (N_11762,N_11135,N_11398);
nand U11763 (N_11763,N_11192,N_11497);
nand U11764 (N_11764,N_11465,N_11037);
xnor U11765 (N_11765,N_11060,N_11342);
nor U11766 (N_11766,N_11074,N_11493);
nor U11767 (N_11767,N_11052,N_11025);
or U11768 (N_11768,N_11354,N_11425);
nor U11769 (N_11769,N_11060,N_11215);
and U11770 (N_11770,N_11194,N_11070);
nand U11771 (N_11771,N_11156,N_11176);
nand U11772 (N_11772,N_11076,N_11057);
or U11773 (N_11773,N_11318,N_11185);
and U11774 (N_11774,N_11319,N_11190);
or U11775 (N_11775,N_11358,N_11220);
nand U11776 (N_11776,N_11355,N_11411);
xor U11777 (N_11777,N_11139,N_11393);
and U11778 (N_11778,N_11463,N_11409);
nor U11779 (N_11779,N_11371,N_11495);
or U11780 (N_11780,N_11339,N_11026);
and U11781 (N_11781,N_11310,N_11218);
nor U11782 (N_11782,N_11042,N_11026);
nand U11783 (N_11783,N_11422,N_11400);
or U11784 (N_11784,N_11492,N_11266);
xnor U11785 (N_11785,N_11026,N_11124);
nand U11786 (N_11786,N_11368,N_11437);
nand U11787 (N_11787,N_11186,N_11334);
and U11788 (N_11788,N_11413,N_11201);
nand U11789 (N_11789,N_11021,N_11250);
xor U11790 (N_11790,N_11048,N_11209);
nand U11791 (N_11791,N_11224,N_11435);
xnor U11792 (N_11792,N_11136,N_11344);
and U11793 (N_11793,N_11216,N_11398);
nor U11794 (N_11794,N_11356,N_11025);
and U11795 (N_11795,N_11414,N_11261);
nand U11796 (N_11796,N_11026,N_11305);
or U11797 (N_11797,N_11485,N_11283);
nor U11798 (N_11798,N_11251,N_11276);
nand U11799 (N_11799,N_11355,N_11107);
or U11800 (N_11800,N_11229,N_11202);
nor U11801 (N_11801,N_11412,N_11351);
xor U11802 (N_11802,N_11189,N_11137);
nand U11803 (N_11803,N_11004,N_11499);
nand U11804 (N_11804,N_11272,N_11154);
and U11805 (N_11805,N_11331,N_11283);
nor U11806 (N_11806,N_11121,N_11015);
nand U11807 (N_11807,N_11061,N_11043);
nor U11808 (N_11808,N_11439,N_11324);
nand U11809 (N_11809,N_11282,N_11344);
nand U11810 (N_11810,N_11192,N_11162);
and U11811 (N_11811,N_11424,N_11348);
xnor U11812 (N_11812,N_11274,N_11087);
or U11813 (N_11813,N_11300,N_11479);
xor U11814 (N_11814,N_11310,N_11373);
and U11815 (N_11815,N_11234,N_11000);
xnor U11816 (N_11816,N_11440,N_11285);
or U11817 (N_11817,N_11304,N_11130);
nand U11818 (N_11818,N_11152,N_11360);
nor U11819 (N_11819,N_11219,N_11468);
and U11820 (N_11820,N_11182,N_11325);
or U11821 (N_11821,N_11470,N_11262);
and U11822 (N_11822,N_11282,N_11202);
xor U11823 (N_11823,N_11253,N_11330);
or U11824 (N_11824,N_11060,N_11248);
and U11825 (N_11825,N_11065,N_11156);
nor U11826 (N_11826,N_11120,N_11380);
or U11827 (N_11827,N_11443,N_11236);
nor U11828 (N_11828,N_11089,N_11482);
nor U11829 (N_11829,N_11090,N_11025);
nand U11830 (N_11830,N_11025,N_11446);
or U11831 (N_11831,N_11311,N_11257);
or U11832 (N_11832,N_11278,N_11450);
nor U11833 (N_11833,N_11122,N_11181);
nand U11834 (N_11834,N_11170,N_11262);
or U11835 (N_11835,N_11409,N_11151);
nand U11836 (N_11836,N_11081,N_11432);
nand U11837 (N_11837,N_11275,N_11313);
and U11838 (N_11838,N_11360,N_11395);
and U11839 (N_11839,N_11134,N_11373);
or U11840 (N_11840,N_11029,N_11482);
or U11841 (N_11841,N_11315,N_11469);
xor U11842 (N_11842,N_11264,N_11112);
or U11843 (N_11843,N_11406,N_11422);
and U11844 (N_11844,N_11009,N_11091);
or U11845 (N_11845,N_11355,N_11057);
or U11846 (N_11846,N_11447,N_11408);
and U11847 (N_11847,N_11302,N_11473);
xnor U11848 (N_11848,N_11374,N_11464);
nor U11849 (N_11849,N_11159,N_11199);
and U11850 (N_11850,N_11096,N_11317);
and U11851 (N_11851,N_11272,N_11101);
xor U11852 (N_11852,N_11447,N_11309);
or U11853 (N_11853,N_11261,N_11392);
nor U11854 (N_11854,N_11359,N_11254);
and U11855 (N_11855,N_11277,N_11295);
nor U11856 (N_11856,N_11187,N_11395);
nand U11857 (N_11857,N_11266,N_11182);
and U11858 (N_11858,N_11184,N_11355);
or U11859 (N_11859,N_11294,N_11490);
and U11860 (N_11860,N_11190,N_11167);
xnor U11861 (N_11861,N_11415,N_11068);
nor U11862 (N_11862,N_11383,N_11261);
nand U11863 (N_11863,N_11340,N_11327);
or U11864 (N_11864,N_11087,N_11308);
nand U11865 (N_11865,N_11433,N_11421);
nand U11866 (N_11866,N_11148,N_11296);
and U11867 (N_11867,N_11005,N_11123);
nand U11868 (N_11868,N_11413,N_11278);
or U11869 (N_11869,N_11433,N_11187);
and U11870 (N_11870,N_11040,N_11280);
and U11871 (N_11871,N_11103,N_11053);
nand U11872 (N_11872,N_11262,N_11176);
or U11873 (N_11873,N_11171,N_11314);
and U11874 (N_11874,N_11139,N_11324);
nor U11875 (N_11875,N_11173,N_11225);
nand U11876 (N_11876,N_11000,N_11308);
nand U11877 (N_11877,N_11035,N_11401);
or U11878 (N_11878,N_11291,N_11039);
nand U11879 (N_11879,N_11338,N_11441);
xor U11880 (N_11880,N_11108,N_11494);
nand U11881 (N_11881,N_11253,N_11153);
and U11882 (N_11882,N_11131,N_11325);
nand U11883 (N_11883,N_11469,N_11344);
or U11884 (N_11884,N_11210,N_11066);
nand U11885 (N_11885,N_11254,N_11181);
and U11886 (N_11886,N_11069,N_11312);
nor U11887 (N_11887,N_11104,N_11379);
nor U11888 (N_11888,N_11000,N_11084);
and U11889 (N_11889,N_11105,N_11017);
or U11890 (N_11890,N_11283,N_11483);
nand U11891 (N_11891,N_11219,N_11138);
and U11892 (N_11892,N_11089,N_11243);
and U11893 (N_11893,N_11126,N_11161);
nand U11894 (N_11894,N_11259,N_11022);
or U11895 (N_11895,N_11084,N_11150);
or U11896 (N_11896,N_11276,N_11327);
nor U11897 (N_11897,N_11446,N_11120);
nand U11898 (N_11898,N_11110,N_11216);
or U11899 (N_11899,N_11365,N_11035);
or U11900 (N_11900,N_11027,N_11036);
nand U11901 (N_11901,N_11247,N_11093);
and U11902 (N_11902,N_11251,N_11266);
nor U11903 (N_11903,N_11470,N_11398);
and U11904 (N_11904,N_11323,N_11302);
xor U11905 (N_11905,N_11454,N_11074);
nor U11906 (N_11906,N_11270,N_11034);
and U11907 (N_11907,N_11494,N_11027);
or U11908 (N_11908,N_11381,N_11343);
nor U11909 (N_11909,N_11489,N_11331);
and U11910 (N_11910,N_11440,N_11428);
and U11911 (N_11911,N_11348,N_11037);
xor U11912 (N_11912,N_11141,N_11430);
nor U11913 (N_11913,N_11420,N_11340);
and U11914 (N_11914,N_11074,N_11172);
nor U11915 (N_11915,N_11336,N_11351);
and U11916 (N_11916,N_11278,N_11053);
xor U11917 (N_11917,N_11139,N_11179);
nor U11918 (N_11918,N_11084,N_11296);
and U11919 (N_11919,N_11180,N_11196);
or U11920 (N_11920,N_11354,N_11024);
nor U11921 (N_11921,N_11383,N_11359);
and U11922 (N_11922,N_11169,N_11174);
or U11923 (N_11923,N_11179,N_11413);
nand U11924 (N_11924,N_11188,N_11220);
and U11925 (N_11925,N_11228,N_11369);
nand U11926 (N_11926,N_11171,N_11386);
and U11927 (N_11927,N_11003,N_11289);
or U11928 (N_11928,N_11261,N_11217);
nor U11929 (N_11929,N_11483,N_11014);
nand U11930 (N_11930,N_11230,N_11028);
nand U11931 (N_11931,N_11021,N_11324);
and U11932 (N_11932,N_11330,N_11388);
nand U11933 (N_11933,N_11015,N_11239);
nand U11934 (N_11934,N_11394,N_11178);
nand U11935 (N_11935,N_11475,N_11178);
or U11936 (N_11936,N_11083,N_11278);
or U11937 (N_11937,N_11294,N_11406);
or U11938 (N_11938,N_11327,N_11412);
and U11939 (N_11939,N_11140,N_11122);
and U11940 (N_11940,N_11073,N_11020);
xor U11941 (N_11941,N_11120,N_11047);
nor U11942 (N_11942,N_11113,N_11337);
xor U11943 (N_11943,N_11161,N_11438);
nor U11944 (N_11944,N_11131,N_11421);
or U11945 (N_11945,N_11235,N_11019);
nor U11946 (N_11946,N_11382,N_11394);
nor U11947 (N_11947,N_11106,N_11415);
nand U11948 (N_11948,N_11177,N_11186);
nor U11949 (N_11949,N_11430,N_11067);
nor U11950 (N_11950,N_11356,N_11267);
and U11951 (N_11951,N_11328,N_11206);
and U11952 (N_11952,N_11283,N_11346);
nand U11953 (N_11953,N_11166,N_11430);
and U11954 (N_11954,N_11234,N_11222);
or U11955 (N_11955,N_11226,N_11090);
nor U11956 (N_11956,N_11063,N_11492);
and U11957 (N_11957,N_11222,N_11260);
nand U11958 (N_11958,N_11495,N_11481);
and U11959 (N_11959,N_11403,N_11494);
and U11960 (N_11960,N_11128,N_11428);
nand U11961 (N_11961,N_11412,N_11008);
and U11962 (N_11962,N_11352,N_11142);
and U11963 (N_11963,N_11231,N_11302);
and U11964 (N_11964,N_11383,N_11070);
nand U11965 (N_11965,N_11396,N_11254);
xnor U11966 (N_11966,N_11019,N_11022);
and U11967 (N_11967,N_11039,N_11289);
nand U11968 (N_11968,N_11472,N_11446);
nor U11969 (N_11969,N_11172,N_11320);
or U11970 (N_11970,N_11125,N_11279);
xnor U11971 (N_11971,N_11459,N_11471);
and U11972 (N_11972,N_11016,N_11373);
nor U11973 (N_11973,N_11084,N_11167);
xnor U11974 (N_11974,N_11050,N_11179);
or U11975 (N_11975,N_11128,N_11449);
nor U11976 (N_11976,N_11005,N_11260);
nor U11977 (N_11977,N_11271,N_11328);
nand U11978 (N_11978,N_11483,N_11485);
nor U11979 (N_11979,N_11327,N_11011);
and U11980 (N_11980,N_11265,N_11373);
and U11981 (N_11981,N_11076,N_11233);
or U11982 (N_11982,N_11237,N_11003);
nor U11983 (N_11983,N_11233,N_11102);
nor U11984 (N_11984,N_11347,N_11182);
and U11985 (N_11985,N_11196,N_11453);
nand U11986 (N_11986,N_11369,N_11279);
nor U11987 (N_11987,N_11170,N_11233);
nor U11988 (N_11988,N_11243,N_11229);
or U11989 (N_11989,N_11497,N_11049);
nor U11990 (N_11990,N_11399,N_11160);
nor U11991 (N_11991,N_11397,N_11096);
nor U11992 (N_11992,N_11061,N_11105);
nor U11993 (N_11993,N_11430,N_11096);
or U11994 (N_11994,N_11317,N_11074);
and U11995 (N_11995,N_11119,N_11495);
or U11996 (N_11996,N_11009,N_11289);
and U11997 (N_11997,N_11341,N_11394);
nand U11998 (N_11998,N_11363,N_11287);
and U11999 (N_11999,N_11037,N_11303);
xnor U12000 (N_12000,N_11617,N_11841);
or U12001 (N_12001,N_11667,N_11625);
and U12002 (N_12002,N_11992,N_11749);
or U12003 (N_12003,N_11912,N_11803);
nand U12004 (N_12004,N_11552,N_11732);
or U12005 (N_12005,N_11895,N_11802);
xnor U12006 (N_12006,N_11850,N_11967);
nand U12007 (N_12007,N_11930,N_11631);
nor U12008 (N_12008,N_11842,N_11534);
and U12009 (N_12009,N_11518,N_11621);
xnor U12010 (N_12010,N_11938,N_11853);
or U12011 (N_12011,N_11604,N_11719);
nand U12012 (N_12012,N_11854,N_11957);
or U12013 (N_12013,N_11596,N_11996);
nand U12014 (N_12014,N_11649,N_11575);
nor U12015 (N_12015,N_11569,N_11834);
and U12016 (N_12016,N_11767,N_11917);
or U12017 (N_12017,N_11859,N_11800);
and U12018 (N_12018,N_11836,N_11861);
nand U12019 (N_12019,N_11580,N_11780);
or U12020 (N_12020,N_11556,N_11900);
and U12021 (N_12021,N_11736,N_11582);
or U12022 (N_12022,N_11528,N_11722);
xor U12023 (N_12023,N_11860,N_11981);
nor U12024 (N_12024,N_11698,N_11638);
xnor U12025 (N_12025,N_11750,N_11738);
xnor U12026 (N_12026,N_11532,N_11971);
and U12027 (N_12027,N_11546,N_11554);
or U12028 (N_12028,N_11947,N_11599);
nand U12029 (N_12029,N_11883,N_11865);
nand U12030 (N_12030,N_11718,N_11729);
nor U12031 (N_12031,N_11687,N_11831);
or U12032 (N_12032,N_11991,N_11624);
nor U12033 (N_12033,N_11796,N_11704);
or U12034 (N_12034,N_11533,N_11504);
or U12035 (N_12035,N_11550,N_11997);
nor U12036 (N_12036,N_11786,N_11821);
nand U12037 (N_12037,N_11746,N_11919);
or U12038 (N_12038,N_11560,N_11657);
nand U12039 (N_12039,N_11665,N_11968);
xor U12040 (N_12040,N_11610,N_11623);
nand U12041 (N_12041,N_11751,N_11990);
nand U12042 (N_12042,N_11586,N_11703);
or U12043 (N_12043,N_11693,N_11619);
and U12044 (N_12044,N_11949,N_11598);
nor U12045 (N_12045,N_11899,N_11512);
nor U12046 (N_12046,N_11727,N_11592);
nand U12047 (N_12047,N_11896,N_11911);
or U12048 (N_12048,N_11568,N_11804);
or U12049 (N_12049,N_11921,N_11678);
and U12050 (N_12050,N_11830,N_11764);
and U12051 (N_12051,N_11634,N_11505);
and U12052 (N_12052,N_11715,N_11956);
or U12053 (N_12053,N_11887,N_11612);
or U12054 (N_12054,N_11812,N_11522);
nand U12055 (N_12055,N_11843,N_11607);
nor U12056 (N_12056,N_11557,N_11666);
nor U12057 (N_12057,N_11794,N_11513);
nand U12058 (N_12058,N_11579,N_11711);
nor U12059 (N_12059,N_11618,N_11869);
or U12060 (N_12060,N_11507,N_11837);
or U12061 (N_12061,N_11888,N_11691);
nand U12062 (N_12062,N_11753,N_11823);
nand U12063 (N_12063,N_11959,N_11614);
or U12064 (N_12064,N_11651,N_11923);
nand U12065 (N_12065,N_11570,N_11526);
and U12066 (N_12066,N_11889,N_11885);
or U12067 (N_12067,N_11673,N_11731);
nand U12068 (N_12068,N_11521,N_11517);
and U12069 (N_12069,N_11960,N_11671);
nand U12070 (N_12070,N_11536,N_11728);
or U12071 (N_12071,N_11725,N_11953);
nor U12072 (N_12072,N_11726,N_11925);
nand U12073 (N_12073,N_11782,N_11581);
xnor U12074 (N_12074,N_11945,N_11656);
or U12075 (N_12075,N_11511,N_11734);
xnor U12076 (N_12076,N_11655,N_11541);
nor U12077 (N_12077,N_11571,N_11892);
and U12078 (N_12078,N_11844,N_11700);
nor U12079 (N_12079,N_11993,N_11578);
or U12080 (N_12080,N_11871,N_11752);
nand U12081 (N_12081,N_11819,N_11975);
and U12082 (N_12082,N_11766,N_11890);
or U12083 (N_12083,N_11792,N_11721);
and U12084 (N_12084,N_11832,N_11606);
nor U12085 (N_12085,N_11774,N_11771);
and U12086 (N_12086,N_11778,N_11998);
nor U12087 (N_12087,N_11795,N_11564);
xor U12088 (N_12088,N_11882,N_11509);
and U12089 (N_12089,N_11745,N_11577);
nand U12090 (N_12090,N_11591,N_11983);
and U12091 (N_12091,N_11547,N_11988);
and U12092 (N_12092,N_11523,N_11926);
nor U12093 (N_12093,N_11877,N_11660);
and U12094 (N_12094,N_11531,N_11668);
or U12095 (N_12095,N_11840,N_11815);
nor U12096 (N_12096,N_11820,N_11540);
xnor U12097 (N_12097,N_11807,N_11519);
nor U12098 (N_12098,N_11626,N_11781);
nand U12099 (N_12099,N_11924,N_11609);
or U12100 (N_12100,N_11566,N_11742);
nor U12101 (N_12101,N_11783,N_11633);
and U12102 (N_12102,N_11894,N_11595);
or U12103 (N_12103,N_11966,N_11674);
nand U12104 (N_12104,N_11669,N_11969);
and U12105 (N_12105,N_11805,N_11797);
nor U12106 (N_12106,N_11791,N_11709);
or U12107 (N_12107,N_11973,N_11948);
nor U12108 (N_12108,N_11628,N_11737);
or U12109 (N_12109,N_11817,N_11874);
nor U12110 (N_12110,N_11645,N_11688);
nand U12111 (N_12111,N_11601,N_11905);
nor U12112 (N_12112,N_11935,N_11961);
nand U12113 (N_12113,N_11701,N_11561);
and U12114 (N_12114,N_11955,N_11733);
nand U12115 (N_12115,N_11931,N_11822);
or U12116 (N_12116,N_11835,N_11755);
nor U12117 (N_12117,N_11567,N_11613);
nor U12118 (N_12118,N_11872,N_11697);
and U12119 (N_12119,N_11989,N_11588);
or U12120 (N_12120,N_11999,N_11644);
nand U12121 (N_12121,N_11724,N_11681);
nand U12122 (N_12122,N_11583,N_11629);
and U12123 (N_12123,N_11806,N_11677);
or U12124 (N_12124,N_11827,N_11542);
and U12125 (N_12125,N_11952,N_11933);
nand U12126 (N_12126,N_11664,N_11984);
xor U12127 (N_12127,N_11713,N_11867);
nor U12128 (N_12128,N_11868,N_11590);
nor U12129 (N_12129,N_11864,N_11809);
xor U12130 (N_12130,N_11574,N_11873);
nor U12131 (N_12131,N_11826,N_11858);
and U12132 (N_12132,N_11608,N_11611);
xnor U12133 (N_12133,N_11941,N_11902);
xor U12134 (N_12134,N_11603,N_11587);
or U12135 (N_12135,N_11863,N_11950);
xor U12136 (N_12136,N_11762,N_11602);
xnor U12137 (N_12137,N_11707,N_11648);
nor U12138 (N_12138,N_11670,N_11879);
nand U12139 (N_12139,N_11849,N_11712);
or U12140 (N_12140,N_11662,N_11916);
nand U12141 (N_12141,N_11747,N_11964);
or U12142 (N_12142,N_11686,N_11636);
nor U12143 (N_12143,N_11754,N_11980);
nand U12144 (N_12144,N_11600,N_11940);
nor U12145 (N_12145,N_11986,N_11920);
or U12146 (N_12146,N_11907,N_11936);
or U12147 (N_12147,N_11741,N_11829);
and U12148 (N_12148,N_11876,N_11878);
or U12149 (N_12149,N_11808,N_11543);
nor U12150 (N_12150,N_11683,N_11685);
nand U12151 (N_12151,N_11520,N_11695);
nor U12152 (N_12152,N_11788,N_11503);
nand U12153 (N_12153,N_11811,N_11632);
and U12154 (N_12154,N_11769,N_11654);
xor U12155 (N_12155,N_11548,N_11994);
and U12156 (N_12156,N_11816,N_11740);
nand U12157 (N_12157,N_11694,N_11846);
and U12158 (N_12158,N_11772,N_11944);
nand U12159 (N_12159,N_11759,N_11530);
nor U12160 (N_12160,N_11717,N_11951);
and U12161 (N_12161,N_11524,N_11965);
nor U12162 (N_12162,N_11775,N_11810);
and U12163 (N_12163,N_11692,N_11615);
nor U12164 (N_12164,N_11875,N_11915);
and U12165 (N_12165,N_11928,N_11539);
and U12166 (N_12166,N_11563,N_11551);
nand U12167 (N_12167,N_11708,N_11801);
and U12168 (N_12168,N_11777,N_11906);
nor U12169 (N_12169,N_11757,N_11855);
and U12170 (N_12170,N_11506,N_11979);
and U12171 (N_12171,N_11839,N_11977);
nand U12172 (N_12172,N_11502,N_11514);
nor U12173 (N_12173,N_11779,N_11643);
or U12174 (N_12174,N_11572,N_11982);
nand U12175 (N_12175,N_11647,N_11642);
or U12176 (N_12176,N_11559,N_11663);
nor U12177 (N_12177,N_11659,N_11639);
or U12178 (N_12178,N_11658,N_11743);
nor U12179 (N_12179,N_11908,N_11787);
or U12180 (N_12180,N_11690,N_11881);
or U12181 (N_12181,N_11825,N_11584);
and U12182 (N_12182,N_11641,N_11635);
or U12183 (N_12183,N_11773,N_11646);
nor U12184 (N_12184,N_11833,N_11744);
and U12185 (N_12185,N_11937,N_11785);
or U12186 (N_12186,N_11963,N_11913);
nor U12187 (N_12187,N_11680,N_11675);
nand U12188 (N_12188,N_11620,N_11880);
xor U12189 (N_12189,N_11515,N_11943);
xor U12190 (N_12190,N_11893,N_11593);
nand U12191 (N_12191,N_11653,N_11932);
nor U12192 (N_12192,N_11838,N_11866);
nor U12193 (N_12193,N_11616,N_11918);
or U12194 (N_12194,N_11553,N_11942);
and U12195 (N_12195,N_11758,N_11974);
nand U12196 (N_12196,N_11723,N_11508);
nor U12197 (N_12197,N_11735,N_11813);
or U12198 (N_12198,N_11985,N_11538);
nand U12199 (N_12199,N_11934,N_11886);
and U12200 (N_12200,N_11954,N_11682);
xor U12201 (N_12201,N_11793,N_11661);
and U12202 (N_12202,N_11760,N_11765);
and U12203 (N_12203,N_11544,N_11776);
xnor U12204 (N_12204,N_11770,N_11558);
and U12205 (N_12205,N_11995,N_11699);
or U12206 (N_12206,N_11976,N_11676);
and U12207 (N_12207,N_11939,N_11914);
xnor U12208 (N_12208,N_11897,N_11555);
nor U12209 (N_12209,N_11904,N_11851);
or U12210 (N_12210,N_11857,N_11500);
and U12211 (N_12211,N_11640,N_11562);
and U12212 (N_12212,N_11545,N_11525);
or U12213 (N_12213,N_11510,N_11799);
nor U12214 (N_12214,N_11501,N_11739);
and U12215 (N_12215,N_11627,N_11637);
and U12216 (N_12216,N_11763,N_11784);
and U12217 (N_12217,N_11565,N_11852);
and U12218 (N_12218,N_11720,N_11605);
and U12219 (N_12219,N_11824,N_11946);
and U12220 (N_12220,N_11535,N_11798);
nand U12221 (N_12221,N_11756,N_11705);
nor U12222 (N_12222,N_11856,N_11597);
or U12223 (N_12223,N_11845,N_11847);
nand U12224 (N_12224,N_11684,N_11891);
nand U12225 (N_12225,N_11630,N_11573);
nand U12226 (N_12226,N_11702,N_11922);
and U12227 (N_12227,N_11650,N_11909);
nand U12228 (N_12228,N_11828,N_11689);
xnor U12229 (N_12229,N_11958,N_11818);
nor U12230 (N_12230,N_11730,N_11903);
nand U12231 (N_12231,N_11790,N_11972);
and U12232 (N_12232,N_11516,N_11927);
xor U12233 (N_12233,N_11706,N_11537);
and U12234 (N_12234,N_11814,N_11672);
xnor U12235 (N_12235,N_11696,N_11901);
nor U12236 (N_12236,N_11848,N_11962);
xor U12237 (N_12237,N_11622,N_11527);
or U12238 (N_12238,N_11929,N_11652);
and U12239 (N_12239,N_11870,N_11594);
nor U12240 (N_12240,N_11748,N_11549);
nand U12241 (N_12241,N_11716,N_11679);
and U12242 (N_12242,N_11789,N_11714);
nor U12243 (N_12243,N_11585,N_11576);
nor U12244 (N_12244,N_11898,N_11978);
nor U12245 (N_12245,N_11710,N_11589);
and U12246 (N_12246,N_11970,N_11862);
and U12247 (N_12247,N_11768,N_11761);
and U12248 (N_12248,N_11910,N_11529);
nand U12249 (N_12249,N_11884,N_11987);
nand U12250 (N_12250,N_11803,N_11659);
and U12251 (N_12251,N_11963,N_11861);
nand U12252 (N_12252,N_11865,N_11564);
nor U12253 (N_12253,N_11558,N_11848);
nand U12254 (N_12254,N_11875,N_11942);
or U12255 (N_12255,N_11502,N_11704);
nor U12256 (N_12256,N_11647,N_11985);
or U12257 (N_12257,N_11806,N_11505);
and U12258 (N_12258,N_11982,N_11788);
nor U12259 (N_12259,N_11858,N_11959);
xor U12260 (N_12260,N_11845,N_11592);
xnor U12261 (N_12261,N_11590,N_11835);
nor U12262 (N_12262,N_11854,N_11604);
and U12263 (N_12263,N_11861,N_11704);
and U12264 (N_12264,N_11705,N_11695);
nor U12265 (N_12265,N_11928,N_11624);
nand U12266 (N_12266,N_11641,N_11678);
nor U12267 (N_12267,N_11622,N_11598);
and U12268 (N_12268,N_11910,N_11641);
nand U12269 (N_12269,N_11814,N_11832);
and U12270 (N_12270,N_11648,N_11858);
nand U12271 (N_12271,N_11552,N_11593);
nor U12272 (N_12272,N_11511,N_11943);
nand U12273 (N_12273,N_11842,N_11699);
nand U12274 (N_12274,N_11819,N_11750);
and U12275 (N_12275,N_11949,N_11516);
nand U12276 (N_12276,N_11714,N_11639);
nor U12277 (N_12277,N_11873,N_11960);
nor U12278 (N_12278,N_11872,N_11727);
or U12279 (N_12279,N_11665,N_11789);
nor U12280 (N_12280,N_11702,N_11872);
and U12281 (N_12281,N_11645,N_11886);
and U12282 (N_12282,N_11790,N_11747);
nand U12283 (N_12283,N_11878,N_11983);
nor U12284 (N_12284,N_11954,N_11511);
or U12285 (N_12285,N_11543,N_11970);
nor U12286 (N_12286,N_11830,N_11745);
or U12287 (N_12287,N_11905,N_11880);
xor U12288 (N_12288,N_11866,N_11519);
or U12289 (N_12289,N_11513,N_11774);
nand U12290 (N_12290,N_11968,N_11523);
xnor U12291 (N_12291,N_11653,N_11771);
nor U12292 (N_12292,N_11805,N_11845);
nor U12293 (N_12293,N_11872,N_11593);
or U12294 (N_12294,N_11755,N_11504);
and U12295 (N_12295,N_11952,N_11616);
nand U12296 (N_12296,N_11593,N_11949);
or U12297 (N_12297,N_11775,N_11883);
nor U12298 (N_12298,N_11734,N_11698);
or U12299 (N_12299,N_11656,N_11535);
nand U12300 (N_12300,N_11880,N_11629);
and U12301 (N_12301,N_11944,N_11745);
nand U12302 (N_12302,N_11825,N_11520);
and U12303 (N_12303,N_11908,N_11715);
nand U12304 (N_12304,N_11503,N_11681);
xnor U12305 (N_12305,N_11713,N_11674);
nand U12306 (N_12306,N_11747,N_11814);
or U12307 (N_12307,N_11782,N_11566);
nand U12308 (N_12308,N_11532,N_11686);
or U12309 (N_12309,N_11805,N_11640);
or U12310 (N_12310,N_11790,N_11950);
nor U12311 (N_12311,N_11650,N_11787);
or U12312 (N_12312,N_11771,N_11911);
nor U12313 (N_12313,N_11961,N_11781);
or U12314 (N_12314,N_11749,N_11881);
or U12315 (N_12315,N_11634,N_11614);
nor U12316 (N_12316,N_11680,N_11837);
and U12317 (N_12317,N_11969,N_11505);
and U12318 (N_12318,N_11794,N_11752);
or U12319 (N_12319,N_11873,N_11613);
and U12320 (N_12320,N_11735,N_11728);
xnor U12321 (N_12321,N_11749,N_11936);
and U12322 (N_12322,N_11769,N_11799);
xor U12323 (N_12323,N_11885,N_11778);
nor U12324 (N_12324,N_11976,N_11576);
nor U12325 (N_12325,N_11594,N_11929);
nand U12326 (N_12326,N_11975,N_11988);
nand U12327 (N_12327,N_11525,N_11728);
or U12328 (N_12328,N_11975,N_11767);
or U12329 (N_12329,N_11922,N_11712);
nand U12330 (N_12330,N_11743,N_11536);
nor U12331 (N_12331,N_11999,N_11582);
or U12332 (N_12332,N_11572,N_11503);
and U12333 (N_12333,N_11885,N_11802);
nand U12334 (N_12334,N_11663,N_11596);
nor U12335 (N_12335,N_11516,N_11710);
nor U12336 (N_12336,N_11678,N_11662);
nor U12337 (N_12337,N_11863,N_11737);
nor U12338 (N_12338,N_11743,N_11561);
nor U12339 (N_12339,N_11530,N_11798);
nor U12340 (N_12340,N_11868,N_11646);
xnor U12341 (N_12341,N_11622,N_11575);
and U12342 (N_12342,N_11779,N_11909);
nand U12343 (N_12343,N_11887,N_11607);
nor U12344 (N_12344,N_11564,N_11765);
and U12345 (N_12345,N_11890,N_11915);
and U12346 (N_12346,N_11915,N_11821);
or U12347 (N_12347,N_11949,N_11500);
nand U12348 (N_12348,N_11878,N_11783);
or U12349 (N_12349,N_11777,N_11685);
xnor U12350 (N_12350,N_11502,N_11716);
nand U12351 (N_12351,N_11575,N_11736);
or U12352 (N_12352,N_11502,N_11927);
nand U12353 (N_12353,N_11549,N_11798);
or U12354 (N_12354,N_11831,N_11664);
nor U12355 (N_12355,N_11774,N_11757);
and U12356 (N_12356,N_11994,N_11646);
xor U12357 (N_12357,N_11559,N_11809);
and U12358 (N_12358,N_11963,N_11828);
or U12359 (N_12359,N_11811,N_11679);
nand U12360 (N_12360,N_11823,N_11946);
nand U12361 (N_12361,N_11910,N_11915);
xnor U12362 (N_12362,N_11586,N_11743);
or U12363 (N_12363,N_11577,N_11919);
nor U12364 (N_12364,N_11838,N_11930);
and U12365 (N_12365,N_11581,N_11537);
and U12366 (N_12366,N_11907,N_11640);
nor U12367 (N_12367,N_11779,N_11846);
xnor U12368 (N_12368,N_11972,N_11603);
or U12369 (N_12369,N_11976,N_11794);
and U12370 (N_12370,N_11570,N_11899);
nor U12371 (N_12371,N_11916,N_11571);
nand U12372 (N_12372,N_11958,N_11799);
nor U12373 (N_12373,N_11716,N_11943);
nand U12374 (N_12374,N_11674,N_11560);
nor U12375 (N_12375,N_11891,N_11597);
nor U12376 (N_12376,N_11552,N_11611);
nor U12377 (N_12377,N_11521,N_11962);
nand U12378 (N_12378,N_11602,N_11538);
nand U12379 (N_12379,N_11821,N_11911);
or U12380 (N_12380,N_11806,N_11635);
or U12381 (N_12381,N_11505,N_11795);
and U12382 (N_12382,N_11994,N_11711);
xnor U12383 (N_12383,N_11700,N_11861);
and U12384 (N_12384,N_11956,N_11643);
nand U12385 (N_12385,N_11977,N_11824);
and U12386 (N_12386,N_11805,N_11556);
or U12387 (N_12387,N_11520,N_11543);
nor U12388 (N_12388,N_11848,N_11878);
xor U12389 (N_12389,N_11691,N_11950);
and U12390 (N_12390,N_11965,N_11511);
and U12391 (N_12391,N_11706,N_11623);
and U12392 (N_12392,N_11669,N_11657);
nand U12393 (N_12393,N_11547,N_11809);
and U12394 (N_12394,N_11812,N_11913);
and U12395 (N_12395,N_11705,N_11575);
nand U12396 (N_12396,N_11930,N_11829);
nand U12397 (N_12397,N_11516,N_11981);
or U12398 (N_12398,N_11520,N_11705);
or U12399 (N_12399,N_11567,N_11576);
or U12400 (N_12400,N_11800,N_11915);
or U12401 (N_12401,N_11875,N_11920);
xor U12402 (N_12402,N_11562,N_11768);
nand U12403 (N_12403,N_11882,N_11619);
nand U12404 (N_12404,N_11869,N_11826);
and U12405 (N_12405,N_11717,N_11576);
nand U12406 (N_12406,N_11583,N_11607);
or U12407 (N_12407,N_11861,N_11993);
or U12408 (N_12408,N_11913,N_11507);
xor U12409 (N_12409,N_11544,N_11572);
or U12410 (N_12410,N_11970,N_11653);
or U12411 (N_12411,N_11901,N_11695);
nor U12412 (N_12412,N_11693,N_11584);
and U12413 (N_12413,N_11834,N_11768);
or U12414 (N_12414,N_11573,N_11964);
nor U12415 (N_12415,N_11921,N_11884);
nor U12416 (N_12416,N_11618,N_11613);
nand U12417 (N_12417,N_11651,N_11786);
nand U12418 (N_12418,N_11593,N_11690);
and U12419 (N_12419,N_11997,N_11545);
or U12420 (N_12420,N_11642,N_11784);
and U12421 (N_12421,N_11732,N_11682);
or U12422 (N_12422,N_11986,N_11741);
xnor U12423 (N_12423,N_11654,N_11563);
nor U12424 (N_12424,N_11725,N_11537);
and U12425 (N_12425,N_11551,N_11627);
nor U12426 (N_12426,N_11979,N_11988);
and U12427 (N_12427,N_11871,N_11933);
and U12428 (N_12428,N_11505,N_11679);
and U12429 (N_12429,N_11537,N_11853);
nand U12430 (N_12430,N_11756,N_11695);
or U12431 (N_12431,N_11941,N_11619);
nand U12432 (N_12432,N_11888,N_11935);
and U12433 (N_12433,N_11685,N_11673);
nand U12434 (N_12434,N_11893,N_11656);
or U12435 (N_12435,N_11584,N_11638);
xnor U12436 (N_12436,N_11786,N_11658);
and U12437 (N_12437,N_11652,N_11887);
and U12438 (N_12438,N_11855,N_11762);
and U12439 (N_12439,N_11824,N_11781);
and U12440 (N_12440,N_11700,N_11785);
nor U12441 (N_12441,N_11830,N_11797);
and U12442 (N_12442,N_11633,N_11665);
or U12443 (N_12443,N_11956,N_11879);
xor U12444 (N_12444,N_11600,N_11584);
and U12445 (N_12445,N_11626,N_11663);
and U12446 (N_12446,N_11613,N_11672);
or U12447 (N_12447,N_11760,N_11856);
nand U12448 (N_12448,N_11675,N_11765);
nand U12449 (N_12449,N_11656,N_11929);
nor U12450 (N_12450,N_11841,N_11964);
nand U12451 (N_12451,N_11874,N_11764);
xor U12452 (N_12452,N_11985,N_11749);
nor U12453 (N_12453,N_11525,N_11805);
or U12454 (N_12454,N_11836,N_11931);
nand U12455 (N_12455,N_11702,N_11795);
and U12456 (N_12456,N_11841,N_11630);
or U12457 (N_12457,N_11943,N_11772);
nor U12458 (N_12458,N_11538,N_11580);
xnor U12459 (N_12459,N_11705,N_11798);
nand U12460 (N_12460,N_11912,N_11737);
or U12461 (N_12461,N_11591,N_11896);
or U12462 (N_12462,N_11647,N_11825);
nor U12463 (N_12463,N_11743,N_11901);
or U12464 (N_12464,N_11990,N_11504);
nor U12465 (N_12465,N_11853,N_11745);
xor U12466 (N_12466,N_11629,N_11916);
and U12467 (N_12467,N_11810,N_11619);
xor U12468 (N_12468,N_11510,N_11953);
nand U12469 (N_12469,N_11615,N_11661);
and U12470 (N_12470,N_11928,N_11603);
and U12471 (N_12471,N_11654,N_11824);
nor U12472 (N_12472,N_11734,N_11897);
or U12473 (N_12473,N_11715,N_11841);
nand U12474 (N_12474,N_11941,N_11710);
and U12475 (N_12475,N_11642,N_11936);
or U12476 (N_12476,N_11919,N_11758);
or U12477 (N_12477,N_11699,N_11879);
or U12478 (N_12478,N_11807,N_11774);
and U12479 (N_12479,N_11658,N_11879);
and U12480 (N_12480,N_11527,N_11941);
nor U12481 (N_12481,N_11748,N_11834);
nor U12482 (N_12482,N_11901,N_11821);
nand U12483 (N_12483,N_11620,N_11518);
nand U12484 (N_12484,N_11688,N_11550);
and U12485 (N_12485,N_11639,N_11957);
or U12486 (N_12486,N_11509,N_11597);
or U12487 (N_12487,N_11547,N_11735);
nor U12488 (N_12488,N_11978,N_11891);
xor U12489 (N_12489,N_11955,N_11907);
or U12490 (N_12490,N_11810,N_11639);
and U12491 (N_12491,N_11907,N_11853);
xnor U12492 (N_12492,N_11934,N_11772);
and U12493 (N_12493,N_11871,N_11658);
nand U12494 (N_12494,N_11557,N_11562);
nand U12495 (N_12495,N_11724,N_11686);
and U12496 (N_12496,N_11594,N_11873);
or U12497 (N_12497,N_11959,N_11532);
or U12498 (N_12498,N_11779,N_11718);
nor U12499 (N_12499,N_11941,N_11722);
nand U12500 (N_12500,N_12387,N_12201);
nor U12501 (N_12501,N_12014,N_12373);
nor U12502 (N_12502,N_12414,N_12382);
and U12503 (N_12503,N_12081,N_12312);
and U12504 (N_12504,N_12249,N_12483);
or U12505 (N_12505,N_12032,N_12429);
xnor U12506 (N_12506,N_12430,N_12401);
and U12507 (N_12507,N_12191,N_12180);
and U12508 (N_12508,N_12303,N_12299);
nand U12509 (N_12509,N_12346,N_12105);
and U12510 (N_12510,N_12051,N_12072);
xnor U12511 (N_12511,N_12017,N_12104);
nand U12512 (N_12512,N_12297,N_12086);
xor U12513 (N_12513,N_12471,N_12124);
xor U12514 (N_12514,N_12481,N_12210);
or U12515 (N_12515,N_12021,N_12093);
nand U12516 (N_12516,N_12155,N_12234);
and U12517 (N_12517,N_12398,N_12241);
or U12518 (N_12518,N_12478,N_12357);
or U12519 (N_12519,N_12018,N_12031);
nand U12520 (N_12520,N_12140,N_12144);
and U12521 (N_12521,N_12150,N_12121);
or U12522 (N_12522,N_12141,N_12385);
nand U12523 (N_12523,N_12146,N_12226);
and U12524 (N_12524,N_12493,N_12045);
nand U12525 (N_12525,N_12125,N_12294);
or U12526 (N_12526,N_12276,N_12351);
nor U12527 (N_12527,N_12211,N_12216);
nor U12528 (N_12528,N_12244,N_12286);
or U12529 (N_12529,N_12280,N_12085);
and U12530 (N_12530,N_12394,N_12477);
or U12531 (N_12531,N_12332,N_12036);
and U12532 (N_12532,N_12412,N_12274);
nand U12533 (N_12533,N_12368,N_12209);
and U12534 (N_12534,N_12247,N_12127);
or U12535 (N_12535,N_12112,N_12050);
nand U12536 (N_12536,N_12006,N_12488);
nand U12537 (N_12537,N_12116,N_12271);
and U12538 (N_12538,N_12070,N_12333);
nor U12539 (N_12539,N_12099,N_12170);
or U12540 (N_12540,N_12298,N_12413);
nand U12541 (N_12541,N_12101,N_12074);
and U12542 (N_12542,N_12388,N_12270);
nand U12543 (N_12543,N_12067,N_12463);
nand U12544 (N_12544,N_12331,N_12371);
xor U12545 (N_12545,N_12453,N_12419);
and U12546 (N_12546,N_12464,N_12143);
or U12547 (N_12547,N_12490,N_12049);
nor U12548 (N_12548,N_12119,N_12054);
nor U12549 (N_12549,N_12120,N_12428);
or U12550 (N_12550,N_12289,N_12082);
nor U12551 (N_12551,N_12160,N_12039);
or U12552 (N_12552,N_12439,N_12052);
nand U12553 (N_12553,N_12433,N_12220);
nor U12554 (N_12554,N_12327,N_12290);
nor U12555 (N_12555,N_12392,N_12041);
xnor U12556 (N_12556,N_12077,N_12405);
xnor U12557 (N_12557,N_12254,N_12213);
nand U12558 (N_12558,N_12171,N_12076);
nand U12559 (N_12559,N_12193,N_12376);
and U12560 (N_12560,N_12059,N_12393);
nand U12561 (N_12561,N_12055,N_12118);
nand U12562 (N_12562,N_12470,N_12338);
or U12563 (N_12563,N_12126,N_12094);
nor U12564 (N_12564,N_12476,N_12361);
or U12565 (N_12565,N_12027,N_12060);
xnor U12566 (N_12566,N_12309,N_12485);
nor U12567 (N_12567,N_12010,N_12396);
nand U12568 (N_12568,N_12240,N_12168);
and U12569 (N_12569,N_12421,N_12314);
xor U12570 (N_12570,N_12305,N_12109);
nor U12571 (N_12571,N_12442,N_12108);
and U12572 (N_12572,N_12250,N_12167);
nand U12573 (N_12573,N_12395,N_12265);
nor U12574 (N_12574,N_12029,N_12106);
nor U12575 (N_12575,N_12472,N_12165);
xor U12576 (N_12576,N_12403,N_12400);
and U12577 (N_12577,N_12443,N_12080);
and U12578 (N_12578,N_12186,N_12353);
and U12579 (N_12579,N_12110,N_12135);
nor U12580 (N_12580,N_12315,N_12425);
and U12581 (N_12581,N_12087,N_12426);
nor U12582 (N_12582,N_12195,N_12480);
nor U12583 (N_12583,N_12179,N_12479);
nand U12584 (N_12584,N_12284,N_12321);
nand U12585 (N_12585,N_12451,N_12206);
and U12586 (N_12586,N_12131,N_12199);
or U12587 (N_12587,N_12374,N_12307);
nand U12588 (N_12588,N_12411,N_12098);
and U12589 (N_12589,N_12103,N_12358);
or U12590 (N_12590,N_12044,N_12448);
and U12591 (N_12591,N_12416,N_12016);
nor U12592 (N_12592,N_12172,N_12013);
and U12593 (N_12593,N_12293,N_12158);
and U12594 (N_12594,N_12200,N_12117);
nand U12595 (N_12595,N_12266,N_12350);
or U12596 (N_12596,N_12415,N_12450);
xor U12597 (N_12597,N_12064,N_12020);
and U12598 (N_12598,N_12324,N_12486);
nand U12599 (N_12599,N_12441,N_12012);
nand U12600 (N_12600,N_12042,N_12408);
and U12601 (N_12601,N_12092,N_12164);
or U12602 (N_12602,N_12188,N_12183);
nand U12603 (N_12603,N_12114,N_12422);
nor U12604 (N_12604,N_12409,N_12192);
nor U12605 (N_12605,N_12467,N_12406);
nor U12606 (N_12606,N_12278,N_12037);
nand U12607 (N_12607,N_12009,N_12214);
or U12608 (N_12608,N_12362,N_12053);
nor U12609 (N_12609,N_12024,N_12465);
nor U12610 (N_12610,N_12107,N_12456);
and U12611 (N_12611,N_12455,N_12198);
or U12612 (N_12612,N_12402,N_12236);
nor U12613 (N_12613,N_12378,N_12469);
and U12614 (N_12614,N_12487,N_12377);
or U12615 (N_12615,N_12022,N_12304);
or U12616 (N_12616,N_12275,N_12034);
nand U12617 (N_12617,N_12475,N_12356);
and U12618 (N_12618,N_12129,N_12173);
nand U12619 (N_12619,N_12218,N_12311);
nor U12620 (N_12620,N_12253,N_12097);
or U12621 (N_12621,N_12499,N_12461);
nor U12622 (N_12622,N_12445,N_12277);
or U12623 (N_12623,N_12313,N_12197);
and U12624 (N_12624,N_12427,N_12288);
or U12625 (N_12625,N_12019,N_12318);
nand U12626 (N_12626,N_12468,N_12420);
or U12627 (N_12627,N_12440,N_12317);
nand U12628 (N_12628,N_12454,N_12163);
nand U12629 (N_12629,N_12256,N_12264);
and U12630 (N_12630,N_12190,N_12056);
nor U12631 (N_12631,N_12496,N_12359);
xnor U12632 (N_12632,N_12484,N_12375);
nand U12633 (N_12633,N_12306,N_12033);
and U12634 (N_12634,N_12437,N_12344);
and U12635 (N_12635,N_12134,N_12147);
nor U12636 (N_12636,N_12272,N_12301);
nor U12637 (N_12637,N_12452,N_12223);
and U12638 (N_12638,N_12038,N_12189);
nand U12639 (N_12639,N_12203,N_12279);
and U12640 (N_12640,N_12404,N_12159);
nand U12641 (N_12641,N_12245,N_12048);
and U12642 (N_12642,N_12025,N_12058);
nor U12643 (N_12643,N_12026,N_12242);
and U12644 (N_12644,N_12326,N_12295);
and U12645 (N_12645,N_12258,N_12418);
and U12646 (N_12646,N_12007,N_12153);
nor U12647 (N_12647,N_12133,N_12340);
nand U12648 (N_12648,N_12325,N_12262);
nor U12649 (N_12649,N_12174,N_12004);
nand U12650 (N_12650,N_12345,N_12498);
and U12651 (N_12651,N_12196,N_12187);
nand U12652 (N_12652,N_12023,N_12335);
or U12653 (N_12653,N_12460,N_12095);
or U12654 (N_12654,N_12128,N_12136);
or U12655 (N_12655,N_12002,N_12255);
and U12656 (N_12656,N_12384,N_12177);
or U12657 (N_12657,N_12156,N_12008);
nand U12658 (N_12658,N_12367,N_12380);
and U12659 (N_12659,N_12111,N_12123);
nand U12660 (N_12660,N_12369,N_12003);
and U12661 (N_12661,N_12248,N_12075);
and U12662 (N_12662,N_12228,N_12497);
nand U12663 (N_12663,N_12329,N_12212);
nand U12664 (N_12664,N_12492,N_12181);
or U12665 (N_12665,N_12142,N_12148);
nand U12666 (N_12666,N_12166,N_12161);
and U12667 (N_12667,N_12348,N_12071);
or U12668 (N_12668,N_12005,N_12176);
and U12669 (N_12669,N_12407,N_12078);
xnor U12670 (N_12670,N_12185,N_12063);
or U12671 (N_12671,N_12444,N_12417);
nor U12672 (N_12672,N_12068,N_12390);
nor U12673 (N_12673,N_12115,N_12316);
nor U12674 (N_12674,N_12269,N_12339);
and U12675 (N_12675,N_12083,N_12438);
nand U12676 (N_12676,N_12035,N_12202);
nor U12677 (N_12677,N_12391,N_12231);
nor U12678 (N_12678,N_12221,N_12222);
nor U12679 (N_12679,N_12084,N_12364);
nand U12680 (N_12680,N_12379,N_12239);
nor U12681 (N_12681,N_12225,N_12273);
nand U12682 (N_12682,N_12073,N_12372);
or U12683 (N_12683,N_12219,N_12491);
nor U12684 (N_12684,N_12137,N_12232);
or U12685 (N_12685,N_12096,N_12263);
and U12686 (N_12686,N_12132,N_12043);
or U12687 (N_12687,N_12113,N_12320);
and U12688 (N_12688,N_12291,N_12061);
nand U12689 (N_12689,N_12162,N_12046);
and U12690 (N_12690,N_12154,N_12296);
and U12691 (N_12691,N_12138,N_12381);
or U12692 (N_12692,N_12057,N_12302);
xor U12693 (N_12693,N_12355,N_12423);
nand U12694 (N_12694,N_12252,N_12238);
and U12695 (N_12695,N_12000,N_12473);
or U12696 (N_12696,N_12011,N_12459);
xor U12697 (N_12697,N_12462,N_12178);
and U12698 (N_12698,N_12466,N_12091);
and U12699 (N_12699,N_12065,N_12474);
nand U12700 (N_12700,N_12431,N_12336);
and U12701 (N_12701,N_12435,N_12233);
and U12702 (N_12702,N_12494,N_12410);
or U12703 (N_12703,N_12334,N_12360);
and U12704 (N_12704,N_12287,N_12323);
or U12705 (N_12705,N_12251,N_12341);
and U12706 (N_12706,N_12157,N_12182);
nand U12707 (N_12707,N_12139,N_12235);
and U12708 (N_12708,N_12363,N_12282);
and U12709 (N_12709,N_12066,N_12285);
and U12710 (N_12710,N_12204,N_12217);
nor U12711 (N_12711,N_12447,N_12227);
or U12712 (N_12712,N_12261,N_12489);
nor U12713 (N_12713,N_12366,N_12328);
and U12714 (N_12714,N_12268,N_12207);
and U12715 (N_12715,N_12257,N_12322);
nor U12716 (N_12716,N_12215,N_12370);
nor U12717 (N_12717,N_12386,N_12337);
xnor U12718 (N_12718,N_12015,N_12436);
and U12719 (N_12719,N_12399,N_12365);
or U12720 (N_12720,N_12281,N_12090);
or U12721 (N_12721,N_12246,N_12458);
and U12722 (N_12722,N_12102,N_12040);
nand U12723 (N_12723,N_12342,N_12028);
and U12724 (N_12724,N_12089,N_12260);
nand U12725 (N_12725,N_12047,N_12319);
nand U12726 (N_12726,N_12308,N_12434);
nor U12727 (N_12727,N_12424,N_12152);
nor U12728 (N_12728,N_12347,N_12243);
or U12729 (N_12729,N_12389,N_12194);
or U12730 (N_12730,N_12330,N_12001);
xor U12731 (N_12731,N_12383,N_12292);
nor U12732 (N_12732,N_12457,N_12267);
nand U12733 (N_12733,N_12100,N_12062);
or U12734 (N_12734,N_12145,N_12205);
and U12735 (N_12735,N_12079,N_12130);
xor U12736 (N_12736,N_12397,N_12151);
or U12737 (N_12737,N_12482,N_12432);
and U12738 (N_12738,N_12237,N_12300);
or U12739 (N_12739,N_12343,N_12175);
or U12740 (N_12740,N_12352,N_12149);
xor U12741 (N_12741,N_12446,N_12259);
nand U12742 (N_12742,N_12122,N_12184);
nor U12743 (N_12743,N_12030,N_12229);
or U12744 (N_12744,N_12088,N_12230);
nor U12745 (N_12745,N_12069,N_12283);
nor U12746 (N_12746,N_12224,N_12354);
nor U12747 (N_12747,N_12310,N_12349);
xor U12748 (N_12748,N_12495,N_12169);
xnor U12749 (N_12749,N_12449,N_12208);
or U12750 (N_12750,N_12433,N_12471);
and U12751 (N_12751,N_12439,N_12232);
nor U12752 (N_12752,N_12057,N_12345);
or U12753 (N_12753,N_12422,N_12341);
nand U12754 (N_12754,N_12065,N_12170);
nor U12755 (N_12755,N_12486,N_12063);
nor U12756 (N_12756,N_12110,N_12166);
and U12757 (N_12757,N_12089,N_12060);
or U12758 (N_12758,N_12037,N_12165);
and U12759 (N_12759,N_12058,N_12087);
and U12760 (N_12760,N_12485,N_12144);
or U12761 (N_12761,N_12262,N_12042);
or U12762 (N_12762,N_12039,N_12117);
or U12763 (N_12763,N_12194,N_12315);
or U12764 (N_12764,N_12216,N_12044);
nor U12765 (N_12765,N_12349,N_12223);
nor U12766 (N_12766,N_12434,N_12496);
nand U12767 (N_12767,N_12086,N_12325);
or U12768 (N_12768,N_12403,N_12347);
nand U12769 (N_12769,N_12480,N_12353);
nor U12770 (N_12770,N_12381,N_12416);
xor U12771 (N_12771,N_12280,N_12466);
and U12772 (N_12772,N_12362,N_12173);
nand U12773 (N_12773,N_12413,N_12072);
or U12774 (N_12774,N_12042,N_12175);
nor U12775 (N_12775,N_12380,N_12151);
or U12776 (N_12776,N_12444,N_12427);
nor U12777 (N_12777,N_12287,N_12377);
xnor U12778 (N_12778,N_12358,N_12463);
and U12779 (N_12779,N_12202,N_12112);
or U12780 (N_12780,N_12494,N_12138);
or U12781 (N_12781,N_12276,N_12149);
and U12782 (N_12782,N_12268,N_12185);
and U12783 (N_12783,N_12367,N_12058);
nor U12784 (N_12784,N_12305,N_12189);
or U12785 (N_12785,N_12457,N_12414);
nand U12786 (N_12786,N_12265,N_12432);
and U12787 (N_12787,N_12181,N_12263);
nand U12788 (N_12788,N_12190,N_12453);
nand U12789 (N_12789,N_12234,N_12360);
nand U12790 (N_12790,N_12339,N_12327);
nand U12791 (N_12791,N_12125,N_12037);
xnor U12792 (N_12792,N_12428,N_12254);
or U12793 (N_12793,N_12065,N_12010);
nor U12794 (N_12794,N_12389,N_12095);
nand U12795 (N_12795,N_12243,N_12305);
nor U12796 (N_12796,N_12177,N_12163);
nor U12797 (N_12797,N_12226,N_12445);
nand U12798 (N_12798,N_12382,N_12152);
xor U12799 (N_12799,N_12080,N_12378);
nor U12800 (N_12800,N_12164,N_12064);
nand U12801 (N_12801,N_12434,N_12411);
nor U12802 (N_12802,N_12020,N_12108);
nor U12803 (N_12803,N_12357,N_12134);
nand U12804 (N_12804,N_12059,N_12321);
or U12805 (N_12805,N_12418,N_12079);
nor U12806 (N_12806,N_12138,N_12356);
and U12807 (N_12807,N_12223,N_12215);
xnor U12808 (N_12808,N_12288,N_12306);
and U12809 (N_12809,N_12362,N_12209);
or U12810 (N_12810,N_12340,N_12390);
or U12811 (N_12811,N_12402,N_12088);
and U12812 (N_12812,N_12333,N_12258);
xor U12813 (N_12813,N_12323,N_12186);
nor U12814 (N_12814,N_12296,N_12064);
and U12815 (N_12815,N_12093,N_12199);
xor U12816 (N_12816,N_12468,N_12321);
or U12817 (N_12817,N_12344,N_12218);
xor U12818 (N_12818,N_12039,N_12195);
nand U12819 (N_12819,N_12416,N_12344);
nand U12820 (N_12820,N_12116,N_12186);
and U12821 (N_12821,N_12109,N_12484);
nand U12822 (N_12822,N_12158,N_12377);
nand U12823 (N_12823,N_12215,N_12156);
and U12824 (N_12824,N_12241,N_12351);
nor U12825 (N_12825,N_12138,N_12427);
and U12826 (N_12826,N_12419,N_12421);
xnor U12827 (N_12827,N_12383,N_12138);
nor U12828 (N_12828,N_12008,N_12048);
nand U12829 (N_12829,N_12279,N_12423);
nor U12830 (N_12830,N_12003,N_12304);
xor U12831 (N_12831,N_12478,N_12188);
and U12832 (N_12832,N_12361,N_12087);
or U12833 (N_12833,N_12286,N_12074);
or U12834 (N_12834,N_12248,N_12324);
nand U12835 (N_12835,N_12267,N_12445);
and U12836 (N_12836,N_12331,N_12239);
nand U12837 (N_12837,N_12049,N_12322);
nor U12838 (N_12838,N_12215,N_12240);
nand U12839 (N_12839,N_12194,N_12163);
nand U12840 (N_12840,N_12018,N_12248);
nor U12841 (N_12841,N_12245,N_12179);
and U12842 (N_12842,N_12309,N_12265);
or U12843 (N_12843,N_12430,N_12375);
xnor U12844 (N_12844,N_12009,N_12163);
nand U12845 (N_12845,N_12346,N_12193);
or U12846 (N_12846,N_12399,N_12491);
and U12847 (N_12847,N_12007,N_12431);
and U12848 (N_12848,N_12356,N_12393);
or U12849 (N_12849,N_12295,N_12038);
or U12850 (N_12850,N_12441,N_12489);
or U12851 (N_12851,N_12356,N_12394);
or U12852 (N_12852,N_12098,N_12030);
and U12853 (N_12853,N_12119,N_12194);
and U12854 (N_12854,N_12147,N_12122);
nand U12855 (N_12855,N_12455,N_12387);
or U12856 (N_12856,N_12232,N_12249);
xor U12857 (N_12857,N_12225,N_12084);
and U12858 (N_12858,N_12403,N_12068);
and U12859 (N_12859,N_12378,N_12412);
or U12860 (N_12860,N_12486,N_12015);
nor U12861 (N_12861,N_12404,N_12117);
nor U12862 (N_12862,N_12048,N_12005);
nor U12863 (N_12863,N_12225,N_12420);
nand U12864 (N_12864,N_12280,N_12258);
nand U12865 (N_12865,N_12382,N_12345);
and U12866 (N_12866,N_12389,N_12415);
nor U12867 (N_12867,N_12458,N_12171);
or U12868 (N_12868,N_12013,N_12214);
or U12869 (N_12869,N_12035,N_12405);
nand U12870 (N_12870,N_12267,N_12381);
and U12871 (N_12871,N_12236,N_12395);
or U12872 (N_12872,N_12080,N_12181);
or U12873 (N_12873,N_12497,N_12422);
xnor U12874 (N_12874,N_12098,N_12384);
xor U12875 (N_12875,N_12443,N_12029);
or U12876 (N_12876,N_12315,N_12045);
xnor U12877 (N_12877,N_12083,N_12047);
nand U12878 (N_12878,N_12007,N_12012);
nor U12879 (N_12879,N_12020,N_12345);
nand U12880 (N_12880,N_12400,N_12034);
nand U12881 (N_12881,N_12311,N_12188);
and U12882 (N_12882,N_12359,N_12346);
nor U12883 (N_12883,N_12396,N_12007);
and U12884 (N_12884,N_12455,N_12010);
or U12885 (N_12885,N_12478,N_12107);
nor U12886 (N_12886,N_12086,N_12072);
xor U12887 (N_12887,N_12305,N_12132);
nand U12888 (N_12888,N_12250,N_12052);
nand U12889 (N_12889,N_12462,N_12475);
or U12890 (N_12890,N_12318,N_12178);
or U12891 (N_12891,N_12239,N_12395);
or U12892 (N_12892,N_12074,N_12285);
nor U12893 (N_12893,N_12370,N_12007);
nand U12894 (N_12894,N_12095,N_12112);
nand U12895 (N_12895,N_12123,N_12396);
or U12896 (N_12896,N_12471,N_12309);
nor U12897 (N_12897,N_12098,N_12160);
nor U12898 (N_12898,N_12117,N_12360);
xnor U12899 (N_12899,N_12003,N_12020);
nand U12900 (N_12900,N_12441,N_12425);
xnor U12901 (N_12901,N_12096,N_12480);
or U12902 (N_12902,N_12363,N_12033);
nand U12903 (N_12903,N_12223,N_12195);
or U12904 (N_12904,N_12159,N_12029);
xnor U12905 (N_12905,N_12384,N_12283);
and U12906 (N_12906,N_12429,N_12329);
nand U12907 (N_12907,N_12300,N_12390);
nor U12908 (N_12908,N_12396,N_12279);
nor U12909 (N_12909,N_12340,N_12265);
or U12910 (N_12910,N_12253,N_12156);
xor U12911 (N_12911,N_12214,N_12379);
and U12912 (N_12912,N_12455,N_12373);
nor U12913 (N_12913,N_12419,N_12342);
and U12914 (N_12914,N_12241,N_12158);
and U12915 (N_12915,N_12498,N_12363);
and U12916 (N_12916,N_12327,N_12416);
or U12917 (N_12917,N_12385,N_12257);
or U12918 (N_12918,N_12311,N_12081);
and U12919 (N_12919,N_12180,N_12177);
xnor U12920 (N_12920,N_12294,N_12465);
nor U12921 (N_12921,N_12103,N_12240);
and U12922 (N_12922,N_12347,N_12049);
and U12923 (N_12923,N_12212,N_12041);
nor U12924 (N_12924,N_12195,N_12412);
or U12925 (N_12925,N_12363,N_12087);
nor U12926 (N_12926,N_12065,N_12002);
or U12927 (N_12927,N_12378,N_12011);
or U12928 (N_12928,N_12133,N_12037);
or U12929 (N_12929,N_12219,N_12139);
nor U12930 (N_12930,N_12463,N_12287);
or U12931 (N_12931,N_12330,N_12374);
or U12932 (N_12932,N_12091,N_12422);
and U12933 (N_12933,N_12398,N_12062);
nor U12934 (N_12934,N_12198,N_12276);
nand U12935 (N_12935,N_12449,N_12498);
nor U12936 (N_12936,N_12294,N_12420);
nor U12937 (N_12937,N_12452,N_12322);
or U12938 (N_12938,N_12082,N_12429);
nand U12939 (N_12939,N_12052,N_12332);
nand U12940 (N_12940,N_12146,N_12244);
or U12941 (N_12941,N_12319,N_12170);
nand U12942 (N_12942,N_12073,N_12379);
and U12943 (N_12943,N_12485,N_12338);
nand U12944 (N_12944,N_12005,N_12423);
nor U12945 (N_12945,N_12437,N_12100);
nand U12946 (N_12946,N_12044,N_12496);
nand U12947 (N_12947,N_12487,N_12167);
nor U12948 (N_12948,N_12239,N_12481);
or U12949 (N_12949,N_12432,N_12164);
or U12950 (N_12950,N_12466,N_12158);
nor U12951 (N_12951,N_12136,N_12038);
or U12952 (N_12952,N_12331,N_12186);
and U12953 (N_12953,N_12154,N_12431);
or U12954 (N_12954,N_12497,N_12165);
and U12955 (N_12955,N_12078,N_12164);
nor U12956 (N_12956,N_12143,N_12296);
nand U12957 (N_12957,N_12254,N_12226);
xnor U12958 (N_12958,N_12263,N_12371);
or U12959 (N_12959,N_12136,N_12434);
or U12960 (N_12960,N_12431,N_12218);
or U12961 (N_12961,N_12458,N_12443);
nor U12962 (N_12962,N_12125,N_12087);
xor U12963 (N_12963,N_12053,N_12391);
nand U12964 (N_12964,N_12027,N_12310);
and U12965 (N_12965,N_12239,N_12216);
nor U12966 (N_12966,N_12483,N_12022);
or U12967 (N_12967,N_12269,N_12255);
or U12968 (N_12968,N_12475,N_12445);
nand U12969 (N_12969,N_12045,N_12389);
and U12970 (N_12970,N_12036,N_12471);
xor U12971 (N_12971,N_12307,N_12409);
nand U12972 (N_12972,N_12340,N_12038);
or U12973 (N_12973,N_12355,N_12339);
nand U12974 (N_12974,N_12382,N_12011);
nor U12975 (N_12975,N_12271,N_12232);
nor U12976 (N_12976,N_12010,N_12188);
or U12977 (N_12977,N_12072,N_12030);
and U12978 (N_12978,N_12186,N_12061);
nand U12979 (N_12979,N_12201,N_12079);
nand U12980 (N_12980,N_12197,N_12428);
or U12981 (N_12981,N_12200,N_12322);
xnor U12982 (N_12982,N_12330,N_12334);
nand U12983 (N_12983,N_12272,N_12481);
or U12984 (N_12984,N_12402,N_12489);
nand U12985 (N_12985,N_12207,N_12141);
or U12986 (N_12986,N_12019,N_12451);
and U12987 (N_12987,N_12043,N_12176);
nor U12988 (N_12988,N_12431,N_12015);
or U12989 (N_12989,N_12384,N_12193);
and U12990 (N_12990,N_12039,N_12203);
or U12991 (N_12991,N_12021,N_12099);
xnor U12992 (N_12992,N_12288,N_12204);
and U12993 (N_12993,N_12123,N_12372);
or U12994 (N_12994,N_12436,N_12206);
and U12995 (N_12995,N_12365,N_12088);
nor U12996 (N_12996,N_12162,N_12192);
and U12997 (N_12997,N_12031,N_12475);
nor U12998 (N_12998,N_12188,N_12051);
nand U12999 (N_12999,N_12037,N_12358);
nor U13000 (N_13000,N_12897,N_12939);
or U13001 (N_13001,N_12928,N_12709);
xnor U13002 (N_13002,N_12557,N_12949);
xnor U13003 (N_13003,N_12951,N_12637);
nand U13004 (N_13004,N_12663,N_12901);
nor U13005 (N_13005,N_12683,N_12684);
and U13006 (N_13006,N_12696,N_12531);
and U13007 (N_13007,N_12769,N_12915);
nor U13008 (N_13008,N_12892,N_12614);
or U13009 (N_13009,N_12802,N_12612);
and U13010 (N_13010,N_12755,N_12941);
nor U13011 (N_13011,N_12877,N_12604);
nor U13012 (N_13012,N_12902,N_12569);
nor U13013 (N_13013,N_12727,N_12729);
or U13014 (N_13014,N_12969,N_12863);
and U13015 (N_13015,N_12946,N_12761);
nor U13016 (N_13016,N_12634,N_12916);
or U13017 (N_13017,N_12717,N_12801);
and U13018 (N_13018,N_12597,N_12811);
and U13019 (N_13019,N_12558,N_12805);
nand U13020 (N_13020,N_12733,N_12918);
nand U13021 (N_13021,N_12615,N_12990);
nand U13022 (N_13022,N_12988,N_12987);
or U13023 (N_13023,N_12803,N_12715);
or U13024 (N_13024,N_12914,N_12925);
nor U13025 (N_13025,N_12705,N_12551);
nand U13026 (N_13026,N_12991,N_12591);
or U13027 (N_13027,N_12593,N_12520);
nand U13028 (N_13028,N_12688,N_12514);
xor U13029 (N_13029,N_12734,N_12828);
nand U13030 (N_13030,N_12837,N_12711);
and U13031 (N_13031,N_12898,N_12701);
and U13032 (N_13032,N_12538,N_12995);
and U13033 (N_13033,N_12876,N_12865);
and U13034 (N_13034,N_12576,N_12840);
nor U13035 (N_13035,N_12697,N_12573);
or U13036 (N_13036,N_12545,N_12555);
nand U13037 (N_13037,N_12799,N_12706);
or U13038 (N_13038,N_12601,N_12605);
or U13039 (N_13039,N_12617,N_12740);
or U13040 (N_13040,N_12971,N_12672);
and U13041 (N_13041,N_12857,N_12927);
and U13042 (N_13042,N_12885,N_12940);
nand U13043 (N_13043,N_12728,N_12750);
xnor U13044 (N_13044,N_12800,N_12689);
nor U13045 (N_13045,N_12638,N_12947);
nand U13046 (N_13046,N_12570,N_12631);
and U13047 (N_13047,N_12838,N_12602);
nor U13048 (N_13048,N_12698,N_12603);
nor U13049 (N_13049,N_12792,N_12513);
and U13050 (N_13050,N_12749,N_12608);
and U13051 (N_13051,N_12607,N_12547);
or U13052 (N_13052,N_12550,N_12599);
nor U13053 (N_13053,N_12894,N_12797);
nand U13054 (N_13054,N_12989,N_12847);
and U13055 (N_13055,N_12537,N_12870);
or U13056 (N_13056,N_12955,N_12624);
and U13057 (N_13057,N_12906,N_12515);
and U13058 (N_13058,N_12850,N_12732);
and U13059 (N_13059,N_12678,N_12950);
nand U13060 (N_13060,N_12977,N_12896);
or U13061 (N_13061,N_12700,N_12763);
and U13062 (N_13062,N_12751,N_12540);
xor U13063 (N_13063,N_12888,N_12726);
nand U13064 (N_13064,N_12543,N_12868);
and U13065 (N_13065,N_12641,N_12767);
nand U13066 (N_13066,N_12835,N_12563);
or U13067 (N_13067,N_12737,N_12996);
xnor U13068 (N_13068,N_12660,N_12534);
nand U13069 (N_13069,N_12845,N_12900);
nand U13070 (N_13070,N_12787,N_12796);
xor U13071 (N_13071,N_12587,N_12775);
xor U13072 (N_13072,N_12772,N_12654);
nor U13073 (N_13073,N_12606,N_12924);
and U13074 (N_13074,N_12699,N_12765);
nor U13075 (N_13075,N_12762,N_12783);
nand U13076 (N_13076,N_12836,N_12610);
and U13077 (N_13077,N_12577,N_12650);
or U13078 (N_13078,N_12964,N_12721);
nor U13079 (N_13079,N_12632,N_12937);
nand U13080 (N_13080,N_12725,N_12708);
or U13081 (N_13081,N_12583,N_12812);
nor U13082 (N_13082,N_12507,N_12829);
nand U13083 (N_13083,N_12776,N_12826);
or U13084 (N_13084,N_12562,N_12856);
nor U13085 (N_13085,N_12667,N_12968);
nand U13086 (N_13086,N_12822,N_12908);
or U13087 (N_13087,N_12975,N_12517);
nor U13088 (N_13088,N_12903,N_12861);
nor U13089 (N_13089,N_12806,N_12756);
and U13090 (N_13090,N_12527,N_12649);
nand U13091 (N_13091,N_12919,N_12773);
nor U13092 (N_13092,N_12702,N_12983);
or U13093 (N_13093,N_12546,N_12665);
and U13094 (N_13094,N_12824,N_12512);
or U13095 (N_13095,N_12798,N_12960);
and U13096 (N_13096,N_12539,N_12578);
nand U13097 (N_13097,N_12895,N_12923);
and U13098 (N_13098,N_12738,N_12674);
or U13099 (N_13099,N_12635,N_12985);
nand U13100 (N_13100,N_12963,N_12646);
and U13101 (N_13101,N_12505,N_12661);
nor U13102 (N_13102,N_12890,N_12613);
nand U13103 (N_13103,N_12619,N_12707);
or U13104 (N_13104,N_12687,N_12973);
xnor U13105 (N_13105,N_12639,N_12851);
xnor U13106 (N_13106,N_12957,N_12848);
and U13107 (N_13107,N_12883,N_12935);
and U13108 (N_13108,N_12759,N_12774);
nand U13109 (N_13109,N_12657,N_12781);
nor U13110 (N_13110,N_12714,N_12766);
nand U13111 (N_13111,N_12817,N_12530);
or U13112 (N_13112,N_12532,N_12735);
and U13113 (N_13113,N_12720,N_12501);
and U13114 (N_13114,N_12712,N_12998);
and U13115 (N_13115,N_12832,N_12926);
xnor U13116 (N_13116,N_12544,N_12757);
nor U13117 (N_13117,N_12743,N_12954);
or U13118 (N_13118,N_12982,N_12967);
nand U13119 (N_13119,N_12907,N_12930);
or U13120 (N_13120,N_12965,N_12535);
or U13121 (N_13121,N_12582,N_12742);
and U13122 (N_13122,N_12536,N_12867);
xnor U13123 (N_13123,N_12986,N_12585);
or U13124 (N_13124,N_12658,N_12655);
nor U13125 (N_13125,N_12815,N_12818);
or U13126 (N_13126,N_12589,N_12600);
nand U13127 (N_13127,N_12913,N_12911);
and U13128 (N_13128,N_12528,N_12859);
xnor U13129 (N_13129,N_12889,N_12872);
xor U13130 (N_13130,N_12575,N_12922);
or U13131 (N_13131,N_12782,N_12640);
nor U13132 (N_13132,N_12652,N_12723);
nor U13133 (N_13133,N_12703,N_12653);
and U13134 (N_13134,N_12970,N_12584);
nor U13135 (N_13135,N_12921,N_12594);
and U13136 (N_13136,N_12521,N_12616);
or U13137 (N_13137,N_12609,N_12580);
nor U13138 (N_13138,N_12526,N_12718);
nor U13139 (N_13139,N_12887,N_12984);
nor U13140 (N_13140,N_12679,N_12938);
and U13141 (N_13141,N_12980,N_12878);
nand U13142 (N_13142,N_12739,N_12814);
nand U13143 (N_13143,N_12785,N_12559);
and U13144 (N_13144,N_12866,N_12636);
or U13145 (N_13145,N_12753,N_12754);
and U13146 (N_13146,N_12588,N_12586);
nor U13147 (N_13147,N_12554,N_12548);
nor U13148 (N_13148,N_12523,N_12692);
nor U13149 (N_13149,N_12959,N_12858);
nor U13150 (N_13150,N_12500,N_12666);
nand U13151 (N_13151,N_12685,N_12849);
xnor U13152 (N_13152,N_12932,N_12552);
and U13153 (N_13153,N_12830,N_12675);
nand U13154 (N_13154,N_12899,N_12936);
nor U13155 (N_13155,N_12966,N_12670);
nor U13156 (N_13156,N_12839,N_12627);
nor U13157 (N_13157,N_12779,N_12522);
or U13158 (N_13158,N_12553,N_12791);
and U13159 (N_13159,N_12869,N_12648);
or U13160 (N_13160,N_12962,N_12778);
nand U13161 (N_13161,N_12997,N_12746);
nor U13162 (N_13162,N_12948,N_12819);
nand U13163 (N_13163,N_12760,N_12904);
xnor U13164 (N_13164,N_12671,N_12506);
or U13165 (N_13165,N_12565,N_12710);
nand U13166 (N_13166,N_12825,N_12647);
and U13167 (N_13167,N_12525,N_12691);
or U13168 (N_13168,N_12579,N_12611);
and U13169 (N_13169,N_12680,N_12677);
nor U13170 (N_13170,N_12854,N_12541);
nor U13171 (N_13171,N_12623,N_12722);
nor U13172 (N_13172,N_12823,N_12626);
nand U13173 (N_13173,N_12944,N_12643);
nor U13174 (N_13174,N_12629,N_12524);
nand U13175 (N_13175,N_12795,N_12716);
or U13176 (N_13176,N_12855,N_12833);
nand U13177 (N_13177,N_12956,N_12846);
nand U13178 (N_13178,N_12644,N_12628);
nor U13179 (N_13179,N_12567,N_12841);
and U13180 (N_13180,N_12503,N_12731);
or U13181 (N_13181,N_12504,N_12695);
nor U13182 (N_13182,N_12862,N_12719);
and U13183 (N_13183,N_12871,N_12912);
or U13184 (N_13184,N_12768,N_12789);
xor U13185 (N_13185,N_12886,N_12917);
xnor U13186 (N_13186,N_12693,N_12518);
nand U13187 (N_13187,N_12744,N_12972);
nor U13188 (N_13188,N_12909,N_12842);
and U13189 (N_13189,N_12809,N_12574);
nand U13190 (N_13190,N_12905,N_12820);
and U13191 (N_13191,N_12929,N_12880);
xnor U13192 (N_13192,N_12549,N_12974);
or U13193 (N_13193,N_12976,N_12808);
nand U13194 (N_13194,N_12943,N_12621);
and U13195 (N_13195,N_12533,N_12999);
nand U13196 (N_13196,N_12981,N_12682);
and U13197 (N_13197,N_12595,N_12879);
or U13198 (N_13198,N_12780,N_12572);
nor U13199 (N_13199,N_12592,N_12669);
nor U13200 (N_13200,N_12843,N_12642);
nand U13201 (N_13201,N_12993,N_12771);
and U13202 (N_13202,N_12724,N_12741);
and U13203 (N_13203,N_12873,N_12560);
and U13204 (N_13204,N_12790,N_12747);
nand U13205 (N_13205,N_12992,N_12786);
and U13206 (N_13206,N_12978,N_12794);
nor U13207 (N_13207,N_12810,N_12953);
and U13208 (N_13208,N_12590,N_12994);
nand U13209 (N_13209,N_12508,N_12681);
and U13210 (N_13210,N_12622,N_12875);
nand U13211 (N_13211,N_12788,N_12686);
and U13212 (N_13212,N_12630,N_12933);
or U13213 (N_13213,N_12910,N_12784);
xor U13214 (N_13214,N_12694,N_12618);
or U13215 (N_13215,N_12568,N_12516);
nand U13216 (N_13216,N_12529,N_12690);
xor U13217 (N_13217,N_12620,N_12511);
xnor U13218 (N_13218,N_12730,N_12668);
or U13219 (N_13219,N_12645,N_12931);
nor U13220 (N_13220,N_12664,N_12745);
nor U13221 (N_13221,N_12566,N_12852);
and U13222 (N_13222,N_12882,N_12571);
and U13223 (N_13223,N_12564,N_12752);
nor U13224 (N_13224,N_12758,N_12625);
xnor U13225 (N_13225,N_12519,N_12598);
and U13226 (N_13226,N_12502,N_12736);
or U13227 (N_13227,N_12673,N_12834);
and U13228 (N_13228,N_12633,N_12945);
and U13229 (N_13229,N_12816,N_12656);
or U13230 (N_13230,N_12893,N_12853);
and U13231 (N_13231,N_12676,N_12844);
and U13232 (N_13232,N_12807,N_12827);
or U13233 (N_13233,N_12864,N_12748);
and U13234 (N_13234,N_12942,N_12561);
nand U13235 (N_13235,N_12958,N_12891);
nor U13236 (N_13236,N_12770,N_12764);
and U13237 (N_13237,N_12831,N_12777);
nor U13238 (N_13238,N_12884,N_12804);
or U13239 (N_13239,N_12662,N_12881);
nand U13240 (N_13240,N_12704,N_12952);
or U13241 (N_13241,N_12509,N_12813);
nand U13242 (N_13242,N_12556,N_12596);
xor U13243 (N_13243,N_12821,N_12793);
and U13244 (N_13244,N_12651,N_12934);
nor U13245 (N_13245,N_12874,N_12542);
and U13246 (N_13246,N_12713,N_12979);
and U13247 (N_13247,N_12860,N_12961);
nand U13248 (N_13248,N_12510,N_12659);
nand U13249 (N_13249,N_12920,N_12581);
or U13250 (N_13250,N_12590,N_12961);
or U13251 (N_13251,N_12555,N_12670);
and U13252 (N_13252,N_12940,N_12732);
nand U13253 (N_13253,N_12561,N_12977);
or U13254 (N_13254,N_12654,N_12596);
nand U13255 (N_13255,N_12938,N_12806);
or U13256 (N_13256,N_12995,N_12788);
or U13257 (N_13257,N_12985,N_12620);
nor U13258 (N_13258,N_12718,N_12790);
nor U13259 (N_13259,N_12522,N_12632);
and U13260 (N_13260,N_12771,N_12893);
or U13261 (N_13261,N_12562,N_12756);
or U13262 (N_13262,N_12872,N_12926);
and U13263 (N_13263,N_12852,N_12743);
or U13264 (N_13264,N_12650,N_12634);
nor U13265 (N_13265,N_12826,N_12660);
xor U13266 (N_13266,N_12625,N_12689);
nor U13267 (N_13267,N_12646,N_12657);
and U13268 (N_13268,N_12769,N_12638);
nor U13269 (N_13269,N_12640,N_12787);
nand U13270 (N_13270,N_12615,N_12660);
and U13271 (N_13271,N_12848,N_12526);
nor U13272 (N_13272,N_12730,N_12688);
nor U13273 (N_13273,N_12779,N_12896);
or U13274 (N_13274,N_12630,N_12723);
nand U13275 (N_13275,N_12687,N_12778);
nand U13276 (N_13276,N_12667,N_12625);
and U13277 (N_13277,N_12967,N_12955);
nor U13278 (N_13278,N_12798,N_12826);
nor U13279 (N_13279,N_12669,N_12586);
nand U13280 (N_13280,N_12642,N_12993);
nand U13281 (N_13281,N_12731,N_12519);
nand U13282 (N_13282,N_12639,N_12879);
nor U13283 (N_13283,N_12744,N_12845);
nor U13284 (N_13284,N_12892,N_12836);
xor U13285 (N_13285,N_12876,N_12780);
and U13286 (N_13286,N_12950,N_12603);
or U13287 (N_13287,N_12915,N_12759);
nor U13288 (N_13288,N_12894,N_12750);
nand U13289 (N_13289,N_12808,N_12970);
and U13290 (N_13290,N_12555,N_12721);
nor U13291 (N_13291,N_12724,N_12836);
xnor U13292 (N_13292,N_12802,N_12540);
and U13293 (N_13293,N_12678,N_12731);
nand U13294 (N_13294,N_12646,N_12944);
xnor U13295 (N_13295,N_12913,N_12738);
or U13296 (N_13296,N_12901,N_12674);
nand U13297 (N_13297,N_12666,N_12709);
xor U13298 (N_13298,N_12631,N_12673);
or U13299 (N_13299,N_12848,N_12524);
nand U13300 (N_13300,N_12529,N_12997);
or U13301 (N_13301,N_12840,N_12754);
and U13302 (N_13302,N_12743,N_12597);
nor U13303 (N_13303,N_12861,N_12957);
or U13304 (N_13304,N_12682,N_12511);
nand U13305 (N_13305,N_12839,N_12812);
nor U13306 (N_13306,N_12550,N_12667);
nand U13307 (N_13307,N_12730,N_12875);
nand U13308 (N_13308,N_12805,N_12864);
nor U13309 (N_13309,N_12838,N_12813);
or U13310 (N_13310,N_12536,N_12750);
nor U13311 (N_13311,N_12930,N_12836);
nor U13312 (N_13312,N_12775,N_12502);
and U13313 (N_13313,N_12528,N_12915);
and U13314 (N_13314,N_12558,N_12755);
nand U13315 (N_13315,N_12519,N_12624);
nand U13316 (N_13316,N_12746,N_12541);
or U13317 (N_13317,N_12832,N_12729);
or U13318 (N_13318,N_12934,N_12535);
xnor U13319 (N_13319,N_12849,N_12654);
nand U13320 (N_13320,N_12733,N_12694);
and U13321 (N_13321,N_12577,N_12552);
nor U13322 (N_13322,N_12773,N_12815);
and U13323 (N_13323,N_12718,N_12633);
and U13324 (N_13324,N_12820,N_12540);
nand U13325 (N_13325,N_12803,N_12885);
and U13326 (N_13326,N_12815,N_12843);
nand U13327 (N_13327,N_12746,N_12821);
or U13328 (N_13328,N_12677,N_12654);
and U13329 (N_13329,N_12876,N_12842);
nand U13330 (N_13330,N_12974,N_12933);
nor U13331 (N_13331,N_12775,N_12578);
or U13332 (N_13332,N_12896,N_12712);
and U13333 (N_13333,N_12509,N_12991);
or U13334 (N_13334,N_12560,N_12578);
nor U13335 (N_13335,N_12843,N_12787);
and U13336 (N_13336,N_12740,N_12558);
and U13337 (N_13337,N_12515,N_12501);
nand U13338 (N_13338,N_12983,N_12724);
nand U13339 (N_13339,N_12886,N_12595);
nor U13340 (N_13340,N_12504,N_12561);
nand U13341 (N_13341,N_12925,N_12640);
xor U13342 (N_13342,N_12737,N_12960);
nand U13343 (N_13343,N_12529,N_12806);
and U13344 (N_13344,N_12628,N_12782);
nand U13345 (N_13345,N_12895,N_12716);
or U13346 (N_13346,N_12699,N_12930);
nor U13347 (N_13347,N_12721,N_12800);
or U13348 (N_13348,N_12906,N_12743);
or U13349 (N_13349,N_12673,N_12867);
and U13350 (N_13350,N_12536,N_12537);
nand U13351 (N_13351,N_12831,N_12958);
or U13352 (N_13352,N_12814,N_12525);
and U13353 (N_13353,N_12621,N_12527);
or U13354 (N_13354,N_12754,N_12525);
or U13355 (N_13355,N_12665,N_12932);
xnor U13356 (N_13356,N_12734,N_12971);
or U13357 (N_13357,N_12971,N_12582);
and U13358 (N_13358,N_12943,N_12922);
or U13359 (N_13359,N_12729,N_12692);
and U13360 (N_13360,N_12580,N_12983);
and U13361 (N_13361,N_12800,N_12993);
nand U13362 (N_13362,N_12770,N_12792);
nand U13363 (N_13363,N_12853,N_12673);
and U13364 (N_13364,N_12735,N_12930);
nand U13365 (N_13365,N_12525,N_12577);
or U13366 (N_13366,N_12703,N_12726);
or U13367 (N_13367,N_12717,N_12766);
nor U13368 (N_13368,N_12620,N_12568);
nor U13369 (N_13369,N_12920,N_12547);
or U13370 (N_13370,N_12692,N_12571);
xnor U13371 (N_13371,N_12967,N_12836);
nand U13372 (N_13372,N_12802,N_12656);
nand U13373 (N_13373,N_12861,N_12920);
nor U13374 (N_13374,N_12816,N_12802);
nor U13375 (N_13375,N_12546,N_12970);
nand U13376 (N_13376,N_12754,N_12994);
nor U13377 (N_13377,N_12554,N_12558);
and U13378 (N_13378,N_12855,N_12580);
or U13379 (N_13379,N_12906,N_12696);
xor U13380 (N_13380,N_12507,N_12791);
nand U13381 (N_13381,N_12550,N_12519);
nor U13382 (N_13382,N_12944,N_12703);
nor U13383 (N_13383,N_12866,N_12845);
or U13384 (N_13384,N_12894,N_12595);
nor U13385 (N_13385,N_12774,N_12621);
or U13386 (N_13386,N_12742,N_12775);
and U13387 (N_13387,N_12617,N_12925);
nor U13388 (N_13388,N_12615,N_12776);
and U13389 (N_13389,N_12947,N_12672);
nor U13390 (N_13390,N_12784,N_12625);
nor U13391 (N_13391,N_12720,N_12841);
and U13392 (N_13392,N_12852,N_12646);
nand U13393 (N_13393,N_12780,N_12518);
and U13394 (N_13394,N_12885,N_12897);
nand U13395 (N_13395,N_12730,N_12624);
and U13396 (N_13396,N_12766,N_12795);
nand U13397 (N_13397,N_12971,N_12756);
or U13398 (N_13398,N_12796,N_12954);
or U13399 (N_13399,N_12613,N_12651);
and U13400 (N_13400,N_12704,N_12931);
or U13401 (N_13401,N_12782,N_12626);
and U13402 (N_13402,N_12680,N_12823);
nor U13403 (N_13403,N_12905,N_12749);
nand U13404 (N_13404,N_12501,N_12929);
nor U13405 (N_13405,N_12945,N_12707);
or U13406 (N_13406,N_12547,N_12564);
or U13407 (N_13407,N_12907,N_12581);
nand U13408 (N_13408,N_12684,N_12537);
or U13409 (N_13409,N_12759,N_12899);
nor U13410 (N_13410,N_12806,N_12538);
or U13411 (N_13411,N_12746,N_12979);
nand U13412 (N_13412,N_12577,N_12932);
and U13413 (N_13413,N_12913,N_12879);
xor U13414 (N_13414,N_12772,N_12955);
nor U13415 (N_13415,N_12913,N_12665);
or U13416 (N_13416,N_12846,N_12694);
and U13417 (N_13417,N_12595,N_12762);
or U13418 (N_13418,N_12679,N_12674);
or U13419 (N_13419,N_12616,N_12774);
or U13420 (N_13420,N_12906,N_12501);
and U13421 (N_13421,N_12523,N_12796);
nand U13422 (N_13422,N_12918,N_12549);
nand U13423 (N_13423,N_12879,N_12855);
or U13424 (N_13424,N_12934,N_12908);
and U13425 (N_13425,N_12877,N_12514);
nor U13426 (N_13426,N_12520,N_12815);
or U13427 (N_13427,N_12601,N_12889);
or U13428 (N_13428,N_12685,N_12833);
or U13429 (N_13429,N_12814,N_12585);
and U13430 (N_13430,N_12693,N_12806);
or U13431 (N_13431,N_12512,N_12542);
xnor U13432 (N_13432,N_12732,N_12561);
nand U13433 (N_13433,N_12574,N_12908);
or U13434 (N_13434,N_12868,N_12928);
or U13435 (N_13435,N_12944,N_12661);
and U13436 (N_13436,N_12557,N_12584);
xnor U13437 (N_13437,N_12597,N_12823);
nor U13438 (N_13438,N_12611,N_12676);
and U13439 (N_13439,N_12813,N_12980);
nand U13440 (N_13440,N_12886,N_12516);
nand U13441 (N_13441,N_12931,N_12519);
or U13442 (N_13442,N_12768,N_12986);
or U13443 (N_13443,N_12984,N_12937);
or U13444 (N_13444,N_12993,N_12790);
nand U13445 (N_13445,N_12692,N_12695);
nand U13446 (N_13446,N_12717,N_12938);
xor U13447 (N_13447,N_12544,N_12752);
xnor U13448 (N_13448,N_12953,N_12600);
xor U13449 (N_13449,N_12587,N_12599);
xor U13450 (N_13450,N_12903,N_12746);
xor U13451 (N_13451,N_12915,N_12525);
nand U13452 (N_13452,N_12537,N_12689);
nor U13453 (N_13453,N_12884,N_12805);
nand U13454 (N_13454,N_12961,N_12830);
and U13455 (N_13455,N_12547,N_12927);
and U13456 (N_13456,N_12766,N_12970);
and U13457 (N_13457,N_12624,N_12892);
nor U13458 (N_13458,N_12504,N_12746);
and U13459 (N_13459,N_12767,N_12523);
nand U13460 (N_13460,N_12954,N_12546);
and U13461 (N_13461,N_12567,N_12652);
or U13462 (N_13462,N_12768,N_12950);
nand U13463 (N_13463,N_12637,N_12936);
and U13464 (N_13464,N_12898,N_12792);
or U13465 (N_13465,N_12897,N_12701);
and U13466 (N_13466,N_12735,N_12526);
and U13467 (N_13467,N_12652,N_12632);
or U13468 (N_13468,N_12776,N_12635);
nand U13469 (N_13469,N_12607,N_12703);
nand U13470 (N_13470,N_12839,N_12906);
nor U13471 (N_13471,N_12989,N_12909);
nand U13472 (N_13472,N_12964,N_12565);
and U13473 (N_13473,N_12885,N_12858);
or U13474 (N_13474,N_12648,N_12797);
nand U13475 (N_13475,N_12643,N_12807);
or U13476 (N_13476,N_12948,N_12991);
nand U13477 (N_13477,N_12950,N_12529);
nor U13478 (N_13478,N_12804,N_12614);
nand U13479 (N_13479,N_12857,N_12874);
nor U13480 (N_13480,N_12848,N_12873);
and U13481 (N_13481,N_12510,N_12899);
nor U13482 (N_13482,N_12736,N_12517);
and U13483 (N_13483,N_12834,N_12549);
and U13484 (N_13484,N_12624,N_12654);
and U13485 (N_13485,N_12970,N_12624);
or U13486 (N_13486,N_12596,N_12512);
and U13487 (N_13487,N_12575,N_12501);
nand U13488 (N_13488,N_12755,N_12902);
and U13489 (N_13489,N_12749,N_12967);
and U13490 (N_13490,N_12612,N_12776);
and U13491 (N_13491,N_12645,N_12607);
nor U13492 (N_13492,N_12580,N_12961);
and U13493 (N_13493,N_12900,N_12600);
nor U13494 (N_13494,N_12538,N_12501);
or U13495 (N_13495,N_12521,N_12817);
nor U13496 (N_13496,N_12581,N_12812);
nor U13497 (N_13497,N_12873,N_12524);
nand U13498 (N_13498,N_12568,N_12549);
nor U13499 (N_13499,N_12936,N_12956);
or U13500 (N_13500,N_13285,N_13374);
and U13501 (N_13501,N_13305,N_13162);
nor U13502 (N_13502,N_13045,N_13340);
and U13503 (N_13503,N_13175,N_13358);
or U13504 (N_13504,N_13221,N_13107);
and U13505 (N_13505,N_13409,N_13327);
nor U13506 (N_13506,N_13313,N_13234);
xnor U13507 (N_13507,N_13365,N_13339);
nand U13508 (N_13508,N_13056,N_13241);
nand U13509 (N_13509,N_13036,N_13255);
or U13510 (N_13510,N_13307,N_13141);
or U13511 (N_13511,N_13033,N_13177);
or U13512 (N_13512,N_13052,N_13247);
nand U13513 (N_13513,N_13455,N_13324);
or U13514 (N_13514,N_13115,N_13316);
nor U13515 (N_13515,N_13135,N_13235);
xnor U13516 (N_13516,N_13207,N_13494);
nor U13517 (N_13517,N_13321,N_13000);
or U13518 (N_13518,N_13481,N_13212);
and U13519 (N_13519,N_13419,N_13144);
or U13520 (N_13520,N_13040,N_13006);
and U13521 (N_13521,N_13399,N_13261);
and U13522 (N_13522,N_13490,N_13079);
or U13523 (N_13523,N_13291,N_13075);
and U13524 (N_13524,N_13354,N_13244);
nand U13525 (N_13525,N_13343,N_13041);
nand U13526 (N_13526,N_13251,N_13472);
nor U13527 (N_13527,N_13427,N_13193);
or U13528 (N_13528,N_13421,N_13088);
nor U13529 (N_13529,N_13403,N_13072);
or U13530 (N_13530,N_13432,N_13347);
nand U13531 (N_13531,N_13065,N_13229);
and U13532 (N_13532,N_13023,N_13043);
nor U13533 (N_13533,N_13466,N_13420);
nor U13534 (N_13534,N_13167,N_13149);
xnor U13535 (N_13535,N_13417,N_13430);
or U13536 (N_13536,N_13287,N_13278);
nand U13537 (N_13537,N_13483,N_13332);
and U13538 (N_13538,N_13414,N_13185);
nor U13539 (N_13539,N_13190,N_13310);
and U13540 (N_13540,N_13388,N_13139);
or U13541 (N_13541,N_13165,N_13487);
xor U13542 (N_13542,N_13413,N_13317);
nand U13543 (N_13543,N_13422,N_13001);
or U13544 (N_13544,N_13326,N_13393);
or U13545 (N_13545,N_13173,N_13094);
nor U13546 (N_13546,N_13395,N_13451);
nand U13547 (N_13547,N_13150,N_13133);
xor U13548 (N_13548,N_13439,N_13122);
and U13549 (N_13549,N_13377,N_13262);
or U13550 (N_13550,N_13136,N_13106);
nand U13551 (N_13551,N_13015,N_13131);
nand U13552 (N_13552,N_13405,N_13265);
and U13553 (N_13553,N_13129,N_13312);
nor U13554 (N_13554,N_13484,N_13461);
or U13555 (N_13555,N_13201,N_13010);
and U13556 (N_13556,N_13458,N_13438);
and U13557 (N_13557,N_13449,N_13205);
nand U13558 (N_13558,N_13329,N_13418);
and U13559 (N_13559,N_13037,N_13157);
and U13560 (N_13560,N_13444,N_13152);
nor U13561 (N_13561,N_13352,N_13441);
xnor U13562 (N_13562,N_13496,N_13266);
nand U13563 (N_13563,N_13019,N_13435);
and U13564 (N_13564,N_13391,N_13465);
nand U13565 (N_13565,N_13448,N_13301);
or U13566 (N_13566,N_13055,N_13140);
or U13567 (N_13567,N_13087,N_13469);
or U13568 (N_13568,N_13192,N_13061);
nor U13569 (N_13569,N_13240,N_13126);
nand U13570 (N_13570,N_13179,N_13191);
and U13571 (N_13571,N_13369,N_13258);
and U13572 (N_13572,N_13263,N_13097);
nand U13573 (N_13573,N_13187,N_13400);
nor U13574 (N_13574,N_13368,N_13463);
nand U13575 (N_13575,N_13223,N_13489);
nand U13576 (N_13576,N_13314,N_13119);
nand U13577 (N_13577,N_13213,N_13308);
nand U13578 (N_13578,N_13289,N_13480);
xnor U13579 (N_13579,N_13154,N_13160);
nor U13580 (N_13580,N_13090,N_13073);
nor U13581 (N_13581,N_13013,N_13074);
and U13582 (N_13582,N_13492,N_13364);
nand U13583 (N_13583,N_13256,N_13357);
nor U13584 (N_13584,N_13415,N_13452);
nor U13585 (N_13585,N_13264,N_13297);
or U13586 (N_13586,N_13274,N_13304);
nand U13587 (N_13587,N_13342,N_13245);
nor U13588 (N_13588,N_13063,N_13467);
nand U13589 (N_13589,N_13086,N_13328);
and U13590 (N_13590,N_13070,N_13066);
or U13591 (N_13591,N_13084,N_13363);
xor U13592 (N_13592,N_13022,N_13170);
and U13593 (N_13593,N_13475,N_13057);
and U13594 (N_13594,N_13273,N_13334);
and U13595 (N_13595,N_13238,N_13159);
nor U13596 (N_13596,N_13294,N_13298);
xnor U13597 (N_13597,N_13302,N_13109);
and U13598 (N_13598,N_13068,N_13450);
and U13599 (N_13599,N_13050,N_13336);
and U13600 (N_13600,N_13279,N_13306);
or U13601 (N_13601,N_13380,N_13491);
nand U13602 (N_13602,N_13268,N_13488);
nor U13603 (N_13603,N_13226,N_13091);
or U13604 (N_13604,N_13424,N_13153);
or U13605 (N_13605,N_13009,N_13431);
nand U13606 (N_13606,N_13004,N_13180);
nor U13607 (N_13607,N_13224,N_13387);
nand U13608 (N_13608,N_13124,N_13186);
and U13609 (N_13609,N_13404,N_13225);
nor U13610 (N_13610,N_13029,N_13398);
or U13611 (N_13611,N_13161,N_13216);
or U13612 (N_13612,N_13411,N_13338);
nand U13613 (N_13613,N_13370,N_13280);
xor U13614 (N_13614,N_13436,N_13486);
nand U13615 (N_13615,N_13242,N_13478);
nor U13616 (N_13616,N_13330,N_13053);
or U13617 (N_13617,N_13098,N_13116);
nor U13618 (N_13618,N_13092,N_13164);
or U13619 (N_13619,N_13323,N_13296);
nand U13620 (N_13620,N_13246,N_13253);
nor U13621 (N_13621,N_13105,N_13027);
nor U13622 (N_13622,N_13456,N_13271);
and U13623 (N_13623,N_13060,N_13189);
nand U13624 (N_13624,N_13209,N_13024);
and U13625 (N_13625,N_13038,N_13104);
nand U13626 (N_13626,N_13231,N_13315);
or U13627 (N_13627,N_13309,N_13046);
and U13628 (N_13628,N_13425,N_13464);
xnor U13629 (N_13629,N_13353,N_13459);
nor U13630 (N_13630,N_13311,N_13171);
xnor U13631 (N_13631,N_13373,N_13151);
xor U13632 (N_13632,N_13345,N_13423);
or U13633 (N_13633,N_13035,N_13386);
or U13634 (N_13634,N_13381,N_13111);
nand U13635 (N_13635,N_13283,N_13300);
nand U13636 (N_13636,N_13290,N_13476);
nand U13637 (N_13637,N_13210,N_13002);
xor U13638 (N_13638,N_13284,N_13206);
nand U13639 (N_13639,N_13292,N_13351);
nand U13640 (N_13640,N_13039,N_13042);
nor U13641 (N_13641,N_13349,N_13099);
nor U13642 (N_13642,N_13078,N_13445);
and U13643 (N_13643,N_13113,N_13341);
xor U13644 (N_13644,N_13434,N_13426);
xor U13645 (N_13645,N_13397,N_13355);
nand U13646 (N_13646,N_13437,N_13457);
or U13647 (N_13647,N_13275,N_13156);
or U13648 (N_13648,N_13453,N_13089);
or U13649 (N_13649,N_13372,N_13401);
or U13650 (N_13650,N_13442,N_13243);
nand U13651 (N_13651,N_13085,N_13394);
and U13652 (N_13652,N_13197,N_13350);
or U13653 (N_13653,N_13371,N_13379);
nand U13654 (N_13654,N_13174,N_13128);
or U13655 (N_13655,N_13101,N_13428);
nand U13656 (N_13656,N_13163,N_13011);
nor U13657 (N_13657,N_13028,N_13120);
nand U13658 (N_13658,N_13277,N_13375);
nor U13659 (N_13659,N_13260,N_13406);
and U13660 (N_13660,N_13183,N_13460);
and U13661 (N_13661,N_13276,N_13454);
or U13662 (N_13662,N_13237,N_13470);
and U13663 (N_13663,N_13026,N_13318);
or U13664 (N_13664,N_13382,N_13477);
and U13665 (N_13665,N_13169,N_13110);
nor U13666 (N_13666,N_13499,N_13474);
nand U13667 (N_13667,N_13054,N_13402);
and U13668 (N_13668,N_13071,N_13408);
nor U13669 (N_13669,N_13250,N_13416);
nor U13670 (N_13670,N_13482,N_13471);
and U13671 (N_13671,N_13007,N_13485);
or U13672 (N_13672,N_13195,N_13146);
nand U13673 (N_13673,N_13337,N_13076);
or U13674 (N_13674,N_13211,N_13137);
and U13675 (N_13675,N_13267,N_13145);
or U13676 (N_13676,N_13443,N_13228);
or U13677 (N_13677,N_13385,N_13016);
and U13678 (N_13678,N_13127,N_13166);
and U13679 (N_13679,N_13208,N_13030);
and U13680 (N_13680,N_13031,N_13272);
or U13681 (N_13681,N_13051,N_13032);
and U13682 (N_13682,N_13198,N_13196);
xor U13683 (N_13683,N_13117,N_13014);
nor U13684 (N_13684,N_13064,N_13252);
nand U13685 (N_13685,N_13044,N_13095);
and U13686 (N_13686,N_13331,N_13259);
nor U13687 (N_13687,N_13067,N_13204);
or U13688 (N_13688,N_13407,N_13429);
nand U13689 (N_13689,N_13012,N_13148);
and U13690 (N_13690,N_13361,N_13093);
or U13691 (N_13691,N_13497,N_13103);
xor U13692 (N_13692,N_13077,N_13286);
xnor U13693 (N_13693,N_13473,N_13081);
nand U13694 (N_13694,N_13003,N_13203);
and U13695 (N_13695,N_13248,N_13378);
nor U13696 (N_13696,N_13138,N_13288);
nor U13697 (N_13697,N_13233,N_13048);
nand U13698 (N_13698,N_13303,N_13390);
and U13699 (N_13699,N_13360,N_13182);
and U13700 (N_13700,N_13114,N_13220);
and U13701 (N_13701,N_13230,N_13155);
or U13702 (N_13702,N_13058,N_13217);
xor U13703 (N_13703,N_13232,N_13299);
nor U13704 (N_13704,N_13005,N_13320);
nand U13705 (N_13705,N_13199,N_13333);
nand U13706 (N_13706,N_13219,N_13392);
nor U13707 (N_13707,N_13389,N_13059);
or U13708 (N_13708,N_13142,N_13254);
nor U13709 (N_13709,N_13194,N_13134);
nand U13710 (N_13710,N_13143,N_13322);
and U13711 (N_13711,N_13034,N_13082);
and U13712 (N_13712,N_13020,N_13158);
nand U13713 (N_13713,N_13412,N_13108);
or U13714 (N_13714,N_13222,N_13440);
or U13715 (N_13715,N_13188,N_13366);
and U13716 (N_13716,N_13123,N_13184);
or U13717 (N_13717,N_13130,N_13495);
and U13718 (N_13718,N_13383,N_13335);
nor U13719 (N_13719,N_13202,N_13396);
nand U13720 (N_13720,N_13362,N_13218);
nand U13721 (N_13721,N_13080,N_13021);
nand U13722 (N_13722,N_13468,N_13462);
and U13723 (N_13723,N_13293,N_13017);
nor U13724 (N_13724,N_13325,N_13083);
nor U13725 (N_13725,N_13121,N_13346);
or U13726 (N_13726,N_13069,N_13348);
nor U13727 (N_13727,N_13281,N_13376);
and U13728 (N_13728,N_13269,N_13493);
nand U13729 (N_13729,N_13227,N_13410);
nand U13730 (N_13730,N_13181,N_13132);
nand U13731 (N_13731,N_13100,N_13176);
xnor U13732 (N_13732,N_13479,N_13047);
nand U13733 (N_13733,N_13344,N_13112);
nand U13734 (N_13734,N_13498,N_13433);
xnor U13735 (N_13735,N_13062,N_13215);
or U13736 (N_13736,N_13096,N_13172);
nor U13737 (N_13737,N_13178,N_13295);
or U13738 (N_13738,N_13446,N_13102);
or U13739 (N_13739,N_13239,N_13236);
nand U13740 (N_13740,N_13356,N_13147);
or U13741 (N_13741,N_13359,N_13200);
or U13742 (N_13742,N_13367,N_13125);
nand U13743 (N_13743,N_13018,N_13319);
nor U13744 (N_13744,N_13008,N_13257);
nand U13745 (N_13745,N_13270,N_13025);
and U13746 (N_13746,N_13049,N_13384);
nand U13747 (N_13747,N_13249,N_13118);
nand U13748 (N_13748,N_13447,N_13214);
nand U13749 (N_13749,N_13168,N_13282);
and U13750 (N_13750,N_13426,N_13080);
nand U13751 (N_13751,N_13384,N_13278);
and U13752 (N_13752,N_13397,N_13275);
nor U13753 (N_13753,N_13339,N_13123);
or U13754 (N_13754,N_13056,N_13219);
and U13755 (N_13755,N_13370,N_13220);
nor U13756 (N_13756,N_13437,N_13455);
or U13757 (N_13757,N_13097,N_13044);
and U13758 (N_13758,N_13311,N_13356);
nor U13759 (N_13759,N_13028,N_13099);
and U13760 (N_13760,N_13005,N_13131);
nand U13761 (N_13761,N_13239,N_13250);
nand U13762 (N_13762,N_13302,N_13238);
xor U13763 (N_13763,N_13216,N_13060);
or U13764 (N_13764,N_13287,N_13308);
or U13765 (N_13765,N_13411,N_13231);
or U13766 (N_13766,N_13370,N_13005);
or U13767 (N_13767,N_13457,N_13103);
and U13768 (N_13768,N_13047,N_13461);
or U13769 (N_13769,N_13087,N_13473);
nor U13770 (N_13770,N_13353,N_13043);
or U13771 (N_13771,N_13467,N_13135);
or U13772 (N_13772,N_13381,N_13414);
nand U13773 (N_13773,N_13109,N_13236);
and U13774 (N_13774,N_13344,N_13176);
nand U13775 (N_13775,N_13268,N_13088);
or U13776 (N_13776,N_13028,N_13043);
nor U13777 (N_13777,N_13225,N_13461);
xnor U13778 (N_13778,N_13211,N_13168);
nor U13779 (N_13779,N_13136,N_13064);
xor U13780 (N_13780,N_13401,N_13229);
nand U13781 (N_13781,N_13286,N_13076);
nor U13782 (N_13782,N_13255,N_13266);
and U13783 (N_13783,N_13387,N_13409);
nor U13784 (N_13784,N_13045,N_13150);
and U13785 (N_13785,N_13206,N_13045);
or U13786 (N_13786,N_13398,N_13367);
or U13787 (N_13787,N_13349,N_13131);
nor U13788 (N_13788,N_13148,N_13303);
nor U13789 (N_13789,N_13408,N_13236);
xnor U13790 (N_13790,N_13046,N_13071);
nor U13791 (N_13791,N_13238,N_13173);
xor U13792 (N_13792,N_13050,N_13350);
xor U13793 (N_13793,N_13105,N_13149);
or U13794 (N_13794,N_13339,N_13069);
nor U13795 (N_13795,N_13388,N_13062);
nor U13796 (N_13796,N_13470,N_13295);
nor U13797 (N_13797,N_13303,N_13431);
or U13798 (N_13798,N_13472,N_13260);
and U13799 (N_13799,N_13351,N_13210);
nand U13800 (N_13800,N_13304,N_13082);
nand U13801 (N_13801,N_13259,N_13117);
nand U13802 (N_13802,N_13394,N_13143);
nand U13803 (N_13803,N_13222,N_13360);
and U13804 (N_13804,N_13026,N_13396);
xor U13805 (N_13805,N_13324,N_13272);
nor U13806 (N_13806,N_13131,N_13285);
and U13807 (N_13807,N_13033,N_13479);
and U13808 (N_13808,N_13342,N_13321);
nand U13809 (N_13809,N_13203,N_13378);
xor U13810 (N_13810,N_13465,N_13364);
nor U13811 (N_13811,N_13444,N_13394);
or U13812 (N_13812,N_13314,N_13095);
or U13813 (N_13813,N_13366,N_13116);
nand U13814 (N_13814,N_13057,N_13322);
nor U13815 (N_13815,N_13236,N_13212);
nand U13816 (N_13816,N_13449,N_13435);
and U13817 (N_13817,N_13175,N_13254);
and U13818 (N_13818,N_13190,N_13456);
and U13819 (N_13819,N_13322,N_13426);
or U13820 (N_13820,N_13411,N_13110);
nand U13821 (N_13821,N_13237,N_13477);
xnor U13822 (N_13822,N_13412,N_13255);
nand U13823 (N_13823,N_13173,N_13148);
and U13824 (N_13824,N_13061,N_13300);
and U13825 (N_13825,N_13267,N_13197);
xor U13826 (N_13826,N_13263,N_13059);
and U13827 (N_13827,N_13380,N_13086);
and U13828 (N_13828,N_13437,N_13472);
xor U13829 (N_13829,N_13160,N_13485);
nand U13830 (N_13830,N_13019,N_13462);
nand U13831 (N_13831,N_13263,N_13447);
nand U13832 (N_13832,N_13139,N_13057);
or U13833 (N_13833,N_13140,N_13096);
and U13834 (N_13834,N_13190,N_13213);
or U13835 (N_13835,N_13369,N_13351);
and U13836 (N_13836,N_13458,N_13019);
or U13837 (N_13837,N_13233,N_13402);
or U13838 (N_13838,N_13304,N_13004);
or U13839 (N_13839,N_13428,N_13491);
nor U13840 (N_13840,N_13410,N_13267);
or U13841 (N_13841,N_13082,N_13462);
or U13842 (N_13842,N_13253,N_13255);
nand U13843 (N_13843,N_13192,N_13346);
nor U13844 (N_13844,N_13481,N_13334);
nand U13845 (N_13845,N_13329,N_13012);
or U13846 (N_13846,N_13128,N_13246);
nor U13847 (N_13847,N_13067,N_13114);
and U13848 (N_13848,N_13304,N_13494);
xor U13849 (N_13849,N_13322,N_13317);
or U13850 (N_13850,N_13491,N_13114);
xnor U13851 (N_13851,N_13386,N_13109);
nor U13852 (N_13852,N_13168,N_13031);
nor U13853 (N_13853,N_13329,N_13041);
nand U13854 (N_13854,N_13205,N_13464);
nand U13855 (N_13855,N_13180,N_13482);
nand U13856 (N_13856,N_13015,N_13251);
nand U13857 (N_13857,N_13416,N_13130);
and U13858 (N_13858,N_13374,N_13453);
nor U13859 (N_13859,N_13443,N_13084);
nand U13860 (N_13860,N_13195,N_13417);
nor U13861 (N_13861,N_13012,N_13101);
or U13862 (N_13862,N_13046,N_13018);
and U13863 (N_13863,N_13236,N_13140);
nand U13864 (N_13864,N_13070,N_13359);
and U13865 (N_13865,N_13098,N_13409);
nor U13866 (N_13866,N_13357,N_13363);
or U13867 (N_13867,N_13248,N_13491);
nor U13868 (N_13868,N_13116,N_13252);
nand U13869 (N_13869,N_13428,N_13448);
or U13870 (N_13870,N_13333,N_13075);
nor U13871 (N_13871,N_13142,N_13038);
or U13872 (N_13872,N_13152,N_13417);
or U13873 (N_13873,N_13404,N_13106);
or U13874 (N_13874,N_13370,N_13367);
and U13875 (N_13875,N_13443,N_13135);
or U13876 (N_13876,N_13323,N_13019);
nand U13877 (N_13877,N_13306,N_13244);
and U13878 (N_13878,N_13416,N_13449);
or U13879 (N_13879,N_13280,N_13467);
nand U13880 (N_13880,N_13161,N_13441);
nor U13881 (N_13881,N_13259,N_13492);
or U13882 (N_13882,N_13299,N_13447);
and U13883 (N_13883,N_13453,N_13019);
and U13884 (N_13884,N_13282,N_13490);
or U13885 (N_13885,N_13246,N_13321);
nor U13886 (N_13886,N_13182,N_13308);
and U13887 (N_13887,N_13437,N_13381);
and U13888 (N_13888,N_13013,N_13444);
nand U13889 (N_13889,N_13166,N_13034);
nand U13890 (N_13890,N_13160,N_13404);
xnor U13891 (N_13891,N_13266,N_13471);
xnor U13892 (N_13892,N_13247,N_13450);
and U13893 (N_13893,N_13440,N_13173);
xnor U13894 (N_13894,N_13406,N_13084);
or U13895 (N_13895,N_13085,N_13320);
or U13896 (N_13896,N_13109,N_13358);
or U13897 (N_13897,N_13035,N_13390);
nand U13898 (N_13898,N_13350,N_13122);
xor U13899 (N_13899,N_13061,N_13109);
and U13900 (N_13900,N_13159,N_13453);
nor U13901 (N_13901,N_13360,N_13086);
or U13902 (N_13902,N_13436,N_13338);
xor U13903 (N_13903,N_13163,N_13242);
nand U13904 (N_13904,N_13278,N_13377);
nor U13905 (N_13905,N_13025,N_13179);
and U13906 (N_13906,N_13148,N_13149);
and U13907 (N_13907,N_13232,N_13229);
nor U13908 (N_13908,N_13228,N_13438);
xor U13909 (N_13909,N_13058,N_13072);
or U13910 (N_13910,N_13328,N_13248);
nand U13911 (N_13911,N_13415,N_13180);
and U13912 (N_13912,N_13369,N_13086);
nand U13913 (N_13913,N_13206,N_13258);
nand U13914 (N_13914,N_13232,N_13007);
nor U13915 (N_13915,N_13237,N_13307);
and U13916 (N_13916,N_13013,N_13033);
or U13917 (N_13917,N_13150,N_13399);
and U13918 (N_13918,N_13323,N_13130);
nand U13919 (N_13919,N_13060,N_13084);
nor U13920 (N_13920,N_13420,N_13347);
or U13921 (N_13921,N_13126,N_13059);
and U13922 (N_13922,N_13079,N_13212);
nor U13923 (N_13923,N_13454,N_13241);
or U13924 (N_13924,N_13251,N_13338);
and U13925 (N_13925,N_13433,N_13412);
and U13926 (N_13926,N_13444,N_13492);
nor U13927 (N_13927,N_13310,N_13170);
nand U13928 (N_13928,N_13281,N_13214);
nor U13929 (N_13929,N_13454,N_13484);
nor U13930 (N_13930,N_13478,N_13092);
nand U13931 (N_13931,N_13202,N_13492);
or U13932 (N_13932,N_13468,N_13492);
nor U13933 (N_13933,N_13070,N_13045);
xnor U13934 (N_13934,N_13245,N_13273);
or U13935 (N_13935,N_13294,N_13153);
and U13936 (N_13936,N_13338,N_13055);
nand U13937 (N_13937,N_13468,N_13249);
nor U13938 (N_13938,N_13265,N_13453);
and U13939 (N_13939,N_13002,N_13484);
xor U13940 (N_13940,N_13303,N_13122);
nand U13941 (N_13941,N_13301,N_13497);
and U13942 (N_13942,N_13423,N_13357);
and U13943 (N_13943,N_13272,N_13052);
or U13944 (N_13944,N_13153,N_13449);
nand U13945 (N_13945,N_13051,N_13035);
or U13946 (N_13946,N_13360,N_13330);
and U13947 (N_13947,N_13482,N_13481);
xor U13948 (N_13948,N_13277,N_13026);
nor U13949 (N_13949,N_13086,N_13354);
nor U13950 (N_13950,N_13295,N_13153);
nor U13951 (N_13951,N_13004,N_13373);
xor U13952 (N_13952,N_13139,N_13408);
or U13953 (N_13953,N_13240,N_13265);
nor U13954 (N_13954,N_13085,N_13040);
nand U13955 (N_13955,N_13397,N_13001);
nor U13956 (N_13956,N_13357,N_13042);
nor U13957 (N_13957,N_13398,N_13358);
nor U13958 (N_13958,N_13393,N_13033);
xor U13959 (N_13959,N_13144,N_13208);
or U13960 (N_13960,N_13183,N_13309);
xor U13961 (N_13961,N_13446,N_13475);
or U13962 (N_13962,N_13032,N_13266);
and U13963 (N_13963,N_13378,N_13099);
nor U13964 (N_13964,N_13446,N_13400);
or U13965 (N_13965,N_13338,N_13280);
nor U13966 (N_13966,N_13387,N_13195);
or U13967 (N_13967,N_13303,N_13147);
nor U13968 (N_13968,N_13478,N_13200);
xnor U13969 (N_13969,N_13404,N_13236);
nand U13970 (N_13970,N_13424,N_13391);
or U13971 (N_13971,N_13077,N_13221);
or U13972 (N_13972,N_13388,N_13314);
nand U13973 (N_13973,N_13033,N_13024);
or U13974 (N_13974,N_13066,N_13092);
and U13975 (N_13975,N_13136,N_13214);
nor U13976 (N_13976,N_13273,N_13380);
or U13977 (N_13977,N_13307,N_13077);
or U13978 (N_13978,N_13478,N_13389);
or U13979 (N_13979,N_13151,N_13069);
xor U13980 (N_13980,N_13096,N_13016);
nor U13981 (N_13981,N_13039,N_13190);
xnor U13982 (N_13982,N_13019,N_13261);
nor U13983 (N_13983,N_13447,N_13471);
or U13984 (N_13984,N_13035,N_13071);
or U13985 (N_13985,N_13173,N_13178);
xnor U13986 (N_13986,N_13487,N_13439);
xor U13987 (N_13987,N_13097,N_13111);
nor U13988 (N_13988,N_13064,N_13200);
nor U13989 (N_13989,N_13004,N_13008);
nor U13990 (N_13990,N_13019,N_13432);
nand U13991 (N_13991,N_13473,N_13025);
or U13992 (N_13992,N_13466,N_13250);
nand U13993 (N_13993,N_13081,N_13335);
nor U13994 (N_13994,N_13322,N_13164);
xor U13995 (N_13995,N_13475,N_13338);
or U13996 (N_13996,N_13289,N_13123);
nor U13997 (N_13997,N_13320,N_13443);
nor U13998 (N_13998,N_13193,N_13218);
nand U13999 (N_13999,N_13476,N_13362);
xnor U14000 (N_14000,N_13911,N_13944);
and U14001 (N_14001,N_13720,N_13607);
xor U14002 (N_14002,N_13792,N_13690);
or U14003 (N_14003,N_13635,N_13500);
nand U14004 (N_14004,N_13817,N_13736);
xor U14005 (N_14005,N_13821,N_13871);
nor U14006 (N_14006,N_13776,N_13676);
or U14007 (N_14007,N_13888,N_13713);
or U14008 (N_14008,N_13518,N_13788);
and U14009 (N_14009,N_13966,N_13722);
xor U14010 (N_14010,N_13598,N_13574);
and U14011 (N_14011,N_13539,N_13924);
or U14012 (N_14012,N_13959,N_13936);
or U14013 (N_14013,N_13809,N_13617);
or U14014 (N_14014,N_13752,N_13850);
nor U14015 (N_14015,N_13648,N_13917);
and U14016 (N_14016,N_13887,N_13560);
nand U14017 (N_14017,N_13655,N_13649);
nand U14018 (N_14018,N_13995,N_13903);
nand U14019 (N_14019,N_13825,N_13775);
nor U14020 (N_14020,N_13869,N_13904);
xor U14021 (N_14021,N_13566,N_13543);
xnor U14022 (N_14022,N_13945,N_13800);
and U14023 (N_14023,N_13663,N_13990);
xor U14024 (N_14024,N_13641,N_13602);
or U14025 (N_14025,N_13643,N_13835);
nand U14026 (N_14026,N_13696,N_13639);
nand U14027 (N_14027,N_13743,N_13831);
xor U14028 (N_14028,N_13734,N_13739);
and U14029 (N_14029,N_13740,N_13544);
nor U14030 (N_14030,N_13787,N_13706);
nand U14031 (N_14031,N_13910,N_13847);
or U14032 (N_14032,N_13731,N_13756);
and U14033 (N_14033,N_13737,N_13719);
nand U14034 (N_14034,N_13926,N_13600);
nand U14035 (N_14035,N_13627,N_13802);
and U14036 (N_14036,N_13953,N_13742);
xor U14037 (N_14037,N_13771,N_13685);
and U14038 (N_14038,N_13630,N_13653);
or U14039 (N_14039,N_13664,N_13813);
nor U14040 (N_14040,N_13625,N_13599);
or U14041 (N_14041,N_13708,N_13781);
or U14042 (N_14042,N_13554,N_13510);
and U14043 (N_14043,N_13662,N_13921);
and U14044 (N_14044,N_13680,N_13609);
nand U14045 (N_14045,N_13986,N_13620);
nand U14046 (N_14046,N_13864,N_13801);
or U14047 (N_14047,N_13933,N_13938);
or U14048 (N_14048,N_13905,N_13750);
or U14049 (N_14049,N_13593,N_13682);
or U14050 (N_14050,N_13583,N_13894);
or U14051 (N_14051,N_13832,N_13795);
and U14052 (N_14052,N_13872,N_13503);
nor U14053 (N_14053,N_13657,N_13533);
nor U14054 (N_14054,N_13928,N_13547);
and U14055 (N_14055,N_13622,N_13614);
nor U14056 (N_14056,N_13803,N_13957);
nor U14057 (N_14057,N_13589,N_13890);
nor U14058 (N_14058,N_13530,N_13954);
and U14059 (N_14059,N_13774,N_13823);
and U14060 (N_14060,N_13666,N_13838);
and U14061 (N_14061,N_13884,N_13816);
and U14062 (N_14062,N_13633,N_13689);
nor U14063 (N_14063,N_13755,N_13845);
or U14064 (N_14064,N_13965,N_13837);
nor U14065 (N_14065,N_13645,N_13853);
or U14066 (N_14066,N_13582,N_13586);
and U14067 (N_14067,N_13697,N_13829);
and U14068 (N_14068,N_13562,N_13519);
and U14069 (N_14069,N_13591,N_13700);
and U14070 (N_14070,N_13857,N_13929);
or U14071 (N_14071,N_13971,N_13947);
and U14072 (N_14072,N_13859,N_13513);
nor U14073 (N_14073,N_13748,N_13906);
and U14074 (N_14074,N_13545,N_13555);
nand U14075 (N_14075,N_13925,N_13727);
and U14076 (N_14076,N_13866,N_13636);
and U14077 (N_14077,N_13932,N_13843);
nor U14078 (N_14078,N_13942,N_13747);
xnor U14079 (N_14079,N_13718,N_13856);
or U14080 (N_14080,N_13794,N_13721);
nand U14081 (N_14081,N_13841,N_13577);
nand U14082 (N_14082,N_13820,N_13749);
and U14083 (N_14083,N_13863,N_13528);
nand U14084 (N_14084,N_13754,N_13671);
and U14085 (N_14085,N_13674,N_13783);
and U14086 (N_14086,N_13818,N_13751);
and U14087 (N_14087,N_13535,N_13652);
and U14088 (N_14088,N_13767,N_13538);
xnor U14089 (N_14089,N_13914,N_13580);
nor U14090 (N_14090,N_13712,N_13879);
nand U14091 (N_14091,N_13961,N_13516);
nor U14092 (N_14092,N_13763,N_13542);
nand U14093 (N_14093,N_13998,N_13684);
and U14094 (N_14094,N_13976,N_13507);
nand U14095 (N_14095,N_13573,N_13908);
nor U14096 (N_14096,N_13793,N_13565);
nor U14097 (N_14097,N_13878,N_13940);
xnor U14098 (N_14098,N_13553,N_13692);
or U14099 (N_14099,N_13753,N_13585);
nor U14100 (N_14100,N_13733,N_13876);
and U14101 (N_14101,N_13806,N_13665);
and U14102 (N_14102,N_13501,N_13717);
xor U14103 (N_14103,N_13515,N_13967);
and U14104 (N_14104,N_13765,N_13812);
xor U14105 (N_14105,N_13670,N_13937);
and U14106 (N_14106,N_13592,N_13564);
nand U14107 (N_14107,N_13703,N_13647);
nor U14108 (N_14108,N_13875,N_13668);
nor U14109 (N_14109,N_13724,N_13999);
nand U14110 (N_14110,N_13907,N_13819);
nand U14111 (N_14111,N_13951,N_13964);
nor U14112 (N_14112,N_13529,N_13939);
nand U14113 (N_14113,N_13993,N_13576);
nor U14114 (N_14114,N_13726,N_13943);
xnor U14115 (N_14115,N_13994,N_13611);
nor U14116 (N_14116,N_13686,N_13968);
nand U14117 (N_14117,N_13842,N_13520);
nand U14118 (N_14118,N_13865,N_13760);
nand U14119 (N_14119,N_13504,N_13891);
nor U14120 (N_14120,N_13658,N_13997);
or U14121 (N_14121,N_13527,N_13762);
and U14122 (N_14122,N_13714,N_13626);
nand U14123 (N_14123,N_13534,N_13672);
xor U14124 (N_14124,N_13561,N_13973);
or U14125 (N_14125,N_13789,N_13766);
nor U14126 (N_14126,N_13855,N_13848);
or U14127 (N_14127,N_13511,N_13950);
nand U14128 (N_14128,N_13590,N_13988);
and U14129 (N_14129,N_13744,N_13930);
xor U14130 (N_14130,N_13764,N_13522);
or U14131 (N_14131,N_13677,N_13741);
nor U14132 (N_14132,N_13920,N_13784);
nor U14133 (N_14133,N_13975,N_13729);
nand U14134 (N_14134,N_13549,N_13735);
or U14135 (N_14135,N_13889,N_13637);
nand U14136 (N_14136,N_13502,N_13579);
and U14137 (N_14137,N_13578,N_13557);
xor U14138 (N_14138,N_13934,N_13524);
nor U14139 (N_14139,N_13723,N_13650);
nand U14140 (N_14140,N_13710,N_13540);
or U14141 (N_14141,N_13667,N_13634);
nor U14142 (N_14142,N_13558,N_13790);
nand U14143 (N_14143,N_13978,N_13769);
nand U14144 (N_14144,N_13517,N_13613);
nand U14145 (N_14145,N_13548,N_13758);
xor U14146 (N_14146,N_13880,N_13615);
nor U14147 (N_14147,N_13526,N_13977);
and U14148 (N_14148,N_13846,N_13605);
nand U14149 (N_14149,N_13892,N_13772);
and U14150 (N_14150,N_13508,N_13777);
nor U14151 (N_14151,N_13900,N_13898);
nand U14152 (N_14152,N_13621,N_13779);
or U14153 (N_14153,N_13631,N_13948);
nand U14154 (N_14154,N_13815,N_13702);
or U14155 (N_14155,N_13509,N_13960);
or U14156 (N_14156,N_13996,N_13824);
and U14157 (N_14157,N_13525,N_13935);
nor U14158 (N_14158,N_13791,N_13985);
nor U14159 (N_14159,N_13551,N_13923);
or U14160 (N_14160,N_13693,N_13572);
nand U14161 (N_14161,N_13896,N_13991);
nor U14162 (N_14162,N_13840,N_13984);
nand U14163 (N_14163,N_13868,N_13883);
nor U14164 (N_14164,N_13646,N_13899);
nand U14165 (N_14165,N_13931,N_13946);
and U14166 (N_14166,N_13567,N_13827);
nand U14167 (N_14167,N_13778,N_13759);
xnor U14168 (N_14168,N_13873,N_13786);
xnor U14169 (N_14169,N_13983,N_13785);
nor U14170 (N_14170,N_13949,N_13808);
nor U14171 (N_14171,N_13974,N_13581);
and U14172 (N_14172,N_13606,N_13707);
and U14173 (N_14173,N_13632,N_13656);
and U14174 (N_14174,N_13955,N_13861);
or U14175 (N_14175,N_13506,N_13768);
or U14176 (N_14176,N_13834,N_13912);
xor U14177 (N_14177,N_13870,N_13698);
or U14178 (N_14178,N_13858,N_13989);
or U14179 (N_14179,N_13669,N_13514);
nor U14180 (N_14180,N_13601,N_13660);
or U14181 (N_14181,N_13862,N_13694);
or U14182 (N_14182,N_13699,N_13780);
nand U14183 (N_14183,N_13550,N_13556);
nand U14184 (N_14184,N_13584,N_13532);
or U14185 (N_14185,N_13570,N_13822);
nand U14186 (N_14186,N_13537,N_13738);
xnor U14187 (N_14187,N_13773,N_13730);
or U14188 (N_14188,N_13716,N_13860);
xor U14189 (N_14189,N_13796,N_13616);
and U14190 (N_14190,N_13770,N_13757);
xor U14191 (N_14191,N_13810,N_13913);
and U14192 (N_14192,N_13597,N_13728);
or U14193 (N_14193,N_13594,N_13797);
nand U14194 (N_14194,N_13987,N_13836);
nand U14195 (N_14195,N_13608,N_13893);
and U14196 (N_14196,N_13683,N_13546);
nor U14197 (N_14197,N_13798,N_13691);
nor U14198 (N_14198,N_13640,N_13512);
or U14199 (N_14199,N_13521,N_13828);
xor U14200 (N_14200,N_13902,N_13732);
nand U14201 (N_14201,N_13575,N_13746);
xnor U14202 (N_14202,N_13814,N_13972);
nand U14203 (N_14203,N_13956,N_13922);
and U14204 (N_14204,N_13919,N_13661);
nand U14205 (N_14205,N_13701,N_13854);
nand U14206 (N_14206,N_13981,N_13624);
nor U14207 (N_14207,N_13619,N_13916);
and U14208 (N_14208,N_13644,N_13839);
or U14209 (N_14209,N_13587,N_13604);
and U14210 (N_14210,N_13612,N_13610);
and U14211 (N_14211,N_13588,N_13963);
nand U14212 (N_14212,N_13895,N_13745);
and U14213 (N_14213,N_13761,N_13688);
nor U14214 (N_14214,N_13559,N_13918);
and U14215 (N_14215,N_13709,N_13886);
nand U14216 (N_14216,N_13958,N_13569);
or U14217 (N_14217,N_13563,N_13941);
nand U14218 (N_14218,N_13830,N_13695);
and U14219 (N_14219,N_13673,N_13711);
and U14220 (N_14220,N_13595,N_13970);
and U14221 (N_14221,N_13603,N_13651);
nor U14222 (N_14222,N_13523,N_13807);
and U14223 (N_14223,N_13629,N_13659);
and U14224 (N_14224,N_13628,N_13505);
nor U14225 (N_14225,N_13867,N_13541);
xnor U14226 (N_14226,N_13571,N_13849);
nand U14227 (N_14227,N_13531,N_13901);
and U14228 (N_14228,N_13799,N_13638);
and U14229 (N_14229,N_13952,N_13852);
nor U14230 (N_14230,N_13704,N_13623);
and U14231 (N_14231,N_13992,N_13678);
and U14232 (N_14232,N_13982,N_13804);
and U14233 (N_14233,N_13654,N_13681);
nand U14234 (N_14234,N_13897,N_13881);
nor U14235 (N_14235,N_13675,N_13874);
nor U14236 (N_14236,N_13536,N_13877);
and U14237 (N_14237,N_13826,N_13882);
and U14238 (N_14238,N_13851,N_13725);
nor U14239 (N_14239,N_13805,N_13642);
and U14240 (N_14240,N_13687,N_13782);
xor U14241 (N_14241,N_13885,N_13844);
nand U14242 (N_14242,N_13927,N_13915);
and U14243 (N_14243,N_13969,N_13552);
nor U14244 (N_14244,N_13811,N_13568);
and U14245 (N_14245,N_13979,N_13618);
or U14246 (N_14246,N_13715,N_13909);
and U14247 (N_14247,N_13962,N_13679);
or U14248 (N_14248,N_13596,N_13705);
and U14249 (N_14249,N_13833,N_13980);
nor U14250 (N_14250,N_13988,N_13547);
nor U14251 (N_14251,N_13623,N_13635);
nand U14252 (N_14252,N_13907,N_13963);
xor U14253 (N_14253,N_13781,N_13501);
nand U14254 (N_14254,N_13955,N_13916);
nor U14255 (N_14255,N_13895,N_13898);
or U14256 (N_14256,N_13909,N_13506);
nand U14257 (N_14257,N_13665,N_13883);
and U14258 (N_14258,N_13651,N_13918);
or U14259 (N_14259,N_13605,N_13899);
nor U14260 (N_14260,N_13781,N_13744);
nand U14261 (N_14261,N_13756,N_13606);
xnor U14262 (N_14262,N_13735,N_13807);
nand U14263 (N_14263,N_13769,N_13665);
or U14264 (N_14264,N_13781,N_13626);
and U14265 (N_14265,N_13752,N_13564);
or U14266 (N_14266,N_13514,N_13602);
xor U14267 (N_14267,N_13980,N_13593);
or U14268 (N_14268,N_13613,N_13707);
nand U14269 (N_14269,N_13903,N_13709);
nand U14270 (N_14270,N_13614,N_13716);
nor U14271 (N_14271,N_13700,N_13545);
xnor U14272 (N_14272,N_13753,N_13584);
and U14273 (N_14273,N_13601,N_13646);
or U14274 (N_14274,N_13521,N_13501);
or U14275 (N_14275,N_13703,N_13852);
and U14276 (N_14276,N_13841,N_13949);
nand U14277 (N_14277,N_13578,N_13584);
and U14278 (N_14278,N_13711,N_13677);
nand U14279 (N_14279,N_13538,N_13937);
and U14280 (N_14280,N_13549,N_13852);
nor U14281 (N_14281,N_13661,N_13625);
and U14282 (N_14282,N_13622,N_13924);
nand U14283 (N_14283,N_13614,N_13962);
nor U14284 (N_14284,N_13694,N_13965);
nand U14285 (N_14285,N_13716,N_13921);
or U14286 (N_14286,N_13953,N_13675);
nor U14287 (N_14287,N_13725,N_13621);
nand U14288 (N_14288,N_13946,N_13512);
nor U14289 (N_14289,N_13792,N_13592);
nand U14290 (N_14290,N_13787,N_13940);
nor U14291 (N_14291,N_13741,N_13711);
nand U14292 (N_14292,N_13717,N_13582);
nor U14293 (N_14293,N_13786,N_13554);
nor U14294 (N_14294,N_13651,N_13878);
nor U14295 (N_14295,N_13754,N_13675);
nand U14296 (N_14296,N_13523,N_13546);
nor U14297 (N_14297,N_13953,N_13939);
and U14298 (N_14298,N_13559,N_13743);
nand U14299 (N_14299,N_13920,N_13516);
nand U14300 (N_14300,N_13826,N_13595);
nand U14301 (N_14301,N_13606,N_13725);
or U14302 (N_14302,N_13617,N_13540);
or U14303 (N_14303,N_13871,N_13560);
and U14304 (N_14304,N_13919,N_13703);
and U14305 (N_14305,N_13524,N_13701);
nor U14306 (N_14306,N_13638,N_13950);
or U14307 (N_14307,N_13616,N_13640);
or U14308 (N_14308,N_13690,N_13563);
or U14309 (N_14309,N_13994,N_13818);
nand U14310 (N_14310,N_13646,N_13678);
nand U14311 (N_14311,N_13749,N_13939);
nor U14312 (N_14312,N_13530,N_13739);
or U14313 (N_14313,N_13667,N_13757);
and U14314 (N_14314,N_13578,N_13742);
or U14315 (N_14315,N_13673,N_13980);
and U14316 (N_14316,N_13557,N_13867);
or U14317 (N_14317,N_13702,N_13708);
or U14318 (N_14318,N_13740,N_13625);
and U14319 (N_14319,N_13608,N_13746);
nor U14320 (N_14320,N_13560,N_13770);
nor U14321 (N_14321,N_13729,N_13585);
and U14322 (N_14322,N_13973,N_13809);
nor U14323 (N_14323,N_13511,N_13895);
or U14324 (N_14324,N_13961,N_13916);
or U14325 (N_14325,N_13771,N_13989);
xor U14326 (N_14326,N_13629,N_13829);
or U14327 (N_14327,N_13505,N_13615);
nor U14328 (N_14328,N_13565,N_13857);
nand U14329 (N_14329,N_13821,N_13697);
nand U14330 (N_14330,N_13809,N_13516);
nor U14331 (N_14331,N_13742,N_13950);
xnor U14332 (N_14332,N_13659,N_13580);
nor U14333 (N_14333,N_13882,N_13538);
and U14334 (N_14334,N_13669,N_13934);
or U14335 (N_14335,N_13556,N_13563);
or U14336 (N_14336,N_13952,N_13788);
xnor U14337 (N_14337,N_13956,N_13994);
or U14338 (N_14338,N_13788,N_13872);
or U14339 (N_14339,N_13745,N_13988);
nor U14340 (N_14340,N_13517,N_13618);
xnor U14341 (N_14341,N_13518,N_13521);
and U14342 (N_14342,N_13928,N_13999);
nor U14343 (N_14343,N_13738,N_13942);
xnor U14344 (N_14344,N_13652,N_13938);
or U14345 (N_14345,N_13611,N_13795);
nor U14346 (N_14346,N_13672,N_13867);
and U14347 (N_14347,N_13559,N_13938);
nand U14348 (N_14348,N_13948,N_13731);
and U14349 (N_14349,N_13515,N_13892);
and U14350 (N_14350,N_13620,N_13904);
or U14351 (N_14351,N_13520,N_13799);
nor U14352 (N_14352,N_13648,N_13729);
or U14353 (N_14353,N_13994,N_13788);
nand U14354 (N_14354,N_13984,N_13952);
or U14355 (N_14355,N_13894,N_13831);
nor U14356 (N_14356,N_13653,N_13800);
nand U14357 (N_14357,N_13611,N_13753);
or U14358 (N_14358,N_13934,N_13816);
nor U14359 (N_14359,N_13560,N_13720);
or U14360 (N_14360,N_13649,N_13876);
xor U14361 (N_14361,N_13858,N_13735);
and U14362 (N_14362,N_13567,N_13690);
nand U14363 (N_14363,N_13723,N_13856);
nor U14364 (N_14364,N_13553,N_13702);
or U14365 (N_14365,N_13893,N_13993);
nand U14366 (N_14366,N_13609,N_13957);
nor U14367 (N_14367,N_13814,N_13614);
or U14368 (N_14368,N_13556,N_13747);
and U14369 (N_14369,N_13887,N_13801);
and U14370 (N_14370,N_13630,N_13700);
xnor U14371 (N_14371,N_13972,N_13989);
and U14372 (N_14372,N_13677,N_13892);
or U14373 (N_14373,N_13619,N_13602);
xnor U14374 (N_14374,N_13850,N_13606);
and U14375 (N_14375,N_13546,N_13947);
nand U14376 (N_14376,N_13936,N_13572);
or U14377 (N_14377,N_13923,N_13566);
nand U14378 (N_14378,N_13624,N_13656);
or U14379 (N_14379,N_13850,N_13904);
nor U14380 (N_14380,N_13729,N_13780);
and U14381 (N_14381,N_13956,N_13619);
nor U14382 (N_14382,N_13693,N_13855);
nand U14383 (N_14383,N_13622,N_13731);
and U14384 (N_14384,N_13911,N_13929);
nor U14385 (N_14385,N_13841,N_13919);
and U14386 (N_14386,N_13786,N_13596);
nor U14387 (N_14387,N_13791,N_13523);
and U14388 (N_14388,N_13955,N_13624);
or U14389 (N_14389,N_13854,N_13839);
nor U14390 (N_14390,N_13723,N_13566);
and U14391 (N_14391,N_13564,N_13964);
nor U14392 (N_14392,N_13858,N_13617);
nor U14393 (N_14393,N_13550,N_13601);
and U14394 (N_14394,N_13777,N_13589);
xnor U14395 (N_14395,N_13956,N_13558);
or U14396 (N_14396,N_13778,N_13584);
and U14397 (N_14397,N_13561,N_13727);
nor U14398 (N_14398,N_13501,N_13853);
or U14399 (N_14399,N_13681,N_13840);
or U14400 (N_14400,N_13822,N_13726);
nand U14401 (N_14401,N_13759,N_13549);
xor U14402 (N_14402,N_13830,N_13988);
and U14403 (N_14403,N_13869,N_13856);
or U14404 (N_14404,N_13893,N_13953);
nand U14405 (N_14405,N_13580,N_13594);
nor U14406 (N_14406,N_13605,N_13520);
and U14407 (N_14407,N_13709,N_13817);
nand U14408 (N_14408,N_13809,N_13695);
nor U14409 (N_14409,N_13702,N_13607);
nand U14410 (N_14410,N_13839,N_13778);
nand U14411 (N_14411,N_13699,N_13537);
nand U14412 (N_14412,N_13739,N_13811);
nand U14413 (N_14413,N_13648,N_13527);
and U14414 (N_14414,N_13803,N_13653);
nand U14415 (N_14415,N_13721,N_13651);
or U14416 (N_14416,N_13542,N_13511);
nand U14417 (N_14417,N_13679,N_13769);
or U14418 (N_14418,N_13760,N_13634);
xnor U14419 (N_14419,N_13939,N_13513);
or U14420 (N_14420,N_13990,N_13830);
nor U14421 (N_14421,N_13881,N_13960);
nand U14422 (N_14422,N_13715,N_13660);
or U14423 (N_14423,N_13609,N_13509);
and U14424 (N_14424,N_13674,N_13827);
nor U14425 (N_14425,N_13514,N_13825);
nand U14426 (N_14426,N_13710,N_13962);
and U14427 (N_14427,N_13977,N_13736);
and U14428 (N_14428,N_13578,N_13561);
and U14429 (N_14429,N_13572,N_13680);
and U14430 (N_14430,N_13775,N_13636);
or U14431 (N_14431,N_13836,N_13848);
or U14432 (N_14432,N_13707,N_13533);
nand U14433 (N_14433,N_13862,N_13839);
or U14434 (N_14434,N_13750,N_13609);
or U14435 (N_14435,N_13982,N_13559);
and U14436 (N_14436,N_13828,N_13596);
or U14437 (N_14437,N_13584,N_13745);
nor U14438 (N_14438,N_13566,N_13812);
nand U14439 (N_14439,N_13540,N_13789);
and U14440 (N_14440,N_13769,N_13681);
nand U14441 (N_14441,N_13777,N_13837);
or U14442 (N_14442,N_13771,N_13870);
and U14443 (N_14443,N_13921,N_13543);
nor U14444 (N_14444,N_13851,N_13835);
and U14445 (N_14445,N_13712,N_13634);
nand U14446 (N_14446,N_13825,N_13609);
and U14447 (N_14447,N_13543,N_13524);
nand U14448 (N_14448,N_13750,N_13956);
or U14449 (N_14449,N_13582,N_13646);
nand U14450 (N_14450,N_13783,N_13550);
nor U14451 (N_14451,N_13790,N_13576);
or U14452 (N_14452,N_13556,N_13629);
nor U14453 (N_14453,N_13574,N_13717);
and U14454 (N_14454,N_13591,N_13742);
nor U14455 (N_14455,N_13508,N_13647);
nor U14456 (N_14456,N_13680,N_13573);
or U14457 (N_14457,N_13762,N_13815);
or U14458 (N_14458,N_13652,N_13624);
and U14459 (N_14459,N_13544,N_13734);
or U14460 (N_14460,N_13633,N_13711);
or U14461 (N_14461,N_13672,N_13763);
or U14462 (N_14462,N_13974,N_13754);
nand U14463 (N_14463,N_13587,N_13730);
and U14464 (N_14464,N_13679,N_13845);
nand U14465 (N_14465,N_13536,N_13691);
xor U14466 (N_14466,N_13715,N_13698);
and U14467 (N_14467,N_13766,N_13980);
xor U14468 (N_14468,N_13601,N_13543);
nor U14469 (N_14469,N_13976,N_13828);
or U14470 (N_14470,N_13935,N_13556);
or U14471 (N_14471,N_13844,N_13736);
xnor U14472 (N_14472,N_13953,N_13760);
or U14473 (N_14473,N_13560,N_13730);
and U14474 (N_14474,N_13672,N_13757);
nor U14475 (N_14475,N_13785,N_13781);
nor U14476 (N_14476,N_13574,N_13894);
nand U14477 (N_14477,N_13706,N_13577);
or U14478 (N_14478,N_13617,N_13584);
nand U14479 (N_14479,N_13823,N_13684);
and U14480 (N_14480,N_13986,N_13916);
nand U14481 (N_14481,N_13643,N_13633);
nand U14482 (N_14482,N_13613,N_13784);
nor U14483 (N_14483,N_13866,N_13796);
nand U14484 (N_14484,N_13526,N_13701);
nand U14485 (N_14485,N_13548,N_13876);
or U14486 (N_14486,N_13800,N_13926);
and U14487 (N_14487,N_13906,N_13505);
nor U14488 (N_14488,N_13972,N_13704);
and U14489 (N_14489,N_13659,N_13911);
xor U14490 (N_14490,N_13684,N_13746);
nand U14491 (N_14491,N_13857,N_13721);
nand U14492 (N_14492,N_13810,N_13875);
nand U14493 (N_14493,N_13534,N_13816);
and U14494 (N_14494,N_13616,N_13988);
and U14495 (N_14495,N_13550,N_13554);
or U14496 (N_14496,N_13840,N_13954);
nor U14497 (N_14497,N_13987,N_13542);
and U14498 (N_14498,N_13925,N_13526);
nand U14499 (N_14499,N_13868,N_13661);
xor U14500 (N_14500,N_14000,N_14308);
or U14501 (N_14501,N_14170,N_14208);
nand U14502 (N_14502,N_14090,N_14388);
nor U14503 (N_14503,N_14318,N_14031);
nand U14504 (N_14504,N_14212,N_14316);
xnor U14505 (N_14505,N_14322,N_14264);
nor U14506 (N_14506,N_14106,N_14013);
nor U14507 (N_14507,N_14156,N_14373);
nor U14508 (N_14508,N_14133,N_14287);
nor U14509 (N_14509,N_14176,N_14047);
nor U14510 (N_14510,N_14074,N_14005);
nand U14511 (N_14511,N_14096,N_14159);
nand U14512 (N_14512,N_14243,N_14128);
xnor U14513 (N_14513,N_14335,N_14069);
xor U14514 (N_14514,N_14481,N_14216);
nand U14515 (N_14515,N_14048,N_14489);
and U14516 (N_14516,N_14344,N_14405);
and U14517 (N_14517,N_14493,N_14366);
nor U14518 (N_14518,N_14068,N_14294);
or U14519 (N_14519,N_14398,N_14153);
nor U14520 (N_14520,N_14122,N_14396);
or U14521 (N_14521,N_14166,N_14129);
and U14522 (N_14522,N_14420,N_14094);
nor U14523 (N_14523,N_14260,N_14435);
nor U14524 (N_14524,N_14228,N_14446);
and U14525 (N_14525,N_14203,N_14223);
nor U14526 (N_14526,N_14175,N_14102);
xnor U14527 (N_14527,N_14340,N_14075);
nand U14528 (N_14528,N_14401,N_14080);
nor U14529 (N_14529,N_14342,N_14281);
nor U14530 (N_14530,N_14444,N_14361);
xor U14531 (N_14531,N_14247,N_14189);
nand U14532 (N_14532,N_14236,N_14311);
or U14533 (N_14533,N_14169,N_14032);
or U14534 (N_14534,N_14227,N_14440);
or U14535 (N_14535,N_14393,N_14462);
or U14536 (N_14536,N_14455,N_14417);
nor U14537 (N_14537,N_14130,N_14015);
and U14538 (N_14538,N_14450,N_14134);
nor U14539 (N_14539,N_14254,N_14055);
or U14540 (N_14540,N_14498,N_14265);
nand U14541 (N_14541,N_14317,N_14154);
and U14542 (N_14542,N_14268,N_14171);
nand U14543 (N_14543,N_14028,N_14418);
nor U14544 (N_14544,N_14306,N_14319);
xor U14545 (N_14545,N_14496,N_14123);
nor U14546 (N_14546,N_14321,N_14365);
or U14547 (N_14547,N_14407,N_14201);
or U14548 (N_14548,N_14249,N_14363);
or U14549 (N_14549,N_14266,N_14488);
nor U14550 (N_14550,N_14165,N_14136);
or U14551 (N_14551,N_14400,N_14109);
nor U14552 (N_14552,N_14390,N_14021);
and U14553 (N_14553,N_14095,N_14379);
nand U14554 (N_14554,N_14395,N_14067);
nor U14555 (N_14555,N_14033,N_14275);
nand U14556 (N_14556,N_14168,N_14486);
nand U14557 (N_14557,N_14235,N_14354);
or U14558 (N_14558,N_14377,N_14037);
or U14559 (N_14559,N_14043,N_14297);
and U14560 (N_14560,N_14160,N_14359);
nor U14561 (N_14561,N_14362,N_14392);
nor U14562 (N_14562,N_14477,N_14060);
or U14563 (N_14563,N_14118,N_14448);
or U14564 (N_14564,N_14066,N_14412);
and U14565 (N_14565,N_14050,N_14052);
and U14566 (N_14566,N_14181,N_14231);
or U14567 (N_14567,N_14424,N_14269);
nor U14568 (N_14568,N_14439,N_14480);
xor U14569 (N_14569,N_14002,N_14022);
or U14570 (N_14570,N_14167,N_14023);
xnor U14571 (N_14571,N_14107,N_14191);
and U14572 (N_14572,N_14332,N_14429);
nand U14573 (N_14573,N_14330,N_14471);
and U14574 (N_14574,N_14177,N_14326);
nor U14575 (N_14575,N_14325,N_14456);
or U14576 (N_14576,N_14045,N_14034);
and U14577 (N_14577,N_14397,N_14183);
and U14578 (N_14578,N_14232,N_14428);
or U14579 (N_14579,N_14084,N_14447);
nor U14580 (N_14580,N_14026,N_14152);
and U14581 (N_14581,N_14125,N_14086);
or U14582 (N_14582,N_14234,N_14105);
and U14583 (N_14583,N_14020,N_14280);
or U14584 (N_14584,N_14196,N_14089);
or U14585 (N_14585,N_14409,N_14229);
and U14586 (N_14586,N_14058,N_14030);
or U14587 (N_14587,N_14327,N_14202);
or U14588 (N_14588,N_14070,N_14441);
nor U14589 (N_14589,N_14483,N_14126);
nand U14590 (N_14590,N_14091,N_14162);
or U14591 (N_14591,N_14082,N_14451);
nand U14592 (N_14592,N_14194,N_14059);
nand U14593 (N_14593,N_14436,N_14230);
nor U14594 (N_14594,N_14193,N_14301);
or U14595 (N_14595,N_14427,N_14284);
nand U14596 (N_14596,N_14348,N_14163);
and U14597 (N_14597,N_14073,N_14346);
or U14598 (N_14598,N_14180,N_14206);
nor U14599 (N_14599,N_14272,N_14256);
or U14600 (N_14600,N_14215,N_14277);
or U14601 (N_14601,N_14367,N_14200);
nor U14602 (N_14602,N_14088,N_14300);
nand U14603 (N_14603,N_14112,N_14410);
nor U14604 (N_14604,N_14357,N_14271);
nand U14605 (N_14605,N_14046,N_14233);
or U14606 (N_14606,N_14380,N_14411);
and U14607 (N_14607,N_14452,N_14083);
nor U14608 (N_14608,N_14298,N_14085);
nand U14609 (N_14609,N_14419,N_14413);
nand U14610 (N_14610,N_14001,N_14328);
or U14611 (N_14611,N_14111,N_14282);
xor U14612 (N_14612,N_14329,N_14484);
or U14613 (N_14613,N_14334,N_14238);
xnor U14614 (N_14614,N_14057,N_14150);
or U14615 (N_14615,N_14053,N_14261);
nand U14616 (N_14616,N_14063,N_14182);
nand U14617 (N_14617,N_14173,N_14278);
or U14618 (N_14618,N_14144,N_14077);
nor U14619 (N_14619,N_14350,N_14101);
or U14620 (N_14620,N_14198,N_14010);
or U14621 (N_14621,N_14119,N_14352);
or U14622 (N_14622,N_14469,N_14376);
or U14623 (N_14623,N_14141,N_14262);
nor U14624 (N_14624,N_14092,N_14197);
nand U14625 (N_14625,N_14437,N_14042);
xor U14626 (N_14626,N_14024,N_14087);
or U14627 (N_14627,N_14104,N_14127);
xnor U14628 (N_14628,N_14039,N_14349);
or U14629 (N_14629,N_14267,N_14474);
nor U14630 (N_14630,N_14360,N_14495);
or U14631 (N_14631,N_14103,N_14185);
or U14632 (N_14632,N_14081,N_14378);
and U14633 (N_14633,N_14382,N_14093);
nor U14634 (N_14634,N_14237,N_14273);
or U14635 (N_14635,N_14078,N_14384);
or U14636 (N_14636,N_14064,N_14072);
nor U14637 (N_14637,N_14252,N_14255);
or U14638 (N_14638,N_14291,N_14218);
nor U14639 (N_14639,N_14210,N_14224);
nand U14640 (N_14640,N_14414,N_14140);
nor U14641 (N_14641,N_14345,N_14178);
nand U14642 (N_14642,N_14394,N_14259);
and U14643 (N_14643,N_14099,N_14009);
or U14644 (N_14644,N_14114,N_14044);
or U14645 (N_14645,N_14290,N_14463);
nor U14646 (N_14646,N_14250,N_14494);
and U14647 (N_14647,N_14475,N_14116);
and U14648 (N_14648,N_14422,N_14131);
and U14649 (N_14649,N_14027,N_14383);
or U14650 (N_14650,N_14460,N_14204);
and U14651 (N_14651,N_14149,N_14312);
nor U14652 (N_14652,N_14399,N_14056);
or U14653 (N_14653,N_14406,N_14161);
and U14654 (N_14654,N_14041,N_14347);
nand U14655 (N_14655,N_14304,N_14097);
and U14656 (N_14656,N_14246,N_14324);
or U14657 (N_14657,N_14192,N_14421);
and U14658 (N_14658,N_14226,N_14211);
or U14659 (N_14659,N_14497,N_14302);
nor U14660 (N_14660,N_14241,N_14184);
and U14661 (N_14661,N_14117,N_14370);
and U14662 (N_14662,N_14222,N_14356);
or U14663 (N_14663,N_14019,N_14295);
nor U14664 (N_14664,N_14214,N_14387);
nor U14665 (N_14665,N_14257,N_14408);
nor U14666 (N_14666,N_14008,N_14479);
nor U14667 (N_14667,N_14458,N_14142);
nor U14668 (N_14668,N_14014,N_14213);
or U14669 (N_14669,N_14016,N_14155);
or U14670 (N_14670,N_14240,N_14485);
nand U14671 (N_14671,N_14385,N_14470);
nor U14672 (N_14672,N_14248,N_14336);
nand U14673 (N_14673,N_14017,N_14425);
nand U14674 (N_14674,N_14431,N_14217);
nor U14675 (N_14675,N_14003,N_14110);
nor U14676 (N_14676,N_14061,N_14416);
nand U14677 (N_14677,N_14006,N_14098);
or U14678 (N_14678,N_14239,N_14415);
nor U14679 (N_14679,N_14279,N_14333);
or U14680 (N_14680,N_14146,N_14369);
or U14681 (N_14681,N_14449,N_14157);
nor U14682 (N_14682,N_14205,N_14179);
nand U14683 (N_14683,N_14432,N_14286);
nand U14684 (N_14684,N_14219,N_14465);
nand U14685 (N_14685,N_14310,N_14358);
or U14686 (N_14686,N_14426,N_14403);
xnor U14687 (N_14687,N_14274,N_14076);
and U14688 (N_14688,N_14423,N_14151);
nor U14689 (N_14689,N_14147,N_14276);
or U14690 (N_14690,N_14468,N_14079);
nor U14691 (N_14691,N_14391,N_14012);
and U14692 (N_14692,N_14476,N_14351);
and U14693 (N_14693,N_14371,N_14386);
nand U14694 (N_14694,N_14338,N_14314);
or U14695 (N_14695,N_14186,N_14018);
nand U14696 (N_14696,N_14374,N_14137);
nor U14697 (N_14697,N_14457,N_14207);
or U14698 (N_14698,N_14195,N_14011);
xor U14699 (N_14699,N_14035,N_14296);
or U14700 (N_14700,N_14158,N_14253);
xor U14701 (N_14701,N_14491,N_14199);
nor U14702 (N_14702,N_14454,N_14364);
and U14703 (N_14703,N_14124,N_14445);
or U14704 (N_14704,N_14375,N_14049);
nor U14705 (N_14705,N_14353,N_14190);
and U14706 (N_14706,N_14453,N_14487);
xor U14707 (N_14707,N_14040,N_14478);
nand U14708 (N_14708,N_14490,N_14289);
nand U14709 (N_14709,N_14341,N_14025);
nand U14710 (N_14710,N_14442,N_14270);
or U14711 (N_14711,N_14389,N_14309);
or U14712 (N_14712,N_14355,N_14120);
nand U14713 (N_14713,N_14292,N_14004);
or U14714 (N_14714,N_14062,N_14138);
xor U14715 (N_14715,N_14293,N_14135);
xnor U14716 (N_14716,N_14473,N_14459);
or U14717 (N_14717,N_14029,N_14434);
or U14718 (N_14718,N_14339,N_14285);
nor U14719 (N_14719,N_14115,N_14404);
and U14720 (N_14720,N_14258,N_14221);
or U14721 (N_14721,N_14172,N_14209);
nor U14722 (N_14722,N_14307,N_14499);
or U14723 (N_14723,N_14121,N_14283);
nand U14724 (N_14724,N_14132,N_14225);
nand U14725 (N_14725,N_14220,N_14472);
xor U14726 (N_14726,N_14461,N_14337);
or U14727 (N_14727,N_14054,N_14164);
nor U14728 (N_14728,N_14482,N_14313);
and U14729 (N_14729,N_14108,N_14036);
nand U14730 (N_14730,N_14242,N_14148);
or U14731 (N_14731,N_14251,N_14343);
nand U14732 (N_14732,N_14433,N_14143);
and U14733 (N_14733,N_14113,N_14305);
and U14734 (N_14734,N_14303,N_14065);
nor U14735 (N_14735,N_14299,N_14139);
and U14736 (N_14736,N_14466,N_14438);
xor U14737 (N_14737,N_14007,N_14372);
or U14738 (N_14738,N_14430,N_14244);
xnor U14739 (N_14739,N_14315,N_14331);
and U14740 (N_14740,N_14381,N_14402);
and U14741 (N_14741,N_14038,N_14174);
nand U14742 (N_14742,N_14492,N_14368);
or U14743 (N_14743,N_14443,N_14320);
nand U14744 (N_14744,N_14288,N_14145);
nor U14745 (N_14745,N_14071,N_14100);
or U14746 (N_14746,N_14188,N_14245);
and U14747 (N_14747,N_14263,N_14467);
and U14748 (N_14748,N_14051,N_14187);
nand U14749 (N_14749,N_14464,N_14323);
or U14750 (N_14750,N_14029,N_14337);
nand U14751 (N_14751,N_14106,N_14104);
xor U14752 (N_14752,N_14079,N_14028);
nor U14753 (N_14753,N_14078,N_14040);
nor U14754 (N_14754,N_14378,N_14004);
nand U14755 (N_14755,N_14077,N_14258);
and U14756 (N_14756,N_14280,N_14039);
and U14757 (N_14757,N_14065,N_14299);
or U14758 (N_14758,N_14374,N_14192);
nor U14759 (N_14759,N_14295,N_14283);
or U14760 (N_14760,N_14010,N_14256);
nor U14761 (N_14761,N_14186,N_14137);
or U14762 (N_14762,N_14148,N_14372);
nand U14763 (N_14763,N_14002,N_14255);
and U14764 (N_14764,N_14033,N_14110);
and U14765 (N_14765,N_14209,N_14085);
nand U14766 (N_14766,N_14324,N_14392);
or U14767 (N_14767,N_14066,N_14395);
and U14768 (N_14768,N_14488,N_14143);
xnor U14769 (N_14769,N_14027,N_14180);
xnor U14770 (N_14770,N_14222,N_14066);
or U14771 (N_14771,N_14107,N_14054);
and U14772 (N_14772,N_14377,N_14178);
nand U14773 (N_14773,N_14403,N_14276);
nand U14774 (N_14774,N_14396,N_14385);
nor U14775 (N_14775,N_14203,N_14293);
xor U14776 (N_14776,N_14438,N_14462);
and U14777 (N_14777,N_14034,N_14303);
nor U14778 (N_14778,N_14011,N_14091);
nor U14779 (N_14779,N_14017,N_14087);
or U14780 (N_14780,N_14443,N_14199);
and U14781 (N_14781,N_14140,N_14126);
and U14782 (N_14782,N_14357,N_14062);
and U14783 (N_14783,N_14467,N_14299);
or U14784 (N_14784,N_14179,N_14242);
nand U14785 (N_14785,N_14413,N_14421);
nor U14786 (N_14786,N_14219,N_14249);
and U14787 (N_14787,N_14422,N_14029);
and U14788 (N_14788,N_14202,N_14034);
or U14789 (N_14789,N_14083,N_14330);
nand U14790 (N_14790,N_14092,N_14051);
and U14791 (N_14791,N_14441,N_14285);
and U14792 (N_14792,N_14499,N_14169);
nor U14793 (N_14793,N_14134,N_14463);
nand U14794 (N_14794,N_14231,N_14461);
nor U14795 (N_14795,N_14103,N_14046);
and U14796 (N_14796,N_14201,N_14196);
and U14797 (N_14797,N_14109,N_14224);
nand U14798 (N_14798,N_14278,N_14003);
nor U14799 (N_14799,N_14293,N_14224);
or U14800 (N_14800,N_14071,N_14316);
and U14801 (N_14801,N_14301,N_14063);
nor U14802 (N_14802,N_14432,N_14124);
nor U14803 (N_14803,N_14007,N_14114);
nand U14804 (N_14804,N_14249,N_14088);
nor U14805 (N_14805,N_14117,N_14263);
and U14806 (N_14806,N_14144,N_14424);
and U14807 (N_14807,N_14450,N_14098);
nand U14808 (N_14808,N_14052,N_14053);
nand U14809 (N_14809,N_14037,N_14066);
and U14810 (N_14810,N_14041,N_14068);
nor U14811 (N_14811,N_14018,N_14215);
xnor U14812 (N_14812,N_14143,N_14096);
and U14813 (N_14813,N_14295,N_14051);
nand U14814 (N_14814,N_14086,N_14149);
xnor U14815 (N_14815,N_14484,N_14295);
and U14816 (N_14816,N_14147,N_14436);
xor U14817 (N_14817,N_14314,N_14429);
xnor U14818 (N_14818,N_14463,N_14250);
nand U14819 (N_14819,N_14283,N_14091);
or U14820 (N_14820,N_14380,N_14227);
or U14821 (N_14821,N_14429,N_14252);
nand U14822 (N_14822,N_14114,N_14288);
xor U14823 (N_14823,N_14075,N_14213);
xnor U14824 (N_14824,N_14004,N_14454);
or U14825 (N_14825,N_14266,N_14064);
nor U14826 (N_14826,N_14278,N_14425);
and U14827 (N_14827,N_14387,N_14004);
nand U14828 (N_14828,N_14083,N_14025);
and U14829 (N_14829,N_14325,N_14218);
nand U14830 (N_14830,N_14289,N_14438);
or U14831 (N_14831,N_14400,N_14163);
and U14832 (N_14832,N_14291,N_14043);
and U14833 (N_14833,N_14103,N_14038);
nor U14834 (N_14834,N_14335,N_14240);
nand U14835 (N_14835,N_14055,N_14092);
nand U14836 (N_14836,N_14166,N_14235);
nand U14837 (N_14837,N_14072,N_14086);
and U14838 (N_14838,N_14249,N_14489);
and U14839 (N_14839,N_14339,N_14363);
and U14840 (N_14840,N_14140,N_14018);
or U14841 (N_14841,N_14401,N_14106);
nor U14842 (N_14842,N_14384,N_14167);
nor U14843 (N_14843,N_14213,N_14438);
nor U14844 (N_14844,N_14054,N_14403);
nand U14845 (N_14845,N_14278,N_14399);
and U14846 (N_14846,N_14495,N_14402);
and U14847 (N_14847,N_14220,N_14484);
nor U14848 (N_14848,N_14146,N_14498);
nor U14849 (N_14849,N_14166,N_14338);
nor U14850 (N_14850,N_14090,N_14178);
nand U14851 (N_14851,N_14215,N_14377);
nand U14852 (N_14852,N_14027,N_14264);
nand U14853 (N_14853,N_14407,N_14047);
and U14854 (N_14854,N_14399,N_14086);
and U14855 (N_14855,N_14407,N_14101);
or U14856 (N_14856,N_14243,N_14497);
nand U14857 (N_14857,N_14059,N_14188);
nor U14858 (N_14858,N_14491,N_14382);
and U14859 (N_14859,N_14128,N_14299);
nor U14860 (N_14860,N_14010,N_14145);
and U14861 (N_14861,N_14008,N_14016);
nor U14862 (N_14862,N_14482,N_14132);
or U14863 (N_14863,N_14445,N_14055);
and U14864 (N_14864,N_14336,N_14005);
and U14865 (N_14865,N_14266,N_14414);
nand U14866 (N_14866,N_14439,N_14098);
or U14867 (N_14867,N_14369,N_14046);
xnor U14868 (N_14868,N_14297,N_14199);
or U14869 (N_14869,N_14253,N_14388);
xnor U14870 (N_14870,N_14050,N_14145);
nand U14871 (N_14871,N_14177,N_14234);
or U14872 (N_14872,N_14247,N_14150);
nor U14873 (N_14873,N_14224,N_14073);
or U14874 (N_14874,N_14468,N_14278);
and U14875 (N_14875,N_14350,N_14134);
and U14876 (N_14876,N_14499,N_14074);
or U14877 (N_14877,N_14155,N_14312);
nand U14878 (N_14878,N_14473,N_14234);
and U14879 (N_14879,N_14240,N_14444);
nand U14880 (N_14880,N_14105,N_14361);
nor U14881 (N_14881,N_14400,N_14030);
nand U14882 (N_14882,N_14295,N_14014);
nand U14883 (N_14883,N_14010,N_14333);
nand U14884 (N_14884,N_14134,N_14412);
xor U14885 (N_14885,N_14468,N_14119);
and U14886 (N_14886,N_14111,N_14197);
nand U14887 (N_14887,N_14139,N_14272);
nand U14888 (N_14888,N_14158,N_14216);
nand U14889 (N_14889,N_14480,N_14450);
nor U14890 (N_14890,N_14027,N_14256);
xor U14891 (N_14891,N_14131,N_14356);
or U14892 (N_14892,N_14416,N_14172);
or U14893 (N_14893,N_14414,N_14420);
and U14894 (N_14894,N_14391,N_14402);
nand U14895 (N_14895,N_14299,N_14328);
or U14896 (N_14896,N_14436,N_14014);
and U14897 (N_14897,N_14005,N_14454);
nor U14898 (N_14898,N_14385,N_14156);
nor U14899 (N_14899,N_14069,N_14382);
and U14900 (N_14900,N_14164,N_14498);
xnor U14901 (N_14901,N_14073,N_14271);
nand U14902 (N_14902,N_14083,N_14343);
xnor U14903 (N_14903,N_14465,N_14442);
nand U14904 (N_14904,N_14345,N_14064);
nand U14905 (N_14905,N_14363,N_14476);
or U14906 (N_14906,N_14330,N_14222);
nand U14907 (N_14907,N_14347,N_14155);
nor U14908 (N_14908,N_14428,N_14197);
and U14909 (N_14909,N_14081,N_14468);
and U14910 (N_14910,N_14327,N_14208);
nand U14911 (N_14911,N_14124,N_14387);
nor U14912 (N_14912,N_14410,N_14190);
or U14913 (N_14913,N_14215,N_14143);
nand U14914 (N_14914,N_14321,N_14076);
nand U14915 (N_14915,N_14357,N_14218);
nor U14916 (N_14916,N_14435,N_14441);
xor U14917 (N_14917,N_14136,N_14234);
nand U14918 (N_14918,N_14364,N_14191);
nor U14919 (N_14919,N_14080,N_14094);
nand U14920 (N_14920,N_14186,N_14158);
or U14921 (N_14921,N_14247,N_14283);
nand U14922 (N_14922,N_14198,N_14372);
and U14923 (N_14923,N_14233,N_14191);
or U14924 (N_14924,N_14221,N_14323);
and U14925 (N_14925,N_14134,N_14348);
and U14926 (N_14926,N_14088,N_14168);
and U14927 (N_14927,N_14087,N_14003);
or U14928 (N_14928,N_14050,N_14249);
nor U14929 (N_14929,N_14262,N_14249);
nor U14930 (N_14930,N_14138,N_14257);
nor U14931 (N_14931,N_14108,N_14349);
or U14932 (N_14932,N_14178,N_14458);
xnor U14933 (N_14933,N_14215,N_14456);
nor U14934 (N_14934,N_14189,N_14121);
or U14935 (N_14935,N_14069,N_14312);
or U14936 (N_14936,N_14005,N_14186);
or U14937 (N_14937,N_14465,N_14431);
nor U14938 (N_14938,N_14390,N_14308);
and U14939 (N_14939,N_14183,N_14495);
nand U14940 (N_14940,N_14051,N_14151);
xnor U14941 (N_14941,N_14358,N_14143);
or U14942 (N_14942,N_14463,N_14477);
or U14943 (N_14943,N_14454,N_14146);
and U14944 (N_14944,N_14231,N_14026);
nor U14945 (N_14945,N_14422,N_14400);
and U14946 (N_14946,N_14086,N_14005);
nor U14947 (N_14947,N_14254,N_14386);
or U14948 (N_14948,N_14020,N_14093);
nand U14949 (N_14949,N_14422,N_14185);
or U14950 (N_14950,N_14441,N_14432);
nor U14951 (N_14951,N_14019,N_14495);
or U14952 (N_14952,N_14128,N_14176);
nand U14953 (N_14953,N_14360,N_14090);
or U14954 (N_14954,N_14201,N_14436);
or U14955 (N_14955,N_14036,N_14223);
nand U14956 (N_14956,N_14328,N_14199);
nor U14957 (N_14957,N_14417,N_14409);
and U14958 (N_14958,N_14378,N_14247);
xnor U14959 (N_14959,N_14186,N_14086);
and U14960 (N_14960,N_14175,N_14208);
and U14961 (N_14961,N_14044,N_14073);
nand U14962 (N_14962,N_14303,N_14082);
or U14963 (N_14963,N_14194,N_14171);
nand U14964 (N_14964,N_14424,N_14498);
nand U14965 (N_14965,N_14046,N_14273);
nor U14966 (N_14966,N_14172,N_14215);
and U14967 (N_14967,N_14361,N_14481);
or U14968 (N_14968,N_14232,N_14299);
nor U14969 (N_14969,N_14065,N_14320);
nor U14970 (N_14970,N_14258,N_14334);
nand U14971 (N_14971,N_14060,N_14282);
nand U14972 (N_14972,N_14395,N_14342);
xnor U14973 (N_14973,N_14374,N_14075);
nand U14974 (N_14974,N_14027,N_14149);
nor U14975 (N_14975,N_14195,N_14364);
xnor U14976 (N_14976,N_14490,N_14011);
nor U14977 (N_14977,N_14078,N_14215);
or U14978 (N_14978,N_14132,N_14416);
nor U14979 (N_14979,N_14232,N_14081);
or U14980 (N_14980,N_14165,N_14051);
and U14981 (N_14981,N_14372,N_14219);
nor U14982 (N_14982,N_14362,N_14295);
and U14983 (N_14983,N_14420,N_14442);
or U14984 (N_14984,N_14150,N_14237);
or U14985 (N_14985,N_14472,N_14014);
and U14986 (N_14986,N_14451,N_14390);
nor U14987 (N_14987,N_14355,N_14130);
nor U14988 (N_14988,N_14074,N_14107);
nand U14989 (N_14989,N_14021,N_14199);
or U14990 (N_14990,N_14259,N_14280);
or U14991 (N_14991,N_14425,N_14476);
nand U14992 (N_14992,N_14296,N_14054);
and U14993 (N_14993,N_14165,N_14493);
and U14994 (N_14994,N_14075,N_14204);
and U14995 (N_14995,N_14451,N_14155);
or U14996 (N_14996,N_14141,N_14072);
and U14997 (N_14997,N_14222,N_14039);
nand U14998 (N_14998,N_14241,N_14030);
and U14999 (N_14999,N_14169,N_14459);
nor U15000 (N_15000,N_14825,N_14884);
or U15001 (N_15001,N_14534,N_14834);
nand U15002 (N_15002,N_14886,N_14805);
or U15003 (N_15003,N_14631,N_14836);
and U15004 (N_15004,N_14863,N_14906);
nor U15005 (N_15005,N_14852,N_14742);
nor U15006 (N_15006,N_14833,N_14804);
and U15007 (N_15007,N_14708,N_14745);
and U15008 (N_15008,N_14890,N_14902);
and U15009 (N_15009,N_14741,N_14983);
and U15010 (N_15010,N_14541,N_14577);
or U15011 (N_15011,N_14506,N_14756);
or U15012 (N_15012,N_14757,N_14823);
nor U15013 (N_15013,N_14963,N_14583);
and U15014 (N_15014,N_14647,N_14965);
and U15015 (N_15015,N_14682,N_14657);
or U15016 (N_15016,N_14513,N_14785);
and U15017 (N_15017,N_14849,N_14750);
nor U15018 (N_15018,N_14775,N_14851);
nor U15019 (N_15019,N_14616,N_14567);
and U15020 (N_15020,N_14699,N_14564);
xor U15021 (N_15021,N_14707,N_14956);
and U15022 (N_15022,N_14720,N_14744);
nand U15023 (N_15023,N_14686,N_14650);
nand U15024 (N_15024,N_14938,N_14710);
or U15025 (N_15025,N_14792,N_14967);
xor U15026 (N_15026,N_14698,N_14611);
xnor U15027 (N_15027,N_14999,N_14571);
or U15028 (N_15028,N_14931,N_14801);
and U15029 (N_15029,N_14576,N_14689);
nand U15030 (N_15030,N_14923,N_14934);
and U15031 (N_15031,N_14525,N_14982);
and U15032 (N_15032,N_14962,N_14843);
nand U15033 (N_15033,N_14865,N_14780);
and U15034 (N_15034,N_14986,N_14837);
and U15035 (N_15035,N_14762,N_14717);
nand U15036 (N_15036,N_14688,N_14747);
nand U15037 (N_15037,N_14526,N_14626);
nand U15038 (N_15038,N_14937,N_14746);
or U15039 (N_15039,N_14822,N_14661);
or U15040 (N_15040,N_14530,N_14909);
and U15041 (N_15041,N_14977,N_14721);
nand U15042 (N_15042,N_14867,N_14592);
nand U15043 (N_15043,N_14531,N_14594);
or U15044 (N_15044,N_14992,N_14892);
nor U15045 (N_15045,N_14544,N_14677);
nor U15046 (N_15046,N_14572,N_14552);
or U15047 (N_15047,N_14697,N_14954);
or U15048 (N_15048,N_14998,N_14809);
nor U15049 (N_15049,N_14927,N_14706);
xnor U15050 (N_15050,N_14591,N_14540);
nand U15051 (N_15051,N_14709,N_14895);
and U15052 (N_15052,N_14939,N_14789);
nand U15053 (N_15053,N_14889,N_14716);
nor U15054 (N_15054,N_14947,N_14946);
or U15055 (N_15055,N_14795,N_14960);
nor U15056 (N_15056,N_14735,N_14918);
or U15057 (N_15057,N_14640,N_14847);
nor U15058 (N_15058,N_14703,N_14700);
or U15059 (N_15059,N_14635,N_14722);
or U15060 (N_15060,N_14578,N_14502);
or U15061 (N_15061,N_14628,N_14959);
or U15062 (N_15062,N_14898,N_14582);
nor U15063 (N_15063,N_14752,N_14821);
and U15064 (N_15064,N_14539,N_14684);
and U15065 (N_15065,N_14812,N_14702);
nor U15066 (N_15066,N_14712,N_14538);
or U15067 (N_15067,N_14632,N_14987);
and U15068 (N_15068,N_14733,N_14951);
or U15069 (N_15069,N_14517,N_14556);
nor U15070 (N_15070,N_14925,N_14674);
or U15071 (N_15071,N_14669,N_14605);
or U15072 (N_15072,N_14738,N_14844);
xnor U15073 (N_15073,N_14759,N_14976);
nand U15074 (N_15074,N_14561,N_14731);
nor U15075 (N_15075,N_14602,N_14520);
nand U15076 (N_15076,N_14830,N_14914);
nand U15077 (N_15077,N_14774,N_14511);
or U15078 (N_15078,N_14672,N_14880);
nand U15079 (N_15079,N_14915,N_14969);
or U15080 (N_15080,N_14877,N_14828);
or U15081 (N_15081,N_14818,N_14781);
or U15082 (N_15082,N_14943,N_14971);
xnor U15083 (N_15083,N_14770,N_14916);
nor U15084 (N_15084,N_14869,N_14569);
nor U15085 (N_15085,N_14715,N_14642);
nor U15086 (N_15086,N_14850,N_14595);
nand U15087 (N_15087,N_14814,N_14664);
nor U15088 (N_15088,N_14793,N_14961);
nand U15089 (N_15089,N_14866,N_14945);
and U15090 (N_15090,N_14760,N_14732);
or U15091 (N_15091,N_14878,N_14797);
xor U15092 (N_15092,N_14656,N_14958);
nand U15093 (N_15093,N_14819,N_14586);
nand U15094 (N_15094,N_14523,N_14758);
nand U15095 (N_15095,N_14769,N_14743);
nand U15096 (N_15096,N_14701,N_14548);
nand U15097 (N_15097,N_14779,N_14996);
nand U15098 (N_15098,N_14871,N_14860);
nor U15099 (N_15099,N_14997,N_14993);
or U15100 (N_15100,N_14719,N_14614);
nor U15101 (N_15101,N_14913,N_14554);
nand U15102 (N_15102,N_14748,N_14585);
or U15103 (N_15103,N_14547,N_14560);
or U15104 (N_15104,N_14562,N_14893);
and U15105 (N_15105,N_14680,N_14806);
nor U15106 (N_15106,N_14876,N_14619);
nand U15107 (N_15107,N_14655,N_14668);
xor U15108 (N_15108,N_14607,N_14535);
and U15109 (N_15109,N_14930,N_14786);
or U15110 (N_15110,N_14533,N_14767);
nor U15111 (N_15111,N_14832,N_14826);
nand U15112 (N_15112,N_14888,N_14675);
or U15113 (N_15113,N_14613,N_14791);
nor U15114 (N_15114,N_14555,N_14799);
xor U15115 (N_15115,N_14776,N_14885);
and U15116 (N_15116,N_14955,N_14581);
and U15117 (N_15117,N_14514,N_14524);
nand U15118 (N_15118,N_14693,N_14536);
or U15119 (N_15119,N_14929,N_14908);
and U15120 (N_15120,N_14597,N_14645);
nand U15121 (N_15121,N_14864,N_14891);
and U15122 (N_15122,N_14573,N_14740);
nor U15123 (N_15123,N_14667,N_14783);
and U15124 (N_15124,N_14978,N_14621);
nor U15125 (N_15125,N_14755,N_14813);
and U15126 (N_15126,N_14553,N_14512);
nor U15127 (N_15127,N_14550,N_14777);
nand U15128 (N_15128,N_14598,N_14790);
xor U15129 (N_15129,N_14824,N_14692);
and U15130 (N_15130,N_14610,N_14521);
nor U15131 (N_15131,N_14728,N_14500);
or U15132 (N_15132,N_14907,N_14985);
nor U15133 (N_15133,N_14690,N_14508);
and U15134 (N_15134,N_14537,N_14570);
nand U15135 (N_15135,N_14634,N_14827);
or U15136 (N_15136,N_14882,N_14545);
nand U15137 (N_15137,N_14988,N_14815);
xnor U15138 (N_15138,N_14899,N_14796);
and U15139 (N_15139,N_14788,N_14516);
or U15140 (N_15140,N_14798,N_14654);
xor U15141 (N_15141,N_14685,N_14639);
or U15142 (N_15142,N_14651,N_14942);
and U15143 (N_15143,N_14881,N_14920);
or U15144 (N_15144,N_14989,N_14665);
nor U15145 (N_15145,N_14768,N_14966);
xnor U15146 (N_15146,N_14563,N_14624);
nor U15147 (N_15147,N_14580,N_14638);
or U15148 (N_15148,N_14948,N_14940);
and U15149 (N_15149,N_14932,N_14858);
or U15150 (N_15150,N_14903,N_14979);
nor U15151 (N_15151,N_14944,N_14687);
nand U15152 (N_15152,N_14507,N_14896);
nand U15153 (N_15153,N_14924,N_14725);
and U15154 (N_15154,N_14991,N_14968);
nor U15155 (N_15155,N_14696,N_14663);
nor U15156 (N_15156,N_14608,N_14764);
nand U15157 (N_15157,N_14620,N_14649);
nand U15158 (N_15158,N_14846,N_14606);
or U15159 (N_15159,N_14970,N_14565);
xor U15160 (N_15160,N_14841,N_14644);
and U15161 (N_15161,N_14623,N_14739);
nor U15162 (N_15162,N_14933,N_14853);
nor U15163 (N_15163,N_14807,N_14673);
and U15164 (N_15164,N_14765,N_14551);
and U15165 (N_15165,N_14676,N_14808);
or U15166 (N_15166,N_14980,N_14782);
nand U15167 (N_15167,N_14839,N_14519);
nand U15168 (N_15168,N_14532,N_14981);
and U15169 (N_15169,N_14599,N_14528);
and U15170 (N_15170,N_14949,N_14928);
or U15171 (N_15171,N_14527,N_14615);
and U15172 (N_15172,N_14800,N_14994);
and U15173 (N_15173,N_14921,N_14727);
or U15174 (N_15174,N_14546,N_14953);
nor U15175 (N_15175,N_14670,N_14622);
nand U15176 (N_15176,N_14840,N_14711);
or U15177 (N_15177,N_14854,N_14603);
nand U15178 (N_15178,N_14671,N_14625);
nand U15179 (N_15179,N_14905,N_14566);
nor U15180 (N_15180,N_14618,N_14723);
nor U15181 (N_15181,N_14952,N_14629);
nor U15182 (N_15182,N_14568,N_14787);
nor U15183 (N_15183,N_14510,N_14505);
and U15184 (N_15184,N_14842,N_14848);
and U15185 (N_15185,N_14643,N_14816);
nand U15186 (N_15186,N_14653,N_14904);
and U15187 (N_15187,N_14666,N_14973);
or U15188 (N_15188,N_14529,N_14509);
and U15189 (N_15189,N_14811,N_14646);
nor U15190 (N_15190,N_14630,N_14990);
and U15191 (N_15191,N_14838,N_14964);
and U15192 (N_15192,N_14590,N_14935);
nand U15193 (N_15193,N_14941,N_14713);
nand U15194 (N_15194,N_14995,N_14660);
nor U15195 (N_15195,N_14974,N_14810);
nand U15196 (N_15196,N_14926,N_14835);
and U15197 (N_15197,N_14600,N_14784);
or U15198 (N_15198,N_14912,N_14831);
nor U15199 (N_15199,N_14636,N_14542);
xor U15200 (N_15200,N_14609,N_14515);
and U15201 (N_15201,N_14857,N_14856);
and U15202 (N_15202,N_14705,N_14936);
xnor U15203 (N_15203,N_14557,N_14771);
or U15204 (N_15204,N_14753,N_14773);
or U15205 (N_15205,N_14901,N_14975);
and U15206 (N_15206,N_14683,N_14589);
nand U15207 (N_15207,N_14872,N_14694);
and U15208 (N_15208,N_14575,N_14549);
nand U15209 (N_15209,N_14718,N_14627);
or U15210 (N_15210,N_14587,N_14503);
and U15211 (N_15211,N_14751,N_14726);
and U15212 (N_15212,N_14829,N_14845);
or U15213 (N_15213,N_14910,N_14820);
and U15214 (N_15214,N_14559,N_14802);
and U15215 (N_15215,N_14887,N_14724);
nand U15216 (N_15216,N_14919,N_14601);
nor U15217 (N_15217,N_14922,N_14859);
or U15218 (N_15218,N_14612,N_14543);
nand U15219 (N_15219,N_14957,N_14817);
nor U15220 (N_15220,N_14803,N_14862);
xor U15221 (N_15221,N_14778,N_14900);
xnor U15222 (N_15222,N_14681,N_14579);
and U15223 (N_15223,N_14855,N_14501);
nand U15224 (N_15224,N_14879,N_14734);
nor U15225 (N_15225,N_14950,N_14749);
and U15226 (N_15226,N_14704,N_14897);
and U15227 (N_15227,N_14870,N_14972);
nand U15228 (N_15228,N_14794,N_14695);
and U15229 (N_15229,N_14730,N_14641);
nand U15230 (N_15230,N_14861,N_14729);
nand U15231 (N_15231,N_14772,N_14558);
nor U15232 (N_15232,N_14504,N_14714);
nor U15233 (N_15233,N_14678,N_14875);
nor U15234 (N_15234,N_14679,N_14648);
xor U15235 (N_15235,N_14652,N_14662);
and U15236 (N_15236,N_14737,N_14868);
or U15237 (N_15237,N_14917,N_14518);
or U15238 (N_15238,N_14604,N_14873);
nand U15239 (N_15239,N_14894,N_14617);
and U15240 (N_15240,N_14984,N_14522);
nor U15241 (N_15241,N_14637,N_14596);
nor U15242 (N_15242,N_14911,N_14763);
and U15243 (N_15243,N_14574,N_14761);
or U15244 (N_15244,N_14659,N_14633);
nor U15245 (N_15245,N_14593,N_14658);
nor U15246 (N_15246,N_14874,N_14691);
nor U15247 (N_15247,N_14766,N_14584);
or U15248 (N_15248,N_14588,N_14736);
and U15249 (N_15249,N_14754,N_14883);
nor U15250 (N_15250,N_14650,N_14830);
or U15251 (N_15251,N_14691,N_14528);
and U15252 (N_15252,N_14548,N_14509);
nand U15253 (N_15253,N_14797,N_14890);
nand U15254 (N_15254,N_14790,N_14583);
and U15255 (N_15255,N_14984,N_14930);
or U15256 (N_15256,N_14747,N_14921);
nand U15257 (N_15257,N_14622,N_14961);
and U15258 (N_15258,N_14813,N_14551);
or U15259 (N_15259,N_14752,N_14861);
and U15260 (N_15260,N_14757,N_14523);
nand U15261 (N_15261,N_14558,N_14751);
and U15262 (N_15262,N_14723,N_14729);
nand U15263 (N_15263,N_14831,N_14875);
nand U15264 (N_15264,N_14861,N_14625);
or U15265 (N_15265,N_14590,N_14646);
nand U15266 (N_15266,N_14679,N_14887);
or U15267 (N_15267,N_14903,N_14847);
nand U15268 (N_15268,N_14753,N_14703);
nand U15269 (N_15269,N_14639,N_14511);
or U15270 (N_15270,N_14771,N_14834);
and U15271 (N_15271,N_14578,N_14662);
or U15272 (N_15272,N_14515,N_14871);
or U15273 (N_15273,N_14710,N_14813);
nand U15274 (N_15274,N_14560,N_14653);
and U15275 (N_15275,N_14994,N_14686);
or U15276 (N_15276,N_14921,N_14501);
nand U15277 (N_15277,N_14954,N_14511);
nand U15278 (N_15278,N_14985,N_14609);
nor U15279 (N_15279,N_14575,N_14939);
nor U15280 (N_15280,N_14965,N_14959);
and U15281 (N_15281,N_14575,N_14867);
nand U15282 (N_15282,N_14958,N_14562);
nand U15283 (N_15283,N_14615,N_14820);
and U15284 (N_15284,N_14774,N_14888);
and U15285 (N_15285,N_14865,N_14776);
nor U15286 (N_15286,N_14755,N_14947);
and U15287 (N_15287,N_14990,N_14585);
or U15288 (N_15288,N_14659,N_14740);
and U15289 (N_15289,N_14995,N_14585);
nor U15290 (N_15290,N_14552,N_14641);
nand U15291 (N_15291,N_14885,N_14854);
nor U15292 (N_15292,N_14830,N_14893);
nor U15293 (N_15293,N_14988,N_14950);
nor U15294 (N_15294,N_14755,N_14730);
xor U15295 (N_15295,N_14957,N_14663);
nand U15296 (N_15296,N_14878,N_14717);
nand U15297 (N_15297,N_14636,N_14730);
nand U15298 (N_15298,N_14955,N_14575);
nor U15299 (N_15299,N_14670,N_14792);
or U15300 (N_15300,N_14754,N_14662);
nand U15301 (N_15301,N_14848,N_14776);
xnor U15302 (N_15302,N_14839,N_14936);
and U15303 (N_15303,N_14989,N_14893);
or U15304 (N_15304,N_14900,N_14582);
nor U15305 (N_15305,N_14868,N_14808);
nand U15306 (N_15306,N_14801,N_14711);
or U15307 (N_15307,N_14841,N_14554);
and U15308 (N_15308,N_14992,N_14821);
nand U15309 (N_15309,N_14531,N_14693);
nand U15310 (N_15310,N_14816,N_14743);
nor U15311 (N_15311,N_14952,N_14910);
nand U15312 (N_15312,N_14643,N_14728);
xor U15313 (N_15313,N_14827,N_14746);
or U15314 (N_15314,N_14606,N_14849);
nor U15315 (N_15315,N_14718,N_14667);
and U15316 (N_15316,N_14645,N_14740);
xnor U15317 (N_15317,N_14557,N_14862);
and U15318 (N_15318,N_14590,N_14950);
and U15319 (N_15319,N_14717,N_14749);
nor U15320 (N_15320,N_14790,N_14863);
or U15321 (N_15321,N_14904,N_14654);
xor U15322 (N_15322,N_14531,N_14828);
xnor U15323 (N_15323,N_14529,N_14605);
nand U15324 (N_15324,N_14934,N_14615);
and U15325 (N_15325,N_14809,N_14567);
or U15326 (N_15326,N_14545,N_14747);
and U15327 (N_15327,N_14647,N_14832);
nor U15328 (N_15328,N_14653,N_14504);
nand U15329 (N_15329,N_14607,N_14609);
or U15330 (N_15330,N_14703,N_14934);
or U15331 (N_15331,N_14839,N_14909);
xnor U15332 (N_15332,N_14804,N_14837);
nand U15333 (N_15333,N_14515,N_14708);
and U15334 (N_15334,N_14799,N_14668);
nand U15335 (N_15335,N_14543,N_14941);
and U15336 (N_15336,N_14822,N_14525);
and U15337 (N_15337,N_14870,N_14601);
nand U15338 (N_15338,N_14735,N_14958);
nor U15339 (N_15339,N_14622,N_14565);
and U15340 (N_15340,N_14832,N_14858);
or U15341 (N_15341,N_14821,N_14596);
nor U15342 (N_15342,N_14911,N_14701);
or U15343 (N_15343,N_14769,N_14710);
xor U15344 (N_15344,N_14700,N_14551);
and U15345 (N_15345,N_14534,N_14901);
and U15346 (N_15346,N_14672,N_14741);
or U15347 (N_15347,N_14721,N_14895);
or U15348 (N_15348,N_14916,N_14822);
or U15349 (N_15349,N_14684,N_14829);
and U15350 (N_15350,N_14908,N_14569);
and U15351 (N_15351,N_14952,N_14732);
and U15352 (N_15352,N_14536,N_14519);
and U15353 (N_15353,N_14970,N_14748);
nor U15354 (N_15354,N_14967,N_14681);
or U15355 (N_15355,N_14972,N_14945);
nand U15356 (N_15356,N_14842,N_14517);
nor U15357 (N_15357,N_14726,N_14786);
nand U15358 (N_15358,N_14729,N_14883);
or U15359 (N_15359,N_14588,N_14901);
nand U15360 (N_15360,N_14770,N_14589);
or U15361 (N_15361,N_14997,N_14943);
and U15362 (N_15362,N_14524,N_14673);
and U15363 (N_15363,N_14910,N_14677);
nor U15364 (N_15364,N_14838,N_14938);
and U15365 (N_15365,N_14718,N_14932);
or U15366 (N_15366,N_14774,N_14768);
nand U15367 (N_15367,N_14853,N_14687);
and U15368 (N_15368,N_14698,N_14548);
xnor U15369 (N_15369,N_14696,N_14815);
or U15370 (N_15370,N_14511,N_14533);
xnor U15371 (N_15371,N_14536,N_14720);
nor U15372 (N_15372,N_14868,N_14520);
nand U15373 (N_15373,N_14517,N_14757);
nor U15374 (N_15374,N_14866,N_14711);
or U15375 (N_15375,N_14765,N_14590);
nand U15376 (N_15376,N_14586,N_14876);
xnor U15377 (N_15377,N_14896,N_14761);
or U15378 (N_15378,N_14658,N_14684);
and U15379 (N_15379,N_14569,N_14755);
xnor U15380 (N_15380,N_14673,N_14730);
nor U15381 (N_15381,N_14919,N_14925);
and U15382 (N_15382,N_14594,N_14583);
or U15383 (N_15383,N_14976,N_14538);
or U15384 (N_15384,N_14506,N_14707);
or U15385 (N_15385,N_14757,N_14736);
or U15386 (N_15386,N_14685,N_14823);
and U15387 (N_15387,N_14818,N_14714);
and U15388 (N_15388,N_14717,N_14784);
and U15389 (N_15389,N_14825,N_14845);
or U15390 (N_15390,N_14544,N_14755);
and U15391 (N_15391,N_14902,N_14788);
nor U15392 (N_15392,N_14788,N_14550);
nor U15393 (N_15393,N_14601,N_14544);
nor U15394 (N_15394,N_14935,N_14852);
nand U15395 (N_15395,N_14824,N_14711);
and U15396 (N_15396,N_14745,N_14955);
nand U15397 (N_15397,N_14678,N_14975);
or U15398 (N_15398,N_14643,N_14580);
and U15399 (N_15399,N_14856,N_14958);
nand U15400 (N_15400,N_14610,N_14538);
nor U15401 (N_15401,N_14775,N_14745);
nor U15402 (N_15402,N_14665,N_14808);
nor U15403 (N_15403,N_14620,N_14731);
or U15404 (N_15404,N_14785,N_14537);
or U15405 (N_15405,N_14703,N_14536);
xnor U15406 (N_15406,N_14887,N_14968);
nor U15407 (N_15407,N_14549,N_14972);
nor U15408 (N_15408,N_14941,N_14650);
xor U15409 (N_15409,N_14974,N_14513);
nor U15410 (N_15410,N_14757,N_14989);
nand U15411 (N_15411,N_14759,N_14733);
and U15412 (N_15412,N_14837,N_14665);
and U15413 (N_15413,N_14761,N_14814);
and U15414 (N_15414,N_14577,N_14945);
and U15415 (N_15415,N_14529,N_14921);
and U15416 (N_15416,N_14944,N_14765);
xnor U15417 (N_15417,N_14822,N_14639);
and U15418 (N_15418,N_14861,N_14772);
xnor U15419 (N_15419,N_14672,N_14685);
or U15420 (N_15420,N_14869,N_14963);
nor U15421 (N_15421,N_14686,N_14983);
nand U15422 (N_15422,N_14635,N_14805);
or U15423 (N_15423,N_14990,N_14999);
or U15424 (N_15424,N_14714,N_14525);
or U15425 (N_15425,N_14526,N_14671);
and U15426 (N_15426,N_14729,N_14761);
nor U15427 (N_15427,N_14758,N_14965);
nor U15428 (N_15428,N_14840,N_14597);
xnor U15429 (N_15429,N_14949,N_14790);
and U15430 (N_15430,N_14535,N_14814);
and U15431 (N_15431,N_14715,N_14509);
nand U15432 (N_15432,N_14570,N_14813);
nor U15433 (N_15433,N_14639,N_14807);
and U15434 (N_15434,N_14604,N_14818);
nor U15435 (N_15435,N_14914,N_14780);
and U15436 (N_15436,N_14658,N_14874);
xor U15437 (N_15437,N_14723,N_14706);
nand U15438 (N_15438,N_14807,N_14830);
xnor U15439 (N_15439,N_14614,N_14830);
and U15440 (N_15440,N_14601,N_14796);
nor U15441 (N_15441,N_14541,N_14908);
or U15442 (N_15442,N_14727,N_14636);
nand U15443 (N_15443,N_14878,N_14958);
nor U15444 (N_15444,N_14644,N_14605);
nor U15445 (N_15445,N_14855,N_14772);
and U15446 (N_15446,N_14524,N_14765);
or U15447 (N_15447,N_14512,N_14503);
or U15448 (N_15448,N_14802,N_14750);
or U15449 (N_15449,N_14866,N_14648);
and U15450 (N_15450,N_14819,N_14814);
or U15451 (N_15451,N_14852,N_14513);
nand U15452 (N_15452,N_14535,N_14893);
and U15453 (N_15453,N_14709,N_14670);
and U15454 (N_15454,N_14812,N_14752);
nand U15455 (N_15455,N_14680,N_14687);
nand U15456 (N_15456,N_14611,N_14936);
nand U15457 (N_15457,N_14646,N_14672);
and U15458 (N_15458,N_14739,N_14898);
and U15459 (N_15459,N_14977,N_14789);
and U15460 (N_15460,N_14791,N_14875);
and U15461 (N_15461,N_14869,N_14829);
nor U15462 (N_15462,N_14601,N_14619);
xor U15463 (N_15463,N_14602,N_14595);
nor U15464 (N_15464,N_14602,N_14646);
nor U15465 (N_15465,N_14891,N_14533);
and U15466 (N_15466,N_14951,N_14699);
and U15467 (N_15467,N_14967,N_14525);
nor U15468 (N_15468,N_14708,N_14936);
nor U15469 (N_15469,N_14750,N_14912);
nor U15470 (N_15470,N_14583,N_14755);
nor U15471 (N_15471,N_14945,N_14757);
nor U15472 (N_15472,N_14797,N_14515);
or U15473 (N_15473,N_14686,N_14526);
or U15474 (N_15474,N_14927,N_14660);
xnor U15475 (N_15475,N_14635,N_14644);
and U15476 (N_15476,N_14906,N_14789);
and U15477 (N_15477,N_14642,N_14893);
nand U15478 (N_15478,N_14787,N_14607);
nor U15479 (N_15479,N_14920,N_14892);
and U15480 (N_15480,N_14564,N_14962);
and U15481 (N_15481,N_14603,N_14866);
and U15482 (N_15482,N_14672,N_14632);
or U15483 (N_15483,N_14955,N_14513);
nand U15484 (N_15484,N_14726,N_14607);
nand U15485 (N_15485,N_14510,N_14646);
nor U15486 (N_15486,N_14879,N_14623);
nor U15487 (N_15487,N_14745,N_14985);
nor U15488 (N_15488,N_14694,N_14987);
xor U15489 (N_15489,N_14643,N_14558);
nand U15490 (N_15490,N_14922,N_14756);
nand U15491 (N_15491,N_14842,N_14859);
nor U15492 (N_15492,N_14709,N_14607);
and U15493 (N_15493,N_14501,N_14851);
nand U15494 (N_15494,N_14853,N_14822);
nand U15495 (N_15495,N_14689,N_14588);
nor U15496 (N_15496,N_14757,N_14919);
or U15497 (N_15497,N_14998,N_14836);
nor U15498 (N_15498,N_14586,N_14813);
nand U15499 (N_15499,N_14887,N_14923);
and U15500 (N_15500,N_15156,N_15258);
xor U15501 (N_15501,N_15346,N_15318);
xor U15502 (N_15502,N_15050,N_15160);
nand U15503 (N_15503,N_15499,N_15158);
nand U15504 (N_15504,N_15034,N_15333);
or U15505 (N_15505,N_15497,N_15039);
or U15506 (N_15506,N_15120,N_15060);
or U15507 (N_15507,N_15047,N_15125);
nor U15508 (N_15508,N_15307,N_15218);
or U15509 (N_15509,N_15486,N_15254);
nor U15510 (N_15510,N_15434,N_15214);
xnor U15511 (N_15511,N_15000,N_15054);
and U15512 (N_15512,N_15243,N_15113);
nand U15513 (N_15513,N_15281,N_15455);
xor U15514 (N_15514,N_15264,N_15429);
xnor U15515 (N_15515,N_15102,N_15454);
and U15516 (N_15516,N_15106,N_15206);
nor U15517 (N_15517,N_15380,N_15262);
nand U15518 (N_15518,N_15256,N_15246);
or U15519 (N_15519,N_15070,N_15362);
xor U15520 (N_15520,N_15456,N_15126);
xnor U15521 (N_15521,N_15231,N_15329);
and U15522 (N_15522,N_15079,N_15285);
nand U15523 (N_15523,N_15229,N_15235);
nand U15524 (N_15524,N_15013,N_15432);
and U15525 (N_15525,N_15419,N_15324);
or U15526 (N_15526,N_15348,N_15320);
or U15527 (N_15527,N_15134,N_15390);
nor U15528 (N_15528,N_15468,N_15321);
nor U15529 (N_15529,N_15452,N_15044);
nor U15530 (N_15530,N_15252,N_15027);
or U15531 (N_15531,N_15467,N_15238);
nor U15532 (N_15532,N_15233,N_15338);
and U15533 (N_15533,N_15301,N_15341);
nor U15534 (N_15534,N_15393,N_15061);
and U15535 (N_15535,N_15314,N_15023);
or U15536 (N_15536,N_15268,N_15353);
nor U15537 (N_15537,N_15477,N_15111);
nor U15538 (N_15538,N_15086,N_15121);
nor U15539 (N_15539,N_15005,N_15396);
or U15540 (N_15540,N_15330,N_15217);
nand U15541 (N_15541,N_15108,N_15479);
nand U15542 (N_15542,N_15397,N_15377);
nor U15543 (N_15543,N_15123,N_15076);
and U15544 (N_15544,N_15412,N_15382);
or U15545 (N_15545,N_15240,N_15310);
and U15546 (N_15546,N_15480,N_15280);
nor U15547 (N_15547,N_15007,N_15275);
nand U15548 (N_15548,N_15265,N_15430);
nor U15549 (N_15549,N_15234,N_15288);
nor U15550 (N_15550,N_15482,N_15300);
and U15551 (N_15551,N_15260,N_15124);
or U15552 (N_15552,N_15127,N_15093);
xor U15553 (N_15553,N_15334,N_15290);
and U15554 (N_15554,N_15196,N_15327);
nand U15555 (N_15555,N_15131,N_15368);
xnor U15556 (N_15556,N_15496,N_15478);
and U15557 (N_15557,N_15161,N_15495);
and U15558 (N_15558,N_15149,N_15431);
or U15559 (N_15559,N_15176,N_15182);
nor U15560 (N_15560,N_15446,N_15272);
nand U15561 (N_15561,N_15177,N_15267);
nand U15562 (N_15562,N_15014,N_15356);
nor U15563 (N_15563,N_15490,N_15114);
and U15564 (N_15564,N_15394,N_15222);
xnor U15565 (N_15565,N_15485,N_15022);
or U15566 (N_15566,N_15194,N_15277);
xnor U15567 (N_15567,N_15067,N_15101);
nand U15568 (N_15568,N_15112,N_15080);
and U15569 (N_15569,N_15019,N_15144);
nor U15570 (N_15570,N_15109,N_15425);
nor U15571 (N_15571,N_15472,N_15029);
and U15572 (N_15572,N_15147,N_15444);
nor U15573 (N_15573,N_15247,N_15219);
xor U15574 (N_15574,N_15033,N_15323);
nand U15575 (N_15575,N_15098,N_15091);
nor U15576 (N_15576,N_15357,N_15132);
and U15577 (N_15577,N_15361,N_15152);
nor U15578 (N_15578,N_15313,N_15483);
nor U15579 (N_15579,N_15458,N_15021);
nor U15580 (N_15580,N_15332,N_15189);
nor U15581 (N_15581,N_15339,N_15306);
and U15582 (N_15582,N_15122,N_15053);
or U15583 (N_15583,N_15178,N_15286);
and U15584 (N_15584,N_15413,N_15175);
nor U15585 (N_15585,N_15433,N_15193);
nand U15586 (N_15586,N_15025,N_15066);
nor U15587 (N_15587,N_15028,N_15464);
and U15588 (N_15588,N_15374,N_15210);
or U15589 (N_15589,N_15351,N_15099);
and U15590 (N_15590,N_15088,N_15403);
and U15591 (N_15591,N_15269,N_15349);
nor U15592 (N_15592,N_15107,N_15011);
nand U15593 (N_15593,N_15045,N_15442);
or U15594 (N_15594,N_15230,N_15414);
nor U15595 (N_15595,N_15354,N_15459);
or U15596 (N_15596,N_15298,N_15063);
and U15597 (N_15597,N_15369,N_15470);
and U15598 (N_15598,N_15450,N_15475);
nand U15599 (N_15599,N_15089,N_15018);
nand U15600 (N_15600,N_15046,N_15469);
and U15601 (N_15601,N_15056,N_15097);
nand U15602 (N_15602,N_15360,N_15407);
or U15603 (N_15603,N_15409,N_15305);
or U15604 (N_15604,N_15365,N_15366);
nand U15605 (N_15605,N_15462,N_15140);
nor U15606 (N_15606,N_15418,N_15162);
xnor U15607 (N_15607,N_15115,N_15183);
nor U15608 (N_15608,N_15103,N_15166);
xnor U15609 (N_15609,N_15116,N_15359);
and U15610 (N_15610,N_15012,N_15040);
xnor U15611 (N_15611,N_15104,N_15173);
or U15612 (N_15612,N_15257,N_15031);
nor U15613 (N_15613,N_15187,N_15170);
nor U15614 (N_15614,N_15026,N_15424);
nor U15615 (N_15615,N_15169,N_15071);
xnor U15616 (N_15616,N_15457,N_15085);
nor U15617 (N_15617,N_15410,N_15335);
nor U15618 (N_15618,N_15367,N_15049);
nor U15619 (N_15619,N_15081,N_15282);
xnor U15620 (N_15620,N_15428,N_15068);
xor U15621 (N_15621,N_15375,N_15271);
nor U15622 (N_15622,N_15498,N_15465);
and U15623 (N_15623,N_15245,N_15100);
or U15624 (N_15624,N_15344,N_15095);
or U15625 (N_15625,N_15092,N_15074);
nand U15626 (N_15626,N_15289,N_15036);
nor U15627 (N_15627,N_15073,N_15266);
nand U15628 (N_15628,N_15057,N_15082);
nor U15629 (N_15629,N_15436,N_15242);
nor U15630 (N_15630,N_15003,N_15388);
xnor U15631 (N_15631,N_15437,N_15315);
or U15632 (N_15632,N_15276,N_15476);
or U15633 (N_15633,N_15096,N_15150);
nand U15634 (N_15634,N_15180,N_15278);
and U15635 (N_15635,N_15408,N_15017);
or U15636 (N_15636,N_15420,N_15445);
and U15637 (N_15637,N_15448,N_15188);
nand U15638 (N_15638,N_15133,N_15328);
nand U15639 (N_15639,N_15211,N_15062);
or U15640 (N_15640,N_15340,N_15201);
and U15641 (N_15641,N_15453,N_15355);
nand U15642 (N_15642,N_15386,N_15051);
and U15643 (N_15643,N_15337,N_15299);
nor U15644 (N_15644,N_15364,N_15325);
nand U15645 (N_15645,N_15208,N_15236);
and U15646 (N_15646,N_15192,N_15378);
nor U15647 (N_15647,N_15226,N_15438);
or U15648 (N_15648,N_15139,N_15241);
nand U15649 (N_15649,N_15381,N_15009);
and U15650 (N_15650,N_15371,N_15004);
xnor U15651 (N_15651,N_15212,N_15261);
and U15652 (N_15652,N_15002,N_15006);
nand U15653 (N_15653,N_15153,N_15148);
and U15654 (N_15654,N_15016,N_15042);
and U15655 (N_15655,N_15461,N_15165);
nand U15656 (N_15656,N_15358,N_15151);
or U15657 (N_15657,N_15020,N_15417);
and U15658 (N_15658,N_15200,N_15317);
xnor U15659 (N_15659,N_15379,N_15041);
and U15660 (N_15660,N_15185,N_15426);
nand U15661 (N_15661,N_15251,N_15345);
nor U15662 (N_15662,N_15473,N_15220);
xnor U15663 (N_15663,N_15263,N_15154);
nor U15664 (N_15664,N_15075,N_15392);
xor U15665 (N_15665,N_15015,N_15399);
nand U15666 (N_15666,N_15032,N_15402);
or U15667 (N_15667,N_15273,N_15312);
nor U15668 (N_15668,N_15463,N_15146);
or U15669 (N_15669,N_15294,N_15443);
or U15670 (N_15670,N_15347,N_15350);
nand U15671 (N_15671,N_15010,N_15376);
nand U15672 (N_15672,N_15205,N_15069);
or U15673 (N_15673,N_15048,N_15471);
or U15674 (N_15674,N_15308,N_15164);
or U15675 (N_15675,N_15439,N_15441);
nand U15676 (N_15676,N_15481,N_15171);
nand U15677 (N_15677,N_15387,N_15415);
nor U15678 (N_15678,N_15225,N_15253);
nor U15679 (N_15679,N_15336,N_15128);
nand U15680 (N_15680,N_15370,N_15215);
nor U15681 (N_15681,N_15174,N_15072);
nor U15682 (N_15682,N_15287,N_15058);
or U15683 (N_15683,N_15302,N_15037);
nand U15684 (N_15684,N_15400,N_15406);
nor U15685 (N_15685,N_15138,N_15384);
and U15686 (N_15686,N_15141,N_15190);
and U15687 (N_15687,N_15391,N_15249);
nand U15688 (N_15688,N_15385,N_15143);
nor U15689 (N_15689,N_15155,N_15421);
xnor U15690 (N_15690,N_15447,N_15159);
or U15691 (N_15691,N_15135,N_15322);
nand U15692 (N_15692,N_15064,N_15239);
and U15693 (N_15693,N_15492,N_15389);
xor U15694 (N_15694,N_15207,N_15493);
nor U15695 (N_15695,N_15343,N_15449);
or U15696 (N_15696,N_15279,N_15422);
nand U15697 (N_15697,N_15297,N_15184);
nand U15698 (N_15698,N_15181,N_15484);
and U15699 (N_15699,N_15427,N_15038);
nor U15700 (N_15700,N_15259,N_15270);
nor U15701 (N_15701,N_15198,N_15030);
xor U15702 (N_15702,N_15232,N_15224);
nand U15703 (N_15703,N_15199,N_15489);
nand U15704 (N_15704,N_15404,N_15311);
and U15705 (N_15705,N_15398,N_15157);
nand U15706 (N_15706,N_15203,N_15078);
and U15707 (N_15707,N_15395,N_15474);
nor U15708 (N_15708,N_15435,N_15087);
nor U15709 (N_15709,N_15142,N_15137);
nand U15710 (N_15710,N_15411,N_15179);
nor U15711 (N_15711,N_15244,N_15237);
nand U15712 (N_15712,N_15204,N_15216);
and U15713 (N_15713,N_15292,N_15283);
nor U15714 (N_15714,N_15105,N_15372);
nand U15715 (N_15715,N_15460,N_15284);
nand U15716 (N_15716,N_15309,N_15001);
or U15717 (N_15717,N_15221,N_15363);
or U15718 (N_15718,N_15250,N_15090);
nor U15719 (N_15719,N_15065,N_15043);
nor U15720 (N_15720,N_15405,N_15255);
and U15721 (N_15721,N_15024,N_15167);
or U15722 (N_15722,N_15191,N_15423);
or U15723 (N_15723,N_15291,N_15296);
xor U15724 (N_15724,N_15195,N_15401);
nor U15725 (N_15725,N_15487,N_15035);
or U15726 (N_15726,N_15440,N_15118);
nor U15727 (N_15727,N_15202,N_15186);
nand U15728 (N_15728,N_15293,N_15168);
and U15729 (N_15729,N_15352,N_15117);
nor U15730 (N_15730,N_15094,N_15055);
nand U15731 (N_15731,N_15209,N_15008);
and U15732 (N_15732,N_15052,N_15228);
nand U15733 (N_15733,N_15373,N_15119);
nor U15734 (N_15734,N_15145,N_15227);
nand U15735 (N_15735,N_15466,N_15331);
xor U15736 (N_15736,N_15248,N_15342);
and U15737 (N_15737,N_15059,N_15223);
or U15738 (N_15738,N_15077,N_15084);
and U15739 (N_15739,N_15491,N_15163);
nor U15740 (N_15740,N_15494,N_15136);
and U15741 (N_15741,N_15295,N_15488);
and U15742 (N_15742,N_15316,N_15304);
and U15743 (N_15743,N_15110,N_15303);
and U15744 (N_15744,N_15319,N_15213);
and U15745 (N_15745,N_15197,N_15383);
nor U15746 (N_15746,N_15083,N_15416);
or U15747 (N_15747,N_15172,N_15130);
nor U15748 (N_15748,N_15451,N_15326);
and U15749 (N_15749,N_15274,N_15129);
and U15750 (N_15750,N_15163,N_15122);
xor U15751 (N_15751,N_15277,N_15363);
or U15752 (N_15752,N_15475,N_15327);
and U15753 (N_15753,N_15286,N_15397);
and U15754 (N_15754,N_15362,N_15065);
xor U15755 (N_15755,N_15043,N_15338);
and U15756 (N_15756,N_15007,N_15095);
or U15757 (N_15757,N_15479,N_15038);
nor U15758 (N_15758,N_15180,N_15173);
and U15759 (N_15759,N_15216,N_15255);
or U15760 (N_15760,N_15266,N_15358);
and U15761 (N_15761,N_15192,N_15340);
and U15762 (N_15762,N_15006,N_15409);
or U15763 (N_15763,N_15174,N_15449);
nand U15764 (N_15764,N_15080,N_15122);
or U15765 (N_15765,N_15220,N_15157);
nand U15766 (N_15766,N_15145,N_15273);
and U15767 (N_15767,N_15353,N_15101);
nor U15768 (N_15768,N_15008,N_15065);
and U15769 (N_15769,N_15155,N_15196);
and U15770 (N_15770,N_15159,N_15227);
nand U15771 (N_15771,N_15421,N_15225);
nor U15772 (N_15772,N_15069,N_15230);
and U15773 (N_15773,N_15255,N_15490);
or U15774 (N_15774,N_15105,N_15419);
and U15775 (N_15775,N_15329,N_15406);
xnor U15776 (N_15776,N_15117,N_15215);
and U15777 (N_15777,N_15082,N_15251);
nor U15778 (N_15778,N_15081,N_15169);
xnor U15779 (N_15779,N_15432,N_15113);
nor U15780 (N_15780,N_15329,N_15367);
nor U15781 (N_15781,N_15105,N_15029);
nor U15782 (N_15782,N_15021,N_15120);
nand U15783 (N_15783,N_15231,N_15085);
nor U15784 (N_15784,N_15122,N_15050);
nor U15785 (N_15785,N_15231,N_15350);
nand U15786 (N_15786,N_15235,N_15494);
and U15787 (N_15787,N_15213,N_15108);
nand U15788 (N_15788,N_15061,N_15260);
or U15789 (N_15789,N_15001,N_15098);
nand U15790 (N_15790,N_15437,N_15068);
nor U15791 (N_15791,N_15103,N_15317);
nand U15792 (N_15792,N_15403,N_15437);
xnor U15793 (N_15793,N_15480,N_15380);
nor U15794 (N_15794,N_15476,N_15410);
nand U15795 (N_15795,N_15381,N_15193);
or U15796 (N_15796,N_15210,N_15490);
xor U15797 (N_15797,N_15017,N_15242);
nand U15798 (N_15798,N_15228,N_15413);
nand U15799 (N_15799,N_15199,N_15289);
nor U15800 (N_15800,N_15003,N_15290);
nand U15801 (N_15801,N_15485,N_15430);
or U15802 (N_15802,N_15201,N_15040);
and U15803 (N_15803,N_15350,N_15474);
nand U15804 (N_15804,N_15228,N_15093);
nand U15805 (N_15805,N_15483,N_15162);
or U15806 (N_15806,N_15210,N_15168);
nand U15807 (N_15807,N_15291,N_15173);
nand U15808 (N_15808,N_15037,N_15183);
or U15809 (N_15809,N_15373,N_15251);
and U15810 (N_15810,N_15273,N_15442);
and U15811 (N_15811,N_15173,N_15396);
nor U15812 (N_15812,N_15022,N_15493);
and U15813 (N_15813,N_15278,N_15435);
and U15814 (N_15814,N_15151,N_15319);
nand U15815 (N_15815,N_15462,N_15005);
or U15816 (N_15816,N_15446,N_15081);
xor U15817 (N_15817,N_15157,N_15294);
nand U15818 (N_15818,N_15146,N_15061);
or U15819 (N_15819,N_15491,N_15252);
and U15820 (N_15820,N_15337,N_15220);
and U15821 (N_15821,N_15430,N_15036);
and U15822 (N_15822,N_15021,N_15129);
nand U15823 (N_15823,N_15350,N_15084);
and U15824 (N_15824,N_15450,N_15061);
or U15825 (N_15825,N_15178,N_15102);
nand U15826 (N_15826,N_15406,N_15316);
or U15827 (N_15827,N_15312,N_15191);
nor U15828 (N_15828,N_15396,N_15307);
nand U15829 (N_15829,N_15360,N_15196);
nand U15830 (N_15830,N_15093,N_15383);
nand U15831 (N_15831,N_15199,N_15350);
nand U15832 (N_15832,N_15355,N_15106);
or U15833 (N_15833,N_15446,N_15133);
or U15834 (N_15834,N_15061,N_15220);
and U15835 (N_15835,N_15321,N_15259);
nor U15836 (N_15836,N_15302,N_15379);
nor U15837 (N_15837,N_15060,N_15239);
or U15838 (N_15838,N_15416,N_15040);
nand U15839 (N_15839,N_15174,N_15048);
nor U15840 (N_15840,N_15460,N_15140);
nor U15841 (N_15841,N_15394,N_15161);
xnor U15842 (N_15842,N_15096,N_15178);
or U15843 (N_15843,N_15028,N_15460);
and U15844 (N_15844,N_15167,N_15225);
nor U15845 (N_15845,N_15256,N_15156);
nand U15846 (N_15846,N_15170,N_15404);
nor U15847 (N_15847,N_15032,N_15298);
or U15848 (N_15848,N_15414,N_15199);
nor U15849 (N_15849,N_15210,N_15482);
nor U15850 (N_15850,N_15269,N_15454);
and U15851 (N_15851,N_15339,N_15225);
or U15852 (N_15852,N_15222,N_15248);
xnor U15853 (N_15853,N_15443,N_15060);
xor U15854 (N_15854,N_15358,N_15064);
or U15855 (N_15855,N_15226,N_15274);
or U15856 (N_15856,N_15209,N_15271);
or U15857 (N_15857,N_15499,N_15190);
nor U15858 (N_15858,N_15401,N_15182);
nor U15859 (N_15859,N_15282,N_15326);
nor U15860 (N_15860,N_15090,N_15195);
or U15861 (N_15861,N_15369,N_15311);
nand U15862 (N_15862,N_15069,N_15070);
xor U15863 (N_15863,N_15190,N_15135);
nand U15864 (N_15864,N_15056,N_15364);
or U15865 (N_15865,N_15154,N_15078);
or U15866 (N_15866,N_15381,N_15276);
or U15867 (N_15867,N_15330,N_15487);
nor U15868 (N_15868,N_15153,N_15146);
nand U15869 (N_15869,N_15207,N_15099);
and U15870 (N_15870,N_15400,N_15338);
nand U15871 (N_15871,N_15052,N_15362);
nand U15872 (N_15872,N_15085,N_15270);
nor U15873 (N_15873,N_15060,N_15014);
and U15874 (N_15874,N_15398,N_15210);
nor U15875 (N_15875,N_15093,N_15447);
or U15876 (N_15876,N_15003,N_15487);
or U15877 (N_15877,N_15238,N_15212);
nor U15878 (N_15878,N_15462,N_15247);
nand U15879 (N_15879,N_15494,N_15077);
nor U15880 (N_15880,N_15106,N_15490);
or U15881 (N_15881,N_15443,N_15202);
xor U15882 (N_15882,N_15307,N_15234);
nand U15883 (N_15883,N_15235,N_15388);
or U15884 (N_15884,N_15328,N_15442);
or U15885 (N_15885,N_15307,N_15066);
and U15886 (N_15886,N_15499,N_15245);
nor U15887 (N_15887,N_15366,N_15460);
nor U15888 (N_15888,N_15451,N_15265);
or U15889 (N_15889,N_15273,N_15065);
nand U15890 (N_15890,N_15124,N_15355);
nand U15891 (N_15891,N_15234,N_15251);
and U15892 (N_15892,N_15179,N_15393);
nor U15893 (N_15893,N_15037,N_15147);
or U15894 (N_15894,N_15388,N_15127);
or U15895 (N_15895,N_15387,N_15071);
nor U15896 (N_15896,N_15035,N_15345);
and U15897 (N_15897,N_15274,N_15035);
and U15898 (N_15898,N_15463,N_15034);
and U15899 (N_15899,N_15402,N_15167);
and U15900 (N_15900,N_15164,N_15417);
nor U15901 (N_15901,N_15481,N_15267);
nor U15902 (N_15902,N_15493,N_15071);
nand U15903 (N_15903,N_15318,N_15194);
nor U15904 (N_15904,N_15088,N_15272);
nand U15905 (N_15905,N_15039,N_15224);
and U15906 (N_15906,N_15493,N_15295);
nor U15907 (N_15907,N_15144,N_15488);
xor U15908 (N_15908,N_15191,N_15157);
xnor U15909 (N_15909,N_15137,N_15068);
and U15910 (N_15910,N_15387,N_15437);
xnor U15911 (N_15911,N_15227,N_15108);
nor U15912 (N_15912,N_15178,N_15291);
and U15913 (N_15913,N_15222,N_15434);
xnor U15914 (N_15914,N_15055,N_15413);
nand U15915 (N_15915,N_15170,N_15139);
nand U15916 (N_15916,N_15313,N_15331);
and U15917 (N_15917,N_15312,N_15458);
and U15918 (N_15918,N_15419,N_15496);
nand U15919 (N_15919,N_15428,N_15153);
nor U15920 (N_15920,N_15159,N_15428);
xor U15921 (N_15921,N_15316,N_15220);
or U15922 (N_15922,N_15007,N_15386);
nor U15923 (N_15923,N_15056,N_15443);
nor U15924 (N_15924,N_15328,N_15224);
and U15925 (N_15925,N_15236,N_15357);
and U15926 (N_15926,N_15477,N_15317);
nor U15927 (N_15927,N_15315,N_15088);
nand U15928 (N_15928,N_15292,N_15157);
and U15929 (N_15929,N_15319,N_15111);
nand U15930 (N_15930,N_15256,N_15106);
nand U15931 (N_15931,N_15107,N_15308);
or U15932 (N_15932,N_15322,N_15323);
nand U15933 (N_15933,N_15399,N_15238);
xor U15934 (N_15934,N_15021,N_15376);
and U15935 (N_15935,N_15369,N_15235);
nor U15936 (N_15936,N_15006,N_15212);
nor U15937 (N_15937,N_15208,N_15428);
nor U15938 (N_15938,N_15439,N_15213);
nand U15939 (N_15939,N_15090,N_15283);
or U15940 (N_15940,N_15226,N_15055);
nor U15941 (N_15941,N_15436,N_15455);
or U15942 (N_15942,N_15280,N_15292);
or U15943 (N_15943,N_15183,N_15432);
and U15944 (N_15944,N_15334,N_15218);
or U15945 (N_15945,N_15277,N_15023);
or U15946 (N_15946,N_15332,N_15109);
or U15947 (N_15947,N_15381,N_15188);
and U15948 (N_15948,N_15304,N_15444);
nand U15949 (N_15949,N_15182,N_15418);
and U15950 (N_15950,N_15471,N_15029);
xor U15951 (N_15951,N_15465,N_15075);
and U15952 (N_15952,N_15261,N_15301);
nor U15953 (N_15953,N_15184,N_15391);
nor U15954 (N_15954,N_15184,N_15449);
and U15955 (N_15955,N_15471,N_15380);
nand U15956 (N_15956,N_15093,N_15368);
nand U15957 (N_15957,N_15157,N_15267);
xor U15958 (N_15958,N_15018,N_15275);
or U15959 (N_15959,N_15028,N_15440);
or U15960 (N_15960,N_15336,N_15491);
or U15961 (N_15961,N_15325,N_15425);
and U15962 (N_15962,N_15090,N_15381);
nand U15963 (N_15963,N_15225,N_15462);
nand U15964 (N_15964,N_15498,N_15343);
or U15965 (N_15965,N_15292,N_15492);
and U15966 (N_15966,N_15351,N_15172);
or U15967 (N_15967,N_15233,N_15450);
nand U15968 (N_15968,N_15209,N_15351);
and U15969 (N_15969,N_15362,N_15421);
and U15970 (N_15970,N_15074,N_15004);
nor U15971 (N_15971,N_15001,N_15352);
nand U15972 (N_15972,N_15169,N_15306);
nand U15973 (N_15973,N_15343,N_15349);
nand U15974 (N_15974,N_15050,N_15235);
nand U15975 (N_15975,N_15040,N_15149);
xor U15976 (N_15976,N_15130,N_15226);
nor U15977 (N_15977,N_15158,N_15263);
or U15978 (N_15978,N_15079,N_15130);
nor U15979 (N_15979,N_15376,N_15280);
xnor U15980 (N_15980,N_15044,N_15041);
nand U15981 (N_15981,N_15401,N_15439);
and U15982 (N_15982,N_15353,N_15371);
nand U15983 (N_15983,N_15317,N_15148);
and U15984 (N_15984,N_15232,N_15348);
nor U15985 (N_15985,N_15150,N_15233);
or U15986 (N_15986,N_15284,N_15494);
xor U15987 (N_15987,N_15496,N_15010);
and U15988 (N_15988,N_15128,N_15075);
and U15989 (N_15989,N_15095,N_15451);
and U15990 (N_15990,N_15375,N_15165);
nor U15991 (N_15991,N_15338,N_15120);
nand U15992 (N_15992,N_15358,N_15237);
nor U15993 (N_15993,N_15082,N_15277);
nand U15994 (N_15994,N_15462,N_15439);
or U15995 (N_15995,N_15139,N_15024);
and U15996 (N_15996,N_15286,N_15245);
or U15997 (N_15997,N_15160,N_15444);
and U15998 (N_15998,N_15213,N_15244);
and U15999 (N_15999,N_15167,N_15276);
or U16000 (N_16000,N_15738,N_15686);
xor U16001 (N_16001,N_15887,N_15943);
nand U16002 (N_16002,N_15962,N_15559);
and U16003 (N_16003,N_15818,N_15938);
or U16004 (N_16004,N_15946,N_15626);
and U16005 (N_16005,N_15699,N_15632);
and U16006 (N_16006,N_15757,N_15950);
xnor U16007 (N_16007,N_15500,N_15915);
and U16008 (N_16008,N_15691,N_15508);
and U16009 (N_16009,N_15720,N_15912);
nor U16010 (N_16010,N_15571,N_15675);
nor U16011 (N_16011,N_15978,N_15521);
or U16012 (N_16012,N_15671,N_15790);
nor U16013 (N_16013,N_15504,N_15722);
xnor U16014 (N_16014,N_15877,N_15983);
xor U16015 (N_16015,N_15808,N_15916);
xor U16016 (N_16016,N_15771,N_15548);
or U16017 (N_16017,N_15893,N_15835);
nor U16018 (N_16018,N_15721,N_15616);
xor U16019 (N_16019,N_15564,N_15824);
nor U16020 (N_16020,N_15768,N_15730);
nor U16021 (N_16021,N_15842,N_15804);
or U16022 (N_16022,N_15595,N_15970);
and U16023 (N_16023,N_15754,N_15641);
nor U16024 (N_16024,N_15655,N_15569);
and U16025 (N_16025,N_15656,N_15693);
or U16026 (N_16026,N_15827,N_15515);
or U16027 (N_16027,N_15690,N_15549);
nand U16028 (N_16028,N_15766,N_15605);
or U16029 (N_16029,N_15914,N_15942);
nor U16030 (N_16030,N_15904,N_15780);
or U16031 (N_16031,N_15960,N_15793);
or U16032 (N_16032,N_15949,N_15861);
nor U16033 (N_16033,N_15939,N_15741);
or U16034 (N_16034,N_15619,N_15697);
nor U16035 (N_16035,N_15849,N_15581);
xor U16036 (N_16036,N_15611,N_15695);
and U16037 (N_16037,N_15816,N_15707);
nor U16038 (N_16038,N_15834,N_15764);
nor U16039 (N_16039,N_15883,N_15734);
or U16040 (N_16040,N_15647,N_15640);
and U16041 (N_16041,N_15737,N_15685);
nor U16042 (N_16042,N_15592,N_15570);
and U16043 (N_16043,N_15567,N_15791);
nor U16044 (N_16044,N_15859,N_15891);
and U16045 (N_16045,N_15858,N_15651);
nor U16046 (N_16046,N_15589,N_15937);
nor U16047 (N_16047,N_15822,N_15782);
and U16048 (N_16048,N_15501,N_15882);
or U16049 (N_16049,N_15586,N_15870);
nand U16050 (N_16050,N_15817,N_15514);
nor U16051 (N_16051,N_15558,N_15667);
and U16052 (N_16052,N_15839,N_15905);
nand U16053 (N_16053,N_15907,N_15840);
nand U16054 (N_16054,N_15958,N_15717);
or U16055 (N_16055,N_15614,N_15853);
or U16056 (N_16056,N_15979,N_15832);
or U16057 (N_16057,N_15638,N_15761);
nand U16058 (N_16058,N_15813,N_15948);
and U16059 (N_16059,N_15980,N_15509);
nor U16060 (N_16060,N_15664,N_15635);
or U16061 (N_16061,N_15799,N_15694);
nor U16062 (N_16062,N_15702,N_15873);
nand U16063 (N_16063,N_15797,N_15518);
and U16064 (N_16064,N_15535,N_15682);
xnor U16065 (N_16065,N_15863,N_15523);
and U16066 (N_16066,N_15673,N_15829);
xor U16067 (N_16067,N_15544,N_15551);
and U16068 (N_16068,N_15617,N_15931);
xor U16069 (N_16069,N_15936,N_15923);
nor U16070 (N_16070,N_15975,N_15927);
nand U16071 (N_16071,N_15781,N_15713);
or U16072 (N_16072,N_15769,N_15926);
or U16073 (N_16073,N_15715,N_15801);
xnor U16074 (N_16074,N_15844,N_15888);
or U16075 (N_16075,N_15908,N_15643);
and U16076 (N_16076,N_15634,N_15653);
or U16077 (N_16077,N_15982,N_15850);
xnor U16078 (N_16078,N_15658,N_15623);
nand U16079 (N_16079,N_15546,N_15711);
nand U16080 (N_16080,N_15510,N_15831);
xor U16081 (N_16081,N_15562,N_15961);
and U16082 (N_16082,N_15716,N_15528);
and U16083 (N_16083,N_15944,N_15867);
or U16084 (N_16084,N_15925,N_15911);
and U16085 (N_16085,N_15973,N_15531);
and U16086 (N_16086,N_15543,N_15806);
xnor U16087 (N_16087,N_15692,N_15725);
nor U16088 (N_16088,N_15807,N_15775);
and U16089 (N_16089,N_15563,N_15770);
nor U16090 (N_16090,N_15630,N_15661);
and U16091 (N_16091,N_15533,N_15989);
or U16092 (N_16092,N_15802,N_15892);
nand U16093 (N_16093,N_15534,N_15852);
nor U16094 (N_16094,N_15609,N_15755);
nand U16095 (N_16095,N_15865,N_15935);
or U16096 (N_16096,N_15557,N_15519);
xnor U16097 (N_16097,N_15959,N_15587);
xnor U16098 (N_16098,N_15968,N_15541);
and U16099 (N_16099,N_15580,N_15718);
xor U16100 (N_16100,N_15669,N_15620);
nor U16101 (N_16101,N_15752,N_15662);
nand U16102 (N_16102,N_15884,N_15810);
or U16103 (N_16103,N_15930,N_15594);
nand U16104 (N_16104,N_15756,N_15659);
or U16105 (N_16105,N_15940,N_15506);
and U16106 (N_16106,N_15706,N_15670);
xor U16107 (N_16107,N_15728,N_15795);
nor U16108 (N_16108,N_15674,N_15712);
or U16109 (N_16109,N_15868,N_15608);
and U16110 (N_16110,N_15872,N_15555);
and U16111 (N_16111,N_15825,N_15999);
nor U16112 (N_16112,N_15837,N_15524);
xnor U16113 (N_16113,N_15800,N_15590);
and U16114 (N_16114,N_15921,N_15507);
nor U16115 (N_16115,N_15941,N_15650);
xor U16116 (N_16116,N_15599,N_15974);
nor U16117 (N_16117,N_15698,N_15540);
and U16118 (N_16118,N_15746,N_15607);
nand U16119 (N_16119,N_15988,N_15951);
and U16120 (N_16120,N_15993,N_15869);
or U16121 (N_16121,N_15815,N_15760);
or U16122 (N_16122,N_15814,N_15646);
nand U16123 (N_16123,N_15919,N_15918);
or U16124 (N_16124,N_15579,N_15753);
nand U16125 (N_16125,N_15991,N_15864);
or U16126 (N_16126,N_15628,N_15847);
or U16127 (N_16127,N_15613,N_15593);
xnor U16128 (N_16128,N_15857,N_15622);
nor U16129 (N_16129,N_15900,N_15909);
or U16130 (N_16130,N_15666,N_15615);
xnor U16131 (N_16131,N_15920,N_15585);
nand U16132 (N_16132,N_15879,N_15739);
nand U16133 (N_16133,N_15560,N_15701);
or U16134 (N_16134,N_15727,N_15917);
nor U16135 (N_16135,N_15588,N_15985);
and U16136 (N_16136,N_15751,N_15724);
xnor U16137 (N_16137,N_15871,N_15583);
nand U16138 (N_16138,N_15803,N_15582);
or U16139 (N_16139,N_15828,N_15966);
and U16140 (N_16140,N_15680,N_15553);
or U16141 (N_16141,N_15789,N_15836);
nor U16142 (N_16142,N_15536,N_15731);
or U16143 (N_16143,N_15986,N_15601);
and U16144 (N_16144,N_15749,N_15934);
nor U16145 (N_16145,N_15826,N_15841);
nor U16146 (N_16146,N_15606,N_15684);
nor U16147 (N_16147,N_15933,N_15894);
nor U16148 (N_16148,N_15575,N_15830);
nand U16149 (N_16149,N_15901,N_15977);
nor U16150 (N_16150,N_15851,N_15767);
nand U16151 (N_16151,N_15689,N_15876);
and U16152 (N_16152,N_15502,N_15805);
and U16153 (N_16153,N_15773,N_15729);
and U16154 (N_16154,N_15537,N_15895);
and U16155 (N_16155,N_15798,N_15704);
nor U16156 (N_16156,N_15644,N_15954);
or U16157 (N_16157,N_15783,N_15965);
and U16158 (N_16158,N_15505,N_15542);
and U16159 (N_16159,N_15838,N_15726);
nand U16160 (N_16160,N_15998,N_15866);
nor U16161 (N_16161,N_15763,N_15772);
or U16162 (N_16162,N_15636,N_15776);
nand U16163 (N_16163,N_15545,N_15723);
or U16164 (N_16164,N_15774,N_15945);
xor U16165 (N_16165,N_15792,N_15994);
nor U16166 (N_16166,N_15902,N_15648);
nand U16167 (N_16167,N_15743,N_15854);
nand U16168 (N_16168,N_15823,N_15565);
or U16169 (N_16169,N_15513,N_15637);
and U16170 (N_16170,N_15657,N_15703);
and U16171 (N_16171,N_15610,N_15631);
or U16172 (N_16172,N_15520,N_15748);
and U16173 (N_16173,N_15922,N_15878);
nor U16174 (N_16174,N_15602,N_15618);
xor U16175 (N_16175,N_15556,N_15969);
nor U16176 (N_16176,N_15976,N_15794);
nor U16177 (N_16177,N_15627,N_15784);
nand U16178 (N_16178,N_15947,N_15732);
or U16179 (N_16179,N_15512,N_15604);
or U16180 (N_16180,N_15603,N_15552);
and U16181 (N_16181,N_15995,N_15677);
nor U16182 (N_16182,N_15516,N_15688);
nand U16183 (N_16183,N_15987,N_15709);
nand U16184 (N_16184,N_15612,N_15788);
xnor U16185 (N_16185,N_15928,N_15621);
nor U16186 (N_16186,N_15668,N_15812);
or U16187 (N_16187,N_15696,N_15809);
nor U16188 (N_16188,N_15511,N_15576);
nand U16189 (N_16189,N_15932,N_15778);
and U16190 (N_16190,N_15719,N_15700);
nand U16191 (N_16191,N_15996,N_15957);
nand U16192 (N_16192,N_15672,N_15963);
xnor U16193 (N_16193,N_15745,N_15759);
nor U16194 (N_16194,N_15903,N_15899);
and U16195 (N_16195,N_15897,N_15896);
or U16196 (N_16196,N_15848,N_15972);
nand U16197 (N_16197,N_15910,N_15708);
or U16198 (N_16198,N_15811,N_15880);
or U16199 (N_16199,N_15913,N_15855);
nand U16200 (N_16200,N_15971,N_15568);
or U16201 (N_16201,N_15624,N_15529);
nand U16202 (N_16202,N_15652,N_15597);
and U16203 (N_16203,N_15779,N_15625);
xnor U16204 (N_16204,N_15875,N_15796);
nand U16205 (N_16205,N_15906,N_15683);
nand U16206 (N_16206,N_15860,N_15679);
xor U16207 (N_16207,N_15740,N_15598);
nand U16208 (N_16208,N_15629,N_15517);
or U16209 (N_16209,N_15956,N_15786);
or U16210 (N_16210,N_15736,N_15539);
nor U16211 (N_16211,N_15642,N_15964);
nand U16212 (N_16212,N_15710,N_15967);
and U16213 (N_16213,N_15561,N_15990);
nor U16214 (N_16214,N_15845,N_15687);
or U16215 (N_16215,N_15762,N_15554);
nand U16216 (N_16216,N_15578,N_15566);
and U16217 (N_16217,N_15885,N_15765);
or U16218 (N_16218,N_15981,N_15889);
xor U16219 (N_16219,N_15952,N_15735);
or U16220 (N_16220,N_15526,N_15633);
or U16221 (N_16221,N_15538,N_15660);
and U16222 (N_16222,N_15525,N_15785);
and U16223 (N_16223,N_15750,N_15890);
or U16224 (N_16224,N_15856,N_15862);
nor U16225 (N_16225,N_15992,N_15929);
xnor U16226 (N_16226,N_15547,N_15705);
or U16227 (N_16227,N_15503,N_15573);
nand U16228 (N_16228,N_15874,N_15819);
and U16229 (N_16229,N_15742,N_15596);
nand U16230 (N_16230,N_15886,N_15663);
nand U16231 (N_16231,N_15665,N_15649);
and U16232 (N_16232,N_15758,N_15676);
nor U16233 (N_16233,N_15955,N_15645);
or U16234 (N_16234,N_15843,N_15833);
nor U16235 (N_16235,N_15681,N_15898);
xor U16236 (N_16236,N_15881,N_15522);
or U16237 (N_16237,N_15747,N_15924);
nand U16238 (N_16238,N_15654,N_15572);
or U16239 (N_16239,N_15733,N_15532);
nand U16240 (N_16240,N_15821,N_15639);
nand U16241 (N_16241,N_15574,N_15584);
nand U16242 (N_16242,N_15550,N_15530);
and U16243 (N_16243,N_15846,N_15714);
nor U16244 (N_16244,N_15577,N_15777);
nand U16245 (N_16245,N_15953,N_15600);
nand U16246 (N_16246,N_15997,N_15527);
and U16247 (N_16247,N_15984,N_15744);
xnor U16248 (N_16248,N_15591,N_15678);
and U16249 (N_16249,N_15820,N_15787);
nand U16250 (N_16250,N_15545,N_15774);
nand U16251 (N_16251,N_15628,N_15780);
or U16252 (N_16252,N_15527,N_15755);
nor U16253 (N_16253,N_15945,N_15573);
or U16254 (N_16254,N_15976,N_15624);
xor U16255 (N_16255,N_15883,N_15827);
or U16256 (N_16256,N_15925,N_15901);
or U16257 (N_16257,N_15984,N_15794);
or U16258 (N_16258,N_15920,N_15706);
or U16259 (N_16259,N_15911,N_15860);
and U16260 (N_16260,N_15589,N_15552);
nor U16261 (N_16261,N_15725,N_15659);
and U16262 (N_16262,N_15783,N_15832);
or U16263 (N_16263,N_15916,N_15519);
xor U16264 (N_16264,N_15753,N_15741);
nor U16265 (N_16265,N_15585,N_15921);
xor U16266 (N_16266,N_15860,N_15942);
nand U16267 (N_16267,N_15781,N_15519);
nor U16268 (N_16268,N_15809,N_15670);
xnor U16269 (N_16269,N_15868,N_15889);
or U16270 (N_16270,N_15579,N_15899);
and U16271 (N_16271,N_15688,N_15864);
nor U16272 (N_16272,N_15865,N_15747);
nor U16273 (N_16273,N_15617,N_15592);
or U16274 (N_16274,N_15843,N_15896);
and U16275 (N_16275,N_15870,N_15691);
xnor U16276 (N_16276,N_15572,N_15722);
or U16277 (N_16277,N_15868,N_15569);
xnor U16278 (N_16278,N_15681,N_15795);
and U16279 (N_16279,N_15670,N_15508);
nand U16280 (N_16280,N_15950,N_15894);
nor U16281 (N_16281,N_15979,N_15790);
xor U16282 (N_16282,N_15584,N_15914);
or U16283 (N_16283,N_15825,N_15534);
or U16284 (N_16284,N_15547,N_15574);
or U16285 (N_16285,N_15877,N_15633);
and U16286 (N_16286,N_15845,N_15979);
and U16287 (N_16287,N_15508,N_15630);
nand U16288 (N_16288,N_15662,N_15524);
and U16289 (N_16289,N_15541,N_15911);
nor U16290 (N_16290,N_15935,N_15580);
and U16291 (N_16291,N_15804,N_15998);
xnor U16292 (N_16292,N_15959,N_15829);
nand U16293 (N_16293,N_15822,N_15841);
or U16294 (N_16294,N_15637,N_15530);
xor U16295 (N_16295,N_15854,N_15532);
xnor U16296 (N_16296,N_15869,N_15519);
nor U16297 (N_16297,N_15794,N_15803);
nor U16298 (N_16298,N_15965,N_15517);
nor U16299 (N_16299,N_15706,N_15604);
nor U16300 (N_16300,N_15530,N_15926);
nor U16301 (N_16301,N_15930,N_15620);
and U16302 (N_16302,N_15824,N_15991);
or U16303 (N_16303,N_15807,N_15929);
nor U16304 (N_16304,N_15899,N_15534);
nand U16305 (N_16305,N_15773,N_15562);
and U16306 (N_16306,N_15980,N_15922);
and U16307 (N_16307,N_15669,N_15709);
nor U16308 (N_16308,N_15557,N_15512);
and U16309 (N_16309,N_15615,N_15916);
or U16310 (N_16310,N_15790,N_15590);
xor U16311 (N_16311,N_15877,N_15645);
nand U16312 (N_16312,N_15604,N_15906);
and U16313 (N_16313,N_15564,N_15549);
nand U16314 (N_16314,N_15874,N_15831);
xor U16315 (N_16315,N_15657,N_15819);
xnor U16316 (N_16316,N_15510,N_15949);
xor U16317 (N_16317,N_15821,N_15853);
nor U16318 (N_16318,N_15605,N_15741);
or U16319 (N_16319,N_15757,N_15845);
or U16320 (N_16320,N_15742,N_15736);
xor U16321 (N_16321,N_15803,N_15713);
nand U16322 (N_16322,N_15784,N_15602);
and U16323 (N_16323,N_15830,N_15523);
nand U16324 (N_16324,N_15859,N_15934);
or U16325 (N_16325,N_15628,N_15957);
nor U16326 (N_16326,N_15582,N_15574);
nor U16327 (N_16327,N_15689,N_15559);
nand U16328 (N_16328,N_15626,N_15938);
nor U16329 (N_16329,N_15570,N_15916);
or U16330 (N_16330,N_15555,N_15785);
nand U16331 (N_16331,N_15675,N_15990);
xnor U16332 (N_16332,N_15917,N_15644);
and U16333 (N_16333,N_15935,N_15599);
or U16334 (N_16334,N_15544,N_15744);
xnor U16335 (N_16335,N_15684,N_15851);
and U16336 (N_16336,N_15531,N_15922);
nor U16337 (N_16337,N_15685,N_15829);
and U16338 (N_16338,N_15933,N_15771);
nor U16339 (N_16339,N_15779,N_15701);
nor U16340 (N_16340,N_15577,N_15861);
nand U16341 (N_16341,N_15524,N_15852);
nor U16342 (N_16342,N_15987,N_15781);
and U16343 (N_16343,N_15758,N_15544);
or U16344 (N_16344,N_15870,N_15575);
or U16345 (N_16345,N_15796,N_15903);
or U16346 (N_16346,N_15557,N_15773);
and U16347 (N_16347,N_15769,N_15750);
nor U16348 (N_16348,N_15854,N_15909);
nor U16349 (N_16349,N_15814,N_15593);
and U16350 (N_16350,N_15569,N_15937);
or U16351 (N_16351,N_15553,N_15806);
and U16352 (N_16352,N_15835,N_15762);
or U16353 (N_16353,N_15505,N_15810);
nand U16354 (N_16354,N_15664,N_15510);
nor U16355 (N_16355,N_15716,N_15606);
xor U16356 (N_16356,N_15967,N_15767);
nand U16357 (N_16357,N_15905,N_15862);
nor U16358 (N_16358,N_15740,N_15791);
nor U16359 (N_16359,N_15802,N_15806);
and U16360 (N_16360,N_15584,N_15649);
xnor U16361 (N_16361,N_15618,N_15613);
xnor U16362 (N_16362,N_15800,N_15988);
and U16363 (N_16363,N_15896,N_15944);
xnor U16364 (N_16364,N_15804,N_15774);
nand U16365 (N_16365,N_15650,N_15711);
nor U16366 (N_16366,N_15783,N_15637);
or U16367 (N_16367,N_15989,N_15560);
xor U16368 (N_16368,N_15681,N_15752);
nand U16369 (N_16369,N_15611,N_15832);
nand U16370 (N_16370,N_15947,N_15639);
and U16371 (N_16371,N_15670,N_15823);
and U16372 (N_16372,N_15895,N_15551);
and U16373 (N_16373,N_15591,N_15687);
nand U16374 (N_16374,N_15506,N_15921);
xor U16375 (N_16375,N_15689,N_15885);
or U16376 (N_16376,N_15692,N_15741);
or U16377 (N_16377,N_15613,N_15530);
and U16378 (N_16378,N_15614,N_15697);
or U16379 (N_16379,N_15756,N_15951);
or U16380 (N_16380,N_15996,N_15876);
or U16381 (N_16381,N_15951,N_15554);
and U16382 (N_16382,N_15986,N_15840);
nand U16383 (N_16383,N_15544,N_15742);
or U16384 (N_16384,N_15738,N_15897);
and U16385 (N_16385,N_15569,N_15612);
nand U16386 (N_16386,N_15781,N_15625);
or U16387 (N_16387,N_15612,N_15986);
nor U16388 (N_16388,N_15766,N_15964);
nor U16389 (N_16389,N_15894,N_15562);
or U16390 (N_16390,N_15846,N_15814);
and U16391 (N_16391,N_15650,N_15906);
and U16392 (N_16392,N_15818,N_15539);
and U16393 (N_16393,N_15523,N_15749);
nor U16394 (N_16394,N_15506,N_15676);
nor U16395 (N_16395,N_15833,N_15792);
and U16396 (N_16396,N_15639,N_15827);
nor U16397 (N_16397,N_15904,N_15821);
nor U16398 (N_16398,N_15998,N_15857);
nor U16399 (N_16399,N_15968,N_15911);
nand U16400 (N_16400,N_15553,N_15534);
nand U16401 (N_16401,N_15597,N_15831);
and U16402 (N_16402,N_15963,N_15598);
nor U16403 (N_16403,N_15812,N_15806);
nor U16404 (N_16404,N_15897,N_15916);
xor U16405 (N_16405,N_15588,N_15505);
or U16406 (N_16406,N_15611,N_15948);
or U16407 (N_16407,N_15651,N_15513);
nor U16408 (N_16408,N_15909,N_15801);
and U16409 (N_16409,N_15974,N_15539);
and U16410 (N_16410,N_15887,N_15683);
nand U16411 (N_16411,N_15735,N_15843);
nand U16412 (N_16412,N_15981,N_15999);
nor U16413 (N_16413,N_15884,N_15626);
nor U16414 (N_16414,N_15863,N_15583);
xnor U16415 (N_16415,N_15969,N_15518);
or U16416 (N_16416,N_15614,N_15711);
or U16417 (N_16417,N_15854,N_15956);
and U16418 (N_16418,N_15904,N_15903);
nand U16419 (N_16419,N_15992,N_15899);
and U16420 (N_16420,N_15734,N_15563);
nand U16421 (N_16421,N_15893,N_15569);
or U16422 (N_16422,N_15912,N_15584);
nor U16423 (N_16423,N_15765,N_15684);
nor U16424 (N_16424,N_15742,N_15941);
and U16425 (N_16425,N_15847,N_15743);
and U16426 (N_16426,N_15579,N_15726);
and U16427 (N_16427,N_15529,N_15940);
nand U16428 (N_16428,N_15591,N_15910);
nor U16429 (N_16429,N_15967,N_15680);
and U16430 (N_16430,N_15707,N_15584);
or U16431 (N_16431,N_15859,N_15615);
nand U16432 (N_16432,N_15619,N_15656);
nand U16433 (N_16433,N_15963,N_15952);
or U16434 (N_16434,N_15670,N_15924);
nor U16435 (N_16435,N_15758,N_15962);
and U16436 (N_16436,N_15567,N_15620);
nor U16437 (N_16437,N_15759,N_15929);
xor U16438 (N_16438,N_15895,N_15658);
nor U16439 (N_16439,N_15507,N_15817);
nand U16440 (N_16440,N_15853,N_15879);
or U16441 (N_16441,N_15595,N_15946);
and U16442 (N_16442,N_15514,N_15755);
nand U16443 (N_16443,N_15766,N_15516);
nand U16444 (N_16444,N_15809,N_15672);
and U16445 (N_16445,N_15898,N_15699);
or U16446 (N_16446,N_15788,N_15843);
and U16447 (N_16447,N_15676,N_15656);
nor U16448 (N_16448,N_15841,N_15584);
and U16449 (N_16449,N_15588,N_15627);
nand U16450 (N_16450,N_15765,N_15601);
nand U16451 (N_16451,N_15603,N_15852);
or U16452 (N_16452,N_15890,N_15522);
nand U16453 (N_16453,N_15847,N_15869);
nor U16454 (N_16454,N_15556,N_15941);
or U16455 (N_16455,N_15613,N_15938);
and U16456 (N_16456,N_15540,N_15896);
xor U16457 (N_16457,N_15762,N_15646);
and U16458 (N_16458,N_15743,N_15619);
or U16459 (N_16459,N_15990,N_15870);
nand U16460 (N_16460,N_15546,N_15513);
nand U16461 (N_16461,N_15550,N_15750);
or U16462 (N_16462,N_15961,N_15638);
xnor U16463 (N_16463,N_15656,N_15737);
nor U16464 (N_16464,N_15864,N_15555);
nand U16465 (N_16465,N_15620,N_15900);
nand U16466 (N_16466,N_15826,N_15600);
nor U16467 (N_16467,N_15899,N_15818);
or U16468 (N_16468,N_15966,N_15690);
nor U16469 (N_16469,N_15727,N_15994);
nor U16470 (N_16470,N_15885,N_15771);
nand U16471 (N_16471,N_15978,N_15667);
and U16472 (N_16472,N_15690,N_15621);
and U16473 (N_16473,N_15788,N_15595);
nand U16474 (N_16474,N_15698,N_15739);
xnor U16475 (N_16475,N_15761,N_15619);
xnor U16476 (N_16476,N_15869,N_15795);
nor U16477 (N_16477,N_15595,N_15949);
nand U16478 (N_16478,N_15673,N_15743);
and U16479 (N_16479,N_15759,N_15580);
and U16480 (N_16480,N_15648,N_15664);
or U16481 (N_16481,N_15728,N_15806);
nor U16482 (N_16482,N_15763,N_15895);
nor U16483 (N_16483,N_15964,N_15817);
nand U16484 (N_16484,N_15688,N_15889);
or U16485 (N_16485,N_15796,N_15739);
nor U16486 (N_16486,N_15853,N_15956);
and U16487 (N_16487,N_15561,N_15832);
nand U16488 (N_16488,N_15888,N_15952);
nand U16489 (N_16489,N_15936,N_15520);
nor U16490 (N_16490,N_15839,N_15726);
or U16491 (N_16491,N_15658,N_15858);
nand U16492 (N_16492,N_15650,N_15673);
nor U16493 (N_16493,N_15850,N_15523);
xnor U16494 (N_16494,N_15872,N_15698);
and U16495 (N_16495,N_15509,N_15916);
or U16496 (N_16496,N_15516,N_15760);
and U16497 (N_16497,N_15775,N_15505);
or U16498 (N_16498,N_15893,N_15639);
nor U16499 (N_16499,N_15514,N_15918);
and U16500 (N_16500,N_16483,N_16030);
and U16501 (N_16501,N_16400,N_16117);
or U16502 (N_16502,N_16396,N_16053);
or U16503 (N_16503,N_16011,N_16160);
nor U16504 (N_16504,N_16312,N_16110);
or U16505 (N_16505,N_16317,N_16135);
nand U16506 (N_16506,N_16029,N_16475);
or U16507 (N_16507,N_16498,N_16299);
and U16508 (N_16508,N_16349,N_16048);
xnor U16509 (N_16509,N_16468,N_16458);
nor U16510 (N_16510,N_16062,N_16066);
nor U16511 (N_16511,N_16284,N_16417);
and U16512 (N_16512,N_16374,N_16385);
nor U16513 (N_16513,N_16454,N_16460);
nand U16514 (N_16514,N_16031,N_16478);
nor U16515 (N_16515,N_16262,N_16094);
nand U16516 (N_16516,N_16184,N_16046);
nor U16517 (N_16517,N_16063,N_16112);
nand U16518 (N_16518,N_16001,N_16490);
and U16519 (N_16519,N_16091,N_16226);
nand U16520 (N_16520,N_16217,N_16166);
nor U16521 (N_16521,N_16336,N_16242);
nor U16522 (N_16522,N_16418,N_16288);
nand U16523 (N_16523,N_16099,N_16311);
nor U16524 (N_16524,N_16174,N_16384);
nor U16525 (N_16525,N_16252,N_16208);
and U16526 (N_16526,N_16370,N_16018);
and U16527 (N_16527,N_16100,N_16143);
xnor U16528 (N_16528,N_16183,N_16363);
nor U16529 (N_16529,N_16213,N_16111);
nor U16530 (N_16530,N_16175,N_16103);
nand U16531 (N_16531,N_16267,N_16399);
and U16532 (N_16532,N_16136,N_16380);
nor U16533 (N_16533,N_16218,N_16153);
nand U16534 (N_16534,N_16192,N_16293);
nand U16535 (N_16535,N_16102,N_16230);
nand U16536 (N_16536,N_16322,N_16301);
or U16537 (N_16537,N_16024,N_16243);
and U16538 (N_16538,N_16133,N_16354);
or U16539 (N_16539,N_16059,N_16321);
nand U16540 (N_16540,N_16274,N_16342);
or U16541 (N_16541,N_16225,N_16351);
or U16542 (N_16542,N_16435,N_16320);
nand U16543 (N_16543,N_16037,N_16403);
nand U16544 (N_16544,N_16087,N_16042);
and U16545 (N_16545,N_16106,N_16497);
nand U16546 (N_16546,N_16357,N_16224);
or U16547 (N_16547,N_16041,N_16255);
or U16548 (N_16548,N_16474,N_16127);
nand U16549 (N_16549,N_16448,N_16486);
or U16550 (N_16550,N_16028,N_16348);
or U16551 (N_16551,N_16236,N_16219);
or U16552 (N_16552,N_16008,N_16169);
and U16553 (N_16553,N_16281,N_16057);
and U16554 (N_16554,N_16114,N_16437);
nand U16555 (N_16555,N_16344,N_16051);
or U16556 (N_16556,N_16198,N_16365);
nand U16557 (N_16557,N_16379,N_16414);
nand U16558 (N_16558,N_16369,N_16356);
nand U16559 (N_16559,N_16350,N_16473);
nor U16560 (N_16560,N_16016,N_16035);
and U16561 (N_16561,N_16347,N_16026);
nand U16562 (N_16562,N_16221,N_16200);
and U16563 (N_16563,N_16196,N_16280);
nor U16564 (N_16564,N_16328,N_16047);
nor U16565 (N_16565,N_16461,N_16378);
nand U16566 (N_16566,N_16150,N_16056);
nor U16567 (N_16567,N_16038,N_16049);
or U16568 (N_16568,N_16382,N_16425);
and U16569 (N_16569,N_16043,N_16431);
or U16570 (N_16570,N_16164,N_16205);
and U16571 (N_16571,N_16426,N_16416);
and U16572 (N_16572,N_16391,N_16427);
and U16573 (N_16573,N_16346,N_16146);
or U16574 (N_16574,N_16089,N_16294);
xor U16575 (N_16575,N_16204,N_16247);
or U16576 (N_16576,N_16251,N_16273);
nand U16577 (N_16577,N_16455,N_16072);
nand U16578 (N_16578,N_16119,N_16450);
or U16579 (N_16579,N_16006,N_16238);
xnor U16580 (N_16580,N_16307,N_16383);
nand U16581 (N_16581,N_16231,N_16408);
nand U16582 (N_16582,N_16093,N_16387);
nor U16583 (N_16583,N_16290,N_16083);
nand U16584 (N_16584,N_16295,N_16085);
and U16585 (N_16585,N_16261,N_16485);
and U16586 (N_16586,N_16096,N_16401);
xor U16587 (N_16587,N_16285,N_16156);
or U16588 (N_16588,N_16256,N_16496);
and U16589 (N_16589,N_16292,N_16209);
or U16590 (N_16590,N_16179,N_16097);
nor U16591 (N_16591,N_16297,N_16118);
nor U16592 (N_16592,N_16173,N_16394);
nand U16593 (N_16593,N_16068,N_16439);
or U16594 (N_16594,N_16142,N_16191);
or U16595 (N_16595,N_16270,N_16181);
nand U16596 (N_16596,N_16442,N_16451);
and U16597 (N_16597,N_16386,N_16278);
nor U16598 (N_16598,N_16163,N_16220);
nand U16599 (N_16599,N_16013,N_16471);
nand U16600 (N_16600,N_16000,N_16177);
or U16601 (N_16601,N_16039,N_16254);
nor U16602 (N_16602,N_16334,N_16176);
or U16603 (N_16603,N_16266,N_16313);
or U16604 (N_16604,N_16206,N_16428);
or U16605 (N_16605,N_16076,N_16190);
nor U16606 (N_16606,N_16055,N_16152);
and U16607 (N_16607,N_16144,N_16429);
and U16608 (N_16608,N_16108,N_16086);
or U16609 (N_16609,N_16159,N_16275);
and U16610 (N_16610,N_16469,N_16263);
or U16611 (N_16611,N_16145,N_16484);
xnor U16612 (N_16612,N_16337,N_16376);
or U16613 (N_16613,N_16023,N_16073);
nor U16614 (N_16614,N_16240,N_16027);
and U16615 (N_16615,N_16185,N_16194);
and U16616 (N_16616,N_16116,N_16113);
or U16617 (N_16617,N_16412,N_16430);
nand U16618 (N_16618,N_16075,N_16132);
nand U16619 (N_16619,N_16147,N_16331);
nor U16620 (N_16620,N_16074,N_16463);
nor U16621 (N_16621,N_16010,N_16434);
nor U16622 (N_16622,N_16241,N_16232);
nand U16623 (N_16623,N_16367,N_16371);
or U16624 (N_16624,N_16419,N_16375);
xor U16625 (N_16625,N_16015,N_16092);
nand U16626 (N_16626,N_16345,N_16202);
and U16627 (N_16627,N_16021,N_16323);
nand U16628 (N_16628,N_16245,N_16197);
nor U16629 (N_16629,N_16361,N_16487);
and U16630 (N_16630,N_16148,N_16466);
and U16631 (N_16631,N_16082,N_16235);
nor U16632 (N_16632,N_16067,N_16137);
nor U16633 (N_16633,N_16012,N_16444);
or U16634 (N_16634,N_16276,N_16207);
xor U16635 (N_16635,N_16339,N_16158);
and U16636 (N_16636,N_16095,N_16129);
and U16637 (N_16637,N_16289,N_16482);
or U16638 (N_16638,N_16186,N_16327);
nor U16639 (N_16639,N_16223,N_16489);
or U16640 (N_16640,N_16338,N_16304);
and U16641 (N_16641,N_16377,N_16310);
nand U16642 (N_16642,N_16362,N_16433);
and U16643 (N_16643,N_16470,N_16101);
nor U16644 (N_16644,N_16324,N_16189);
xor U16645 (N_16645,N_16054,N_16341);
and U16646 (N_16646,N_16305,N_16171);
nand U16647 (N_16647,N_16115,N_16123);
nand U16648 (N_16648,N_16303,N_16343);
nand U16649 (N_16649,N_16413,N_16456);
xnor U16650 (N_16650,N_16269,N_16022);
nor U16651 (N_16651,N_16494,N_16332);
and U16652 (N_16652,N_16033,N_16260);
and U16653 (N_16653,N_16335,N_16286);
nor U16654 (N_16654,N_16277,N_16193);
and U16655 (N_16655,N_16003,N_16229);
xnor U16656 (N_16656,N_16239,N_16464);
or U16657 (N_16657,N_16228,N_16329);
nand U16658 (N_16658,N_16415,N_16488);
or U16659 (N_16659,N_16271,N_16034);
nand U16660 (N_16660,N_16014,N_16032);
nand U16661 (N_16661,N_16170,N_16180);
xor U16662 (N_16662,N_16476,N_16154);
nor U16663 (N_16663,N_16017,N_16222);
nand U16664 (N_16664,N_16420,N_16234);
and U16665 (N_16665,N_16090,N_16407);
or U16666 (N_16666,N_16314,N_16125);
or U16667 (N_16667,N_16199,N_16326);
nor U16668 (N_16668,N_16259,N_16452);
or U16669 (N_16669,N_16465,N_16104);
nor U16670 (N_16670,N_16019,N_16162);
or U16671 (N_16671,N_16172,N_16315);
or U16672 (N_16672,N_16402,N_16447);
nand U16673 (N_16673,N_16355,N_16257);
and U16674 (N_16674,N_16318,N_16495);
nand U16675 (N_16675,N_16203,N_16409);
or U16676 (N_16676,N_16364,N_16005);
nor U16677 (N_16677,N_16368,N_16155);
or U16678 (N_16678,N_16268,N_16025);
and U16679 (N_16679,N_16250,N_16080);
nor U16680 (N_16680,N_16330,N_16134);
nor U16681 (N_16681,N_16440,N_16359);
and U16682 (N_16682,N_16406,N_16107);
or U16683 (N_16683,N_16366,N_16388);
nand U16684 (N_16684,N_16065,N_16405);
or U16685 (N_16685,N_16467,N_16045);
or U16686 (N_16686,N_16353,N_16462);
nand U16687 (N_16687,N_16128,N_16390);
and U16688 (N_16688,N_16493,N_16404);
nand U16689 (N_16689,N_16161,N_16167);
and U16690 (N_16690,N_16201,N_16248);
or U16691 (N_16691,N_16122,N_16453);
nand U16692 (N_16692,N_16050,N_16410);
and U16693 (N_16693,N_16071,N_16139);
nand U16694 (N_16694,N_16004,N_16149);
or U16695 (N_16695,N_16393,N_16397);
nand U16696 (N_16696,N_16084,N_16061);
xnor U16697 (N_16697,N_16436,N_16079);
and U16698 (N_16698,N_16237,N_16105);
and U16699 (N_16699,N_16306,N_16088);
nand U16700 (N_16700,N_16216,N_16296);
or U16701 (N_16701,N_16264,N_16165);
xor U16702 (N_16702,N_16126,N_16441);
and U16703 (N_16703,N_16492,N_16178);
nor U16704 (N_16704,N_16060,N_16443);
or U16705 (N_16705,N_16121,N_16141);
and U16706 (N_16706,N_16233,N_16389);
and U16707 (N_16707,N_16044,N_16477);
and U16708 (N_16708,N_16195,N_16373);
and U16709 (N_16709,N_16077,N_16265);
or U16710 (N_16710,N_16352,N_16182);
and U16711 (N_16711,N_16282,N_16446);
nand U16712 (N_16712,N_16283,N_16308);
and U16713 (N_16713,N_16020,N_16372);
and U16714 (N_16714,N_16479,N_16432);
nand U16715 (N_16715,N_16438,N_16358);
nand U16716 (N_16716,N_16298,N_16210);
or U16717 (N_16717,N_16212,N_16246);
nor U16718 (N_16718,N_16272,N_16291);
nand U16719 (N_16719,N_16424,N_16411);
or U16720 (N_16720,N_16002,N_16491);
nand U16721 (N_16721,N_16215,N_16392);
and U16722 (N_16722,N_16052,N_16445);
or U16723 (N_16723,N_16459,N_16258);
nor U16724 (N_16724,N_16287,N_16421);
nand U16725 (N_16725,N_16381,N_16070);
or U16726 (N_16726,N_16151,N_16481);
nand U16727 (N_16727,N_16398,N_16138);
nand U16728 (N_16728,N_16227,N_16058);
or U16729 (N_16729,N_16098,N_16157);
nand U16730 (N_16730,N_16472,N_16064);
xnor U16731 (N_16731,N_16130,N_16325);
and U16732 (N_16732,N_16319,N_16187);
nor U16733 (N_16733,N_16253,N_16069);
or U16734 (N_16734,N_16120,N_16131);
or U16735 (N_16735,N_16211,N_16168);
nor U16736 (N_16736,N_16188,N_16140);
nand U16737 (N_16737,N_16395,N_16244);
or U16738 (N_16738,N_16109,N_16078);
nor U16739 (N_16739,N_16316,N_16302);
or U16740 (N_16740,N_16300,N_16009);
nand U16741 (N_16741,N_16499,N_16457);
nand U16742 (N_16742,N_16449,N_16214);
nor U16743 (N_16743,N_16124,N_16081);
nor U16744 (N_16744,N_16340,N_16480);
and U16745 (N_16745,N_16279,N_16423);
and U16746 (N_16746,N_16333,N_16036);
and U16747 (N_16747,N_16007,N_16249);
nor U16748 (N_16748,N_16040,N_16360);
xnor U16749 (N_16749,N_16422,N_16309);
and U16750 (N_16750,N_16488,N_16329);
xnor U16751 (N_16751,N_16027,N_16451);
and U16752 (N_16752,N_16018,N_16365);
nor U16753 (N_16753,N_16211,N_16398);
nand U16754 (N_16754,N_16487,N_16472);
or U16755 (N_16755,N_16215,N_16126);
nand U16756 (N_16756,N_16411,N_16155);
nor U16757 (N_16757,N_16176,N_16219);
and U16758 (N_16758,N_16315,N_16456);
nor U16759 (N_16759,N_16253,N_16035);
and U16760 (N_16760,N_16399,N_16322);
nor U16761 (N_16761,N_16492,N_16481);
nand U16762 (N_16762,N_16471,N_16496);
nor U16763 (N_16763,N_16176,N_16139);
or U16764 (N_16764,N_16120,N_16250);
nor U16765 (N_16765,N_16171,N_16023);
nor U16766 (N_16766,N_16251,N_16142);
xnor U16767 (N_16767,N_16134,N_16025);
and U16768 (N_16768,N_16193,N_16453);
nand U16769 (N_16769,N_16406,N_16039);
nand U16770 (N_16770,N_16112,N_16010);
xnor U16771 (N_16771,N_16179,N_16319);
or U16772 (N_16772,N_16000,N_16373);
xnor U16773 (N_16773,N_16226,N_16243);
or U16774 (N_16774,N_16092,N_16115);
nand U16775 (N_16775,N_16333,N_16062);
nand U16776 (N_16776,N_16389,N_16460);
nand U16777 (N_16777,N_16160,N_16239);
and U16778 (N_16778,N_16174,N_16220);
xnor U16779 (N_16779,N_16080,N_16469);
and U16780 (N_16780,N_16334,N_16359);
nand U16781 (N_16781,N_16289,N_16399);
nand U16782 (N_16782,N_16253,N_16335);
nor U16783 (N_16783,N_16116,N_16299);
nor U16784 (N_16784,N_16040,N_16383);
and U16785 (N_16785,N_16373,N_16129);
nand U16786 (N_16786,N_16259,N_16291);
and U16787 (N_16787,N_16456,N_16311);
xnor U16788 (N_16788,N_16014,N_16152);
nand U16789 (N_16789,N_16306,N_16278);
or U16790 (N_16790,N_16232,N_16450);
or U16791 (N_16791,N_16408,N_16214);
nor U16792 (N_16792,N_16443,N_16066);
nor U16793 (N_16793,N_16284,N_16061);
nand U16794 (N_16794,N_16439,N_16157);
nor U16795 (N_16795,N_16090,N_16210);
and U16796 (N_16796,N_16365,N_16256);
and U16797 (N_16797,N_16367,N_16240);
nand U16798 (N_16798,N_16343,N_16328);
xnor U16799 (N_16799,N_16016,N_16428);
and U16800 (N_16800,N_16167,N_16077);
and U16801 (N_16801,N_16024,N_16270);
and U16802 (N_16802,N_16316,N_16016);
nand U16803 (N_16803,N_16471,N_16440);
and U16804 (N_16804,N_16125,N_16129);
and U16805 (N_16805,N_16110,N_16275);
and U16806 (N_16806,N_16180,N_16330);
or U16807 (N_16807,N_16036,N_16125);
nand U16808 (N_16808,N_16186,N_16318);
nor U16809 (N_16809,N_16034,N_16103);
nand U16810 (N_16810,N_16235,N_16323);
nor U16811 (N_16811,N_16360,N_16163);
xor U16812 (N_16812,N_16078,N_16288);
and U16813 (N_16813,N_16364,N_16400);
or U16814 (N_16814,N_16301,N_16158);
nand U16815 (N_16815,N_16101,N_16195);
nor U16816 (N_16816,N_16234,N_16139);
nor U16817 (N_16817,N_16411,N_16097);
nand U16818 (N_16818,N_16309,N_16171);
nand U16819 (N_16819,N_16303,N_16288);
or U16820 (N_16820,N_16217,N_16028);
and U16821 (N_16821,N_16141,N_16005);
and U16822 (N_16822,N_16052,N_16454);
or U16823 (N_16823,N_16352,N_16411);
and U16824 (N_16824,N_16381,N_16410);
nand U16825 (N_16825,N_16192,N_16232);
xor U16826 (N_16826,N_16261,N_16043);
nor U16827 (N_16827,N_16108,N_16371);
or U16828 (N_16828,N_16053,N_16019);
xnor U16829 (N_16829,N_16247,N_16437);
or U16830 (N_16830,N_16464,N_16152);
nand U16831 (N_16831,N_16003,N_16108);
xnor U16832 (N_16832,N_16369,N_16340);
nor U16833 (N_16833,N_16219,N_16028);
xor U16834 (N_16834,N_16400,N_16081);
and U16835 (N_16835,N_16430,N_16470);
and U16836 (N_16836,N_16233,N_16223);
nor U16837 (N_16837,N_16057,N_16171);
nand U16838 (N_16838,N_16459,N_16142);
xor U16839 (N_16839,N_16452,N_16398);
nand U16840 (N_16840,N_16368,N_16256);
xor U16841 (N_16841,N_16243,N_16398);
and U16842 (N_16842,N_16063,N_16376);
nand U16843 (N_16843,N_16406,N_16121);
or U16844 (N_16844,N_16237,N_16398);
nand U16845 (N_16845,N_16393,N_16105);
nor U16846 (N_16846,N_16416,N_16322);
and U16847 (N_16847,N_16360,N_16067);
nor U16848 (N_16848,N_16150,N_16355);
and U16849 (N_16849,N_16134,N_16057);
nor U16850 (N_16850,N_16411,N_16026);
xor U16851 (N_16851,N_16276,N_16418);
or U16852 (N_16852,N_16455,N_16179);
nand U16853 (N_16853,N_16346,N_16284);
and U16854 (N_16854,N_16462,N_16320);
nor U16855 (N_16855,N_16432,N_16053);
or U16856 (N_16856,N_16410,N_16320);
or U16857 (N_16857,N_16185,N_16445);
and U16858 (N_16858,N_16267,N_16316);
or U16859 (N_16859,N_16166,N_16340);
nor U16860 (N_16860,N_16338,N_16379);
xnor U16861 (N_16861,N_16063,N_16194);
xnor U16862 (N_16862,N_16424,N_16468);
nor U16863 (N_16863,N_16463,N_16392);
nor U16864 (N_16864,N_16436,N_16058);
and U16865 (N_16865,N_16440,N_16206);
xor U16866 (N_16866,N_16120,N_16221);
and U16867 (N_16867,N_16265,N_16086);
and U16868 (N_16868,N_16356,N_16106);
and U16869 (N_16869,N_16201,N_16260);
or U16870 (N_16870,N_16260,N_16466);
nor U16871 (N_16871,N_16100,N_16134);
or U16872 (N_16872,N_16484,N_16354);
and U16873 (N_16873,N_16440,N_16152);
nand U16874 (N_16874,N_16002,N_16433);
nor U16875 (N_16875,N_16251,N_16237);
nand U16876 (N_16876,N_16388,N_16234);
nor U16877 (N_16877,N_16266,N_16149);
nand U16878 (N_16878,N_16214,N_16028);
and U16879 (N_16879,N_16287,N_16458);
nor U16880 (N_16880,N_16416,N_16374);
or U16881 (N_16881,N_16357,N_16033);
nor U16882 (N_16882,N_16333,N_16088);
or U16883 (N_16883,N_16385,N_16473);
nor U16884 (N_16884,N_16154,N_16039);
nor U16885 (N_16885,N_16470,N_16121);
or U16886 (N_16886,N_16062,N_16415);
nand U16887 (N_16887,N_16313,N_16450);
xor U16888 (N_16888,N_16128,N_16115);
and U16889 (N_16889,N_16433,N_16396);
or U16890 (N_16890,N_16045,N_16127);
or U16891 (N_16891,N_16148,N_16013);
nand U16892 (N_16892,N_16206,N_16047);
nor U16893 (N_16893,N_16386,N_16406);
and U16894 (N_16894,N_16175,N_16369);
and U16895 (N_16895,N_16154,N_16272);
and U16896 (N_16896,N_16050,N_16465);
and U16897 (N_16897,N_16294,N_16137);
and U16898 (N_16898,N_16458,N_16022);
and U16899 (N_16899,N_16097,N_16240);
or U16900 (N_16900,N_16138,N_16210);
and U16901 (N_16901,N_16096,N_16425);
or U16902 (N_16902,N_16482,N_16408);
nor U16903 (N_16903,N_16294,N_16414);
nand U16904 (N_16904,N_16101,N_16093);
nor U16905 (N_16905,N_16011,N_16086);
or U16906 (N_16906,N_16457,N_16444);
and U16907 (N_16907,N_16373,N_16189);
xor U16908 (N_16908,N_16075,N_16185);
or U16909 (N_16909,N_16209,N_16449);
or U16910 (N_16910,N_16201,N_16008);
nand U16911 (N_16911,N_16239,N_16452);
nand U16912 (N_16912,N_16285,N_16206);
and U16913 (N_16913,N_16141,N_16107);
and U16914 (N_16914,N_16124,N_16267);
and U16915 (N_16915,N_16403,N_16170);
or U16916 (N_16916,N_16168,N_16477);
nor U16917 (N_16917,N_16482,N_16421);
or U16918 (N_16918,N_16178,N_16470);
nor U16919 (N_16919,N_16340,N_16036);
or U16920 (N_16920,N_16175,N_16065);
nor U16921 (N_16921,N_16298,N_16321);
xor U16922 (N_16922,N_16157,N_16136);
and U16923 (N_16923,N_16387,N_16194);
nor U16924 (N_16924,N_16060,N_16344);
nand U16925 (N_16925,N_16413,N_16034);
or U16926 (N_16926,N_16236,N_16066);
xnor U16927 (N_16927,N_16026,N_16088);
nor U16928 (N_16928,N_16086,N_16016);
nor U16929 (N_16929,N_16374,N_16077);
or U16930 (N_16930,N_16105,N_16339);
nor U16931 (N_16931,N_16365,N_16210);
nor U16932 (N_16932,N_16301,N_16235);
and U16933 (N_16933,N_16368,N_16247);
nand U16934 (N_16934,N_16310,N_16466);
nand U16935 (N_16935,N_16148,N_16150);
nor U16936 (N_16936,N_16066,N_16127);
or U16937 (N_16937,N_16170,N_16037);
nand U16938 (N_16938,N_16163,N_16011);
and U16939 (N_16939,N_16340,N_16439);
nor U16940 (N_16940,N_16105,N_16351);
nor U16941 (N_16941,N_16148,N_16003);
xor U16942 (N_16942,N_16285,N_16069);
nand U16943 (N_16943,N_16206,N_16198);
nand U16944 (N_16944,N_16363,N_16395);
nand U16945 (N_16945,N_16483,N_16356);
or U16946 (N_16946,N_16221,N_16246);
nor U16947 (N_16947,N_16032,N_16223);
or U16948 (N_16948,N_16088,N_16216);
xnor U16949 (N_16949,N_16082,N_16179);
nand U16950 (N_16950,N_16411,N_16180);
nand U16951 (N_16951,N_16217,N_16048);
and U16952 (N_16952,N_16256,N_16435);
or U16953 (N_16953,N_16296,N_16423);
xor U16954 (N_16954,N_16488,N_16317);
nand U16955 (N_16955,N_16285,N_16411);
xor U16956 (N_16956,N_16254,N_16301);
nor U16957 (N_16957,N_16374,N_16290);
and U16958 (N_16958,N_16320,N_16170);
nand U16959 (N_16959,N_16091,N_16010);
nand U16960 (N_16960,N_16134,N_16198);
nand U16961 (N_16961,N_16059,N_16176);
nand U16962 (N_16962,N_16384,N_16239);
nor U16963 (N_16963,N_16206,N_16409);
nand U16964 (N_16964,N_16071,N_16197);
and U16965 (N_16965,N_16150,N_16163);
nand U16966 (N_16966,N_16160,N_16278);
nor U16967 (N_16967,N_16422,N_16370);
and U16968 (N_16968,N_16076,N_16014);
nand U16969 (N_16969,N_16016,N_16156);
nand U16970 (N_16970,N_16431,N_16252);
or U16971 (N_16971,N_16094,N_16444);
nand U16972 (N_16972,N_16050,N_16252);
and U16973 (N_16973,N_16301,N_16382);
nand U16974 (N_16974,N_16071,N_16310);
and U16975 (N_16975,N_16414,N_16035);
nand U16976 (N_16976,N_16095,N_16126);
nor U16977 (N_16977,N_16461,N_16255);
and U16978 (N_16978,N_16450,N_16071);
and U16979 (N_16979,N_16234,N_16205);
nor U16980 (N_16980,N_16412,N_16465);
nand U16981 (N_16981,N_16204,N_16336);
and U16982 (N_16982,N_16291,N_16072);
or U16983 (N_16983,N_16285,N_16419);
nor U16984 (N_16984,N_16033,N_16324);
nand U16985 (N_16985,N_16281,N_16208);
nor U16986 (N_16986,N_16284,N_16354);
nor U16987 (N_16987,N_16315,N_16120);
nand U16988 (N_16988,N_16368,N_16430);
nor U16989 (N_16989,N_16486,N_16081);
or U16990 (N_16990,N_16079,N_16367);
nor U16991 (N_16991,N_16073,N_16016);
and U16992 (N_16992,N_16388,N_16349);
or U16993 (N_16993,N_16442,N_16177);
or U16994 (N_16994,N_16051,N_16229);
or U16995 (N_16995,N_16299,N_16118);
or U16996 (N_16996,N_16489,N_16237);
and U16997 (N_16997,N_16409,N_16482);
nand U16998 (N_16998,N_16113,N_16286);
or U16999 (N_16999,N_16468,N_16170);
or U17000 (N_17000,N_16795,N_16960);
nor U17001 (N_17001,N_16609,N_16754);
nand U17002 (N_17002,N_16798,N_16781);
nand U17003 (N_17003,N_16921,N_16610);
nand U17004 (N_17004,N_16592,N_16856);
nand U17005 (N_17005,N_16737,N_16603);
and U17006 (N_17006,N_16615,N_16863);
nor U17007 (N_17007,N_16529,N_16706);
nand U17008 (N_17008,N_16952,N_16812);
and U17009 (N_17009,N_16837,N_16702);
and U17010 (N_17010,N_16721,N_16792);
and U17011 (N_17011,N_16848,N_16855);
or U17012 (N_17012,N_16885,N_16653);
and U17013 (N_17013,N_16690,N_16916);
nand U17014 (N_17014,N_16934,N_16540);
nand U17015 (N_17015,N_16555,N_16849);
xor U17016 (N_17016,N_16749,N_16973);
and U17017 (N_17017,N_16533,N_16753);
nor U17018 (N_17018,N_16810,N_16931);
nor U17019 (N_17019,N_16865,N_16731);
nor U17020 (N_17020,N_16878,N_16707);
nand U17021 (N_17021,N_16532,N_16995);
and U17022 (N_17022,N_16616,N_16694);
nor U17023 (N_17023,N_16606,N_16709);
nor U17024 (N_17024,N_16806,N_16770);
nand U17025 (N_17025,N_16791,N_16745);
nor U17026 (N_17026,N_16773,N_16646);
or U17027 (N_17027,N_16583,N_16826);
and U17028 (N_17028,N_16612,N_16638);
nor U17029 (N_17029,N_16501,N_16539);
nand U17030 (N_17030,N_16752,N_16652);
nor U17031 (N_17031,N_16777,N_16663);
and U17032 (N_17032,N_16534,N_16516);
xor U17033 (N_17033,N_16824,N_16624);
or U17034 (N_17034,N_16928,N_16665);
or U17035 (N_17035,N_16695,N_16667);
nor U17036 (N_17036,N_16966,N_16743);
or U17037 (N_17037,N_16608,N_16808);
or U17038 (N_17038,N_16658,N_16935);
nand U17039 (N_17039,N_16988,N_16860);
nor U17040 (N_17040,N_16922,N_16760);
nor U17041 (N_17041,N_16799,N_16835);
nor U17042 (N_17042,N_16957,N_16677);
and U17043 (N_17043,N_16660,N_16746);
or U17044 (N_17044,N_16984,N_16953);
and U17045 (N_17045,N_16742,N_16593);
nand U17046 (N_17046,N_16871,N_16989);
or U17047 (N_17047,N_16940,N_16767);
nand U17048 (N_17048,N_16523,N_16979);
and U17049 (N_17049,N_16589,N_16904);
nor U17050 (N_17050,N_16570,N_16964);
or U17051 (N_17051,N_16599,N_16802);
or U17052 (N_17052,N_16554,N_16967);
nor U17053 (N_17053,N_16897,N_16633);
nand U17054 (N_17054,N_16733,N_16869);
nand U17055 (N_17055,N_16821,N_16634);
nand U17056 (N_17056,N_16669,N_16977);
and U17057 (N_17057,N_16951,N_16990);
and U17058 (N_17058,N_16873,N_16668);
nor U17059 (N_17059,N_16672,N_16684);
nand U17060 (N_17060,N_16854,N_16825);
or U17061 (N_17061,N_16582,N_16775);
nor U17062 (N_17062,N_16870,N_16755);
nor U17063 (N_17063,N_16794,N_16561);
or U17064 (N_17064,N_16576,N_16717);
xnor U17065 (N_17065,N_16783,N_16866);
xor U17066 (N_17066,N_16628,N_16782);
nand U17067 (N_17067,N_16963,N_16600);
and U17068 (N_17068,N_16585,N_16632);
or U17069 (N_17069,N_16759,N_16840);
nand U17070 (N_17070,N_16649,N_16828);
nand U17071 (N_17071,N_16899,N_16574);
or U17072 (N_17072,N_16772,N_16903);
and U17073 (N_17073,N_16682,N_16568);
or U17074 (N_17074,N_16542,N_16898);
or U17075 (N_17075,N_16722,N_16734);
and U17076 (N_17076,N_16862,N_16919);
nor U17077 (N_17077,N_16641,N_16565);
nand U17078 (N_17078,N_16937,N_16617);
and U17079 (N_17079,N_16836,N_16738);
and U17080 (N_17080,N_16805,N_16933);
xnor U17081 (N_17081,N_16572,N_16506);
nor U17082 (N_17082,N_16502,N_16605);
or U17083 (N_17083,N_16685,N_16528);
nand U17084 (N_17084,N_16732,N_16526);
nand U17085 (N_17085,N_16908,N_16689);
xnor U17086 (N_17086,N_16882,N_16673);
nor U17087 (N_17087,N_16947,N_16710);
or U17088 (N_17088,N_16842,N_16822);
xor U17089 (N_17089,N_16944,N_16776);
nand U17090 (N_17090,N_16699,N_16939);
and U17091 (N_17091,N_16946,N_16573);
or U17092 (N_17092,N_16861,N_16591);
or U17093 (N_17093,N_16728,N_16942);
nand U17094 (N_17094,N_16906,N_16962);
xor U17095 (N_17095,N_16761,N_16692);
or U17096 (N_17096,N_16705,N_16851);
or U17097 (N_17097,N_16588,N_16793);
nand U17098 (N_17098,N_16981,N_16896);
or U17099 (N_17099,N_16748,N_16510);
nor U17100 (N_17100,N_16744,N_16713);
xor U17101 (N_17101,N_16872,N_16567);
nor U17102 (N_17102,N_16718,N_16549);
and U17103 (N_17103,N_16558,N_16530);
nand U17104 (N_17104,N_16521,N_16762);
xnor U17105 (N_17105,N_16524,N_16954);
nor U17106 (N_17106,N_16676,N_16971);
nor U17107 (N_17107,N_16881,N_16618);
nand U17108 (N_17108,N_16643,N_16726);
nand U17109 (N_17109,N_16535,N_16790);
nor U17110 (N_17110,N_16587,N_16531);
nand U17111 (N_17111,N_16843,N_16804);
nand U17112 (N_17112,N_16562,N_16985);
or U17113 (N_17113,N_16635,N_16581);
nand U17114 (N_17114,N_16938,N_16846);
nand U17115 (N_17115,N_16723,N_16893);
and U17116 (N_17116,N_16758,N_16509);
nand U17117 (N_17117,N_16703,N_16980);
nor U17118 (N_17118,N_16797,N_16719);
nor U17119 (N_17119,N_16818,N_16909);
or U17120 (N_17120,N_16575,N_16642);
nor U17121 (N_17121,N_16974,N_16890);
or U17122 (N_17122,N_16820,N_16864);
nand U17123 (N_17123,N_16785,N_16912);
nand U17124 (N_17124,N_16675,N_16997);
xor U17125 (N_17125,N_16538,N_16936);
nor U17126 (N_17126,N_16994,N_16858);
or U17127 (N_17127,N_16741,N_16780);
or U17128 (N_17128,N_16730,N_16827);
nor U17129 (N_17129,N_16522,N_16630);
nand U17130 (N_17130,N_16640,N_16815);
nand U17131 (N_17131,N_16811,N_16800);
and U17132 (N_17132,N_16739,N_16894);
nor U17133 (N_17133,N_16626,N_16832);
nor U17134 (N_17134,N_16631,N_16704);
xnor U17135 (N_17135,N_16786,N_16902);
and U17136 (N_17136,N_16886,N_16647);
nand U17137 (N_17137,N_16735,N_16596);
nand U17138 (N_17138,N_16648,N_16955);
nand U17139 (N_17139,N_16883,N_16779);
xor U17140 (N_17140,N_16627,N_16801);
and U17141 (N_17141,N_16680,N_16838);
xnor U17142 (N_17142,N_16765,N_16740);
nand U17143 (N_17143,N_16519,N_16578);
and U17144 (N_17144,N_16504,N_16943);
and U17145 (N_17145,N_16662,N_16517);
and U17146 (N_17146,N_16661,N_16819);
nand U17147 (N_17147,N_16888,N_16978);
nand U17148 (N_17148,N_16725,N_16637);
and U17149 (N_17149,N_16857,N_16545);
or U17150 (N_17150,N_16927,N_16543);
or U17151 (N_17151,N_16945,N_16691);
and U17152 (N_17152,N_16727,N_16859);
nand U17153 (N_17153,N_16715,N_16604);
nand U17154 (N_17154,N_16999,N_16751);
and U17155 (N_17155,N_16518,N_16625);
and U17156 (N_17156,N_16551,N_16507);
or U17157 (N_17157,N_16500,N_16674);
xor U17158 (N_17158,N_16907,N_16756);
nand U17159 (N_17159,N_16602,N_16678);
nor U17160 (N_17160,N_16544,N_16830);
nand U17161 (N_17161,N_16564,N_16853);
nor U17162 (N_17162,N_16763,N_16569);
nor U17163 (N_17163,N_16993,N_16693);
or U17164 (N_17164,N_16619,N_16900);
xor U17165 (N_17165,N_16956,N_16764);
nor U17166 (N_17166,N_16926,N_16918);
or U17167 (N_17167,N_16959,N_16976);
xor U17168 (N_17168,N_16813,N_16520);
and U17169 (N_17169,N_16852,N_16525);
or U17170 (N_17170,N_16586,N_16829);
and U17171 (N_17171,N_16910,N_16670);
or U17172 (N_17172,N_16914,N_16948);
nand U17173 (N_17173,N_16823,N_16636);
nand U17174 (N_17174,N_16778,N_16874);
or U17175 (N_17175,N_16996,N_16654);
nand U17176 (N_17176,N_16972,N_16867);
nor U17177 (N_17177,N_16560,N_16503);
or U17178 (N_17178,N_16716,N_16879);
and U17179 (N_17179,N_16789,N_16803);
nor U17180 (N_17180,N_16766,N_16969);
nor U17181 (N_17181,N_16708,N_16548);
nor U17182 (N_17182,N_16563,N_16998);
nand U17183 (N_17183,N_16650,N_16831);
nor U17184 (N_17184,N_16712,N_16924);
nor U17185 (N_17185,N_16970,N_16657);
nand U17186 (N_17186,N_16769,N_16687);
nand U17187 (N_17187,N_16511,N_16887);
nor U17188 (N_17188,N_16913,N_16788);
nand U17189 (N_17189,N_16991,N_16736);
nor U17190 (N_17190,N_16553,N_16697);
and U17191 (N_17191,N_16850,N_16590);
nand U17192 (N_17192,N_16537,N_16527);
or U17193 (N_17193,N_16556,N_16639);
xnor U17194 (N_17194,N_16929,N_16714);
or U17195 (N_17195,N_16536,N_16958);
nor U17196 (N_17196,N_16645,N_16659);
xnor U17197 (N_17197,N_16941,N_16598);
nor U17198 (N_17198,N_16513,N_16774);
and U17199 (N_17199,N_16750,N_16514);
and U17200 (N_17200,N_16546,N_16656);
and U17201 (N_17201,N_16949,N_16688);
nor U17202 (N_17202,N_16595,N_16986);
nand U17203 (N_17203,N_16877,N_16584);
and U17204 (N_17204,N_16796,N_16920);
xor U17205 (N_17205,N_16757,N_16925);
and U17206 (N_17206,N_16620,N_16629);
nand U17207 (N_17207,N_16845,N_16968);
or U17208 (N_17208,N_16839,N_16901);
nor U17209 (N_17209,N_16601,N_16817);
nand U17210 (N_17210,N_16550,N_16607);
nand U17211 (N_17211,N_16559,N_16580);
nand U17212 (N_17212,N_16505,N_16983);
or U17213 (N_17213,N_16784,N_16681);
and U17214 (N_17214,N_16891,N_16579);
or U17215 (N_17215,N_16923,N_16622);
or U17216 (N_17216,N_16787,N_16847);
nor U17217 (N_17217,N_16679,N_16651);
and U17218 (N_17218,N_16686,N_16597);
nor U17219 (N_17219,N_16720,N_16992);
nand U17220 (N_17220,N_16771,N_16594);
nor U17221 (N_17221,N_16698,N_16809);
nand U17222 (N_17222,N_16950,N_16930);
nor U17223 (N_17223,N_16768,N_16700);
nor U17224 (N_17224,N_16889,N_16621);
nor U17225 (N_17225,N_16932,N_16729);
nand U17226 (N_17226,N_16987,N_16844);
and U17227 (N_17227,N_16613,N_16814);
and U17228 (N_17228,N_16611,N_16975);
nor U17229 (N_17229,N_16961,N_16868);
and U17230 (N_17230,N_16696,N_16683);
nand U17231 (N_17231,N_16833,N_16515);
and U17232 (N_17232,N_16884,N_16905);
nor U17233 (N_17233,N_16701,N_16747);
xnor U17234 (N_17234,N_16911,N_16552);
nor U17235 (N_17235,N_16547,N_16724);
nor U17236 (N_17236,N_16982,N_16965);
nand U17237 (N_17237,N_16711,N_16614);
xor U17238 (N_17238,N_16644,N_16816);
or U17239 (N_17239,N_16566,N_16571);
nor U17240 (N_17240,N_16508,N_16557);
nor U17241 (N_17241,N_16892,N_16577);
nand U17242 (N_17242,N_16915,N_16666);
nand U17243 (N_17243,N_16541,N_16917);
nor U17244 (N_17244,N_16876,N_16895);
nand U17245 (N_17245,N_16841,N_16623);
nor U17246 (N_17246,N_16655,N_16880);
xnor U17247 (N_17247,N_16664,N_16512);
or U17248 (N_17248,N_16807,N_16834);
or U17249 (N_17249,N_16875,N_16671);
and U17250 (N_17250,N_16981,N_16941);
or U17251 (N_17251,N_16573,N_16774);
or U17252 (N_17252,N_16772,N_16672);
or U17253 (N_17253,N_16632,N_16807);
or U17254 (N_17254,N_16728,N_16788);
or U17255 (N_17255,N_16935,N_16694);
nor U17256 (N_17256,N_16677,N_16844);
nor U17257 (N_17257,N_16805,N_16618);
xor U17258 (N_17258,N_16622,N_16649);
or U17259 (N_17259,N_16505,N_16674);
nor U17260 (N_17260,N_16672,N_16850);
or U17261 (N_17261,N_16595,N_16560);
nor U17262 (N_17262,N_16777,N_16771);
and U17263 (N_17263,N_16972,N_16625);
nor U17264 (N_17264,N_16572,N_16897);
and U17265 (N_17265,N_16762,N_16953);
nand U17266 (N_17266,N_16728,N_16779);
or U17267 (N_17267,N_16543,N_16728);
nand U17268 (N_17268,N_16948,N_16902);
nand U17269 (N_17269,N_16550,N_16609);
nand U17270 (N_17270,N_16574,N_16941);
or U17271 (N_17271,N_16576,N_16533);
nand U17272 (N_17272,N_16510,N_16828);
and U17273 (N_17273,N_16578,N_16680);
or U17274 (N_17274,N_16789,N_16864);
nor U17275 (N_17275,N_16581,N_16965);
nor U17276 (N_17276,N_16604,N_16642);
nor U17277 (N_17277,N_16952,N_16822);
and U17278 (N_17278,N_16821,N_16745);
or U17279 (N_17279,N_16741,N_16581);
or U17280 (N_17280,N_16961,N_16582);
xor U17281 (N_17281,N_16898,N_16958);
xnor U17282 (N_17282,N_16940,N_16952);
xnor U17283 (N_17283,N_16735,N_16532);
nand U17284 (N_17284,N_16508,N_16881);
nand U17285 (N_17285,N_16635,N_16853);
and U17286 (N_17286,N_16532,N_16779);
nand U17287 (N_17287,N_16505,N_16863);
nand U17288 (N_17288,N_16821,N_16670);
nor U17289 (N_17289,N_16916,N_16914);
or U17290 (N_17290,N_16738,N_16750);
or U17291 (N_17291,N_16667,N_16753);
or U17292 (N_17292,N_16514,N_16507);
or U17293 (N_17293,N_16947,N_16856);
nand U17294 (N_17294,N_16630,N_16856);
nand U17295 (N_17295,N_16754,N_16544);
and U17296 (N_17296,N_16517,N_16726);
and U17297 (N_17297,N_16531,N_16751);
and U17298 (N_17298,N_16654,N_16881);
nor U17299 (N_17299,N_16555,N_16693);
nand U17300 (N_17300,N_16751,N_16514);
nor U17301 (N_17301,N_16821,N_16831);
or U17302 (N_17302,N_16757,N_16559);
nor U17303 (N_17303,N_16923,N_16566);
xnor U17304 (N_17304,N_16921,N_16669);
or U17305 (N_17305,N_16924,N_16505);
or U17306 (N_17306,N_16556,N_16991);
xnor U17307 (N_17307,N_16914,N_16742);
and U17308 (N_17308,N_16932,N_16684);
xnor U17309 (N_17309,N_16707,N_16714);
nand U17310 (N_17310,N_16653,N_16509);
nand U17311 (N_17311,N_16818,N_16554);
nor U17312 (N_17312,N_16993,N_16813);
nor U17313 (N_17313,N_16512,N_16543);
and U17314 (N_17314,N_16731,N_16886);
and U17315 (N_17315,N_16952,N_16730);
nand U17316 (N_17316,N_16694,N_16583);
nor U17317 (N_17317,N_16777,N_16957);
nand U17318 (N_17318,N_16730,N_16762);
nand U17319 (N_17319,N_16792,N_16848);
and U17320 (N_17320,N_16844,N_16970);
nand U17321 (N_17321,N_16519,N_16989);
and U17322 (N_17322,N_16779,N_16639);
or U17323 (N_17323,N_16542,N_16980);
nand U17324 (N_17324,N_16525,N_16567);
or U17325 (N_17325,N_16747,N_16975);
nor U17326 (N_17326,N_16884,N_16533);
xnor U17327 (N_17327,N_16997,N_16886);
or U17328 (N_17328,N_16634,N_16746);
nor U17329 (N_17329,N_16924,N_16948);
and U17330 (N_17330,N_16841,N_16848);
or U17331 (N_17331,N_16694,N_16837);
or U17332 (N_17332,N_16788,N_16623);
and U17333 (N_17333,N_16744,N_16676);
or U17334 (N_17334,N_16648,N_16613);
nor U17335 (N_17335,N_16793,N_16777);
xor U17336 (N_17336,N_16887,N_16741);
nand U17337 (N_17337,N_16596,N_16584);
nand U17338 (N_17338,N_16511,N_16551);
nand U17339 (N_17339,N_16811,N_16803);
or U17340 (N_17340,N_16919,N_16518);
and U17341 (N_17341,N_16530,N_16553);
and U17342 (N_17342,N_16977,N_16748);
xor U17343 (N_17343,N_16641,N_16798);
xnor U17344 (N_17344,N_16917,N_16767);
or U17345 (N_17345,N_16950,N_16998);
nand U17346 (N_17346,N_16952,N_16830);
and U17347 (N_17347,N_16948,N_16539);
nand U17348 (N_17348,N_16723,N_16724);
nor U17349 (N_17349,N_16897,N_16716);
or U17350 (N_17350,N_16757,N_16804);
nor U17351 (N_17351,N_16973,N_16610);
nor U17352 (N_17352,N_16553,N_16983);
xor U17353 (N_17353,N_16698,N_16777);
and U17354 (N_17354,N_16680,N_16556);
and U17355 (N_17355,N_16560,N_16786);
nand U17356 (N_17356,N_16884,N_16873);
xnor U17357 (N_17357,N_16733,N_16780);
nor U17358 (N_17358,N_16540,N_16730);
nand U17359 (N_17359,N_16604,N_16618);
nand U17360 (N_17360,N_16558,N_16937);
or U17361 (N_17361,N_16860,N_16896);
and U17362 (N_17362,N_16820,N_16980);
nand U17363 (N_17363,N_16990,N_16511);
nor U17364 (N_17364,N_16536,N_16534);
xor U17365 (N_17365,N_16532,N_16596);
nor U17366 (N_17366,N_16706,N_16525);
and U17367 (N_17367,N_16526,N_16877);
nand U17368 (N_17368,N_16991,N_16808);
xnor U17369 (N_17369,N_16819,N_16791);
nor U17370 (N_17370,N_16891,N_16743);
nor U17371 (N_17371,N_16675,N_16593);
nand U17372 (N_17372,N_16682,N_16541);
nand U17373 (N_17373,N_16878,N_16999);
nand U17374 (N_17374,N_16804,N_16719);
nor U17375 (N_17375,N_16892,N_16833);
nand U17376 (N_17376,N_16868,N_16662);
xor U17377 (N_17377,N_16870,N_16685);
and U17378 (N_17378,N_16839,N_16974);
nor U17379 (N_17379,N_16785,N_16906);
nand U17380 (N_17380,N_16758,N_16558);
nand U17381 (N_17381,N_16548,N_16969);
and U17382 (N_17382,N_16975,N_16650);
xor U17383 (N_17383,N_16887,N_16737);
nor U17384 (N_17384,N_16597,N_16809);
nand U17385 (N_17385,N_16838,N_16989);
nand U17386 (N_17386,N_16957,N_16575);
or U17387 (N_17387,N_16676,N_16637);
nor U17388 (N_17388,N_16572,N_16566);
nor U17389 (N_17389,N_16759,N_16657);
xnor U17390 (N_17390,N_16899,N_16898);
or U17391 (N_17391,N_16752,N_16571);
nor U17392 (N_17392,N_16661,N_16856);
xor U17393 (N_17393,N_16821,N_16581);
nor U17394 (N_17394,N_16801,N_16951);
nor U17395 (N_17395,N_16658,N_16508);
nor U17396 (N_17396,N_16910,N_16691);
xor U17397 (N_17397,N_16633,N_16504);
and U17398 (N_17398,N_16751,N_16710);
xnor U17399 (N_17399,N_16794,N_16873);
xnor U17400 (N_17400,N_16741,N_16858);
nor U17401 (N_17401,N_16764,N_16671);
nor U17402 (N_17402,N_16708,N_16897);
nor U17403 (N_17403,N_16911,N_16577);
or U17404 (N_17404,N_16537,N_16600);
and U17405 (N_17405,N_16932,N_16840);
nand U17406 (N_17406,N_16693,N_16848);
nand U17407 (N_17407,N_16749,N_16606);
and U17408 (N_17408,N_16765,N_16616);
nor U17409 (N_17409,N_16977,N_16611);
and U17410 (N_17410,N_16960,N_16917);
nand U17411 (N_17411,N_16992,N_16595);
nor U17412 (N_17412,N_16851,N_16770);
or U17413 (N_17413,N_16641,N_16719);
nand U17414 (N_17414,N_16638,N_16884);
or U17415 (N_17415,N_16505,N_16860);
nand U17416 (N_17416,N_16568,N_16839);
xor U17417 (N_17417,N_16957,N_16572);
or U17418 (N_17418,N_16969,N_16695);
nand U17419 (N_17419,N_16639,N_16586);
xnor U17420 (N_17420,N_16962,N_16539);
xor U17421 (N_17421,N_16845,N_16792);
nor U17422 (N_17422,N_16918,N_16792);
nor U17423 (N_17423,N_16536,N_16895);
nor U17424 (N_17424,N_16823,N_16511);
nor U17425 (N_17425,N_16737,N_16676);
xor U17426 (N_17426,N_16802,N_16778);
nor U17427 (N_17427,N_16559,N_16805);
nand U17428 (N_17428,N_16740,N_16694);
or U17429 (N_17429,N_16847,N_16749);
nor U17430 (N_17430,N_16858,N_16558);
nor U17431 (N_17431,N_16968,N_16854);
and U17432 (N_17432,N_16880,N_16992);
nand U17433 (N_17433,N_16793,N_16840);
nand U17434 (N_17434,N_16958,N_16860);
nand U17435 (N_17435,N_16820,N_16829);
and U17436 (N_17436,N_16677,N_16716);
nand U17437 (N_17437,N_16718,N_16544);
or U17438 (N_17438,N_16847,N_16654);
or U17439 (N_17439,N_16830,N_16837);
and U17440 (N_17440,N_16856,N_16727);
and U17441 (N_17441,N_16903,N_16769);
or U17442 (N_17442,N_16579,N_16906);
or U17443 (N_17443,N_16985,N_16519);
and U17444 (N_17444,N_16882,N_16730);
nand U17445 (N_17445,N_16567,N_16652);
and U17446 (N_17446,N_16978,N_16919);
or U17447 (N_17447,N_16739,N_16944);
nor U17448 (N_17448,N_16917,N_16970);
xnor U17449 (N_17449,N_16974,N_16838);
and U17450 (N_17450,N_16505,N_16914);
nor U17451 (N_17451,N_16755,N_16876);
and U17452 (N_17452,N_16506,N_16871);
nand U17453 (N_17453,N_16976,N_16633);
nand U17454 (N_17454,N_16873,N_16587);
and U17455 (N_17455,N_16901,N_16982);
nand U17456 (N_17456,N_16699,N_16629);
or U17457 (N_17457,N_16727,N_16555);
nand U17458 (N_17458,N_16568,N_16587);
or U17459 (N_17459,N_16984,N_16908);
nand U17460 (N_17460,N_16677,N_16988);
nor U17461 (N_17461,N_16550,N_16818);
nor U17462 (N_17462,N_16942,N_16972);
nor U17463 (N_17463,N_16833,N_16823);
and U17464 (N_17464,N_16554,N_16532);
or U17465 (N_17465,N_16570,N_16772);
nand U17466 (N_17466,N_16982,N_16778);
and U17467 (N_17467,N_16903,N_16619);
or U17468 (N_17468,N_16931,N_16643);
nor U17469 (N_17469,N_16644,N_16713);
nand U17470 (N_17470,N_16768,N_16618);
or U17471 (N_17471,N_16715,N_16928);
nand U17472 (N_17472,N_16895,N_16838);
nor U17473 (N_17473,N_16651,N_16984);
nand U17474 (N_17474,N_16993,N_16819);
or U17475 (N_17475,N_16928,N_16673);
or U17476 (N_17476,N_16750,N_16948);
nand U17477 (N_17477,N_16528,N_16655);
or U17478 (N_17478,N_16580,N_16687);
nor U17479 (N_17479,N_16737,N_16641);
nand U17480 (N_17480,N_16837,N_16613);
nand U17481 (N_17481,N_16514,N_16973);
nor U17482 (N_17482,N_16668,N_16538);
nor U17483 (N_17483,N_16734,N_16838);
xor U17484 (N_17484,N_16827,N_16818);
and U17485 (N_17485,N_16641,N_16904);
nand U17486 (N_17486,N_16876,N_16829);
nor U17487 (N_17487,N_16996,N_16644);
xor U17488 (N_17488,N_16741,N_16542);
nand U17489 (N_17489,N_16829,N_16601);
and U17490 (N_17490,N_16864,N_16924);
nand U17491 (N_17491,N_16973,N_16995);
and U17492 (N_17492,N_16989,N_16987);
nor U17493 (N_17493,N_16669,N_16794);
xor U17494 (N_17494,N_16732,N_16563);
and U17495 (N_17495,N_16893,N_16838);
nand U17496 (N_17496,N_16710,N_16954);
xor U17497 (N_17497,N_16799,N_16682);
or U17498 (N_17498,N_16846,N_16698);
or U17499 (N_17499,N_16897,N_16744);
nor U17500 (N_17500,N_17089,N_17252);
and U17501 (N_17501,N_17295,N_17406);
xnor U17502 (N_17502,N_17018,N_17444);
or U17503 (N_17503,N_17293,N_17477);
and U17504 (N_17504,N_17200,N_17288);
nand U17505 (N_17505,N_17178,N_17365);
or U17506 (N_17506,N_17117,N_17268);
or U17507 (N_17507,N_17425,N_17185);
nor U17508 (N_17508,N_17161,N_17375);
nand U17509 (N_17509,N_17186,N_17013);
or U17510 (N_17510,N_17048,N_17120);
xnor U17511 (N_17511,N_17448,N_17203);
or U17512 (N_17512,N_17064,N_17134);
nand U17513 (N_17513,N_17164,N_17224);
and U17514 (N_17514,N_17231,N_17033);
and U17515 (N_17515,N_17184,N_17328);
xnor U17516 (N_17516,N_17223,N_17196);
or U17517 (N_17517,N_17142,N_17286);
nor U17518 (N_17518,N_17060,N_17315);
or U17519 (N_17519,N_17097,N_17219);
nor U17520 (N_17520,N_17449,N_17370);
and U17521 (N_17521,N_17218,N_17266);
nand U17522 (N_17522,N_17055,N_17119);
and U17523 (N_17523,N_17190,N_17020);
and U17524 (N_17524,N_17367,N_17355);
nand U17525 (N_17525,N_17182,N_17150);
nand U17526 (N_17526,N_17351,N_17232);
or U17527 (N_17527,N_17452,N_17007);
or U17528 (N_17528,N_17475,N_17024);
xor U17529 (N_17529,N_17363,N_17493);
xor U17530 (N_17530,N_17366,N_17297);
or U17531 (N_17531,N_17310,N_17095);
nor U17532 (N_17532,N_17377,N_17222);
and U17533 (N_17533,N_17239,N_17245);
or U17534 (N_17534,N_17459,N_17220);
and U17535 (N_17535,N_17430,N_17472);
nor U17536 (N_17536,N_17061,N_17225);
or U17537 (N_17537,N_17262,N_17210);
and U17538 (N_17538,N_17382,N_17454);
and U17539 (N_17539,N_17088,N_17299);
and U17540 (N_17540,N_17306,N_17198);
nand U17541 (N_17541,N_17353,N_17156);
nor U17542 (N_17542,N_17063,N_17499);
xnor U17543 (N_17543,N_17346,N_17169);
and U17544 (N_17544,N_17079,N_17254);
or U17545 (N_17545,N_17285,N_17443);
xor U17546 (N_17546,N_17412,N_17418);
nor U17547 (N_17547,N_17364,N_17241);
nor U17548 (N_17548,N_17374,N_17298);
and U17549 (N_17549,N_17140,N_17307);
nand U17550 (N_17550,N_17221,N_17453);
and U17551 (N_17551,N_17311,N_17162);
nor U17552 (N_17552,N_17242,N_17331);
and U17553 (N_17553,N_17276,N_17300);
and U17554 (N_17554,N_17204,N_17483);
or U17555 (N_17555,N_17442,N_17436);
nand U17556 (N_17556,N_17282,N_17101);
and U17557 (N_17557,N_17209,N_17361);
and U17558 (N_17558,N_17342,N_17168);
and U17559 (N_17559,N_17409,N_17283);
nor U17560 (N_17560,N_17216,N_17113);
or U17561 (N_17561,N_17424,N_17423);
nand U17562 (N_17562,N_17484,N_17265);
and U17563 (N_17563,N_17270,N_17338);
and U17564 (N_17564,N_17093,N_17143);
nand U17565 (N_17565,N_17130,N_17320);
nor U17566 (N_17566,N_17108,N_17133);
nor U17567 (N_17567,N_17422,N_17301);
and U17568 (N_17568,N_17460,N_17012);
and U17569 (N_17569,N_17352,N_17359);
and U17570 (N_17570,N_17098,N_17481);
or U17571 (N_17571,N_17487,N_17376);
nor U17572 (N_17572,N_17362,N_17014);
and U17573 (N_17573,N_17076,N_17465);
and U17574 (N_17574,N_17492,N_17416);
or U17575 (N_17575,N_17305,N_17255);
and U17576 (N_17576,N_17102,N_17144);
nor U17577 (N_17577,N_17358,N_17135);
or U17578 (N_17578,N_17263,N_17159);
and U17579 (N_17579,N_17006,N_17138);
nand U17580 (N_17580,N_17432,N_17345);
and U17581 (N_17581,N_17466,N_17287);
and U17582 (N_17582,N_17294,N_17165);
nor U17583 (N_17583,N_17148,N_17128);
or U17584 (N_17584,N_17371,N_17404);
nand U17585 (N_17585,N_17399,N_17435);
and U17586 (N_17586,N_17084,N_17433);
xnor U17587 (N_17587,N_17304,N_17495);
nor U17588 (N_17588,N_17136,N_17032);
and U17589 (N_17589,N_17192,N_17170);
nor U17590 (N_17590,N_17261,N_17314);
and U17591 (N_17591,N_17176,N_17105);
or U17592 (N_17592,N_17208,N_17290);
and U17593 (N_17593,N_17395,N_17118);
nor U17594 (N_17594,N_17217,N_17236);
xnor U17595 (N_17595,N_17193,N_17405);
or U17596 (N_17596,N_17498,N_17129);
and U17597 (N_17597,N_17446,N_17147);
nand U17598 (N_17598,N_17327,N_17440);
nor U17599 (N_17599,N_17066,N_17330);
nor U17600 (N_17600,N_17069,N_17166);
and U17601 (N_17601,N_17380,N_17271);
nor U17602 (N_17602,N_17302,N_17384);
and U17603 (N_17603,N_17116,N_17123);
and U17604 (N_17604,N_17083,N_17075);
and U17605 (N_17605,N_17068,N_17090);
or U17606 (N_17606,N_17397,N_17378);
or U17607 (N_17607,N_17030,N_17212);
or U17608 (N_17608,N_17078,N_17388);
or U17609 (N_17609,N_17008,N_17369);
nor U17610 (N_17610,N_17158,N_17016);
xor U17611 (N_17611,N_17468,N_17341);
nor U17612 (N_17612,N_17227,N_17189);
xor U17613 (N_17613,N_17272,N_17122);
nand U17614 (N_17614,N_17322,N_17126);
nor U17615 (N_17615,N_17072,N_17277);
and U17616 (N_17616,N_17426,N_17046);
nand U17617 (N_17617,N_17188,N_17009);
nand U17618 (N_17618,N_17321,N_17044);
or U17619 (N_17619,N_17230,N_17039);
nand U17620 (N_17620,N_17031,N_17028);
nand U17621 (N_17621,N_17333,N_17256);
nand U17622 (N_17622,N_17467,N_17050);
xor U17623 (N_17623,N_17368,N_17206);
nand U17624 (N_17624,N_17141,N_17110);
nand U17625 (N_17625,N_17396,N_17323);
or U17626 (N_17626,N_17348,N_17004);
and U17627 (N_17627,N_17478,N_17127);
nand U17628 (N_17628,N_17356,N_17100);
or U17629 (N_17629,N_17260,N_17393);
or U17630 (N_17630,N_17464,N_17211);
or U17631 (N_17631,N_17497,N_17407);
nand U17632 (N_17632,N_17336,N_17002);
or U17633 (N_17633,N_17439,N_17458);
and U17634 (N_17634,N_17146,N_17421);
or U17635 (N_17635,N_17428,N_17080);
nor U17636 (N_17636,N_17427,N_17106);
and U17637 (N_17637,N_17248,N_17480);
nand U17638 (N_17638,N_17081,N_17181);
nor U17639 (N_17639,N_17281,N_17233);
nor U17640 (N_17640,N_17052,N_17434);
or U17641 (N_17641,N_17383,N_17035);
nand U17642 (N_17642,N_17447,N_17099);
or U17643 (N_17643,N_17247,N_17347);
or U17644 (N_17644,N_17019,N_17390);
and U17645 (N_17645,N_17461,N_17034);
or U17646 (N_17646,N_17086,N_17114);
nand U17647 (N_17647,N_17022,N_17400);
or U17648 (N_17648,N_17470,N_17235);
nor U17649 (N_17649,N_17308,N_17091);
and U17650 (N_17650,N_17036,N_17160);
nand U17651 (N_17651,N_17474,N_17414);
and U17652 (N_17652,N_17010,N_17387);
nand U17653 (N_17653,N_17056,N_17391);
and U17654 (N_17654,N_17037,N_17155);
and U17655 (N_17655,N_17386,N_17213);
or U17656 (N_17656,N_17417,N_17462);
and U17657 (N_17657,N_17469,N_17275);
or U17658 (N_17658,N_17456,N_17103);
and U17659 (N_17659,N_17051,N_17175);
nor U17660 (N_17660,N_17372,N_17408);
and U17661 (N_17661,N_17058,N_17292);
and U17662 (N_17662,N_17403,N_17243);
and U17663 (N_17663,N_17071,N_17445);
nand U17664 (N_17664,N_17455,N_17157);
or U17665 (N_17665,N_17049,N_17131);
nor U17666 (N_17666,N_17339,N_17074);
or U17667 (N_17667,N_17488,N_17043);
or U17668 (N_17668,N_17420,N_17023);
or U17669 (N_17669,N_17325,N_17451);
xnor U17670 (N_17670,N_17438,N_17485);
nand U17671 (N_17671,N_17003,N_17429);
or U17672 (N_17672,N_17163,N_17240);
or U17673 (N_17673,N_17017,N_17494);
nand U17674 (N_17674,N_17202,N_17229);
nor U17675 (N_17675,N_17177,N_17179);
nor U17676 (N_17676,N_17154,N_17389);
or U17677 (N_17677,N_17057,N_17350);
and U17678 (N_17678,N_17228,N_17096);
and U17679 (N_17679,N_17324,N_17253);
and U17680 (N_17680,N_17152,N_17332);
nand U17681 (N_17681,N_17289,N_17053);
and U17682 (N_17682,N_17250,N_17145);
nor U17683 (N_17683,N_17385,N_17410);
or U17684 (N_17684,N_17171,N_17392);
or U17685 (N_17685,N_17234,N_17087);
nand U17686 (N_17686,N_17226,N_17278);
nand U17687 (N_17687,N_17137,N_17000);
nand U17688 (N_17688,N_17379,N_17476);
nand U17689 (N_17689,N_17047,N_17038);
and U17690 (N_17690,N_17257,N_17199);
or U17691 (N_17691,N_17174,N_17041);
nor U17692 (N_17692,N_17496,N_17279);
nor U17693 (N_17693,N_17344,N_17490);
nand U17694 (N_17694,N_17360,N_17011);
nand U17695 (N_17695,N_17381,N_17402);
or U17696 (N_17696,N_17132,N_17437);
and U17697 (N_17697,N_17411,N_17045);
nand U17698 (N_17698,N_17197,N_17029);
nor U17699 (N_17699,N_17001,N_17349);
or U17700 (N_17700,N_17025,N_17173);
nor U17701 (N_17701,N_17398,N_17267);
nand U17702 (N_17702,N_17482,N_17062);
nand U17703 (N_17703,N_17191,N_17065);
nand U17704 (N_17704,N_17194,N_17077);
nor U17705 (N_17705,N_17394,N_17104);
and U17706 (N_17706,N_17153,N_17040);
nor U17707 (N_17707,N_17021,N_17115);
xor U17708 (N_17708,N_17172,N_17303);
and U17709 (N_17709,N_17167,N_17258);
nand U17710 (N_17710,N_17246,N_17296);
nand U17711 (N_17711,N_17082,N_17214);
nand U17712 (N_17712,N_17026,N_17251);
nand U17713 (N_17713,N_17085,N_17094);
and U17714 (N_17714,N_17149,N_17431);
or U17715 (N_17715,N_17180,N_17070);
nor U17716 (N_17716,N_17092,N_17124);
nor U17717 (N_17717,N_17054,N_17318);
xnor U17718 (N_17718,N_17357,N_17264);
and U17719 (N_17719,N_17259,N_17015);
or U17720 (N_17720,N_17125,N_17340);
nor U17721 (N_17721,N_17489,N_17269);
xor U17722 (N_17722,N_17413,N_17273);
nand U17723 (N_17723,N_17207,N_17309);
nand U17724 (N_17724,N_17457,N_17354);
nand U17725 (N_17725,N_17316,N_17244);
and U17726 (N_17726,N_17473,N_17042);
and U17727 (N_17727,N_17151,N_17312);
nand U17728 (N_17728,N_17486,N_17326);
nand U17729 (N_17729,N_17334,N_17111);
xor U17730 (N_17730,N_17479,N_17249);
nand U17731 (N_17731,N_17471,N_17280);
or U17732 (N_17732,N_17139,N_17284);
xnor U17733 (N_17733,N_17291,N_17373);
xor U17734 (N_17734,N_17027,N_17005);
nor U17735 (N_17735,N_17183,N_17073);
nor U17736 (N_17736,N_17463,N_17274);
or U17737 (N_17737,N_17059,N_17109);
xnor U17738 (N_17738,N_17450,N_17238);
xnor U17739 (N_17739,N_17337,N_17415);
xor U17740 (N_17740,N_17121,N_17195);
nand U17741 (N_17741,N_17107,N_17201);
and U17742 (N_17742,N_17205,N_17067);
nor U17743 (N_17743,N_17187,N_17329);
and U17744 (N_17744,N_17441,N_17419);
nand U17745 (N_17745,N_17317,N_17237);
nand U17746 (N_17746,N_17313,N_17401);
nand U17747 (N_17747,N_17343,N_17112);
nor U17748 (N_17748,N_17335,N_17491);
and U17749 (N_17749,N_17215,N_17319);
nand U17750 (N_17750,N_17084,N_17201);
nor U17751 (N_17751,N_17009,N_17477);
nand U17752 (N_17752,N_17090,N_17044);
nor U17753 (N_17753,N_17006,N_17089);
or U17754 (N_17754,N_17046,N_17090);
nand U17755 (N_17755,N_17448,N_17343);
or U17756 (N_17756,N_17016,N_17095);
nand U17757 (N_17757,N_17329,N_17029);
nor U17758 (N_17758,N_17351,N_17470);
or U17759 (N_17759,N_17014,N_17265);
and U17760 (N_17760,N_17209,N_17066);
nand U17761 (N_17761,N_17066,N_17367);
and U17762 (N_17762,N_17211,N_17485);
and U17763 (N_17763,N_17255,N_17489);
and U17764 (N_17764,N_17182,N_17165);
nor U17765 (N_17765,N_17372,N_17326);
or U17766 (N_17766,N_17439,N_17030);
xor U17767 (N_17767,N_17233,N_17128);
nand U17768 (N_17768,N_17490,N_17358);
or U17769 (N_17769,N_17319,N_17444);
and U17770 (N_17770,N_17264,N_17164);
nor U17771 (N_17771,N_17131,N_17426);
or U17772 (N_17772,N_17213,N_17303);
and U17773 (N_17773,N_17022,N_17386);
nor U17774 (N_17774,N_17430,N_17440);
xnor U17775 (N_17775,N_17017,N_17287);
and U17776 (N_17776,N_17402,N_17357);
or U17777 (N_17777,N_17028,N_17097);
or U17778 (N_17778,N_17093,N_17214);
nor U17779 (N_17779,N_17209,N_17331);
or U17780 (N_17780,N_17074,N_17331);
and U17781 (N_17781,N_17026,N_17025);
xnor U17782 (N_17782,N_17036,N_17395);
xnor U17783 (N_17783,N_17234,N_17446);
or U17784 (N_17784,N_17119,N_17347);
nor U17785 (N_17785,N_17158,N_17407);
or U17786 (N_17786,N_17429,N_17031);
or U17787 (N_17787,N_17131,N_17314);
or U17788 (N_17788,N_17160,N_17087);
or U17789 (N_17789,N_17008,N_17373);
or U17790 (N_17790,N_17431,N_17391);
and U17791 (N_17791,N_17423,N_17206);
nor U17792 (N_17792,N_17271,N_17245);
xnor U17793 (N_17793,N_17315,N_17178);
nand U17794 (N_17794,N_17175,N_17371);
xnor U17795 (N_17795,N_17229,N_17265);
xnor U17796 (N_17796,N_17197,N_17039);
nand U17797 (N_17797,N_17263,N_17064);
xor U17798 (N_17798,N_17327,N_17468);
or U17799 (N_17799,N_17268,N_17295);
or U17800 (N_17800,N_17236,N_17242);
and U17801 (N_17801,N_17300,N_17415);
and U17802 (N_17802,N_17062,N_17378);
and U17803 (N_17803,N_17352,N_17032);
and U17804 (N_17804,N_17298,N_17190);
and U17805 (N_17805,N_17478,N_17254);
nor U17806 (N_17806,N_17445,N_17107);
nand U17807 (N_17807,N_17044,N_17216);
and U17808 (N_17808,N_17043,N_17113);
nand U17809 (N_17809,N_17182,N_17114);
nor U17810 (N_17810,N_17159,N_17196);
and U17811 (N_17811,N_17052,N_17157);
nand U17812 (N_17812,N_17266,N_17154);
nand U17813 (N_17813,N_17365,N_17004);
nand U17814 (N_17814,N_17403,N_17286);
xor U17815 (N_17815,N_17253,N_17430);
or U17816 (N_17816,N_17431,N_17193);
nor U17817 (N_17817,N_17427,N_17498);
nand U17818 (N_17818,N_17090,N_17407);
nand U17819 (N_17819,N_17085,N_17320);
nor U17820 (N_17820,N_17068,N_17377);
or U17821 (N_17821,N_17469,N_17064);
or U17822 (N_17822,N_17391,N_17275);
nand U17823 (N_17823,N_17154,N_17130);
xnor U17824 (N_17824,N_17228,N_17116);
nand U17825 (N_17825,N_17477,N_17429);
xnor U17826 (N_17826,N_17203,N_17498);
xor U17827 (N_17827,N_17405,N_17492);
nand U17828 (N_17828,N_17322,N_17296);
nor U17829 (N_17829,N_17480,N_17214);
nor U17830 (N_17830,N_17498,N_17140);
nand U17831 (N_17831,N_17490,N_17160);
nand U17832 (N_17832,N_17061,N_17350);
or U17833 (N_17833,N_17425,N_17478);
and U17834 (N_17834,N_17394,N_17461);
nand U17835 (N_17835,N_17074,N_17428);
nand U17836 (N_17836,N_17291,N_17478);
or U17837 (N_17837,N_17454,N_17054);
and U17838 (N_17838,N_17259,N_17457);
nor U17839 (N_17839,N_17295,N_17205);
or U17840 (N_17840,N_17489,N_17149);
and U17841 (N_17841,N_17188,N_17121);
nor U17842 (N_17842,N_17302,N_17404);
nor U17843 (N_17843,N_17223,N_17231);
nand U17844 (N_17844,N_17015,N_17212);
and U17845 (N_17845,N_17029,N_17142);
or U17846 (N_17846,N_17149,N_17343);
and U17847 (N_17847,N_17193,N_17336);
nand U17848 (N_17848,N_17392,N_17167);
or U17849 (N_17849,N_17210,N_17264);
xor U17850 (N_17850,N_17306,N_17349);
nand U17851 (N_17851,N_17149,N_17368);
or U17852 (N_17852,N_17480,N_17397);
or U17853 (N_17853,N_17014,N_17452);
nand U17854 (N_17854,N_17317,N_17294);
or U17855 (N_17855,N_17206,N_17456);
xnor U17856 (N_17856,N_17064,N_17262);
nand U17857 (N_17857,N_17358,N_17107);
nand U17858 (N_17858,N_17371,N_17066);
and U17859 (N_17859,N_17492,N_17420);
nor U17860 (N_17860,N_17222,N_17219);
xor U17861 (N_17861,N_17122,N_17134);
and U17862 (N_17862,N_17443,N_17178);
nand U17863 (N_17863,N_17280,N_17349);
xnor U17864 (N_17864,N_17366,N_17076);
nand U17865 (N_17865,N_17054,N_17075);
and U17866 (N_17866,N_17360,N_17307);
or U17867 (N_17867,N_17008,N_17004);
or U17868 (N_17868,N_17475,N_17020);
and U17869 (N_17869,N_17349,N_17340);
or U17870 (N_17870,N_17059,N_17239);
and U17871 (N_17871,N_17070,N_17186);
nor U17872 (N_17872,N_17014,N_17101);
nor U17873 (N_17873,N_17387,N_17033);
nor U17874 (N_17874,N_17140,N_17009);
xor U17875 (N_17875,N_17262,N_17214);
or U17876 (N_17876,N_17030,N_17169);
and U17877 (N_17877,N_17174,N_17288);
xor U17878 (N_17878,N_17187,N_17161);
and U17879 (N_17879,N_17236,N_17173);
nand U17880 (N_17880,N_17256,N_17484);
or U17881 (N_17881,N_17051,N_17475);
or U17882 (N_17882,N_17428,N_17177);
and U17883 (N_17883,N_17182,N_17121);
nor U17884 (N_17884,N_17453,N_17280);
nor U17885 (N_17885,N_17403,N_17276);
xor U17886 (N_17886,N_17189,N_17279);
xor U17887 (N_17887,N_17412,N_17423);
nor U17888 (N_17888,N_17443,N_17389);
nand U17889 (N_17889,N_17457,N_17083);
xnor U17890 (N_17890,N_17021,N_17407);
nand U17891 (N_17891,N_17230,N_17070);
and U17892 (N_17892,N_17474,N_17124);
or U17893 (N_17893,N_17245,N_17248);
or U17894 (N_17894,N_17032,N_17390);
nor U17895 (N_17895,N_17484,N_17385);
nor U17896 (N_17896,N_17081,N_17225);
and U17897 (N_17897,N_17446,N_17213);
or U17898 (N_17898,N_17197,N_17033);
nor U17899 (N_17899,N_17474,N_17093);
or U17900 (N_17900,N_17307,N_17314);
nand U17901 (N_17901,N_17438,N_17253);
and U17902 (N_17902,N_17216,N_17215);
nor U17903 (N_17903,N_17252,N_17103);
and U17904 (N_17904,N_17169,N_17360);
nor U17905 (N_17905,N_17433,N_17460);
and U17906 (N_17906,N_17484,N_17069);
nor U17907 (N_17907,N_17365,N_17418);
xor U17908 (N_17908,N_17149,N_17445);
or U17909 (N_17909,N_17403,N_17221);
nand U17910 (N_17910,N_17038,N_17252);
and U17911 (N_17911,N_17495,N_17009);
and U17912 (N_17912,N_17322,N_17088);
or U17913 (N_17913,N_17363,N_17240);
or U17914 (N_17914,N_17349,N_17242);
nand U17915 (N_17915,N_17361,N_17341);
and U17916 (N_17916,N_17338,N_17131);
and U17917 (N_17917,N_17156,N_17439);
and U17918 (N_17918,N_17032,N_17158);
or U17919 (N_17919,N_17468,N_17299);
xnor U17920 (N_17920,N_17416,N_17222);
nor U17921 (N_17921,N_17384,N_17472);
nand U17922 (N_17922,N_17316,N_17479);
and U17923 (N_17923,N_17284,N_17022);
and U17924 (N_17924,N_17233,N_17331);
or U17925 (N_17925,N_17424,N_17160);
xor U17926 (N_17926,N_17276,N_17399);
xor U17927 (N_17927,N_17269,N_17155);
or U17928 (N_17928,N_17178,N_17289);
xor U17929 (N_17929,N_17250,N_17044);
or U17930 (N_17930,N_17276,N_17482);
or U17931 (N_17931,N_17001,N_17050);
nor U17932 (N_17932,N_17462,N_17469);
nor U17933 (N_17933,N_17429,N_17380);
and U17934 (N_17934,N_17058,N_17269);
or U17935 (N_17935,N_17020,N_17073);
nor U17936 (N_17936,N_17347,N_17387);
nand U17937 (N_17937,N_17358,N_17290);
nand U17938 (N_17938,N_17060,N_17427);
nor U17939 (N_17939,N_17497,N_17447);
nor U17940 (N_17940,N_17285,N_17148);
nor U17941 (N_17941,N_17347,N_17069);
xor U17942 (N_17942,N_17133,N_17087);
nor U17943 (N_17943,N_17050,N_17403);
nand U17944 (N_17944,N_17254,N_17388);
and U17945 (N_17945,N_17460,N_17091);
and U17946 (N_17946,N_17305,N_17164);
nor U17947 (N_17947,N_17108,N_17348);
or U17948 (N_17948,N_17430,N_17331);
and U17949 (N_17949,N_17462,N_17135);
nand U17950 (N_17950,N_17013,N_17114);
nand U17951 (N_17951,N_17121,N_17441);
or U17952 (N_17952,N_17416,N_17195);
and U17953 (N_17953,N_17434,N_17462);
xnor U17954 (N_17954,N_17122,N_17201);
or U17955 (N_17955,N_17199,N_17352);
and U17956 (N_17956,N_17015,N_17322);
nand U17957 (N_17957,N_17171,N_17362);
or U17958 (N_17958,N_17347,N_17486);
nor U17959 (N_17959,N_17316,N_17124);
nor U17960 (N_17960,N_17288,N_17065);
nand U17961 (N_17961,N_17345,N_17371);
xnor U17962 (N_17962,N_17472,N_17466);
nor U17963 (N_17963,N_17051,N_17196);
nor U17964 (N_17964,N_17183,N_17195);
xor U17965 (N_17965,N_17436,N_17004);
nor U17966 (N_17966,N_17075,N_17069);
nor U17967 (N_17967,N_17468,N_17374);
xor U17968 (N_17968,N_17242,N_17347);
xnor U17969 (N_17969,N_17218,N_17398);
xor U17970 (N_17970,N_17428,N_17286);
nand U17971 (N_17971,N_17301,N_17253);
nor U17972 (N_17972,N_17339,N_17205);
nor U17973 (N_17973,N_17171,N_17225);
or U17974 (N_17974,N_17397,N_17315);
or U17975 (N_17975,N_17455,N_17363);
and U17976 (N_17976,N_17335,N_17186);
and U17977 (N_17977,N_17467,N_17148);
nor U17978 (N_17978,N_17192,N_17237);
nand U17979 (N_17979,N_17108,N_17322);
nand U17980 (N_17980,N_17286,N_17161);
nand U17981 (N_17981,N_17180,N_17402);
and U17982 (N_17982,N_17381,N_17275);
or U17983 (N_17983,N_17398,N_17193);
and U17984 (N_17984,N_17435,N_17340);
nor U17985 (N_17985,N_17019,N_17382);
nand U17986 (N_17986,N_17013,N_17252);
nor U17987 (N_17987,N_17168,N_17082);
nand U17988 (N_17988,N_17281,N_17405);
nor U17989 (N_17989,N_17275,N_17335);
and U17990 (N_17990,N_17249,N_17279);
xnor U17991 (N_17991,N_17174,N_17038);
or U17992 (N_17992,N_17076,N_17205);
nor U17993 (N_17993,N_17198,N_17272);
nor U17994 (N_17994,N_17135,N_17312);
nand U17995 (N_17995,N_17304,N_17251);
nor U17996 (N_17996,N_17054,N_17476);
nand U17997 (N_17997,N_17082,N_17152);
or U17998 (N_17998,N_17386,N_17013);
nand U17999 (N_17999,N_17480,N_17061);
xnor U18000 (N_18000,N_17596,N_17810);
nor U18001 (N_18001,N_17687,N_17824);
nor U18002 (N_18002,N_17736,N_17768);
xnor U18003 (N_18003,N_17528,N_17922);
or U18004 (N_18004,N_17983,N_17599);
or U18005 (N_18005,N_17785,N_17849);
or U18006 (N_18006,N_17550,N_17733);
and U18007 (N_18007,N_17924,N_17981);
nor U18008 (N_18008,N_17717,N_17794);
nor U18009 (N_18009,N_17813,N_17882);
nor U18010 (N_18010,N_17720,N_17713);
and U18011 (N_18011,N_17923,N_17704);
nand U18012 (N_18012,N_17762,N_17759);
or U18013 (N_18013,N_17827,N_17769);
nand U18014 (N_18014,N_17513,N_17754);
nor U18015 (N_18015,N_17594,N_17626);
and U18016 (N_18016,N_17820,N_17862);
nor U18017 (N_18017,N_17531,N_17699);
xor U18018 (N_18018,N_17905,N_17995);
nor U18019 (N_18019,N_17669,N_17556);
nand U18020 (N_18020,N_17685,N_17823);
nand U18021 (N_18021,N_17635,N_17637);
nand U18022 (N_18022,N_17700,N_17741);
nand U18023 (N_18023,N_17865,N_17872);
nor U18024 (N_18024,N_17600,N_17544);
nor U18025 (N_18025,N_17642,N_17623);
or U18026 (N_18026,N_17707,N_17737);
or U18027 (N_18027,N_17653,N_17962);
or U18028 (N_18028,N_17634,N_17994);
xnor U18029 (N_18029,N_17886,N_17791);
nand U18030 (N_18030,N_17691,N_17927);
and U18031 (N_18031,N_17690,N_17801);
and U18032 (N_18032,N_17795,N_17848);
and U18033 (N_18033,N_17566,N_17870);
nand U18034 (N_18034,N_17775,N_17940);
nand U18035 (N_18035,N_17518,N_17842);
and U18036 (N_18036,N_17672,N_17765);
or U18037 (N_18037,N_17627,N_17752);
or U18038 (N_18038,N_17776,N_17818);
and U18039 (N_18039,N_17638,N_17658);
xor U18040 (N_18040,N_17773,N_17861);
and U18041 (N_18041,N_17763,N_17722);
or U18042 (N_18042,N_17656,N_17931);
nor U18043 (N_18043,N_17784,N_17705);
and U18044 (N_18044,N_17807,N_17540);
or U18045 (N_18045,N_17515,N_17547);
and U18046 (N_18046,N_17972,N_17702);
and U18047 (N_18047,N_17790,N_17788);
nand U18048 (N_18048,N_17977,N_17682);
nand U18049 (N_18049,N_17680,N_17667);
nand U18050 (N_18050,N_17555,N_17783);
and U18051 (N_18051,N_17947,N_17615);
nand U18052 (N_18052,N_17628,N_17595);
xnor U18053 (N_18053,N_17739,N_17884);
and U18054 (N_18054,N_17673,N_17616);
or U18055 (N_18055,N_17891,N_17529);
and U18056 (N_18056,N_17944,N_17975);
nand U18057 (N_18057,N_17636,N_17614);
or U18058 (N_18058,N_17799,N_17876);
nor U18059 (N_18059,N_17949,N_17689);
or U18060 (N_18060,N_17693,N_17878);
nand U18061 (N_18061,N_17959,N_17805);
nor U18062 (N_18062,N_17561,N_17661);
or U18063 (N_18063,N_17777,N_17694);
nor U18064 (N_18064,N_17665,N_17582);
nor U18065 (N_18065,N_17679,N_17514);
nand U18066 (N_18066,N_17917,N_17605);
and U18067 (N_18067,N_17979,N_17883);
nand U18068 (N_18068,N_17964,N_17557);
nand U18069 (N_18069,N_17649,N_17630);
or U18070 (N_18070,N_17527,N_17918);
nand U18071 (N_18071,N_17710,N_17703);
or U18072 (N_18072,N_17817,N_17538);
xnor U18073 (N_18073,N_17660,N_17552);
nor U18074 (N_18074,N_17512,N_17934);
or U18075 (N_18075,N_17684,N_17816);
nor U18076 (N_18076,N_17915,N_17901);
and U18077 (N_18077,N_17639,N_17879);
and U18078 (N_18078,N_17569,N_17778);
nand U18079 (N_18079,N_17906,N_17802);
and U18080 (N_18080,N_17937,N_17888);
nor U18081 (N_18081,N_17617,N_17952);
nand U18082 (N_18082,N_17902,N_17970);
nor U18083 (N_18083,N_17911,N_17648);
or U18084 (N_18084,N_17900,N_17604);
nor U18085 (N_18085,N_17757,N_17867);
nand U18086 (N_18086,N_17579,N_17892);
nor U18087 (N_18087,N_17852,N_17572);
and U18088 (N_18088,N_17747,N_17504);
nor U18089 (N_18089,N_17521,N_17697);
or U18090 (N_18090,N_17880,N_17958);
nand U18091 (N_18091,N_17945,N_17798);
or U18092 (N_18092,N_17898,N_17771);
or U18093 (N_18093,N_17522,N_17620);
nor U18094 (N_18094,N_17534,N_17991);
nand U18095 (N_18095,N_17845,N_17973);
or U18096 (N_18096,N_17965,N_17612);
and U18097 (N_18097,N_17812,N_17779);
or U18098 (N_18098,N_17701,N_17837);
or U18099 (N_18099,N_17930,N_17986);
nand U18100 (N_18100,N_17920,N_17908);
nor U18101 (N_18101,N_17575,N_17734);
nand U18102 (N_18102,N_17766,N_17863);
nand U18103 (N_18103,N_17897,N_17933);
nor U18104 (N_18104,N_17568,N_17619);
nand U18105 (N_18105,N_17858,N_17645);
and U18106 (N_18106,N_17834,N_17881);
and U18107 (N_18107,N_17588,N_17866);
xor U18108 (N_18108,N_17811,N_17729);
nor U18109 (N_18109,N_17893,N_17559);
nand U18110 (N_18110,N_17738,N_17692);
and U18111 (N_18111,N_17726,N_17592);
nor U18112 (N_18112,N_17815,N_17909);
and U18113 (N_18113,N_17618,N_17871);
and U18114 (N_18114,N_17647,N_17610);
and U18115 (N_18115,N_17963,N_17990);
nor U18116 (N_18116,N_17657,N_17758);
nand U18117 (N_18117,N_17681,N_17953);
or U18118 (N_18118,N_17553,N_17686);
nand U18119 (N_18119,N_17537,N_17974);
nand U18120 (N_18120,N_17868,N_17590);
nor U18121 (N_18121,N_17708,N_17706);
nand U18122 (N_18122,N_17804,N_17742);
nor U18123 (N_18123,N_17800,N_17532);
xnor U18124 (N_18124,N_17885,N_17519);
xor U18125 (N_18125,N_17786,N_17516);
and U18126 (N_18126,N_17980,N_17960);
nor U18127 (N_18127,N_17510,N_17652);
nand U18128 (N_18128,N_17764,N_17854);
nand U18129 (N_18129,N_17961,N_17601);
and U18130 (N_18130,N_17782,N_17535);
or U18131 (N_18131,N_17536,N_17997);
and U18132 (N_18132,N_17524,N_17928);
and U18133 (N_18133,N_17641,N_17695);
xnor U18134 (N_18134,N_17743,N_17814);
nor U18135 (N_18135,N_17567,N_17509);
and U18136 (N_18136,N_17573,N_17844);
nor U18137 (N_18137,N_17502,N_17929);
nor U18138 (N_18138,N_17608,N_17939);
xnor U18139 (N_18139,N_17853,N_17654);
nor U18140 (N_18140,N_17753,N_17602);
or U18141 (N_18141,N_17830,N_17840);
nor U18142 (N_18142,N_17621,N_17640);
nand U18143 (N_18143,N_17542,N_17677);
nor U18144 (N_18144,N_17749,N_17533);
and U18145 (N_18145,N_17584,N_17761);
nor U18146 (N_18146,N_17857,N_17951);
nand U18147 (N_18147,N_17921,N_17716);
nand U18148 (N_18148,N_17833,N_17526);
and U18149 (N_18149,N_17718,N_17789);
nand U18150 (N_18150,N_17819,N_17668);
nand U18151 (N_18151,N_17910,N_17916);
nor U18152 (N_18152,N_17731,N_17832);
or U18153 (N_18153,N_17676,N_17698);
xor U18154 (N_18154,N_17822,N_17523);
nor U18155 (N_18155,N_17606,N_17926);
xor U18156 (N_18156,N_17996,N_17808);
and U18157 (N_18157,N_17750,N_17622);
nor U18158 (N_18158,N_17554,N_17992);
xnor U18159 (N_18159,N_17803,N_17548);
and U18160 (N_18160,N_17683,N_17506);
nand U18161 (N_18161,N_17755,N_17770);
and U18162 (N_18162,N_17663,N_17580);
nor U18163 (N_18163,N_17745,N_17793);
xor U18164 (N_18164,N_17987,N_17511);
nand U18165 (N_18165,N_17941,N_17877);
nand U18166 (N_18166,N_17760,N_17586);
and U18167 (N_18167,N_17651,N_17631);
or U18168 (N_18168,N_17887,N_17525);
nor U18169 (N_18169,N_17501,N_17919);
nand U18170 (N_18170,N_17570,N_17792);
and U18171 (N_18171,N_17856,N_17577);
nand U18172 (N_18172,N_17890,N_17574);
xor U18173 (N_18173,N_17583,N_17869);
nor U18174 (N_18174,N_17632,N_17774);
xor U18175 (N_18175,N_17751,N_17925);
or U18176 (N_18176,N_17912,N_17625);
nand U18177 (N_18177,N_17831,N_17978);
nor U18178 (N_18178,N_17781,N_17855);
nor U18179 (N_18179,N_17549,N_17727);
nand U18180 (N_18180,N_17571,N_17563);
and U18181 (N_18181,N_17539,N_17675);
nand U18182 (N_18182,N_17957,N_17719);
or U18183 (N_18183,N_17936,N_17598);
nor U18184 (N_18184,N_17730,N_17581);
and U18185 (N_18185,N_17838,N_17825);
nor U18186 (N_18186,N_17907,N_17603);
and U18187 (N_18187,N_17889,N_17913);
nand U18188 (N_18188,N_17993,N_17659);
xnor U18189 (N_18189,N_17896,N_17688);
or U18190 (N_18190,N_17797,N_17725);
and U18191 (N_18191,N_17976,N_17895);
or U18192 (N_18192,N_17633,N_17674);
or U18193 (N_18193,N_17999,N_17841);
nor U18194 (N_18194,N_17740,N_17587);
xnor U18195 (N_18195,N_17748,N_17709);
or U18196 (N_18196,N_17806,N_17715);
and U18197 (N_18197,N_17984,N_17517);
or U18198 (N_18198,N_17988,N_17696);
or U18199 (N_18199,N_17543,N_17530);
and U18200 (N_18200,N_17578,N_17500);
nand U18201 (N_18201,N_17711,N_17950);
and U18202 (N_18202,N_17943,N_17966);
and U18203 (N_18203,N_17505,N_17732);
nand U18204 (N_18204,N_17597,N_17545);
and U18205 (N_18205,N_17956,N_17968);
or U18206 (N_18206,N_17851,N_17503);
and U18207 (N_18207,N_17666,N_17809);
nand U18208 (N_18208,N_17678,N_17564);
or U18209 (N_18209,N_17875,N_17836);
or U18210 (N_18210,N_17655,N_17756);
or U18211 (N_18211,N_17846,N_17507);
nor U18212 (N_18212,N_17723,N_17985);
xor U18213 (N_18213,N_17829,N_17938);
and U18214 (N_18214,N_17826,N_17611);
nand U18215 (N_18215,N_17998,N_17560);
xnor U18216 (N_18216,N_17873,N_17576);
and U18217 (N_18217,N_17558,N_17828);
xor U18218 (N_18218,N_17562,N_17894);
or U18219 (N_18219,N_17967,N_17864);
xnor U18220 (N_18220,N_17843,N_17948);
or U18221 (N_18221,N_17565,N_17714);
nor U18222 (N_18222,N_17767,N_17585);
nand U18223 (N_18223,N_17646,N_17914);
nor U18224 (N_18224,N_17821,N_17591);
or U18225 (N_18225,N_17932,N_17796);
nor U18226 (N_18226,N_17835,N_17903);
and U18227 (N_18227,N_17860,N_17746);
or U18228 (N_18228,N_17874,N_17551);
nor U18229 (N_18229,N_17607,N_17847);
nor U18230 (N_18230,N_17662,N_17643);
nand U18231 (N_18231,N_17969,N_17989);
nand U18232 (N_18232,N_17712,N_17850);
or U18233 (N_18233,N_17508,N_17609);
or U18234 (N_18234,N_17971,N_17721);
and U18235 (N_18235,N_17546,N_17589);
nand U18236 (N_18236,N_17671,N_17664);
or U18237 (N_18237,N_17946,N_17787);
and U18238 (N_18238,N_17744,N_17613);
nor U18239 (N_18239,N_17859,N_17670);
and U18240 (N_18240,N_17520,N_17772);
and U18241 (N_18241,N_17541,N_17629);
and U18242 (N_18242,N_17624,N_17593);
nor U18243 (N_18243,N_17650,N_17942);
nand U18244 (N_18244,N_17982,N_17935);
nor U18245 (N_18245,N_17724,N_17954);
and U18246 (N_18246,N_17728,N_17839);
and U18247 (N_18247,N_17735,N_17904);
nor U18248 (N_18248,N_17780,N_17899);
or U18249 (N_18249,N_17955,N_17644);
or U18250 (N_18250,N_17989,N_17914);
nor U18251 (N_18251,N_17898,N_17920);
or U18252 (N_18252,N_17659,N_17592);
or U18253 (N_18253,N_17889,N_17512);
xor U18254 (N_18254,N_17661,N_17906);
nand U18255 (N_18255,N_17613,N_17730);
or U18256 (N_18256,N_17946,N_17698);
nor U18257 (N_18257,N_17845,N_17992);
xor U18258 (N_18258,N_17671,N_17642);
nand U18259 (N_18259,N_17648,N_17888);
and U18260 (N_18260,N_17669,N_17512);
nor U18261 (N_18261,N_17583,N_17654);
or U18262 (N_18262,N_17864,N_17866);
nor U18263 (N_18263,N_17762,N_17544);
nor U18264 (N_18264,N_17755,N_17750);
and U18265 (N_18265,N_17604,N_17749);
and U18266 (N_18266,N_17868,N_17822);
or U18267 (N_18267,N_17968,N_17685);
nand U18268 (N_18268,N_17622,N_17903);
nand U18269 (N_18269,N_17753,N_17763);
or U18270 (N_18270,N_17990,N_17857);
nand U18271 (N_18271,N_17506,N_17714);
or U18272 (N_18272,N_17873,N_17807);
or U18273 (N_18273,N_17669,N_17807);
nor U18274 (N_18274,N_17667,N_17785);
nand U18275 (N_18275,N_17775,N_17615);
or U18276 (N_18276,N_17500,N_17894);
and U18277 (N_18277,N_17560,N_17867);
or U18278 (N_18278,N_17775,N_17559);
nand U18279 (N_18279,N_17979,N_17900);
xnor U18280 (N_18280,N_17683,N_17594);
or U18281 (N_18281,N_17663,N_17573);
xnor U18282 (N_18282,N_17757,N_17871);
and U18283 (N_18283,N_17600,N_17929);
or U18284 (N_18284,N_17906,N_17993);
nand U18285 (N_18285,N_17645,N_17568);
and U18286 (N_18286,N_17792,N_17883);
nand U18287 (N_18287,N_17989,N_17661);
or U18288 (N_18288,N_17720,N_17963);
nor U18289 (N_18289,N_17678,N_17907);
and U18290 (N_18290,N_17879,N_17813);
and U18291 (N_18291,N_17638,N_17600);
and U18292 (N_18292,N_17861,N_17971);
or U18293 (N_18293,N_17619,N_17518);
nand U18294 (N_18294,N_17607,N_17560);
and U18295 (N_18295,N_17741,N_17528);
nand U18296 (N_18296,N_17725,N_17759);
nand U18297 (N_18297,N_17884,N_17548);
nor U18298 (N_18298,N_17618,N_17704);
and U18299 (N_18299,N_17803,N_17629);
and U18300 (N_18300,N_17666,N_17760);
xor U18301 (N_18301,N_17792,N_17614);
nor U18302 (N_18302,N_17849,N_17593);
and U18303 (N_18303,N_17798,N_17553);
xnor U18304 (N_18304,N_17765,N_17536);
nand U18305 (N_18305,N_17885,N_17573);
and U18306 (N_18306,N_17695,N_17955);
nand U18307 (N_18307,N_17579,N_17992);
nor U18308 (N_18308,N_17516,N_17986);
xnor U18309 (N_18309,N_17641,N_17508);
nand U18310 (N_18310,N_17825,N_17860);
and U18311 (N_18311,N_17998,N_17602);
nor U18312 (N_18312,N_17859,N_17600);
xnor U18313 (N_18313,N_17667,N_17769);
nor U18314 (N_18314,N_17508,N_17709);
and U18315 (N_18315,N_17736,N_17852);
nand U18316 (N_18316,N_17577,N_17865);
nor U18317 (N_18317,N_17894,N_17529);
or U18318 (N_18318,N_17711,N_17677);
and U18319 (N_18319,N_17616,N_17523);
and U18320 (N_18320,N_17546,N_17815);
nand U18321 (N_18321,N_17766,N_17509);
or U18322 (N_18322,N_17785,N_17753);
xnor U18323 (N_18323,N_17850,N_17886);
nand U18324 (N_18324,N_17814,N_17921);
or U18325 (N_18325,N_17740,N_17981);
and U18326 (N_18326,N_17960,N_17873);
and U18327 (N_18327,N_17640,N_17588);
and U18328 (N_18328,N_17660,N_17675);
or U18329 (N_18329,N_17779,N_17923);
or U18330 (N_18330,N_17799,N_17776);
nand U18331 (N_18331,N_17736,N_17554);
nor U18332 (N_18332,N_17742,N_17912);
or U18333 (N_18333,N_17992,N_17908);
nor U18334 (N_18334,N_17876,N_17712);
nor U18335 (N_18335,N_17630,N_17887);
or U18336 (N_18336,N_17503,N_17578);
nor U18337 (N_18337,N_17603,N_17996);
nor U18338 (N_18338,N_17995,N_17534);
and U18339 (N_18339,N_17575,N_17663);
nand U18340 (N_18340,N_17540,N_17701);
or U18341 (N_18341,N_17597,N_17972);
and U18342 (N_18342,N_17908,N_17871);
and U18343 (N_18343,N_17601,N_17714);
or U18344 (N_18344,N_17535,N_17790);
and U18345 (N_18345,N_17610,N_17884);
or U18346 (N_18346,N_17762,N_17735);
xnor U18347 (N_18347,N_17871,N_17705);
and U18348 (N_18348,N_17687,N_17711);
nor U18349 (N_18349,N_17842,N_17759);
nor U18350 (N_18350,N_17913,N_17944);
nor U18351 (N_18351,N_17852,N_17851);
and U18352 (N_18352,N_17964,N_17739);
or U18353 (N_18353,N_17762,N_17707);
nand U18354 (N_18354,N_17593,N_17763);
nor U18355 (N_18355,N_17501,N_17524);
and U18356 (N_18356,N_17653,N_17672);
nor U18357 (N_18357,N_17615,N_17743);
nand U18358 (N_18358,N_17958,N_17948);
or U18359 (N_18359,N_17990,N_17900);
or U18360 (N_18360,N_17908,N_17568);
nand U18361 (N_18361,N_17998,N_17514);
or U18362 (N_18362,N_17682,N_17945);
xor U18363 (N_18363,N_17617,N_17982);
or U18364 (N_18364,N_17800,N_17662);
or U18365 (N_18365,N_17764,N_17713);
nand U18366 (N_18366,N_17947,N_17661);
nand U18367 (N_18367,N_17856,N_17936);
and U18368 (N_18368,N_17887,N_17551);
nand U18369 (N_18369,N_17521,N_17584);
nand U18370 (N_18370,N_17681,N_17647);
nor U18371 (N_18371,N_17579,N_17850);
xor U18372 (N_18372,N_17775,N_17742);
or U18373 (N_18373,N_17889,N_17684);
and U18374 (N_18374,N_17685,N_17802);
xor U18375 (N_18375,N_17656,N_17722);
or U18376 (N_18376,N_17875,N_17844);
or U18377 (N_18377,N_17862,N_17786);
nand U18378 (N_18378,N_17832,N_17988);
and U18379 (N_18379,N_17797,N_17806);
and U18380 (N_18380,N_17647,N_17508);
xor U18381 (N_18381,N_17821,N_17639);
nand U18382 (N_18382,N_17503,N_17720);
or U18383 (N_18383,N_17941,N_17772);
nand U18384 (N_18384,N_17733,N_17671);
or U18385 (N_18385,N_17531,N_17500);
xnor U18386 (N_18386,N_17673,N_17580);
nor U18387 (N_18387,N_17883,N_17815);
and U18388 (N_18388,N_17719,N_17775);
nand U18389 (N_18389,N_17974,N_17796);
and U18390 (N_18390,N_17692,N_17584);
nor U18391 (N_18391,N_17553,N_17848);
and U18392 (N_18392,N_17688,N_17555);
nand U18393 (N_18393,N_17582,N_17972);
nor U18394 (N_18394,N_17807,N_17751);
nand U18395 (N_18395,N_17936,N_17986);
nand U18396 (N_18396,N_17887,N_17712);
nand U18397 (N_18397,N_17569,N_17534);
nand U18398 (N_18398,N_17719,N_17998);
nand U18399 (N_18399,N_17946,N_17565);
nor U18400 (N_18400,N_17696,N_17503);
nand U18401 (N_18401,N_17648,N_17594);
nand U18402 (N_18402,N_17588,N_17927);
xnor U18403 (N_18403,N_17609,N_17606);
nand U18404 (N_18404,N_17821,N_17817);
nand U18405 (N_18405,N_17796,N_17651);
nor U18406 (N_18406,N_17897,N_17542);
nor U18407 (N_18407,N_17500,N_17692);
xor U18408 (N_18408,N_17574,N_17792);
xnor U18409 (N_18409,N_17820,N_17692);
or U18410 (N_18410,N_17682,N_17866);
nor U18411 (N_18411,N_17535,N_17824);
nor U18412 (N_18412,N_17568,N_17823);
nor U18413 (N_18413,N_17568,N_17829);
or U18414 (N_18414,N_17830,N_17846);
nand U18415 (N_18415,N_17681,N_17704);
nand U18416 (N_18416,N_17778,N_17721);
or U18417 (N_18417,N_17793,N_17699);
nor U18418 (N_18418,N_17892,N_17541);
and U18419 (N_18419,N_17745,N_17652);
nor U18420 (N_18420,N_17835,N_17921);
or U18421 (N_18421,N_17553,N_17703);
nand U18422 (N_18422,N_17820,N_17656);
and U18423 (N_18423,N_17729,N_17563);
nand U18424 (N_18424,N_17853,N_17967);
nor U18425 (N_18425,N_17580,N_17671);
nor U18426 (N_18426,N_17713,N_17590);
nand U18427 (N_18427,N_17833,N_17656);
and U18428 (N_18428,N_17601,N_17570);
nand U18429 (N_18429,N_17677,N_17636);
nand U18430 (N_18430,N_17873,N_17842);
xnor U18431 (N_18431,N_17913,N_17878);
nand U18432 (N_18432,N_17770,N_17662);
nor U18433 (N_18433,N_17851,N_17548);
nand U18434 (N_18434,N_17661,N_17998);
nand U18435 (N_18435,N_17697,N_17604);
xor U18436 (N_18436,N_17823,N_17936);
nand U18437 (N_18437,N_17841,N_17505);
and U18438 (N_18438,N_17526,N_17748);
or U18439 (N_18439,N_17746,N_17782);
nor U18440 (N_18440,N_17512,N_17856);
nor U18441 (N_18441,N_17871,N_17640);
nor U18442 (N_18442,N_17895,N_17644);
xnor U18443 (N_18443,N_17820,N_17699);
and U18444 (N_18444,N_17561,N_17604);
and U18445 (N_18445,N_17741,N_17584);
and U18446 (N_18446,N_17756,N_17728);
nand U18447 (N_18447,N_17951,N_17836);
and U18448 (N_18448,N_17753,N_17774);
or U18449 (N_18449,N_17760,N_17689);
and U18450 (N_18450,N_17575,N_17944);
xor U18451 (N_18451,N_17818,N_17972);
nand U18452 (N_18452,N_17674,N_17803);
or U18453 (N_18453,N_17917,N_17830);
or U18454 (N_18454,N_17815,N_17764);
and U18455 (N_18455,N_17880,N_17691);
and U18456 (N_18456,N_17859,N_17653);
and U18457 (N_18457,N_17933,N_17686);
and U18458 (N_18458,N_17811,N_17651);
or U18459 (N_18459,N_17812,N_17882);
and U18460 (N_18460,N_17810,N_17787);
xor U18461 (N_18461,N_17910,N_17579);
and U18462 (N_18462,N_17744,N_17632);
nand U18463 (N_18463,N_17798,N_17875);
nand U18464 (N_18464,N_17890,N_17677);
nand U18465 (N_18465,N_17857,N_17508);
and U18466 (N_18466,N_17941,N_17917);
or U18467 (N_18467,N_17503,N_17743);
nor U18468 (N_18468,N_17768,N_17663);
or U18469 (N_18469,N_17726,N_17682);
nor U18470 (N_18470,N_17774,N_17997);
nand U18471 (N_18471,N_17792,N_17973);
or U18472 (N_18472,N_17794,N_17708);
nand U18473 (N_18473,N_17895,N_17882);
nor U18474 (N_18474,N_17850,N_17748);
nor U18475 (N_18475,N_17679,N_17841);
or U18476 (N_18476,N_17771,N_17882);
or U18477 (N_18477,N_17741,N_17600);
xor U18478 (N_18478,N_17796,N_17510);
xor U18479 (N_18479,N_17764,N_17662);
nand U18480 (N_18480,N_17722,N_17623);
or U18481 (N_18481,N_17976,N_17560);
nand U18482 (N_18482,N_17635,N_17629);
and U18483 (N_18483,N_17584,N_17528);
nor U18484 (N_18484,N_17929,N_17824);
nor U18485 (N_18485,N_17517,N_17660);
xor U18486 (N_18486,N_17513,N_17941);
or U18487 (N_18487,N_17885,N_17714);
nand U18488 (N_18488,N_17945,N_17789);
and U18489 (N_18489,N_17967,N_17608);
and U18490 (N_18490,N_17581,N_17923);
nand U18491 (N_18491,N_17791,N_17982);
nand U18492 (N_18492,N_17542,N_17768);
xnor U18493 (N_18493,N_17708,N_17628);
and U18494 (N_18494,N_17953,N_17878);
nor U18495 (N_18495,N_17506,N_17644);
or U18496 (N_18496,N_17621,N_17604);
nand U18497 (N_18497,N_17899,N_17800);
nor U18498 (N_18498,N_17839,N_17971);
and U18499 (N_18499,N_17943,N_17791);
and U18500 (N_18500,N_18457,N_18478);
nor U18501 (N_18501,N_18169,N_18105);
xor U18502 (N_18502,N_18438,N_18026);
xor U18503 (N_18503,N_18160,N_18029);
xor U18504 (N_18504,N_18393,N_18408);
nor U18505 (N_18505,N_18031,N_18234);
or U18506 (N_18506,N_18313,N_18086);
and U18507 (N_18507,N_18197,N_18278);
nand U18508 (N_18508,N_18145,N_18286);
or U18509 (N_18509,N_18180,N_18335);
and U18510 (N_18510,N_18125,N_18304);
or U18511 (N_18511,N_18370,N_18373);
and U18512 (N_18512,N_18298,N_18441);
nand U18513 (N_18513,N_18281,N_18415);
and U18514 (N_18514,N_18480,N_18171);
nand U18515 (N_18515,N_18109,N_18052);
or U18516 (N_18516,N_18194,N_18091);
or U18517 (N_18517,N_18132,N_18096);
nand U18518 (N_18518,N_18292,N_18252);
or U18519 (N_18519,N_18092,N_18230);
or U18520 (N_18520,N_18233,N_18210);
or U18521 (N_18521,N_18128,N_18030);
nand U18522 (N_18522,N_18253,N_18306);
xnor U18523 (N_18523,N_18452,N_18100);
or U18524 (N_18524,N_18003,N_18463);
or U18525 (N_18525,N_18356,N_18085);
and U18526 (N_18526,N_18146,N_18187);
and U18527 (N_18527,N_18449,N_18069);
and U18528 (N_18528,N_18458,N_18349);
or U18529 (N_18529,N_18191,N_18468);
xnor U18530 (N_18530,N_18222,N_18073);
and U18531 (N_18531,N_18017,N_18106);
nand U18532 (N_18532,N_18305,N_18414);
nand U18533 (N_18533,N_18032,N_18243);
nand U18534 (N_18534,N_18061,N_18063);
nor U18535 (N_18535,N_18070,N_18156);
nand U18536 (N_18536,N_18176,N_18422);
nor U18537 (N_18537,N_18260,N_18406);
nand U18538 (N_18538,N_18440,N_18251);
nand U18539 (N_18539,N_18483,N_18444);
and U18540 (N_18540,N_18228,N_18258);
and U18541 (N_18541,N_18332,N_18144);
or U18542 (N_18542,N_18172,N_18110);
nand U18543 (N_18543,N_18072,N_18163);
nand U18544 (N_18544,N_18377,N_18418);
or U18545 (N_18545,N_18235,N_18357);
nor U18546 (N_18546,N_18192,N_18365);
or U18547 (N_18547,N_18376,N_18208);
nor U18548 (N_18548,N_18445,N_18189);
or U18549 (N_18549,N_18333,N_18093);
and U18550 (N_18550,N_18436,N_18329);
or U18551 (N_18551,N_18198,N_18301);
nor U18552 (N_18552,N_18257,N_18202);
and U18553 (N_18553,N_18394,N_18159);
nor U18554 (N_18554,N_18124,N_18450);
xnor U18555 (N_18555,N_18469,N_18212);
and U18556 (N_18556,N_18007,N_18255);
xor U18557 (N_18557,N_18261,N_18411);
nor U18558 (N_18558,N_18337,N_18479);
nand U18559 (N_18559,N_18225,N_18114);
nor U18560 (N_18560,N_18379,N_18434);
and U18561 (N_18561,N_18204,N_18446);
nor U18562 (N_18562,N_18161,N_18164);
or U18563 (N_18563,N_18283,N_18390);
nand U18564 (N_18564,N_18244,N_18407);
nor U18565 (N_18565,N_18268,N_18201);
nor U18566 (N_18566,N_18001,N_18389);
nand U18567 (N_18567,N_18167,N_18274);
nand U18568 (N_18568,N_18203,N_18447);
xnor U18569 (N_18569,N_18477,N_18020);
nor U18570 (N_18570,N_18350,N_18325);
and U18571 (N_18571,N_18015,N_18012);
or U18572 (N_18572,N_18419,N_18060);
nand U18573 (N_18573,N_18123,N_18439);
xor U18574 (N_18574,N_18303,N_18428);
and U18575 (N_18575,N_18249,N_18471);
nor U18576 (N_18576,N_18147,N_18402);
and U18577 (N_18577,N_18143,N_18104);
and U18578 (N_18578,N_18018,N_18388);
nand U18579 (N_18579,N_18416,N_18182);
xor U18580 (N_18580,N_18273,N_18443);
nor U18581 (N_18581,N_18068,N_18089);
and U18582 (N_18582,N_18359,N_18098);
nor U18583 (N_18583,N_18195,N_18276);
or U18584 (N_18584,N_18067,N_18316);
nor U18585 (N_18585,N_18046,N_18364);
nor U18586 (N_18586,N_18430,N_18429);
nor U18587 (N_18587,N_18213,N_18417);
nor U18588 (N_18588,N_18177,N_18473);
and U18589 (N_18589,N_18088,N_18395);
nor U18590 (N_18590,N_18295,N_18102);
nand U18591 (N_18591,N_18053,N_18118);
nand U18592 (N_18592,N_18499,N_18300);
nand U18593 (N_18593,N_18453,N_18385);
xor U18594 (N_18594,N_18308,N_18340);
nand U18595 (N_18595,N_18410,N_18165);
and U18596 (N_18596,N_18004,N_18232);
and U18597 (N_18597,N_18490,N_18310);
nand U18598 (N_18598,N_18384,N_18279);
nand U18599 (N_18599,N_18022,N_18448);
or U18600 (N_18600,N_18263,N_18339);
or U18601 (N_18601,N_18207,N_18327);
nand U18602 (N_18602,N_18248,N_18162);
nor U18603 (N_18603,N_18178,N_18285);
xor U18604 (N_18604,N_18374,N_18078);
nor U18605 (N_18605,N_18014,N_18497);
nor U18606 (N_18606,N_18367,N_18013);
xnor U18607 (N_18607,N_18223,N_18269);
nand U18608 (N_18608,N_18037,N_18183);
and U18609 (N_18609,N_18034,N_18076);
and U18610 (N_18610,N_18351,N_18371);
and U18611 (N_18611,N_18050,N_18464);
and U18612 (N_18612,N_18000,N_18116);
or U18613 (N_18613,N_18433,N_18461);
or U18614 (N_18614,N_18215,N_18141);
nor U18615 (N_18615,N_18318,N_18391);
and U18616 (N_18616,N_18309,N_18271);
nand U18617 (N_18617,N_18056,N_18467);
nand U18618 (N_18618,N_18264,N_18019);
and U18619 (N_18619,N_18470,N_18082);
nor U18620 (N_18620,N_18342,N_18107);
nand U18621 (N_18621,N_18314,N_18080);
and U18622 (N_18622,N_18361,N_18129);
nand U18623 (N_18623,N_18140,N_18299);
and U18624 (N_18624,N_18220,N_18287);
or U18625 (N_18625,N_18035,N_18288);
or U18626 (N_18626,N_18154,N_18319);
and U18627 (N_18627,N_18113,N_18262);
and U18628 (N_18628,N_18038,N_18117);
or U18629 (N_18629,N_18239,N_18135);
nor U18630 (N_18630,N_18087,N_18343);
or U18631 (N_18631,N_18231,N_18083);
nor U18632 (N_18632,N_18033,N_18168);
nand U18633 (N_18633,N_18250,N_18023);
and U18634 (N_18634,N_18101,N_18294);
nand U18635 (N_18635,N_18055,N_18016);
xnor U18636 (N_18636,N_18041,N_18297);
or U18637 (N_18637,N_18427,N_18413);
and U18638 (N_18638,N_18491,N_18284);
or U18639 (N_18639,N_18226,N_18188);
and U18640 (N_18640,N_18227,N_18133);
or U18641 (N_18641,N_18148,N_18238);
xnor U18642 (N_18642,N_18175,N_18472);
or U18643 (N_18643,N_18360,N_18420);
nand U18644 (N_18644,N_18272,N_18366);
and U18645 (N_18645,N_18307,N_18302);
nor U18646 (N_18646,N_18328,N_18174);
nand U18647 (N_18647,N_18435,N_18216);
nor U18648 (N_18648,N_18081,N_18206);
and U18649 (N_18649,N_18494,N_18462);
nor U18650 (N_18650,N_18256,N_18369);
xor U18651 (N_18651,N_18331,N_18387);
or U18652 (N_18652,N_18153,N_18010);
and U18653 (N_18653,N_18240,N_18242);
or U18654 (N_18654,N_18465,N_18084);
nor U18655 (N_18655,N_18496,N_18059);
xnor U18656 (N_18656,N_18437,N_18064);
nand U18657 (N_18657,N_18345,N_18150);
and U18658 (N_18658,N_18138,N_18094);
or U18659 (N_18659,N_18399,N_18259);
or U18660 (N_18660,N_18265,N_18071);
nand U18661 (N_18661,N_18336,N_18451);
nor U18662 (N_18662,N_18179,N_18484);
and U18663 (N_18663,N_18121,N_18044);
and U18664 (N_18664,N_18205,N_18122);
or U18665 (N_18665,N_18266,N_18454);
xnor U18666 (N_18666,N_18456,N_18347);
nor U18667 (N_18667,N_18152,N_18344);
and U18668 (N_18668,N_18466,N_18139);
nand U18669 (N_18669,N_18200,N_18186);
nor U18670 (N_18670,N_18011,N_18119);
nor U18671 (N_18671,N_18224,N_18024);
nand U18672 (N_18672,N_18049,N_18120);
or U18673 (N_18673,N_18323,N_18282);
nor U18674 (N_18674,N_18403,N_18131);
nand U18675 (N_18675,N_18066,N_18425);
and U18676 (N_18676,N_18311,N_18352);
nor U18677 (N_18677,N_18039,N_18383);
nand U18678 (N_18678,N_18396,N_18363);
nor U18679 (N_18679,N_18378,N_18021);
nand U18680 (N_18680,N_18199,N_18398);
xor U18681 (N_18681,N_18341,N_18289);
and U18682 (N_18682,N_18209,N_18047);
nand U18683 (N_18683,N_18404,N_18170);
or U18684 (N_18684,N_18112,N_18397);
nor U18685 (N_18685,N_18334,N_18320);
nand U18686 (N_18686,N_18291,N_18412);
nor U18687 (N_18687,N_18002,N_18079);
or U18688 (N_18688,N_18405,N_18108);
xnor U18689 (N_18689,N_18158,N_18214);
and U18690 (N_18690,N_18442,N_18057);
nand U18691 (N_18691,N_18027,N_18090);
and U18692 (N_18692,N_18151,N_18275);
and U18693 (N_18693,N_18043,N_18317);
and U18694 (N_18694,N_18368,N_18221);
or U18695 (N_18695,N_18293,N_18254);
and U18696 (N_18696,N_18184,N_18267);
and U18697 (N_18697,N_18381,N_18115);
nor U18698 (N_18698,N_18103,N_18423);
nor U18699 (N_18699,N_18028,N_18246);
and U18700 (N_18700,N_18354,N_18111);
nand U18701 (N_18701,N_18355,N_18040);
nand U18702 (N_18702,N_18489,N_18421);
and U18703 (N_18703,N_18353,N_18326);
or U18704 (N_18704,N_18062,N_18190);
nand U18705 (N_18705,N_18097,N_18136);
and U18706 (N_18706,N_18474,N_18481);
and U18707 (N_18707,N_18095,N_18280);
and U18708 (N_18708,N_18487,N_18426);
nand U18709 (N_18709,N_18338,N_18045);
or U18710 (N_18710,N_18245,N_18382);
nor U18711 (N_18711,N_18130,N_18358);
nor U18712 (N_18712,N_18431,N_18372);
nand U18713 (N_18713,N_18127,N_18492);
and U18714 (N_18714,N_18482,N_18142);
nor U18715 (N_18715,N_18185,N_18270);
nor U18716 (N_18716,N_18241,N_18362);
and U18717 (N_18717,N_18005,N_18346);
and U18718 (N_18718,N_18048,N_18476);
and U18719 (N_18719,N_18065,N_18401);
nand U18720 (N_18720,N_18058,N_18042);
nor U18721 (N_18721,N_18409,N_18424);
nor U18722 (N_18722,N_18149,N_18217);
nand U18723 (N_18723,N_18460,N_18488);
nor U18724 (N_18724,N_18277,N_18455);
nand U18725 (N_18725,N_18025,N_18006);
or U18726 (N_18726,N_18051,N_18485);
nor U18727 (N_18727,N_18036,N_18074);
or U18728 (N_18728,N_18375,N_18322);
nand U18729 (N_18729,N_18475,N_18400);
and U18730 (N_18730,N_18173,N_18181);
or U18731 (N_18731,N_18008,N_18495);
and U18732 (N_18732,N_18312,N_18196);
nand U18733 (N_18733,N_18137,N_18321);
nand U18734 (N_18734,N_18126,N_18330);
and U18735 (N_18735,N_18380,N_18229);
nor U18736 (N_18736,N_18054,N_18236);
nor U18737 (N_18737,N_18290,N_18493);
nand U18738 (N_18738,N_18134,N_18392);
and U18739 (N_18739,N_18237,N_18157);
and U18740 (N_18740,N_18193,N_18218);
and U18741 (N_18741,N_18324,N_18486);
nor U18742 (N_18742,N_18315,N_18498);
nand U18743 (N_18743,N_18432,N_18247);
and U18744 (N_18744,N_18099,N_18296);
or U18745 (N_18745,N_18386,N_18077);
and U18746 (N_18746,N_18166,N_18459);
nor U18747 (N_18747,N_18219,N_18075);
and U18748 (N_18748,N_18211,N_18009);
and U18749 (N_18749,N_18348,N_18155);
xor U18750 (N_18750,N_18260,N_18063);
and U18751 (N_18751,N_18036,N_18477);
and U18752 (N_18752,N_18068,N_18440);
and U18753 (N_18753,N_18344,N_18057);
nor U18754 (N_18754,N_18269,N_18199);
nor U18755 (N_18755,N_18150,N_18335);
or U18756 (N_18756,N_18229,N_18043);
and U18757 (N_18757,N_18226,N_18057);
nand U18758 (N_18758,N_18474,N_18380);
or U18759 (N_18759,N_18457,N_18448);
or U18760 (N_18760,N_18224,N_18201);
and U18761 (N_18761,N_18222,N_18490);
or U18762 (N_18762,N_18046,N_18223);
and U18763 (N_18763,N_18467,N_18117);
nor U18764 (N_18764,N_18019,N_18152);
nand U18765 (N_18765,N_18475,N_18148);
xnor U18766 (N_18766,N_18233,N_18006);
nand U18767 (N_18767,N_18328,N_18140);
or U18768 (N_18768,N_18341,N_18397);
and U18769 (N_18769,N_18031,N_18211);
nand U18770 (N_18770,N_18280,N_18498);
or U18771 (N_18771,N_18404,N_18371);
nor U18772 (N_18772,N_18299,N_18450);
nor U18773 (N_18773,N_18204,N_18020);
nor U18774 (N_18774,N_18207,N_18185);
and U18775 (N_18775,N_18477,N_18201);
nor U18776 (N_18776,N_18154,N_18288);
or U18777 (N_18777,N_18052,N_18469);
and U18778 (N_18778,N_18390,N_18466);
nand U18779 (N_18779,N_18350,N_18460);
nand U18780 (N_18780,N_18032,N_18175);
or U18781 (N_18781,N_18429,N_18034);
nor U18782 (N_18782,N_18093,N_18043);
nor U18783 (N_18783,N_18249,N_18346);
nor U18784 (N_18784,N_18196,N_18228);
nor U18785 (N_18785,N_18144,N_18082);
or U18786 (N_18786,N_18230,N_18410);
or U18787 (N_18787,N_18309,N_18175);
and U18788 (N_18788,N_18255,N_18234);
or U18789 (N_18789,N_18150,N_18368);
xor U18790 (N_18790,N_18351,N_18428);
and U18791 (N_18791,N_18308,N_18065);
or U18792 (N_18792,N_18317,N_18190);
nand U18793 (N_18793,N_18470,N_18144);
and U18794 (N_18794,N_18273,N_18152);
nand U18795 (N_18795,N_18186,N_18044);
nand U18796 (N_18796,N_18342,N_18003);
and U18797 (N_18797,N_18062,N_18347);
or U18798 (N_18798,N_18175,N_18194);
or U18799 (N_18799,N_18406,N_18311);
nand U18800 (N_18800,N_18212,N_18126);
nand U18801 (N_18801,N_18116,N_18442);
nand U18802 (N_18802,N_18028,N_18041);
and U18803 (N_18803,N_18132,N_18351);
and U18804 (N_18804,N_18211,N_18242);
nor U18805 (N_18805,N_18450,N_18109);
and U18806 (N_18806,N_18324,N_18293);
nand U18807 (N_18807,N_18100,N_18206);
or U18808 (N_18808,N_18499,N_18228);
nor U18809 (N_18809,N_18034,N_18221);
or U18810 (N_18810,N_18355,N_18493);
and U18811 (N_18811,N_18400,N_18496);
and U18812 (N_18812,N_18151,N_18408);
nor U18813 (N_18813,N_18005,N_18366);
xnor U18814 (N_18814,N_18177,N_18116);
nand U18815 (N_18815,N_18050,N_18494);
xor U18816 (N_18816,N_18168,N_18141);
xor U18817 (N_18817,N_18371,N_18296);
or U18818 (N_18818,N_18380,N_18108);
nand U18819 (N_18819,N_18229,N_18193);
nand U18820 (N_18820,N_18110,N_18441);
and U18821 (N_18821,N_18125,N_18109);
nand U18822 (N_18822,N_18217,N_18082);
or U18823 (N_18823,N_18037,N_18443);
nor U18824 (N_18824,N_18350,N_18324);
and U18825 (N_18825,N_18123,N_18250);
and U18826 (N_18826,N_18422,N_18288);
xnor U18827 (N_18827,N_18326,N_18271);
and U18828 (N_18828,N_18072,N_18084);
nor U18829 (N_18829,N_18288,N_18374);
xnor U18830 (N_18830,N_18289,N_18131);
or U18831 (N_18831,N_18484,N_18250);
xnor U18832 (N_18832,N_18194,N_18465);
nand U18833 (N_18833,N_18373,N_18131);
or U18834 (N_18834,N_18289,N_18236);
and U18835 (N_18835,N_18304,N_18077);
nand U18836 (N_18836,N_18007,N_18318);
nor U18837 (N_18837,N_18010,N_18121);
nor U18838 (N_18838,N_18423,N_18447);
nor U18839 (N_18839,N_18329,N_18111);
xnor U18840 (N_18840,N_18227,N_18420);
nand U18841 (N_18841,N_18346,N_18411);
nor U18842 (N_18842,N_18435,N_18200);
nand U18843 (N_18843,N_18308,N_18474);
or U18844 (N_18844,N_18042,N_18341);
and U18845 (N_18845,N_18493,N_18397);
nor U18846 (N_18846,N_18348,N_18402);
and U18847 (N_18847,N_18366,N_18171);
nor U18848 (N_18848,N_18202,N_18272);
nor U18849 (N_18849,N_18291,N_18108);
or U18850 (N_18850,N_18335,N_18268);
nand U18851 (N_18851,N_18007,N_18053);
nor U18852 (N_18852,N_18474,N_18014);
or U18853 (N_18853,N_18027,N_18254);
nand U18854 (N_18854,N_18324,N_18095);
xor U18855 (N_18855,N_18267,N_18441);
or U18856 (N_18856,N_18469,N_18168);
or U18857 (N_18857,N_18482,N_18475);
nand U18858 (N_18858,N_18192,N_18429);
nor U18859 (N_18859,N_18249,N_18468);
nor U18860 (N_18860,N_18119,N_18374);
and U18861 (N_18861,N_18211,N_18203);
nor U18862 (N_18862,N_18331,N_18437);
and U18863 (N_18863,N_18186,N_18173);
nand U18864 (N_18864,N_18253,N_18190);
or U18865 (N_18865,N_18258,N_18170);
xor U18866 (N_18866,N_18412,N_18014);
and U18867 (N_18867,N_18449,N_18309);
nand U18868 (N_18868,N_18455,N_18008);
nor U18869 (N_18869,N_18078,N_18409);
nand U18870 (N_18870,N_18084,N_18013);
and U18871 (N_18871,N_18161,N_18018);
nand U18872 (N_18872,N_18337,N_18116);
and U18873 (N_18873,N_18483,N_18174);
or U18874 (N_18874,N_18019,N_18298);
nand U18875 (N_18875,N_18029,N_18279);
nor U18876 (N_18876,N_18442,N_18105);
nor U18877 (N_18877,N_18406,N_18468);
or U18878 (N_18878,N_18287,N_18094);
nand U18879 (N_18879,N_18084,N_18111);
xor U18880 (N_18880,N_18024,N_18474);
nand U18881 (N_18881,N_18367,N_18297);
or U18882 (N_18882,N_18031,N_18357);
xor U18883 (N_18883,N_18206,N_18174);
nand U18884 (N_18884,N_18432,N_18391);
or U18885 (N_18885,N_18330,N_18136);
nand U18886 (N_18886,N_18094,N_18303);
nand U18887 (N_18887,N_18182,N_18429);
xnor U18888 (N_18888,N_18018,N_18240);
and U18889 (N_18889,N_18220,N_18312);
and U18890 (N_18890,N_18132,N_18150);
nor U18891 (N_18891,N_18142,N_18059);
nor U18892 (N_18892,N_18266,N_18203);
nor U18893 (N_18893,N_18473,N_18269);
and U18894 (N_18894,N_18017,N_18480);
nand U18895 (N_18895,N_18011,N_18434);
or U18896 (N_18896,N_18473,N_18287);
xnor U18897 (N_18897,N_18444,N_18400);
nor U18898 (N_18898,N_18130,N_18233);
or U18899 (N_18899,N_18416,N_18201);
nor U18900 (N_18900,N_18259,N_18449);
nor U18901 (N_18901,N_18400,N_18394);
nor U18902 (N_18902,N_18207,N_18402);
nand U18903 (N_18903,N_18404,N_18053);
and U18904 (N_18904,N_18341,N_18339);
and U18905 (N_18905,N_18132,N_18008);
or U18906 (N_18906,N_18196,N_18199);
nor U18907 (N_18907,N_18483,N_18121);
or U18908 (N_18908,N_18037,N_18475);
and U18909 (N_18909,N_18208,N_18308);
nor U18910 (N_18910,N_18152,N_18106);
nand U18911 (N_18911,N_18082,N_18131);
or U18912 (N_18912,N_18015,N_18292);
nand U18913 (N_18913,N_18258,N_18479);
and U18914 (N_18914,N_18169,N_18255);
nand U18915 (N_18915,N_18144,N_18093);
or U18916 (N_18916,N_18084,N_18147);
nand U18917 (N_18917,N_18008,N_18141);
xor U18918 (N_18918,N_18140,N_18211);
or U18919 (N_18919,N_18206,N_18331);
and U18920 (N_18920,N_18018,N_18404);
xnor U18921 (N_18921,N_18128,N_18141);
or U18922 (N_18922,N_18316,N_18023);
nor U18923 (N_18923,N_18323,N_18135);
nor U18924 (N_18924,N_18457,N_18480);
and U18925 (N_18925,N_18429,N_18210);
or U18926 (N_18926,N_18454,N_18396);
nand U18927 (N_18927,N_18007,N_18261);
or U18928 (N_18928,N_18459,N_18357);
or U18929 (N_18929,N_18083,N_18094);
and U18930 (N_18930,N_18112,N_18240);
nor U18931 (N_18931,N_18395,N_18151);
and U18932 (N_18932,N_18118,N_18084);
and U18933 (N_18933,N_18075,N_18216);
or U18934 (N_18934,N_18188,N_18075);
xnor U18935 (N_18935,N_18402,N_18268);
xnor U18936 (N_18936,N_18277,N_18173);
and U18937 (N_18937,N_18485,N_18003);
or U18938 (N_18938,N_18276,N_18370);
nand U18939 (N_18939,N_18411,N_18300);
nand U18940 (N_18940,N_18095,N_18420);
xor U18941 (N_18941,N_18448,N_18149);
nor U18942 (N_18942,N_18474,N_18253);
or U18943 (N_18943,N_18198,N_18328);
and U18944 (N_18944,N_18340,N_18334);
nor U18945 (N_18945,N_18391,N_18282);
nand U18946 (N_18946,N_18363,N_18133);
and U18947 (N_18947,N_18439,N_18001);
and U18948 (N_18948,N_18489,N_18204);
nor U18949 (N_18949,N_18468,N_18357);
and U18950 (N_18950,N_18063,N_18004);
or U18951 (N_18951,N_18331,N_18235);
nand U18952 (N_18952,N_18473,N_18404);
nor U18953 (N_18953,N_18366,N_18037);
nand U18954 (N_18954,N_18156,N_18263);
or U18955 (N_18955,N_18251,N_18069);
nor U18956 (N_18956,N_18480,N_18198);
and U18957 (N_18957,N_18122,N_18223);
nor U18958 (N_18958,N_18275,N_18203);
nor U18959 (N_18959,N_18187,N_18005);
nand U18960 (N_18960,N_18377,N_18028);
nand U18961 (N_18961,N_18393,N_18327);
nor U18962 (N_18962,N_18191,N_18313);
and U18963 (N_18963,N_18355,N_18417);
nor U18964 (N_18964,N_18018,N_18147);
nor U18965 (N_18965,N_18406,N_18331);
nor U18966 (N_18966,N_18128,N_18227);
or U18967 (N_18967,N_18333,N_18167);
nand U18968 (N_18968,N_18002,N_18138);
or U18969 (N_18969,N_18068,N_18400);
and U18970 (N_18970,N_18442,N_18432);
or U18971 (N_18971,N_18153,N_18151);
nand U18972 (N_18972,N_18364,N_18012);
nor U18973 (N_18973,N_18159,N_18203);
and U18974 (N_18974,N_18207,N_18311);
nor U18975 (N_18975,N_18440,N_18466);
and U18976 (N_18976,N_18454,N_18033);
xnor U18977 (N_18977,N_18325,N_18273);
nor U18978 (N_18978,N_18488,N_18462);
and U18979 (N_18979,N_18112,N_18201);
nand U18980 (N_18980,N_18186,N_18205);
nand U18981 (N_18981,N_18055,N_18374);
or U18982 (N_18982,N_18114,N_18207);
nor U18983 (N_18983,N_18348,N_18176);
or U18984 (N_18984,N_18297,N_18303);
and U18985 (N_18985,N_18088,N_18252);
or U18986 (N_18986,N_18479,N_18351);
nor U18987 (N_18987,N_18128,N_18463);
or U18988 (N_18988,N_18333,N_18446);
and U18989 (N_18989,N_18334,N_18213);
or U18990 (N_18990,N_18472,N_18165);
and U18991 (N_18991,N_18374,N_18422);
nand U18992 (N_18992,N_18394,N_18423);
nor U18993 (N_18993,N_18296,N_18460);
and U18994 (N_18994,N_18008,N_18036);
nor U18995 (N_18995,N_18207,N_18383);
and U18996 (N_18996,N_18343,N_18182);
or U18997 (N_18997,N_18135,N_18493);
and U18998 (N_18998,N_18335,N_18062);
nand U18999 (N_18999,N_18494,N_18315);
nand U19000 (N_19000,N_18660,N_18888);
nor U19001 (N_19001,N_18739,N_18634);
nor U19002 (N_19002,N_18591,N_18930);
and U19003 (N_19003,N_18706,N_18869);
nor U19004 (N_19004,N_18673,N_18843);
and U19005 (N_19005,N_18893,N_18607);
and U19006 (N_19006,N_18664,N_18854);
and U19007 (N_19007,N_18880,N_18518);
nor U19008 (N_19008,N_18517,N_18697);
or U19009 (N_19009,N_18862,N_18501);
or U19010 (N_19010,N_18514,N_18506);
or U19011 (N_19011,N_18729,N_18910);
nand U19012 (N_19012,N_18923,N_18771);
nand U19013 (N_19013,N_18709,N_18875);
nor U19014 (N_19014,N_18655,N_18887);
and U19015 (N_19015,N_18554,N_18928);
nand U19016 (N_19016,N_18998,N_18553);
nand U19017 (N_19017,N_18797,N_18909);
nor U19018 (N_19018,N_18754,N_18650);
and U19019 (N_19019,N_18544,N_18595);
nand U19020 (N_19020,N_18939,N_18870);
or U19021 (N_19021,N_18704,N_18953);
or U19022 (N_19022,N_18750,N_18512);
nand U19023 (N_19023,N_18614,N_18565);
and U19024 (N_19024,N_18977,N_18736);
or U19025 (N_19025,N_18959,N_18938);
xnor U19026 (N_19026,N_18895,N_18728);
xnor U19027 (N_19027,N_18992,N_18804);
nor U19028 (N_19028,N_18513,N_18916);
nor U19029 (N_19029,N_18999,N_18738);
nor U19030 (N_19030,N_18502,N_18897);
and U19031 (N_19031,N_18546,N_18950);
nor U19032 (N_19032,N_18511,N_18759);
and U19033 (N_19033,N_18883,N_18906);
or U19034 (N_19034,N_18568,N_18859);
and U19035 (N_19035,N_18594,N_18646);
nor U19036 (N_19036,N_18925,N_18872);
and U19037 (N_19037,N_18791,N_18816);
or U19038 (N_19038,N_18764,N_18948);
or U19039 (N_19039,N_18809,N_18579);
or U19040 (N_19040,N_18683,N_18878);
nand U19041 (N_19041,N_18636,N_18629);
nand U19042 (N_19042,N_18719,N_18752);
and U19043 (N_19043,N_18631,N_18756);
xor U19044 (N_19044,N_18755,N_18725);
nor U19045 (N_19045,N_18724,N_18734);
and U19046 (N_19046,N_18622,N_18576);
or U19047 (N_19047,N_18812,N_18933);
or U19048 (N_19048,N_18603,N_18831);
nor U19049 (N_19049,N_18885,N_18913);
xnor U19050 (N_19050,N_18600,N_18991);
nand U19051 (N_19051,N_18645,N_18896);
nand U19052 (N_19052,N_18879,N_18856);
nand U19053 (N_19053,N_18747,N_18765);
nand U19054 (N_19054,N_18860,N_18661);
and U19055 (N_19055,N_18621,N_18592);
and U19056 (N_19056,N_18627,N_18943);
and U19057 (N_19057,N_18782,N_18929);
nor U19058 (N_19058,N_18796,N_18753);
nor U19059 (N_19059,N_18931,N_18882);
xnor U19060 (N_19060,N_18708,N_18844);
and U19061 (N_19061,N_18618,N_18640);
and U19062 (N_19062,N_18767,N_18612);
and U19063 (N_19063,N_18761,N_18902);
and U19064 (N_19064,N_18973,N_18651);
xnor U19065 (N_19065,N_18528,N_18680);
nand U19066 (N_19066,N_18868,N_18996);
nor U19067 (N_19067,N_18519,N_18601);
nor U19068 (N_19068,N_18585,N_18571);
and U19069 (N_19069,N_18714,N_18588);
nor U19070 (N_19070,N_18596,N_18638);
nand U19071 (N_19071,N_18994,N_18965);
nand U19072 (N_19072,N_18670,N_18821);
nor U19073 (N_19073,N_18785,N_18891);
or U19074 (N_19074,N_18707,N_18671);
and U19075 (N_19075,N_18836,N_18881);
and U19076 (N_19076,N_18637,N_18656);
or U19077 (N_19077,N_18749,N_18905);
and U19078 (N_19078,N_18717,N_18962);
nand U19079 (N_19079,N_18613,N_18848);
and U19080 (N_19080,N_18510,N_18907);
or U19081 (N_19081,N_18975,N_18803);
or U19082 (N_19082,N_18653,N_18525);
xnor U19083 (N_19083,N_18863,N_18917);
nor U19084 (N_19084,N_18694,N_18963);
or U19085 (N_19085,N_18847,N_18508);
or U19086 (N_19086,N_18556,N_18572);
nor U19087 (N_19087,N_18827,N_18711);
or U19088 (N_19088,N_18780,N_18951);
nor U19089 (N_19089,N_18678,N_18966);
nand U19090 (N_19090,N_18945,N_18702);
nor U19091 (N_19091,N_18551,N_18699);
nand U19092 (N_19092,N_18985,N_18526);
nor U19093 (N_19093,N_18924,N_18904);
or U19094 (N_19094,N_18609,N_18641);
nor U19095 (N_19095,N_18851,N_18842);
and U19096 (N_19096,N_18748,N_18976);
nor U19097 (N_19097,N_18997,N_18643);
nand U19098 (N_19098,N_18813,N_18871);
nand U19099 (N_19099,N_18583,N_18516);
and U19100 (N_19100,N_18818,N_18611);
and U19101 (N_19101,N_18674,N_18876);
and U19102 (N_19102,N_18632,N_18967);
nor U19103 (N_19103,N_18733,N_18986);
and U19104 (N_19104,N_18838,N_18577);
nor U19105 (N_19105,N_18772,N_18620);
nor U19106 (N_19106,N_18520,N_18690);
or U19107 (N_19107,N_18806,N_18538);
and U19108 (N_19108,N_18777,N_18825);
nand U19109 (N_19109,N_18540,N_18549);
nor U19110 (N_19110,N_18586,N_18988);
nand U19111 (N_19111,N_18617,N_18606);
xor U19112 (N_19112,N_18584,N_18961);
nor U19113 (N_19113,N_18841,N_18555);
nand U19114 (N_19114,N_18679,N_18901);
nand U19115 (N_19115,N_18944,N_18574);
and U19116 (N_19116,N_18658,N_18597);
nand U19117 (N_19117,N_18980,N_18826);
or U19118 (N_19118,N_18745,N_18857);
nor U19119 (N_19119,N_18995,N_18635);
and U19120 (N_19120,N_18539,N_18698);
nor U19121 (N_19121,N_18558,N_18770);
nand U19122 (N_19122,N_18587,N_18846);
or U19123 (N_19123,N_18927,N_18830);
nor U19124 (N_19124,N_18548,N_18524);
or U19125 (N_19125,N_18751,N_18769);
and U19126 (N_19126,N_18937,N_18530);
or U19127 (N_19127,N_18758,N_18908);
or U19128 (N_19128,N_18783,N_18582);
nand U19129 (N_19129,N_18884,N_18919);
and U19130 (N_19130,N_18914,N_18786);
nor U19131 (N_19131,N_18720,N_18956);
and U19132 (N_19132,N_18763,N_18853);
or U19133 (N_19133,N_18993,N_18958);
xnor U19134 (N_19134,N_18529,N_18682);
or U19135 (N_19135,N_18776,N_18955);
and U19136 (N_19136,N_18981,N_18936);
and U19137 (N_19137,N_18760,N_18542);
nor U19138 (N_19138,N_18675,N_18787);
or U19139 (N_19139,N_18799,N_18663);
nor U19140 (N_19140,N_18817,N_18649);
or U19141 (N_19141,N_18504,N_18949);
nor U19142 (N_19142,N_18590,N_18989);
or U19143 (N_19143,N_18899,N_18537);
nand U19144 (N_19144,N_18625,N_18952);
and U19145 (N_19145,N_18811,N_18543);
nor U19146 (N_19146,N_18833,N_18726);
nand U19147 (N_19147,N_18718,N_18766);
xnor U19148 (N_19148,N_18768,N_18557);
nor U19149 (N_19149,N_18560,N_18515);
xnor U19150 (N_19150,N_18805,N_18639);
nand U19151 (N_19151,N_18987,N_18974);
or U19152 (N_19152,N_18500,N_18503);
and U19153 (N_19153,N_18864,N_18969);
nand U19154 (N_19154,N_18834,N_18722);
or U19155 (N_19155,N_18982,N_18934);
xor U19156 (N_19156,N_18795,N_18693);
or U19157 (N_19157,N_18657,N_18593);
nand U19158 (N_19158,N_18781,N_18731);
nor U19159 (N_19159,N_18940,N_18630);
xor U19160 (N_19160,N_18522,N_18921);
xor U19161 (N_19161,N_18866,N_18685);
nor U19162 (N_19162,N_18935,N_18861);
and U19163 (N_19163,N_18608,N_18573);
or U19164 (N_19164,N_18788,N_18835);
nand U19165 (N_19165,N_18903,N_18886);
nor U19166 (N_19166,N_18954,N_18889);
xor U19167 (N_19167,N_18665,N_18941);
or U19168 (N_19168,N_18533,N_18604);
nor U19169 (N_19169,N_18983,N_18534);
nor U19170 (N_19170,N_18695,N_18692);
nor U19171 (N_19171,N_18824,N_18605);
nand U19172 (N_19172,N_18920,N_18915);
nand U19173 (N_19173,N_18688,N_18521);
nand U19174 (N_19174,N_18898,N_18654);
and U19175 (N_19175,N_18561,N_18578);
and U19176 (N_19176,N_18509,N_18684);
or U19177 (N_19177,N_18784,N_18531);
and U19178 (N_19178,N_18648,N_18602);
nand U19179 (N_19179,N_18610,N_18802);
or U19180 (N_19180,N_18662,N_18922);
and U19181 (N_19181,N_18523,N_18800);
nand U19182 (N_19182,N_18822,N_18858);
xnor U19183 (N_19183,N_18840,N_18687);
nand U19184 (N_19184,N_18569,N_18647);
nor U19185 (N_19185,N_18911,N_18735);
nand U19186 (N_19186,N_18689,N_18972);
or U19187 (N_19187,N_18960,N_18918);
nor U19188 (N_19188,N_18676,N_18823);
nor U19189 (N_19189,N_18742,N_18716);
nand U19190 (N_19190,N_18712,N_18740);
nand U19191 (N_19191,N_18723,N_18721);
or U19192 (N_19192,N_18667,N_18743);
or U19193 (N_19193,N_18894,N_18681);
nor U19194 (N_19194,N_18633,N_18810);
and U19195 (N_19195,N_18642,N_18978);
nand U19196 (N_19196,N_18946,N_18652);
and U19197 (N_19197,N_18947,N_18547);
and U19198 (N_19198,N_18527,N_18757);
nor U19199 (N_19199,N_18892,N_18798);
or U19200 (N_19200,N_18552,N_18774);
nand U19201 (N_19201,N_18644,N_18926);
and U19202 (N_19202,N_18619,N_18715);
or U19203 (N_19203,N_18599,N_18626);
nor U19204 (N_19204,N_18666,N_18874);
nand U19205 (N_19205,N_18668,N_18819);
and U19206 (N_19206,N_18705,N_18710);
and U19207 (N_19207,N_18912,N_18775);
and U19208 (N_19208,N_18727,N_18700);
and U19209 (N_19209,N_18900,N_18628);
or U19210 (N_19210,N_18984,N_18794);
xnor U19211 (N_19211,N_18507,N_18616);
or U19212 (N_19212,N_18793,N_18696);
nand U19213 (N_19213,N_18581,N_18566);
nor U19214 (N_19214,N_18762,N_18814);
nor U19215 (N_19215,N_18532,N_18686);
and U19216 (N_19216,N_18580,N_18832);
and U19217 (N_19217,N_18970,N_18541);
or U19218 (N_19218,N_18971,N_18942);
or U19219 (N_19219,N_18563,N_18701);
nor U19220 (N_19220,N_18615,N_18575);
nor U19221 (N_19221,N_18829,N_18850);
and U19222 (N_19222,N_18564,N_18505);
nand U19223 (N_19223,N_18691,N_18932);
nor U19224 (N_19224,N_18659,N_18845);
and U19225 (N_19225,N_18852,N_18623);
nor U19226 (N_19226,N_18815,N_18773);
nor U19227 (N_19227,N_18808,N_18746);
and U19228 (N_19228,N_18672,N_18598);
or U19229 (N_19229,N_18535,N_18545);
nor U19230 (N_19230,N_18828,N_18677);
and U19231 (N_19231,N_18801,N_18867);
nor U19232 (N_19232,N_18669,N_18744);
and U19233 (N_19233,N_18713,N_18839);
and U19234 (N_19234,N_18890,N_18624);
and U19235 (N_19235,N_18741,N_18550);
or U19236 (N_19236,N_18570,N_18807);
nor U19237 (N_19237,N_18778,N_18849);
nand U19238 (N_19238,N_18737,N_18567);
nand U19239 (N_19239,N_18792,N_18790);
and U19240 (N_19240,N_18837,N_18979);
nor U19241 (N_19241,N_18703,N_18877);
nor U19242 (N_19242,N_18779,N_18964);
nor U19243 (N_19243,N_18865,N_18730);
nor U19244 (N_19244,N_18789,N_18957);
nand U19245 (N_19245,N_18855,N_18559);
and U19246 (N_19246,N_18536,N_18990);
and U19247 (N_19247,N_18562,N_18820);
or U19248 (N_19248,N_18732,N_18589);
or U19249 (N_19249,N_18873,N_18968);
or U19250 (N_19250,N_18774,N_18558);
nor U19251 (N_19251,N_18806,N_18574);
and U19252 (N_19252,N_18953,N_18803);
nor U19253 (N_19253,N_18688,N_18967);
and U19254 (N_19254,N_18731,N_18594);
and U19255 (N_19255,N_18838,N_18955);
and U19256 (N_19256,N_18759,N_18531);
or U19257 (N_19257,N_18790,N_18626);
or U19258 (N_19258,N_18974,N_18892);
or U19259 (N_19259,N_18895,N_18846);
nor U19260 (N_19260,N_18592,N_18942);
and U19261 (N_19261,N_18580,N_18672);
nor U19262 (N_19262,N_18773,N_18572);
nand U19263 (N_19263,N_18690,N_18629);
nand U19264 (N_19264,N_18950,N_18975);
nor U19265 (N_19265,N_18987,N_18669);
nand U19266 (N_19266,N_18868,N_18520);
and U19267 (N_19267,N_18739,N_18863);
nand U19268 (N_19268,N_18592,N_18709);
nor U19269 (N_19269,N_18677,N_18734);
xnor U19270 (N_19270,N_18545,N_18757);
and U19271 (N_19271,N_18760,N_18899);
xnor U19272 (N_19272,N_18689,N_18847);
nand U19273 (N_19273,N_18613,N_18765);
and U19274 (N_19274,N_18795,N_18792);
nor U19275 (N_19275,N_18716,N_18704);
and U19276 (N_19276,N_18794,N_18840);
nor U19277 (N_19277,N_18524,N_18869);
and U19278 (N_19278,N_18782,N_18625);
and U19279 (N_19279,N_18674,N_18757);
or U19280 (N_19280,N_18810,N_18986);
and U19281 (N_19281,N_18661,N_18603);
or U19282 (N_19282,N_18892,N_18934);
or U19283 (N_19283,N_18700,N_18567);
nand U19284 (N_19284,N_18616,N_18708);
xnor U19285 (N_19285,N_18599,N_18529);
xor U19286 (N_19286,N_18769,N_18577);
or U19287 (N_19287,N_18559,N_18935);
or U19288 (N_19288,N_18910,N_18678);
nor U19289 (N_19289,N_18806,N_18847);
nand U19290 (N_19290,N_18893,N_18947);
xor U19291 (N_19291,N_18752,N_18880);
nand U19292 (N_19292,N_18910,N_18575);
nor U19293 (N_19293,N_18733,N_18926);
nor U19294 (N_19294,N_18964,N_18930);
nand U19295 (N_19295,N_18663,N_18843);
and U19296 (N_19296,N_18638,N_18735);
or U19297 (N_19297,N_18709,N_18728);
nand U19298 (N_19298,N_18808,N_18523);
nand U19299 (N_19299,N_18769,N_18715);
and U19300 (N_19300,N_18891,N_18743);
nor U19301 (N_19301,N_18759,N_18949);
nor U19302 (N_19302,N_18540,N_18836);
nor U19303 (N_19303,N_18737,N_18875);
xor U19304 (N_19304,N_18934,N_18963);
nand U19305 (N_19305,N_18875,N_18690);
and U19306 (N_19306,N_18508,N_18900);
nand U19307 (N_19307,N_18715,N_18571);
or U19308 (N_19308,N_18894,N_18751);
and U19309 (N_19309,N_18615,N_18955);
and U19310 (N_19310,N_18693,N_18606);
nand U19311 (N_19311,N_18881,N_18591);
nor U19312 (N_19312,N_18514,N_18787);
or U19313 (N_19313,N_18881,N_18900);
nor U19314 (N_19314,N_18681,N_18800);
nand U19315 (N_19315,N_18742,N_18643);
nor U19316 (N_19316,N_18956,N_18820);
nand U19317 (N_19317,N_18702,N_18795);
nor U19318 (N_19318,N_18907,N_18640);
or U19319 (N_19319,N_18857,N_18660);
nor U19320 (N_19320,N_18584,N_18519);
nor U19321 (N_19321,N_18793,N_18640);
nand U19322 (N_19322,N_18743,N_18714);
nand U19323 (N_19323,N_18765,N_18781);
or U19324 (N_19324,N_18568,N_18536);
nor U19325 (N_19325,N_18755,N_18686);
nor U19326 (N_19326,N_18690,N_18649);
xnor U19327 (N_19327,N_18608,N_18889);
xnor U19328 (N_19328,N_18956,N_18536);
xnor U19329 (N_19329,N_18583,N_18813);
nand U19330 (N_19330,N_18985,N_18732);
and U19331 (N_19331,N_18857,N_18545);
nand U19332 (N_19332,N_18540,N_18919);
and U19333 (N_19333,N_18928,N_18994);
nor U19334 (N_19334,N_18519,N_18735);
nand U19335 (N_19335,N_18552,N_18955);
nor U19336 (N_19336,N_18556,N_18936);
and U19337 (N_19337,N_18808,N_18948);
and U19338 (N_19338,N_18922,N_18878);
nor U19339 (N_19339,N_18820,N_18701);
and U19340 (N_19340,N_18823,N_18825);
nor U19341 (N_19341,N_18770,N_18950);
or U19342 (N_19342,N_18998,N_18988);
nor U19343 (N_19343,N_18614,N_18668);
nor U19344 (N_19344,N_18717,N_18525);
xor U19345 (N_19345,N_18736,N_18610);
nand U19346 (N_19346,N_18555,N_18956);
and U19347 (N_19347,N_18547,N_18815);
nor U19348 (N_19348,N_18806,N_18707);
nand U19349 (N_19349,N_18681,N_18597);
or U19350 (N_19350,N_18873,N_18963);
or U19351 (N_19351,N_18878,N_18883);
or U19352 (N_19352,N_18898,N_18953);
nor U19353 (N_19353,N_18805,N_18594);
nor U19354 (N_19354,N_18792,N_18589);
or U19355 (N_19355,N_18886,N_18536);
and U19356 (N_19356,N_18812,N_18840);
or U19357 (N_19357,N_18904,N_18926);
nand U19358 (N_19358,N_18732,N_18714);
or U19359 (N_19359,N_18882,N_18642);
nor U19360 (N_19360,N_18877,N_18652);
or U19361 (N_19361,N_18590,N_18686);
and U19362 (N_19362,N_18876,N_18806);
and U19363 (N_19363,N_18687,N_18893);
nand U19364 (N_19364,N_18574,N_18690);
nor U19365 (N_19365,N_18522,N_18969);
and U19366 (N_19366,N_18972,N_18799);
nor U19367 (N_19367,N_18837,N_18618);
xor U19368 (N_19368,N_18794,N_18709);
nand U19369 (N_19369,N_18912,N_18782);
nor U19370 (N_19370,N_18968,N_18708);
and U19371 (N_19371,N_18929,N_18765);
and U19372 (N_19372,N_18860,N_18666);
and U19373 (N_19373,N_18628,N_18940);
nor U19374 (N_19374,N_18575,N_18902);
nor U19375 (N_19375,N_18673,N_18927);
and U19376 (N_19376,N_18518,N_18991);
or U19377 (N_19377,N_18565,N_18510);
nand U19378 (N_19378,N_18681,N_18885);
nand U19379 (N_19379,N_18790,N_18545);
and U19380 (N_19380,N_18905,N_18584);
nand U19381 (N_19381,N_18515,N_18723);
or U19382 (N_19382,N_18580,N_18978);
and U19383 (N_19383,N_18592,N_18830);
or U19384 (N_19384,N_18642,N_18632);
and U19385 (N_19385,N_18839,N_18551);
nand U19386 (N_19386,N_18894,N_18667);
or U19387 (N_19387,N_18737,N_18508);
or U19388 (N_19388,N_18802,N_18703);
and U19389 (N_19389,N_18791,N_18830);
nor U19390 (N_19390,N_18536,N_18713);
nor U19391 (N_19391,N_18613,N_18616);
nand U19392 (N_19392,N_18911,N_18764);
nor U19393 (N_19393,N_18858,N_18604);
nor U19394 (N_19394,N_18688,N_18824);
nand U19395 (N_19395,N_18558,N_18568);
and U19396 (N_19396,N_18768,N_18739);
and U19397 (N_19397,N_18710,N_18635);
and U19398 (N_19398,N_18576,N_18961);
or U19399 (N_19399,N_18936,N_18619);
nand U19400 (N_19400,N_18918,N_18752);
and U19401 (N_19401,N_18814,N_18606);
or U19402 (N_19402,N_18586,N_18727);
nor U19403 (N_19403,N_18857,N_18549);
xnor U19404 (N_19404,N_18745,N_18748);
nand U19405 (N_19405,N_18765,N_18502);
nor U19406 (N_19406,N_18665,N_18839);
or U19407 (N_19407,N_18888,N_18787);
and U19408 (N_19408,N_18785,N_18532);
or U19409 (N_19409,N_18762,N_18936);
nor U19410 (N_19410,N_18534,N_18518);
and U19411 (N_19411,N_18981,N_18995);
and U19412 (N_19412,N_18909,N_18629);
nand U19413 (N_19413,N_18547,N_18901);
nand U19414 (N_19414,N_18723,N_18650);
and U19415 (N_19415,N_18836,N_18797);
or U19416 (N_19416,N_18743,N_18615);
nor U19417 (N_19417,N_18675,N_18951);
and U19418 (N_19418,N_18588,N_18827);
and U19419 (N_19419,N_18911,N_18700);
or U19420 (N_19420,N_18645,N_18915);
nand U19421 (N_19421,N_18974,N_18767);
nand U19422 (N_19422,N_18946,N_18545);
nor U19423 (N_19423,N_18601,N_18681);
nor U19424 (N_19424,N_18859,N_18788);
xor U19425 (N_19425,N_18695,N_18503);
xor U19426 (N_19426,N_18668,N_18743);
and U19427 (N_19427,N_18918,N_18591);
nand U19428 (N_19428,N_18571,N_18986);
xor U19429 (N_19429,N_18919,N_18783);
xnor U19430 (N_19430,N_18713,N_18803);
and U19431 (N_19431,N_18746,N_18660);
nand U19432 (N_19432,N_18733,N_18571);
or U19433 (N_19433,N_18943,N_18822);
nor U19434 (N_19434,N_18750,N_18955);
or U19435 (N_19435,N_18585,N_18860);
and U19436 (N_19436,N_18722,N_18849);
nor U19437 (N_19437,N_18876,N_18655);
and U19438 (N_19438,N_18804,N_18827);
or U19439 (N_19439,N_18728,N_18977);
or U19440 (N_19440,N_18604,N_18504);
xnor U19441 (N_19441,N_18858,N_18806);
nor U19442 (N_19442,N_18982,N_18614);
nor U19443 (N_19443,N_18682,N_18821);
and U19444 (N_19444,N_18978,N_18799);
and U19445 (N_19445,N_18696,N_18953);
and U19446 (N_19446,N_18956,N_18972);
and U19447 (N_19447,N_18561,N_18931);
nand U19448 (N_19448,N_18922,N_18709);
xnor U19449 (N_19449,N_18670,N_18825);
and U19450 (N_19450,N_18657,N_18553);
nand U19451 (N_19451,N_18993,N_18550);
or U19452 (N_19452,N_18762,N_18993);
or U19453 (N_19453,N_18792,N_18752);
nand U19454 (N_19454,N_18896,N_18589);
nor U19455 (N_19455,N_18537,N_18672);
nor U19456 (N_19456,N_18786,N_18989);
or U19457 (N_19457,N_18864,N_18881);
or U19458 (N_19458,N_18546,N_18984);
nor U19459 (N_19459,N_18769,N_18948);
or U19460 (N_19460,N_18661,N_18867);
or U19461 (N_19461,N_18731,N_18710);
nand U19462 (N_19462,N_18582,N_18798);
nand U19463 (N_19463,N_18561,N_18656);
or U19464 (N_19464,N_18906,N_18582);
and U19465 (N_19465,N_18911,N_18528);
and U19466 (N_19466,N_18842,N_18771);
or U19467 (N_19467,N_18552,N_18894);
and U19468 (N_19468,N_18685,N_18869);
nand U19469 (N_19469,N_18640,N_18916);
and U19470 (N_19470,N_18920,N_18856);
nor U19471 (N_19471,N_18859,N_18939);
nor U19472 (N_19472,N_18778,N_18730);
or U19473 (N_19473,N_18834,N_18901);
nor U19474 (N_19474,N_18713,N_18661);
xnor U19475 (N_19475,N_18700,N_18507);
or U19476 (N_19476,N_18531,N_18537);
or U19477 (N_19477,N_18629,N_18674);
nand U19478 (N_19478,N_18780,N_18678);
nor U19479 (N_19479,N_18845,N_18627);
xor U19480 (N_19480,N_18749,N_18812);
or U19481 (N_19481,N_18719,N_18502);
or U19482 (N_19482,N_18755,N_18652);
nand U19483 (N_19483,N_18743,N_18594);
or U19484 (N_19484,N_18620,N_18696);
nand U19485 (N_19485,N_18800,N_18810);
nand U19486 (N_19486,N_18957,N_18712);
nor U19487 (N_19487,N_18549,N_18780);
nor U19488 (N_19488,N_18524,N_18599);
xnor U19489 (N_19489,N_18951,N_18600);
nand U19490 (N_19490,N_18883,N_18786);
and U19491 (N_19491,N_18593,N_18515);
and U19492 (N_19492,N_18504,N_18906);
nand U19493 (N_19493,N_18832,N_18723);
and U19494 (N_19494,N_18526,N_18751);
nor U19495 (N_19495,N_18626,N_18535);
and U19496 (N_19496,N_18953,N_18989);
and U19497 (N_19497,N_18668,N_18511);
or U19498 (N_19498,N_18901,N_18707);
and U19499 (N_19499,N_18933,N_18666);
nand U19500 (N_19500,N_19278,N_19053);
and U19501 (N_19501,N_19200,N_19319);
nor U19502 (N_19502,N_19494,N_19490);
and U19503 (N_19503,N_19339,N_19499);
xor U19504 (N_19504,N_19195,N_19017);
or U19505 (N_19505,N_19299,N_19227);
and U19506 (N_19506,N_19420,N_19435);
and U19507 (N_19507,N_19259,N_19488);
and U19508 (N_19508,N_19140,N_19412);
nor U19509 (N_19509,N_19433,N_19461);
or U19510 (N_19510,N_19325,N_19457);
nor U19511 (N_19511,N_19192,N_19437);
xnor U19512 (N_19512,N_19027,N_19024);
nor U19513 (N_19513,N_19197,N_19374);
nor U19514 (N_19514,N_19038,N_19232);
and U19515 (N_19515,N_19392,N_19328);
nor U19516 (N_19516,N_19052,N_19338);
nor U19517 (N_19517,N_19079,N_19403);
nor U19518 (N_19518,N_19343,N_19284);
and U19519 (N_19519,N_19096,N_19137);
or U19520 (N_19520,N_19029,N_19005);
or U19521 (N_19521,N_19093,N_19275);
nand U19522 (N_19522,N_19453,N_19240);
nor U19523 (N_19523,N_19154,N_19382);
or U19524 (N_19524,N_19478,N_19318);
and U19525 (N_19525,N_19445,N_19156);
or U19526 (N_19526,N_19273,N_19064);
nand U19527 (N_19527,N_19134,N_19489);
or U19528 (N_19528,N_19250,N_19108);
nor U19529 (N_19529,N_19400,N_19257);
and U19530 (N_19530,N_19495,N_19071);
or U19531 (N_19531,N_19062,N_19237);
or U19532 (N_19532,N_19394,N_19133);
or U19533 (N_19533,N_19158,N_19149);
nand U19534 (N_19534,N_19280,N_19235);
and U19535 (N_19535,N_19363,N_19212);
xor U19536 (N_19536,N_19407,N_19182);
and U19537 (N_19537,N_19152,N_19123);
nand U19538 (N_19538,N_19099,N_19268);
or U19539 (N_19539,N_19039,N_19314);
and U19540 (N_19540,N_19308,N_19312);
nand U19541 (N_19541,N_19463,N_19146);
or U19542 (N_19542,N_19413,N_19411);
nand U19543 (N_19543,N_19124,N_19417);
nor U19544 (N_19544,N_19387,N_19467);
or U19545 (N_19545,N_19384,N_19443);
nor U19546 (N_19546,N_19393,N_19125);
nand U19547 (N_19547,N_19160,N_19065);
nand U19548 (N_19548,N_19132,N_19444);
and U19549 (N_19549,N_19277,N_19342);
xor U19550 (N_19550,N_19440,N_19239);
nor U19551 (N_19551,N_19205,N_19150);
and U19552 (N_19552,N_19424,N_19097);
or U19553 (N_19553,N_19088,N_19317);
nand U19554 (N_19554,N_19376,N_19370);
and U19555 (N_19555,N_19247,N_19470);
xor U19556 (N_19556,N_19050,N_19094);
and U19557 (N_19557,N_19040,N_19196);
nor U19558 (N_19558,N_19448,N_19310);
and U19559 (N_19559,N_19429,N_19341);
nand U19560 (N_19560,N_19270,N_19077);
and U19561 (N_19561,N_19436,N_19164);
nor U19562 (N_19562,N_19049,N_19054);
nand U19563 (N_19563,N_19383,N_19224);
nand U19564 (N_19564,N_19110,N_19352);
or U19565 (N_19565,N_19203,N_19207);
and U19566 (N_19566,N_19476,N_19129);
or U19567 (N_19567,N_19460,N_19036);
nand U19568 (N_19568,N_19191,N_19416);
or U19569 (N_19569,N_19183,N_19324);
nand U19570 (N_19570,N_19210,N_19114);
and U19571 (N_19571,N_19090,N_19174);
or U19572 (N_19572,N_19288,N_19332);
and U19573 (N_19573,N_19431,N_19037);
nand U19574 (N_19574,N_19218,N_19272);
and U19575 (N_19575,N_19209,N_19215);
or U19576 (N_19576,N_19241,N_19472);
nor U19577 (N_19577,N_19311,N_19464);
xnor U19578 (N_19578,N_19087,N_19139);
or U19579 (N_19579,N_19320,N_19057);
and U19580 (N_19580,N_19131,N_19035);
and U19581 (N_19581,N_19377,N_19153);
nor U19582 (N_19582,N_19373,N_19439);
or U19583 (N_19583,N_19419,N_19059);
and U19584 (N_19584,N_19135,N_19089);
and U19585 (N_19585,N_19178,N_19327);
or U19586 (N_19586,N_19006,N_19043);
nand U19587 (N_19587,N_19186,N_19009);
nand U19588 (N_19588,N_19402,N_19010);
nor U19589 (N_19589,N_19347,N_19300);
or U19590 (N_19590,N_19265,N_19034);
nand U19591 (N_19591,N_19198,N_19348);
xnor U19592 (N_19592,N_19112,N_19078);
or U19593 (N_19593,N_19172,N_19161);
or U19594 (N_19594,N_19000,N_19386);
and U19595 (N_19595,N_19359,N_19001);
nand U19596 (N_19596,N_19408,N_19122);
and U19597 (N_19597,N_19498,N_19331);
or U19598 (N_19598,N_19365,N_19118);
nor U19599 (N_19599,N_19244,N_19107);
nor U19600 (N_19600,N_19362,N_19167);
nand U19601 (N_19601,N_19350,N_19111);
and U19602 (N_19602,N_19143,N_19165);
or U19603 (N_19603,N_19357,N_19014);
nand U19604 (N_19604,N_19345,N_19313);
nor U19605 (N_19605,N_19441,N_19261);
and U19606 (N_19606,N_19294,N_19217);
or U19607 (N_19607,N_19260,N_19126);
nand U19608 (N_19608,N_19222,N_19425);
and U19609 (N_19609,N_19011,N_19199);
nand U19610 (N_19610,N_19423,N_19296);
nand U19611 (N_19611,N_19041,N_19105);
nor U19612 (N_19612,N_19303,N_19354);
nor U19613 (N_19613,N_19360,N_19026);
or U19614 (N_19614,N_19101,N_19058);
nand U19615 (N_19615,N_19389,N_19381);
or U19616 (N_19616,N_19283,N_19493);
nor U19617 (N_19617,N_19368,N_19007);
nor U19618 (N_19618,N_19475,N_19030);
and U19619 (N_19619,N_19100,N_19166);
nand U19620 (N_19620,N_19204,N_19072);
xnor U19621 (N_19621,N_19438,N_19267);
nand U19622 (N_19622,N_19119,N_19144);
nand U19623 (N_19623,N_19432,N_19208);
nand U19624 (N_19624,N_19349,N_19371);
or U19625 (N_19625,N_19255,N_19206);
and U19626 (N_19626,N_19379,N_19086);
nor U19627 (N_19627,N_19301,N_19326);
nor U19628 (N_19628,N_19292,N_19388);
and U19629 (N_19629,N_19455,N_19117);
nand U19630 (N_19630,N_19397,N_19449);
xor U19631 (N_19631,N_19015,N_19102);
xnor U19632 (N_19632,N_19194,N_19337);
nor U19633 (N_19633,N_19002,N_19375);
or U19634 (N_19634,N_19290,N_19075);
nor U19635 (N_19635,N_19462,N_19142);
nand U19636 (N_19636,N_19098,N_19080);
nand U19637 (N_19637,N_19391,N_19287);
and U19638 (N_19638,N_19378,N_19297);
nand U19639 (N_19639,N_19266,N_19473);
nor U19640 (N_19640,N_19229,N_19155);
and U19641 (N_19641,N_19068,N_19380);
nor U19642 (N_19642,N_19390,N_19019);
nand U19643 (N_19643,N_19016,N_19447);
and U19644 (N_19644,N_19483,N_19056);
nand U19645 (N_19645,N_19293,N_19279);
nand U19646 (N_19646,N_19410,N_19151);
or U19647 (N_19647,N_19091,N_19334);
or U19648 (N_19648,N_19329,N_19055);
nor U19649 (N_19649,N_19022,N_19282);
or U19650 (N_19650,N_19095,N_19415);
nor U19651 (N_19651,N_19385,N_19076);
and U19652 (N_19652,N_19304,N_19451);
and U19653 (N_19653,N_19487,N_19236);
nor U19654 (N_19654,N_19248,N_19398);
nor U19655 (N_19655,N_19092,N_19231);
nor U19656 (N_19656,N_19477,N_19193);
or U19657 (N_19657,N_19061,N_19262);
nor U19658 (N_19658,N_19322,N_19169);
nor U19659 (N_19659,N_19456,N_19189);
and U19660 (N_19660,N_19335,N_19213);
and U19661 (N_19661,N_19033,N_19221);
or U19662 (N_19662,N_19353,N_19175);
nand U19663 (N_19663,N_19163,N_19276);
nand U19664 (N_19664,N_19289,N_19471);
nand U19665 (N_19665,N_19228,N_19474);
and U19666 (N_19666,N_19021,N_19285);
and U19667 (N_19667,N_19246,N_19252);
and U19668 (N_19668,N_19426,N_19253);
nor U19669 (N_19669,N_19355,N_19148);
nand U19670 (N_19670,N_19184,N_19047);
nor U19671 (N_19671,N_19269,N_19004);
xor U19672 (N_19672,N_19031,N_19136);
or U19673 (N_19673,N_19177,N_19109);
nor U19674 (N_19674,N_19141,N_19067);
and U19675 (N_19675,N_19323,N_19168);
nor U19676 (N_19676,N_19020,N_19083);
and U19677 (N_19677,N_19251,N_19295);
or U19678 (N_19678,N_19263,N_19344);
and U19679 (N_19679,N_19286,N_19220);
nor U19680 (N_19680,N_19333,N_19216);
or U19681 (N_19681,N_19479,N_19316);
nand U19682 (N_19682,N_19045,N_19181);
nand U19683 (N_19683,N_19446,N_19185);
and U19684 (N_19684,N_19482,N_19306);
nand U19685 (N_19685,N_19302,N_19157);
xor U19686 (N_19686,N_19115,N_19491);
nor U19687 (N_19687,N_19104,N_19060);
or U19688 (N_19688,N_19340,N_19361);
or U19689 (N_19689,N_19048,N_19082);
nor U19690 (N_19690,N_19013,N_19330);
nand U19691 (N_19691,N_19234,N_19271);
and U19692 (N_19692,N_19452,N_19414);
xnor U19693 (N_19693,N_19305,N_19046);
nor U19694 (N_19694,N_19147,N_19492);
nor U19695 (N_19695,N_19063,N_19480);
nand U19696 (N_19696,N_19214,N_19485);
and U19697 (N_19697,N_19066,N_19405);
or U19698 (N_19698,N_19138,N_19409);
nor U19699 (N_19699,N_19187,N_19434);
and U19700 (N_19700,N_19003,N_19442);
nand U19701 (N_19701,N_19226,N_19481);
xor U19702 (N_19702,N_19298,N_19404);
and U19703 (N_19703,N_19421,N_19202);
nor U19704 (N_19704,N_19008,N_19012);
or U19705 (N_19705,N_19372,N_19070);
nand U19706 (N_19706,N_19084,N_19256);
and U19707 (N_19707,N_19468,N_19291);
nand U19708 (N_19708,N_19121,N_19309);
nor U19709 (N_19709,N_19281,N_19025);
or U19710 (N_19710,N_19127,N_19497);
nand U19711 (N_19711,N_19106,N_19116);
and U19712 (N_19712,N_19085,N_19179);
nand U19713 (N_19713,N_19395,N_19336);
nor U19714 (N_19714,N_19364,N_19170);
xor U19715 (N_19715,N_19230,N_19428);
xor U19716 (N_19716,N_19018,N_19238);
nand U19717 (N_19717,N_19358,N_19346);
nor U19718 (N_19718,N_19351,N_19307);
or U19719 (N_19719,N_19465,N_19450);
nand U19720 (N_19720,N_19315,N_19249);
xnor U19721 (N_19721,N_19225,N_19173);
and U19722 (N_19722,N_19171,N_19254);
or U19723 (N_19723,N_19113,N_19176);
and U19724 (N_19724,N_19396,N_19130);
and U19725 (N_19725,N_19044,N_19103);
nand U19726 (N_19726,N_19128,N_19369);
nand U19727 (N_19727,N_19399,N_19023);
and U19728 (N_19728,N_19120,N_19274);
nand U19729 (N_19729,N_19454,N_19243);
nand U19730 (N_19730,N_19258,N_19430);
nand U19731 (N_19731,N_19401,N_19145);
or U19732 (N_19732,N_19486,N_19418);
nand U19733 (N_19733,N_19422,N_19081);
nor U19734 (N_19734,N_19042,N_19245);
nor U19735 (N_19735,N_19223,N_19201);
or U19736 (N_19736,N_19233,N_19406);
and U19737 (N_19737,N_19484,N_19264);
or U19738 (N_19738,N_19074,N_19356);
or U19739 (N_19739,N_19367,N_19051);
nand U19740 (N_19740,N_19219,N_19466);
xor U19741 (N_19741,N_19458,N_19028);
nand U19742 (N_19742,N_19032,N_19427);
or U19743 (N_19743,N_19069,N_19190);
xor U19744 (N_19744,N_19073,N_19496);
nor U19745 (N_19745,N_19180,N_19211);
and U19746 (N_19746,N_19188,N_19366);
xnor U19747 (N_19747,N_19162,N_19459);
and U19748 (N_19748,N_19242,N_19321);
or U19749 (N_19749,N_19469,N_19159);
xor U19750 (N_19750,N_19491,N_19125);
and U19751 (N_19751,N_19030,N_19321);
and U19752 (N_19752,N_19209,N_19290);
and U19753 (N_19753,N_19008,N_19451);
nand U19754 (N_19754,N_19227,N_19201);
or U19755 (N_19755,N_19270,N_19021);
nand U19756 (N_19756,N_19262,N_19297);
xnor U19757 (N_19757,N_19263,N_19019);
nor U19758 (N_19758,N_19192,N_19306);
xor U19759 (N_19759,N_19301,N_19291);
nand U19760 (N_19760,N_19050,N_19412);
nor U19761 (N_19761,N_19462,N_19266);
or U19762 (N_19762,N_19280,N_19392);
and U19763 (N_19763,N_19124,N_19173);
nand U19764 (N_19764,N_19336,N_19021);
nand U19765 (N_19765,N_19390,N_19418);
nor U19766 (N_19766,N_19093,N_19290);
and U19767 (N_19767,N_19267,N_19345);
nand U19768 (N_19768,N_19276,N_19424);
nand U19769 (N_19769,N_19498,N_19075);
nand U19770 (N_19770,N_19174,N_19016);
xnor U19771 (N_19771,N_19001,N_19209);
and U19772 (N_19772,N_19021,N_19182);
and U19773 (N_19773,N_19422,N_19380);
and U19774 (N_19774,N_19180,N_19051);
or U19775 (N_19775,N_19128,N_19130);
and U19776 (N_19776,N_19330,N_19035);
nor U19777 (N_19777,N_19471,N_19337);
or U19778 (N_19778,N_19473,N_19420);
and U19779 (N_19779,N_19410,N_19271);
or U19780 (N_19780,N_19303,N_19056);
and U19781 (N_19781,N_19437,N_19442);
or U19782 (N_19782,N_19204,N_19367);
nor U19783 (N_19783,N_19061,N_19067);
nor U19784 (N_19784,N_19084,N_19468);
and U19785 (N_19785,N_19092,N_19322);
nand U19786 (N_19786,N_19341,N_19377);
nand U19787 (N_19787,N_19333,N_19484);
and U19788 (N_19788,N_19071,N_19414);
nor U19789 (N_19789,N_19299,N_19473);
or U19790 (N_19790,N_19390,N_19436);
and U19791 (N_19791,N_19289,N_19383);
nor U19792 (N_19792,N_19058,N_19001);
nand U19793 (N_19793,N_19102,N_19113);
nand U19794 (N_19794,N_19418,N_19292);
nor U19795 (N_19795,N_19328,N_19120);
and U19796 (N_19796,N_19418,N_19065);
xor U19797 (N_19797,N_19399,N_19132);
nor U19798 (N_19798,N_19155,N_19032);
xor U19799 (N_19799,N_19121,N_19141);
nor U19800 (N_19800,N_19383,N_19275);
and U19801 (N_19801,N_19117,N_19032);
and U19802 (N_19802,N_19484,N_19385);
or U19803 (N_19803,N_19153,N_19292);
or U19804 (N_19804,N_19090,N_19437);
and U19805 (N_19805,N_19032,N_19336);
and U19806 (N_19806,N_19445,N_19125);
or U19807 (N_19807,N_19258,N_19009);
nand U19808 (N_19808,N_19125,N_19105);
nor U19809 (N_19809,N_19471,N_19221);
nor U19810 (N_19810,N_19325,N_19009);
nor U19811 (N_19811,N_19489,N_19442);
nand U19812 (N_19812,N_19325,N_19413);
nand U19813 (N_19813,N_19139,N_19218);
xor U19814 (N_19814,N_19178,N_19083);
or U19815 (N_19815,N_19411,N_19010);
or U19816 (N_19816,N_19139,N_19041);
and U19817 (N_19817,N_19338,N_19219);
nor U19818 (N_19818,N_19283,N_19440);
or U19819 (N_19819,N_19254,N_19218);
nor U19820 (N_19820,N_19436,N_19342);
and U19821 (N_19821,N_19493,N_19490);
and U19822 (N_19822,N_19393,N_19387);
nor U19823 (N_19823,N_19476,N_19270);
or U19824 (N_19824,N_19352,N_19135);
or U19825 (N_19825,N_19103,N_19039);
nand U19826 (N_19826,N_19340,N_19101);
nor U19827 (N_19827,N_19325,N_19274);
nand U19828 (N_19828,N_19436,N_19137);
xor U19829 (N_19829,N_19058,N_19402);
and U19830 (N_19830,N_19409,N_19494);
nand U19831 (N_19831,N_19006,N_19250);
nor U19832 (N_19832,N_19379,N_19465);
and U19833 (N_19833,N_19174,N_19192);
nand U19834 (N_19834,N_19497,N_19307);
and U19835 (N_19835,N_19092,N_19317);
or U19836 (N_19836,N_19409,N_19402);
nand U19837 (N_19837,N_19266,N_19121);
and U19838 (N_19838,N_19442,N_19091);
nor U19839 (N_19839,N_19226,N_19113);
and U19840 (N_19840,N_19128,N_19028);
xnor U19841 (N_19841,N_19343,N_19345);
or U19842 (N_19842,N_19225,N_19172);
and U19843 (N_19843,N_19311,N_19235);
and U19844 (N_19844,N_19067,N_19302);
nand U19845 (N_19845,N_19235,N_19061);
or U19846 (N_19846,N_19297,N_19337);
xor U19847 (N_19847,N_19164,N_19348);
and U19848 (N_19848,N_19218,N_19135);
or U19849 (N_19849,N_19271,N_19306);
or U19850 (N_19850,N_19279,N_19163);
nor U19851 (N_19851,N_19030,N_19055);
nor U19852 (N_19852,N_19279,N_19286);
and U19853 (N_19853,N_19024,N_19367);
nor U19854 (N_19854,N_19066,N_19211);
or U19855 (N_19855,N_19301,N_19104);
nor U19856 (N_19856,N_19001,N_19364);
nand U19857 (N_19857,N_19329,N_19380);
or U19858 (N_19858,N_19199,N_19020);
nor U19859 (N_19859,N_19395,N_19387);
nand U19860 (N_19860,N_19453,N_19082);
and U19861 (N_19861,N_19101,N_19160);
or U19862 (N_19862,N_19236,N_19300);
or U19863 (N_19863,N_19275,N_19251);
nand U19864 (N_19864,N_19148,N_19130);
or U19865 (N_19865,N_19206,N_19099);
and U19866 (N_19866,N_19304,N_19193);
nor U19867 (N_19867,N_19351,N_19150);
or U19868 (N_19868,N_19343,N_19370);
or U19869 (N_19869,N_19103,N_19181);
and U19870 (N_19870,N_19450,N_19284);
xnor U19871 (N_19871,N_19199,N_19126);
nand U19872 (N_19872,N_19068,N_19030);
nand U19873 (N_19873,N_19141,N_19378);
nor U19874 (N_19874,N_19136,N_19377);
nand U19875 (N_19875,N_19370,N_19085);
nor U19876 (N_19876,N_19314,N_19249);
or U19877 (N_19877,N_19188,N_19364);
nand U19878 (N_19878,N_19230,N_19476);
and U19879 (N_19879,N_19386,N_19183);
nand U19880 (N_19880,N_19243,N_19052);
nand U19881 (N_19881,N_19268,N_19394);
and U19882 (N_19882,N_19186,N_19287);
nand U19883 (N_19883,N_19289,N_19181);
nor U19884 (N_19884,N_19071,N_19332);
nand U19885 (N_19885,N_19206,N_19307);
or U19886 (N_19886,N_19427,N_19480);
nand U19887 (N_19887,N_19285,N_19332);
and U19888 (N_19888,N_19136,N_19400);
or U19889 (N_19889,N_19306,N_19010);
nand U19890 (N_19890,N_19235,N_19123);
and U19891 (N_19891,N_19353,N_19477);
nand U19892 (N_19892,N_19211,N_19256);
nand U19893 (N_19893,N_19001,N_19400);
nor U19894 (N_19894,N_19314,N_19142);
and U19895 (N_19895,N_19143,N_19021);
and U19896 (N_19896,N_19227,N_19074);
or U19897 (N_19897,N_19487,N_19467);
and U19898 (N_19898,N_19017,N_19008);
nand U19899 (N_19899,N_19365,N_19109);
nand U19900 (N_19900,N_19488,N_19124);
or U19901 (N_19901,N_19027,N_19063);
xor U19902 (N_19902,N_19369,N_19380);
nand U19903 (N_19903,N_19283,N_19103);
xnor U19904 (N_19904,N_19493,N_19461);
and U19905 (N_19905,N_19029,N_19292);
and U19906 (N_19906,N_19400,N_19029);
or U19907 (N_19907,N_19022,N_19333);
and U19908 (N_19908,N_19347,N_19150);
or U19909 (N_19909,N_19437,N_19355);
and U19910 (N_19910,N_19091,N_19378);
or U19911 (N_19911,N_19353,N_19448);
and U19912 (N_19912,N_19375,N_19119);
nor U19913 (N_19913,N_19382,N_19156);
nor U19914 (N_19914,N_19144,N_19459);
or U19915 (N_19915,N_19340,N_19403);
nand U19916 (N_19916,N_19472,N_19483);
and U19917 (N_19917,N_19092,N_19254);
and U19918 (N_19918,N_19001,N_19450);
or U19919 (N_19919,N_19133,N_19084);
and U19920 (N_19920,N_19178,N_19038);
or U19921 (N_19921,N_19018,N_19388);
and U19922 (N_19922,N_19433,N_19160);
nand U19923 (N_19923,N_19228,N_19321);
nand U19924 (N_19924,N_19384,N_19297);
and U19925 (N_19925,N_19009,N_19406);
nor U19926 (N_19926,N_19248,N_19352);
nand U19927 (N_19927,N_19485,N_19035);
nand U19928 (N_19928,N_19290,N_19137);
xor U19929 (N_19929,N_19333,N_19228);
nand U19930 (N_19930,N_19336,N_19231);
or U19931 (N_19931,N_19064,N_19450);
xnor U19932 (N_19932,N_19079,N_19035);
nand U19933 (N_19933,N_19188,N_19355);
xnor U19934 (N_19934,N_19245,N_19428);
or U19935 (N_19935,N_19310,N_19097);
and U19936 (N_19936,N_19334,N_19481);
nor U19937 (N_19937,N_19415,N_19145);
or U19938 (N_19938,N_19328,N_19215);
nor U19939 (N_19939,N_19433,N_19140);
or U19940 (N_19940,N_19319,N_19213);
or U19941 (N_19941,N_19065,N_19369);
and U19942 (N_19942,N_19485,N_19216);
nor U19943 (N_19943,N_19485,N_19164);
nor U19944 (N_19944,N_19086,N_19459);
nand U19945 (N_19945,N_19273,N_19062);
nand U19946 (N_19946,N_19422,N_19449);
or U19947 (N_19947,N_19384,N_19399);
or U19948 (N_19948,N_19442,N_19009);
or U19949 (N_19949,N_19109,N_19165);
xor U19950 (N_19950,N_19164,N_19014);
and U19951 (N_19951,N_19395,N_19268);
xor U19952 (N_19952,N_19493,N_19142);
nand U19953 (N_19953,N_19478,N_19311);
or U19954 (N_19954,N_19275,N_19050);
or U19955 (N_19955,N_19152,N_19415);
nor U19956 (N_19956,N_19219,N_19396);
or U19957 (N_19957,N_19150,N_19284);
or U19958 (N_19958,N_19167,N_19437);
nor U19959 (N_19959,N_19429,N_19306);
or U19960 (N_19960,N_19484,N_19026);
or U19961 (N_19961,N_19293,N_19456);
and U19962 (N_19962,N_19099,N_19111);
nand U19963 (N_19963,N_19253,N_19457);
xnor U19964 (N_19964,N_19068,N_19104);
xnor U19965 (N_19965,N_19289,N_19331);
nor U19966 (N_19966,N_19349,N_19121);
nand U19967 (N_19967,N_19433,N_19273);
xor U19968 (N_19968,N_19024,N_19461);
nand U19969 (N_19969,N_19084,N_19116);
nor U19970 (N_19970,N_19459,N_19372);
nor U19971 (N_19971,N_19229,N_19393);
or U19972 (N_19972,N_19271,N_19332);
and U19973 (N_19973,N_19391,N_19195);
nand U19974 (N_19974,N_19174,N_19277);
or U19975 (N_19975,N_19255,N_19346);
and U19976 (N_19976,N_19407,N_19128);
nor U19977 (N_19977,N_19360,N_19326);
or U19978 (N_19978,N_19447,N_19388);
xor U19979 (N_19979,N_19337,N_19141);
nor U19980 (N_19980,N_19150,N_19499);
nand U19981 (N_19981,N_19327,N_19127);
and U19982 (N_19982,N_19217,N_19152);
nor U19983 (N_19983,N_19428,N_19316);
nand U19984 (N_19984,N_19375,N_19241);
or U19985 (N_19985,N_19477,N_19127);
or U19986 (N_19986,N_19088,N_19448);
or U19987 (N_19987,N_19181,N_19159);
nor U19988 (N_19988,N_19256,N_19400);
or U19989 (N_19989,N_19454,N_19158);
and U19990 (N_19990,N_19468,N_19393);
or U19991 (N_19991,N_19365,N_19481);
xnor U19992 (N_19992,N_19279,N_19220);
nand U19993 (N_19993,N_19281,N_19470);
or U19994 (N_19994,N_19241,N_19227);
or U19995 (N_19995,N_19354,N_19158);
or U19996 (N_19996,N_19242,N_19059);
nor U19997 (N_19997,N_19276,N_19182);
and U19998 (N_19998,N_19371,N_19331);
and U19999 (N_19999,N_19205,N_19480);
nor UO_0 (O_0,N_19857,N_19502);
and UO_1 (O_1,N_19988,N_19706);
and UO_2 (O_2,N_19916,N_19518);
and UO_3 (O_3,N_19892,N_19925);
xor UO_4 (O_4,N_19727,N_19555);
nand UO_5 (O_5,N_19508,N_19985);
xor UO_6 (O_6,N_19658,N_19500);
or UO_7 (O_7,N_19789,N_19901);
nor UO_8 (O_8,N_19694,N_19856);
or UO_9 (O_9,N_19757,N_19840);
nand UO_10 (O_10,N_19955,N_19854);
nor UO_11 (O_11,N_19516,N_19534);
and UO_12 (O_12,N_19963,N_19893);
nand UO_13 (O_13,N_19818,N_19728);
nand UO_14 (O_14,N_19725,N_19790);
and UO_15 (O_15,N_19842,N_19866);
and UO_16 (O_16,N_19904,N_19792);
and UO_17 (O_17,N_19646,N_19689);
and UO_18 (O_18,N_19519,N_19768);
and UO_19 (O_19,N_19656,N_19505);
nand UO_20 (O_20,N_19585,N_19573);
nand UO_21 (O_21,N_19870,N_19816);
xnor UO_22 (O_22,N_19962,N_19619);
nand UO_23 (O_23,N_19843,N_19948);
nor UO_24 (O_24,N_19788,N_19986);
or UO_25 (O_25,N_19859,N_19543);
nor UO_26 (O_26,N_19588,N_19660);
or UO_27 (O_27,N_19596,N_19874);
nor UO_28 (O_28,N_19635,N_19592);
or UO_29 (O_29,N_19535,N_19864);
or UO_30 (O_30,N_19993,N_19712);
or UO_31 (O_31,N_19702,N_19742);
xnor UO_32 (O_32,N_19616,N_19614);
and UO_33 (O_33,N_19610,N_19553);
nand UO_34 (O_34,N_19591,N_19775);
nand UO_35 (O_35,N_19523,N_19629);
and UO_36 (O_36,N_19741,N_19883);
nand UO_37 (O_37,N_19997,N_19782);
nor UO_38 (O_38,N_19525,N_19644);
or UO_39 (O_39,N_19559,N_19894);
nor UO_40 (O_40,N_19922,N_19888);
and UO_41 (O_41,N_19846,N_19550);
nand UO_42 (O_42,N_19514,N_19618);
and UO_43 (O_43,N_19628,N_19708);
xnor UO_44 (O_44,N_19544,N_19670);
nor UO_45 (O_45,N_19839,N_19510);
and UO_46 (O_46,N_19957,N_19785);
nor UO_47 (O_47,N_19806,N_19504);
nand UO_48 (O_48,N_19528,N_19717);
or UO_49 (O_49,N_19898,N_19969);
and UO_50 (O_50,N_19677,N_19844);
nand UO_51 (O_51,N_19736,N_19719);
and UO_52 (O_52,N_19675,N_19795);
nor UO_53 (O_53,N_19624,N_19587);
or UO_54 (O_54,N_19650,N_19828);
and UO_55 (O_55,N_19581,N_19820);
nor UO_56 (O_56,N_19853,N_19756);
and UO_57 (O_57,N_19873,N_19762);
or UO_58 (O_58,N_19634,N_19990);
nor UO_59 (O_59,N_19558,N_19776);
nand UO_60 (O_60,N_19620,N_19590);
and UO_61 (O_61,N_19529,N_19766);
xnor UO_62 (O_62,N_19750,N_19944);
nor UO_63 (O_63,N_19917,N_19851);
xor UO_64 (O_64,N_19765,N_19819);
nand UO_65 (O_65,N_19810,N_19815);
xnor UO_66 (O_66,N_19764,N_19907);
or UO_67 (O_67,N_19729,N_19684);
nor UO_68 (O_68,N_19976,N_19730);
nor UO_69 (O_69,N_19982,N_19805);
or UO_70 (O_70,N_19605,N_19556);
and UO_71 (O_71,N_19784,N_19511);
nor UO_72 (O_72,N_19902,N_19950);
nand UO_73 (O_73,N_19512,N_19759);
nor UO_74 (O_74,N_19612,N_19509);
nor UO_75 (O_75,N_19603,N_19974);
xnor UO_76 (O_76,N_19699,N_19723);
or UO_77 (O_77,N_19769,N_19631);
and UO_78 (O_78,N_19632,N_19659);
nand UO_79 (O_79,N_19607,N_19623);
nor UO_80 (O_80,N_19935,N_19606);
xnor UO_81 (O_81,N_19862,N_19771);
nor UO_82 (O_82,N_19696,N_19520);
or UO_83 (O_83,N_19597,N_19928);
nand UO_84 (O_84,N_19536,N_19869);
or UO_85 (O_85,N_19823,N_19897);
nor UO_86 (O_86,N_19995,N_19682);
and UO_87 (O_87,N_19945,N_19919);
or UO_88 (O_88,N_19680,N_19861);
or UO_89 (O_89,N_19633,N_19895);
nand UO_90 (O_90,N_19979,N_19927);
nand UO_91 (O_91,N_19664,N_19994);
nand UO_92 (O_92,N_19551,N_19726);
and UO_93 (O_93,N_19887,N_19686);
nand UO_94 (O_94,N_19942,N_19989);
or UO_95 (O_95,N_19651,N_19630);
nand UO_96 (O_96,N_19754,N_19731);
nor UO_97 (O_97,N_19662,N_19787);
xnor UO_98 (O_98,N_19875,N_19809);
nor UO_99 (O_99,N_19714,N_19746);
nor UO_100 (O_100,N_19586,N_19937);
or UO_101 (O_101,N_19931,N_19999);
and UO_102 (O_102,N_19733,N_19740);
and UO_103 (O_103,N_19913,N_19835);
xnor UO_104 (O_104,N_19577,N_19625);
and UO_105 (O_105,N_19817,N_19583);
and UO_106 (O_106,N_19705,N_19745);
xnor UO_107 (O_107,N_19517,N_19698);
xor UO_108 (O_108,N_19896,N_19802);
and UO_109 (O_109,N_19506,N_19540);
or UO_110 (O_110,N_19803,N_19710);
or UO_111 (O_111,N_19949,N_19753);
xor UO_112 (O_112,N_19552,N_19831);
nand UO_113 (O_113,N_19991,N_19739);
nand UO_114 (O_114,N_19911,N_19565);
and UO_115 (O_115,N_19539,N_19983);
nor UO_116 (O_116,N_19637,N_19568);
nor UO_117 (O_117,N_19882,N_19527);
xnor UO_118 (O_118,N_19977,N_19665);
nor UO_119 (O_119,N_19779,N_19821);
xnor UO_120 (O_120,N_19563,N_19915);
nand UO_121 (O_121,N_19910,N_19700);
nand UO_122 (O_122,N_19829,N_19538);
nand UO_123 (O_123,N_19797,N_19521);
xor UO_124 (O_124,N_19501,N_19826);
or UO_125 (O_125,N_19643,N_19626);
and UO_126 (O_126,N_19681,N_19669);
or UO_127 (O_127,N_19807,N_19661);
nor UO_128 (O_128,N_19960,N_19780);
nand UO_129 (O_129,N_19713,N_19560);
and UO_130 (O_130,N_19971,N_19691);
nor UO_131 (O_131,N_19751,N_19783);
or UO_132 (O_132,N_19732,N_19621);
or UO_133 (O_133,N_19611,N_19881);
xnor UO_134 (O_134,N_19777,N_19852);
nor UO_135 (O_135,N_19940,N_19956);
nand UO_136 (O_136,N_19522,N_19825);
nand UO_137 (O_137,N_19668,N_19965);
nor UO_138 (O_138,N_19758,N_19532);
or UO_139 (O_139,N_19721,N_19655);
or UO_140 (O_140,N_19570,N_19770);
nand UO_141 (O_141,N_19755,N_19834);
and UO_142 (O_142,N_19947,N_19863);
or UO_143 (O_143,N_19930,N_19526);
nand UO_144 (O_144,N_19791,N_19921);
nor UO_145 (O_145,N_19918,N_19850);
nand UO_146 (O_146,N_19871,N_19608);
xor UO_147 (O_147,N_19647,N_19934);
nand UO_148 (O_148,N_19545,N_19849);
nor UO_149 (O_149,N_19679,N_19830);
nor UO_150 (O_150,N_19941,N_19980);
nor UO_151 (O_151,N_19507,N_19760);
and UO_152 (O_152,N_19909,N_19613);
or UO_153 (O_153,N_19879,N_19649);
and UO_154 (O_154,N_19808,N_19672);
nor UO_155 (O_155,N_19833,N_19752);
or UO_156 (O_156,N_19800,N_19533);
nor UO_157 (O_157,N_19569,N_19848);
and UO_158 (O_158,N_19878,N_19709);
and UO_159 (O_159,N_19822,N_19798);
or UO_160 (O_160,N_19813,N_19767);
nand UO_161 (O_161,N_19636,N_19781);
xor UO_162 (O_162,N_19796,N_19695);
and UO_163 (O_163,N_19541,N_19604);
or UO_164 (O_164,N_19811,N_19987);
nand UO_165 (O_165,N_19860,N_19641);
nor UO_166 (O_166,N_19654,N_19761);
nor UO_167 (O_167,N_19687,N_19557);
and UO_168 (O_168,N_19954,N_19899);
or UO_169 (O_169,N_19967,N_19503);
or UO_170 (O_170,N_19598,N_19858);
nand UO_171 (O_171,N_19973,N_19744);
nor UO_172 (O_172,N_19599,N_19537);
or UO_173 (O_173,N_19734,N_19972);
nor UO_174 (O_174,N_19959,N_19580);
nor UO_175 (O_175,N_19653,N_19738);
or UO_176 (O_176,N_19673,N_19737);
nor UO_177 (O_177,N_19932,N_19838);
or UO_178 (O_178,N_19515,N_19953);
nor UO_179 (O_179,N_19743,N_19584);
nor UO_180 (O_180,N_19594,N_19880);
nand UO_181 (O_181,N_19567,N_19992);
nand UO_182 (O_182,N_19867,N_19958);
and UO_183 (O_183,N_19884,N_19774);
nand UO_184 (O_184,N_19841,N_19926);
and UO_185 (O_185,N_19793,N_19827);
and UO_186 (O_186,N_19975,N_19749);
and UO_187 (O_187,N_19693,N_19998);
or UO_188 (O_188,N_19933,N_19978);
and UO_189 (O_189,N_19697,N_19578);
nand UO_190 (O_190,N_19772,N_19601);
nor UO_191 (O_191,N_19877,N_19716);
and UO_192 (O_192,N_19964,N_19929);
and UO_193 (O_193,N_19923,N_19683);
nor UO_194 (O_194,N_19914,N_19524);
nand UO_195 (O_195,N_19801,N_19575);
nand UO_196 (O_196,N_19824,N_19707);
and UO_197 (O_197,N_19836,N_19627);
nor UO_198 (O_198,N_19685,N_19778);
and UO_199 (O_199,N_19938,N_19576);
nor UO_200 (O_200,N_19952,N_19804);
xnor UO_201 (O_201,N_19688,N_19786);
nand UO_202 (O_202,N_19645,N_19666);
or UO_203 (O_203,N_19720,N_19622);
and UO_204 (O_204,N_19747,N_19549);
or UO_205 (O_205,N_19574,N_19600);
nand UO_206 (O_206,N_19885,N_19663);
nand UO_207 (O_207,N_19724,N_19886);
nor UO_208 (O_208,N_19547,N_19905);
and UO_209 (O_209,N_19722,N_19900);
nand UO_210 (O_210,N_19562,N_19554);
xor UO_211 (O_211,N_19903,N_19970);
or UO_212 (O_212,N_19984,N_19638);
and UO_213 (O_213,N_19855,N_19531);
nand UO_214 (O_214,N_19981,N_19961);
or UO_215 (O_215,N_19617,N_19674);
xnor UO_216 (O_216,N_19837,N_19996);
and UO_217 (O_217,N_19845,N_19609);
nor UO_218 (O_218,N_19943,N_19690);
and UO_219 (O_219,N_19571,N_19924);
xor UO_220 (O_220,N_19703,N_19912);
or UO_221 (O_221,N_19566,N_19890);
or UO_222 (O_222,N_19735,N_19968);
nor UO_223 (O_223,N_19572,N_19847);
nand UO_224 (O_224,N_19564,N_19920);
xnor UO_225 (O_225,N_19748,N_19865);
and UO_226 (O_226,N_19799,N_19872);
xnor UO_227 (O_227,N_19579,N_19530);
or UO_228 (O_228,N_19906,N_19642);
nor UO_229 (O_229,N_19966,N_19812);
or UO_230 (O_230,N_19615,N_19946);
nor UO_231 (O_231,N_19640,N_19589);
nand UO_232 (O_232,N_19676,N_19667);
and UO_233 (O_233,N_19701,N_19595);
or UO_234 (O_234,N_19657,N_19832);
xor UO_235 (O_235,N_19704,N_19889);
or UO_236 (O_236,N_19711,N_19548);
nor UO_237 (O_237,N_19593,N_19814);
nor UO_238 (O_238,N_19639,N_19891);
and UO_239 (O_239,N_19652,N_19794);
or UO_240 (O_240,N_19951,N_19678);
nor UO_241 (O_241,N_19939,N_19582);
nor UO_242 (O_242,N_19602,N_19718);
and UO_243 (O_243,N_19671,N_19648);
and UO_244 (O_244,N_19715,N_19936);
nor UO_245 (O_245,N_19513,N_19908);
nor UO_246 (O_246,N_19561,N_19546);
or UO_247 (O_247,N_19763,N_19542);
or UO_248 (O_248,N_19773,N_19868);
xor UO_249 (O_249,N_19876,N_19692);
or UO_250 (O_250,N_19777,N_19586);
xor UO_251 (O_251,N_19878,N_19590);
and UO_252 (O_252,N_19677,N_19590);
nor UO_253 (O_253,N_19692,N_19886);
xor UO_254 (O_254,N_19794,N_19831);
nor UO_255 (O_255,N_19508,N_19636);
nor UO_256 (O_256,N_19704,N_19965);
and UO_257 (O_257,N_19533,N_19660);
nor UO_258 (O_258,N_19765,N_19754);
nor UO_259 (O_259,N_19899,N_19537);
nand UO_260 (O_260,N_19974,N_19814);
or UO_261 (O_261,N_19671,N_19688);
nor UO_262 (O_262,N_19699,N_19843);
or UO_263 (O_263,N_19971,N_19544);
or UO_264 (O_264,N_19743,N_19631);
xor UO_265 (O_265,N_19620,N_19737);
nand UO_266 (O_266,N_19843,N_19683);
and UO_267 (O_267,N_19843,N_19514);
or UO_268 (O_268,N_19854,N_19644);
and UO_269 (O_269,N_19776,N_19652);
xnor UO_270 (O_270,N_19740,N_19963);
and UO_271 (O_271,N_19945,N_19795);
nor UO_272 (O_272,N_19891,N_19987);
nand UO_273 (O_273,N_19907,N_19994);
nor UO_274 (O_274,N_19680,N_19629);
or UO_275 (O_275,N_19595,N_19929);
nor UO_276 (O_276,N_19827,N_19893);
or UO_277 (O_277,N_19984,N_19764);
nor UO_278 (O_278,N_19880,N_19583);
and UO_279 (O_279,N_19774,N_19706);
and UO_280 (O_280,N_19584,N_19741);
or UO_281 (O_281,N_19510,N_19555);
and UO_282 (O_282,N_19694,N_19626);
or UO_283 (O_283,N_19902,N_19818);
and UO_284 (O_284,N_19680,N_19890);
and UO_285 (O_285,N_19525,N_19849);
nor UO_286 (O_286,N_19631,N_19931);
nand UO_287 (O_287,N_19639,N_19681);
or UO_288 (O_288,N_19842,N_19912);
or UO_289 (O_289,N_19522,N_19645);
nor UO_290 (O_290,N_19526,N_19915);
nor UO_291 (O_291,N_19547,N_19598);
nor UO_292 (O_292,N_19916,N_19749);
and UO_293 (O_293,N_19766,N_19983);
or UO_294 (O_294,N_19599,N_19774);
or UO_295 (O_295,N_19917,N_19568);
and UO_296 (O_296,N_19870,N_19948);
and UO_297 (O_297,N_19791,N_19747);
and UO_298 (O_298,N_19957,N_19877);
nor UO_299 (O_299,N_19702,N_19632);
xor UO_300 (O_300,N_19674,N_19940);
and UO_301 (O_301,N_19775,N_19719);
and UO_302 (O_302,N_19571,N_19563);
nand UO_303 (O_303,N_19656,N_19756);
nor UO_304 (O_304,N_19596,N_19882);
nor UO_305 (O_305,N_19875,N_19605);
nand UO_306 (O_306,N_19989,N_19822);
nand UO_307 (O_307,N_19705,N_19732);
nand UO_308 (O_308,N_19703,N_19546);
and UO_309 (O_309,N_19712,N_19866);
xor UO_310 (O_310,N_19728,N_19875);
xor UO_311 (O_311,N_19977,N_19654);
nor UO_312 (O_312,N_19865,N_19982);
and UO_313 (O_313,N_19614,N_19593);
nor UO_314 (O_314,N_19523,N_19544);
nor UO_315 (O_315,N_19732,N_19794);
nand UO_316 (O_316,N_19813,N_19728);
and UO_317 (O_317,N_19652,N_19596);
nor UO_318 (O_318,N_19978,N_19969);
or UO_319 (O_319,N_19701,N_19807);
and UO_320 (O_320,N_19835,N_19627);
and UO_321 (O_321,N_19681,N_19772);
or UO_322 (O_322,N_19636,N_19558);
and UO_323 (O_323,N_19539,N_19571);
nand UO_324 (O_324,N_19747,N_19518);
or UO_325 (O_325,N_19609,N_19902);
nand UO_326 (O_326,N_19906,N_19660);
and UO_327 (O_327,N_19735,N_19742);
and UO_328 (O_328,N_19703,N_19878);
and UO_329 (O_329,N_19663,N_19723);
nand UO_330 (O_330,N_19568,N_19880);
nor UO_331 (O_331,N_19801,N_19855);
nor UO_332 (O_332,N_19736,N_19813);
nand UO_333 (O_333,N_19700,N_19772);
nor UO_334 (O_334,N_19739,N_19919);
or UO_335 (O_335,N_19593,N_19973);
nand UO_336 (O_336,N_19534,N_19504);
nand UO_337 (O_337,N_19834,N_19671);
and UO_338 (O_338,N_19824,N_19768);
or UO_339 (O_339,N_19669,N_19906);
nor UO_340 (O_340,N_19766,N_19545);
nor UO_341 (O_341,N_19671,N_19731);
xnor UO_342 (O_342,N_19730,N_19985);
and UO_343 (O_343,N_19788,N_19589);
nor UO_344 (O_344,N_19979,N_19850);
nor UO_345 (O_345,N_19801,N_19589);
or UO_346 (O_346,N_19975,N_19573);
nand UO_347 (O_347,N_19874,N_19753);
nor UO_348 (O_348,N_19969,N_19637);
and UO_349 (O_349,N_19661,N_19764);
nor UO_350 (O_350,N_19830,N_19577);
or UO_351 (O_351,N_19723,N_19923);
or UO_352 (O_352,N_19532,N_19593);
nand UO_353 (O_353,N_19727,N_19726);
nand UO_354 (O_354,N_19740,N_19981);
and UO_355 (O_355,N_19864,N_19689);
nor UO_356 (O_356,N_19704,N_19778);
and UO_357 (O_357,N_19504,N_19505);
nor UO_358 (O_358,N_19987,N_19989);
or UO_359 (O_359,N_19729,N_19738);
nand UO_360 (O_360,N_19783,N_19538);
and UO_361 (O_361,N_19646,N_19606);
and UO_362 (O_362,N_19553,N_19782);
and UO_363 (O_363,N_19962,N_19724);
nor UO_364 (O_364,N_19752,N_19886);
or UO_365 (O_365,N_19765,N_19541);
or UO_366 (O_366,N_19782,N_19627);
nand UO_367 (O_367,N_19985,N_19600);
and UO_368 (O_368,N_19832,N_19523);
or UO_369 (O_369,N_19844,N_19799);
nand UO_370 (O_370,N_19863,N_19807);
nor UO_371 (O_371,N_19563,N_19668);
or UO_372 (O_372,N_19613,N_19829);
nand UO_373 (O_373,N_19742,N_19836);
or UO_374 (O_374,N_19721,N_19894);
or UO_375 (O_375,N_19804,N_19854);
or UO_376 (O_376,N_19967,N_19739);
nor UO_377 (O_377,N_19529,N_19969);
nand UO_378 (O_378,N_19961,N_19586);
or UO_379 (O_379,N_19776,N_19955);
nor UO_380 (O_380,N_19610,N_19563);
or UO_381 (O_381,N_19908,N_19671);
xor UO_382 (O_382,N_19896,N_19581);
nand UO_383 (O_383,N_19767,N_19823);
nand UO_384 (O_384,N_19620,N_19720);
nand UO_385 (O_385,N_19717,N_19913);
nor UO_386 (O_386,N_19595,N_19557);
or UO_387 (O_387,N_19878,N_19950);
nor UO_388 (O_388,N_19569,N_19600);
nand UO_389 (O_389,N_19925,N_19838);
nand UO_390 (O_390,N_19506,N_19504);
xor UO_391 (O_391,N_19798,N_19738);
or UO_392 (O_392,N_19869,N_19604);
nor UO_393 (O_393,N_19761,N_19833);
nand UO_394 (O_394,N_19566,N_19854);
nand UO_395 (O_395,N_19775,N_19684);
or UO_396 (O_396,N_19508,N_19683);
nand UO_397 (O_397,N_19879,N_19524);
nor UO_398 (O_398,N_19613,N_19914);
or UO_399 (O_399,N_19756,N_19538);
xnor UO_400 (O_400,N_19995,N_19669);
nand UO_401 (O_401,N_19541,N_19844);
nor UO_402 (O_402,N_19938,N_19658);
or UO_403 (O_403,N_19634,N_19618);
and UO_404 (O_404,N_19867,N_19581);
and UO_405 (O_405,N_19912,N_19797);
or UO_406 (O_406,N_19687,N_19646);
nand UO_407 (O_407,N_19686,N_19836);
and UO_408 (O_408,N_19775,N_19516);
and UO_409 (O_409,N_19885,N_19502);
and UO_410 (O_410,N_19794,N_19670);
nand UO_411 (O_411,N_19573,N_19728);
and UO_412 (O_412,N_19828,N_19655);
or UO_413 (O_413,N_19801,N_19914);
nor UO_414 (O_414,N_19511,N_19547);
or UO_415 (O_415,N_19913,N_19698);
or UO_416 (O_416,N_19785,N_19996);
nor UO_417 (O_417,N_19785,N_19729);
or UO_418 (O_418,N_19878,N_19895);
and UO_419 (O_419,N_19597,N_19622);
xor UO_420 (O_420,N_19538,N_19510);
and UO_421 (O_421,N_19728,N_19735);
nand UO_422 (O_422,N_19948,N_19860);
xnor UO_423 (O_423,N_19601,N_19782);
nand UO_424 (O_424,N_19941,N_19880);
or UO_425 (O_425,N_19930,N_19908);
and UO_426 (O_426,N_19955,N_19675);
xor UO_427 (O_427,N_19665,N_19601);
xnor UO_428 (O_428,N_19951,N_19601);
nor UO_429 (O_429,N_19691,N_19689);
or UO_430 (O_430,N_19582,N_19775);
or UO_431 (O_431,N_19736,N_19741);
or UO_432 (O_432,N_19784,N_19575);
or UO_433 (O_433,N_19924,N_19535);
or UO_434 (O_434,N_19648,N_19530);
nand UO_435 (O_435,N_19571,N_19721);
and UO_436 (O_436,N_19690,N_19951);
or UO_437 (O_437,N_19856,N_19861);
nand UO_438 (O_438,N_19534,N_19529);
and UO_439 (O_439,N_19997,N_19905);
or UO_440 (O_440,N_19583,N_19621);
nor UO_441 (O_441,N_19958,N_19612);
nand UO_442 (O_442,N_19881,N_19571);
nand UO_443 (O_443,N_19528,N_19840);
nor UO_444 (O_444,N_19899,N_19909);
or UO_445 (O_445,N_19738,N_19934);
xor UO_446 (O_446,N_19674,N_19596);
nand UO_447 (O_447,N_19647,N_19994);
or UO_448 (O_448,N_19830,N_19788);
nand UO_449 (O_449,N_19925,N_19519);
or UO_450 (O_450,N_19946,N_19712);
and UO_451 (O_451,N_19707,N_19871);
nand UO_452 (O_452,N_19681,N_19932);
or UO_453 (O_453,N_19589,N_19632);
and UO_454 (O_454,N_19519,N_19546);
nor UO_455 (O_455,N_19977,N_19744);
nand UO_456 (O_456,N_19937,N_19834);
nor UO_457 (O_457,N_19538,N_19801);
nand UO_458 (O_458,N_19979,N_19645);
or UO_459 (O_459,N_19771,N_19817);
nor UO_460 (O_460,N_19797,N_19839);
nand UO_461 (O_461,N_19711,N_19856);
nand UO_462 (O_462,N_19616,N_19758);
nand UO_463 (O_463,N_19867,N_19714);
nand UO_464 (O_464,N_19674,N_19651);
nor UO_465 (O_465,N_19600,N_19788);
and UO_466 (O_466,N_19751,N_19558);
nand UO_467 (O_467,N_19666,N_19974);
nand UO_468 (O_468,N_19689,N_19709);
xnor UO_469 (O_469,N_19686,N_19507);
nor UO_470 (O_470,N_19896,N_19595);
nand UO_471 (O_471,N_19583,N_19750);
and UO_472 (O_472,N_19857,N_19958);
xor UO_473 (O_473,N_19999,N_19704);
or UO_474 (O_474,N_19746,N_19519);
nand UO_475 (O_475,N_19697,N_19693);
nand UO_476 (O_476,N_19819,N_19876);
nand UO_477 (O_477,N_19708,N_19802);
nand UO_478 (O_478,N_19796,N_19671);
or UO_479 (O_479,N_19779,N_19850);
nor UO_480 (O_480,N_19988,N_19781);
nand UO_481 (O_481,N_19678,N_19995);
nor UO_482 (O_482,N_19675,N_19781);
nand UO_483 (O_483,N_19765,N_19559);
xnor UO_484 (O_484,N_19684,N_19578);
nor UO_485 (O_485,N_19838,N_19660);
or UO_486 (O_486,N_19814,N_19748);
nor UO_487 (O_487,N_19855,N_19836);
or UO_488 (O_488,N_19801,N_19996);
or UO_489 (O_489,N_19720,N_19805);
and UO_490 (O_490,N_19676,N_19678);
nand UO_491 (O_491,N_19973,N_19935);
nor UO_492 (O_492,N_19921,N_19777);
or UO_493 (O_493,N_19930,N_19873);
nand UO_494 (O_494,N_19544,N_19787);
xnor UO_495 (O_495,N_19999,N_19961);
and UO_496 (O_496,N_19753,N_19775);
nand UO_497 (O_497,N_19666,N_19562);
and UO_498 (O_498,N_19933,N_19802);
and UO_499 (O_499,N_19666,N_19540);
nand UO_500 (O_500,N_19575,N_19713);
nand UO_501 (O_501,N_19534,N_19641);
xnor UO_502 (O_502,N_19678,N_19513);
nand UO_503 (O_503,N_19937,N_19788);
nor UO_504 (O_504,N_19833,N_19617);
and UO_505 (O_505,N_19779,N_19585);
nand UO_506 (O_506,N_19511,N_19505);
nand UO_507 (O_507,N_19522,N_19571);
or UO_508 (O_508,N_19519,N_19930);
and UO_509 (O_509,N_19747,N_19534);
and UO_510 (O_510,N_19738,N_19959);
nand UO_511 (O_511,N_19635,N_19864);
nand UO_512 (O_512,N_19670,N_19781);
and UO_513 (O_513,N_19673,N_19670);
or UO_514 (O_514,N_19692,N_19518);
nand UO_515 (O_515,N_19861,N_19915);
or UO_516 (O_516,N_19980,N_19869);
nor UO_517 (O_517,N_19690,N_19987);
nor UO_518 (O_518,N_19748,N_19945);
nor UO_519 (O_519,N_19976,N_19616);
and UO_520 (O_520,N_19569,N_19760);
nand UO_521 (O_521,N_19896,N_19709);
or UO_522 (O_522,N_19907,N_19863);
and UO_523 (O_523,N_19781,N_19911);
and UO_524 (O_524,N_19925,N_19993);
or UO_525 (O_525,N_19792,N_19830);
or UO_526 (O_526,N_19514,N_19662);
nand UO_527 (O_527,N_19570,N_19826);
xor UO_528 (O_528,N_19964,N_19595);
and UO_529 (O_529,N_19686,N_19803);
and UO_530 (O_530,N_19681,N_19568);
or UO_531 (O_531,N_19749,N_19682);
nand UO_532 (O_532,N_19930,N_19994);
nor UO_533 (O_533,N_19623,N_19739);
and UO_534 (O_534,N_19818,N_19509);
and UO_535 (O_535,N_19929,N_19594);
xor UO_536 (O_536,N_19785,N_19621);
xnor UO_537 (O_537,N_19737,N_19733);
nor UO_538 (O_538,N_19658,N_19556);
nor UO_539 (O_539,N_19933,N_19822);
or UO_540 (O_540,N_19586,N_19903);
nor UO_541 (O_541,N_19739,N_19952);
nand UO_542 (O_542,N_19670,N_19865);
xor UO_543 (O_543,N_19560,N_19721);
nor UO_544 (O_544,N_19589,N_19979);
and UO_545 (O_545,N_19826,N_19508);
and UO_546 (O_546,N_19559,N_19732);
and UO_547 (O_547,N_19988,N_19742);
nor UO_548 (O_548,N_19717,N_19872);
nand UO_549 (O_549,N_19834,N_19657);
and UO_550 (O_550,N_19880,N_19758);
or UO_551 (O_551,N_19700,N_19669);
or UO_552 (O_552,N_19861,N_19988);
nand UO_553 (O_553,N_19881,N_19912);
or UO_554 (O_554,N_19731,N_19815);
or UO_555 (O_555,N_19674,N_19539);
nor UO_556 (O_556,N_19644,N_19557);
or UO_557 (O_557,N_19503,N_19517);
nand UO_558 (O_558,N_19571,N_19895);
nand UO_559 (O_559,N_19896,N_19597);
nand UO_560 (O_560,N_19841,N_19994);
xor UO_561 (O_561,N_19520,N_19724);
nor UO_562 (O_562,N_19906,N_19610);
and UO_563 (O_563,N_19795,N_19692);
or UO_564 (O_564,N_19820,N_19809);
nand UO_565 (O_565,N_19622,N_19811);
and UO_566 (O_566,N_19645,N_19832);
xnor UO_567 (O_567,N_19809,N_19958);
nand UO_568 (O_568,N_19814,N_19933);
or UO_569 (O_569,N_19666,N_19767);
or UO_570 (O_570,N_19626,N_19527);
nor UO_571 (O_571,N_19721,N_19973);
and UO_572 (O_572,N_19520,N_19882);
and UO_573 (O_573,N_19752,N_19768);
and UO_574 (O_574,N_19824,N_19571);
or UO_575 (O_575,N_19801,N_19569);
nand UO_576 (O_576,N_19644,N_19930);
and UO_577 (O_577,N_19904,N_19552);
nand UO_578 (O_578,N_19660,N_19513);
and UO_579 (O_579,N_19665,N_19785);
nand UO_580 (O_580,N_19972,N_19796);
nor UO_581 (O_581,N_19977,N_19707);
nor UO_582 (O_582,N_19748,N_19861);
xnor UO_583 (O_583,N_19648,N_19718);
or UO_584 (O_584,N_19798,N_19532);
and UO_585 (O_585,N_19729,N_19560);
nand UO_586 (O_586,N_19670,N_19746);
and UO_587 (O_587,N_19894,N_19555);
nor UO_588 (O_588,N_19683,N_19665);
or UO_589 (O_589,N_19954,N_19911);
and UO_590 (O_590,N_19869,N_19572);
and UO_591 (O_591,N_19662,N_19612);
and UO_592 (O_592,N_19621,N_19574);
nor UO_593 (O_593,N_19840,N_19605);
nor UO_594 (O_594,N_19647,N_19501);
or UO_595 (O_595,N_19584,N_19868);
or UO_596 (O_596,N_19678,N_19957);
and UO_597 (O_597,N_19564,N_19811);
nor UO_598 (O_598,N_19659,N_19686);
nor UO_599 (O_599,N_19528,N_19979);
and UO_600 (O_600,N_19976,N_19797);
nor UO_601 (O_601,N_19929,N_19513);
or UO_602 (O_602,N_19576,N_19631);
or UO_603 (O_603,N_19582,N_19820);
nand UO_604 (O_604,N_19809,N_19765);
nand UO_605 (O_605,N_19813,N_19811);
xnor UO_606 (O_606,N_19739,N_19710);
and UO_607 (O_607,N_19515,N_19813);
nor UO_608 (O_608,N_19831,N_19850);
nand UO_609 (O_609,N_19700,N_19735);
or UO_610 (O_610,N_19530,N_19915);
nor UO_611 (O_611,N_19623,N_19961);
nand UO_612 (O_612,N_19561,N_19782);
nor UO_613 (O_613,N_19905,N_19754);
nand UO_614 (O_614,N_19880,N_19786);
or UO_615 (O_615,N_19955,N_19893);
xor UO_616 (O_616,N_19870,N_19538);
and UO_617 (O_617,N_19961,N_19916);
nand UO_618 (O_618,N_19955,N_19631);
nand UO_619 (O_619,N_19686,N_19791);
nand UO_620 (O_620,N_19973,N_19694);
xor UO_621 (O_621,N_19578,N_19777);
nor UO_622 (O_622,N_19503,N_19723);
nand UO_623 (O_623,N_19814,N_19573);
nand UO_624 (O_624,N_19728,N_19550);
nand UO_625 (O_625,N_19513,N_19759);
nand UO_626 (O_626,N_19932,N_19783);
and UO_627 (O_627,N_19923,N_19515);
or UO_628 (O_628,N_19593,N_19718);
and UO_629 (O_629,N_19773,N_19880);
nor UO_630 (O_630,N_19675,N_19626);
nor UO_631 (O_631,N_19915,N_19908);
or UO_632 (O_632,N_19651,N_19675);
nor UO_633 (O_633,N_19638,N_19615);
nand UO_634 (O_634,N_19621,N_19561);
and UO_635 (O_635,N_19528,N_19674);
nor UO_636 (O_636,N_19781,N_19587);
nor UO_637 (O_637,N_19900,N_19635);
or UO_638 (O_638,N_19716,N_19572);
or UO_639 (O_639,N_19747,N_19883);
and UO_640 (O_640,N_19668,N_19905);
or UO_641 (O_641,N_19691,N_19947);
or UO_642 (O_642,N_19968,N_19633);
nand UO_643 (O_643,N_19965,N_19711);
nor UO_644 (O_644,N_19856,N_19543);
or UO_645 (O_645,N_19598,N_19809);
or UO_646 (O_646,N_19911,N_19719);
nand UO_647 (O_647,N_19777,N_19787);
nor UO_648 (O_648,N_19974,N_19614);
or UO_649 (O_649,N_19504,N_19844);
nand UO_650 (O_650,N_19730,N_19627);
nand UO_651 (O_651,N_19718,N_19591);
nand UO_652 (O_652,N_19547,N_19938);
nand UO_653 (O_653,N_19591,N_19684);
and UO_654 (O_654,N_19879,N_19978);
nand UO_655 (O_655,N_19537,N_19692);
or UO_656 (O_656,N_19990,N_19955);
and UO_657 (O_657,N_19944,N_19653);
and UO_658 (O_658,N_19580,N_19922);
nand UO_659 (O_659,N_19696,N_19903);
or UO_660 (O_660,N_19741,N_19899);
nand UO_661 (O_661,N_19727,N_19859);
and UO_662 (O_662,N_19864,N_19781);
xor UO_663 (O_663,N_19816,N_19592);
and UO_664 (O_664,N_19792,N_19942);
and UO_665 (O_665,N_19522,N_19701);
nand UO_666 (O_666,N_19770,N_19644);
and UO_667 (O_667,N_19790,N_19867);
nor UO_668 (O_668,N_19729,N_19853);
and UO_669 (O_669,N_19518,N_19803);
and UO_670 (O_670,N_19926,N_19617);
or UO_671 (O_671,N_19904,N_19632);
nand UO_672 (O_672,N_19816,N_19715);
or UO_673 (O_673,N_19719,N_19588);
and UO_674 (O_674,N_19865,N_19825);
xnor UO_675 (O_675,N_19753,N_19687);
xor UO_676 (O_676,N_19956,N_19780);
or UO_677 (O_677,N_19754,N_19873);
nand UO_678 (O_678,N_19803,N_19746);
nor UO_679 (O_679,N_19887,N_19514);
or UO_680 (O_680,N_19713,N_19725);
and UO_681 (O_681,N_19641,N_19890);
and UO_682 (O_682,N_19825,N_19944);
and UO_683 (O_683,N_19582,N_19734);
and UO_684 (O_684,N_19635,N_19937);
nand UO_685 (O_685,N_19693,N_19663);
nand UO_686 (O_686,N_19884,N_19545);
or UO_687 (O_687,N_19857,N_19591);
or UO_688 (O_688,N_19625,N_19939);
and UO_689 (O_689,N_19845,N_19597);
or UO_690 (O_690,N_19868,N_19534);
nand UO_691 (O_691,N_19898,N_19862);
nor UO_692 (O_692,N_19931,N_19799);
nor UO_693 (O_693,N_19852,N_19980);
and UO_694 (O_694,N_19700,N_19838);
or UO_695 (O_695,N_19743,N_19961);
and UO_696 (O_696,N_19824,N_19845);
xnor UO_697 (O_697,N_19827,N_19511);
and UO_698 (O_698,N_19948,N_19782);
or UO_699 (O_699,N_19954,N_19688);
and UO_700 (O_700,N_19515,N_19597);
xnor UO_701 (O_701,N_19575,N_19921);
or UO_702 (O_702,N_19581,N_19617);
nor UO_703 (O_703,N_19757,N_19654);
and UO_704 (O_704,N_19876,N_19866);
and UO_705 (O_705,N_19785,N_19899);
or UO_706 (O_706,N_19781,N_19531);
or UO_707 (O_707,N_19543,N_19506);
nor UO_708 (O_708,N_19863,N_19828);
nor UO_709 (O_709,N_19545,N_19727);
nand UO_710 (O_710,N_19966,N_19848);
xnor UO_711 (O_711,N_19998,N_19807);
nor UO_712 (O_712,N_19901,N_19596);
xor UO_713 (O_713,N_19758,N_19595);
nand UO_714 (O_714,N_19809,N_19973);
nor UO_715 (O_715,N_19814,N_19775);
xor UO_716 (O_716,N_19875,N_19854);
nor UO_717 (O_717,N_19831,N_19813);
nand UO_718 (O_718,N_19676,N_19509);
nand UO_719 (O_719,N_19902,N_19618);
or UO_720 (O_720,N_19513,N_19698);
nand UO_721 (O_721,N_19578,N_19855);
nor UO_722 (O_722,N_19833,N_19570);
nand UO_723 (O_723,N_19673,N_19868);
or UO_724 (O_724,N_19657,N_19632);
or UO_725 (O_725,N_19750,N_19539);
and UO_726 (O_726,N_19599,N_19986);
xnor UO_727 (O_727,N_19514,N_19581);
and UO_728 (O_728,N_19579,N_19575);
or UO_729 (O_729,N_19776,N_19713);
and UO_730 (O_730,N_19911,N_19838);
or UO_731 (O_731,N_19779,N_19890);
nor UO_732 (O_732,N_19741,N_19765);
and UO_733 (O_733,N_19766,N_19561);
nor UO_734 (O_734,N_19598,N_19527);
or UO_735 (O_735,N_19988,N_19729);
and UO_736 (O_736,N_19956,N_19727);
and UO_737 (O_737,N_19800,N_19808);
or UO_738 (O_738,N_19537,N_19592);
nor UO_739 (O_739,N_19761,N_19947);
nand UO_740 (O_740,N_19740,N_19666);
or UO_741 (O_741,N_19739,N_19757);
nor UO_742 (O_742,N_19625,N_19692);
xor UO_743 (O_743,N_19948,N_19990);
nand UO_744 (O_744,N_19920,N_19965);
or UO_745 (O_745,N_19527,N_19608);
or UO_746 (O_746,N_19820,N_19613);
or UO_747 (O_747,N_19644,N_19874);
nor UO_748 (O_748,N_19610,N_19924);
nor UO_749 (O_749,N_19747,N_19832);
xor UO_750 (O_750,N_19943,N_19670);
nor UO_751 (O_751,N_19539,N_19645);
xor UO_752 (O_752,N_19743,N_19589);
nor UO_753 (O_753,N_19999,N_19702);
nand UO_754 (O_754,N_19891,N_19644);
and UO_755 (O_755,N_19768,N_19683);
nand UO_756 (O_756,N_19961,N_19670);
nor UO_757 (O_757,N_19512,N_19835);
or UO_758 (O_758,N_19602,N_19777);
nand UO_759 (O_759,N_19647,N_19818);
nor UO_760 (O_760,N_19715,N_19556);
and UO_761 (O_761,N_19885,N_19956);
nand UO_762 (O_762,N_19657,N_19755);
and UO_763 (O_763,N_19750,N_19950);
xor UO_764 (O_764,N_19995,N_19772);
nand UO_765 (O_765,N_19536,N_19855);
nand UO_766 (O_766,N_19567,N_19561);
or UO_767 (O_767,N_19663,N_19947);
xnor UO_768 (O_768,N_19688,N_19545);
nor UO_769 (O_769,N_19739,N_19686);
nor UO_770 (O_770,N_19647,N_19802);
nor UO_771 (O_771,N_19736,N_19984);
nor UO_772 (O_772,N_19761,N_19671);
nand UO_773 (O_773,N_19574,N_19909);
nor UO_774 (O_774,N_19519,N_19936);
or UO_775 (O_775,N_19895,N_19998);
or UO_776 (O_776,N_19688,N_19826);
nand UO_777 (O_777,N_19968,N_19944);
or UO_778 (O_778,N_19523,N_19893);
nor UO_779 (O_779,N_19856,N_19922);
and UO_780 (O_780,N_19699,N_19934);
xnor UO_781 (O_781,N_19760,N_19911);
and UO_782 (O_782,N_19515,N_19780);
nor UO_783 (O_783,N_19757,N_19628);
xor UO_784 (O_784,N_19889,N_19571);
nor UO_785 (O_785,N_19632,N_19775);
and UO_786 (O_786,N_19579,N_19625);
or UO_787 (O_787,N_19743,N_19780);
nand UO_788 (O_788,N_19539,N_19515);
nand UO_789 (O_789,N_19737,N_19969);
or UO_790 (O_790,N_19596,N_19701);
nand UO_791 (O_791,N_19784,N_19692);
nand UO_792 (O_792,N_19827,N_19723);
nand UO_793 (O_793,N_19570,N_19517);
nor UO_794 (O_794,N_19879,N_19581);
xnor UO_795 (O_795,N_19656,N_19904);
or UO_796 (O_796,N_19938,N_19885);
and UO_797 (O_797,N_19661,N_19714);
xnor UO_798 (O_798,N_19614,N_19769);
or UO_799 (O_799,N_19927,N_19945);
and UO_800 (O_800,N_19980,N_19730);
or UO_801 (O_801,N_19855,N_19631);
or UO_802 (O_802,N_19829,N_19949);
nor UO_803 (O_803,N_19525,N_19999);
and UO_804 (O_804,N_19612,N_19954);
nor UO_805 (O_805,N_19819,N_19803);
or UO_806 (O_806,N_19746,N_19572);
or UO_807 (O_807,N_19824,N_19682);
nor UO_808 (O_808,N_19907,N_19815);
or UO_809 (O_809,N_19789,N_19968);
xor UO_810 (O_810,N_19925,N_19865);
or UO_811 (O_811,N_19816,N_19504);
nand UO_812 (O_812,N_19514,N_19785);
or UO_813 (O_813,N_19965,N_19824);
nor UO_814 (O_814,N_19985,N_19825);
xor UO_815 (O_815,N_19956,N_19947);
and UO_816 (O_816,N_19547,N_19871);
and UO_817 (O_817,N_19598,N_19641);
nand UO_818 (O_818,N_19527,N_19979);
or UO_819 (O_819,N_19587,N_19958);
and UO_820 (O_820,N_19944,N_19624);
or UO_821 (O_821,N_19963,N_19624);
xor UO_822 (O_822,N_19920,N_19529);
or UO_823 (O_823,N_19742,N_19699);
nand UO_824 (O_824,N_19898,N_19793);
nand UO_825 (O_825,N_19865,N_19556);
nand UO_826 (O_826,N_19562,N_19980);
or UO_827 (O_827,N_19825,N_19811);
nand UO_828 (O_828,N_19569,N_19636);
nand UO_829 (O_829,N_19930,N_19548);
nor UO_830 (O_830,N_19954,N_19544);
nor UO_831 (O_831,N_19976,N_19767);
or UO_832 (O_832,N_19521,N_19671);
and UO_833 (O_833,N_19969,N_19789);
and UO_834 (O_834,N_19994,N_19629);
and UO_835 (O_835,N_19824,N_19758);
xor UO_836 (O_836,N_19971,N_19501);
xnor UO_837 (O_837,N_19710,N_19962);
nor UO_838 (O_838,N_19691,N_19706);
xor UO_839 (O_839,N_19614,N_19584);
xnor UO_840 (O_840,N_19560,N_19974);
or UO_841 (O_841,N_19598,N_19870);
nand UO_842 (O_842,N_19776,N_19858);
and UO_843 (O_843,N_19805,N_19671);
and UO_844 (O_844,N_19708,N_19502);
nand UO_845 (O_845,N_19691,N_19500);
nor UO_846 (O_846,N_19570,N_19588);
nand UO_847 (O_847,N_19737,N_19887);
nand UO_848 (O_848,N_19995,N_19910);
xor UO_849 (O_849,N_19962,N_19637);
nor UO_850 (O_850,N_19543,N_19724);
and UO_851 (O_851,N_19903,N_19958);
nand UO_852 (O_852,N_19535,N_19882);
nand UO_853 (O_853,N_19621,N_19886);
or UO_854 (O_854,N_19900,N_19889);
nand UO_855 (O_855,N_19979,N_19572);
xnor UO_856 (O_856,N_19825,N_19693);
or UO_857 (O_857,N_19540,N_19824);
and UO_858 (O_858,N_19967,N_19943);
and UO_859 (O_859,N_19696,N_19524);
or UO_860 (O_860,N_19560,N_19916);
nor UO_861 (O_861,N_19721,N_19796);
nand UO_862 (O_862,N_19682,N_19710);
nand UO_863 (O_863,N_19944,N_19922);
or UO_864 (O_864,N_19845,N_19861);
nor UO_865 (O_865,N_19719,N_19561);
nand UO_866 (O_866,N_19823,N_19614);
nand UO_867 (O_867,N_19817,N_19603);
and UO_868 (O_868,N_19719,N_19644);
or UO_869 (O_869,N_19748,N_19712);
nand UO_870 (O_870,N_19908,N_19833);
nor UO_871 (O_871,N_19801,N_19813);
nor UO_872 (O_872,N_19980,N_19728);
and UO_873 (O_873,N_19980,N_19837);
nor UO_874 (O_874,N_19858,N_19832);
nor UO_875 (O_875,N_19893,N_19536);
nand UO_876 (O_876,N_19558,N_19694);
xor UO_877 (O_877,N_19846,N_19554);
or UO_878 (O_878,N_19733,N_19616);
and UO_879 (O_879,N_19589,N_19519);
and UO_880 (O_880,N_19539,N_19685);
and UO_881 (O_881,N_19570,N_19568);
xor UO_882 (O_882,N_19536,N_19577);
nand UO_883 (O_883,N_19986,N_19801);
nor UO_884 (O_884,N_19752,N_19826);
and UO_885 (O_885,N_19564,N_19863);
nand UO_886 (O_886,N_19737,N_19660);
nor UO_887 (O_887,N_19986,N_19708);
nand UO_888 (O_888,N_19832,N_19843);
nor UO_889 (O_889,N_19643,N_19682);
and UO_890 (O_890,N_19944,N_19901);
nand UO_891 (O_891,N_19828,N_19932);
or UO_892 (O_892,N_19691,N_19870);
and UO_893 (O_893,N_19838,N_19973);
nor UO_894 (O_894,N_19531,N_19980);
or UO_895 (O_895,N_19746,N_19880);
or UO_896 (O_896,N_19621,N_19810);
nand UO_897 (O_897,N_19722,N_19672);
nand UO_898 (O_898,N_19683,N_19620);
or UO_899 (O_899,N_19994,N_19803);
and UO_900 (O_900,N_19724,N_19712);
or UO_901 (O_901,N_19637,N_19837);
xor UO_902 (O_902,N_19504,N_19943);
or UO_903 (O_903,N_19720,N_19893);
nand UO_904 (O_904,N_19814,N_19776);
or UO_905 (O_905,N_19588,N_19846);
and UO_906 (O_906,N_19545,N_19990);
or UO_907 (O_907,N_19586,N_19953);
nor UO_908 (O_908,N_19609,N_19882);
nor UO_909 (O_909,N_19685,N_19633);
nor UO_910 (O_910,N_19622,N_19571);
or UO_911 (O_911,N_19844,N_19733);
nand UO_912 (O_912,N_19562,N_19648);
and UO_913 (O_913,N_19989,N_19747);
nand UO_914 (O_914,N_19982,N_19525);
nor UO_915 (O_915,N_19640,N_19921);
nor UO_916 (O_916,N_19708,N_19741);
nor UO_917 (O_917,N_19658,N_19987);
and UO_918 (O_918,N_19535,N_19792);
nor UO_919 (O_919,N_19870,N_19796);
nor UO_920 (O_920,N_19866,N_19952);
or UO_921 (O_921,N_19798,N_19599);
xnor UO_922 (O_922,N_19984,N_19990);
or UO_923 (O_923,N_19651,N_19798);
or UO_924 (O_924,N_19741,N_19656);
nand UO_925 (O_925,N_19606,N_19513);
or UO_926 (O_926,N_19701,N_19887);
nand UO_927 (O_927,N_19736,N_19833);
nor UO_928 (O_928,N_19844,N_19930);
or UO_929 (O_929,N_19836,N_19892);
and UO_930 (O_930,N_19668,N_19639);
and UO_931 (O_931,N_19630,N_19500);
xor UO_932 (O_932,N_19508,N_19679);
nor UO_933 (O_933,N_19756,N_19858);
or UO_934 (O_934,N_19898,N_19765);
or UO_935 (O_935,N_19710,N_19776);
nor UO_936 (O_936,N_19593,N_19855);
or UO_937 (O_937,N_19885,N_19733);
nor UO_938 (O_938,N_19570,N_19777);
and UO_939 (O_939,N_19695,N_19646);
or UO_940 (O_940,N_19970,N_19901);
and UO_941 (O_941,N_19586,N_19908);
nand UO_942 (O_942,N_19914,N_19815);
or UO_943 (O_943,N_19527,N_19823);
and UO_944 (O_944,N_19511,N_19990);
nand UO_945 (O_945,N_19996,N_19968);
nor UO_946 (O_946,N_19714,N_19552);
and UO_947 (O_947,N_19930,N_19890);
xor UO_948 (O_948,N_19701,N_19569);
nor UO_949 (O_949,N_19589,N_19730);
nor UO_950 (O_950,N_19588,N_19836);
nand UO_951 (O_951,N_19651,N_19892);
nor UO_952 (O_952,N_19757,N_19960);
or UO_953 (O_953,N_19791,N_19711);
xnor UO_954 (O_954,N_19622,N_19924);
or UO_955 (O_955,N_19578,N_19905);
nor UO_956 (O_956,N_19742,N_19588);
and UO_957 (O_957,N_19679,N_19864);
and UO_958 (O_958,N_19814,N_19590);
or UO_959 (O_959,N_19865,N_19707);
and UO_960 (O_960,N_19752,N_19974);
nor UO_961 (O_961,N_19663,N_19591);
nor UO_962 (O_962,N_19771,N_19934);
or UO_963 (O_963,N_19896,N_19913);
nand UO_964 (O_964,N_19655,N_19823);
or UO_965 (O_965,N_19884,N_19560);
nor UO_966 (O_966,N_19951,N_19821);
or UO_967 (O_967,N_19695,N_19881);
nor UO_968 (O_968,N_19914,N_19954);
nand UO_969 (O_969,N_19752,N_19809);
and UO_970 (O_970,N_19783,N_19799);
nand UO_971 (O_971,N_19926,N_19697);
and UO_972 (O_972,N_19588,N_19531);
and UO_973 (O_973,N_19814,N_19665);
and UO_974 (O_974,N_19621,N_19995);
and UO_975 (O_975,N_19578,N_19860);
nand UO_976 (O_976,N_19533,N_19707);
and UO_977 (O_977,N_19689,N_19783);
or UO_978 (O_978,N_19627,N_19510);
or UO_979 (O_979,N_19709,N_19665);
or UO_980 (O_980,N_19534,N_19970);
and UO_981 (O_981,N_19629,N_19763);
nand UO_982 (O_982,N_19913,N_19811);
nand UO_983 (O_983,N_19844,N_19994);
xnor UO_984 (O_984,N_19634,N_19753);
or UO_985 (O_985,N_19550,N_19617);
nand UO_986 (O_986,N_19864,N_19760);
or UO_987 (O_987,N_19568,N_19668);
xnor UO_988 (O_988,N_19878,N_19968);
or UO_989 (O_989,N_19910,N_19946);
xnor UO_990 (O_990,N_19822,N_19742);
xnor UO_991 (O_991,N_19572,N_19580);
nand UO_992 (O_992,N_19606,N_19883);
or UO_993 (O_993,N_19874,N_19861);
or UO_994 (O_994,N_19710,N_19529);
nor UO_995 (O_995,N_19719,N_19931);
and UO_996 (O_996,N_19650,N_19994);
and UO_997 (O_997,N_19865,N_19819);
or UO_998 (O_998,N_19689,N_19640);
and UO_999 (O_999,N_19662,N_19509);
or UO_1000 (O_1000,N_19635,N_19717);
and UO_1001 (O_1001,N_19558,N_19807);
and UO_1002 (O_1002,N_19710,N_19658);
and UO_1003 (O_1003,N_19684,N_19891);
xor UO_1004 (O_1004,N_19664,N_19763);
nor UO_1005 (O_1005,N_19586,N_19881);
and UO_1006 (O_1006,N_19759,N_19971);
or UO_1007 (O_1007,N_19787,N_19972);
and UO_1008 (O_1008,N_19993,N_19861);
nor UO_1009 (O_1009,N_19528,N_19649);
nor UO_1010 (O_1010,N_19799,N_19843);
nand UO_1011 (O_1011,N_19586,N_19990);
nor UO_1012 (O_1012,N_19733,N_19963);
nand UO_1013 (O_1013,N_19708,N_19604);
nand UO_1014 (O_1014,N_19851,N_19896);
nand UO_1015 (O_1015,N_19599,N_19581);
nand UO_1016 (O_1016,N_19923,N_19758);
and UO_1017 (O_1017,N_19829,N_19507);
nor UO_1018 (O_1018,N_19727,N_19952);
or UO_1019 (O_1019,N_19713,N_19515);
nand UO_1020 (O_1020,N_19926,N_19886);
nand UO_1021 (O_1021,N_19584,N_19943);
xnor UO_1022 (O_1022,N_19848,N_19870);
and UO_1023 (O_1023,N_19738,N_19643);
nand UO_1024 (O_1024,N_19773,N_19632);
nand UO_1025 (O_1025,N_19716,N_19529);
nor UO_1026 (O_1026,N_19870,N_19710);
nor UO_1027 (O_1027,N_19623,N_19838);
nand UO_1028 (O_1028,N_19884,N_19810);
and UO_1029 (O_1029,N_19916,N_19886);
and UO_1030 (O_1030,N_19639,N_19602);
nand UO_1031 (O_1031,N_19670,N_19648);
nand UO_1032 (O_1032,N_19877,N_19868);
nand UO_1033 (O_1033,N_19663,N_19603);
or UO_1034 (O_1034,N_19892,N_19720);
or UO_1035 (O_1035,N_19930,N_19978);
and UO_1036 (O_1036,N_19898,N_19850);
xnor UO_1037 (O_1037,N_19717,N_19804);
nor UO_1038 (O_1038,N_19967,N_19616);
and UO_1039 (O_1039,N_19918,N_19653);
and UO_1040 (O_1040,N_19798,N_19513);
and UO_1041 (O_1041,N_19858,N_19946);
or UO_1042 (O_1042,N_19714,N_19562);
nand UO_1043 (O_1043,N_19792,N_19765);
nand UO_1044 (O_1044,N_19958,N_19907);
xor UO_1045 (O_1045,N_19524,N_19669);
and UO_1046 (O_1046,N_19547,N_19630);
and UO_1047 (O_1047,N_19921,N_19806);
or UO_1048 (O_1048,N_19953,N_19906);
or UO_1049 (O_1049,N_19746,N_19978);
nor UO_1050 (O_1050,N_19759,N_19706);
nor UO_1051 (O_1051,N_19665,N_19820);
xor UO_1052 (O_1052,N_19837,N_19997);
nor UO_1053 (O_1053,N_19617,N_19731);
or UO_1054 (O_1054,N_19975,N_19872);
or UO_1055 (O_1055,N_19713,N_19693);
nor UO_1056 (O_1056,N_19762,N_19514);
and UO_1057 (O_1057,N_19658,N_19962);
and UO_1058 (O_1058,N_19834,N_19913);
or UO_1059 (O_1059,N_19612,N_19568);
or UO_1060 (O_1060,N_19625,N_19600);
nor UO_1061 (O_1061,N_19651,N_19939);
nand UO_1062 (O_1062,N_19588,N_19614);
and UO_1063 (O_1063,N_19922,N_19816);
nor UO_1064 (O_1064,N_19993,N_19803);
xor UO_1065 (O_1065,N_19619,N_19932);
or UO_1066 (O_1066,N_19946,N_19918);
or UO_1067 (O_1067,N_19827,N_19888);
nor UO_1068 (O_1068,N_19838,N_19972);
or UO_1069 (O_1069,N_19898,N_19726);
nand UO_1070 (O_1070,N_19958,N_19991);
xnor UO_1071 (O_1071,N_19763,N_19983);
nor UO_1072 (O_1072,N_19847,N_19900);
or UO_1073 (O_1073,N_19802,N_19506);
or UO_1074 (O_1074,N_19535,N_19877);
and UO_1075 (O_1075,N_19860,N_19843);
and UO_1076 (O_1076,N_19977,N_19877);
and UO_1077 (O_1077,N_19571,N_19978);
nand UO_1078 (O_1078,N_19763,N_19760);
and UO_1079 (O_1079,N_19568,N_19504);
and UO_1080 (O_1080,N_19862,N_19921);
or UO_1081 (O_1081,N_19814,N_19767);
nand UO_1082 (O_1082,N_19894,N_19734);
and UO_1083 (O_1083,N_19798,N_19561);
nand UO_1084 (O_1084,N_19748,N_19792);
xnor UO_1085 (O_1085,N_19553,N_19907);
and UO_1086 (O_1086,N_19520,N_19620);
or UO_1087 (O_1087,N_19861,N_19611);
nor UO_1088 (O_1088,N_19766,N_19777);
and UO_1089 (O_1089,N_19600,N_19521);
or UO_1090 (O_1090,N_19617,N_19707);
or UO_1091 (O_1091,N_19784,N_19991);
or UO_1092 (O_1092,N_19539,N_19696);
or UO_1093 (O_1093,N_19920,N_19575);
or UO_1094 (O_1094,N_19584,N_19560);
nand UO_1095 (O_1095,N_19621,N_19508);
or UO_1096 (O_1096,N_19891,N_19887);
and UO_1097 (O_1097,N_19552,N_19920);
or UO_1098 (O_1098,N_19571,N_19590);
nand UO_1099 (O_1099,N_19639,N_19949);
and UO_1100 (O_1100,N_19516,N_19866);
or UO_1101 (O_1101,N_19875,N_19502);
nor UO_1102 (O_1102,N_19606,N_19927);
or UO_1103 (O_1103,N_19874,N_19833);
and UO_1104 (O_1104,N_19686,N_19896);
nand UO_1105 (O_1105,N_19754,N_19822);
or UO_1106 (O_1106,N_19513,N_19872);
nor UO_1107 (O_1107,N_19830,N_19893);
nand UO_1108 (O_1108,N_19808,N_19552);
xnor UO_1109 (O_1109,N_19984,N_19693);
nor UO_1110 (O_1110,N_19603,N_19894);
or UO_1111 (O_1111,N_19992,N_19741);
or UO_1112 (O_1112,N_19570,N_19569);
nand UO_1113 (O_1113,N_19788,N_19761);
and UO_1114 (O_1114,N_19802,N_19783);
or UO_1115 (O_1115,N_19597,N_19692);
or UO_1116 (O_1116,N_19920,N_19533);
and UO_1117 (O_1117,N_19739,N_19837);
or UO_1118 (O_1118,N_19685,N_19552);
nor UO_1119 (O_1119,N_19625,N_19673);
nand UO_1120 (O_1120,N_19516,N_19733);
or UO_1121 (O_1121,N_19963,N_19890);
or UO_1122 (O_1122,N_19873,N_19572);
nor UO_1123 (O_1123,N_19544,N_19669);
and UO_1124 (O_1124,N_19943,N_19755);
and UO_1125 (O_1125,N_19727,N_19941);
nor UO_1126 (O_1126,N_19645,N_19883);
or UO_1127 (O_1127,N_19593,N_19556);
or UO_1128 (O_1128,N_19819,N_19591);
nand UO_1129 (O_1129,N_19909,N_19701);
and UO_1130 (O_1130,N_19754,N_19536);
or UO_1131 (O_1131,N_19604,N_19632);
or UO_1132 (O_1132,N_19662,N_19666);
xor UO_1133 (O_1133,N_19847,N_19706);
nor UO_1134 (O_1134,N_19732,N_19555);
or UO_1135 (O_1135,N_19644,N_19833);
and UO_1136 (O_1136,N_19680,N_19955);
xor UO_1137 (O_1137,N_19991,N_19840);
and UO_1138 (O_1138,N_19579,N_19582);
nand UO_1139 (O_1139,N_19825,N_19987);
and UO_1140 (O_1140,N_19811,N_19735);
and UO_1141 (O_1141,N_19905,N_19925);
or UO_1142 (O_1142,N_19529,N_19992);
nor UO_1143 (O_1143,N_19799,N_19779);
and UO_1144 (O_1144,N_19699,N_19802);
or UO_1145 (O_1145,N_19911,N_19873);
or UO_1146 (O_1146,N_19796,N_19687);
xnor UO_1147 (O_1147,N_19921,N_19509);
and UO_1148 (O_1148,N_19596,N_19972);
and UO_1149 (O_1149,N_19600,N_19969);
nor UO_1150 (O_1150,N_19592,N_19791);
xnor UO_1151 (O_1151,N_19816,N_19833);
nor UO_1152 (O_1152,N_19695,N_19746);
nand UO_1153 (O_1153,N_19826,N_19738);
and UO_1154 (O_1154,N_19610,N_19904);
nand UO_1155 (O_1155,N_19933,N_19610);
or UO_1156 (O_1156,N_19623,N_19635);
nor UO_1157 (O_1157,N_19730,N_19734);
and UO_1158 (O_1158,N_19723,N_19557);
nor UO_1159 (O_1159,N_19903,N_19523);
xnor UO_1160 (O_1160,N_19979,N_19642);
or UO_1161 (O_1161,N_19692,N_19797);
nand UO_1162 (O_1162,N_19547,N_19987);
or UO_1163 (O_1163,N_19610,N_19686);
and UO_1164 (O_1164,N_19510,N_19516);
nor UO_1165 (O_1165,N_19815,N_19840);
or UO_1166 (O_1166,N_19997,N_19936);
nor UO_1167 (O_1167,N_19637,N_19788);
nor UO_1168 (O_1168,N_19951,N_19563);
or UO_1169 (O_1169,N_19819,N_19920);
and UO_1170 (O_1170,N_19979,N_19740);
nor UO_1171 (O_1171,N_19943,N_19777);
or UO_1172 (O_1172,N_19547,N_19650);
and UO_1173 (O_1173,N_19734,N_19844);
xor UO_1174 (O_1174,N_19693,N_19596);
or UO_1175 (O_1175,N_19794,N_19511);
nand UO_1176 (O_1176,N_19587,N_19956);
and UO_1177 (O_1177,N_19507,N_19521);
and UO_1178 (O_1178,N_19829,N_19752);
nor UO_1179 (O_1179,N_19663,N_19718);
and UO_1180 (O_1180,N_19717,N_19809);
or UO_1181 (O_1181,N_19509,N_19945);
nand UO_1182 (O_1182,N_19802,N_19938);
nor UO_1183 (O_1183,N_19896,N_19945);
nor UO_1184 (O_1184,N_19990,N_19805);
nor UO_1185 (O_1185,N_19705,N_19624);
xnor UO_1186 (O_1186,N_19771,N_19572);
nor UO_1187 (O_1187,N_19889,N_19785);
nor UO_1188 (O_1188,N_19822,N_19631);
or UO_1189 (O_1189,N_19912,N_19917);
xnor UO_1190 (O_1190,N_19522,N_19886);
nand UO_1191 (O_1191,N_19548,N_19644);
and UO_1192 (O_1192,N_19611,N_19931);
or UO_1193 (O_1193,N_19666,N_19973);
and UO_1194 (O_1194,N_19716,N_19675);
or UO_1195 (O_1195,N_19908,N_19595);
or UO_1196 (O_1196,N_19913,N_19582);
nor UO_1197 (O_1197,N_19788,N_19731);
or UO_1198 (O_1198,N_19609,N_19549);
nor UO_1199 (O_1199,N_19501,N_19995);
xnor UO_1200 (O_1200,N_19558,N_19704);
and UO_1201 (O_1201,N_19706,N_19638);
and UO_1202 (O_1202,N_19775,N_19791);
or UO_1203 (O_1203,N_19879,N_19940);
or UO_1204 (O_1204,N_19643,N_19826);
and UO_1205 (O_1205,N_19936,N_19594);
and UO_1206 (O_1206,N_19940,N_19977);
nand UO_1207 (O_1207,N_19697,N_19918);
and UO_1208 (O_1208,N_19947,N_19905);
and UO_1209 (O_1209,N_19879,N_19561);
and UO_1210 (O_1210,N_19811,N_19591);
nand UO_1211 (O_1211,N_19846,N_19700);
nor UO_1212 (O_1212,N_19788,N_19820);
nand UO_1213 (O_1213,N_19629,N_19934);
or UO_1214 (O_1214,N_19503,N_19887);
and UO_1215 (O_1215,N_19795,N_19837);
or UO_1216 (O_1216,N_19812,N_19627);
or UO_1217 (O_1217,N_19790,N_19772);
nor UO_1218 (O_1218,N_19970,N_19849);
xor UO_1219 (O_1219,N_19940,N_19556);
and UO_1220 (O_1220,N_19691,N_19973);
or UO_1221 (O_1221,N_19755,N_19947);
nand UO_1222 (O_1222,N_19939,N_19544);
nor UO_1223 (O_1223,N_19855,N_19669);
nor UO_1224 (O_1224,N_19823,N_19979);
nand UO_1225 (O_1225,N_19611,N_19592);
nand UO_1226 (O_1226,N_19713,N_19889);
or UO_1227 (O_1227,N_19673,N_19618);
and UO_1228 (O_1228,N_19733,N_19788);
or UO_1229 (O_1229,N_19862,N_19916);
xor UO_1230 (O_1230,N_19787,N_19695);
nor UO_1231 (O_1231,N_19531,N_19996);
or UO_1232 (O_1232,N_19748,N_19784);
nand UO_1233 (O_1233,N_19873,N_19923);
nor UO_1234 (O_1234,N_19881,N_19817);
and UO_1235 (O_1235,N_19672,N_19744);
or UO_1236 (O_1236,N_19537,N_19888);
or UO_1237 (O_1237,N_19828,N_19722);
nand UO_1238 (O_1238,N_19541,N_19643);
and UO_1239 (O_1239,N_19824,N_19812);
and UO_1240 (O_1240,N_19998,N_19870);
nor UO_1241 (O_1241,N_19797,N_19694);
and UO_1242 (O_1242,N_19595,N_19546);
or UO_1243 (O_1243,N_19573,N_19916);
nand UO_1244 (O_1244,N_19673,N_19587);
and UO_1245 (O_1245,N_19649,N_19804);
and UO_1246 (O_1246,N_19956,N_19684);
or UO_1247 (O_1247,N_19603,N_19703);
and UO_1248 (O_1248,N_19507,N_19594);
or UO_1249 (O_1249,N_19559,N_19720);
nor UO_1250 (O_1250,N_19950,N_19507);
nand UO_1251 (O_1251,N_19782,N_19915);
and UO_1252 (O_1252,N_19937,N_19709);
xnor UO_1253 (O_1253,N_19628,N_19791);
or UO_1254 (O_1254,N_19909,N_19628);
and UO_1255 (O_1255,N_19794,N_19505);
nand UO_1256 (O_1256,N_19968,N_19801);
nor UO_1257 (O_1257,N_19970,N_19827);
nor UO_1258 (O_1258,N_19937,N_19754);
xor UO_1259 (O_1259,N_19813,N_19641);
nor UO_1260 (O_1260,N_19602,N_19641);
or UO_1261 (O_1261,N_19810,N_19963);
or UO_1262 (O_1262,N_19958,N_19541);
nor UO_1263 (O_1263,N_19776,N_19972);
nor UO_1264 (O_1264,N_19992,N_19919);
and UO_1265 (O_1265,N_19977,N_19838);
nor UO_1266 (O_1266,N_19783,N_19815);
or UO_1267 (O_1267,N_19871,N_19795);
or UO_1268 (O_1268,N_19585,N_19664);
nand UO_1269 (O_1269,N_19768,N_19818);
nand UO_1270 (O_1270,N_19842,N_19776);
or UO_1271 (O_1271,N_19513,N_19525);
xor UO_1272 (O_1272,N_19686,N_19664);
nand UO_1273 (O_1273,N_19978,N_19944);
or UO_1274 (O_1274,N_19742,N_19657);
nor UO_1275 (O_1275,N_19549,N_19990);
or UO_1276 (O_1276,N_19598,N_19903);
or UO_1277 (O_1277,N_19616,N_19552);
nor UO_1278 (O_1278,N_19959,N_19814);
and UO_1279 (O_1279,N_19519,N_19509);
and UO_1280 (O_1280,N_19684,N_19666);
or UO_1281 (O_1281,N_19881,N_19816);
and UO_1282 (O_1282,N_19658,N_19660);
or UO_1283 (O_1283,N_19977,N_19593);
nor UO_1284 (O_1284,N_19502,N_19771);
or UO_1285 (O_1285,N_19887,N_19968);
and UO_1286 (O_1286,N_19932,N_19780);
xor UO_1287 (O_1287,N_19936,N_19881);
nand UO_1288 (O_1288,N_19909,N_19836);
nand UO_1289 (O_1289,N_19724,N_19912);
xor UO_1290 (O_1290,N_19711,N_19592);
nor UO_1291 (O_1291,N_19684,N_19952);
nor UO_1292 (O_1292,N_19748,N_19621);
or UO_1293 (O_1293,N_19585,N_19969);
nand UO_1294 (O_1294,N_19566,N_19821);
and UO_1295 (O_1295,N_19710,N_19986);
nor UO_1296 (O_1296,N_19536,N_19790);
and UO_1297 (O_1297,N_19527,N_19822);
and UO_1298 (O_1298,N_19926,N_19946);
and UO_1299 (O_1299,N_19620,N_19945);
nand UO_1300 (O_1300,N_19972,N_19722);
and UO_1301 (O_1301,N_19932,N_19763);
and UO_1302 (O_1302,N_19559,N_19871);
or UO_1303 (O_1303,N_19829,N_19725);
or UO_1304 (O_1304,N_19753,N_19774);
nor UO_1305 (O_1305,N_19923,N_19570);
and UO_1306 (O_1306,N_19510,N_19655);
nand UO_1307 (O_1307,N_19959,N_19932);
nor UO_1308 (O_1308,N_19703,N_19501);
or UO_1309 (O_1309,N_19721,N_19767);
nor UO_1310 (O_1310,N_19701,N_19868);
nand UO_1311 (O_1311,N_19756,N_19539);
and UO_1312 (O_1312,N_19814,N_19595);
and UO_1313 (O_1313,N_19612,N_19730);
or UO_1314 (O_1314,N_19900,N_19899);
or UO_1315 (O_1315,N_19602,N_19833);
nand UO_1316 (O_1316,N_19655,N_19598);
nor UO_1317 (O_1317,N_19964,N_19908);
nand UO_1318 (O_1318,N_19620,N_19786);
nand UO_1319 (O_1319,N_19951,N_19794);
and UO_1320 (O_1320,N_19578,N_19965);
xnor UO_1321 (O_1321,N_19884,N_19603);
or UO_1322 (O_1322,N_19995,N_19868);
and UO_1323 (O_1323,N_19501,N_19911);
nand UO_1324 (O_1324,N_19854,N_19649);
or UO_1325 (O_1325,N_19780,N_19829);
and UO_1326 (O_1326,N_19693,N_19629);
nor UO_1327 (O_1327,N_19636,N_19873);
or UO_1328 (O_1328,N_19686,N_19720);
and UO_1329 (O_1329,N_19559,N_19869);
and UO_1330 (O_1330,N_19890,N_19829);
or UO_1331 (O_1331,N_19615,N_19862);
nand UO_1332 (O_1332,N_19703,N_19629);
nand UO_1333 (O_1333,N_19895,N_19692);
nor UO_1334 (O_1334,N_19554,N_19524);
nor UO_1335 (O_1335,N_19832,N_19791);
or UO_1336 (O_1336,N_19665,N_19795);
or UO_1337 (O_1337,N_19592,N_19575);
xnor UO_1338 (O_1338,N_19557,N_19923);
nor UO_1339 (O_1339,N_19599,N_19751);
or UO_1340 (O_1340,N_19648,N_19911);
or UO_1341 (O_1341,N_19723,N_19515);
nand UO_1342 (O_1342,N_19630,N_19944);
or UO_1343 (O_1343,N_19622,N_19675);
nand UO_1344 (O_1344,N_19703,N_19747);
nand UO_1345 (O_1345,N_19943,N_19569);
nand UO_1346 (O_1346,N_19881,N_19678);
and UO_1347 (O_1347,N_19595,N_19554);
nand UO_1348 (O_1348,N_19962,N_19536);
nand UO_1349 (O_1349,N_19991,N_19687);
or UO_1350 (O_1350,N_19920,N_19962);
and UO_1351 (O_1351,N_19920,N_19576);
and UO_1352 (O_1352,N_19981,N_19877);
and UO_1353 (O_1353,N_19550,N_19801);
and UO_1354 (O_1354,N_19629,N_19696);
and UO_1355 (O_1355,N_19640,N_19660);
nor UO_1356 (O_1356,N_19562,N_19662);
xnor UO_1357 (O_1357,N_19996,N_19953);
nor UO_1358 (O_1358,N_19977,N_19705);
or UO_1359 (O_1359,N_19978,N_19501);
nor UO_1360 (O_1360,N_19774,N_19981);
xnor UO_1361 (O_1361,N_19827,N_19617);
or UO_1362 (O_1362,N_19973,N_19817);
nor UO_1363 (O_1363,N_19827,N_19751);
xnor UO_1364 (O_1364,N_19582,N_19888);
or UO_1365 (O_1365,N_19792,N_19680);
nor UO_1366 (O_1366,N_19832,N_19618);
or UO_1367 (O_1367,N_19653,N_19569);
and UO_1368 (O_1368,N_19986,N_19899);
nand UO_1369 (O_1369,N_19844,N_19918);
xor UO_1370 (O_1370,N_19761,N_19624);
nor UO_1371 (O_1371,N_19660,N_19789);
and UO_1372 (O_1372,N_19870,N_19818);
xor UO_1373 (O_1373,N_19875,N_19748);
or UO_1374 (O_1374,N_19569,N_19604);
nand UO_1375 (O_1375,N_19802,N_19675);
nand UO_1376 (O_1376,N_19613,N_19823);
and UO_1377 (O_1377,N_19515,N_19852);
and UO_1378 (O_1378,N_19921,N_19997);
nor UO_1379 (O_1379,N_19954,N_19546);
and UO_1380 (O_1380,N_19698,N_19911);
or UO_1381 (O_1381,N_19755,N_19763);
nand UO_1382 (O_1382,N_19505,N_19674);
nor UO_1383 (O_1383,N_19898,N_19652);
or UO_1384 (O_1384,N_19597,N_19892);
and UO_1385 (O_1385,N_19599,N_19785);
nor UO_1386 (O_1386,N_19514,N_19894);
or UO_1387 (O_1387,N_19800,N_19801);
or UO_1388 (O_1388,N_19728,N_19748);
nor UO_1389 (O_1389,N_19858,N_19698);
and UO_1390 (O_1390,N_19793,N_19643);
or UO_1391 (O_1391,N_19637,N_19830);
nand UO_1392 (O_1392,N_19974,N_19630);
and UO_1393 (O_1393,N_19829,N_19962);
nand UO_1394 (O_1394,N_19844,N_19724);
xnor UO_1395 (O_1395,N_19674,N_19816);
or UO_1396 (O_1396,N_19646,N_19678);
and UO_1397 (O_1397,N_19651,N_19993);
or UO_1398 (O_1398,N_19778,N_19780);
and UO_1399 (O_1399,N_19818,N_19719);
or UO_1400 (O_1400,N_19668,N_19781);
xnor UO_1401 (O_1401,N_19957,N_19537);
nor UO_1402 (O_1402,N_19840,N_19759);
and UO_1403 (O_1403,N_19590,N_19599);
nor UO_1404 (O_1404,N_19734,N_19976);
nand UO_1405 (O_1405,N_19928,N_19708);
or UO_1406 (O_1406,N_19687,N_19982);
or UO_1407 (O_1407,N_19616,N_19634);
and UO_1408 (O_1408,N_19889,N_19710);
or UO_1409 (O_1409,N_19565,N_19688);
nor UO_1410 (O_1410,N_19644,N_19790);
nand UO_1411 (O_1411,N_19630,N_19767);
or UO_1412 (O_1412,N_19918,N_19749);
nor UO_1413 (O_1413,N_19706,N_19732);
and UO_1414 (O_1414,N_19973,N_19876);
or UO_1415 (O_1415,N_19745,N_19737);
nor UO_1416 (O_1416,N_19573,N_19943);
xor UO_1417 (O_1417,N_19832,N_19955);
and UO_1418 (O_1418,N_19526,N_19906);
nor UO_1419 (O_1419,N_19670,N_19710);
nor UO_1420 (O_1420,N_19715,N_19582);
nor UO_1421 (O_1421,N_19565,N_19896);
or UO_1422 (O_1422,N_19845,N_19551);
xnor UO_1423 (O_1423,N_19975,N_19763);
nand UO_1424 (O_1424,N_19731,N_19790);
or UO_1425 (O_1425,N_19885,N_19973);
and UO_1426 (O_1426,N_19728,N_19903);
nand UO_1427 (O_1427,N_19695,N_19902);
or UO_1428 (O_1428,N_19660,N_19527);
nand UO_1429 (O_1429,N_19782,N_19909);
nand UO_1430 (O_1430,N_19822,N_19613);
nand UO_1431 (O_1431,N_19786,N_19820);
or UO_1432 (O_1432,N_19520,N_19769);
nor UO_1433 (O_1433,N_19703,N_19576);
nand UO_1434 (O_1434,N_19929,N_19569);
nor UO_1435 (O_1435,N_19742,N_19734);
nor UO_1436 (O_1436,N_19515,N_19940);
nand UO_1437 (O_1437,N_19550,N_19856);
xnor UO_1438 (O_1438,N_19789,N_19609);
nand UO_1439 (O_1439,N_19909,N_19612);
nand UO_1440 (O_1440,N_19628,N_19519);
xnor UO_1441 (O_1441,N_19766,N_19652);
and UO_1442 (O_1442,N_19911,N_19938);
and UO_1443 (O_1443,N_19747,N_19501);
nor UO_1444 (O_1444,N_19840,N_19923);
xor UO_1445 (O_1445,N_19661,N_19686);
or UO_1446 (O_1446,N_19880,N_19625);
nand UO_1447 (O_1447,N_19525,N_19725);
and UO_1448 (O_1448,N_19648,N_19903);
xnor UO_1449 (O_1449,N_19991,N_19834);
and UO_1450 (O_1450,N_19534,N_19622);
nand UO_1451 (O_1451,N_19578,N_19800);
and UO_1452 (O_1452,N_19838,N_19979);
nor UO_1453 (O_1453,N_19810,N_19803);
nand UO_1454 (O_1454,N_19552,N_19584);
xor UO_1455 (O_1455,N_19701,N_19752);
nand UO_1456 (O_1456,N_19678,N_19642);
nor UO_1457 (O_1457,N_19838,N_19918);
and UO_1458 (O_1458,N_19814,N_19856);
nor UO_1459 (O_1459,N_19964,N_19668);
and UO_1460 (O_1460,N_19552,N_19579);
nor UO_1461 (O_1461,N_19930,N_19527);
nand UO_1462 (O_1462,N_19751,N_19984);
xor UO_1463 (O_1463,N_19616,N_19765);
or UO_1464 (O_1464,N_19547,N_19751);
nand UO_1465 (O_1465,N_19789,N_19938);
nor UO_1466 (O_1466,N_19831,N_19525);
nor UO_1467 (O_1467,N_19593,N_19940);
or UO_1468 (O_1468,N_19939,N_19895);
nand UO_1469 (O_1469,N_19511,N_19810);
and UO_1470 (O_1470,N_19580,N_19883);
and UO_1471 (O_1471,N_19668,N_19947);
and UO_1472 (O_1472,N_19618,N_19542);
nor UO_1473 (O_1473,N_19750,N_19827);
and UO_1474 (O_1474,N_19525,N_19701);
xnor UO_1475 (O_1475,N_19527,N_19595);
xnor UO_1476 (O_1476,N_19597,N_19858);
nand UO_1477 (O_1477,N_19573,N_19998);
nand UO_1478 (O_1478,N_19681,N_19894);
nor UO_1479 (O_1479,N_19771,N_19649);
xor UO_1480 (O_1480,N_19670,N_19965);
or UO_1481 (O_1481,N_19527,N_19751);
nor UO_1482 (O_1482,N_19584,N_19530);
or UO_1483 (O_1483,N_19748,N_19783);
nand UO_1484 (O_1484,N_19811,N_19632);
nor UO_1485 (O_1485,N_19714,N_19846);
nand UO_1486 (O_1486,N_19650,N_19815);
or UO_1487 (O_1487,N_19535,N_19976);
or UO_1488 (O_1488,N_19847,N_19659);
xnor UO_1489 (O_1489,N_19730,N_19707);
or UO_1490 (O_1490,N_19977,N_19530);
and UO_1491 (O_1491,N_19623,N_19698);
or UO_1492 (O_1492,N_19879,N_19580);
and UO_1493 (O_1493,N_19567,N_19622);
nor UO_1494 (O_1494,N_19947,N_19560);
or UO_1495 (O_1495,N_19731,N_19993);
nor UO_1496 (O_1496,N_19952,N_19895);
and UO_1497 (O_1497,N_19915,N_19550);
or UO_1498 (O_1498,N_19971,N_19733);
nand UO_1499 (O_1499,N_19561,N_19704);
nor UO_1500 (O_1500,N_19728,N_19894);
or UO_1501 (O_1501,N_19919,N_19852);
or UO_1502 (O_1502,N_19719,N_19638);
nor UO_1503 (O_1503,N_19811,N_19531);
nor UO_1504 (O_1504,N_19818,N_19677);
nand UO_1505 (O_1505,N_19959,N_19669);
and UO_1506 (O_1506,N_19866,N_19720);
and UO_1507 (O_1507,N_19975,N_19577);
nand UO_1508 (O_1508,N_19524,N_19762);
xnor UO_1509 (O_1509,N_19831,N_19645);
or UO_1510 (O_1510,N_19871,N_19619);
xnor UO_1511 (O_1511,N_19672,N_19715);
nand UO_1512 (O_1512,N_19562,N_19509);
xnor UO_1513 (O_1513,N_19630,N_19958);
nor UO_1514 (O_1514,N_19816,N_19918);
nand UO_1515 (O_1515,N_19710,N_19743);
and UO_1516 (O_1516,N_19628,N_19802);
nand UO_1517 (O_1517,N_19657,N_19668);
or UO_1518 (O_1518,N_19770,N_19882);
and UO_1519 (O_1519,N_19553,N_19871);
and UO_1520 (O_1520,N_19714,N_19588);
nor UO_1521 (O_1521,N_19920,N_19590);
nor UO_1522 (O_1522,N_19711,N_19786);
xnor UO_1523 (O_1523,N_19694,N_19621);
nand UO_1524 (O_1524,N_19751,N_19917);
or UO_1525 (O_1525,N_19510,N_19909);
xnor UO_1526 (O_1526,N_19715,N_19821);
and UO_1527 (O_1527,N_19928,N_19632);
nor UO_1528 (O_1528,N_19850,N_19893);
nor UO_1529 (O_1529,N_19864,N_19916);
xnor UO_1530 (O_1530,N_19607,N_19744);
and UO_1531 (O_1531,N_19757,N_19673);
xor UO_1532 (O_1532,N_19848,N_19863);
nor UO_1533 (O_1533,N_19874,N_19757);
or UO_1534 (O_1534,N_19881,N_19675);
nand UO_1535 (O_1535,N_19649,N_19748);
or UO_1536 (O_1536,N_19563,N_19651);
nor UO_1537 (O_1537,N_19804,N_19793);
or UO_1538 (O_1538,N_19602,N_19930);
nand UO_1539 (O_1539,N_19794,N_19646);
and UO_1540 (O_1540,N_19549,N_19630);
xnor UO_1541 (O_1541,N_19687,N_19587);
or UO_1542 (O_1542,N_19525,N_19510);
nand UO_1543 (O_1543,N_19841,N_19887);
or UO_1544 (O_1544,N_19559,N_19700);
nor UO_1545 (O_1545,N_19737,N_19530);
nor UO_1546 (O_1546,N_19666,N_19926);
nor UO_1547 (O_1547,N_19639,N_19779);
xnor UO_1548 (O_1548,N_19802,N_19549);
or UO_1549 (O_1549,N_19729,N_19862);
nor UO_1550 (O_1550,N_19618,N_19862);
nor UO_1551 (O_1551,N_19842,N_19777);
and UO_1552 (O_1552,N_19540,N_19621);
or UO_1553 (O_1553,N_19590,N_19655);
and UO_1554 (O_1554,N_19750,N_19912);
nand UO_1555 (O_1555,N_19919,N_19627);
or UO_1556 (O_1556,N_19714,N_19508);
nand UO_1557 (O_1557,N_19975,N_19871);
and UO_1558 (O_1558,N_19811,N_19598);
nor UO_1559 (O_1559,N_19814,N_19988);
xor UO_1560 (O_1560,N_19809,N_19604);
nand UO_1561 (O_1561,N_19933,N_19795);
or UO_1562 (O_1562,N_19667,N_19917);
nor UO_1563 (O_1563,N_19835,N_19549);
or UO_1564 (O_1564,N_19966,N_19879);
nand UO_1565 (O_1565,N_19941,N_19990);
nand UO_1566 (O_1566,N_19966,N_19653);
or UO_1567 (O_1567,N_19929,N_19523);
or UO_1568 (O_1568,N_19627,N_19988);
xor UO_1569 (O_1569,N_19676,N_19746);
nand UO_1570 (O_1570,N_19655,N_19799);
nand UO_1571 (O_1571,N_19596,N_19682);
nand UO_1572 (O_1572,N_19981,N_19859);
and UO_1573 (O_1573,N_19580,N_19520);
or UO_1574 (O_1574,N_19749,N_19706);
nor UO_1575 (O_1575,N_19582,N_19765);
xnor UO_1576 (O_1576,N_19894,N_19805);
or UO_1577 (O_1577,N_19771,N_19511);
or UO_1578 (O_1578,N_19901,N_19871);
and UO_1579 (O_1579,N_19596,N_19520);
nor UO_1580 (O_1580,N_19607,N_19799);
or UO_1581 (O_1581,N_19940,N_19880);
nand UO_1582 (O_1582,N_19707,N_19772);
and UO_1583 (O_1583,N_19727,N_19633);
nor UO_1584 (O_1584,N_19797,N_19560);
or UO_1585 (O_1585,N_19813,N_19850);
nor UO_1586 (O_1586,N_19769,N_19755);
xnor UO_1587 (O_1587,N_19709,N_19526);
or UO_1588 (O_1588,N_19941,N_19747);
nor UO_1589 (O_1589,N_19665,N_19680);
and UO_1590 (O_1590,N_19904,N_19570);
nor UO_1591 (O_1591,N_19510,N_19884);
nor UO_1592 (O_1592,N_19929,N_19657);
or UO_1593 (O_1593,N_19744,N_19586);
nor UO_1594 (O_1594,N_19974,N_19745);
and UO_1595 (O_1595,N_19586,N_19732);
nor UO_1596 (O_1596,N_19682,N_19946);
and UO_1597 (O_1597,N_19515,N_19552);
nand UO_1598 (O_1598,N_19824,N_19742);
nand UO_1599 (O_1599,N_19981,N_19939);
nand UO_1600 (O_1600,N_19603,N_19713);
or UO_1601 (O_1601,N_19650,N_19930);
nand UO_1602 (O_1602,N_19579,N_19874);
nand UO_1603 (O_1603,N_19987,N_19948);
or UO_1604 (O_1604,N_19671,N_19951);
or UO_1605 (O_1605,N_19566,N_19532);
and UO_1606 (O_1606,N_19531,N_19582);
nor UO_1607 (O_1607,N_19722,N_19802);
and UO_1608 (O_1608,N_19666,N_19661);
or UO_1609 (O_1609,N_19955,N_19803);
xnor UO_1610 (O_1610,N_19904,N_19967);
and UO_1611 (O_1611,N_19931,N_19641);
nand UO_1612 (O_1612,N_19608,N_19545);
xor UO_1613 (O_1613,N_19921,N_19722);
or UO_1614 (O_1614,N_19981,N_19923);
nand UO_1615 (O_1615,N_19664,N_19592);
nor UO_1616 (O_1616,N_19908,N_19875);
nor UO_1617 (O_1617,N_19804,N_19581);
nor UO_1618 (O_1618,N_19673,N_19738);
nor UO_1619 (O_1619,N_19568,N_19626);
nor UO_1620 (O_1620,N_19742,N_19643);
and UO_1621 (O_1621,N_19883,N_19533);
or UO_1622 (O_1622,N_19948,N_19781);
nor UO_1623 (O_1623,N_19716,N_19861);
nand UO_1624 (O_1624,N_19527,N_19879);
or UO_1625 (O_1625,N_19587,N_19607);
nor UO_1626 (O_1626,N_19786,N_19651);
nor UO_1627 (O_1627,N_19728,N_19539);
or UO_1628 (O_1628,N_19866,N_19678);
or UO_1629 (O_1629,N_19895,N_19834);
and UO_1630 (O_1630,N_19655,N_19931);
nand UO_1631 (O_1631,N_19911,N_19958);
and UO_1632 (O_1632,N_19597,N_19638);
or UO_1633 (O_1633,N_19860,N_19646);
nand UO_1634 (O_1634,N_19829,N_19993);
nor UO_1635 (O_1635,N_19816,N_19835);
nand UO_1636 (O_1636,N_19647,N_19538);
nand UO_1637 (O_1637,N_19591,N_19631);
nand UO_1638 (O_1638,N_19981,N_19869);
nor UO_1639 (O_1639,N_19680,N_19579);
nor UO_1640 (O_1640,N_19858,N_19745);
or UO_1641 (O_1641,N_19771,N_19886);
and UO_1642 (O_1642,N_19984,N_19665);
or UO_1643 (O_1643,N_19794,N_19575);
and UO_1644 (O_1644,N_19763,N_19650);
nand UO_1645 (O_1645,N_19689,N_19899);
and UO_1646 (O_1646,N_19607,N_19614);
nor UO_1647 (O_1647,N_19932,N_19792);
or UO_1648 (O_1648,N_19595,N_19877);
nor UO_1649 (O_1649,N_19994,N_19536);
nor UO_1650 (O_1650,N_19750,N_19638);
or UO_1651 (O_1651,N_19854,N_19695);
nor UO_1652 (O_1652,N_19599,N_19565);
or UO_1653 (O_1653,N_19579,N_19809);
or UO_1654 (O_1654,N_19954,N_19878);
or UO_1655 (O_1655,N_19605,N_19906);
and UO_1656 (O_1656,N_19969,N_19608);
nand UO_1657 (O_1657,N_19952,N_19594);
nand UO_1658 (O_1658,N_19890,N_19523);
nand UO_1659 (O_1659,N_19551,N_19500);
nand UO_1660 (O_1660,N_19601,N_19757);
nand UO_1661 (O_1661,N_19914,N_19980);
nor UO_1662 (O_1662,N_19671,N_19831);
nand UO_1663 (O_1663,N_19519,N_19629);
or UO_1664 (O_1664,N_19766,N_19754);
and UO_1665 (O_1665,N_19617,N_19625);
or UO_1666 (O_1666,N_19812,N_19766);
or UO_1667 (O_1667,N_19778,N_19566);
or UO_1668 (O_1668,N_19651,N_19511);
nand UO_1669 (O_1669,N_19819,N_19521);
and UO_1670 (O_1670,N_19678,N_19582);
nor UO_1671 (O_1671,N_19578,N_19778);
and UO_1672 (O_1672,N_19659,N_19932);
nand UO_1673 (O_1673,N_19708,N_19686);
nand UO_1674 (O_1674,N_19575,N_19689);
or UO_1675 (O_1675,N_19914,N_19893);
and UO_1676 (O_1676,N_19860,N_19777);
nand UO_1677 (O_1677,N_19643,N_19892);
and UO_1678 (O_1678,N_19954,N_19562);
or UO_1679 (O_1679,N_19713,N_19899);
and UO_1680 (O_1680,N_19676,N_19947);
nand UO_1681 (O_1681,N_19976,N_19930);
and UO_1682 (O_1682,N_19891,N_19626);
nor UO_1683 (O_1683,N_19891,N_19900);
nand UO_1684 (O_1684,N_19812,N_19532);
or UO_1685 (O_1685,N_19808,N_19747);
or UO_1686 (O_1686,N_19552,N_19641);
nor UO_1687 (O_1687,N_19659,N_19639);
nand UO_1688 (O_1688,N_19964,N_19716);
and UO_1689 (O_1689,N_19979,N_19640);
or UO_1690 (O_1690,N_19956,N_19622);
or UO_1691 (O_1691,N_19641,N_19589);
nand UO_1692 (O_1692,N_19916,N_19848);
or UO_1693 (O_1693,N_19783,N_19864);
nor UO_1694 (O_1694,N_19689,N_19948);
or UO_1695 (O_1695,N_19533,N_19625);
nor UO_1696 (O_1696,N_19988,N_19807);
nor UO_1697 (O_1697,N_19757,N_19729);
or UO_1698 (O_1698,N_19966,N_19850);
nor UO_1699 (O_1699,N_19973,N_19702);
xnor UO_1700 (O_1700,N_19885,N_19677);
nand UO_1701 (O_1701,N_19745,N_19580);
nand UO_1702 (O_1702,N_19884,N_19741);
or UO_1703 (O_1703,N_19531,N_19623);
or UO_1704 (O_1704,N_19987,N_19924);
and UO_1705 (O_1705,N_19699,N_19950);
or UO_1706 (O_1706,N_19608,N_19996);
and UO_1707 (O_1707,N_19654,N_19855);
xor UO_1708 (O_1708,N_19550,N_19737);
nor UO_1709 (O_1709,N_19728,N_19639);
nand UO_1710 (O_1710,N_19621,N_19848);
nor UO_1711 (O_1711,N_19867,N_19672);
nor UO_1712 (O_1712,N_19889,N_19999);
and UO_1713 (O_1713,N_19713,N_19783);
nor UO_1714 (O_1714,N_19628,N_19882);
or UO_1715 (O_1715,N_19972,N_19547);
nor UO_1716 (O_1716,N_19708,N_19583);
or UO_1717 (O_1717,N_19581,N_19629);
and UO_1718 (O_1718,N_19845,N_19503);
or UO_1719 (O_1719,N_19931,N_19854);
nand UO_1720 (O_1720,N_19996,N_19570);
nand UO_1721 (O_1721,N_19867,N_19891);
nor UO_1722 (O_1722,N_19806,N_19839);
or UO_1723 (O_1723,N_19729,N_19655);
nand UO_1724 (O_1724,N_19596,N_19599);
nor UO_1725 (O_1725,N_19751,N_19688);
nor UO_1726 (O_1726,N_19707,N_19582);
xor UO_1727 (O_1727,N_19511,N_19705);
nand UO_1728 (O_1728,N_19730,N_19756);
or UO_1729 (O_1729,N_19783,N_19842);
nor UO_1730 (O_1730,N_19722,N_19604);
nand UO_1731 (O_1731,N_19746,N_19502);
or UO_1732 (O_1732,N_19640,N_19647);
or UO_1733 (O_1733,N_19946,N_19772);
and UO_1734 (O_1734,N_19566,N_19948);
or UO_1735 (O_1735,N_19747,N_19894);
and UO_1736 (O_1736,N_19745,N_19907);
or UO_1737 (O_1737,N_19667,N_19693);
nand UO_1738 (O_1738,N_19820,N_19833);
or UO_1739 (O_1739,N_19541,N_19910);
nand UO_1740 (O_1740,N_19659,N_19593);
xor UO_1741 (O_1741,N_19987,N_19728);
xnor UO_1742 (O_1742,N_19613,N_19619);
or UO_1743 (O_1743,N_19868,N_19529);
or UO_1744 (O_1744,N_19806,N_19882);
xor UO_1745 (O_1745,N_19932,N_19563);
nand UO_1746 (O_1746,N_19520,N_19708);
nand UO_1747 (O_1747,N_19591,N_19525);
and UO_1748 (O_1748,N_19922,N_19844);
xnor UO_1749 (O_1749,N_19757,N_19952);
or UO_1750 (O_1750,N_19511,N_19533);
nand UO_1751 (O_1751,N_19593,N_19951);
and UO_1752 (O_1752,N_19883,N_19919);
or UO_1753 (O_1753,N_19876,N_19988);
or UO_1754 (O_1754,N_19950,N_19732);
nand UO_1755 (O_1755,N_19799,N_19573);
or UO_1756 (O_1756,N_19549,N_19704);
nand UO_1757 (O_1757,N_19874,N_19793);
and UO_1758 (O_1758,N_19841,N_19524);
nor UO_1759 (O_1759,N_19732,N_19900);
and UO_1760 (O_1760,N_19861,N_19550);
and UO_1761 (O_1761,N_19880,N_19809);
and UO_1762 (O_1762,N_19759,N_19644);
nand UO_1763 (O_1763,N_19542,N_19839);
nand UO_1764 (O_1764,N_19702,N_19505);
nand UO_1765 (O_1765,N_19896,N_19683);
and UO_1766 (O_1766,N_19590,N_19644);
nor UO_1767 (O_1767,N_19999,N_19828);
or UO_1768 (O_1768,N_19504,N_19743);
or UO_1769 (O_1769,N_19822,N_19737);
nor UO_1770 (O_1770,N_19574,N_19633);
and UO_1771 (O_1771,N_19553,N_19675);
and UO_1772 (O_1772,N_19709,N_19940);
nor UO_1773 (O_1773,N_19919,N_19854);
nor UO_1774 (O_1774,N_19823,N_19594);
or UO_1775 (O_1775,N_19595,N_19800);
nand UO_1776 (O_1776,N_19800,N_19609);
nand UO_1777 (O_1777,N_19769,N_19650);
nand UO_1778 (O_1778,N_19619,N_19535);
or UO_1779 (O_1779,N_19537,N_19796);
nor UO_1780 (O_1780,N_19652,N_19892);
and UO_1781 (O_1781,N_19751,N_19671);
xnor UO_1782 (O_1782,N_19930,N_19523);
or UO_1783 (O_1783,N_19759,N_19797);
or UO_1784 (O_1784,N_19902,N_19890);
and UO_1785 (O_1785,N_19554,N_19973);
xor UO_1786 (O_1786,N_19876,N_19541);
nand UO_1787 (O_1787,N_19794,N_19671);
nor UO_1788 (O_1788,N_19704,N_19845);
and UO_1789 (O_1789,N_19976,N_19638);
and UO_1790 (O_1790,N_19700,N_19827);
nor UO_1791 (O_1791,N_19763,N_19742);
nor UO_1792 (O_1792,N_19805,N_19618);
nor UO_1793 (O_1793,N_19902,N_19993);
and UO_1794 (O_1794,N_19668,N_19911);
nand UO_1795 (O_1795,N_19558,N_19608);
nand UO_1796 (O_1796,N_19854,N_19918);
or UO_1797 (O_1797,N_19806,N_19525);
nand UO_1798 (O_1798,N_19674,N_19568);
and UO_1799 (O_1799,N_19982,N_19913);
or UO_1800 (O_1800,N_19805,N_19737);
xor UO_1801 (O_1801,N_19812,N_19695);
and UO_1802 (O_1802,N_19578,N_19788);
nor UO_1803 (O_1803,N_19640,N_19784);
nor UO_1804 (O_1804,N_19567,N_19861);
xor UO_1805 (O_1805,N_19934,N_19773);
and UO_1806 (O_1806,N_19961,N_19835);
and UO_1807 (O_1807,N_19817,N_19533);
nand UO_1808 (O_1808,N_19788,N_19847);
nand UO_1809 (O_1809,N_19856,N_19695);
or UO_1810 (O_1810,N_19973,N_19708);
or UO_1811 (O_1811,N_19581,N_19582);
nand UO_1812 (O_1812,N_19913,N_19592);
nand UO_1813 (O_1813,N_19810,N_19549);
and UO_1814 (O_1814,N_19510,N_19864);
and UO_1815 (O_1815,N_19792,N_19533);
and UO_1816 (O_1816,N_19742,N_19777);
nand UO_1817 (O_1817,N_19730,N_19995);
nand UO_1818 (O_1818,N_19546,N_19621);
and UO_1819 (O_1819,N_19672,N_19677);
nor UO_1820 (O_1820,N_19931,N_19807);
nor UO_1821 (O_1821,N_19972,N_19950);
nand UO_1822 (O_1822,N_19838,N_19888);
nor UO_1823 (O_1823,N_19536,N_19753);
xor UO_1824 (O_1824,N_19798,N_19720);
nand UO_1825 (O_1825,N_19800,N_19792);
nand UO_1826 (O_1826,N_19986,N_19835);
or UO_1827 (O_1827,N_19638,N_19816);
and UO_1828 (O_1828,N_19860,N_19686);
and UO_1829 (O_1829,N_19747,N_19908);
nor UO_1830 (O_1830,N_19656,N_19977);
nor UO_1831 (O_1831,N_19604,N_19874);
or UO_1832 (O_1832,N_19519,N_19657);
nand UO_1833 (O_1833,N_19828,N_19890);
nand UO_1834 (O_1834,N_19848,N_19512);
and UO_1835 (O_1835,N_19875,N_19929);
or UO_1836 (O_1836,N_19678,N_19901);
or UO_1837 (O_1837,N_19619,N_19519);
nor UO_1838 (O_1838,N_19609,N_19828);
or UO_1839 (O_1839,N_19640,N_19788);
nor UO_1840 (O_1840,N_19731,N_19670);
or UO_1841 (O_1841,N_19965,N_19865);
and UO_1842 (O_1842,N_19940,N_19688);
or UO_1843 (O_1843,N_19740,N_19813);
nand UO_1844 (O_1844,N_19602,N_19800);
nand UO_1845 (O_1845,N_19993,N_19728);
and UO_1846 (O_1846,N_19728,N_19921);
xnor UO_1847 (O_1847,N_19567,N_19560);
or UO_1848 (O_1848,N_19903,N_19854);
or UO_1849 (O_1849,N_19729,N_19786);
and UO_1850 (O_1850,N_19972,N_19990);
nand UO_1851 (O_1851,N_19953,N_19635);
xnor UO_1852 (O_1852,N_19755,N_19952);
nor UO_1853 (O_1853,N_19907,N_19940);
or UO_1854 (O_1854,N_19749,N_19542);
xor UO_1855 (O_1855,N_19549,N_19988);
nor UO_1856 (O_1856,N_19718,N_19548);
or UO_1857 (O_1857,N_19560,N_19683);
nand UO_1858 (O_1858,N_19890,N_19506);
nor UO_1859 (O_1859,N_19935,N_19524);
or UO_1860 (O_1860,N_19869,N_19610);
or UO_1861 (O_1861,N_19866,N_19680);
or UO_1862 (O_1862,N_19516,N_19987);
nand UO_1863 (O_1863,N_19631,N_19954);
nor UO_1864 (O_1864,N_19683,N_19573);
and UO_1865 (O_1865,N_19549,N_19852);
xnor UO_1866 (O_1866,N_19831,N_19777);
or UO_1867 (O_1867,N_19588,N_19993);
nor UO_1868 (O_1868,N_19614,N_19877);
nand UO_1869 (O_1869,N_19825,N_19933);
or UO_1870 (O_1870,N_19986,N_19858);
or UO_1871 (O_1871,N_19934,N_19958);
and UO_1872 (O_1872,N_19703,N_19954);
and UO_1873 (O_1873,N_19819,N_19922);
and UO_1874 (O_1874,N_19746,N_19795);
and UO_1875 (O_1875,N_19613,N_19712);
xor UO_1876 (O_1876,N_19610,N_19983);
xnor UO_1877 (O_1877,N_19528,N_19793);
or UO_1878 (O_1878,N_19865,N_19915);
and UO_1879 (O_1879,N_19674,N_19591);
or UO_1880 (O_1880,N_19985,N_19972);
and UO_1881 (O_1881,N_19747,N_19952);
nor UO_1882 (O_1882,N_19817,N_19618);
or UO_1883 (O_1883,N_19622,N_19797);
and UO_1884 (O_1884,N_19667,N_19683);
nand UO_1885 (O_1885,N_19829,N_19926);
or UO_1886 (O_1886,N_19769,N_19941);
xnor UO_1887 (O_1887,N_19579,N_19936);
nand UO_1888 (O_1888,N_19664,N_19509);
xor UO_1889 (O_1889,N_19617,N_19968);
nand UO_1890 (O_1890,N_19791,N_19730);
nand UO_1891 (O_1891,N_19881,N_19573);
or UO_1892 (O_1892,N_19865,N_19920);
nor UO_1893 (O_1893,N_19537,N_19714);
and UO_1894 (O_1894,N_19834,N_19534);
nand UO_1895 (O_1895,N_19653,N_19568);
nor UO_1896 (O_1896,N_19916,N_19550);
nand UO_1897 (O_1897,N_19904,N_19858);
nand UO_1898 (O_1898,N_19963,N_19546);
nand UO_1899 (O_1899,N_19906,N_19854);
xor UO_1900 (O_1900,N_19984,N_19603);
and UO_1901 (O_1901,N_19783,N_19876);
nand UO_1902 (O_1902,N_19540,N_19637);
or UO_1903 (O_1903,N_19809,N_19581);
and UO_1904 (O_1904,N_19801,N_19629);
nor UO_1905 (O_1905,N_19987,N_19580);
xnor UO_1906 (O_1906,N_19588,N_19692);
nor UO_1907 (O_1907,N_19544,N_19983);
nor UO_1908 (O_1908,N_19605,N_19984);
nor UO_1909 (O_1909,N_19793,N_19900);
nor UO_1910 (O_1910,N_19659,N_19975);
or UO_1911 (O_1911,N_19910,N_19756);
nor UO_1912 (O_1912,N_19882,N_19850);
nor UO_1913 (O_1913,N_19558,N_19562);
and UO_1914 (O_1914,N_19697,N_19864);
and UO_1915 (O_1915,N_19588,N_19883);
or UO_1916 (O_1916,N_19708,N_19703);
and UO_1917 (O_1917,N_19677,N_19975);
xnor UO_1918 (O_1918,N_19529,N_19656);
nand UO_1919 (O_1919,N_19873,N_19943);
xor UO_1920 (O_1920,N_19899,N_19959);
nor UO_1921 (O_1921,N_19740,N_19715);
nor UO_1922 (O_1922,N_19754,N_19783);
xnor UO_1923 (O_1923,N_19786,N_19701);
nor UO_1924 (O_1924,N_19666,N_19822);
nand UO_1925 (O_1925,N_19773,N_19919);
or UO_1926 (O_1926,N_19579,N_19615);
xor UO_1927 (O_1927,N_19921,N_19861);
nor UO_1928 (O_1928,N_19964,N_19859);
nor UO_1929 (O_1929,N_19563,N_19823);
nand UO_1930 (O_1930,N_19603,N_19934);
nand UO_1931 (O_1931,N_19847,N_19902);
nand UO_1932 (O_1932,N_19899,N_19830);
and UO_1933 (O_1933,N_19845,N_19631);
and UO_1934 (O_1934,N_19774,N_19722);
and UO_1935 (O_1935,N_19793,N_19521);
xor UO_1936 (O_1936,N_19770,N_19933);
nor UO_1937 (O_1937,N_19816,N_19880);
nand UO_1938 (O_1938,N_19822,N_19804);
and UO_1939 (O_1939,N_19978,N_19831);
and UO_1940 (O_1940,N_19624,N_19701);
nor UO_1941 (O_1941,N_19711,N_19912);
nor UO_1942 (O_1942,N_19555,N_19509);
and UO_1943 (O_1943,N_19941,N_19505);
nor UO_1944 (O_1944,N_19847,N_19824);
nand UO_1945 (O_1945,N_19917,N_19717);
and UO_1946 (O_1946,N_19646,N_19621);
nand UO_1947 (O_1947,N_19946,N_19648);
and UO_1948 (O_1948,N_19741,N_19988);
and UO_1949 (O_1949,N_19618,N_19718);
nand UO_1950 (O_1950,N_19676,N_19817);
and UO_1951 (O_1951,N_19975,N_19629);
or UO_1952 (O_1952,N_19933,N_19882);
nand UO_1953 (O_1953,N_19978,N_19710);
nor UO_1954 (O_1954,N_19519,N_19639);
nor UO_1955 (O_1955,N_19721,N_19729);
nand UO_1956 (O_1956,N_19909,N_19756);
or UO_1957 (O_1957,N_19782,N_19892);
and UO_1958 (O_1958,N_19880,N_19790);
or UO_1959 (O_1959,N_19849,N_19605);
nand UO_1960 (O_1960,N_19631,N_19676);
xnor UO_1961 (O_1961,N_19806,N_19579);
and UO_1962 (O_1962,N_19571,N_19962);
nor UO_1963 (O_1963,N_19519,N_19796);
nor UO_1964 (O_1964,N_19699,N_19856);
and UO_1965 (O_1965,N_19768,N_19651);
or UO_1966 (O_1966,N_19533,N_19664);
nand UO_1967 (O_1967,N_19914,N_19663);
nand UO_1968 (O_1968,N_19949,N_19681);
nor UO_1969 (O_1969,N_19851,N_19592);
or UO_1970 (O_1970,N_19965,N_19580);
nand UO_1971 (O_1971,N_19570,N_19712);
or UO_1972 (O_1972,N_19637,N_19544);
or UO_1973 (O_1973,N_19831,N_19534);
or UO_1974 (O_1974,N_19894,N_19534);
nor UO_1975 (O_1975,N_19510,N_19635);
and UO_1976 (O_1976,N_19918,N_19631);
nor UO_1977 (O_1977,N_19932,N_19626);
nand UO_1978 (O_1978,N_19835,N_19666);
or UO_1979 (O_1979,N_19791,N_19856);
and UO_1980 (O_1980,N_19781,N_19892);
nand UO_1981 (O_1981,N_19798,N_19621);
and UO_1982 (O_1982,N_19955,N_19962);
nand UO_1983 (O_1983,N_19668,N_19761);
or UO_1984 (O_1984,N_19632,N_19649);
or UO_1985 (O_1985,N_19765,N_19990);
and UO_1986 (O_1986,N_19861,N_19819);
nand UO_1987 (O_1987,N_19640,N_19541);
nand UO_1988 (O_1988,N_19517,N_19818);
xnor UO_1989 (O_1989,N_19739,N_19621);
and UO_1990 (O_1990,N_19633,N_19983);
or UO_1991 (O_1991,N_19833,N_19506);
nor UO_1992 (O_1992,N_19937,N_19964);
nor UO_1993 (O_1993,N_19699,N_19683);
or UO_1994 (O_1994,N_19516,N_19579);
nor UO_1995 (O_1995,N_19836,N_19723);
and UO_1996 (O_1996,N_19959,N_19600);
nand UO_1997 (O_1997,N_19720,N_19678);
or UO_1998 (O_1998,N_19592,N_19808);
or UO_1999 (O_1999,N_19722,N_19790);
xor UO_2000 (O_2000,N_19520,N_19868);
nand UO_2001 (O_2001,N_19830,N_19716);
nand UO_2002 (O_2002,N_19727,N_19709);
xor UO_2003 (O_2003,N_19882,N_19902);
or UO_2004 (O_2004,N_19921,N_19780);
nand UO_2005 (O_2005,N_19912,N_19699);
or UO_2006 (O_2006,N_19638,N_19739);
or UO_2007 (O_2007,N_19730,N_19554);
or UO_2008 (O_2008,N_19895,N_19681);
nor UO_2009 (O_2009,N_19719,N_19516);
or UO_2010 (O_2010,N_19544,N_19984);
or UO_2011 (O_2011,N_19578,N_19706);
nand UO_2012 (O_2012,N_19599,N_19851);
or UO_2013 (O_2013,N_19980,N_19946);
nor UO_2014 (O_2014,N_19701,N_19825);
nand UO_2015 (O_2015,N_19536,N_19842);
nand UO_2016 (O_2016,N_19939,N_19729);
nand UO_2017 (O_2017,N_19546,N_19530);
and UO_2018 (O_2018,N_19661,N_19941);
xnor UO_2019 (O_2019,N_19755,N_19799);
and UO_2020 (O_2020,N_19800,N_19617);
nand UO_2021 (O_2021,N_19691,N_19929);
nand UO_2022 (O_2022,N_19977,N_19505);
or UO_2023 (O_2023,N_19865,N_19772);
nor UO_2024 (O_2024,N_19753,N_19794);
nor UO_2025 (O_2025,N_19765,N_19565);
nor UO_2026 (O_2026,N_19518,N_19824);
and UO_2027 (O_2027,N_19728,N_19667);
and UO_2028 (O_2028,N_19603,N_19883);
or UO_2029 (O_2029,N_19918,N_19635);
or UO_2030 (O_2030,N_19915,N_19745);
nand UO_2031 (O_2031,N_19886,N_19591);
xor UO_2032 (O_2032,N_19923,N_19579);
or UO_2033 (O_2033,N_19900,N_19629);
or UO_2034 (O_2034,N_19982,N_19740);
nand UO_2035 (O_2035,N_19635,N_19882);
xnor UO_2036 (O_2036,N_19792,N_19768);
and UO_2037 (O_2037,N_19770,N_19849);
and UO_2038 (O_2038,N_19694,N_19775);
and UO_2039 (O_2039,N_19695,N_19626);
nand UO_2040 (O_2040,N_19607,N_19874);
and UO_2041 (O_2041,N_19895,N_19635);
or UO_2042 (O_2042,N_19969,N_19603);
xor UO_2043 (O_2043,N_19514,N_19673);
and UO_2044 (O_2044,N_19585,N_19504);
nor UO_2045 (O_2045,N_19778,N_19577);
and UO_2046 (O_2046,N_19591,N_19522);
or UO_2047 (O_2047,N_19891,N_19745);
nor UO_2048 (O_2048,N_19764,N_19998);
or UO_2049 (O_2049,N_19576,N_19989);
or UO_2050 (O_2050,N_19566,N_19965);
and UO_2051 (O_2051,N_19669,N_19710);
nand UO_2052 (O_2052,N_19571,N_19558);
nor UO_2053 (O_2053,N_19962,N_19531);
and UO_2054 (O_2054,N_19784,N_19716);
or UO_2055 (O_2055,N_19697,N_19831);
or UO_2056 (O_2056,N_19546,N_19808);
and UO_2057 (O_2057,N_19770,N_19607);
and UO_2058 (O_2058,N_19837,N_19876);
nor UO_2059 (O_2059,N_19890,N_19807);
or UO_2060 (O_2060,N_19820,N_19753);
nand UO_2061 (O_2061,N_19698,N_19919);
nand UO_2062 (O_2062,N_19637,N_19659);
nor UO_2063 (O_2063,N_19939,N_19958);
nor UO_2064 (O_2064,N_19761,N_19815);
or UO_2065 (O_2065,N_19994,N_19632);
nand UO_2066 (O_2066,N_19865,N_19917);
and UO_2067 (O_2067,N_19681,N_19555);
and UO_2068 (O_2068,N_19568,N_19761);
nand UO_2069 (O_2069,N_19766,N_19589);
and UO_2070 (O_2070,N_19963,N_19895);
nand UO_2071 (O_2071,N_19665,N_19911);
nor UO_2072 (O_2072,N_19598,N_19891);
or UO_2073 (O_2073,N_19987,N_19846);
xor UO_2074 (O_2074,N_19674,N_19894);
nor UO_2075 (O_2075,N_19544,N_19740);
or UO_2076 (O_2076,N_19982,N_19999);
and UO_2077 (O_2077,N_19810,N_19990);
or UO_2078 (O_2078,N_19982,N_19862);
or UO_2079 (O_2079,N_19817,N_19895);
xnor UO_2080 (O_2080,N_19536,N_19886);
nand UO_2081 (O_2081,N_19623,N_19855);
and UO_2082 (O_2082,N_19965,N_19846);
nor UO_2083 (O_2083,N_19956,N_19821);
nand UO_2084 (O_2084,N_19877,N_19690);
nand UO_2085 (O_2085,N_19862,N_19941);
and UO_2086 (O_2086,N_19821,N_19783);
or UO_2087 (O_2087,N_19520,N_19943);
or UO_2088 (O_2088,N_19947,N_19652);
nor UO_2089 (O_2089,N_19533,N_19520);
nand UO_2090 (O_2090,N_19750,N_19832);
or UO_2091 (O_2091,N_19920,N_19852);
nand UO_2092 (O_2092,N_19570,N_19906);
xor UO_2093 (O_2093,N_19770,N_19852);
or UO_2094 (O_2094,N_19861,N_19815);
or UO_2095 (O_2095,N_19926,N_19608);
or UO_2096 (O_2096,N_19883,N_19607);
xnor UO_2097 (O_2097,N_19722,N_19700);
and UO_2098 (O_2098,N_19784,N_19806);
xor UO_2099 (O_2099,N_19769,N_19578);
and UO_2100 (O_2100,N_19996,N_19554);
and UO_2101 (O_2101,N_19659,N_19703);
nand UO_2102 (O_2102,N_19740,N_19793);
nor UO_2103 (O_2103,N_19582,N_19945);
or UO_2104 (O_2104,N_19987,N_19501);
nand UO_2105 (O_2105,N_19591,N_19957);
xnor UO_2106 (O_2106,N_19731,N_19946);
and UO_2107 (O_2107,N_19910,N_19845);
nand UO_2108 (O_2108,N_19861,N_19756);
or UO_2109 (O_2109,N_19788,N_19605);
or UO_2110 (O_2110,N_19791,N_19824);
or UO_2111 (O_2111,N_19586,N_19776);
and UO_2112 (O_2112,N_19692,N_19589);
nor UO_2113 (O_2113,N_19937,N_19609);
nand UO_2114 (O_2114,N_19789,N_19773);
nand UO_2115 (O_2115,N_19623,N_19512);
nand UO_2116 (O_2116,N_19894,N_19956);
nand UO_2117 (O_2117,N_19896,N_19769);
and UO_2118 (O_2118,N_19502,N_19640);
nand UO_2119 (O_2119,N_19654,N_19612);
and UO_2120 (O_2120,N_19674,N_19878);
nand UO_2121 (O_2121,N_19689,N_19543);
nand UO_2122 (O_2122,N_19661,N_19846);
nand UO_2123 (O_2123,N_19509,N_19752);
and UO_2124 (O_2124,N_19879,N_19550);
xnor UO_2125 (O_2125,N_19569,N_19599);
nand UO_2126 (O_2126,N_19721,N_19530);
nor UO_2127 (O_2127,N_19652,N_19979);
nand UO_2128 (O_2128,N_19714,N_19808);
and UO_2129 (O_2129,N_19965,N_19684);
or UO_2130 (O_2130,N_19722,N_19734);
nor UO_2131 (O_2131,N_19527,N_19670);
and UO_2132 (O_2132,N_19707,N_19727);
xnor UO_2133 (O_2133,N_19994,N_19522);
or UO_2134 (O_2134,N_19615,N_19766);
nand UO_2135 (O_2135,N_19872,N_19807);
or UO_2136 (O_2136,N_19740,N_19532);
nor UO_2137 (O_2137,N_19596,N_19884);
nand UO_2138 (O_2138,N_19640,N_19953);
or UO_2139 (O_2139,N_19937,N_19886);
or UO_2140 (O_2140,N_19962,N_19844);
and UO_2141 (O_2141,N_19987,N_19513);
and UO_2142 (O_2142,N_19658,N_19805);
and UO_2143 (O_2143,N_19993,N_19963);
nand UO_2144 (O_2144,N_19882,N_19555);
nand UO_2145 (O_2145,N_19605,N_19862);
nand UO_2146 (O_2146,N_19925,N_19858);
nand UO_2147 (O_2147,N_19620,N_19949);
and UO_2148 (O_2148,N_19505,N_19909);
xor UO_2149 (O_2149,N_19561,N_19552);
nand UO_2150 (O_2150,N_19855,N_19510);
nand UO_2151 (O_2151,N_19668,N_19714);
nor UO_2152 (O_2152,N_19960,N_19699);
xor UO_2153 (O_2153,N_19509,N_19558);
or UO_2154 (O_2154,N_19985,N_19816);
nor UO_2155 (O_2155,N_19971,N_19863);
nand UO_2156 (O_2156,N_19929,N_19861);
xnor UO_2157 (O_2157,N_19840,N_19628);
or UO_2158 (O_2158,N_19893,N_19817);
nor UO_2159 (O_2159,N_19968,N_19825);
or UO_2160 (O_2160,N_19589,N_19790);
nand UO_2161 (O_2161,N_19537,N_19656);
nor UO_2162 (O_2162,N_19686,N_19963);
and UO_2163 (O_2163,N_19827,N_19729);
or UO_2164 (O_2164,N_19845,N_19737);
and UO_2165 (O_2165,N_19806,N_19946);
or UO_2166 (O_2166,N_19507,N_19901);
nor UO_2167 (O_2167,N_19634,N_19938);
nor UO_2168 (O_2168,N_19599,N_19824);
xnor UO_2169 (O_2169,N_19862,N_19590);
nand UO_2170 (O_2170,N_19693,N_19859);
nor UO_2171 (O_2171,N_19675,N_19944);
and UO_2172 (O_2172,N_19891,N_19612);
nor UO_2173 (O_2173,N_19634,N_19711);
nor UO_2174 (O_2174,N_19937,N_19631);
nor UO_2175 (O_2175,N_19505,N_19569);
nand UO_2176 (O_2176,N_19558,N_19743);
nor UO_2177 (O_2177,N_19647,N_19853);
or UO_2178 (O_2178,N_19584,N_19528);
nor UO_2179 (O_2179,N_19991,N_19911);
nand UO_2180 (O_2180,N_19942,N_19894);
or UO_2181 (O_2181,N_19693,N_19876);
or UO_2182 (O_2182,N_19596,N_19553);
nor UO_2183 (O_2183,N_19850,N_19957);
and UO_2184 (O_2184,N_19676,N_19643);
nor UO_2185 (O_2185,N_19583,N_19674);
nor UO_2186 (O_2186,N_19500,N_19913);
and UO_2187 (O_2187,N_19549,N_19791);
or UO_2188 (O_2188,N_19536,N_19732);
and UO_2189 (O_2189,N_19973,N_19998);
or UO_2190 (O_2190,N_19936,N_19765);
nor UO_2191 (O_2191,N_19860,N_19649);
nand UO_2192 (O_2192,N_19664,N_19849);
or UO_2193 (O_2193,N_19572,N_19653);
nor UO_2194 (O_2194,N_19594,N_19776);
or UO_2195 (O_2195,N_19819,N_19746);
nor UO_2196 (O_2196,N_19968,N_19715);
or UO_2197 (O_2197,N_19798,N_19823);
nor UO_2198 (O_2198,N_19534,N_19505);
nand UO_2199 (O_2199,N_19680,N_19874);
or UO_2200 (O_2200,N_19746,N_19526);
or UO_2201 (O_2201,N_19525,N_19572);
nor UO_2202 (O_2202,N_19904,N_19626);
and UO_2203 (O_2203,N_19684,N_19646);
nand UO_2204 (O_2204,N_19526,N_19722);
nand UO_2205 (O_2205,N_19961,N_19596);
nor UO_2206 (O_2206,N_19891,N_19956);
nand UO_2207 (O_2207,N_19561,N_19835);
and UO_2208 (O_2208,N_19925,N_19949);
nor UO_2209 (O_2209,N_19955,N_19870);
or UO_2210 (O_2210,N_19917,N_19849);
nand UO_2211 (O_2211,N_19932,N_19554);
nor UO_2212 (O_2212,N_19555,N_19819);
nor UO_2213 (O_2213,N_19550,N_19992);
or UO_2214 (O_2214,N_19786,N_19830);
nand UO_2215 (O_2215,N_19613,N_19666);
nand UO_2216 (O_2216,N_19598,N_19938);
nor UO_2217 (O_2217,N_19709,N_19918);
nor UO_2218 (O_2218,N_19720,N_19907);
or UO_2219 (O_2219,N_19564,N_19826);
nand UO_2220 (O_2220,N_19537,N_19759);
and UO_2221 (O_2221,N_19611,N_19947);
nand UO_2222 (O_2222,N_19988,N_19582);
or UO_2223 (O_2223,N_19677,N_19641);
and UO_2224 (O_2224,N_19678,N_19734);
xor UO_2225 (O_2225,N_19959,N_19816);
xnor UO_2226 (O_2226,N_19933,N_19983);
nor UO_2227 (O_2227,N_19928,N_19788);
nor UO_2228 (O_2228,N_19639,N_19854);
or UO_2229 (O_2229,N_19680,N_19759);
nor UO_2230 (O_2230,N_19806,N_19676);
nand UO_2231 (O_2231,N_19894,N_19940);
or UO_2232 (O_2232,N_19583,N_19785);
and UO_2233 (O_2233,N_19738,N_19705);
nand UO_2234 (O_2234,N_19782,N_19568);
nand UO_2235 (O_2235,N_19615,N_19730);
nand UO_2236 (O_2236,N_19542,N_19696);
nor UO_2237 (O_2237,N_19979,N_19774);
or UO_2238 (O_2238,N_19522,N_19835);
nand UO_2239 (O_2239,N_19577,N_19645);
nor UO_2240 (O_2240,N_19584,N_19949);
xnor UO_2241 (O_2241,N_19672,N_19759);
or UO_2242 (O_2242,N_19735,N_19789);
nand UO_2243 (O_2243,N_19660,N_19671);
nor UO_2244 (O_2244,N_19746,N_19661);
nand UO_2245 (O_2245,N_19719,N_19806);
nor UO_2246 (O_2246,N_19722,N_19777);
and UO_2247 (O_2247,N_19626,N_19782);
nor UO_2248 (O_2248,N_19637,N_19772);
nand UO_2249 (O_2249,N_19875,N_19998);
and UO_2250 (O_2250,N_19513,N_19860);
and UO_2251 (O_2251,N_19995,N_19586);
nor UO_2252 (O_2252,N_19942,N_19949);
and UO_2253 (O_2253,N_19931,N_19793);
nand UO_2254 (O_2254,N_19950,N_19593);
nor UO_2255 (O_2255,N_19831,N_19511);
nor UO_2256 (O_2256,N_19511,N_19852);
nand UO_2257 (O_2257,N_19936,N_19793);
and UO_2258 (O_2258,N_19782,N_19615);
or UO_2259 (O_2259,N_19981,N_19599);
nand UO_2260 (O_2260,N_19812,N_19709);
and UO_2261 (O_2261,N_19865,N_19659);
xnor UO_2262 (O_2262,N_19925,N_19673);
or UO_2263 (O_2263,N_19658,N_19677);
and UO_2264 (O_2264,N_19770,N_19556);
xnor UO_2265 (O_2265,N_19883,N_19759);
nand UO_2266 (O_2266,N_19526,N_19678);
nand UO_2267 (O_2267,N_19865,N_19553);
nor UO_2268 (O_2268,N_19815,N_19759);
and UO_2269 (O_2269,N_19559,N_19545);
xor UO_2270 (O_2270,N_19583,N_19698);
nor UO_2271 (O_2271,N_19668,N_19958);
nor UO_2272 (O_2272,N_19514,N_19544);
nor UO_2273 (O_2273,N_19627,N_19793);
or UO_2274 (O_2274,N_19672,N_19729);
or UO_2275 (O_2275,N_19695,N_19988);
nand UO_2276 (O_2276,N_19642,N_19831);
and UO_2277 (O_2277,N_19900,N_19617);
and UO_2278 (O_2278,N_19884,N_19613);
nor UO_2279 (O_2279,N_19774,N_19839);
nor UO_2280 (O_2280,N_19756,N_19700);
nor UO_2281 (O_2281,N_19872,N_19952);
or UO_2282 (O_2282,N_19720,N_19781);
nor UO_2283 (O_2283,N_19521,N_19803);
and UO_2284 (O_2284,N_19842,N_19711);
xnor UO_2285 (O_2285,N_19801,N_19597);
or UO_2286 (O_2286,N_19660,N_19812);
and UO_2287 (O_2287,N_19801,N_19924);
or UO_2288 (O_2288,N_19618,N_19798);
nand UO_2289 (O_2289,N_19716,N_19868);
and UO_2290 (O_2290,N_19726,N_19855);
and UO_2291 (O_2291,N_19940,N_19891);
nor UO_2292 (O_2292,N_19714,N_19733);
nand UO_2293 (O_2293,N_19597,N_19877);
or UO_2294 (O_2294,N_19639,N_19850);
nor UO_2295 (O_2295,N_19857,N_19954);
or UO_2296 (O_2296,N_19663,N_19698);
xnor UO_2297 (O_2297,N_19943,N_19713);
or UO_2298 (O_2298,N_19814,N_19964);
nor UO_2299 (O_2299,N_19907,N_19744);
or UO_2300 (O_2300,N_19604,N_19537);
and UO_2301 (O_2301,N_19547,N_19657);
and UO_2302 (O_2302,N_19956,N_19515);
and UO_2303 (O_2303,N_19854,N_19745);
and UO_2304 (O_2304,N_19834,N_19716);
or UO_2305 (O_2305,N_19803,N_19544);
or UO_2306 (O_2306,N_19967,N_19671);
nor UO_2307 (O_2307,N_19669,N_19832);
xnor UO_2308 (O_2308,N_19706,N_19934);
xnor UO_2309 (O_2309,N_19558,N_19829);
nand UO_2310 (O_2310,N_19942,N_19755);
and UO_2311 (O_2311,N_19817,N_19849);
nor UO_2312 (O_2312,N_19896,N_19731);
and UO_2313 (O_2313,N_19901,N_19761);
and UO_2314 (O_2314,N_19984,N_19958);
or UO_2315 (O_2315,N_19710,N_19619);
nor UO_2316 (O_2316,N_19778,N_19797);
and UO_2317 (O_2317,N_19625,N_19569);
and UO_2318 (O_2318,N_19820,N_19734);
or UO_2319 (O_2319,N_19686,N_19533);
nor UO_2320 (O_2320,N_19795,N_19976);
nand UO_2321 (O_2321,N_19866,N_19753);
xor UO_2322 (O_2322,N_19531,N_19971);
nor UO_2323 (O_2323,N_19748,N_19951);
nand UO_2324 (O_2324,N_19843,N_19723);
nor UO_2325 (O_2325,N_19955,N_19665);
or UO_2326 (O_2326,N_19957,N_19523);
nand UO_2327 (O_2327,N_19832,N_19829);
xor UO_2328 (O_2328,N_19893,N_19959);
nand UO_2329 (O_2329,N_19823,N_19894);
nand UO_2330 (O_2330,N_19955,N_19963);
and UO_2331 (O_2331,N_19972,N_19555);
and UO_2332 (O_2332,N_19660,N_19603);
nand UO_2333 (O_2333,N_19840,N_19654);
nand UO_2334 (O_2334,N_19898,N_19654);
nand UO_2335 (O_2335,N_19654,N_19702);
xnor UO_2336 (O_2336,N_19506,N_19889);
nor UO_2337 (O_2337,N_19995,N_19804);
nor UO_2338 (O_2338,N_19595,N_19840);
nor UO_2339 (O_2339,N_19960,N_19942);
nor UO_2340 (O_2340,N_19682,N_19941);
nor UO_2341 (O_2341,N_19521,N_19758);
nor UO_2342 (O_2342,N_19837,N_19546);
and UO_2343 (O_2343,N_19730,N_19830);
and UO_2344 (O_2344,N_19944,N_19538);
nand UO_2345 (O_2345,N_19633,N_19623);
or UO_2346 (O_2346,N_19555,N_19797);
and UO_2347 (O_2347,N_19893,N_19925);
nand UO_2348 (O_2348,N_19835,N_19837);
nor UO_2349 (O_2349,N_19716,N_19974);
and UO_2350 (O_2350,N_19695,N_19661);
and UO_2351 (O_2351,N_19642,N_19762);
nor UO_2352 (O_2352,N_19537,N_19549);
and UO_2353 (O_2353,N_19938,N_19920);
nor UO_2354 (O_2354,N_19712,N_19848);
and UO_2355 (O_2355,N_19743,N_19752);
and UO_2356 (O_2356,N_19569,N_19821);
or UO_2357 (O_2357,N_19933,N_19643);
and UO_2358 (O_2358,N_19722,N_19511);
or UO_2359 (O_2359,N_19873,N_19597);
or UO_2360 (O_2360,N_19905,N_19865);
nor UO_2361 (O_2361,N_19772,N_19828);
or UO_2362 (O_2362,N_19806,N_19942);
xnor UO_2363 (O_2363,N_19699,N_19739);
nand UO_2364 (O_2364,N_19728,N_19990);
nor UO_2365 (O_2365,N_19836,N_19930);
and UO_2366 (O_2366,N_19614,N_19662);
nor UO_2367 (O_2367,N_19724,N_19527);
nand UO_2368 (O_2368,N_19778,N_19676);
nand UO_2369 (O_2369,N_19857,N_19886);
or UO_2370 (O_2370,N_19902,N_19546);
nand UO_2371 (O_2371,N_19906,N_19800);
xnor UO_2372 (O_2372,N_19753,N_19970);
nand UO_2373 (O_2373,N_19817,N_19773);
nor UO_2374 (O_2374,N_19732,N_19659);
xnor UO_2375 (O_2375,N_19798,N_19818);
nor UO_2376 (O_2376,N_19730,N_19624);
nor UO_2377 (O_2377,N_19942,N_19713);
nor UO_2378 (O_2378,N_19744,N_19598);
nand UO_2379 (O_2379,N_19836,N_19749);
nand UO_2380 (O_2380,N_19777,N_19779);
nor UO_2381 (O_2381,N_19655,N_19877);
and UO_2382 (O_2382,N_19834,N_19785);
or UO_2383 (O_2383,N_19981,N_19709);
nor UO_2384 (O_2384,N_19556,N_19834);
nor UO_2385 (O_2385,N_19908,N_19881);
or UO_2386 (O_2386,N_19502,N_19779);
and UO_2387 (O_2387,N_19647,N_19867);
nor UO_2388 (O_2388,N_19783,N_19774);
and UO_2389 (O_2389,N_19680,N_19935);
or UO_2390 (O_2390,N_19982,N_19605);
nand UO_2391 (O_2391,N_19920,N_19897);
nor UO_2392 (O_2392,N_19948,N_19840);
nand UO_2393 (O_2393,N_19881,N_19546);
nor UO_2394 (O_2394,N_19561,N_19952);
and UO_2395 (O_2395,N_19596,N_19515);
or UO_2396 (O_2396,N_19940,N_19608);
nor UO_2397 (O_2397,N_19567,N_19559);
xor UO_2398 (O_2398,N_19660,N_19623);
and UO_2399 (O_2399,N_19822,N_19659);
nor UO_2400 (O_2400,N_19932,N_19760);
or UO_2401 (O_2401,N_19555,N_19846);
and UO_2402 (O_2402,N_19889,N_19698);
xnor UO_2403 (O_2403,N_19858,N_19666);
xor UO_2404 (O_2404,N_19578,N_19502);
or UO_2405 (O_2405,N_19726,N_19623);
nor UO_2406 (O_2406,N_19537,N_19532);
xnor UO_2407 (O_2407,N_19776,N_19889);
and UO_2408 (O_2408,N_19983,N_19622);
nand UO_2409 (O_2409,N_19711,N_19626);
and UO_2410 (O_2410,N_19676,N_19839);
or UO_2411 (O_2411,N_19941,N_19526);
or UO_2412 (O_2412,N_19613,N_19977);
nor UO_2413 (O_2413,N_19647,N_19653);
and UO_2414 (O_2414,N_19722,N_19975);
xor UO_2415 (O_2415,N_19929,N_19966);
xnor UO_2416 (O_2416,N_19685,N_19868);
and UO_2417 (O_2417,N_19594,N_19783);
nand UO_2418 (O_2418,N_19713,N_19852);
or UO_2419 (O_2419,N_19705,N_19920);
or UO_2420 (O_2420,N_19642,N_19956);
nand UO_2421 (O_2421,N_19869,N_19525);
and UO_2422 (O_2422,N_19722,N_19665);
or UO_2423 (O_2423,N_19572,N_19626);
and UO_2424 (O_2424,N_19528,N_19883);
or UO_2425 (O_2425,N_19673,N_19619);
nand UO_2426 (O_2426,N_19670,N_19905);
nor UO_2427 (O_2427,N_19899,N_19755);
nor UO_2428 (O_2428,N_19655,N_19734);
nor UO_2429 (O_2429,N_19760,N_19656);
nor UO_2430 (O_2430,N_19858,N_19608);
xor UO_2431 (O_2431,N_19771,N_19605);
or UO_2432 (O_2432,N_19970,N_19796);
or UO_2433 (O_2433,N_19798,N_19957);
nand UO_2434 (O_2434,N_19936,N_19913);
nor UO_2435 (O_2435,N_19533,N_19617);
nor UO_2436 (O_2436,N_19699,N_19805);
nor UO_2437 (O_2437,N_19545,N_19557);
xnor UO_2438 (O_2438,N_19910,N_19912);
nor UO_2439 (O_2439,N_19774,N_19841);
nor UO_2440 (O_2440,N_19785,N_19735);
xor UO_2441 (O_2441,N_19971,N_19815);
nor UO_2442 (O_2442,N_19717,N_19943);
nand UO_2443 (O_2443,N_19909,N_19917);
and UO_2444 (O_2444,N_19922,N_19678);
or UO_2445 (O_2445,N_19861,N_19505);
nand UO_2446 (O_2446,N_19686,N_19544);
nand UO_2447 (O_2447,N_19963,N_19990);
or UO_2448 (O_2448,N_19557,N_19885);
or UO_2449 (O_2449,N_19652,N_19941);
nand UO_2450 (O_2450,N_19529,N_19640);
or UO_2451 (O_2451,N_19753,N_19676);
xor UO_2452 (O_2452,N_19548,N_19541);
nand UO_2453 (O_2453,N_19682,N_19862);
nor UO_2454 (O_2454,N_19868,N_19791);
or UO_2455 (O_2455,N_19543,N_19729);
nand UO_2456 (O_2456,N_19946,N_19532);
or UO_2457 (O_2457,N_19742,N_19788);
nor UO_2458 (O_2458,N_19885,N_19604);
and UO_2459 (O_2459,N_19870,N_19918);
xnor UO_2460 (O_2460,N_19911,N_19531);
or UO_2461 (O_2461,N_19754,N_19643);
or UO_2462 (O_2462,N_19656,N_19786);
and UO_2463 (O_2463,N_19528,N_19539);
or UO_2464 (O_2464,N_19526,N_19895);
nand UO_2465 (O_2465,N_19685,N_19586);
nor UO_2466 (O_2466,N_19968,N_19504);
nor UO_2467 (O_2467,N_19573,N_19768);
or UO_2468 (O_2468,N_19918,N_19981);
xor UO_2469 (O_2469,N_19574,N_19635);
nand UO_2470 (O_2470,N_19993,N_19656);
or UO_2471 (O_2471,N_19730,N_19744);
nor UO_2472 (O_2472,N_19918,N_19729);
or UO_2473 (O_2473,N_19752,N_19876);
xnor UO_2474 (O_2474,N_19835,N_19924);
or UO_2475 (O_2475,N_19567,N_19803);
or UO_2476 (O_2476,N_19565,N_19777);
nand UO_2477 (O_2477,N_19592,N_19570);
nand UO_2478 (O_2478,N_19612,N_19613);
nor UO_2479 (O_2479,N_19729,N_19724);
and UO_2480 (O_2480,N_19638,N_19581);
xor UO_2481 (O_2481,N_19531,N_19777);
nor UO_2482 (O_2482,N_19513,N_19804);
nand UO_2483 (O_2483,N_19586,N_19897);
nand UO_2484 (O_2484,N_19980,N_19796);
and UO_2485 (O_2485,N_19820,N_19927);
and UO_2486 (O_2486,N_19505,N_19613);
or UO_2487 (O_2487,N_19585,N_19767);
nand UO_2488 (O_2488,N_19733,N_19749);
or UO_2489 (O_2489,N_19725,N_19638);
nand UO_2490 (O_2490,N_19768,N_19716);
xnor UO_2491 (O_2491,N_19800,N_19690);
and UO_2492 (O_2492,N_19777,N_19532);
nand UO_2493 (O_2493,N_19752,N_19760);
and UO_2494 (O_2494,N_19679,N_19960);
nand UO_2495 (O_2495,N_19639,N_19852);
and UO_2496 (O_2496,N_19773,N_19960);
xnor UO_2497 (O_2497,N_19704,N_19576);
nor UO_2498 (O_2498,N_19799,N_19645);
and UO_2499 (O_2499,N_19556,N_19583);
endmodule