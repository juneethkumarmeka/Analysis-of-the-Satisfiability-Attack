module basic_1000_10000_1500_10_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_701,In_642);
nor U1 (N_1,In_706,In_837);
xnor U2 (N_2,In_789,In_371);
nand U3 (N_3,In_657,In_806);
xor U4 (N_4,In_704,In_717);
nand U5 (N_5,In_303,In_690);
nor U6 (N_6,In_253,In_297);
and U7 (N_7,In_815,In_425);
nor U8 (N_8,In_902,In_75);
nand U9 (N_9,In_278,In_0);
nand U10 (N_10,In_80,In_218);
and U11 (N_11,In_46,In_621);
and U12 (N_12,In_664,In_613);
nor U13 (N_13,In_810,In_333);
xnor U14 (N_14,In_381,In_460);
nand U15 (N_15,In_391,In_928);
nand U16 (N_16,In_796,In_399);
nand U17 (N_17,In_968,In_211);
nor U18 (N_18,In_615,In_42);
xnor U19 (N_19,In_554,In_597);
xnor U20 (N_20,In_485,In_186);
or U21 (N_21,In_936,In_343);
or U22 (N_22,In_572,In_667);
or U23 (N_23,In_834,In_188);
and U24 (N_24,In_49,In_752);
xnor U25 (N_25,In_405,In_937);
and U26 (N_26,In_67,In_130);
and U27 (N_27,In_892,In_941);
or U28 (N_28,In_248,In_808);
xor U29 (N_29,In_935,In_675);
or U30 (N_30,In_279,In_52);
and U31 (N_31,In_756,In_584);
nand U32 (N_32,In_511,In_13);
and U33 (N_33,In_659,In_955);
xor U34 (N_34,In_417,In_816);
nor U35 (N_35,In_821,In_22);
and U36 (N_36,In_848,In_838);
xnor U37 (N_37,In_727,In_880);
and U38 (N_38,In_385,In_576);
nor U39 (N_39,In_787,In_889);
nand U40 (N_40,In_54,In_366);
and U41 (N_41,In_660,In_392);
xor U42 (N_42,In_703,In_341);
or U43 (N_43,In_369,In_940);
nor U44 (N_44,In_166,In_770);
nor U45 (N_45,In_488,In_35);
nor U46 (N_46,In_709,In_643);
nor U47 (N_47,In_846,In_550);
nor U48 (N_48,In_823,In_145);
or U49 (N_49,In_463,In_11);
nor U50 (N_50,In_670,In_931);
and U51 (N_51,In_612,In_869);
nand U52 (N_52,In_68,In_975);
nor U53 (N_53,In_626,In_595);
xnor U54 (N_54,In_534,In_541);
or U55 (N_55,In_714,In_114);
xnor U56 (N_56,In_991,In_436);
or U57 (N_57,In_88,In_396);
or U58 (N_58,In_339,In_547);
xor U59 (N_59,In_990,In_627);
nor U60 (N_60,In_348,In_895);
and U61 (N_61,In_546,In_687);
or U62 (N_62,In_241,In_216);
nand U63 (N_63,In_799,In_750);
or U64 (N_64,In_645,In_607);
and U65 (N_65,In_143,In_331);
and U66 (N_66,In_144,In_450);
nor U67 (N_67,In_454,In_977);
or U68 (N_68,In_411,In_212);
nand U69 (N_69,In_938,In_61);
nor U70 (N_70,In_428,In_592);
or U71 (N_71,In_281,In_220);
nor U72 (N_72,In_581,In_555);
or U73 (N_73,In_978,In_908);
nand U74 (N_74,In_679,In_693);
and U75 (N_75,In_844,In_833);
nor U76 (N_76,In_89,In_668);
nor U77 (N_77,In_8,In_324);
nand U78 (N_78,In_422,In_329);
xnor U79 (N_79,In_539,In_876);
xor U80 (N_80,In_110,In_301);
or U81 (N_81,In_338,In_50);
or U82 (N_82,In_85,In_138);
nand U83 (N_83,In_256,In_711);
xnor U84 (N_84,In_367,In_856);
nor U85 (N_85,In_774,In_912);
xnor U86 (N_86,In_408,In_420);
xnor U87 (N_87,In_24,In_947);
xnor U88 (N_88,In_618,In_20);
xor U89 (N_89,In_307,In_589);
nor U90 (N_90,In_872,In_743);
xnor U91 (N_91,In_115,In_309);
nor U92 (N_92,In_536,In_429);
xor U93 (N_93,In_854,In_374);
nand U94 (N_94,In_364,In_865);
and U95 (N_95,In_721,In_171);
nor U96 (N_96,In_793,In_363);
xor U97 (N_97,In_795,In_406);
or U98 (N_98,In_82,In_780);
nor U99 (N_99,In_2,In_655);
and U100 (N_100,In_305,In_802);
or U101 (N_101,In_580,In_244);
or U102 (N_102,In_404,In_55);
and U103 (N_103,In_773,In_861);
nand U104 (N_104,In_632,In_337);
and U105 (N_105,In_499,In_261);
xnor U106 (N_106,In_21,In_432);
nand U107 (N_107,In_317,In_263);
nand U108 (N_108,In_150,In_974);
nand U109 (N_109,In_735,In_830);
nor U110 (N_110,In_782,In_163);
xor U111 (N_111,In_335,In_493);
xor U112 (N_112,In_72,In_243);
nand U113 (N_113,In_433,In_585);
nor U114 (N_114,In_828,In_684);
or U115 (N_115,In_918,In_972);
nand U116 (N_116,In_416,In_287);
or U117 (N_117,In_268,In_291);
xor U118 (N_118,In_386,In_131);
xor U119 (N_119,In_40,In_683);
nand U120 (N_120,In_376,In_122);
xnor U121 (N_121,In_781,In_598);
or U122 (N_122,In_982,In_790);
or U123 (N_123,In_739,In_707);
xor U124 (N_124,In_622,In_112);
or U125 (N_125,In_206,In_356);
xor U126 (N_126,In_151,In_71);
or U127 (N_127,In_956,In_702);
nor U128 (N_128,In_853,In_258);
and U129 (N_129,In_923,In_473);
nand U130 (N_130,In_898,In_847);
nor U131 (N_131,In_304,In_201);
nor U132 (N_132,In_540,In_987);
and U133 (N_133,In_323,In_45);
and U134 (N_134,In_820,In_299);
and U135 (N_135,In_93,In_108);
or U136 (N_136,In_639,In_440);
and U137 (N_137,In_885,In_360);
or U138 (N_138,In_564,In_202);
or U139 (N_139,In_601,In_219);
nor U140 (N_140,In_934,In_894);
nor U141 (N_141,In_867,In_456);
or U142 (N_142,In_855,In_183);
xnor U143 (N_143,In_388,In_357);
nor U144 (N_144,In_728,In_916);
and U145 (N_145,In_373,In_538);
nand U146 (N_146,In_311,In_284);
xor U147 (N_147,In_494,In_650);
nor U148 (N_148,In_868,In_298);
and U149 (N_149,In_749,In_768);
xnor U150 (N_150,In_905,In_181);
nand U151 (N_151,In_497,In_678);
and U152 (N_152,In_101,In_48);
xor U153 (N_153,In_226,In_33);
nor U154 (N_154,In_361,In_575);
nand U155 (N_155,In_187,In_302);
or U156 (N_156,In_467,In_992);
nor U157 (N_157,In_553,In_345);
xnor U158 (N_158,In_322,In_648);
and U159 (N_159,In_142,In_843);
nand U160 (N_160,In_772,In_958);
xor U161 (N_161,In_930,In_97);
nor U162 (N_162,In_259,In_353);
and U163 (N_163,In_686,In_746);
and U164 (N_164,In_507,In_198);
and U165 (N_165,In_634,In_496);
or U166 (N_166,In_63,In_368);
nand U167 (N_167,In_922,In_141);
xor U168 (N_168,In_321,In_246);
or U169 (N_169,In_451,In_633);
nand U170 (N_170,In_383,In_3);
xor U171 (N_171,In_194,In_953);
nor U172 (N_172,In_280,In_441);
nor U173 (N_173,In_6,In_822);
xnor U174 (N_174,In_290,In_751);
or U175 (N_175,In_168,In_900);
xnor U176 (N_176,In_736,In_119);
xnor U177 (N_177,In_545,In_177);
xnor U178 (N_178,In_740,In_677);
nand U179 (N_179,In_235,In_443);
xnor U180 (N_180,In_242,In_608);
xnor U181 (N_181,In_980,In_897);
or U182 (N_182,In_225,In_695);
xnor U183 (N_183,In_124,In_53);
or U184 (N_184,In_999,In_901);
nand U185 (N_185,In_9,In_951);
xor U186 (N_186,In_51,In_334);
or U187 (N_187,In_34,In_245);
and U188 (N_188,In_336,In_609);
nand U189 (N_189,In_884,In_556);
nand U190 (N_190,In_676,In_891);
nand U191 (N_191,In_566,In_669);
and U192 (N_192,In_824,In_407);
and U193 (N_193,In_641,In_73);
nor U194 (N_194,In_102,In_207);
xor U195 (N_195,In_74,In_427);
or U196 (N_196,In_267,In_380);
nor U197 (N_197,In_689,In_691);
xnor U198 (N_198,In_66,In_529);
or U199 (N_199,In_478,In_758);
nor U200 (N_200,In_926,In_996);
nand U201 (N_201,In_924,In_510);
nor U202 (N_202,In_41,In_172);
or U203 (N_203,In_535,In_994);
nand U204 (N_204,In_221,In_447);
and U205 (N_205,In_91,In_710);
xor U206 (N_206,In_92,In_995);
and U207 (N_207,In_520,In_104);
and U208 (N_208,In_197,In_176);
xnor U209 (N_209,In_43,In_31);
nor U210 (N_210,In_182,In_811);
nor U211 (N_211,In_969,In_631);
and U212 (N_212,In_763,In_504);
or U213 (N_213,In_505,In_685);
nand U214 (N_214,In_984,In_573);
nor U215 (N_215,In_475,In_306);
or U216 (N_216,In_674,In_814);
nor U217 (N_217,In_439,In_526);
xor U218 (N_218,In_588,In_503);
or U219 (N_219,In_552,In_946);
or U220 (N_220,In_149,In_522);
and U221 (N_221,In_81,In_954);
nor U222 (N_222,In_285,In_841);
xor U223 (N_223,In_582,In_77);
or U224 (N_224,In_379,In_753);
nor U225 (N_225,In_318,In_402);
nor U226 (N_226,In_136,In_647);
or U227 (N_227,In_459,In_827);
nor U228 (N_228,In_418,In_875);
nand U229 (N_229,In_779,In_989);
nor U230 (N_230,In_903,In_312);
and U231 (N_231,In_965,In_195);
or U232 (N_232,In_542,In_730);
nor U233 (N_233,In_44,In_314);
xor U234 (N_234,In_160,In_874);
or U235 (N_235,In_568,In_680);
xnor U236 (N_236,In_277,In_389);
xor U237 (N_237,In_185,In_755);
and U238 (N_238,In_489,In_530);
or U239 (N_239,In_169,In_126);
and U240 (N_240,In_184,In_286);
or U241 (N_241,In_313,In_58);
nand U242 (N_242,In_656,In_771);
or U243 (N_243,In_466,In_269);
and U244 (N_244,In_320,In_435);
or U245 (N_245,In_403,In_121);
and U246 (N_246,In_860,In_914);
or U247 (N_247,In_156,In_105);
nor U248 (N_248,In_325,In_118);
nor U249 (N_249,In_733,In_512);
nor U250 (N_250,In_797,In_579);
nand U251 (N_251,In_986,In_490);
and U252 (N_252,In_103,In_296);
nor U253 (N_253,In_962,In_794);
nor U254 (N_254,In_879,In_646);
nand U255 (N_255,In_665,In_154);
nor U256 (N_256,In_264,In_557);
nand U257 (N_257,In_250,In_100);
nor U258 (N_258,In_351,In_382);
nand U259 (N_259,In_696,In_178);
nor U260 (N_260,In_559,In_393);
and U261 (N_261,In_18,In_583);
nor U262 (N_262,In_574,In_531);
nand U263 (N_263,In_508,In_516);
or U264 (N_264,In_319,In_533);
nor U265 (N_265,In_434,In_948);
nor U266 (N_266,In_839,In_94);
nand U267 (N_267,In_921,In_59);
nor U268 (N_268,In_113,In_205);
or U269 (N_269,In_358,In_604);
nand U270 (N_270,In_893,In_826);
nand U271 (N_271,In_699,In_69);
nor U272 (N_272,In_39,In_25);
xor U273 (N_273,In_973,In_890);
xnor U274 (N_274,In_596,In_593);
nor U275 (N_275,In_845,In_487);
nand U276 (N_276,In_716,In_481);
xnor U277 (N_277,In_945,In_801);
or U278 (N_278,In_64,In_62);
or U279 (N_279,In_179,In_340);
or U280 (N_280,In_378,In_708);
and U281 (N_281,In_448,In_222);
xor U282 (N_282,In_798,In_754);
nand U283 (N_283,In_84,In_653);
and U284 (N_284,In_273,In_140);
nor U285 (N_285,In_56,In_330);
nor U286 (N_286,In_370,In_759);
nand U287 (N_287,In_180,In_997);
and U288 (N_288,In_161,In_464);
nand U289 (N_289,In_944,In_227);
nor U290 (N_290,In_785,In_217);
or U291 (N_291,In_725,In_492);
nor U292 (N_292,In_159,In_431);
nor U293 (N_293,In_300,In_272);
nor U294 (N_294,In_199,In_37);
and U295 (N_295,In_471,In_1);
or U296 (N_296,In_332,In_784);
or U297 (N_297,In_681,In_476);
and U298 (N_298,In_671,In_619);
nand U299 (N_299,In_95,In_594);
nand U300 (N_300,In_352,In_423);
xnor U301 (N_301,In_672,In_929);
and U302 (N_302,In_629,In_342);
nor U303 (N_303,In_375,In_409);
and U304 (N_304,In_882,In_36);
and U305 (N_305,In_726,In_863);
nor U306 (N_306,In_398,In_524);
nor U307 (N_307,In_807,In_229);
and U308 (N_308,In_359,In_57);
nor U309 (N_309,In_294,In_254);
nand U310 (N_310,In_240,In_792);
nand U311 (N_311,In_548,In_742);
xor U312 (N_312,In_831,In_462);
nor U313 (N_313,In_734,In_457);
xnor U314 (N_314,In_486,In_355);
nor U315 (N_315,In_560,In_230);
or U316 (N_316,In_265,In_967);
nand U317 (N_317,In_663,In_135);
nor U318 (N_318,In_617,In_146);
or U319 (N_319,In_959,In_413);
or U320 (N_320,In_964,In_887);
nand U321 (N_321,In_233,In_237);
xnor U322 (N_322,In_26,In_139);
xor U323 (N_323,In_765,In_7);
and U324 (N_324,In_362,In_791);
nor U325 (N_325,In_204,In_482);
or U326 (N_326,In_569,In_979);
xor U327 (N_327,In_116,In_514);
xnor U328 (N_328,In_106,In_917);
nor U329 (N_329,In_12,In_705);
and U330 (N_330,In_697,In_76);
nand U331 (N_331,In_748,In_173);
or U332 (N_332,In_682,In_453);
and U333 (N_333,In_600,In_800);
nand U334 (N_334,In_741,In_911);
nand U335 (N_335,In_939,In_852);
nor U336 (N_336,In_426,In_981);
or U337 (N_337,In_532,In_805);
nand U338 (N_338,In_465,In_630);
nor U339 (N_339,In_117,In_480);
or U340 (N_340,In_38,In_328);
nor U341 (N_341,In_551,In_518);
xor U342 (N_342,In_764,In_698);
nand U343 (N_343,In_495,In_347);
or U344 (N_344,In_558,In_904);
xor U345 (N_345,In_387,In_952);
xnor U346 (N_346,In_603,In_127);
xnor U347 (N_347,In_778,In_189);
and U348 (N_348,In_829,In_910);
or U349 (N_349,In_477,In_652);
nor U350 (N_350,In_79,In_175);
and U351 (N_351,In_424,In_983);
nand U352 (N_352,In_658,In_210);
xor U353 (N_353,In_636,In_731);
xor U354 (N_354,In_17,In_501);
nor U355 (N_355,In_577,In_228);
or U356 (N_356,In_153,In_134);
nor U357 (N_357,In_744,In_27);
nand U358 (N_358,In_111,In_170);
nor U359 (N_359,In_236,In_769);
nand U360 (N_360,In_919,In_616);
nand U361 (N_361,In_346,In_419);
nand U362 (N_362,In_60,In_213);
nor U363 (N_363,In_165,In_513);
and U364 (N_364,In_775,In_32);
nor U365 (N_365,In_896,In_410);
nand U366 (N_366,In_442,In_19);
xnor U367 (N_367,In_906,In_637);
and U368 (N_368,In_760,In_208);
and U369 (N_369,In_283,In_851);
nor U370 (N_370,In_960,In_293);
and U371 (N_371,In_715,In_850);
or U372 (N_372,In_966,In_129);
and U373 (N_373,In_638,In_223);
or U374 (N_374,In_498,In_523);
nand U375 (N_375,In_719,In_635);
nand U376 (N_376,In_238,In_502);
and U377 (N_377,In_517,In_614);
nor U378 (N_378,In_812,In_158);
xnor U379 (N_379,In_909,In_430);
or U380 (N_380,In_942,In_437);
nand U381 (N_381,In_563,In_78);
xnor U382 (N_382,In_993,In_927);
or U383 (N_383,In_803,In_155);
nor U384 (N_384,In_190,In_777);
and U385 (N_385,In_125,In_472);
and U386 (N_386,In_587,In_15);
nand U387 (N_387,In_315,In_832);
nor U388 (N_388,In_862,In_120);
and U389 (N_389,In_817,In_444);
nor U390 (N_390,In_196,In_761);
or U391 (N_391,In_354,In_786);
nor U392 (N_392,In_390,In_109);
nor U393 (N_393,In_762,In_694);
xor U394 (N_394,In_722,In_251);
or U395 (N_395,In_474,In_28);
nand U396 (N_396,In_412,In_907);
nand U397 (N_397,In_836,In_625);
or U398 (N_398,In_943,In_191);
nor U399 (N_399,In_107,In_365);
nor U400 (N_400,In_644,In_414);
nand U401 (N_401,In_819,In_723);
nand U402 (N_402,In_718,In_10);
nor U403 (N_403,In_271,In_963);
or U404 (N_404,In_737,In_455);
xnor U405 (N_405,In_350,In_415);
nor U406 (N_406,In_65,In_866);
nand U407 (N_407,In_96,In_961);
and U408 (N_408,In_519,In_87);
and U409 (N_409,In_661,In_804);
xor U410 (N_410,In_720,In_83);
xnor U411 (N_411,In_152,In_835);
nor U412 (N_412,In_888,In_232);
nand U413 (N_413,In_590,In_295);
nand U414 (N_414,In_326,In_469);
nand U415 (N_415,In_767,In_276);
or U416 (N_416,In_157,In_724);
nor U417 (N_417,In_713,In_950);
nand U418 (N_418,In_813,In_132);
nand U419 (N_419,In_174,In_483);
nor U420 (N_420,In_458,In_327);
nor U421 (N_421,In_521,In_452);
nand U422 (N_422,In_605,In_249);
and U423 (N_423,In_877,In_857);
nor U424 (N_424,In_214,In_732);
or U425 (N_425,In_747,In_395);
xnor U426 (N_426,In_224,In_401);
nor U427 (N_427,In_858,In_970);
or U428 (N_428,In_282,In_570);
or U429 (N_429,In_29,In_565);
and U430 (N_430,In_591,In_509);
nand U431 (N_431,In_640,In_257);
or U432 (N_432,In_468,In_445);
nand U433 (N_433,In_446,In_920);
xor U434 (N_434,In_871,In_611);
nor U435 (N_435,In_649,In_30);
xor U436 (N_436,In_840,In_788);
and U437 (N_437,In_515,In_825);
nor U438 (N_438,In_729,In_776);
nand U439 (N_439,In_270,In_491);
xor U440 (N_440,In_998,In_167);
xnor U441 (N_441,In_349,In_461);
xnor U442 (N_442,In_628,In_200);
nand U443 (N_443,In_16,In_932);
xor U444 (N_444,In_234,In_985);
xor U445 (N_445,In_610,In_602);
nand U446 (N_446,In_438,In_712);
xor U447 (N_447,In_544,In_400);
or U448 (N_448,In_571,In_543);
nand U449 (N_449,In_500,In_933);
or U450 (N_450,In_292,In_479);
or U451 (N_451,In_549,In_147);
and U452 (N_452,In_870,In_98);
nor U453 (N_453,In_203,In_651);
or U454 (N_454,In_859,In_745);
xor U455 (N_455,In_586,In_673);
and U456 (N_456,In_231,In_484);
xor U457 (N_457,In_873,In_377);
xnor U458 (N_458,In_384,In_957);
or U459 (N_459,In_700,In_394);
and U460 (N_460,In_899,In_266);
nor U461 (N_461,In_849,In_14);
nor U462 (N_462,In_215,In_949);
or U463 (N_463,In_164,In_537);
nand U464 (N_464,In_123,In_133);
xor U465 (N_465,In_23,In_262);
nor U466 (N_466,In_148,In_971);
xor U467 (N_467,In_162,In_193);
or U468 (N_468,In_562,In_90);
or U469 (N_469,In_128,In_606);
and U470 (N_470,In_449,In_654);
or U471 (N_471,In_567,In_988);
nor U472 (N_472,In_86,In_525);
xor U473 (N_473,In_561,In_976);
xnor U474 (N_474,In_209,In_666);
nor U475 (N_475,In_578,In_757);
xnor U476 (N_476,In_288,In_809);
nand U477 (N_477,In_421,In_864);
nand U478 (N_478,In_137,In_881);
and U479 (N_479,In_255,In_766);
nand U480 (N_480,In_925,In_5);
nand U481 (N_481,In_527,In_623);
or U482 (N_482,In_372,In_692);
or U483 (N_483,In_886,In_662);
or U484 (N_484,In_344,In_783);
nand U485 (N_485,In_818,In_506);
xor U486 (N_486,In_528,In_624);
xnor U487 (N_487,In_308,In_913);
nor U488 (N_488,In_842,In_70);
and U489 (N_489,In_878,In_252);
nor U490 (N_490,In_239,In_310);
or U491 (N_491,In_260,In_289);
nand U492 (N_492,In_397,In_688);
or U493 (N_493,In_47,In_738);
xor U494 (N_494,In_316,In_620);
and U495 (N_495,In_192,In_599);
and U496 (N_496,In_99,In_274);
xnor U497 (N_497,In_470,In_883);
and U498 (N_498,In_915,In_275);
and U499 (N_499,In_247,In_4);
xor U500 (N_500,In_297,In_237);
nand U501 (N_501,In_535,In_261);
xnor U502 (N_502,In_351,In_711);
nor U503 (N_503,In_237,In_609);
nor U504 (N_504,In_306,In_558);
or U505 (N_505,In_301,In_605);
or U506 (N_506,In_757,In_382);
or U507 (N_507,In_96,In_115);
xnor U508 (N_508,In_523,In_531);
nand U509 (N_509,In_563,In_187);
nand U510 (N_510,In_711,In_503);
xnor U511 (N_511,In_43,In_823);
and U512 (N_512,In_872,In_346);
nand U513 (N_513,In_515,In_136);
and U514 (N_514,In_824,In_280);
and U515 (N_515,In_796,In_359);
xor U516 (N_516,In_989,In_110);
or U517 (N_517,In_127,In_974);
and U518 (N_518,In_468,In_991);
nor U519 (N_519,In_992,In_611);
nand U520 (N_520,In_474,In_5);
xor U521 (N_521,In_494,In_637);
nand U522 (N_522,In_140,In_739);
xnor U523 (N_523,In_51,In_111);
or U524 (N_524,In_108,In_430);
and U525 (N_525,In_133,In_597);
or U526 (N_526,In_958,In_818);
and U527 (N_527,In_636,In_600);
nand U528 (N_528,In_479,In_343);
nand U529 (N_529,In_871,In_545);
or U530 (N_530,In_129,In_995);
or U531 (N_531,In_392,In_947);
or U532 (N_532,In_514,In_441);
nor U533 (N_533,In_742,In_184);
and U534 (N_534,In_154,In_67);
or U535 (N_535,In_519,In_950);
or U536 (N_536,In_844,In_504);
or U537 (N_537,In_247,In_623);
nor U538 (N_538,In_738,In_780);
or U539 (N_539,In_587,In_541);
xnor U540 (N_540,In_307,In_751);
xnor U541 (N_541,In_526,In_464);
and U542 (N_542,In_824,In_403);
or U543 (N_543,In_413,In_896);
xnor U544 (N_544,In_890,In_598);
nand U545 (N_545,In_612,In_516);
xor U546 (N_546,In_860,In_77);
and U547 (N_547,In_65,In_753);
xor U548 (N_548,In_385,In_2);
and U549 (N_549,In_806,In_691);
or U550 (N_550,In_340,In_317);
or U551 (N_551,In_864,In_126);
or U552 (N_552,In_798,In_724);
nor U553 (N_553,In_701,In_450);
nand U554 (N_554,In_383,In_162);
nand U555 (N_555,In_187,In_833);
or U556 (N_556,In_841,In_927);
and U557 (N_557,In_196,In_283);
nand U558 (N_558,In_801,In_971);
and U559 (N_559,In_382,In_393);
and U560 (N_560,In_465,In_390);
nor U561 (N_561,In_887,In_65);
and U562 (N_562,In_766,In_940);
or U563 (N_563,In_373,In_54);
xor U564 (N_564,In_932,In_460);
nand U565 (N_565,In_92,In_225);
xnor U566 (N_566,In_764,In_628);
nor U567 (N_567,In_717,In_312);
and U568 (N_568,In_27,In_181);
or U569 (N_569,In_731,In_901);
or U570 (N_570,In_558,In_400);
and U571 (N_571,In_728,In_646);
or U572 (N_572,In_989,In_289);
nor U573 (N_573,In_526,In_240);
xor U574 (N_574,In_103,In_917);
nand U575 (N_575,In_438,In_772);
xor U576 (N_576,In_956,In_745);
or U577 (N_577,In_936,In_895);
or U578 (N_578,In_843,In_562);
and U579 (N_579,In_950,In_119);
nand U580 (N_580,In_886,In_354);
or U581 (N_581,In_975,In_448);
xnor U582 (N_582,In_158,In_370);
and U583 (N_583,In_526,In_131);
nor U584 (N_584,In_538,In_619);
xor U585 (N_585,In_781,In_57);
nand U586 (N_586,In_883,In_986);
xnor U587 (N_587,In_22,In_462);
or U588 (N_588,In_117,In_481);
nand U589 (N_589,In_597,In_972);
or U590 (N_590,In_301,In_135);
or U591 (N_591,In_211,In_869);
nor U592 (N_592,In_657,In_762);
and U593 (N_593,In_561,In_368);
nor U594 (N_594,In_190,In_177);
xnor U595 (N_595,In_51,In_778);
nand U596 (N_596,In_211,In_74);
xor U597 (N_597,In_384,In_577);
and U598 (N_598,In_117,In_985);
nand U599 (N_599,In_889,In_182);
or U600 (N_600,In_398,In_454);
nand U601 (N_601,In_671,In_321);
xor U602 (N_602,In_534,In_648);
xnor U603 (N_603,In_199,In_866);
xor U604 (N_604,In_70,In_432);
and U605 (N_605,In_466,In_797);
and U606 (N_606,In_11,In_778);
and U607 (N_607,In_970,In_702);
nand U608 (N_608,In_717,In_287);
or U609 (N_609,In_328,In_223);
nand U610 (N_610,In_872,In_270);
or U611 (N_611,In_730,In_150);
xor U612 (N_612,In_118,In_33);
nor U613 (N_613,In_347,In_134);
and U614 (N_614,In_781,In_875);
or U615 (N_615,In_275,In_891);
nor U616 (N_616,In_805,In_850);
nor U617 (N_617,In_24,In_295);
or U618 (N_618,In_48,In_959);
nor U619 (N_619,In_431,In_55);
nor U620 (N_620,In_77,In_697);
or U621 (N_621,In_982,In_240);
nor U622 (N_622,In_985,In_761);
xor U623 (N_623,In_927,In_755);
nor U624 (N_624,In_318,In_98);
nor U625 (N_625,In_403,In_980);
and U626 (N_626,In_544,In_129);
and U627 (N_627,In_901,In_485);
xnor U628 (N_628,In_538,In_600);
nor U629 (N_629,In_824,In_230);
and U630 (N_630,In_620,In_144);
nor U631 (N_631,In_583,In_77);
xnor U632 (N_632,In_477,In_404);
xor U633 (N_633,In_1,In_205);
and U634 (N_634,In_554,In_111);
or U635 (N_635,In_741,In_506);
nor U636 (N_636,In_259,In_308);
or U637 (N_637,In_354,In_901);
xor U638 (N_638,In_324,In_163);
nor U639 (N_639,In_112,In_643);
nor U640 (N_640,In_706,In_741);
or U641 (N_641,In_218,In_497);
nand U642 (N_642,In_935,In_365);
nor U643 (N_643,In_5,In_139);
and U644 (N_644,In_128,In_995);
nor U645 (N_645,In_389,In_393);
nor U646 (N_646,In_671,In_4);
xor U647 (N_647,In_919,In_657);
and U648 (N_648,In_351,In_183);
nand U649 (N_649,In_714,In_226);
or U650 (N_650,In_688,In_379);
and U651 (N_651,In_557,In_532);
and U652 (N_652,In_211,In_445);
xnor U653 (N_653,In_692,In_353);
xnor U654 (N_654,In_280,In_382);
and U655 (N_655,In_157,In_260);
nor U656 (N_656,In_613,In_939);
and U657 (N_657,In_292,In_585);
and U658 (N_658,In_698,In_451);
and U659 (N_659,In_421,In_919);
nand U660 (N_660,In_37,In_896);
xnor U661 (N_661,In_652,In_449);
and U662 (N_662,In_183,In_395);
xnor U663 (N_663,In_720,In_748);
xnor U664 (N_664,In_471,In_44);
or U665 (N_665,In_105,In_753);
nor U666 (N_666,In_352,In_320);
nand U667 (N_667,In_683,In_327);
xnor U668 (N_668,In_747,In_934);
and U669 (N_669,In_429,In_77);
and U670 (N_670,In_63,In_808);
or U671 (N_671,In_304,In_114);
nor U672 (N_672,In_883,In_321);
nand U673 (N_673,In_358,In_209);
or U674 (N_674,In_152,In_330);
nor U675 (N_675,In_295,In_568);
nor U676 (N_676,In_228,In_466);
xor U677 (N_677,In_953,In_120);
nand U678 (N_678,In_476,In_95);
nor U679 (N_679,In_283,In_798);
and U680 (N_680,In_336,In_927);
or U681 (N_681,In_840,In_391);
and U682 (N_682,In_199,In_76);
or U683 (N_683,In_343,In_753);
xnor U684 (N_684,In_658,In_130);
nand U685 (N_685,In_653,In_896);
and U686 (N_686,In_663,In_683);
nand U687 (N_687,In_987,In_602);
xor U688 (N_688,In_860,In_753);
and U689 (N_689,In_786,In_109);
and U690 (N_690,In_30,In_505);
and U691 (N_691,In_783,In_914);
nor U692 (N_692,In_769,In_407);
or U693 (N_693,In_842,In_689);
nand U694 (N_694,In_679,In_887);
nor U695 (N_695,In_546,In_424);
xnor U696 (N_696,In_190,In_385);
and U697 (N_697,In_871,In_424);
nand U698 (N_698,In_163,In_62);
nor U699 (N_699,In_217,In_385);
and U700 (N_700,In_760,In_874);
xor U701 (N_701,In_43,In_526);
or U702 (N_702,In_97,In_236);
and U703 (N_703,In_722,In_391);
and U704 (N_704,In_901,In_83);
and U705 (N_705,In_843,In_247);
and U706 (N_706,In_793,In_336);
xor U707 (N_707,In_310,In_634);
nand U708 (N_708,In_591,In_536);
nand U709 (N_709,In_708,In_749);
nor U710 (N_710,In_528,In_130);
nand U711 (N_711,In_551,In_648);
or U712 (N_712,In_521,In_560);
xnor U713 (N_713,In_592,In_380);
nor U714 (N_714,In_433,In_949);
nor U715 (N_715,In_663,In_691);
nand U716 (N_716,In_852,In_771);
xor U717 (N_717,In_495,In_768);
nand U718 (N_718,In_726,In_482);
nor U719 (N_719,In_711,In_196);
nand U720 (N_720,In_907,In_630);
nor U721 (N_721,In_970,In_216);
nor U722 (N_722,In_788,In_870);
nand U723 (N_723,In_164,In_449);
nor U724 (N_724,In_56,In_432);
or U725 (N_725,In_61,In_659);
nand U726 (N_726,In_476,In_8);
nand U727 (N_727,In_448,In_173);
and U728 (N_728,In_376,In_875);
xnor U729 (N_729,In_449,In_313);
and U730 (N_730,In_17,In_272);
and U731 (N_731,In_985,In_539);
nand U732 (N_732,In_173,In_779);
nand U733 (N_733,In_679,In_708);
or U734 (N_734,In_136,In_147);
nor U735 (N_735,In_771,In_786);
or U736 (N_736,In_376,In_104);
xnor U737 (N_737,In_574,In_432);
or U738 (N_738,In_720,In_112);
nor U739 (N_739,In_553,In_420);
or U740 (N_740,In_553,In_362);
xor U741 (N_741,In_28,In_884);
or U742 (N_742,In_466,In_908);
and U743 (N_743,In_730,In_732);
and U744 (N_744,In_121,In_337);
nor U745 (N_745,In_591,In_92);
nor U746 (N_746,In_370,In_392);
or U747 (N_747,In_94,In_633);
nand U748 (N_748,In_396,In_793);
or U749 (N_749,In_38,In_599);
xor U750 (N_750,In_268,In_116);
nand U751 (N_751,In_187,In_526);
nand U752 (N_752,In_734,In_53);
nor U753 (N_753,In_927,In_162);
nor U754 (N_754,In_43,In_379);
nand U755 (N_755,In_243,In_993);
or U756 (N_756,In_595,In_782);
nand U757 (N_757,In_737,In_591);
xnor U758 (N_758,In_454,In_437);
or U759 (N_759,In_125,In_934);
nand U760 (N_760,In_734,In_537);
or U761 (N_761,In_78,In_514);
nor U762 (N_762,In_786,In_642);
nor U763 (N_763,In_339,In_840);
or U764 (N_764,In_919,In_67);
or U765 (N_765,In_478,In_107);
and U766 (N_766,In_330,In_928);
or U767 (N_767,In_917,In_279);
xnor U768 (N_768,In_623,In_443);
xnor U769 (N_769,In_765,In_131);
and U770 (N_770,In_423,In_547);
xnor U771 (N_771,In_572,In_374);
or U772 (N_772,In_15,In_164);
or U773 (N_773,In_674,In_541);
or U774 (N_774,In_287,In_514);
nor U775 (N_775,In_235,In_693);
and U776 (N_776,In_291,In_464);
and U777 (N_777,In_161,In_28);
nor U778 (N_778,In_932,In_782);
or U779 (N_779,In_19,In_759);
nand U780 (N_780,In_783,In_94);
xnor U781 (N_781,In_947,In_590);
nand U782 (N_782,In_585,In_520);
and U783 (N_783,In_60,In_718);
nor U784 (N_784,In_281,In_898);
nor U785 (N_785,In_277,In_274);
xor U786 (N_786,In_933,In_792);
or U787 (N_787,In_293,In_871);
or U788 (N_788,In_772,In_563);
and U789 (N_789,In_887,In_180);
or U790 (N_790,In_923,In_977);
xnor U791 (N_791,In_716,In_13);
nand U792 (N_792,In_791,In_152);
xor U793 (N_793,In_344,In_276);
and U794 (N_794,In_522,In_850);
nor U795 (N_795,In_987,In_33);
and U796 (N_796,In_91,In_886);
or U797 (N_797,In_837,In_341);
nor U798 (N_798,In_545,In_377);
xor U799 (N_799,In_354,In_16);
xnor U800 (N_800,In_20,In_647);
or U801 (N_801,In_615,In_392);
xor U802 (N_802,In_971,In_606);
nor U803 (N_803,In_481,In_511);
and U804 (N_804,In_862,In_964);
and U805 (N_805,In_143,In_35);
nor U806 (N_806,In_933,In_814);
xor U807 (N_807,In_188,In_653);
xor U808 (N_808,In_77,In_676);
nand U809 (N_809,In_736,In_30);
or U810 (N_810,In_888,In_860);
or U811 (N_811,In_17,In_724);
xor U812 (N_812,In_266,In_213);
xnor U813 (N_813,In_598,In_602);
xor U814 (N_814,In_33,In_352);
and U815 (N_815,In_207,In_629);
nor U816 (N_816,In_613,In_232);
or U817 (N_817,In_720,In_29);
xor U818 (N_818,In_368,In_793);
or U819 (N_819,In_735,In_667);
nor U820 (N_820,In_658,In_593);
or U821 (N_821,In_978,In_734);
nand U822 (N_822,In_719,In_841);
or U823 (N_823,In_154,In_421);
or U824 (N_824,In_204,In_122);
or U825 (N_825,In_530,In_131);
nor U826 (N_826,In_989,In_519);
xnor U827 (N_827,In_705,In_925);
nand U828 (N_828,In_191,In_240);
and U829 (N_829,In_576,In_663);
xnor U830 (N_830,In_862,In_546);
xnor U831 (N_831,In_854,In_94);
nor U832 (N_832,In_610,In_863);
nand U833 (N_833,In_278,In_353);
nand U834 (N_834,In_976,In_750);
or U835 (N_835,In_264,In_504);
or U836 (N_836,In_277,In_238);
nor U837 (N_837,In_35,In_582);
nand U838 (N_838,In_109,In_27);
or U839 (N_839,In_121,In_596);
xor U840 (N_840,In_316,In_141);
and U841 (N_841,In_617,In_96);
nand U842 (N_842,In_994,In_941);
or U843 (N_843,In_382,In_75);
and U844 (N_844,In_750,In_241);
and U845 (N_845,In_584,In_546);
xor U846 (N_846,In_973,In_129);
and U847 (N_847,In_391,In_843);
nand U848 (N_848,In_747,In_916);
nand U849 (N_849,In_468,In_439);
nor U850 (N_850,In_73,In_655);
or U851 (N_851,In_757,In_968);
nand U852 (N_852,In_626,In_756);
and U853 (N_853,In_918,In_381);
and U854 (N_854,In_723,In_440);
xnor U855 (N_855,In_924,In_709);
nand U856 (N_856,In_825,In_838);
and U857 (N_857,In_273,In_290);
or U858 (N_858,In_394,In_966);
nor U859 (N_859,In_790,In_356);
nand U860 (N_860,In_757,In_735);
and U861 (N_861,In_694,In_308);
nand U862 (N_862,In_609,In_57);
nor U863 (N_863,In_666,In_647);
and U864 (N_864,In_574,In_263);
xnor U865 (N_865,In_273,In_352);
xnor U866 (N_866,In_319,In_517);
or U867 (N_867,In_434,In_241);
or U868 (N_868,In_432,In_169);
nand U869 (N_869,In_286,In_704);
xnor U870 (N_870,In_606,In_310);
or U871 (N_871,In_553,In_10);
nor U872 (N_872,In_695,In_256);
and U873 (N_873,In_529,In_663);
xor U874 (N_874,In_22,In_528);
nand U875 (N_875,In_123,In_420);
or U876 (N_876,In_109,In_458);
and U877 (N_877,In_620,In_103);
nand U878 (N_878,In_266,In_301);
nor U879 (N_879,In_649,In_777);
or U880 (N_880,In_949,In_18);
xnor U881 (N_881,In_540,In_937);
xor U882 (N_882,In_43,In_1);
or U883 (N_883,In_405,In_479);
and U884 (N_884,In_479,In_955);
or U885 (N_885,In_874,In_637);
and U886 (N_886,In_288,In_2);
xor U887 (N_887,In_269,In_600);
nor U888 (N_888,In_33,In_256);
or U889 (N_889,In_885,In_883);
and U890 (N_890,In_873,In_823);
or U891 (N_891,In_116,In_925);
xnor U892 (N_892,In_995,In_979);
nand U893 (N_893,In_806,In_437);
nor U894 (N_894,In_626,In_699);
and U895 (N_895,In_861,In_407);
nand U896 (N_896,In_704,In_556);
nand U897 (N_897,In_954,In_965);
and U898 (N_898,In_582,In_325);
nand U899 (N_899,In_412,In_103);
or U900 (N_900,In_516,In_159);
and U901 (N_901,In_496,In_131);
or U902 (N_902,In_487,In_492);
xor U903 (N_903,In_230,In_126);
xnor U904 (N_904,In_98,In_510);
or U905 (N_905,In_639,In_533);
nor U906 (N_906,In_99,In_273);
and U907 (N_907,In_370,In_765);
xor U908 (N_908,In_906,In_141);
nor U909 (N_909,In_86,In_365);
xor U910 (N_910,In_621,In_532);
nand U911 (N_911,In_784,In_599);
nor U912 (N_912,In_309,In_919);
and U913 (N_913,In_642,In_659);
nand U914 (N_914,In_605,In_697);
nor U915 (N_915,In_122,In_551);
nand U916 (N_916,In_958,In_324);
or U917 (N_917,In_263,In_514);
and U918 (N_918,In_631,In_722);
nand U919 (N_919,In_748,In_617);
or U920 (N_920,In_96,In_338);
nor U921 (N_921,In_905,In_199);
nand U922 (N_922,In_363,In_376);
nand U923 (N_923,In_476,In_67);
or U924 (N_924,In_136,In_565);
xnor U925 (N_925,In_487,In_905);
and U926 (N_926,In_947,In_984);
and U927 (N_927,In_855,In_526);
xnor U928 (N_928,In_966,In_566);
nor U929 (N_929,In_854,In_717);
nand U930 (N_930,In_483,In_668);
nor U931 (N_931,In_420,In_915);
nand U932 (N_932,In_95,In_428);
and U933 (N_933,In_215,In_749);
xnor U934 (N_934,In_169,In_896);
or U935 (N_935,In_479,In_173);
or U936 (N_936,In_818,In_778);
and U937 (N_937,In_152,In_214);
nor U938 (N_938,In_960,In_688);
nor U939 (N_939,In_263,In_303);
nor U940 (N_940,In_172,In_908);
xnor U941 (N_941,In_251,In_471);
nand U942 (N_942,In_209,In_575);
xor U943 (N_943,In_745,In_954);
nand U944 (N_944,In_814,In_145);
and U945 (N_945,In_42,In_644);
nor U946 (N_946,In_556,In_837);
or U947 (N_947,In_903,In_262);
or U948 (N_948,In_300,In_52);
and U949 (N_949,In_681,In_46);
nor U950 (N_950,In_687,In_215);
or U951 (N_951,In_921,In_956);
and U952 (N_952,In_831,In_914);
and U953 (N_953,In_67,In_751);
xor U954 (N_954,In_837,In_826);
or U955 (N_955,In_73,In_711);
nor U956 (N_956,In_389,In_49);
xor U957 (N_957,In_863,In_847);
and U958 (N_958,In_879,In_57);
nand U959 (N_959,In_922,In_499);
nand U960 (N_960,In_98,In_91);
nor U961 (N_961,In_131,In_775);
xor U962 (N_962,In_315,In_546);
or U963 (N_963,In_801,In_700);
or U964 (N_964,In_77,In_883);
or U965 (N_965,In_496,In_631);
xnor U966 (N_966,In_51,In_133);
nand U967 (N_967,In_306,In_690);
and U968 (N_968,In_18,In_56);
or U969 (N_969,In_62,In_288);
nor U970 (N_970,In_821,In_757);
xor U971 (N_971,In_45,In_378);
nand U972 (N_972,In_3,In_794);
or U973 (N_973,In_664,In_107);
nor U974 (N_974,In_87,In_969);
or U975 (N_975,In_699,In_438);
nand U976 (N_976,In_499,In_669);
xnor U977 (N_977,In_558,In_425);
nor U978 (N_978,In_746,In_884);
nand U979 (N_979,In_849,In_23);
xnor U980 (N_980,In_122,In_769);
or U981 (N_981,In_609,In_464);
xor U982 (N_982,In_722,In_759);
xor U983 (N_983,In_184,In_540);
or U984 (N_984,In_481,In_256);
and U985 (N_985,In_161,In_790);
nand U986 (N_986,In_222,In_921);
xor U987 (N_987,In_704,In_737);
or U988 (N_988,In_187,In_509);
nor U989 (N_989,In_471,In_946);
or U990 (N_990,In_665,In_362);
nand U991 (N_991,In_622,In_544);
or U992 (N_992,In_39,In_786);
xor U993 (N_993,In_751,In_485);
nand U994 (N_994,In_565,In_304);
nand U995 (N_995,In_47,In_739);
nor U996 (N_996,In_356,In_216);
nand U997 (N_997,In_371,In_967);
or U998 (N_998,In_31,In_197);
nand U999 (N_999,In_570,In_606);
and U1000 (N_1000,N_700,N_292);
nor U1001 (N_1001,N_870,N_629);
xnor U1002 (N_1002,N_798,N_876);
nand U1003 (N_1003,N_571,N_432);
or U1004 (N_1004,N_163,N_557);
nand U1005 (N_1005,N_827,N_142);
xor U1006 (N_1006,N_754,N_134);
and U1007 (N_1007,N_31,N_608);
or U1008 (N_1008,N_200,N_756);
xor U1009 (N_1009,N_941,N_990);
nor U1010 (N_1010,N_179,N_121);
nor U1011 (N_1011,N_467,N_901);
xor U1012 (N_1012,N_935,N_391);
xnor U1013 (N_1013,N_795,N_581);
nor U1014 (N_1014,N_528,N_748);
and U1015 (N_1015,N_372,N_466);
or U1016 (N_1016,N_360,N_994);
and U1017 (N_1017,N_989,N_757);
nor U1018 (N_1018,N_797,N_921);
xnor U1019 (N_1019,N_423,N_913);
and U1020 (N_1020,N_553,N_868);
or U1021 (N_1021,N_667,N_633);
nor U1022 (N_1022,N_185,N_957);
nand U1023 (N_1023,N_315,N_118);
nand U1024 (N_1024,N_353,N_916);
xnor U1025 (N_1025,N_461,N_894);
and U1026 (N_1026,N_739,N_320);
or U1027 (N_1027,N_44,N_815);
or U1028 (N_1028,N_129,N_313);
or U1029 (N_1029,N_279,N_7);
nor U1030 (N_1030,N_49,N_211);
and U1031 (N_1031,N_769,N_305);
nor U1032 (N_1032,N_25,N_672);
and U1033 (N_1033,N_737,N_294);
nand U1034 (N_1034,N_144,N_693);
nor U1035 (N_1035,N_782,N_920);
xnor U1036 (N_1036,N_540,N_763);
nand U1037 (N_1037,N_176,N_366);
or U1038 (N_1038,N_61,N_337);
xor U1039 (N_1039,N_70,N_555);
nand U1040 (N_1040,N_60,N_310);
or U1041 (N_1041,N_548,N_250);
and U1042 (N_1042,N_547,N_848);
nand U1043 (N_1043,N_900,N_355);
or U1044 (N_1044,N_114,N_836);
nor U1045 (N_1045,N_962,N_233);
or U1046 (N_1046,N_945,N_488);
xnor U1047 (N_1047,N_450,N_597);
and U1048 (N_1048,N_460,N_860);
and U1049 (N_1049,N_733,N_958);
or U1050 (N_1050,N_1,N_255);
nand U1051 (N_1051,N_172,N_568);
nand U1052 (N_1052,N_10,N_670);
xor U1053 (N_1053,N_59,N_646);
or U1054 (N_1054,N_671,N_569);
or U1055 (N_1055,N_874,N_277);
nor U1056 (N_1056,N_83,N_468);
xnor U1057 (N_1057,N_253,N_993);
xnor U1058 (N_1058,N_194,N_768);
nand U1059 (N_1059,N_418,N_611);
and U1060 (N_1060,N_58,N_985);
nand U1061 (N_1061,N_19,N_486);
nand U1062 (N_1062,N_284,N_231);
and U1063 (N_1063,N_412,N_323);
and U1064 (N_1064,N_834,N_546);
and U1065 (N_1065,N_377,N_598);
nand U1066 (N_1066,N_524,N_496);
or U1067 (N_1067,N_765,N_147);
nor U1068 (N_1068,N_724,N_708);
nor U1069 (N_1069,N_182,N_838);
and U1070 (N_1070,N_312,N_544);
and U1071 (N_1071,N_531,N_186);
and U1072 (N_1072,N_961,N_203);
xnor U1073 (N_1073,N_744,N_12);
nand U1074 (N_1074,N_3,N_660);
xor U1075 (N_1075,N_183,N_793);
xnor U1076 (N_1076,N_862,N_959);
nand U1077 (N_1077,N_923,N_563);
xnor U1078 (N_1078,N_878,N_518);
xor U1079 (N_1079,N_499,N_251);
or U1080 (N_1080,N_706,N_191);
and U1081 (N_1081,N_813,N_394);
and U1082 (N_1082,N_601,N_615);
or U1083 (N_1083,N_164,N_529);
nand U1084 (N_1084,N_302,N_583);
and U1085 (N_1085,N_227,N_324);
or U1086 (N_1086,N_88,N_367);
nor U1087 (N_1087,N_566,N_788);
nor U1088 (N_1088,N_833,N_866);
or U1089 (N_1089,N_831,N_687);
and U1090 (N_1090,N_462,N_967);
and U1091 (N_1091,N_770,N_791);
xnor U1092 (N_1092,N_396,N_623);
xnor U1093 (N_1093,N_287,N_382);
nor U1094 (N_1094,N_283,N_910);
nor U1095 (N_1095,N_802,N_361);
xnor U1096 (N_1096,N_812,N_30);
nor U1097 (N_1097,N_398,N_713);
nand U1098 (N_1098,N_475,N_166);
nor U1099 (N_1099,N_86,N_966);
nand U1100 (N_1100,N_71,N_95);
or U1101 (N_1101,N_861,N_259);
nor U1102 (N_1102,N_918,N_573);
and U1103 (N_1103,N_123,N_787);
nor U1104 (N_1104,N_170,N_112);
xnor U1105 (N_1105,N_663,N_556);
or U1106 (N_1106,N_652,N_120);
nor U1107 (N_1107,N_839,N_18);
nor U1108 (N_1108,N_968,N_909);
xor U1109 (N_1109,N_697,N_371);
nor U1110 (N_1110,N_998,N_469);
nand U1111 (N_1111,N_976,N_745);
xor U1112 (N_1112,N_425,N_258);
xor U1113 (N_1113,N_606,N_657);
and U1114 (N_1114,N_677,N_773);
or U1115 (N_1115,N_380,N_806);
nand U1116 (N_1116,N_932,N_110);
nor U1117 (N_1117,N_379,N_4);
or U1118 (N_1118,N_722,N_109);
xnor U1119 (N_1119,N_960,N_479);
xnor U1120 (N_1120,N_193,N_625);
nand U1121 (N_1121,N_665,N_300);
and U1122 (N_1122,N_175,N_607);
nor U1123 (N_1123,N_153,N_133);
nor U1124 (N_1124,N_94,N_810);
and U1125 (N_1125,N_653,N_429);
xnor U1126 (N_1126,N_593,N_707);
and U1127 (N_1127,N_942,N_232);
or U1128 (N_1128,N_319,N_991);
and U1129 (N_1129,N_458,N_220);
and U1130 (N_1130,N_871,N_330);
or U1131 (N_1131,N_326,N_113);
or U1132 (N_1132,N_456,N_442);
or U1133 (N_1133,N_417,N_214);
xnor U1134 (N_1134,N_198,N_638);
nor U1135 (N_1135,N_542,N_634);
and U1136 (N_1136,N_914,N_406);
or U1137 (N_1137,N_775,N_507);
and U1138 (N_1138,N_244,N_883);
nor U1139 (N_1139,N_24,N_951);
xor U1140 (N_1140,N_459,N_222);
nand U1141 (N_1141,N_753,N_619);
xnor U1142 (N_1142,N_735,N_141);
nand U1143 (N_1143,N_307,N_599);
or U1144 (N_1144,N_241,N_221);
and U1145 (N_1145,N_579,N_308);
xor U1146 (N_1146,N_558,N_661);
or U1147 (N_1147,N_26,N_872);
nand U1148 (N_1148,N_216,N_481);
xnor U1149 (N_1149,N_627,N_239);
nor U1150 (N_1150,N_23,N_851);
or U1151 (N_1151,N_595,N_956);
or U1152 (N_1152,N_74,N_201);
xnor U1153 (N_1153,N_946,N_45);
nand U1154 (N_1154,N_158,N_917);
nor U1155 (N_1155,N_281,N_487);
and U1156 (N_1156,N_290,N_13);
nor U1157 (N_1157,N_699,N_195);
nor U1158 (N_1158,N_617,N_602);
xor U1159 (N_1159,N_14,N_694);
nand U1160 (N_1160,N_386,N_342);
nand U1161 (N_1161,N_730,N_40);
and U1162 (N_1162,N_919,N_6);
xnor U1163 (N_1163,N_647,N_322);
xnor U1164 (N_1164,N_63,N_278);
nor U1165 (N_1165,N_20,N_740);
xnor U1166 (N_1166,N_734,N_64);
and U1167 (N_1167,N_422,N_226);
nor U1168 (N_1168,N_156,N_676);
nand U1169 (N_1169,N_902,N_38);
or U1170 (N_1170,N_410,N_952);
nor U1171 (N_1171,N_750,N_317);
or U1172 (N_1172,N_318,N_280);
or U1173 (N_1173,N_344,N_424);
nor U1174 (N_1174,N_438,N_115);
xnor U1175 (N_1175,N_476,N_718);
nand U1176 (N_1176,N_828,N_329);
xnor U1177 (N_1177,N_760,N_364);
and U1178 (N_1178,N_349,N_358);
nor U1179 (N_1179,N_137,N_580);
and U1180 (N_1180,N_35,N_297);
and U1181 (N_1181,N_403,N_247);
nor U1182 (N_1182,N_855,N_873);
nor U1183 (N_1183,N_685,N_983);
and U1184 (N_1184,N_65,N_347);
or U1185 (N_1185,N_149,N_173);
nand U1186 (N_1186,N_41,N_345);
nand U1187 (N_1187,N_363,N_373);
xnor U1188 (N_1188,N_965,N_435);
nand U1189 (N_1189,N_314,N_742);
or U1190 (N_1190,N_774,N_844);
xnor U1191 (N_1191,N_343,N_260);
xnor U1192 (N_1192,N_464,N_949);
and U1193 (N_1193,N_446,N_819);
and U1194 (N_1194,N_0,N_645);
or U1195 (N_1195,N_354,N_911);
xnor U1196 (N_1196,N_263,N_511);
nand U1197 (N_1197,N_230,N_554);
nor U1198 (N_1198,N_891,N_440);
xor U1199 (N_1199,N_882,N_881);
or U1200 (N_1200,N_289,N_180);
xor U1201 (N_1201,N_631,N_275);
nand U1202 (N_1202,N_189,N_513);
nor U1203 (N_1203,N_493,N_605);
xor U1204 (N_1204,N_937,N_789);
nand U1205 (N_1205,N_817,N_145);
or U1206 (N_1206,N_545,N_178);
and U1207 (N_1207,N_659,N_565);
nor U1208 (N_1208,N_161,N_8);
or U1209 (N_1209,N_421,N_577);
nor U1210 (N_1210,N_784,N_519);
nand U1211 (N_1211,N_217,N_254);
xor U1212 (N_1212,N_332,N_96);
xor U1213 (N_1213,N_840,N_471);
nand U1214 (N_1214,N_111,N_779);
or U1215 (N_1215,N_311,N_738);
nor U1216 (N_1216,N_240,N_76);
nand U1217 (N_1217,N_262,N_726);
nor U1218 (N_1218,N_139,N_155);
and U1219 (N_1219,N_944,N_29);
nor U1220 (N_1220,N_494,N_437);
or U1221 (N_1221,N_22,N_538);
xor U1222 (N_1222,N_15,N_288);
xnor U1223 (N_1223,N_490,N_441);
nand U1224 (N_1224,N_751,N_979);
or U1225 (N_1225,N_238,N_741);
nand U1226 (N_1226,N_613,N_954);
xnor U1227 (N_1227,N_395,N_409);
nor U1228 (N_1228,N_904,N_624);
nand U1229 (N_1229,N_808,N_703);
nand U1230 (N_1230,N_209,N_841);
nand U1231 (N_1231,N_340,N_938);
xnor U1232 (N_1232,N_37,N_357);
nand U1233 (N_1233,N_626,N_430);
xor U1234 (N_1234,N_167,N_886);
nand U1235 (N_1235,N_505,N_451);
or U1236 (N_1236,N_963,N_261);
nand U1237 (N_1237,N_341,N_333);
nor U1238 (N_1238,N_835,N_489);
nor U1239 (N_1239,N_478,N_912);
nor U1240 (N_1240,N_400,N_809);
nor U1241 (N_1241,N_375,N_897);
xor U1242 (N_1242,N_522,N_541);
nor U1243 (N_1243,N_614,N_272);
nor U1244 (N_1244,N_908,N_483);
xor U1245 (N_1245,N_778,N_235);
nor U1246 (N_1246,N_717,N_397);
and U1247 (N_1247,N_591,N_863);
and U1248 (N_1248,N_427,N_526);
nand U1249 (N_1249,N_82,N_887);
and U1250 (N_1250,N_762,N_160);
nand U1251 (N_1251,N_445,N_621);
and U1252 (N_1252,N_560,N_858);
nand U1253 (N_1253,N_732,N_925);
nor U1254 (N_1254,N_759,N_184);
or U1255 (N_1255,N_299,N_130);
nand U1256 (N_1256,N_316,N_950);
xor U1257 (N_1257,N_953,N_169);
and U1258 (N_1258,N_727,N_988);
and U1259 (N_1259,N_271,N_236);
and U1260 (N_1260,N_504,N_704);
nor U1261 (N_1261,N_684,N_245);
xnor U1262 (N_1262,N_673,N_492);
nand U1263 (N_1263,N_721,N_895);
and U1264 (N_1264,N_80,N_928);
xor U1265 (N_1265,N_594,N_924);
nor U1266 (N_1266,N_470,N_69);
and U1267 (N_1267,N_55,N_482);
or U1268 (N_1268,N_87,N_208);
or U1269 (N_1269,N_196,N_274);
or U1270 (N_1270,N_36,N_68);
nor U1271 (N_1271,N_535,N_890);
xnor U1272 (N_1272,N_777,N_749);
or U1273 (N_1273,N_800,N_273);
nor U1274 (N_1274,N_683,N_512);
and U1275 (N_1275,N_766,N_413);
nand U1276 (N_1276,N_402,N_509);
nor U1277 (N_1277,N_502,N_365);
and U1278 (N_1278,N_119,N_869);
nor U1279 (N_1279,N_428,N_306);
nor U1280 (N_1280,N_567,N_335);
nand U1281 (N_1281,N_643,N_92);
or U1282 (N_1282,N_596,N_588);
xnor U1283 (N_1283,N_856,N_688);
nor U1284 (N_1284,N_472,N_501);
and U1285 (N_1285,N_640,N_885);
or U1286 (N_1286,N_690,N_116);
and U1287 (N_1287,N_215,N_62);
nor U1288 (N_1288,N_162,N_151);
xnor U1289 (N_1289,N_709,N_830);
xor U1290 (N_1290,N_39,N_219);
or U1291 (N_1291,N_971,N_140);
or U1292 (N_1292,N_651,N_586);
or U1293 (N_1293,N_257,N_552);
nand U1294 (N_1294,N_204,N_940);
xor U1295 (N_1295,N_934,N_414);
or U1296 (N_1296,N_896,N_117);
and U1297 (N_1297,N_843,N_992);
or U1298 (N_1298,N_525,N_712);
or U1299 (N_1299,N_385,N_801);
nand U1300 (N_1300,N_491,N_33);
nand U1301 (N_1301,N_845,N_783);
nand U1302 (N_1302,N_237,N_936);
or U1303 (N_1303,N_575,N_54);
nand U1304 (N_1304,N_407,N_411);
and U1305 (N_1305,N_105,N_996);
and U1306 (N_1306,N_269,N_537);
and U1307 (N_1307,N_678,N_658);
nand U1308 (N_1308,N_559,N_223);
nand U1309 (N_1309,N_229,N_197);
nor U1310 (N_1310,N_85,N_202);
xnor U1311 (N_1311,N_81,N_346);
xnor U1312 (N_1312,N_212,N_867);
nor U1313 (N_1313,N_649,N_154);
and U1314 (N_1314,N_695,N_419);
nor U1315 (N_1315,N_943,N_587);
nor U1316 (N_1316,N_510,N_715);
and U1317 (N_1317,N_561,N_157);
xor U1318 (N_1318,N_136,N_731);
nand U1319 (N_1319,N_929,N_285);
or U1320 (N_1320,N_11,N_906);
xnor U1321 (N_1321,N_321,N_293);
xor U1322 (N_1322,N_656,N_820);
nor U1323 (N_1323,N_648,N_523);
nor U1324 (N_1324,N_102,N_73);
nor U1325 (N_1325,N_234,N_600);
and U1326 (N_1326,N_439,N_997);
nand U1327 (N_1327,N_837,N_388);
nor U1328 (N_1328,N_101,N_381);
nand U1329 (N_1329,N_348,N_865);
nand U1330 (N_1330,N_148,N_691);
xnor U1331 (N_1331,N_705,N_804);
and U1332 (N_1332,N_662,N_852);
nor U1333 (N_1333,N_805,N_97);
xor U1334 (N_1334,N_696,N_228);
nand U1335 (N_1335,N_609,N_964);
nand U1336 (N_1336,N_449,N_604);
and U1337 (N_1337,N_893,N_256);
nor U1338 (N_1338,N_986,N_666);
xor U1339 (N_1339,N_796,N_584);
nor U1340 (N_1340,N_108,N_159);
or U1341 (N_1341,N_821,N_453);
nand U1342 (N_1342,N_53,N_521);
nor U1343 (N_1343,N_826,N_17);
and U1344 (N_1344,N_686,N_905);
or U1345 (N_1345,N_814,N_399);
nand U1346 (N_1346,N_444,N_455);
xor U1347 (N_1347,N_420,N_104);
nand U1348 (N_1348,N_84,N_811);
nand U1349 (N_1349,N_714,N_338);
xor U1350 (N_1350,N_824,N_125);
or U1351 (N_1351,N_150,N_792);
nand U1352 (N_1352,N_295,N_847);
and U1353 (N_1353,N_850,N_463);
or U1354 (N_1354,N_79,N_574);
nor U1355 (N_1355,N_99,N_100);
nand U1356 (N_1356,N_374,N_975);
nand U1357 (N_1357,N_34,N_842);
or U1358 (N_1358,N_589,N_880);
or U1359 (N_1359,N_131,N_630);
or U1360 (N_1360,N_276,N_576);
nand U1361 (N_1361,N_642,N_972);
and U1362 (N_1362,N_761,N_127);
nand U1363 (N_1363,N_610,N_978);
nand U1364 (N_1364,N_508,N_415);
nand U1365 (N_1365,N_585,N_416);
nor U1366 (N_1366,N_447,N_889);
xor U1367 (N_1367,N_701,N_551);
xnor U1368 (N_1368,N_168,N_359);
nor U1369 (N_1369,N_764,N_785);
nand U1370 (N_1370,N_454,N_165);
or U1371 (N_1371,N_426,N_75);
and U1372 (N_1372,N_644,N_225);
xor U1373 (N_1373,N_641,N_362);
nand U1374 (N_1374,N_875,N_915);
and U1375 (N_1375,N_816,N_803);
nand U1376 (N_1376,N_78,N_864);
xor U1377 (N_1377,N_603,N_698);
xnor U1378 (N_1378,N_533,N_72);
nor U1379 (N_1379,N_368,N_128);
and U1380 (N_1380,N_689,N_632);
and U1381 (N_1381,N_922,N_590);
nand U1382 (N_1382,N_520,N_46);
nor U1383 (N_1383,N_190,N_433);
or U1384 (N_1384,N_434,N_387);
nand U1385 (N_1385,N_794,N_243);
xor U1386 (N_1386,N_16,N_825);
nor U1387 (N_1387,N_723,N_622);
xnor U1388 (N_1388,N_484,N_664);
and U1389 (N_1389,N_199,N_242);
nor U1390 (N_1390,N_654,N_296);
xor U1391 (N_1391,N_171,N_376);
or U1392 (N_1392,N_716,N_47);
nand U1393 (N_1393,N_530,N_669);
and U1394 (N_1394,N_77,N_500);
nand U1395 (N_1395,N_452,N_485);
xnor U1396 (N_1396,N_974,N_680);
nand U1397 (N_1397,N_729,N_970);
nand U1398 (N_1398,N_350,N_668);
or U1399 (N_1399,N_213,N_618);
xnor U1400 (N_1400,N_246,N_331);
or U1401 (N_1401,N_582,N_532);
and U1402 (N_1402,N_612,N_877);
xnor U1403 (N_1403,N_383,N_857);
or U1404 (N_1404,N_752,N_898);
xnor U1405 (N_1405,N_899,N_549);
xnor U1406 (N_1406,N_67,N_517);
nand U1407 (N_1407,N_572,N_931);
xnor U1408 (N_1408,N_27,N_93);
nor U1409 (N_1409,N_465,N_772);
or U1410 (N_1410,N_682,N_408);
or U1411 (N_1411,N_564,N_736);
nand U1412 (N_1412,N_720,N_135);
or U1413 (N_1413,N_301,N_635);
or U1414 (N_1414,N_431,N_152);
xor U1415 (N_1415,N_981,N_710);
and U1416 (N_1416,N_448,N_252);
and U1417 (N_1417,N_270,N_9);
or U1418 (N_1418,N_711,N_980);
xnor U1419 (N_1419,N_205,N_639);
nor U1420 (N_1420,N_401,N_702);
or U1421 (N_1421,N_473,N_771);
nand U1422 (N_1422,N_98,N_674);
nand U1423 (N_1423,N_933,N_90);
nand U1424 (N_1424,N_999,N_309);
nand U1425 (N_1425,N_984,N_282);
nor U1426 (N_1426,N_498,N_336);
and U1427 (N_1427,N_743,N_210);
nand U1428 (N_1428,N_298,N_495);
or U1429 (N_1429,N_352,N_822);
and U1430 (N_1430,N_370,N_405);
nor U1431 (N_1431,N_977,N_903);
or U1432 (N_1432,N_268,N_267);
xnor U1433 (N_1433,N_188,N_807);
nor U1434 (N_1434,N_955,N_248);
nor U1435 (N_1435,N_143,N_28);
xnor U1436 (N_1436,N_786,N_107);
xor U1437 (N_1437,N_728,N_393);
or U1438 (N_1438,N_206,N_303);
xor U1439 (N_1439,N_5,N_832);
or U1440 (N_1440,N_43,N_21);
or U1441 (N_1441,N_679,N_390);
and U1442 (N_1442,N_879,N_457);
and U1443 (N_1443,N_746,N_369);
nand U1444 (N_1444,N_799,N_146);
or U1445 (N_1445,N_536,N_973);
nand U1446 (N_1446,N_218,N_356);
xnor U1447 (N_1447,N_888,N_42);
nor U1448 (N_1448,N_747,N_52);
xnor U1449 (N_1449,N_907,N_132);
or U1450 (N_1450,N_91,N_692);
and U1451 (N_1451,N_550,N_474);
and U1452 (N_1452,N_2,N_948);
nand U1453 (N_1453,N_719,N_181);
nor U1454 (N_1454,N_404,N_304);
or U1455 (N_1455,N_818,N_334);
and U1456 (N_1456,N_939,N_637);
and U1457 (N_1457,N_534,N_384);
nand U1458 (N_1458,N_514,N_539);
xor U1459 (N_1459,N_655,N_291);
xnor U1460 (N_1460,N_327,N_995);
nand U1461 (N_1461,N_174,N_392);
or U1462 (N_1462,N_325,N_767);
and U1463 (N_1463,N_286,N_628);
nor U1464 (N_1464,N_264,N_378);
or U1465 (N_1465,N_650,N_266);
and U1466 (N_1466,N_497,N_616);
nand U1467 (N_1467,N_106,N_339);
nand U1468 (N_1468,N_829,N_636);
and U1469 (N_1469,N_56,N_477);
nand U1470 (N_1470,N_122,N_562);
or U1471 (N_1471,N_592,N_328);
xnor U1472 (N_1472,N_50,N_138);
and U1473 (N_1473,N_48,N_776);
or U1474 (N_1474,N_681,N_207);
xor U1475 (N_1475,N_480,N_124);
and U1476 (N_1476,N_51,N_436);
or U1477 (N_1477,N_755,N_192);
and U1478 (N_1478,N_947,N_892);
and U1479 (N_1479,N_351,N_823);
and U1480 (N_1480,N_126,N_506);
nor U1481 (N_1481,N_849,N_570);
xnor U1482 (N_1482,N_969,N_790);
xnor U1483 (N_1483,N_89,N_57);
or U1484 (N_1484,N_265,N_853);
xor U1485 (N_1485,N_884,N_854);
nor U1486 (N_1486,N_249,N_503);
and U1487 (N_1487,N_846,N_926);
or U1488 (N_1488,N_515,N_927);
and U1489 (N_1489,N_224,N_177);
nor U1490 (N_1490,N_930,N_725);
or U1491 (N_1491,N_859,N_758);
or U1492 (N_1492,N_516,N_780);
and U1493 (N_1493,N_66,N_187);
and U1494 (N_1494,N_543,N_32);
or U1495 (N_1495,N_389,N_527);
xnor U1496 (N_1496,N_675,N_443);
nor U1497 (N_1497,N_982,N_578);
and U1498 (N_1498,N_781,N_620);
or U1499 (N_1499,N_103,N_987);
or U1500 (N_1500,N_123,N_85);
and U1501 (N_1501,N_255,N_693);
or U1502 (N_1502,N_300,N_361);
nor U1503 (N_1503,N_284,N_361);
nand U1504 (N_1504,N_240,N_970);
or U1505 (N_1505,N_224,N_23);
and U1506 (N_1506,N_302,N_670);
and U1507 (N_1507,N_484,N_341);
or U1508 (N_1508,N_403,N_314);
and U1509 (N_1509,N_149,N_221);
nor U1510 (N_1510,N_540,N_450);
or U1511 (N_1511,N_600,N_971);
nor U1512 (N_1512,N_858,N_698);
nand U1513 (N_1513,N_705,N_780);
xnor U1514 (N_1514,N_505,N_904);
and U1515 (N_1515,N_406,N_224);
or U1516 (N_1516,N_393,N_596);
and U1517 (N_1517,N_22,N_117);
nor U1518 (N_1518,N_33,N_138);
and U1519 (N_1519,N_449,N_458);
nor U1520 (N_1520,N_628,N_126);
nand U1521 (N_1521,N_249,N_24);
or U1522 (N_1522,N_766,N_556);
or U1523 (N_1523,N_199,N_339);
xnor U1524 (N_1524,N_962,N_546);
xnor U1525 (N_1525,N_856,N_598);
nor U1526 (N_1526,N_388,N_622);
or U1527 (N_1527,N_611,N_525);
or U1528 (N_1528,N_586,N_483);
xnor U1529 (N_1529,N_422,N_118);
xnor U1530 (N_1530,N_167,N_54);
nand U1531 (N_1531,N_308,N_552);
nor U1532 (N_1532,N_764,N_997);
xnor U1533 (N_1533,N_570,N_46);
nand U1534 (N_1534,N_209,N_183);
xor U1535 (N_1535,N_746,N_403);
nand U1536 (N_1536,N_691,N_329);
or U1537 (N_1537,N_84,N_936);
nor U1538 (N_1538,N_192,N_716);
xor U1539 (N_1539,N_666,N_723);
nor U1540 (N_1540,N_316,N_2);
nor U1541 (N_1541,N_894,N_703);
nand U1542 (N_1542,N_75,N_388);
nor U1543 (N_1543,N_860,N_642);
nand U1544 (N_1544,N_552,N_563);
and U1545 (N_1545,N_416,N_293);
xnor U1546 (N_1546,N_98,N_177);
nand U1547 (N_1547,N_916,N_278);
or U1548 (N_1548,N_38,N_225);
or U1549 (N_1549,N_609,N_101);
xor U1550 (N_1550,N_784,N_832);
xnor U1551 (N_1551,N_53,N_866);
nand U1552 (N_1552,N_109,N_861);
or U1553 (N_1553,N_781,N_88);
and U1554 (N_1554,N_772,N_602);
and U1555 (N_1555,N_976,N_798);
and U1556 (N_1556,N_626,N_665);
or U1557 (N_1557,N_605,N_472);
or U1558 (N_1558,N_225,N_597);
or U1559 (N_1559,N_296,N_268);
and U1560 (N_1560,N_362,N_866);
nor U1561 (N_1561,N_253,N_827);
nand U1562 (N_1562,N_107,N_422);
nor U1563 (N_1563,N_694,N_883);
or U1564 (N_1564,N_472,N_77);
nor U1565 (N_1565,N_531,N_446);
nand U1566 (N_1566,N_272,N_857);
xor U1567 (N_1567,N_78,N_86);
xor U1568 (N_1568,N_930,N_436);
nand U1569 (N_1569,N_880,N_381);
nand U1570 (N_1570,N_702,N_515);
or U1571 (N_1571,N_994,N_462);
and U1572 (N_1572,N_80,N_459);
or U1573 (N_1573,N_120,N_758);
xnor U1574 (N_1574,N_801,N_498);
nor U1575 (N_1575,N_308,N_164);
and U1576 (N_1576,N_818,N_288);
nor U1577 (N_1577,N_300,N_576);
xor U1578 (N_1578,N_491,N_996);
xnor U1579 (N_1579,N_69,N_605);
or U1580 (N_1580,N_934,N_136);
or U1581 (N_1581,N_268,N_913);
and U1582 (N_1582,N_450,N_362);
or U1583 (N_1583,N_417,N_466);
xor U1584 (N_1584,N_978,N_907);
and U1585 (N_1585,N_268,N_721);
xor U1586 (N_1586,N_639,N_953);
nor U1587 (N_1587,N_919,N_374);
and U1588 (N_1588,N_81,N_114);
nor U1589 (N_1589,N_450,N_946);
and U1590 (N_1590,N_311,N_706);
or U1591 (N_1591,N_405,N_658);
and U1592 (N_1592,N_169,N_283);
and U1593 (N_1593,N_719,N_510);
or U1594 (N_1594,N_129,N_89);
and U1595 (N_1595,N_405,N_286);
nand U1596 (N_1596,N_488,N_192);
nor U1597 (N_1597,N_33,N_362);
or U1598 (N_1598,N_182,N_124);
or U1599 (N_1599,N_628,N_387);
nor U1600 (N_1600,N_811,N_674);
xor U1601 (N_1601,N_747,N_589);
or U1602 (N_1602,N_579,N_950);
nor U1603 (N_1603,N_501,N_752);
xor U1604 (N_1604,N_815,N_382);
nor U1605 (N_1605,N_892,N_119);
and U1606 (N_1606,N_852,N_325);
or U1607 (N_1607,N_988,N_869);
or U1608 (N_1608,N_505,N_792);
nand U1609 (N_1609,N_897,N_873);
nand U1610 (N_1610,N_981,N_14);
nor U1611 (N_1611,N_365,N_274);
and U1612 (N_1612,N_209,N_553);
nand U1613 (N_1613,N_332,N_92);
and U1614 (N_1614,N_613,N_365);
or U1615 (N_1615,N_907,N_375);
or U1616 (N_1616,N_692,N_787);
nor U1617 (N_1617,N_441,N_236);
and U1618 (N_1618,N_456,N_199);
nand U1619 (N_1619,N_383,N_579);
and U1620 (N_1620,N_830,N_421);
xor U1621 (N_1621,N_683,N_604);
or U1622 (N_1622,N_397,N_945);
or U1623 (N_1623,N_954,N_644);
xnor U1624 (N_1624,N_397,N_152);
nor U1625 (N_1625,N_937,N_622);
and U1626 (N_1626,N_563,N_545);
nor U1627 (N_1627,N_721,N_915);
and U1628 (N_1628,N_233,N_234);
nand U1629 (N_1629,N_605,N_156);
or U1630 (N_1630,N_482,N_663);
and U1631 (N_1631,N_91,N_931);
xor U1632 (N_1632,N_947,N_562);
xor U1633 (N_1633,N_427,N_443);
nand U1634 (N_1634,N_737,N_953);
or U1635 (N_1635,N_549,N_160);
xor U1636 (N_1636,N_921,N_68);
and U1637 (N_1637,N_40,N_556);
xnor U1638 (N_1638,N_869,N_302);
or U1639 (N_1639,N_478,N_474);
nand U1640 (N_1640,N_249,N_190);
or U1641 (N_1641,N_958,N_364);
nor U1642 (N_1642,N_373,N_777);
xnor U1643 (N_1643,N_359,N_319);
or U1644 (N_1644,N_410,N_942);
nand U1645 (N_1645,N_70,N_981);
nand U1646 (N_1646,N_178,N_843);
nand U1647 (N_1647,N_81,N_672);
xnor U1648 (N_1648,N_709,N_58);
xnor U1649 (N_1649,N_583,N_840);
xnor U1650 (N_1650,N_598,N_442);
nor U1651 (N_1651,N_499,N_189);
xnor U1652 (N_1652,N_258,N_454);
and U1653 (N_1653,N_974,N_907);
or U1654 (N_1654,N_266,N_394);
or U1655 (N_1655,N_746,N_320);
xnor U1656 (N_1656,N_672,N_865);
nand U1657 (N_1657,N_898,N_665);
nor U1658 (N_1658,N_28,N_373);
or U1659 (N_1659,N_469,N_922);
nand U1660 (N_1660,N_345,N_786);
nor U1661 (N_1661,N_921,N_298);
nor U1662 (N_1662,N_154,N_519);
and U1663 (N_1663,N_295,N_278);
nand U1664 (N_1664,N_679,N_887);
and U1665 (N_1665,N_655,N_251);
or U1666 (N_1666,N_575,N_431);
xor U1667 (N_1667,N_280,N_114);
xor U1668 (N_1668,N_445,N_811);
nor U1669 (N_1669,N_129,N_485);
and U1670 (N_1670,N_198,N_17);
nor U1671 (N_1671,N_252,N_87);
or U1672 (N_1672,N_419,N_698);
nand U1673 (N_1673,N_734,N_54);
nand U1674 (N_1674,N_431,N_367);
nand U1675 (N_1675,N_308,N_916);
nand U1676 (N_1676,N_559,N_534);
nor U1677 (N_1677,N_174,N_908);
xnor U1678 (N_1678,N_656,N_584);
nand U1679 (N_1679,N_521,N_381);
nand U1680 (N_1680,N_713,N_924);
nor U1681 (N_1681,N_423,N_155);
xnor U1682 (N_1682,N_994,N_916);
and U1683 (N_1683,N_916,N_580);
and U1684 (N_1684,N_601,N_953);
nor U1685 (N_1685,N_376,N_873);
and U1686 (N_1686,N_746,N_297);
xor U1687 (N_1687,N_134,N_485);
or U1688 (N_1688,N_924,N_214);
or U1689 (N_1689,N_129,N_160);
xnor U1690 (N_1690,N_876,N_73);
nand U1691 (N_1691,N_129,N_999);
or U1692 (N_1692,N_93,N_293);
xnor U1693 (N_1693,N_891,N_352);
nor U1694 (N_1694,N_357,N_222);
xnor U1695 (N_1695,N_931,N_242);
and U1696 (N_1696,N_297,N_28);
nor U1697 (N_1697,N_696,N_562);
xnor U1698 (N_1698,N_694,N_479);
xor U1699 (N_1699,N_195,N_519);
or U1700 (N_1700,N_661,N_561);
or U1701 (N_1701,N_384,N_122);
nor U1702 (N_1702,N_354,N_727);
nand U1703 (N_1703,N_84,N_836);
nand U1704 (N_1704,N_296,N_564);
or U1705 (N_1705,N_4,N_84);
xnor U1706 (N_1706,N_183,N_978);
xor U1707 (N_1707,N_951,N_298);
xnor U1708 (N_1708,N_753,N_472);
or U1709 (N_1709,N_951,N_764);
or U1710 (N_1710,N_325,N_787);
nor U1711 (N_1711,N_599,N_184);
nand U1712 (N_1712,N_717,N_553);
or U1713 (N_1713,N_53,N_333);
xnor U1714 (N_1714,N_725,N_114);
xnor U1715 (N_1715,N_857,N_587);
or U1716 (N_1716,N_564,N_963);
xnor U1717 (N_1717,N_451,N_591);
nor U1718 (N_1718,N_547,N_98);
nand U1719 (N_1719,N_469,N_276);
nand U1720 (N_1720,N_658,N_953);
nor U1721 (N_1721,N_531,N_733);
or U1722 (N_1722,N_136,N_407);
nand U1723 (N_1723,N_390,N_778);
xor U1724 (N_1724,N_469,N_83);
and U1725 (N_1725,N_453,N_63);
and U1726 (N_1726,N_634,N_352);
or U1727 (N_1727,N_892,N_513);
and U1728 (N_1728,N_384,N_39);
or U1729 (N_1729,N_899,N_907);
nand U1730 (N_1730,N_421,N_222);
and U1731 (N_1731,N_1,N_454);
xor U1732 (N_1732,N_766,N_954);
nand U1733 (N_1733,N_237,N_245);
or U1734 (N_1734,N_456,N_341);
nand U1735 (N_1735,N_227,N_313);
nand U1736 (N_1736,N_447,N_788);
nor U1737 (N_1737,N_704,N_824);
and U1738 (N_1738,N_428,N_790);
nor U1739 (N_1739,N_21,N_649);
or U1740 (N_1740,N_976,N_501);
nand U1741 (N_1741,N_207,N_423);
nor U1742 (N_1742,N_116,N_905);
and U1743 (N_1743,N_613,N_819);
nor U1744 (N_1744,N_167,N_312);
xor U1745 (N_1745,N_615,N_241);
nor U1746 (N_1746,N_562,N_351);
nor U1747 (N_1747,N_35,N_963);
and U1748 (N_1748,N_684,N_396);
nand U1749 (N_1749,N_280,N_868);
or U1750 (N_1750,N_136,N_576);
nor U1751 (N_1751,N_918,N_586);
or U1752 (N_1752,N_848,N_135);
or U1753 (N_1753,N_225,N_56);
nand U1754 (N_1754,N_91,N_522);
nand U1755 (N_1755,N_920,N_248);
and U1756 (N_1756,N_420,N_916);
or U1757 (N_1757,N_545,N_512);
xnor U1758 (N_1758,N_652,N_779);
or U1759 (N_1759,N_946,N_396);
xor U1760 (N_1760,N_222,N_600);
or U1761 (N_1761,N_13,N_815);
nand U1762 (N_1762,N_546,N_751);
and U1763 (N_1763,N_551,N_41);
nor U1764 (N_1764,N_678,N_737);
nand U1765 (N_1765,N_522,N_68);
and U1766 (N_1766,N_629,N_420);
xor U1767 (N_1767,N_858,N_880);
nand U1768 (N_1768,N_408,N_894);
and U1769 (N_1769,N_854,N_858);
nand U1770 (N_1770,N_920,N_798);
xor U1771 (N_1771,N_92,N_383);
and U1772 (N_1772,N_571,N_760);
or U1773 (N_1773,N_303,N_470);
xnor U1774 (N_1774,N_336,N_361);
and U1775 (N_1775,N_716,N_386);
or U1776 (N_1776,N_528,N_938);
and U1777 (N_1777,N_246,N_640);
and U1778 (N_1778,N_401,N_300);
and U1779 (N_1779,N_362,N_848);
and U1780 (N_1780,N_451,N_205);
nand U1781 (N_1781,N_529,N_579);
nand U1782 (N_1782,N_513,N_357);
nand U1783 (N_1783,N_73,N_737);
nor U1784 (N_1784,N_163,N_152);
and U1785 (N_1785,N_579,N_707);
nand U1786 (N_1786,N_127,N_996);
nor U1787 (N_1787,N_111,N_923);
or U1788 (N_1788,N_267,N_478);
nand U1789 (N_1789,N_340,N_831);
or U1790 (N_1790,N_875,N_439);
nor U1791 (N_1791,N_931,N_704);
and U1792 (N_1792,N_966,N_292);
and U1793 (N_1793,N_790,N_206);
and U1794 (N_1794,N_946,N_596);
and U1795 (N_1795,N_695,N_723);
nand U1796 (N_1796,N_539,N_446);
or U1797 (N_1797,N_780,N_570);
nor U1798 (N_1798,N_907,N_15);
nand U1799 (N_1799,N_790,N_150);
nor U1800 (N_1800,N_469,N_54);
nand U1801 (N_1801,N_15,N_792);
or U1802 (N_1802,N_873,N_943);
or U1803 (N_1803,N_141,N_482);
nor U1804 (N_1804,N_621,N_319);
nand U1805 (N_1805,N_149,N_756);
or U1806 (N_1806,N_786,N_443);
nand U1807 (N_1807,N_714,N_393);
nor U1808 (N_1808,N_304,N_318);
and U1809 (N_1809,N_209,N_162);
nand U1810 (N_1810,N_565,N_898);
nor U1811 (N_1811,N_216,N_974);
nor U1812 (N_1812,N_558,N_646);
or U1813 (N_1813,N_95,N_617);
nor U1814 (N_1814,N_826,N_508);
xor U1815 (N_1815,N_262,N_434);
and U1816 (N_1816,N_881,N_738);
or U1817 (N_1817,N_961,N_478);
nor U1818 (N_1818,N_449,N_833);
nand U1819 (N_1819,N_401,N_473);
and U1820 (N_1820,N_333,N_36);
or U1821 (N_1821,N_724,N_925);
nand U1822 (N_1822,N_839,N_760);
nor U1823 (N_1823,N_266,N_138);
nand U1824 (N_1824,N_849,N_254);
nor U1825 (N_1825,N_410,N_788);
nand U1826 (N_1826,N_483,N_212);
or U1827 (N_1827,N_615,N_474);
nand U1828 (N_1828,N_656,N_355);
xor U1829 (N_1829,N_397,N_810);
xor U1830 (N_1830,N_71,N_340);
or U1831 (N_1831,N_953,N_423);
nand U1832 (N_1832,N_657,N_317);
nand U1833 (N_1833,N_631,N_135);
and U1834 (N_1834,N_763,N_341);
or U1835 (N_1835,N_906,N_978);
nor U1836 (N_1836,N_581,N_224);
or U1837 (N_1837,N_23,N_276);
nand U1838 (N_1838,N_394,N_995);
xor U1839 (N_1839,N_115,N_961);
nand U1840 (N_1840,N_203,N_902);
nor U1841 (N_1841,N_550,N_655);
xnor U1842 (N_1842,N_217,N_665);
nor U1843 (N_1843,N_391,N_674);
or U1844 (N_1844,N_22,N_849);
or U1845 (N_1845,N_747,N_184);
or U1846 (N_1846,N_999,N_216);
nor U1847 (N_1847,N_555,N_111);
and U1848 (N_1848,N_66,N_346);
nand U1849 (N_1849,N_355,N_135);
xor U1850 (N_1850,N_927,N_470);
nand U1851 (N_1851,N_871,N_117);
nand U1852 (N_1852,N_449,N_26);
and U1853 (N_1853,N_343,N_683);
nor U1854 (N_1854,N_988,N_35);
nand U1855 (N_1855,N_591,N_376);
xor U1856 (N_1856,N_953,N_732);
xnor U1857 (N_1857,N_646,N_474);
xnor U1858 (N_1858,N_981,N_836);
nor U1859 (N_1859,N_897,N_426);
and U1860 (N_1860,N_479,N_701);
or U1861 (N_1861,N_357,N_392);
nand U1862 (N_1862,N_123,N_916);
and U1863 (N_1863,N_995,N_745);
or U1864 (N_1864,N_585,N_162);
nor U1865 (N_1865,N_361,N_429);
nand U1866 (N_1866,N_990,N_889);
nor U1867 (N_1867,N_725,N_833);
or U1868 (N_1868,N_852,N_508);
xnor U1869 (N_1869,N_59,N_984);
xnor U1870 (N_1870,N_11,N_17);
or U1871 (N_1871,N_177,N_807);
nor U1872 (N_1872,N_89,N_196);
nor U1873 (N_1873,N_909,N_724);
and U1874 (N_1874,N_68,N_817);
nand U1875 (N_1875,N_207,N_858);
and U1876 (N_1876,N_371,N_955);
or U1877 (N_1877,N_554,N_687);
xnor U1878 (N_1878,N_148,N_419);
nand U1879 (N_1879,N_536,N_350);
or U1880 (N_1880,N_402,N_308);
nand U1881 (N_1881,N_359,N_900);
xor U1882 (N_1882,N_243,N_911);
or U1883 (N_1883,N_622,N_599);
nor U1884 (N_1884,N_180,N_373);
and U1885 (N_1885,N_337,N_812);
nand U1886 (N_1886,N_353,N_760);
nand U1887 (N_1887,N_534,N_722);
or U1888 (N_1888,N_520,N_58);
and U1889 (N_1889,N_261,N_649);
nand U1890 (N_1890,N_215,N_316);
nor U1891 (N_1891,N_693,N_642);
xor U1892 (N_1892,N_752,N_226);
nor U1893 (N_1893,N_532,N_185);
nor U1894 (N_1894,N_684,N_200);
nand U1895 (N_1895,N_581,N_96);
xnor U1896 (N_1896,N_946,N_731);
xnor U1897 (N_1897,N_160,N_104);
nor U1898 (N_1898,N_66,N_93);
and U1899 (N_1899,N_426,N_319);
nand U1900 (N_1900,N_381,N_632);
xnor U1901 (N_1901,N_983,N_596);
nand U1902 (N_1902,N_553,N_92);
or U1903 (N_1903,N_181,N_78);
nand U1904 (N_1904,N_10,N_796);
nand U1905 (N_1905,N_378,N_621);
xnor U1906 (N_1906,N_779,N_684);
nand U1907 (N_1907,N_208,N_482);
or U1908 (N_1908,N_142,N_647);
or U1909 (N_1909,N_155,N_733);
xor U1910 (N_1910,N_368,N_819);
or U1911 (N_1911,N_475,N_384);
xnor U1912 (N_1912,N_435,N_572);
nand U1913 (N_1913,N_502,N_210);
or U1914 (N_1914,N_822,N_107);
nor U1915 (N_1915,N_614,N_231);
nor U1916 (N_1916,N_303,N_608);
or U1917 (N_1917,N_389,N_729);
nand U1918 (N_1918,N_188,N_960);
or U1919 (N_1919,N_876,N_357);
and U1920 (N_1920,N_320,N_691);
xor U1921 (N_1921,N_238,N_281);
and U1922 (N_1922,N_640,N_42);
nand U1923 (N_1923,N_941,N_106);
nor U1924 (N_1924,N_38,N_462);
or U1925 (N_1925,N_275,N_66);
xor U1926 (N_1926,N_26,N_366);
nor U1927 (N_1927,N_416,N_314);
nor U1928 (N_1928,N_581,N_903);
or U1929 (N_1929,N_928,N_302);
nor U1930 (N_1930,N_876,N_533);
nand U1931 (N_1931,N_481,N_342);
or U1932 (N_1932,N_660,N_491);
and U1933 (N_1933,N_929,N_24);
or U1934 (N_1934,N_776,N_571);
or U1935 (N_1935,N_166,N_246);
nor U1936 (N_1936,N_33,N_898);
and U1937 (N_1937,N_941,N_856);
and U1938 (N_1938,N_748,N_934);
nor U1939 (N_1939,N_737,N_890);
nand U1940 (N_1940,N_918,N_510);
xor U1941 (N_1941,N_902,N_816);
or U1942 (N_1942,N_482,N_780);
and U1943 (N_1943,N_545,N_89);
nand U1944 (N_1944,N_132,N_978);
or U1945 (N_1945,N_936,N_100);
or U1946 (N_1946,N_412,N_322);
and U1947 (N_1947,N_82,N_876);
or U1948 (N_1948,N_7,N_787);
nand U1949 (N_1949,N_394,N_233);
xnor U1950 (N_1950,N_76,N_854);
xnor U1951 (N_1951,N_17,N_389);
and U1952 (N_1952,N_255,N_831);
xor U1953 (N_1953,N_795,N_192);
nor U1954 (N_1954,N_442,N_44);
or U1955 (N_1955,N_944,N_307);
and U1956 (N_1956,N_749,N_837);
nor U1957 (N_1957,N_505,N_778);
nand U1958 (N_1958,N_384,N_235);
or U1959 (N_1959,N_875,N_942);
nor U1960 (N_1960,N_982,N_818);
and U1961 (N_1961,N_493,N_79);
and U1962 (N_1962,N_584,N_670);
and U1963 (N_1963,N_210,N_372);
or U1964 (N_1964,N_303,N_639);
nand U1965 (N_1965,N_777,N_710);
nor U1966 (N_1966,N_597,N_976);
xor U1967 (N_1967,N_836,N_640);
or U1968 (N_1968,N_352,N_954);
and U1969 (N_1969,N_562,N_500);
and U1970 (N_1970,N_577,N_736);
xnor U1971 (N_1971,N_295,N_873);
and U1972 (N_1972,N_453,N_846);
or U1973 (N_1973,N_242,N_401);
nor U1974 (N_1974,N_217,N_931);
nor U1975 (N_1975,N_457,N_246);
or U1976 (N_1976,N_332,N_792);
nand U1977 (N_1977,N_891,N_184);
nand U1978 (N_1978,N_269,N_288);
xor U1979 (N_1979,N_219,N_46);
xor U1980 (N_1980,N_715,N_878);
nand U1981 (N_1981,N_555,N_129);
and U1982 (N_1982,N_425,N_82);
xnor U1983 (N_1983,N_289,N_338);
nand U1984 (N_1984,N_288,N_308);
xnor U1985 (N_1985,N_388,N_309);
xnor U1986 (N_1986,N_410,N_511);
nand U1987 (N_1987,N_354,N_529);
nor U1988 (N_1988,N_848,N_235);
and U1989 (N_1989,N_480,N_947);
nor U1990 (N_1990,N_11,N_985);
or U1991 (N_1991,N_792,N_67);
nor U1992 (N_1992,N_276,N_892);
nand U1993 (N_1993,N_172,N_443);
nor U1994 (N_1994,N_284,N_226);
and U1995 (N_1995,N_213,N_818);
or U1996 (N_1996,N_890,N_577);
nor U1997 (N_1997,N_650,N_949);
or U1998 (N_1998,N_939,N_900);
or U1999 (N_1999,N_617,N_693);
nand U2000 (N_2000,N_1608,N_1383);
nor U2001 (N_2001,N_1355,N_1899);
or U2002 (N_2002,N_1915,N_1120);
xnor U2003 (N_2003,N_1087,N_1560);
and U2004 (N_2004,N_1512,N_1907);
xnor U2005 (N_2005,N_1689,N_1146);
nand U2006 (N_2006,N_1211,N_1766);
xor U2007 (N_2007,N_1350,N_1949);
nor U2008 (N_2008,N_1836,N_1820);
and U2009 (N_2009,N_1500,N_1777);
xnor U2010 (N_2010,N_1156,N_1534);
nor U2011 (N_2011,N_1171,N_1433);
nor U2012 (N_2012,N_1053,N_1154);
nor U2013 (N_2013,N_1417,N_1672);
nand U2014 (N_2014,N_1405,N_1660);
nor U2015 (N_2015,N_1056,N_1546);
nand U2016 (N_2016,N_1853,N_1765);
nand U2017 (N_2017,N_1070,N_1467);
xnor U2018 (N_2018,N_1522,N_1014);
or U2019 (N_2019,N_1860,N_1451);
xor U2020 (N_2020,N_1513,N_1113);
nand U2021 (N_2021,N_1695,N_1835);
or U2022 (N_2022,N_1391,N_1166);
nand U2023 (N_2023,N_1091,N_1665);
or U2024 (N_2024,N_1484,N_1948);
xnor U2025 (N_2025,N_1128,N_1914);
nor U2026 (N_2026,N_1668,N_1478);
or U2027 (N_2027,N_1844,N_1790);
nand U2028 (N_2028,N_1325,N_1928);
or U2029 (N_2029,N_1531,N_1293);
or U2030 (N_2030,N_1228,N_1382);
nand U2031 (N_2031,N_1252,N_1047);
nor U2032 (N_2032,N_1872,N_1328);
or U2033 (N_2033,N_1038,N_1498);
nor U2034 (N_2034,N_1728,N_1549);
and U2035 (N_2035,N_1842,N_1739);
nor U2036 (N_2036,N_1438,N_1487);
and U2037 (N_2037,N_1023,N_1138);
and U2038 (N_2038,N_1753,N_1002);
xnor U2039 (N_2039,N_1155,N_1468);
xor U2040 (N_2040,N_1351,N_1840);
or U2041 (N_2041,N_1197,N_1568);
nand U2042 (N_2042,N_1745,N_1116);
or U2043 (N_2043,N_1241,N_1266);
nor U2044 (N_2044,N_1910,N_1401);
nor U2045 (N_2045,N_1551,N_1400);
and U2046 (N_2046,N_1804,N_1664);
or U2047 (N_2047,N_1800,N_1571);
or U2048 (N_2048,N_1951,N_1063);
and U2049 (N_2049,N_1707,N_1989);
nand U2050 (N_2050,N_1258,N_1598);
or U2051 (N_2051,N_1843,N_1801);
or U2052 (N_2052,N_1286,N_1912);
xor U2053 (N_2053,N_1191,N_1494);
xor U2054 (N_2054,N_1363,N_1524);
xnor U2055 (N_2055,N_1260,N_1505);
xor U2056 (N_2056,N_1388,N_1812);
xor U2057 (N_2057,N_1666,N_1802);
nor U2058 (N_2058,N_1845,N_1719);
nand U2059 (N_2059,N_1394,N_1082);
and U2060 (N_2060,N_1327,N_1413);
nor U2061 (N_2061,N_1003,N_1779);
or U2062 (N_2062,N_1673,N_1204);
and U2063 (N_2063,N_1480,N_1538);
nor U2064 (N_2064,N_1396,N_1490);
and U2065 (N_2065,N_1376,N_1445);
nor U2066 (N_2066,N_1593,N_1220);
or U2067 (N_2067,N_1065,N_1318);
nand U2068 (N_2068,N_1297,N_1878);
nand U2069 (N_2069,N_1752,N_1595);
or U2070 (N_2070,N_1127,N_1424);
and U2071 (N_2071,N_1261,N_1435);
nor U2072 (N_2072,N_1074,N_1353);
nor U2073 (N_2073,N_1580,N_1039);
or U2074 (N_2074,N_1570,N_1028);
or U2075 (N_2075,N_1964,N_1436);
nand U2076 (N_2076,N_1557,N_1681);
or U2077 (N_2077,N_1939,N_1723);
or U2078 (N_2078,N_1221,N_1886);
xnor U2079 (N_2079,N_1345,N_1900);
and U2080 (N_2080,N_1320,N_1309);
nand U2081 (N_2081,N_1817,N_1540);
and U2082 (N_2082,N_1868,N_1193);
nand U2083 (N_2083,N_1958,N_1810);
and U2084 (N_2084,N_1930,N_1234);
or U2085 (N_2085,N_1602,N_1970);
nand U2086 (N_2086,N_1257,N_1620);
nor U2087 (N_2087,N_1049,N_1052);
xnor U2088 (N_2088,N_1877,N_1903);
nor U2089 (N_2089,N_1893,N_1225);
or U2090 (N_2090,N_1447,N_1663);
nand U2091 (N_2091,N_1541,N_1306);
and U2092 (N_2092,N_1690,N_1461);
and U2093 (N_2093,N_1167,N_1215);
or U2094 (N_2094,N_1352,N_1576);
nand U2095 (N_2095,N_1996,N_1890);
or U2096 (N_2096,N_1050,N_1129);
and U2097 (N_2097,N_1760,N_1302);
or U2098 (N_2098,N_1624,N_1709);
or U2099 (N_2099,N_1343,N_1040);
xnor U2100 (N_2100,N_1605,N_1873);
nand U2101 (N_2101,N_1937,N_1575);
and U2102 (N_2102,N_1239,N_1969);
nor U2103 (N_2103,N_1294,N_1313);
nor U2104 (N_2104,N_1710,N_1251);
nand U2105 (N_2105,N_1264,N_1150);
nor U2106 (N_2106,N_1242,N_1863);
nor U2107 (N_2107,N_1096,N_1621);
nor U2108 (N_2108,N_1532,N_1094);
xor U2109 (N_2109,N_1832,N_1420);
xnor U2110 (N_2110,N_1861,N_1960);
xor U2111 (N_2111,N_1566,N_1644);
or U2112 (N_2112,N_1004,N_1975);
nand U2113 (N_2113,N_1418,N_1961);
and U2114 (N_2114,N_1983,N_1013);
or U2115 (N_2115,N_1229,N_1462);
nand U2116 (N_2116,N_1616,N_1392);
or U2117 (N_2117,N_1591,N_1677);
xnor U2118 (N_2118,N_1667,N_1332);
xnor U2119 (N_2119,N_1730,N_1651);
nand U2120 (N_2120,N_1527,N_1785);
xor U2121 (N_2121,N_1315,N_1354);
nand U2122 (N_2122,N_1153,N_1543);
nand U2123 (N_2123,N_1963,N_1411);
or U2124 (N_2124,N_1083,N_1629);
nand U2125 (N_2125,N_1323,N_1387);
nor U2126 (N_2126,N_1278,N_1465);
xor U2127 (N_2127,N_1680,N_1669);
or U2128 (N_2128,N_1579,N_1972);
xnor U2129 (N_2129,N_1539,N_1290);
nor U2130 (N_2130,N_1713,N_1272);
or U2131 (N_2131,N_1104,N_1578);
and U2132 (N_2132,N_1636,N_1122);
or U2133 (N_2133,N_1992,N_1279);
or U2134 (N_2134,N_1881,N_1995);
nand U2135 (N_2135,N_1043,N_1255);
nand U2136 (N_2136,N_1604,N_1235);
nor U2137 (N_2137,N_1654,N_1131);
xnor U2138 (N_2138,N_1699,N_1757);
and U2139 (N_2139,N_1712,N_1750);
nand U2140 (N_2140,N_1559,N_1922);
or U2141 (N_2141,N_1112,N_1725);
or U2142 (N_2142,N_1657,N_1022);
and U2143 (N_2143,N_1941,N_1045);
and U2144 (N_2144,N_1170,N_1476);
and U2145 (N_2145,N_1909,N_1419);
nand U2146 (N_2146,N_1208,N_1178);
or U2147 (N_2147,N_1175,N_1249);
or U2148 (N_2148,N_1796,N_1068);
xor U2149 (N_2149,N_1622,N_1100);
nand U2150 (N_2150,N_1600,N_1942);
nand U2151 (N_2151,N_1870,N_1823);
nand U2152 (N_2152,N_1130,N_1032);
xnor U2153 (N_2153,N_1316,N_1997);
nor U2154 (N_2154,N_1289,N_1837);
xor U2155 (N_2155,N_1784,N_1535);
nand U2156 (N_2156,N_1805,N_1212);
or U2157 (N_2157,N_1923,N_1731);
nand U2158 (N_2158,N_1188,N_1301);
xnor U2159 (N_2159,N_1062,N_1377);
nand U2160 (N_2160,N_1361,N_1517);
or U2161 (N_2161,N_1523,N_1691);
and U2162 (N_2162,N_1510,N_1986);
and U2163 (N_2163,N_1459,N_1847);
nand U2164 (N_2164,N_1727,N_1917);
xnor U2165 (N_2165,N_1601,N_1846);
and U2166 (N_2166,N_1230,N_1545);
and U2167 (N_2167,N_1299,N_1107);
nand U2168 (N_2168,N_1428,N_1213);
xor U2169 (N_2169,N_1288,N_1764);
xor U2170 (N_2170,N_1019,N_1256);
xnor U2171 (N_2171,N_1051,N_1612);
nand U2172 (N_2172,N_1555,N_1947);
nand U2173 (N_2173,N_1184,N_1123);
and U2174 (N_2174,N_1811,N_1422);
or U2175 (N_2175,N_1645,N_1618);
or U2176 (N_2176,N_1953,N_1493);
xnor U2177 (N_2177,N_1714,N_1359);
or U2178 (N_2178,N_1702,N_1862);
or U2179 (N_2179,N_1203,N_1009);
and U2180 (N_2180,N_1838,N_1815);
nor U2181 (N_2181,N_1375,N_1913);
xnor U2182 (N_2182,N_1277,N_1464);
nor U2183 (N_2183,N_1304,N_1058);
or U2184 (N_2184,N_1086,N_1895);
nand U2185 (N_2185,N_1275,N_1207);
nand U2186 (N_2186,N_1305,N_1483);
nor U2187 (N_2187,N_1037,N_1874);
or U2188 (N_2188,N_1652,N_1147);
and U2189 (N_2189,N_1768,N_1084);
and U2190 (N_2190,N_1630,N_1296);
xnor U2191 (N_2191,N_1974,N_1973);
nor U2192 (N_2192,N_1233,N_1427);
or U2193 (N_2193,N_1341,N_1735);
and U2194 (N_2194,N_1029,N_1158);
and U2195 (N_2195,N_1945,N_1816);
xor U2196 (N_2196,N_1477,N_1456);
nor U2197 (N_2197,N_1268,N_1044);
nor U2198 (N_2198,N_1430,N_1581);
nor U2199 (N_2199,N_1916,N_1446);
or U2200 (N_2200,N_1993,N_1773);
nor U2201 (N_2201,N_1888,N_1499);
and U2202 (N_2202,N_1340,N_1504);
nand U2203 (N_2203,N_1181,N_1530);
xor U2204 (N_2204,N_1988,N_1190);
and U2205 (N_2205,N_1747,N_1001);
and U2206 (N_2206,N_1187,N_1693);
nand U2207 (N_2207,N_1911,N_1717);
and U2208 (N_2208,N_1000,N_1834);
xor U2209 (N_2209,N_1108,N_1423);
or U2210 (N_2210,N_1807,N_1679);
nor U2211 (N_2211,N_1139,N_1390);
or U2212 (N_2212,N_1414,N_1650);
nand U2213 (N_2213,N_1470,N_1011);
nand U2214 (N_2214,N_1236,N_1226);
nand U2215 (N_2215,N_1788,N_1245);
nor U2216 (N_2216,N_1936,N_1463);
xor U2217 (N_2217,N_1199,N_1615);
or U2218 (N_2218,N_1926,N_1080);
nand U2219 (N_2219,N_1059,N_1143);
nand U2220 (N_2220,N_1851,N_1751);
nand U2221 (N_2221,N_1173,N_1165);
nor U2222 (N_2222,N_1440,N_1659);
xnor U2223 (N_2223,N_1298,N_1865);
or U2224 (N_2224,N_1253,N_1339);
xor U2225 (N_2225,N_1018,N_1168);
nor U2226 (N_2226,N_1761,N_1572);
nand U2227 (N_2227,N_1101,N_1415);
nand U2228 (N_2228,N_1584,N_1871);
nor U2229 (N_2229,N_1283,N_1932);
and U2230 (N_2230,N_1473,N_1908);
nand U2231 (N_2231,N_1491,N_1329);
and U2232 (N_2232,N_1088,N_1267);
or U2233 (N_2233,N_1090,N_1262);
nand U2234 (N_2234,N_1831,N_1824);
nand U2235 (N_2235,N_1778,N_1406);
nor U2236 (N_2236,N_1330,N_1854);
and U2237 (N_2237,N_1946,N_1347);
nor U2238 (N_2238,N_1696,N_1643);
or U2239 (N_2239,N_1326,N_1250);
nand U2240 (N_2240,N_1894,N_1386);
nand U2241 (N_2241,N_1133,N_1148);
xnor U2242 (N_2242,N_1061,N_1829);
and U2243 (N_2243,N_1639,N_1182);
or U2244 (N_2244,N_1076,N_1554);
or U2245 (N_2245,N_1337,N_1295);
or U2246 (N_2246,N_1736,N_1426);
or U2247 (N_2247,N_1030,N_1869);
nor U2248 (N_2248,N_1592,N_1688);
xor U2249 (N_2249,N_1136,N_1626);
and U2250 (N_2250,N_1176,N_1515);
or U2251 (N_2251,N_1164,N_1991);
xor U2252 (N_2252,N_1378,N_1635);
and U2253 (N_2253,N_1486,N_1925);
and U2254 (N_2254,N_1927,N_1850);
or U2255 (N_2255,N_1611,N_1111);
or U2256 (N_2256,N_1799,N_1317);
nand U2257 (N_2257,N_1981,N_1619);
and U2258 (N_2258,N_1222,N_1533);
or U2259 (N_2259,N_1075,N_1403);
xnor U2260 (N_2260,N_1548,N_1021);
xor U2261 (N_2261,N_1733,N_1274);
xnor U2262 (N_2262,N_1209,N_1310);
nor U2263 (N_2263,N_1887,N_1469);
xnor U2264 (N_2264,N_1159,N_1806);
xor U2265 (N_2265,N_1743,N_1357);
or U2266 (N_2266,N_1360,N_1008);
and U2267 (N_2267,N_1526,N_1471);
xor U2268 (N_2268,N_1185,N_1244);
xnor U2269 (N_2269,N_1569,N_1511);
nand U2270 (N_2270,N_1152,N_1919);
or U2271 (N_2271,N_1017,N_1587);
or U2272 (N_2272,N_1749,N_1334);
nand U2273 (N_2273,N_1640,N_1726);
xor U2274 (N_2274,N_1085,N_1588);
and U2275 (N_2275,N_1827,N_1333);
nand U2276 (N_2276,N_1786,N_1756);
nor U2277 (N_2277,N_1976,N_1161);
nor U2278 (N_2278,N_1819,N_1867);
nand U2279 (N_2279,N_1603,N_1586);
or U2280 (N_2280,N_1782,N_1738);
xor U2281 (N_2281,N_1662,N_1453);
xnor U2282 (N_2282,N_1706,N_1367);
nand U2283 (N_2283,N_1631,N_1567);
nor U2284 (N_2284,N_1118,N_1194);
nor U2285 (N_2285,N_1454,N_1125);
nor U2286 (N_2286,N_1771,N_1322);
or U2287 (N_2287,N_1905,N_1787);
and U2288 (N_2288,N_1006,N_1921);
and U2289 (N_2289,N_1271,N_1195);
xor U2290 (N_2290,N_1321,N_1553);
and U2291 (N_2291,N_1521,N_1449);
and U2292 (N_2292,N_1319,N_1781);
nand U2293 (N_2293,N_1982,N_1384);
nor U2294 (N_2294,N_1506,N_1623);
and U2295 (N_2295,N_1825,N_1685);
nand U2296 (N_2296,N_1774,N_1783);
or U2297 (N_2297,N_1791,N_1966);
or U2298 (N_2298,N_1589,N_1336);
nor U2299 (N_2299,N_1550,N_1859);
nor U2300 (N_2300,N_1495,N_1189);
xor U2301 (N_2301,N_1617,N_1206);
or U2302 (N_2302,N_1775,N_1081);
or U2303 (N_2303,N_1496,N_1016);
or U2304 (N_2304,N_1770,N_1520);
nor U2305 (N_2305,N_1931,N_1795);
nor U2306 (N_2306,N_1421,N_1965);
nor U2307 (N_2307,N_1186,N_1458);
and U2308 (N_2308,N_1882,N_1431);
xor U2309 (N_2309,N_1759,N_1649);
or U2310 (N_2310,N_1280,N_1231);
nor U2311 (N_2311,N_1169,N_1448);
or U2312 (N_2312,N_1897,N_1722);
and U2313 (N_2313,N_1134,N_1744);
xor U2314 (N_2314,N_1552,N_1254);
nand U2315 (N_2315,N_1507,N_1303);
and U2316 (N_2316,N_1105,N_1482);
xor U2317 (N_2317,N_1174,N_1026);
or U2318 (N_2318,N_1682,N_1078);
and U2319 (N_2319,N_1944,N_1833);
or U2320 (N_2320,N_1647,N_1940);
nand U2321 (N_2321,N_1072,N_1346);
and U2322 (N_2322,N_1007,N_1977);
or U2323 (N_2323,N_1704,N_1711);
or U2324 (N_2324,N_1055,N_1140);
xor U2325 (N_2325,N_1410,N_1848);
and U2326 (N_2326,N_1599,N_1701);
nor U2327 (N_2327,N_1219,N_1938);
nand U2328 (N_2328,N_1518,N_1514);
nand U2329 (N_2329,N_1889,N_1641);
and U2330 (N_2330,N_1634,N_1042);
or U2331 (N_2331,N_1412,N_1232);
or U2332 (N_2332,N_1324,N_1822);
xor U2333 (N_2333,N_1489,N_1281);
nand U2334 (N_2334,N_1998,N_1661);
nor U2335 (N_2335,N_1980,N_1089);
nand U2336 (N_2336,N_1920,N_1607);
and U2337 (N_2337,N_1025,N_1124);
nand U2338 (N_2338,N_1071,N_1852);
or U2339 (N_2339,N_1067,N_1767);
nand U2340 (N_2340,N_1876,N_1223);
or U2341 (N_2341,N_1385,N_1671);
nor U2342 (N_2342,N_1374,N_1734);
nor U2343 (N_2343,N_1935,N_1857);
xnor U2344 (N_2344,N_1999,N_1240);
or U2345 (N_2345,N_1676,N_1425);
xor U2346 (N_2346,N_1609,N_1183);
nand U2347 (N_2347,N_1192,N_1117);
nor U2348 (N_2348,N_1460,N_1814);
nand U2349 (N_2349,N_1179,N_1808);
and U2350 (N_2350,N_1632,N_1457);
or U2351 (N_2351,N_1162,N_1628);
xor U2352 (N_2352,N_1046,N_1481);
nor U2353 (N_2353,N_1762,N_1344);
and U2354 (N_2354,N_1763,N_1012);
or U2355 (N_2355,N_1959,N_1311);
nand U2356 (N_2356,N_1536,N_1472);
nand U2357 (N_2357,N_1144,N_1248);
or U2358 (N_2358,N_1439,N_1102);
nor U2359 (N_2359,N_1633,N_1441);
nand U2360 (N_2360,N_1389,N_1674);
nand U2361 (N_2361,N_1813,N_1892);
xnor U2362 (N_2362,N_1364,N_1141);
or U2363 (N_2363,N_1409,N_1338);
and U2364 (N_2364,N_1542,N_1048);
xnor U2365 (N_2365,N_1729,N_1115);
nor U2366 (N_2366,N_1700,N_1529);
nand U2367 (N_2367,N_1793,N_1402);
nand U2368 (N_2368,N_1160,N_1379);
nand U2369 (N_2369,N_1263,N_1349);
and U2370 (N_2370,N_1821,N_1285);
or U2371 (N_2371,N_1740,N_1404);
and U2372 (N_2372,N_1748,N_1196);
nand U2373 (N_2373,N_1918,N_1797);
and U2374 (N_2374,N_1891,N_1794);
and U2375 (N_2375,N_1577,N_1606);
nand U2376 (N_2376,N_1742,N_1841);
nand U2377 (N_2377,N_1830,N_1408);
xnor U2378 (N_2378,N_1119,N_1904);
or U2379 (N_2379,N_1054,N_1955);
nor U2380 (N_2380,N_1202,N_1528);
nand U2381 (N_2381,N_1432,N_1269);
xor U2382 (N_2382,N_1137,N_1561);
nand U2383 (N_2383,N_1502,N_1180);
and U2384 (N_2384,N_1563,N_1474);
or U2385 (N_2385,N_1097,N_1151);
and U2386 (N_2386,N_1715,N_1670);
and U2387 (N_2387,N_1314,N_1492);
and U2388 (N_2388,N_1142,N_1653);
or U2389 (N_2389,N_1519,N_1292);
xor U2390 (N_2390,N_1866,N_1933);
and U2391 (N_2391,N_1901,N_1466);
nor U2392 (N_2392,N_1198,N_1638);
and U2393 (N_2393,N_1686,N_1721);
or U2394 (N_2394,N_1564,N_1342);
nand U2395 (N_2395,N_1683,N_1826);
nand U2396 (N_2396,N_1596,N_1434);
or U2397 (N_2397,N_1849,N_1985);
xnor U2398 (N_2398,N_1246,N_1380);
or U2399 (N_2399,N_1858,N_1655);
and U2400 (N_2400,N_1365,N_1307);
nand U2401 (N_2401,N_1362,N_1809);
xnor U2402 (N_2402,N_1537,N_1373);
and U2403 (N_2403,N_1718,N_1979);
nor U2404 (N_2404,N_1218,N_1145);
xor U2405 (N_2405,N_1746,N_1109);
nor U2406 (N_2406,N_1443,N_1590);
or U2407 (N_2407,N_1395,N_1792);
and U2408 (N_2408,N_1776,N_1348);
or U2409 (N_2409,N_1429,N_1994);
xor U2410 (N_2410,N_1312,N_1381);
nor U2411 (N_2411,N_1210,N_1034);
nor U2412 (N_2412,N_1934,N_1335);
xor U2413 (N_2413,N_1929,N_1488);
nor U2414 (N_2414,N_1358,N_1839);
or U2415 (N_2415,N_1273,N_1027);
nand U2416 (N_2416,N_1902,N_1444);
nor U2417 (N_2417,N_1393,N_1227);
or U2418 (N_2418,N_1163,N_1287);
and U2419 (N_2419,N_1216,N_1031);
and U2420 (N_2420,N_1452,N_1508);
or U2421 (N_2421,N_1177,N_1224);
nand U2422 (N_2422,N_1789,N_1132);
nand U2423 (N_2423,N_1399,N_1201);
nor U2424 (N_2424,N_1978,N_1967);
nor U2425 (N_2425,N_1583,N_1990);
or U2426 (N_2426,N_1556,N_1366);
xnor U2427 (N_2427,N_1300,N_1954);
nor U2428 (N_2428,N_1724,N_1237);
and U2429 (N_2429,N_1121,N_1574);
nor U2430 (N_2430,N_1407,N_1648);
nor U2431 (N_2431,N_1597,N_1703);
or U2432 (N_2432,N_1036,N_1885);
and U2433 (N_2433,N_1708,N_1755);
nand U2434 (N_2434,N_1883,N_1656);
nand U2435 (N_2435,N_1884,N_1758);
and U2436 (N_2436,N_1547,N_1398);
xnor U2437 (N_2437,N_1135,N_1372);
nor U2438 (N_2438,N_1525,N_1020);
or U2439 (N_2439,N_1015,N_1694);
xor U2440 (N_2440,N_1060,N_1875);
and U2441 (N_2441,N_1093,N_1247);
xor U2442 (N_2442,N_1437,N_1754);
xor U2443 (N_2443,N_1033,N_1968);
nor U2444 (N_2444,N_1041,N_1172);
and U2445 (N_2445,N_1818,N_1698);
nor U2446 (N_2446,N_1217,N_1095);
and U2447 (N_2447,N_1906,N_1716);
or U2448 (N_2448,N_1069,N_1610);
and U2449 (N_2449,N_1126,N_1585);
nor U2450 (N_2450,N_1772,N_1331);
nor U2451 (N_2451,N_1956,N_1501);
nor U2452 (N_2452,N_1642,N_1625);
nor U2453 (N_2453,N_1503,N_1855);
or U2454 (N_2454,N_1957,N_1024);
xnor U2455 (N_2455,N_1106,N_1950);
and U2456 (N_2456,N_1684,N_1971);
and U2457 (N_2457,N_1614,N_1594);
xor U2458 (N_2458,N_1064,N_1276);
xnor U2459 (N_2459,N_1798,N_1803);
or U2460 (N_2460,N_1485,N_1416);
nor U2461 (N_2461,N_1544,N_1697);
nor U2462 (N_2462,N_1962,N_1705);
and U2463 (N_2463,N_1562,N_1450);
xnor U2464 (N_2464,N_1265,N_1369);
and U2465 (N_2465,N_1509,N_1479);
nand U2466 (N_2466,N_1259,N_1356);
and U2467 (N_2467,N_1157,N_1720);
and U2468 (N_2468,N_1200,N_1687);
nand U2469 (N_2469,N_1678,N_1114);
xor U2470 (N_2470,N_1952,N_1582);
nand U2471 (N_2471,N_1573,N_1455);
and U2472 (N_2472,N_1658,N_1737);
or U2473 (N_2473,N_1497,N_1284);
and U2474 (N_2474,N_1864,N_1646);
and U2475 (N_2475,N_1092,N_1098);
xnor U2476 (N_2476,N_1516,N_1984);
xor U2477 (N_2477,N_1924,N_1099);
xor U2478 (N_2478,N_1370,N_1565);
nand U2479 (N_2479,N_1282,N_1243);
nor U2480 (N_2480,N_1397,N_1073);
nand U2481 (N_2481,N_1010,N_1879);
nor U2482 (N_2482,N_1627,N_1943);
nor U2483 (N_2483,N_1308,N_1692);
and U2484 (N_2484,N_1035,N_1442);
nor U2485 (N_2485,N_1371,N_1675);
or U2486 (N_2486,N_1880,N_1270);
or U2487 (N_2487,N_1110,N_1214);
and U2488 (N_2488,N_1103,N_1005);
and U2489 (N_2489,N_1637,N_1475);
and U2490 (N_2490,N_1769,N_1741);
and U2491 (N_2491,N_1368,N_1828);
nand U2492 (N_2492,N_1856,N_1896);
and U2493 (N_2493,N_1898,N_1238);
nor U2494 (N_2494,N_1613,N_1079);
and U2495 (N_2495,N_1558,N_1149);
and U2496 (N_2496,N_1780,N_1066);
xor U2497 (N_2497,N_1057,N_1291);
nand U2498 (N_2498,N_1077,N_1987);
nor U2499 (N_2499,N_1205,N_1732);
nand U2500 (N_2500,N_1497,N_1536);
nor U2501 (N_2501,N_1208,N_1531);
or U2502 (N_2502,N_1441,N_1446);
nand U2503 (N_2503,N_1078,N_1673);
xor U2504 (N_2504,N_1192,N_1677);
or U2505 (N_2505,N_1388,N_1694);
nor U2506 (N_2506,N_1256,N_1598);
xor U2507 (N_2507,N_1564,N_1749);
nor U2508 (N_2508,N_1894,N_1257);
xnor U2509 (N_2509,N_1709,N_1619);
xnor U2510 (N_2510,N_1157,N_1764);
nor U2511 (N_2511,N_1432,N_1947);
nand U2512 (N_2512,N_1315,N_1963);
and U2513 (N_2513,N_1847,N_1652);
nor U2514 (N_2514,N_1822,N_1848);
and U2515 (N_2515,N_1021,N_1248);
and U2516 (N_2516,N_1320,N_1803);
nor U2517 (N_2517,N_1142,N_1723);
nand U2518 (N_2518,N_1427,N_1886);
nor U2519 (N_2519,N_1709,N_1304);
nor U2520 (N_2520,N_1393,N_1020);
nand U2521 (N_2521,N_1489,N_1444);
or U2522 (N_2522,N_1484,N_1048);
nand U2523 (N_2523,N_1608,N_1832);
and U2524 (N_2524,N_1736,N_1514);
nor U2525 (N_2525,N_1524,N_1572);
and U2526 (N_2526,N_1688,N_1961);
and U2527 (N_2527,N_1201,N_1485);
xnor U2528 (N_2528,N_1582,N_1470);
or U2529 (N_2529,N_1175,N_1185);
nor U2530 (N_2530,N_1971,N_1989);
xnor U2531 (N_2531,N_1418,N_1597);
or U2532 (N_2532,N_1416,N_1183);
and U2533 (N_2533,N_1770,N_1550);
and U2534 (N_2534,N_1961,N_1592);
nand U2535 (N_2535,N_1199,N_1815);
and U2536 (N_2536,N_1407,N_1072);
nand U2537 (N_2537,N_1857,N_1129);
nand U2538 (N_2538,N_1611,N_1644);
nand U2539 (N_2539,N_1807,N_1924);
and U2540 (N_2540,N_1676,N_1886);
nor U2541 (N_2541,N_1519,N_1542);
and U2542 (N_2542,N_1870,N_1189);
and U2543 (N_2543,N_1062,N_1407);
or U2544 (N_2544,N_1185,N_1984);
nor U2545 (N_2545,N_1896,N_1940);
nor U2546 (N_2546,N_1360,N_1721);
and U2547 (N_2547,N_1113,N_1190);
and U2548 (N_2548,N_1956,N_1265);
nand U2549 (N_2549,N_1751,N_1635);
nor U2550 (N_2550,N_1438,N_1536);
xnor U2551 (N_2551,N_1117,N_1381);
and U2552 (N_2552,N_1100,N_1413);
nand U2553 (N_2553,N_1506,N_1988);
and U2554 (N_2554,N_1481,N_1269);
nor U2555 (N_2555,N_1119,N_1726);
xor U2556 (N_2556,N_1695,N_1919);
xor U2557 (N_2557,N_1335,N_1056);
xnor U2558 (N_2558,N_1647,N_1330);
nand U2559 (N_2559,N_1629,N_1135);
or U2560 (N_2560,N_1495,N_1048);
and U2561 (N_2561,N_1749,N_1415);
and U2562 (N_2562,N_1863,N_1667);
and U2563 (N_2563,N_1904,N_1525);
nor U2564 (N_2564,N_1289,N_1729);
nor U2565 (N_2565,N_1544,N_1518);
xnor U2566 (N_2566,N_1253,N_1239);
xnor U2567 (N_2567,N_1908,N_1370);
and U2568 (N_2568,N_1206,N_1845);
nand U2569 (N_2569,N_1054,N_1563);
xor U2570 (N_2570,N_1835,N_1794);
and U2571 (N_2571,N_1921,N_1314);
xor U2572 (N_2572,N_1171,N_1387);
or U2573 (N_2573,N_1769,N_1114);
nand U2574 (N_2574,N_1790,N_1106);
xor U2575 (N_2575,N_1168,N_1306);
and U2576 (N_2576,N_1850,N_1054);
and U2577 (N_2577,N_1955,N_1941);
nand U2578 (N_2578,N_1647,N_1381);
or U2579 (N_2579,N_1058,N_1745);
xor U2580 (N_2580,N_1915,N_1380);
nor U2581 (N_2581,N_1706,N_1939);
or U2582 (N_2582,N_1012,N_1436);
or U2583 (N_2583,N_1375,N_1122);
or U2584 (N_2584,N_1772,N_1750);
xor U2585 (N_2585,N_1097,N_1428);
and U2586 (N_2586,N_1858,N_1970);
nand U2587 (N_2587,N_1187,N_1882);
or U2588 (N_2588,N_1883,N_1815);
and U2589 (N_2589,N_1603,N_1330);
or U2590 (N_2590,N_1091,N_1057);
nand U2591 (N_2591,N_1862,N_1141);
nand U2592 (N_2592,N_1758,N_1589);
and U2593 (N_2593,N_1215,N_1435);
xor U2594 (N_2594,N_1379,N_1211);
or U2595 (N_2595,N_1995,N_1060);
nor U2596 (N_2596,N_1216,N_1394);
nor U2597 (N_2597,N_1266,N_1170);
or U2598 (N_2598,N_1567,N_1695);
nor U2599 (N_2599,N_1207,N_1940);
and U2600 (N_2600,N_1181,N_1134);
nor U2601 (N_2601,N_1070,N_1944);
and U2602 (N_2602,N_1860,N_1893);
or U2603 (N_2603,N_1667,N_1167);
nor U2604 (N_2604,N_1259,N_1304);
and U2605 (N_2605,N_1448,N_1722);
nor U2606 (N_2606,N_1224,N_1334);
nor U2607 (N_2607,N_1312,N_1540);
nor U2608 (N_2608,N_1850,N_1504);
or U2609 (N_2609,N_1776,N_1622);
and U2610 (N_2610,N_1347,N_1401);
and U2611 (N_2611,N_1709,N_1582);
nand U2612 (N_2612,N_1432,N_1150);
nand U2613 (N_2613,N_1153,N_1495);
nand U2614 (N_2614,N_1077,N_1276);
nand U2615 (N_2615,N_1605,N_1649);
nand U2616 (N_2616,N_1428,N_1435);
or U2617 (N_2617,N_1042,N_1789);
or U2618 (N_2618,N_1304,N_1537);
or U2619 (N_2619,N_1016,N_1976);
and U2620 (N_2620,N_1189,N_1260);
xor U2621 (N_2621,N_1258,N_1345);
xnor U2622 (N_2622,N_1187,N_1071);
or U2623 (N_2623,N_1275,N_1889);
nand U2624 (N_2624,N_1532,N_1761);
nand U2625 (N_2625,N_1622,N_1402);
and U2626 (N_2626,N_1583,N_1446);
and U2627 (N_2627,N_1835,N_1715);
xor U2628 (N_2628,N_1899,N_1299);
nand U2629 (N_2629,N_1973,N_1339);
nor U2630 (N_2630,N_1657,N_1943);
or U2631 (N_2631,N_1496,N_1220);
xnor U2632 (N_2632,N_1126,N_1804);
and U2633 (N_2633,N_1521,N_1524);
nor U2634 (N_2634,N_1189,N_1226);
xnor U2635 (N_2635,N_1173,N_1965);
or U2636 (N_2636,N_1469,N_1494);
nand U2637 (N_2637,N_1583,N_1440);
nor U2638 (N_2638,N_1962,N_1491);
nor U2639 (N_2639,N_1683,N_1526);
or U2640 (N_2640,N_1977,N_1204);
nand U2641 (N_2641,N_1719,N_1264);
nand U2642 (N_2642,N_1494,N_1939);
or U2643 (N_2643,N_1407,N_1054);
nand U2644 (N_2644,N_1434,N_1538);
nand U2645 (N_2645,N_1758,N_1616);
and U2646 (N_2646,N_1895,N_1448);
nand U2647 (N_2647,N_1250,N_1213);
nand U2648 (N_2648,N_1196,N_1878);
and U2649 (N_2649,N_1497,N_1383);
and U2650 (N_2650,N_1252,N_1902);
nand U2651 (N_2651,N_1416,N_1873);
xor U2652 (N_2652,N_1563,N_1767);
or U2653 (N_2653,N_1474,N_1285);
or U2654 (N_2654,N_1102,N_1623);
xor U2655 (N_2655,N_1548,N_1216);
and U2656 (N_2656,N_1332,N_1442);
and U2657 (N_2657,N_1035,N_1319);
or U2658 (N_2658,N_1349,N_1007);
and U2659 (N_2659,N_1303,N_1867);
nand U2660 (N_2660,N_1242,N_1119);
nor U2661 (N_2661,N_1531,N_1987);
or U2662 (N_2662,N_1571,N_1252);
xor U2663 (N_2663,N_1887,N_1729);
and U2664 (N_2664,N_1837,N_1243);
nand U2665 (N_2665,N_1008,N_1428);
nand U2666 (N_2666,N_1919,N_1696);
nor U2667 (N_2667,N_1072,N_1706);
and U2668 (N_2668,N_1392,N_1005);
or U2669 (N_2669,N_1650,N_1615);
and U2670 (N_2670,N_1780,N_1557);
nand U2671 (N_2671,N_1799,N_1715);
nor U2672 (N_2672,N_1852,N_1114);
nor U2673 (N_2673,N_1613,N_1110);
nor U2674 (N_2674,N_1731,N_1788);
and U2675 (N_2675,N_1781,N_1692);
or U2676 (N_2676,N_1763,N_1728);
or U2677 (N_2677,N_1372,N_1637);
nor U2678 (N_2678,N_1247,N_1668);
nand U2679 (N_2679,N_1757,N_1622);
and U2680 (N_2680,N_1883,N_1236);
or U2681 (N_2681,N_1907,N_1464);
nor U2682 (N_2682,N_1170,N_1276);
nor U2683 (N_2683,N_1966,N_1084);
or U2684 (N_2684,N_1701,N_1730);
xnor U2685 (N_2685,N_1440,N_1133);
xor U2686 (N_2686,N_1719,N_1542);
nor U2687 (N_2687,N_1726,N_1019);
xnor U2688 (N_2688,N_1903,N_1021);
and U2689 (N_2689,N_1619,N_1038);
and U2690 (N_2690,N_1767,N_1926);
xnor U2691 (N_2691,N_1178,N_1800);
and U2692 (N_2692,N_1031,N_1900);
or U2693 (N_2693,N_1587,N_1127);
or U2694 (N_2694,N_1986,N_1172);
nor U2695 (N_2695,N_1510,N_1319);
or U2696 (N_2696,N_1469,N_1976);
nand U2697 (N_2697,N_1217,N_1607);
xnor U2698 (N_2698,N_1131,N_1262);
nand U2699 (N_2699,N_1626,N_1192);
and U2700 (N_2700,N_1223,N_1977);
xnor U2701 (N_2701,N_1994,N_1441);
xor U2702 (N_2702,N_1658,N_1464);
nor U2703 (N_2703,N_1697,N_1519);
xnor U2704 (N_2704,N_1419,N_1847);
and U2705 (N_2705,N_1726,N_1635);
nand U2706 (N_2706,N_1220,N_1452);
and U2707 (N_2707,N_1226,N_1445);
or U2708 (N_2708,N_1615,N_1304);
xnor U2709 (N_2709,N_1951,N_1467);
xor U2710 (N_2710,N_1495,N_1169);
nand U2711 (N_2711,N_1344,N_1282);
and U2712 (N_2712,N_1815,N_1824);
nand U2713 (N_2713,N_1771,N_1527);
nand U2714 (N_2714,N_1125,N_1769);
or U2715 (N_2715,N_1796,N_1202);
xnor U2716 (N_2716,N_1044,N_1741);
and U2717 (N_2717,N_1018,N_1884);
nand U2718 (N_2718,N_1108,N_1859);
nor U2719 (N_2719,N_1403,N_1801);
or U2720 (N_2720,N_1517,N_1882);
xnor U2721 (N_2721,N_1546,N_1068);
nand U2722 (N_2722,N_1446,N_1419);
or U2723 (N_2723,N_1160,N_1592);
xnor U2724 (N_2724,N_1977,N_1051);
and U2725 (N_2725,N_1208,N_1183);
and U2726 (N_2726,N_1369,N_1918);
or U2727 (N_2727,N_1769,N_1799);
nand U2728 (N_2728,N_1010,N_1353);
or U2729 (N_2729,N_1477,N_1164);
nor U2730 (N_2730,N_1882,N_1095);
nand U2731 (N_2731,N_1379,N_1512);
nor U2732 (N_2732,N_1709,N_1177);
and U2733 (N_2733,N_1486,N_1358);
or U2734 (N_2734,N_1964,N_1489);
nand U2735 (N_2735,N_1149,N_1866);
nand U2736 (N_2736,N_1952,N_1469);
and U2737 (N_2737,N_1768,N_1091);
xor U2738 (N_2738,N_1212,N_1553);
and U2739 (N_2739,N_1170,N_1314);
nand U2740 (N_2740,N_1577,N_1297);
and U2741 (N_2741,N_1187,N_1624);
xor U2742 (N_2742,N_1955,N_1240);
or U2743 (N_2743,N_1608,N_1710);
and U2744 (N_2744,N_1800,N_1044);
nand U2745 (N_2745,N_1063,N_1441);
and U2746 (N_2746,N_1418,N_1217);
nand U2747 (N_2747,N_1282,N_1987);
xnor U2748 (N_2748,N_1263,N_1510);
nand U2749 (N_2749,N_1317,N_1632);
and U2750 (N_2750,N_1188,N_1613);
or U2751 (N_2751,N_1611,N_1173);
nand U2752 (N_2752,N_1958,N_1715);
nand U2753 (N_2753,N_1351,N_1581);
and U2754 (N_2754,N_1679,N_1837);
xnor U2755 (N_2755,N_1554,N_1958);
and U2756 (N_2756,N_1086,N_1863);
and U2757 (N_2757,N_1202,N_1766);
xor U2758 (N_2758,N_1958,N_1211);
xnor U2759 (N_2759,N_1640,N_1167);
nor U2760 (N_2760,N_1383,N_1881);
xnor U2761 (N_2761,N_1912,N_1677);
and U2762 (N_2762,N_1707,N_1304);
and U2763 (N_2763,N_1171,N_1849);
and U2764 (N_2764,N_1934,N_1773);
nand U2765 (N_2765,N_1935,N_1433);
and U2766 (N_2766,N_1164,N_1497);
and U2767 (N_2767,N_1031,N_1647);
nand U2768 (N_2768,N_1523,N_1663);
nand U2769 (N_2769,N_1422,N_1494);
or U2770 (N_2770,N_1746,N_1559);
nand U2771 (N_2771,N_1171,N_1794);
nor U2772 (N_2772,N_1188,N_1064);
nor U2773 (N_2773,N_1689,N_1489);
nand U2774 (N_2774,N_1566,N_1025);
xnor U2775 (N_2775,N_1967,N_1429);
or U2776 (N_2776,N_1308,N_1242);
xnor U2777 (N_2777,N_1693,N_1827);
and U2778 (N_2778,N_1327,N_1906);
or U2779 (N_2779,N_1230,N_1840);
nand U2780 (N_2780,N_1117,N_1048);
xor U2781 (N_2781,N_1399,N_1144);
and U2782 (N_2782,N_1014,N_1802);
nor U2783 (N_2783,N_1712,N_1402);
xnor U2784 (N_2784,N_1990,N_1960);
nor U2785 (N_2785,N_1973,N_1710);
nor U2786 (N_2786,N_1337,N_1700);
or U2787 (N_2787,N_1990,N_1399);
and U2788 (N_2788,N_1406,N_1242);
xor U2789 (N_2789,N_1726,N_1323);
nand U2790 (N_2790,N_1921,N_1387);
and U2791 (N_2791,N_1171,N_1568);
or U2792 (N_2792,N_1671,N_1606);
nor U2793 (N_2793,N_1357,N_1364);
nor U2794 (N_2794,N_1951,N_1991);
or U2795 (N_2795,N_1399,N_1880);
xnor U2796 (N_2796,N_1984,N_1026);
and U2797 (N_2797,N_1708,N_1675);
xor U2798 (N_2798,N_1465,N_1456);
nor U2799 (N_2799,N_1309,N_1970);
or U2800 (N_2800,N_1032,N_1279);
or U2801 (N_2801,N_1703,N_1640);
nor U2802 (N_2802,N_1383,N_1361);
xnor U2803 (N_2803,N_1655,N_1813);
xnor U2804 (N_2804,N_1646,N_1412);
and U2805 (N_2805,N_1080,N_1654);
or U2806 (N_2806,N_1186,N_1162);
xnor U2807 (N_2807,N_1305,N_1004);
nor U2808 (N_2808,N_1158,N_1172);
or U2809 (N_2809,N_1601,N_1194);
xnor U2810 (N_2810,N_1627,N_1583);
or U2811 (N_2811,N_1170,N_1404);
or U2812 (N_2812,N_1417,N_1923);
xnor U2813 (N_2813,N_1095,N_1201);
nand U2814 (N_2814,N_1939,N_1048);
nor U2815 (N_2815,N_1262,N_1603);
xnor U2816 (N_2816,N_1738,N_1492);
xor U2817 (N_2817,N_1239,N_1075);
or U2818 (N_2818,N_1765,N_1520);
or U2819 (N_2819,N_1841,N_1097);
nor U2820 (N_2820,N_1744,N_1410);
xor U2821 (N_2821,N_1568,N_1480);
xnor U2822 (N_2822,N_1273,N_1629);
nor U2823 (N_2823,N_1903,N_1714);
or U2824 (N_2824,N_1379,N_1540);
and U2825 (N_2825,N_1408,N_1088);
and U2826 (N_2826,N_1038,N_1978);
nor U2827 (N_2827,N_1363,N_1352);
xnor U2828 (N_2828,N_1932,N_1144);
xor U2829 (N_2829,N_1327,N_1929);
nor U2830 (N_2830,N_1852,N_1390);
xnor U2831 (N_2831,N_1940,N_1578);
xnor U2832 (N_2832,N_1924,N_1690);
or U2833 (N_2833,N_1648,N_1671);
and U2834 (N_2834,N_1264,N_1703);
nand U2835 (N_2835,N_1482,N_1786);
nand U2836 (N_2836,N_1242,N_1292);
nor U2837 (N_2837,N_1066,N_1878);
nand U2838 (N_2838,N_1525,N_1133);
nand U2839 (N_2839,N_1953,N_1456);
nor U2840 (N_2840,N_1404,N_1783);
and U2841 (N_2841,N_1893,N_1946);
or U2842 (N_2842,N_1228,N_1093);
or U2843 (N_2843,N_1532,N_1459);
and U2844 (N_2844,N_1170,N_1285);
and U2845 (N_2845,N_1760,N_1566);
nand U2846 (N_2846,N_1825,N_1692);
or U2847 (N_2847,N_1853,N_1654);
or U2848 (N_2848,N_1626,N_1045);
nand U2849 (N_2849,N_1648,N_1196);
nor U2850 (N_2850,N_1403,N_1142);
or U2851 (N_2851,N_1019,N_1291);
or U2852 (N_2852,N_1399,N_1511);
and U2853 (N_2853,N_1589,N_1854);
or U2854 (N_2854,N_1217,N_1372);
xnor U2855 (N_2855,N_1990,N_1173);
nor U2856 (N_2856,N_1249,N_1670);
nor U2857 (N_2857,N_1850,N_1034);
and U2858 (N_2858,N_1888,N_1120);
or U2859 (N_2859,N_1697,N_1174);
xor U2860 (N_2860,N_1482,N_1684);
xor U2861 (N_2861,N_1070,N_1299);
nand U2862 (N_2862,N_1442,N_1217);
or U2863 (N_2863,N_1699,N_1032);
and U2864 (N_2864,N_1520,N_1258);
and U2865 (N_2865,N_1074,N_1588);
xnor U2866 (N_2866,N_1068,N_1367);
nor U2867 (N_2867,N_1884,N_1215);
and U2868 (N_2868,N_1123,N_1848);
or U2869 (N_2869,N_1358,N_1923);
nor U2870 (N_2870,N_1600,N_1249);
and U2871 (N_2871,N_1679,N_1634);
nand U2872 (N_2872,N_1947,N_1554);
xor U2873 (N_2873,N_1597,N_1439);
nand U2874 (N_2874,N_1000,N_1445);
xor U2875 (N_2875,N_1980,N_1850);
nor U2876 (N_2876,N_1551,N_1076);
nor U2877 (N_2877,N_1804,N_1418);
nand U2878 (N_2878,N_1984,N_1195);
or U2879 (N_2879,N_1857,N_1231);
or U2880 (N_2880,N_1905,N_1191);
and U2881 (N_2881,N_1120,N_1765);
nor U2882 (N_2882,N_1727,N_1155);
nor U2883 (N_2883,N_1664,N_1570);
or U2884 (N_2884,N_1605,N_1117);
xnor U2885 (N_2885,N_1043,N_1655);
xnor U2886 (N_2886,N_1473,N_1515);
xnor U2887 (N_2887,N_1192,N_1483);
nor U2888 (N_2888,N_1324,N_1508);
nor U2889 (N_2889,N_1865,N_1573);
nor U2890 (N_2890,N_1152,N_1758);
nand U2891 (N_2891,N_1902,N_1334);
nor U2892 (N_2892,N_1158,N_1339);
nand U2893 (N_2893,N_1318,N_1754);
xnor U2894 (N_2894,N_1320,N_1914);
xor U2895 (N_2895,N_1706,N_1687);
nand U2896 (N_2896,N_1551,N_1124);
and U2897 (N_2897,N_1198,N_1248);
nand U2898 (N_2898,N_1536,N_1847);
and U2899 (N_2899,N_1036,N_1049);
xor U2900 (N_2900,N_1495,N_1818);
nand U2901 (N_2901,N_1458,N_1460);
xnor U2902 (N_2902,N_1791,N_1302);
nor U2903 (N_2903,N_1927,N_1879);
nor U2904 (N_2904,N_1746,N_1316);
or U2905 (N_2905,N_1810,N_1380);
nor U2906 (N_2906,N_1908,N_1180);
nor U2907 (N_2907,N_1022,N_1763);
xnor U2908 (N_2908,N_1922,N_1903);
nor U2909 (N_2909,N_1076,N_1531);
nand U2910 (N_2910,N_1984,N_1993);
or U2911 (N_2911,N_1517,N_1923);
nor U2912 (N_2912,N_1009,N_1846);
and U2913 (N_2913,N_1310,N_1294);
and U2914 (N_2914,N_1791,N_1475);
and U2915 (N_2915,N_1323,N_1048);
or U2916 (N_2916,N_1878,N_1291);
and U2917 (N_2917,N_1575,N_1553);
or U2918 (N_2918,N_1976,N_1078);
and U2919 (N_2919,N_1818,N_1454);
or U2920 (N_2920,N_1248,N_1417);
or U2921 (N_2921,N_1460,N_1764);
and U2922 (N_2922,N_1815,N_1652);
xnor U2923 (N_2923,N_1213,N_1706);
and U2924 (N_2924,N_1104,N_1219);
nand U2925 (N_2925,N_1158,N_1247);
and U2926 (N_2926,N_1646,N_1374);
and U2927 (N_2927,N_1682,N_1806);
nand U2928 (N_2928,N_1177,N_1902);
and U2929 (N_2929,N_1366,N_1126);
or U2930 (N_2930,N_1746,N_1544);
xnor U2931 (N_2931,N_1307,N_1154);
nor U2932 (N_2932,N_1021,N_1080);
nand U2933 (N_2933,N_1231,N_1139);
xnor U2934 (N_2934,N_1637,N_1814);
xnor U2935 (N_2935,N_1922,N_1830);
nand U2936 (N_2936,N_1938,N_1300);
and U2937 (N_2937,N_1974,N_1361);
and U2938 (N_2938,N_1847,N_1528);
nand U2939 (N_2939,N_1725,N_1623);
or U2940 (N_2940,N_1768,N_1378);
nor U2941 (N_2941,N_1673,N_1266);
nor U2942 (N_2942,N_1277,N_1640);
nor U2943 (N_2943,N_1058,N_1352);
and U2944 (N_2944,N_1532,N_1612);
xor U2945 (N_2945,N_1380,N_1962);
or U2946 (N_2946,N_1940,N_1266);
and U2947 (N_2947,N_1095,N_1701);
xor U2948 (N_2948,N_1201,N_1763);
xor U2949 (N_2949,N_1074,N_1243);
and U2950 (N_2950,N_1383,N_1223);
nand U2951 (N_2951,N_1594,N_1220);
xnor U2952 (N_2952,N_1442,N_1358);
xnor U2953 (N_2953,N_1001,N_1368);
or U2954 (N_2954,N_1360,N_1214);
nand U2955 (N_2955,N_1297,N_1156);
xnor U2956 (N_2956,N_1963,N_1149);
nor U2957 (N_2957,N_1523,N_1217);
nand U2958 (N_2958,N_1553,N_1125);
nand U2959 (N_2959,N_1026,N_1762);
nand U2960 (N_2960,N_1722,N_1468);
or U2961 (N_2961,N_1379,N_1393);
and U2962 (N_2962,N_1518,N_1834);
xor U2963 (N_2963,N_1065,N_1806);
nor U2964 (N_2964,N_1455,N_1124);
and U2965 (N_2965,N_1498,N_1586);
nor U2966 (N_2966,N_1595,N_1724);
xor U2967 (N_2967,N_1246,N_1112);
nand U2968 (N_2968,N_1443,N_1824);
xor U2969 (N_2969,N_1853,N_1234);
xnor U2970 (N_2970,N_1379,N_1187);
xnor U2971 (N_2971,N_1968,N_1938);
and U2972 (N_2972,N_1433,N_1896);
nand U2973 (N_2973,N_1188,N_1136);
xor U2974 (N_2974,N_1120,N_1621);
nor U2975 (N_2975,N_1277,N_1611);
or U2976 (N_2976,N_1593,N_1407);
xnor U2977 (N_2977,N_1139,N_1451);
or U2978 (N_2978,N_1598,N_1520);
nand U2979 (N_2979,N_1258,N_1891);
and U2980 (N_2980,N_1406,N_1862);
nand U2981 (N_2981,N_1379,N_1626);
or U2982 (N_2982,N_1792,N_1483);
xor U2983 (N_2983,N_1819,N_1256);
nor U2984 (N_2984,N_1111,N_1545);
or U2985 (N_2985,N_1706,N_1659);
or U2986 (N_2986,N_1522,N_1060);
nand U2987 (N_2987,N_1909,N_1785);
xnor U2988 (N_2988,N_1978,N_1547);
and U2989 (N_2989,N_1356,N_1349);
nand U2990 (N_2990,N_1111,N_1137);
nand U2991 (N_2991,N_1628,N_1888);
and U2992 (N_2992,N_1348,N_1877);
and U2993 (N_2993,N_1626,N_1163);
and U2994 (N_2994,N_1901,N_1443);
or U2995 (N_2995,N_1348,N_1398);
or U2996 (N_2996,N_1404,N_1704);
or U2997 (N_2997,N_1294,N_1380);
and U2998 (N_2998,N_1451,N_1211);
or U2999 (N_2999,N_1675,N_1831);
or U3000 (N_3000,N_2566,N_2121);
and U3001 (N_3001,N_2657,N_2791);
xor U3002 (N_3002,N_2222,N_2495);
nand U3003 (N_3003,N_2689,N_2831);
and U3004 (N_3004,N_2843,N_2888);
nor U3005 (N_3005,N_2771,N_2329);
nor U3006 (N_3006,N_2612,N_2517);
or U3007 (N_3007,N_2340,N_2110);
xor U3008 (N_3008,N_2536,N_2950);
nor U3009 (N_3009,N_2932,N_2377);
or U3010 (N_3010,N_2840,N_2181);
and U3011 (N_3011,N_2993,N_2907);
nand U3012 (N_3012,N_2025,N_2698);
nand U3013 (N_3013,N_2618,N_2113);
nand U3014 (N_3014,N_2229,N_2451);
xor U3015 (N_3015,N_2708,N_2572);
or U3016 (N_3016,N_2453,N_2974);
nor U3017 (N_3017,N_2449,N_2728);
nand U3018 (N_3018,N_2962,N_2189);
nor U3019 (N_3019,N_2382,N_2366);
xnor U3020 (N_3020,N_2992,N_2802);
nand U3021 (N_3021,N_2349,N_2193);
nand U3022 (N_3022,N_2529,N_2481);
nand U3023 (N_3023,N_2159,N_2763);
xnor U3024 (N_3024,N_2626,N_2887);
and U3025 (N_3025,N_2872,N_2239);
xnor U3026 (N_3026,N_2119,N_2798);
nand U3027 (N_3027,N_2910,N_2716);
and U3028 (N_3028,N_2849,N_2639);
nand U3029 (N_3029,N_2278,N_2635);
xor U3030 (N_3030,N_2866,N_2851);
nand U3031 (N_3031,N_2498,N_2174);
nor U3032 (N_3032,N_2939,N_2770);
nor U3033 (N_3033,N_2331,N_2833);
nand U3034 (N_3034,N_2800,N_2961);
nor U3035 (N_3035,N_2075,N_2394);
nand U3036 (N_3036,N_2345,N_2531);
nand U3037 (N_3037,N_2196,N_2376);
and U3038 (N_3038,N_2880,N_2282);
nor U3039 (N_3039,N_2699,N_2839);
nand U3040 (N_3040,N_2631,N_2818);
nor U3041 (N_3041,N_2805,N_2867);
or U3042 (N_3042,N_2368,N_2646);
and U3043 (N_3043,N_2494,N_2504);
and U3044 (N_3044,N_2623,N_2673);
xnor U3045 (N_3045,N_2984,N_2560);
or U3046 (N_3046,N_2314,N_2985);
nor U3047 (N_3047,N_2172,N_2287);
and U3048 (N_3048,N_2408,N_2948);
nor U3049 (N_3049,N_2968,N_2107);
xnor U3050 (N_3050,N_2393,N_2319);
or U3051 (N_3051,N_2885,N_2938);
nor U3052 (N_3052,N_2123,N_2485);
or U3053 (N_3053,N_2564,N_2445);
and U3054 (N_3054,N_2252,N_2004);
nor U3055 (N_3055,N_2773,N_2343);
nor U3056 (N_3056,N_2064,N_2803);
xor U3057 (N_3057,N_2078,N_2098);
nand U3058 (N_3058,N_2459,N_2940);
or U3059 (N_3059,N_2778,N_2898);
and U3060 (N_3060,N_2678,N_2761);
and U3061 (N_3061,N_2999,N_2783);
nand U3062 (N_3062,N_2593,N_2295);
xor U3063 (N_3063,N_2475,N_2914);
or U3064 (N_3064,N_2916,N_2093);
nand U3065 (N_3065,N_2378,N_2836);
or U3066 (N_3066,N_2488,N_2160);
xnor U3067 (N_3067,N_2620,N_2071);
or U3068 (N_3068,N_2362,N_2302);
and U3069 (N_3069,N_2801,N_2288);
nor U3070 (N_3070,N_2500,N_2554);
nor U3071 (N_3071,N_2884,N_2232);
nand U3072 (N_3072,N_2212,N_2365);
nor U3073 (N_3073,N_2541,N_2662);
and U3074 (N_3074,N_2403,N_2902);
xnor U3075 (N_3075,N_2519,N_2118);
or U3076 (N_3076,N_2289,N_2081);
or U3077 (N_3077,N_2019,N_2129);
nand U3078 (N_3078,N_2431,N_2260);
nand U3079 (N_3079,N_2311,N_2591);
or U3080 (N_3080,N_2934,N_2469);
or U3081 (N_3081,N_2949,N_2268);
nand U3082 (N_3082,N_2061,N_2178);
xnor U3083 (N_3083,N_2850,N_2161);
nand U3084 (N_3084,N_2419,N_2234);
or U3085 (N_3085,N_2294,N_2450);
nand U3086 (N_3086,N_2757,N_2779);
and U3087 (N_3087,N_2751,N_2398);
nand U3088 (N_3088,N_2503,N_2165);
or U3089 (N_3089,N_2055,N_2405);
or U3090 (N_3090,N_2069,N_2003);
nor U3091 (N_3091,N_2520,N_2957);
nand U3092 (N_3092,N_2052,N_2972);
and U3093 (N_3093,N_2223,N_2760);
nand U3094 (N_3094,N_2447,N_2556);
nand U3095 (N_3095,N_2568,N_2058);
or U3096 (N_3096,N_2651,N_2099);
xor U3097 (N_3097,N_2354,N_2236);
or U3098 (N_3098,N_2417,N_2927);
nor U3099 (N_3099,N_2404,N_2086);
nor U3100 (N_3100,N_2273,N_2685);
or U3101 (N_3101,N_2891,N_2175);
and U3102 (N_3102,N_2956,N_2277);
nand U3103 (N_3103,N_2243,N_2903);
and U3104 (N_3104,N_2442,N_2266);
or U3105 (N_3105,N_2913,N_2045);
nand U3106 (N_3106,N_2307,N_2952);
xnor U3107 (N_3107,N_2544,N_2870);
and U3108 (N_3108,N_2894,N_2518);
or U3109 (N_3109,N_2561,N_2996);
nand U3110 (N_3110,N_2293,N_2258);
and U3111 (N_3111,N_2422,N_2309);
nand U3112 (N_3112,N_2000,N_2039);
nor U3113 (N_3113,N_2753,N_2549);
or U3114 (N_3114,N_2043,N_2983);
xnor U3115 (N_3115,N_2653,N_2524);
and U3116 (N_3116,N_2721,N_2718);
nor U3117 (N_3117,N_2599,N_2477);
and U3118 (N_3118,N_2158,N_2216);
nor U3119 (N_3119,N_2144,N_2040);
nand U3120 (N_3120,N_2603,N_2318);
nand U3121 (N_3121,N_2490,N_2690);
xnor U3122 (N_3122,N_2863,N_2660);
nand U3123 (N_3123,N_2946,N_2614);
and U3124 (N_3124,N_2316,N_2912);
or U3125 (N_3125,N_2242,N_2512);
nor U3126 (N_3126,N_2100,N_2929);
or U3127 (N_3127,N_2901,N_2248);
nand U3128 (N_3128,N_2649,N_2820);
nand U3129 (N_3129,N_2767,N_2346);
xor U3130 (N_3130,N_2251,N_2135);
and U3131 (N_3131,N_2363,N_2947);
nor U3132 (N_3132,N_2575,N_2875);
or U3133 (N_3133,N_2748,N_2226);
nor U3134 (N_3134,N_2864,N_2579);
nor U3135 (N_3135,N_2204,N_2672);
nor U3136 (N_3136,N_2819,N_2238);
nand U3137 (N_3137,N_2816,N_2067);
and U3138 (N_3138,N_2457,N_2571);
nor U3139 (N_3139,N_2857,N_2131);
nand U3140 (N_3140,N_2070,N_2637);
xor U3141 (N_3141,N_2513,N_2641);
and U3142 (N_3142,N_2928,N_2326);
xnor U3143 (N_3143,N_2177,N_2682);
nor U3144 (N_3144,N_2908,N_2303);
nand U3145 (N_3145,N_2976,N_2923);
nor U3146 (N_3146,N_2528,N_2465);
nand U3147 (N_3147,N_2925,N_2522);
or U3148 (N_3148,N_2942,N_2291);
nor U3149 (N_3149,N_2742,N_2876);
nand U3150 (N_3150,N_2979,N_2994);
xnor U3151 (N_3151,N_2730,N_2227);
nand U3152 (N_3152,N_2693,N_2815);
and U3153 (N_3153,N_2301,N_2665);
xnor U3154 (N_3154,N_2407,N_2640);
nand U3155 (N_3155,N_2900,N_2374);
and U3156 (N_3156,N_2991,N_2735);
nor U3157 (N_3157,N_2588,N_2023);
nor U3158 (N_3158,N_2497,N_2899);
or U3159 (N_3159,N_2625,N_2194);
nand U3160 (N_3160,N_2466,N_2713);
and U3161 (N_3161,N_2995,N_2214);
xnor U3162 (N_3162,N_2063,N_2147);
nand U3163 (N_3163,N_2677,N_2036);
xnor U3164 (N_3164,N_2480,N_2463);
nand U3165 (N_3165,N_2122,N_2022);
nor U3166 (N_3166,N_2132,N_2796);
nand U3167 (N_3167,N_2245,N_2250);
nor U3168 (N_3168,N_2590,N_2435);
xor U3169 (N_3169,N_2478,N_2842);
xor U3170 (N_3170,N_2370,N_2595);
nand U3171 (N_3171,N_2681,N_2613);
nor U3172 (N_3172,N_2854,N_2364);
and U3173 (N_3173,N_2941,N_2338);
and U3174 (N_3174,N_2281,N_2521);
or U3175 (N_3175,N_2719,N_2654);
and U3176 (N_3176,N_2010,N_2084);
or U3177 (N_3177,N_2874,N_2198);
nand U3178 (N_3178,N_2254,N_2171);
and U3179 (N_3179,N_2511,N_2146);
nand U3180 (N_3180,N_2967,N_2987);
and U3181 (N_3181,N_2865,N_2601);
and U3182 (N_3182,N_2632,N_2986);
nor U3183 (N_3183,N_2199,N_2200);
or U3184 (N_3184,N_2548,N_2026);
xor U3185 (N_3185,N_2090,N_2482);
nor U3186 (N_3186,N_2711,N_2016);
or U3187 (N_3187,N_2028,N_2697);
nor U3188 (N_3188,N_2889,N_2608);
and U3189 (N_3189,N_2822,N_2674);
xor U3190 (N_3190,N_2904,N_2412);
and U3191 (N_3191,N_2092,N_2797);
nor U3192 (N_3192,N_2104,N_2552);
or U3193 (N_3193,N_2249,N_2873);
and U3194 (N_3194,N_2809,N_2072);
or U3195 (N_3195,N_2013,N_2051);
or U3196 (N_3196,N_2461,N_2211);
or U3197 (N_3197,N_2562,N_2179);
xnor U3198 (N_3198,N_2335,N_2551);
or U3199 (N_3199,N_2397,N_2811);
nand U3200 (N_3200,N_2306,N_2415);
nand U3201 (N_3201,N_2452,N_2321);
or U3202 (N_3202,N_2464,N_2691);
and U3203 (N_3203,N_2731,N_2741);
nand U3204 (N_3204,N_2484,N_2031);
nand U3205 (N_3205,N_2675,N_2772);
and U3206 (N_3206,N_2642,N_2710);
xnor U3207 (N_3207,N_2184,N_2073);
or U3208 (N_3208,N_2953,N_2387);
xor U3209 (N_3209,N_2759,N_2082);
xor U3210 (N_3210,N_2844,N_2024);
or U3211 (N_3211,N_2380,N_2703);
or U3212 (N_3212,N_2333,N_2943);
and U3213 (N_3213,N_2539,N_2788);
nor U3214 (N_3214,N_2656,N_2433);
or U3215 (N_3215,N_2269,N_2421);
and U3216 (N_3216,N_2299,N_2777);
nand U3217 (N_3217,N_2297,N_2205);
nand U3218 (N_3218,N_2154,N_2074);
nor U3219 (N_3219,N_2963,N_2032);
and U3220 (N_3220,N_2758,N_2821);
nor U3221 (N_3221,N_2667,N_2565);
or U3222 (N_3222,N_2356,N_2997);
and U3223 (N_3223,N_2666,N_2807);
nand U3224 (N_3224,N_2392,N_2337);
nor U3225 (N_3225,N_2180,N_2853);
xnor U3226 (N_3226,N_2810,N_2806);
nand U3227 (N_3227,N_2203,N_2438);
nand U3228 (N_3228,N_2707,N_2592);
and U3229 (N_3229,N_2128,N_2347);
nand U3230 (N_3230,N_2722,N_2046);
nand U3231 (N_3231,N_2041,N_2095);
nand U3232 (N_3232,N_2091,N_2372);
nand U3233 (N_3233,N_2510,N_2396);
nand U3234 (N_3234,N_2155,N_2162);
and U3235 (N_3235,N_2430,N_2823);
xor U3236 (N_3236,N_2755,N_2924);
nor U3237 (N_3237,N_2555,N_2877);
or U3238 (N_3238,N_2706,N_2395);
and U3239 (N_3239,N_2279,N_2780);
xor U3240 (N_3240,N_2576,N_2259);
or U3241 (N_3241,N_2785,N_2182);
nor U3242 (N_3242,N_2018,N_2835);
or U3243 (N_3243,N_2582,N_2501);
xor U3244 (N_3244,N_2225,N_2813);
and U3245 (N_3245,N_2076,N_2327);
and U3246 (N_3246,N_2506,N_2507);
nor U3247 (N_3247,N_2587,N_2633);
nor U3248 (N_3248,N_2607,N_2879);
nand U3249 (N_3249,N_2208,N_2097);
or U3250 (N_3250,N_2786,N_2508);
xor U3251 (N_3251,N_2683,N_2153);
xor U3252 (N_3252,N_2729,N_2400);
or U3253 (N_3253,N_2460,N_2765);
xor U3254 (N_3254,N_2604,N_2926);
nand U3255 (N_3255,N_2817,N_2784);
or U3256 (N_3256,N_2381,N_2176);
nand U3257 (N_3257,N_2643,N_2661);
or U3258 (N_3258,N_2860,N_2700);
nor U3259 (N_3259,N_2149,N_2971);
or U3260 (N_3260,N_2261,N_2066);
xor U3261 (N_3261,N_2896,N_2109);
or U3262 (N_3262,N_2411,N_2265);
nand U3263 (N_3263,N_2157,N_2695);
or U3264 (N_3264,N_2136,N_2371);
or U3265 (N_3265,N_2402,N_2322);
nor U3266 (N_3266,N_2726,N_2933);
nand U3267 (N_3267,N_2712,N_2606);
and U3268 (N_3268,N_2824,N_2325);
nand U3269 (N_3269,N_2351,N_2312);
or U3270 (N_3270,N_2334,N_2627);
nand U3271 (N_3271,N_2183,N_2304);
nand U3272 (N_3272,N_2424,N_2859);
and U3273 (N_3273,N_2692,N_2483);
xor U3274 (N_3274,N_2112,N_2862);
nor U3275 (N_3275,N_2652,N_2298);
and U3276 (N_3276,N_2981,N_2848);
nor U3277 (N_3277,N_2472,N_2747);
nor U3278 (N_3278,N_2516,N_2878);
nor U3279 (N_3279,N_2704,N_2578);
and U3280 (N_3280,N_2882,N_2137);
or U3281 (N_3281,N_2399,N_2423);
nor U3282 (N_3282,N_2740,N_2909);
nor U3283 (N_3283,N_2057,N_2534);
xor U3284 (N_3284,N_2305,N_2630);
and U3285 (N_3285,N_2969,N_2414);
nand U3286 (N_3286,N_2530,N_2008);
nand U3287 (N_3287,N_2474,N_2317);
nor U3288 (N_3288,N_2829,N_2124);
nor U3289 (N_3289,N_2493,N_2341);
nor U3290 (N_3290,N_2663,N_2367);
nor U3291 (N_3291,N_2622,N_2869);
nand U3292 (N_3292,N_2496,N_2830);
xor U3293 (N_3293,N_2655,N_2492);
nand U3294 (N_3294,N_2585,N_2982);
or U3295 (N_3295,N_2426,N_2794);
nand U3296 (N_3296,N_2197,N_2744);
or U3297 (N_3297,N_2228,N_2042);
and U3298 (N_3298,N_2033,N_2456);
xnor U3299 (N_3299,N_2920,N_2284);
or U3300 (N_3300,N_2537,N_2418);
xor U3301 (N_3301,N_2733,N_2218);
or U3302 (N_3302,N_2436,N_2192);
xor U3303 (N_3303,N_2388,N_2958);
xnor U3304 (N_3304,N_2955,N_2975);
and U3305 (N_3305,N_2120,N_2355);
xnor U3306 (N_3306,N_2114,N_2115);
nor U3307 (N_3307,N_2776,N_2049);
nor U3308 (N_3308,N_2659,N_2668);
nor U3309 (N_3309,N_2454,N_2286);
and U3310 (N_3310,N_2702,N_2964);
nor U3311 (N_3311,N_2812,N_2473);
or U3312 (N_3312,N_2257,N_2001);
or U3313 (N_3313,N_2557,N_2201);
xnor U3314 (N_3314,N_2906,N_2077);
or U3315 (N_3315,N_2832,N_2737);
nand U3316 (N_3316,N_2068,N_2389);
or U3317 (N_3317,N_2413,N_2650);
or U3318 (N_3318,N_2116,N_2169);
nor U3319 (N_3319,N_2714,N_2240);
nor U3320 (N_3320,N_2684,N_2434);
or U3321 (N_3321,N_2002,N_2883);
and U3322 (N_3322,N_2837,N_2687);
or U3323 (N_3323,N_2267,N_2515);
nand U3324 (N_3324,N_2847,N_2029);
xor U3325 (N_3325,N_2296,N_2053);
or U3326 (N_3326,N_2550,N_2905);
nand U3327 (N_3327,N_2247,N_2416);
xnor U3328 (N_3328,N_2375,N_2038);
nand U3329 (N_3329,N_2750,N_2486);
or U3330 (N_3330,N_2237,N_2202);
or U3331 (N_3331,N_2918,N_2012);
or U3332 (N_3332,N_2432,N_2709);
nand U3333 (N_3333,N_2256,N_2523);
nor U3334 (N_3334,N_2315,N_2547);
and U3335 (N_3335,N_2369,N_2213);
or U3336 (N_3336,N_2930,N_2525);
nor U3337 (N_3337,N_2756,N_2152);
or U3338 (N_3338,N_2782,N_2921);
and U3339 (N_3339,N_2441,N_2117);
nand U3340 (N_3340,N_2059,N_2543);
nand U3341 (N_3341,N_2130,N_2330);
nor U3342 (N_3342,N_2108,N_2085);
or U3343 (N_3343,N_2998,N_2215);
nor U3344 (N_3344,N_2808,N_2954);
and U3345 (N_3345,N_2079,N_2616);
nand U3346 (N_3346,N_2060,N_2828);
and U3347 (N_3347,N_2479,N_2262);
or U3348 (N_3348,N_2006,N_2826);
nand U3349 (N_3349,N_2502,N_2186);
and U3350 (N_3350,N_2532,N_2580);
nor U3351 (N_3351,N_2007,N_2443);
xnor U3352 (N_3352,N_2037,N_2960);
xor U3353 (N_3353,N_2361,N_2209);
nor U3354 (N_3354,N_2336,N_2589);
xnor U3355 (N_3355,N_2409,N_2664);
or U3356 (N_3356,N_2283,N_2762);
or U3357 (N_3357,N_2644,N_2723);
and U3358 (N_3358,N_2035,N_2357);
or U3359 (N_3359,N_2720,N_2545);
nor U3360 (N_3360,N_2491,N_2044);
nand U3361 (N_3361,N_2233,N_2648);
and U3362 (N_3362,N_2384,N_2163);
xnor U3363 (N_3363,N_2080,N_2391);
and U3364 (N_3364,N_2936,N_2538);
nor U3365 (N_3365,N_2308,N_2636);
and U3366 (N_3366,N_2429,N_2439);
and U3367 (N_3367,N_2017,N_2246);
and U3368 (N_3368,N_2724,N_2094);
and U3369 (N_3369,N_2140,N_2944);
xnor U3370 (N_3370,N_2166,N_2138);
and U3371 (N_3371,N_2103,N_2795);
xor U3372 (N_3372,N_2792,N_2255);
nand U3373 (N_3373,N_2271,N_2386);
or U3374 (N_3374,N_2919,N_2977);
and U3375 (N_3375,N_2669,N_2970);
nand U3376 (N_3376,N_2126,N_2594);
or U3377 (N_3377,N_2263,N_2634);
xor U3378 (N_3378,N_2034,N_2280);
nand U3379 (N_3379,N_2359,N_2645);
xnor U3380 (N_3380,N_2527,N_2814);
and U3381 (N_3381,N_2567,N_2143);
or U3382 (N_3382,N_2168,N_2789);
xnor U3383 (N_3383,N_2696,N_2420);
or U3384 (N_3384,N_2127,N_2231);
and U3385 (N_3385,N_2047,N_2324);
and U3386 (N_3386,N_2185,N_2133);
and U3387 (N_3387,N_2945,N_2440);
xor U3388 (N_3388,N_2546,N_2509);
nor U3389 (N_3389,N_2111,N_2005);
and U3390 (N_3390,N_2581,N_2540);
nor U3391 (N_3391,N_2390,N_2360);
nor U3392 (N_3392,N_2573,N_2917);
and U3393 (N_3393,N_2980,N_2775);
xnor U3394 (N_3394,N_2272,N_2358);
nor U3395 (N_3395,N_2738,N_2385);
nor U3396 (N_3396,N_2804,N_2868);
or U3397 (N_3397,N_2027,N_2089);
nor U3398 (N_3398,N_2574,N_2734);
nor U3399 (N_3399,N_2526,N_2629);
nor U3400 (N_3400,N_2141,N_2332);
xor U3401 (N_3401,N_2951,N_2088);
nand U3402 (N_3402,N_2164,N_2167);
xnor U3403 (N_3403,N_2892,N_2766);
and U3404 (N_3404,N_2746,N_2739);
or U3405 (N_3405,N_2373,N_2990);
xor U3406 (N_3406,N_2609,N_2427);
and U3407 (N_3407,N_2310,N_2244);
xnor U3408 (N_3408,N_2106,N_2569);
nor U3409 (N_3409,N_2715,N_2241);
and U3410 (N_3410,N_2754,N_2893);
xor U3411 (N_3411,N_2009,N_2535);
or U3412 (N_3412,N_2015,N_2087);
or U3413 (N_3413,N_2671,N_2342);
nand U3414 (N_3414,N_2151,N_2841);
or U3415 (N_3415,N_2725,N_2647);
xnor U3416 (N_3416,N_2455,N_2827);
xor U3417 (N_3417,N_2628,N_2102);
nor U3418 (N_3418,N_2978,N_2558);
and U3419 (N_3419,N_2348,N_2030);
or U3420 (N_3420,N_2658,N_2602);
nor U3421 (N_3421,N_2467,N_2444);
nor U3422 (N_3422,N_2769,N_2676);
xor U3423 (N_3423,N_2458,N_2586);
xnor U3424 (N_3424,N_2021,N_2959);
nand U3425 (N_3425,N_2230,N_2353);
and U3426 (N_3426,N_2062,N_2965);
and U3427 (N_3427,N_2056,N_2570);
or U3428 (N_3428,N_2886,N_2065);
or U3429 (N_3429,N_2705,N_2858);
or U3430 (N_3430,N_2191,N_2749);
and U3431 (N_3431,N_2313,N_2727);
nor U3432 (N_3432,N_2328,N_2217);
and U3433 (N_3433,N_2605,N_2600);
nand U3434 (N_3434,N_2619,N_2871);
xor U3435 (N_3435,N_2290,N_2425);
xnor U3436 (N_3436,N_2014,N_2210);
or U3437 (N_3437,N_2988,N_2834);
or U3438 (N_3438,N_2470,N_2768);
and U3439 (N_3439,N_2134,N_2881);
xor U3440 (N_3440,N_2597,N_2406);
and U3441 (N_3441,N_2274,N_2221);
or U3442 (N_3442,N_2054,N_2989);
and U3443 (N_3443,N_2895,N_2897);
or U3444 (N_3444,N_2344,N_2101);
and U3445 (N_3445,N_2966,N_2610);
xnor U3446 (N_3446,N_2292,N_2688);
nand U3447 (N_3447,N_2489,N_2437);
or U3448 (N_3448,N_2235,N_2468);
nor U3449 (N_3449,N_2011,N_2320);
nand U3450 (N_3450,N_2825,N_2476);
nor U3451 (N_3451,N_2220,N_2621);
nand U3452 (N_3452,N_2148,N_2615);
nor U3453 (N_3453,N_2680,N_2577);
nor U3454 (N_3454,N_2584,N_2188);
xor U3455 (N_3455,N_2764,N_2890);
nand U3456 (N_3456,N_2048,N_2142);
xnor U3457 (N_3457,N_2446,N_2195);
xor U3458 (N_3458,N_2150,N_2276);
or U3459 (N_3459,N_2596,N_2774);
xor U3460 (N_3460,N_2670,N_2170);
and U3461 (N_3461,N_2383,N_2743);
xnor U3462 (N_3462,N_2838,N_2083);
or U3463 (N_3463,N_2542,N_2937);
nor U3464 (N_3464,N_2352,N_2206);
nand U3465 (N_3465,N_2935,N_2173);
and U3466 (N_3466,N_2611,N_2285);
xor U3467 (N_3467,N_2583,N_2533);
xor U3468 (N_3468,N_2846,N_2617);
or U3469 (N_3469,N_2736,N_2270);
nor U3470 (N_3470,N_2732,N_2187);
or U3471 (N_3471,N_2514,N_2781);
or U3472 (N_3472,N_2275,N_2139);
nor U3473 (N_3473,N_2745,N_2638);
or U3474 (N_3474,N_2852,N_2253);
and U3475 (N_3475,N_2339,N_2915);
nor U3476 (N_3476,N_2323,N_2922);
and U3477 (N_3477,N_2694,N_2145);
or U3478 (N_3478,N_2499,N_2861);
and U3479 (N_3479,N_2207,N_2379);
xor U3480 (N_3480,N_2752,N_2717);
and U3481 (N_3481,N_2559,N_2448);
xor U3482 (N_3482,N_2105,N_2410);
nor U3483 (N_3483,N_2462,N_2845);
or U3484 (N_3484,N_2793,N_2428);
or U3485 (N_3485,N_2125,N_2096);
xnor U3486 (N_3486,N_2190,N_2219);
and U3487 (N_3487,N_2487,N_2931);
or U3488 (N_3488,N_2624,N_2856);
xnor U3489 (N_3489,N_2799,N_2401);
or U3490 (N_3490,N_2598,N_2224);
nor U3491 (N_3491,N_2350,N_2471);
or U3492 (N_3492,N_2505,N_2264);
xor U3493 (N_3493,N_2855,N_2300);
xor U3494 (N_3494,N_2701,N_2911);
and U3495 (N_3495,N_2156,N_2553);
nand U3496 (N_3496,N_2050,N_2679);
nor U3497 (N_3497,N_2790,N_2973);
nand U3498 (N_3498,N_2020,N_2686);
nor U3499 (N_3499,N_2563,N_2787);
nor U3500 (N_3500,N_2319,N_2620);
xor U3501 (N_3501,N_2584,N_2233);
and U3502 (N_3502,N_2305,N_2319);
or U3503 (N_3503,N_2105,N_2405);
or U3504 (N_3504,N_2409,N_2631);
nor U3505 (N_3505,N_2130,N_2234);
or U3506 (N_3506,N_2663,N_2807);
or U3507 (N_3507,N_2177,N_2533);
nor U3508 (N_3508,N_2614,N_2977);
nand U3509 (N_3509,N_2369,N_2418);
and U3510 (N_3510,N_2621,N_2311);
nand U3511 (N_3511,N_2191,N_2473);
or U3512 (N_3512,N_2256,N_2177);
or U3513 (N_3513,N_2313,N_2722);
nor U3514 (N_3514,N_2666,N_2878);
or U3515 (N_3515,N_2478,N_2539);
nor U3516 (N_3516,N_2555,N_2647);
nand U3517 (N_3517,N_2650,N_2663);
nand U3518 (N_3518,N_2775,N_2026);
xnor U3519 (N_3519,N_2562,N_2743);
or U3520 (N_3520,N_2866,N_2968);
nor U3521 (N_3521,N_2332,N_2265);
nor U3522 (N_3522,N_2597,N_2605);
xnor U3523 (N_3523,N_2953,N_2756);
nor U3524 (N_3524,N_2919,N_2089);
xor U3525 (N_3525,N_2556,N_2126);
and U3526 (N_3526,N_2113,N_2432);
and U3527 (N_3527,N_2862,N_2034);
xor U3528 (N_3528,N_2536,N_2831);
and U3529 (N_3529,N_2878,N_2339);
xor U3530 (N_3530,N_2838,N_2618);
or U3531 (N_3531,N_2945,N_2181);
or U3532 (N_3532,N_2354,N_2370);
nand U3533 (N_3533,N_2905,N_2818);
and U3534 (N_3534,N_2625,N_2118);
xor U3535 (N_3535,N_2363,N_2782);
or U3536 (N_3536,N_2344,N_2006);
xor U3537 (N_3537,N_2263,N_2361);
nand U3538 (N_3538,N_2445,N_2819);
xor U3539 (N_3539,N_2001,N_2629);
or U3540 (N_3540,N_2976,N_2008);
or U3541 (N_3541,N_2810,N_2723);
or U3542 (N_3542,N_2727,N_2100);
and U3543 (N_3543,N_2696,N_2651);
or U3544 (N_3544,N_2552,N_2958);
or U3545 (N_3545,N_2122,N_2604);
nand U3546 (N_3546,N_2312,N_2442);
and U3547 (N_3547,N_2880,N_2200);
nand U3548 (N_3548,N_2267,N_2099);
xor U3549 (N_3549,N_2061,N_2369);
or U3550 (N_3550,N_2368,N_2474);
xnor U3551 (N_3551,N_2317,N_2990);
xnor U3552 (N_3552,N_2322,N_2593);
nand U3553 (N_3553,N_2344,N_2267);
nand U3554 (N_3554,N_2190,N_2860);
nor U3555 (N_3555,N_2443,N_2660);
xnor U3556 (N_3556,N_2995,N_2367);
nand U3557 (N_3557,N_2709,N_2113);
nand U3558 (N_3558,N_2708,N_2175);
nor U3559 (N_3559,N_2179,N_2329);
or U3560 (N_3560,N_2797,N_2260);
xnor U3561 (N_3561,N_2675,N_2936);
nand U3562 (N_3562,N_2801,N_2229);
nand U3563 (N_3563,N_2075,N_2680);
xor U3564 (N_3564,N_2583,N_2705);
xnor U3565 (N_3565,N_2533,N_2513);
nor U3566 (N_3566,N_2526,N_2857);
xnor U3567 (N_3567,N_2673,N_2939);
or U3568 (N_3568,N_2366,N_2295);
xnor U3569 (N_3569,N_2328,N_2720);
xor U3570 (N_3570,N_2279,N_2951);
and U3571 (N_3571,N_2221,N_2090);
xnor U3572 (N_3572,N_2490,N_2483);
nand U3573 (N_3573,N_2870,N_2017);
nand U3574 (N_3574,N_2842,N_2741);
nor U3575 (N_3575,N_2093,N_2088);
nor U3576 (N_3576,N_2571,N_2378);
xnor U3577 (N_3577,N_2213,N_2143);
nor U3578 (N_3578,N_2203,N_2671);
xnor U3579 (N_3579,N_2271,N_2751);
and U3580 (N_3580,N_2006,N_2934);
nor U3581 (N_3581,N_2570,N_2441);
xnor U3582 (N_3582,N_2661,N_2457);
and U3583 (N_3583,N_2408,N_2498);
and U3584 (N_3584,N_2789,N_2009);
or U3585 (N_3585,N_2482,N_2310);
nor U3586 (N_3586,N_2003,N_2940);
and U3587 (N_3587,N_2136,N_2953);
and U3588 (N_3588,N_2065,N_2865);
and U3589 (N_3589,N_2553,N_2801);
nor U3590 (N_3590,N_2300,N_2345);
or U3591 (N_3591,N_2677,N_2531);
and U3592 (N_3592,N_2638,N_2292);
xnor U3593 (N_3593,N_2457,N_2756);
xnor U3594 (N_3594,N_2655,N_2509);
nor U3595 (N_3595,N_2417,N_2969);
xor U3596 (N_3596,N_2667,N_2391);
and U3597 (N_3597,N_2026,N_2890);
nor U3598 (N_3598,N_2832,N_2133);
or U3599 (N_3599,N_2787,N_2419);
xnor U3600 (N_3600,N_2917,N_2995);
nor U3601 (N_3601,N_2971,N_2593);
nor U3602 (N_3602,N_2192,N_2122);
nor U3603 (N_3603,N_2283,N_2199);
nand U3604 (N_3604,N_2595,N_2818);
xor U3605 (N_3605,N_2074,N_2599);
and U3606 (N_3606,N_2903,N_2675);
and U3607 (N_3607,N_2390,N_2275);
nand U3608 (N_3608,N_2364,N_2932);
xnor U3609 (N_3609,N_2775,N_2821);
xor U3610 (N_3610,N_2928,N_2644);
and U3611 (N_3611,N_2871,N_2989);
nand U3612 (N_3612,N_2467,N_2923);
nor U3613 (N_3613,N_2261,N_2383);
nand U3614 (N_3614,N_2740,N_2833);
xnor U3615 (N_3615,N_2610,N_2063);
or U3616 (N_3616,N_2693,N_2339);
or U3617 (N_3617,N_2401,N_2862);
nor U3618 (N_3618,N_2624,N_2857);
and U3619 (N_3619,N_2177,N_2402);
nor U3620 (N_3620,N_2480,N_2315);
nor U3621 (N_3621,N_2241,N_2127);
xnor U3622 (N_3622,N_2826,N_2666);
nor U3623 (N_3623,N_2546,N_2958);
and U3624 (N_3624,N_2750,N_2436);
nand U3625 (N_3625,N_2244,N_2081);
nor U3626 (N_3626,N_2417,N_2838);
nor U3627 (N_3627,N_2035,N_2309);
xnor U3628 (N_3628,N_2748,N_2731);
xor U3629 (N_3629,N_2953,N_2309);
xor U3630 (N_3630,N_2713,N_2808);
xnor U3631 (N_3631,N_2955,N_2459);
or U3632 (N_3632,N_2985,N_2026);
xor U3633 (N_3633,N_2126,N_2624);
nand U3634 (N_3634,N_2268,N_2382);
or U3635 (N_3635,N_2297,N_2508);
or U3636 (N_3636,N_2696,N_2094);
nand U3637 (N_3637,N_2425,N_2012);
nand U3638 (N_3638,N_2600,N_2043);
nand U3639 (N_3639,N_2994,N_2312);
nor U3640 (N_3640,N_2339,N_2454);
xnor U3641 (N_3641,N_2694,N_2321);
nor U3642 (N_3642,N_2638,N_2511);
nor U3643 (N_3643,N_2400,N_2732);
nand U3644 (N_3644,N_2184,N_2702);
nor U3645 (N_3645,N_2815,N_2785);
nand U3646 (N_3646,N_2319,N_2663);
and U3647 (N_3647,N_2237,N_2719);
or U3648 (N_3648,N_2884,N_2621);
or U3649 (N_3649,N_2897,N_2959);
xnor U3650 (N_3650,N_2888,N_2935);
nand U3651 (N_3651,N_2437,N_2625);
or U3652 (N_3652,N_2506,N_2531);
nor U3653 (N_3653,N_2344,N_2172);
nor U3654 (N_3654,N_2798,N_2020);
nand U3655 (N_3655,N_2667,N_2062);
and U3656 (N_3656,N_2674,N_2875);
xor U3657 (N_3657,N_2268,N_2700);
nand U3658 (N_3658,N_2192,N_2532);
nor U3659 (N_3659,N_2316,N_2813);
and U3660 (N_3660,N_2043,N_2321);
xnor U3661 (N_3661,N_2611,N_2240);
xnor U3662 (N_3662,N_2019,N_2999);
and U3663 (N_3663,N_2063,N_2132);
nand U3664 (N_3664,N_2010,N_2620);
nand U3665 (N_3665,N_2706,N_2491);
or U3666 (N_3666,N_2666,N_2181);
or U3667 (N_3667,N_2648,N_2017);
or U3668 (N_3668,N_2420,N_2177);
or U3669 (N_3669,N_2813,N_2512);
nand U3670 (N_3670,N_2278,N_2515);
or U3671 (N_3671,N_2537,N_2567);
and U3672 (N_3672,N_2827,N_2721);
and U3673 (N_3673,N_2581,N_2167);
or U3674 (N_3674,N_2842,N_2117);
nand U3675 (N_3675,N_2565,N_2370);
nor U3676 (N_3676,N_2574,N_2563);
or U3677 (N_3677,N_2989,N_2785);
xnor U3678 (N_3678,N_2859,N_2602);
and U3679 (N_3679,N_2876,N_2003);
xnor U3680 (N_3680,N_2093,N_2535);
or U3681 (N_3681,N_2383,N_2806);
xor U3682 (N_3682,N_2418,N_2666);
nor U3683 (N_3683,N_2056,N_2781);
nand U3684 (N_3684,N_2253,N_2073);
nor U3685 (N_3685,N_2773,N_2782);
nor U3686 (N_3686,N_2958,N_2436);
and U3687 (N_3687,N_2960,N_2598);
xor U3688 (N_3688,N_2709,N_2779);
nand U3689 (N_3689,N_2460,N_2053);
nor U3690 (N_3690,N_2309,N_2915);
nor U3691 (N_3691,N_2388,N_2265);
nand U3692 (N_3692,N_2585,N_2127);
xor U3693 (N_3693,N_2801,N_2749);
and U3694 (N_3694,N_2730,N_2895);
xor U3695 (N_3695,N_2782,N_2804);
xnor U3696 (N_3696,N_2210,N_2007);
nand U3697 (N_3697,N_2368,N_2920);
xnor U3698 (N_3698,N_2031,N_2628);
xor U3699 (N_3699,N_2980,N_2771);
nor U3700 (N_3700,N_2800,N_2994);
and U3701 (N_3701,N_2867,N_2153);
nand U3702 (N_3702,N_2630,N_2966);
nor U3703 (N_3703,N_2391,N_2887);
or U3704 (N_3704,N_2417,N_2132);
nand U3705 (N_3705,N_2531,N_2538);
nand U3706 (N_3706,N_2358,N_2437);
nand U3707 (N_3707,N_2600,N_2144);
xnor U3708 (N_3708,N_2860,N_2606);
or U3709 (N_3709,N_2760,N_2222);
or U3710 (N_3710,N_2143,N_2295);
and U3711 (N_3711,N_2041,N_2130);
and U3712 (N_3712,N_2342,N_2164);
nor U3713 (N_3713,N_2512,N_2825);
and U3714 (N_3714,N_2855,N_2181);
nor U3715 (N_3715,N_2454,N_2474);
nor U3716 (N_3716,N_2608,N_2490);
nor U3717 (N_3717,N_2814,N_2634);
nor U3718 (N_3718,N_2541,N_2478);
nand U3719 (N_3719,N_2886,N_2552);
or U3720 (N_3720,N_2535,N_2898);
or U3721 (N_3721,N_2094,N_2510);
nor U3722 (N_3722,N_2740,N_2005);
nor U3723 (N_3723,N_2381,N_2811);
or U3724 (N_3724,N_2505,N_2219);
nand U3725 (N_3725,N_2504,N_2415);
xnor U3726 (N_3726,N_2721,N_2338);
or U3727 (N_3727,N_2439,N_2131);
xor U3728 (N_3728,N_2028,N_2526);
and U3729 (N_3729,N_2651,N_2776);
nor U3730 (N_3730,N_2339,N_2034);
nand U3731 (N_3731,N_2526,N_2333);
nor U3732 (N_3732,N_2909,N_2164);
and U3733 (N_3733,N_2934,N_2304);
and U3734 (N_3734,N_2221,N_2650);
or U3735 (N_3735,N_2120,N_2351);
and U3736 (N_3736,N_2305,N_2723);
or U3737 (N_3737,N_2403,N_2924);
or U3738 (N_3738,N_2145,N_2287);
and U3739 (N_3739,N_2753,N_2037);
nor U3740 (N_3740,N_2529,N_2110);
nor U3741 (N_3741,N_2254,N_2064);
nor U3742 (N_3742,N_2127,N_2569);
nand U3743 (N_3743,N_2187,N_2198);
xnor U3744 (N_3744,N_2676,N_2460);
and U3745 (N_3745,N_2537,N_2873);
nor U3746 (N_3746,N_2371,N_2094);
nor U3747 (N_3747,N_2127,N_2249);
xnor U3748 (N_3748,N_2336,N_2230);
and U3749 (N_3749,N_2463,N_2802);
and U3750 (N_3750,N_2676,N_2467);
and U3751 (N_3751,N_2620,N_2329);
xnor U3752 (N_3752,N_2819,N_2603);
nand U3753 (N_3753,N_2750,N_2926);
nor U3754 (N_3754,N_2165,N_2921);
xor U3755 (N_3755,N_2794,N_2746);
xor U3756 (N_3756,N_2781,N_2940);
and U3757 (N_3757,N_2257,N_2366);
nand U3758 (N_3758,N_2554,N_2638);
or U3759 (N_3759,N_2075,N_2856);
or U3760 (N_3760,N_2883,N_2363);
xor U3761 (N_3761,N_2307,N_2584);
nor U3762 (N_3762,N_2829,N_2613);
nor U3763 (N_3763,N_2120,N_2507);
or U3764 (N_3764,N_2702,N_2316);
xnor U3765 (N_3765,N_2984,N_2060);
nor U3766 (N_3766,N_2514,N_2844);
or U3767 (N_3767,N_2054,N_2954);
xnor U3768 (N_3768,N_2480,N_2566);
and U3769 (N_3769,N_2899,N_2366);
nand U3770 (N_3770,N_2621,N_2377);
or U3771 (N_3771,N_2875,N_2058);
nor U3772 (N_3772,N_2062,N_2181);
and U3773 (N_3773,N_2557,N_2384);
nand U3774 (N_3774,N_2689,N_2703);
nor U3775 (N_3775,N_2432,N_2637);
xor U3776 (N_3776,N_2284,N_2151);
nand U3777 (N_3777,N_2581,N_2550);
nor U3778 (N_3778,N_2670,N_2642);
or U3779 (N_3779,N_2062,N_2954);
nor U3780 (N_3780,N_2076,N_2108);
nor U3781 (N_3781,N_2766,N_2889);
or U3782 (N_3782,N_2008,N_2262);
or U3783 (N_3783,N_2340,N_2749);
and U3784 (N_3784,N_2689,N_2826);
xnor U3785 (N_3785,N_2892,N_2299);
nand U3786 (N_3786,N_2849,N_2573);
nor U3787 (N_3787,N_2729,N_2410);
or U3788 (N_3788,N_2883,N_2997);
xor U3789 (N_3789,N_2110,N_2015);
or U3790 (N_3790,N_2828,N_2667);
nor U3791 (N_3791,N_2474,N_2896);
nor U3792 (N_3792,N_2303,N_2467);
or U3793 (N_3793,N_2335,N_2758);
xnor U3794 (N_3794,N_2768,N_2820);
nand U3795 (N_3795,N_2255,N_2613);
and U3796 (N_3796,N_2702,N_2839);
and U3797 (N_3797,N_2426,N_2101);
and U3798 (N_3798,N_2593,N_2054);
nor U3799 (N_3799,N_2044,N_2587);
nor U3800 (N_3800,N_2868,N_2798);
or U3801 (N_3801,N_2368,N_2084);
nand U3802 (N_3802,N_2262,N_2842);
and U3803 (N_3803,N_2924,N_2184);
nand U3804 (N_3804,N_2092,N_2749);
nor U3805 (N_3805,N_2631,N_2531);
xor U3806 (N_3806,N_2387,N_2370);
and U3807 (N_3807,N_2181,N_2835);
nand U3808 (N_3808,N_2630,N_2977);
nand U3809 (N_3809,N_2849,N_2357);
and U3810 (N_3810,N_2360,N_2709);
and U3811 (N_3811,N_2589,N_2319);
and U3812 (N_3812,N_2417,N_2493);
nor U3813 (N_3813,N_2439,N_2402);
and U3814 (N_3814,N_2359,N_2767);
xor U3815 (N_3815,N_2751,N_2022);
or U3816 (N_3816,N_2566,N_2022);
and U3817 (N_3817,N_2167,N_2551);
nor U3818 (N_3818,N_2965,N_2338);
and U3819 (N_3819,N_2434,N_2712);
and U3820 (N_3820,N_2497,N_2651);
or U3821 (N_3821,N_2840,N_2347);
nand U3822 (N_3822,N_2235,N_2509);
xor U3823 (N_3823,N_2193,N_2485);
or U3824 (N_3824,N_2499,N_2015);
nor U3825 (N_3825,N_2275,N_2759);
or U3826 (N_3826,N_2094,N_2772);
xnor U3827 (N_3827,N_2473,N_2243);
or U3828 (N_3828,N_2152,N_2275);
nand U3829 (N_3829,N_2653,N_2754);
xnor U3830 (N_3830,N_2507,N_2652);
or U3831 (N_3831,N_2481,N_2971);
and U3832 (N_3832,N_2153,N_2655);
nor U3833 (N_3833,N_2737,N_2582);
nor U3834 (N_3834,N_2143,N_2715);
nand U3835 (N_3835,N_2275,N_2484);
or U3836 (N_3836,N_2012,N_2052);
nand U3837 (N_3837,N_2958,N_2058);
nor U3838 (N_3838,N_2163,N_2270);
and U3839 (N_3839,N_2925,N_2823);
xor U3840 (N_3840,N_2775,N_2877);
or U3841 (N_3841,N_2811,N_2570);
nand U3842 (N_3842,N_2887,N_2572);
nand U3843 (N_3843,N_2244,N_2495);
xnor U3844 (N_3844,N_2969,N_2024);
nor U3845 (N_3845,N_2987,N_2518);
xor U3846 (N_3846,N_2401,N_2608);
or U3847 (N_3847,N_2778,N_2872);
or U3848 (N_3848,N_2295,N_2308);
nand U3849 (N_3849,N_2815,N_2869);
nand U3850 (N_3850,N_2817,N_2606);
xor U3851 (N_3851,N_2654,N_2091);
nand U3852 (N_3852,N_2919,N_2889);
xor U3853 (N_3853,N_2668,N_2389);
nor U3854 (N_3854,N_2310,N_2137);
or U3855 (N_3855,N_2564,N_2787);
or U3856 (N_3856,N_2704,N_2858);
or U3857 (N_3857,N_2906,N_2857);
nand U3858 (N_3858,N_2334,N_2848);
nor U3859 (N_3859,N_2318,N_2419);
and U3860 (N_3860,N_2594,N_2131);
nand U3861 (N_3861,N_2043,N_2880);
nor U3862 (N_3862,N_2551,N_2807);
nor U3863 (N_3863,N_2997,N_2073);
xnor U3864 (N_3864,N_2262,N_2247);
and U3865 (N_3865,N_2047,N_2645);
and U3866 (N_3866,N_2562,N_2054);
nand U3867 (N_3867,N_2303,N_2311);
or U3868 (N_3868,N_2112,N_2710);
or U3869 (N_3869,N_2669,N_2453);
and U3870 (N_3870,N_2215,N_2642);
or U3871 (N_3871,N_2191,N_2316);
xnor U3872 (N_3872,N_2459,N_2428);
xor U3873 (N_3873,N_2949,N_2330);
or U3874 (N_3874,N_2075,N_2294);
nand U3875 (N_3875,N_2299,N_2568);
nor U3876 (N_3876,N_2807,N_2568);
xor U3877 (N_3877,N_2646,N_2641);
nand U3878 (N_3878,N_2991,N_2738);
and U3879 (N_3879,N_2393,N_2143);
nand U3880 (N_3880,N_2851,N_2824);
nor U3881 (N_3881,N_2499,N_2509);
nand U3882 (N_3882,N_2249,N_2172);
and U3883 (N_3883,N_2770,N_2262);
or U3884 (N_3884,N_2139,N_2065);
xor U3885 (N_3885,N_2979,N_2996);
or U3886 (N_3886,N_2654,N_2057);
xor U3887 (N_3887,N_2972,N_2736);
and U3888 (N_3888,N_2421,N_2866);
nand U3889 (N_3889,N_2155,N_2932);
xnor U3890 (N_3890,N_2797,N_2057);
xor U3891 (N_3891,N_2519,N_2664);
or U3892 (N_3892,N_2903,N_2051);
or U3893 (N_3893,N_2627,N_2986);
nor U3894 (N_3894,N_2855,N_2761);
xnor U3895 (N_3895,N_2678,N_2042);
nand U3896 (N_3896,N_2604,N_2244);
nor U3897 (N_3897,N_2098,N_2796);
nand U3898 (N_3898,N_2184,N_2805);
xor U3899 (N_3899,N_2542,N_2783);
nor U3900 (N_3900,N_2277,N_2993);
nand U3901 (N_3901,N_2774,N_2798);
nand U3902 (N_3902,N_2663,N_2535);
and U3903 (N_3903,N_2489,N_2311);
and U3904 (N_3904,N_2513,N_2922);
or U3905 (N_3905,N_2623,N_2475);
and U3906 (N_3906,N_2342,N_2113);
xor U3907 (N_3907,N_2772,N_2145);
nor U3908 (N_3908,N_2085,N_2904);
nor U3909 (N_3909,N_2514,N_2068);
nand U3910 (N_3910,N_2369,N_2574);
nand U3911 (N_3911,N_2868,N_2915);
or U3912 (N_3912,N_2993,N_2660);
and U3913 (N_3913,N_2589,N_2724);
and U3914 (N_3914,N_2811,N_2689);
and U3915 (N_3915,N_2693,N_2169);
nand U3916 (N_3916,N_2872,N_2666);
nor U3917 (N_3917,N_2330,N_2482);
xnor U3918 (N_3918,N_2908,N_2024);
nor U3919 (N_3919,N_2798,N_2308);
nand U3920 (N_3920,N_2614,N_2729);
or U3921 (N_3921,N_2494,N_2930);
or U3922 (N_3922,N_2456,N_2549);
or U3923 (N_3923,N_2922,N_2443);
xor U3924 (N_3924,N_2764,N_2758);
nand U3925 (N_3925,N_2399,N_2102);
xnor U3926 (N_3926,N_2258,N_2934);
xnor U3927 (N_3927,N_2085,N_2842);
xor U3928 (N_3928,N_2339,N_2925);
nand U3929 (N_3929,N_2114,N_2117);
or U3930 (N_3930,N_2770,N_2314);
xor U3931 (N_3931,N_2565,N_2555);
nor U3932 (N_3932,N_2347,N_2204);
and U3933 (N_3933,N_2712,N_2149);
nand U3934 (N_3934,N_2875,N_2331);
nand U3935 (N_3935,N_2697,N_2754);
and U3936 (N_3936,N_2073,N_2745);
xnor U3937 (N_3937,N_2280,N_2938);
nand U3938 (N_3938,N_2770,N_2463);
or U3939 (N_3939,N_2231,N_2242);
and U3940 (N_3940,N_2341,N_2914);
nor U3941 (N_3941,N_2132,N_2027);
nand U3942 (N_3942,N_2052,N_2936);
and U3943 (N_3943,N_2667,N_2642);
or U3944 (N_3944,N_2534,N_2974);
nor U3945 (N_3945,N_2676,N_2475);
and U3946 (N_3946,N_2539,N_2225);
and U3947 (N_3947,N_2859,N_2277);
and U3948 (N_3948,N_2863,N_2058);
nand U3949 (N_3949,N_2648,N_2103);
nor U3950 (N_3950,N_2663,N_2546);
and U3951 (N_3951,N_2229,N_2253);
and U3952 (N_3952,N_2398,N_2654);
nand U3953 (N_3953,N_2850,N_2801);
nand U3954 (N_3954,N_2068,N_2880);
or U3955 (N_3955,N_2779,N_2900);
nand U3956 (N_3956,N_2673,N_2545);
xor U3957 (N_3957,N_2734,N_2345);
or U3958 (N_3958,N_2945,N_2220);
nand U3959 (N_3959,N_2589,N_2198);
and U3960 (N_3960,N_2327,N_2854);
nor U3961 (N_3961,N_2878,N_2827);
or U3962 (N_3962,N_2815,N_2580);
or U3963 (N_3963,N_2607,N_2638);
nand U3964 (N_3964,N_2199,N_2117);
and U3965 (N_3965,N_2697,N_2205);
nand U3966 (N_3966,N_2040,N_2842);
nand U3967 (N_3967,N_2668,N_2579);
and U3968 (N_3968,N_2751,N_2362);
nand U3969 (N_3969,N_2900,N_2101);
xor U3970 (N_3970,N_2941,N_2875);
nor U3971 (N_3971,N_2517,N_2583);
xnor U3972 (N_3972,N_2144,N_2490);
xor U3973 (N_3973,N_2551,N_2148);
or U3974 (N_3974,N_2497,N_2639);
or U3975 (N_3975,N_2520,N_2113);
xnor U3976 (N_3976,N_2065,N_2949);
and U3977 (N_3977,N_2886,N_2391);
nand U3978 (N_3978,N_2969,N_2753);
and U3979 (N_3979,N_2420,N_2405);
nor U3980 (N_3980,N_2622,N_2621);
or U3981 (N_3981,N_2134,N_2431);
nand U3982 (N_3982,N_2240,N_2168);
nand U3983 (N_3983,N_2617,N_2053);
or U3984 (N_3984,N_2490,N_2178);
xnor U3985 (N_3985,N_2921,N_2558);
nor U3986 (N_3986,N_2666,N_2510);
nand U3987 (N_3987,N_2493,N_2678);
nand U3988 (N_3988,N_2006,N_2907);
and U3989 (N_3989,N_2297,N_2282);
nor U3990 (N_3990,N_2180,N_2705);
and U3991 (N_3991,N_2068,N_2380);
xor U3992 (N_3992,N_2805,N_2161);
xnor U3993 (N_3993,N_2565,N_2417);
xnor U3994 (N_3994,N_2829,N_2249);
xor U3995 (N_3995,N_2022,N_2902);
and U3996 (N_3996,N_2583,N_2278);
and U3997 (N_3997,N_2835,N_2436);
xor U3998 (N_3998,N_2706,N_2819);
xor U3999 (N_3999,N_2574,N_2899);
nor U4000 (N_4000,N_3920,N_3584);
nor U4001 (N_4001,N_3376,N_3131);
and U4002 (N_4002,N_3554,N_3424);
nand U4003 (N_4003,N_3243,N_3578);
nand U4004 (N_4004,N_3629,N_3053);
xor U4005 (N_4005,N_3322,N_3445);
and U4006 (N_4006,N_3603,N_3472);
nor U4007 (N_4007,N_3992,N_3836);
and U4008 (N_4008,N_3972,N_3655);
or U4009 (N_4009,N_3160,N_3174);
and U4010 (N_4010,N_3264,N_3870);
nand U4011 (N_4011,N_3503,N_3499);
nand U4012 (N_4012,N_3446,N_3394);
or U4013 (N_4013,N_3268,N_3671);
or U4014 (N_4014,N_3813,N_3539);
nor U4015 (N_4015,N_3095,N_3052);
nor U4016 (N_4016,N_3789,N_3207);
xor U4017 (N_4017,N_3638,N_3215);
or U4018 (N_4018,N_3777,N_3509);
or U4019 (N_4019,N_3974,N_3469);
nand U4020 (N_4020,N_3919,N_3019);
and U4021 (N_4021,N_3352,N_3328);
or U4022 (N_4022,N_3871,N_3916);
or U4023 (N_4023,N_3959,N_3627);
xnor U4024 (N_4024,N_3912,N_3094);
and U4025 (N_4025,N_3193,N_3156);
and U4026 (N_4026,N_3184,N_3764);
nor U4027 (N_4027,N_3489,N_3716);
and U4028 (N_4028,N_3295,N_3534);
nand U4029 (N_4029,N_3712,N_3928);
xor U4030 (N_4030,N_3946,N_3435);
and U4031 (N_4031,N_3548,N_3206);
or U4032 (N_4032,N_3795,N_3700);
xnor U4033 (N_4033,N_3456,N_3988);
or U4034 (N_4034,N_3382,N_3632);
and U4035 (N_4035,N_3581,N_3693);
xor U4036 (N_4036,N_3375,N_3484);
nand U4037 (N_4037,N_3252,N_3560);
xnor U4038 (N_4038,N_3758,N_3579);
nand U4039 (N_4039,N_3396,N_3099);
nand U4040 (N_4040,N_3075,N_3773);
nor U4041 (N_4041,N_3146,N_3824);
nor U4042 (N_4042,N_3312,N_3267);
nor U4043 (N_4043,N_3620,N_3236);
and U4044 (N_4044,N_3601,N_3894);
or U4045 (N_4045,N_3676,N_3705);
xor U4046 (N_4046,N_3205,N_3204);
nand U4047 (N_4047,N_3513,N_3426);
nand U4048 (N_4048,N_3029,N_3355);
xor U4049 (N_4049,N_3540,N_3185);
nor U4050 (N_4050,N_3796,N_3129);
nor U4051 (N_4051,N_3544,N_3457);
and U4052 (N_4052,N_3470,N_3161);
xnor U4053 (N_4053,N_3454,N_3985);
xnor U4054 (N_4054,N_3944,N_3187);
nand U4055 (N_4055,N_3464,N_3440);
or U4056 (N_4056,N_3820,N_3171);
or U4057 (N_4057,N_3324,N_3719);
and U4058 (N_4058,N_3128,N_3844);
nand U4059 (N_4059,N_3222,N_3877);
nand U4060 (N_4060,N_3388,N_3049);
nor U4061 (N_4061,N_3882,N_3884);
nor U4062 (N_4062,N_3814,N_3754);
or U4063 (N_4063,N_3904,N_3090);
nor U4064 (N_4064,N_3197,N_3771);
xor U4065 (N_4065,N_3315,N_3317);
and U4066 (N_4066,N_3432,N_3888);
and U4067 (N_4067,N_3084,N_3559);
and U4068 (N_4068,N_3865,N_3311);
and U4069 (N_4069,N_3833,N_3731);
or U4070 (N_4070,N_3044,N_3073);
nor U4071 (N_4071,N_3014,N_3990);
and U4072 (N_4072,N_3144,N_3872);
nand U4073 (N_4073,N_3168,N_3492);
nor U4074 (N_4074,N_3176,N_3493);
and U4075 (N_4075,N_3209,N_3338);
xnor U4076 (N_4076,N_3610,N_3588);
xnor U4077 (N_4077,N_3428,N_3068);
xor U4078 (N_4078,N_3203,N_3093);
xor U4079 (N_4079,N_3361,N_3648);
nand U4080 (N_4080,N_3483,N_3346);
nor U4081 (N_4081,N_3092,N_3859);
nand U4082 (N_4082,N_3728,N_3466);
xor U4083 (N_4083,N_3337,N_3862);
or U4084 (N_4084,N_3040,N_3098);
xnor U4085 (N_4085,N_3518,N_3977);
nor U4086 (N_4086,N_3109,N_3002);
and U4087 (N_4087,N_3310,N_3351);
or U4088 (N_4088,N_3682,N_3050);
or U4089 (N_4089,N_3656,N_3890);
nand U4090 (N_4090,N_3221,N_3138);
xor U4091 (N_4091,N_3347,N_3213);
and U4092 (N_4092,N_3506,N_3850);
nor U4093 (N_4093,N_3231,N_3158);
nor U4094 (N_4094,N_3232,N_3962);
xnor U4095 (N_4095,N_3122,N_3399);
xor U4096 (N_4096,N_3886,N_3551);
nand U4097 (N_4097,N_3153,N_3798);
nand U4098 (N_4098,N_3443,N_3327);
or U4099 (N_4099,N_3032,N_3063);
and U4100 (N_4100,N_3653,N_3616);
or U4101 (N_4101,N_3590,N_3699);
and U4102 (N_4102,N_3415,N_3255);
nand U4103 (N_4103,N_3812,N_3697);
and U4104 (N_4104,N_3150,N_3298);
and U4105 (N_4105,N_3574,N_3439);
nand U4106 (N_4106,N_3909,N_3172);
or U4107 (N_4107,N_3940,N_3949);
or U4108 (N_4108,N_3247,N_3971);
nor U4109 (N_4109,N_3634,N_3757);
nor U4110 (N_4110,N_3323,N_3933);
and U4111 (N_4111,N_3643,N_3058);
or U4112 (N_4112,N_3026,N_3490);
and U4113 (N_4113,N_3975,N_3937);
or U4114 (N_4114,N_3856,N_3104);
and U4115 (N_4115,N_3594,N_3725);
or U4116 (N_4116,N_3462,N_3720);
or U4117 (N_4117,N_3956,N_3006);
and U4118 (N_4118,N_3300,N_3386);
nand U4119 (N_4119,N_3233,N_3167);
xor U4120 (N_4120,N_3288,N_3597);
and U4121 (N_4121,N_3143,N_3111);
and U4122 (N_4122,N_3746,N_3216);
and U4123 (N_4123,N_3430,N_3807);
nor U4124 (N_4124,N_3639,N_3163);
or U4125 (N_4125,N_3285,N_3645);
xnor U4126 (N_4126,N_3733,N_3786);
nand U4127 (N_4127,N_3291,N_3970);
nor U4128 (N_4128,N_3722,N_3091);
and U4129 (N_4129,N_3265,N_3692);
nor U4130 (N_4130,N_3417,N_3599);
and U4131 (N_4131,N_3917,N_3076);
nor U4132 (N_4132,N_3628,N_3984);
or U4133 (N_4133,N_3874,N_3114);
or U4134 (N_4134,N_3250,N_3748);
or U4135 (N_4135,N_3377,N_3791);
and U4136 (N_4136,N_3670,N_3476);
and U4137 (N_4137,N_3561,N_3309);
nand U4138 (N_4138,N_3303,N_3902);
and U4139 (N_4139,N_3071,N_3826);
or U4140 (N_4140,N_3704,N_3792);
nor U4141 (N_4141,N_3418,N_3926);
xor U4142 (N_4142,N_3522,N_3938);
nor U4143 (N_4143,N_3048,N_3967);
and U4144 (N_4144,N_3305,N_3065);
or U4145 (N_4145,N_3686,N_3819);
nor U4146 (N_4146,N_3169,N_3625);
and U4147 (N_4147,N_3296,N_3393);
xnor U4148 (N_4148,N_3431,N_3342);
xor U4149 (N_4149,N_3955,N_3212);
or U4150 (N_4150,N_3107,N_3448);
nor U4151 (N_4151,N_3465,N_3307);
nor U4152 (N_4152,N_3525,N_3681);
nand U4153 (N_4153,N_3897,N_3553);
nor U4154 (N_4154,N_3593,N_3838);
or U4155 (N_4155,N_3289,N_3196);
xor U4156 (N_4156,N_3766,N_3330);
and U4157 (N_4157,N_3649,N_3921);
nand U4158 (N_4158,N_3242,N_3459);
nor U4159 (N_4159,N_3367,N_3414);
xnor U4160 (N_4160,N_3982,N_3781);
xor U4161 (N_4161,N_3117,N_3318);
xor U4162 (N_4162,N_3517,N_3732);
nand U4163 (N_4163,N_3069,N_3140);
nand U4164 (N_4164,N_3793,N_3701);
nand U4165 (N_4165,N_3478,N_3673);
and U4166 (N_4166,N_3239,N_3570);
nand U4167 (N_4167,N_3360,N_3966);
nand U4168 (N_4168,N_3861,N_3316);
or U4169 (N_4169,N_3384,N_3362);
nor U4170 (N_4170,N_3060,N_3190);
xor U4171 (N_4171,N_3979,N_3723);
nand U4172 (N_4172,N_3467,N_3282);
and U4173 (N_4173,N_3321,N_3392);
or U4174 (N_4174,N_3302,N_3219);
nand U4175 (N_4175,N_3875,N_3945);
nand U4176 (N_4176,N_3519,N_3986);
nand U4177 (N_4177,N_3779,N_3078);
nor U4178 (N_4178,N_3918,N_3381);
nand U4179 (N_4179,N_3501,N_3112);
or U4180 (N_4180,N_3591,N_3261);
xor U4181 (N_4181,N_3911,N_3101);
or U4182 (N_4182,N_3567,N_3314);
and U4183 (N_4183,N_3313,N_3121);
nor U4184 (N_4184,N_3441,N_3349);
or U4185 (N_4185,N_3976,N_3743);
or U4186 (N_4186,N_3741,N_3370);
or U4187 (N_4187,N_3334,N_3198);
and U4188 (N_4188,N_3429,N_3925);
xor U4189 (N_4189,N_3915,N_3552);
and U4190 (N_4190,N_3669,N_3595);
xor U4191 (N_4191,N_3989,N_3016);
or U4192 (N_4192,N_3684,N_3840);
nor U4193 (N_4193,N_3822,N_3834);
or U4194 (N_4194,N_3279,N_3283);
nand U4195 (N_4195,N_3088,N_3849);
xnor U4196 (N_4196,N_3654,N_3046);
nor U4197 (N_4197,N_3652,N_3287);
nor U4198 (N_4198,N_3433,N_3054);
and U4199 (N_4199,N_3450,N_3857);
xor U4200 (N_4200,N_3170,N_3718);
xor U4201 (N_4201,N_3508,N_3404);
and U4202 (N_4202,N_3502,N_3041);
nand U4203 (N_4203,N_3278,N_3745);
and U4204 (N_4204,N_3566,N_3408);
nor U4205 (N_4205,N_3677,N_3948);
nor U4206 (N_4206,N_3858,N_3775);
nand U4207 (N_4207,N_3740,N_3043);
nor U4208 (N_4208,N_3407,N_3229);
xor U4209 (N_4209,N_3706,N_3854);
xnor U4210 (N_4210,N_3621,N_3262);
nand U4211 (N_4211,N_3931,N_3123);
and U4212 (N_4212,N_3973,N_3934);
or U4213 (N_4213,N_3017,N_3660);
nand U4214 (N_4214,N_3770,N_3301);
or U4215 (N_4215,N_3617,N_3935);
and U4216 (N_4216,N_3225,N_3175);
nand U4217 (N_4217,N_3390,N_3864);
and U4218 (N_4218,N_3411,N_3378);
or U4219 (N_4219,N_3800,N_3217);
and U4220 (N_4220,N_3531,N_3344);
xnor U4221 (N_4221,N_3406,N_3710);
or U4222 (N_4222,N_3753,N_3845);
nor U4223 (N_4223,N_3113,N_3269);
and U4224 (N_4224,N_3855,N_3332);
or U4225 (N_4225,N_3208,N_3274);
nor U4226 (N_4226,N_3852,N_3115);
or U4227 (N_4227,N_3577,N_3964);
and U4228 (N_4228,N_3007,N_3943);
or U4229 (N_4229,N_3319,N_3905);
xnor U4230 (N_4230,N_3846,N_3132);
xor U4231 (N_4231,N_3817,N_3734);
nand U4232 (N_4232,N_3618,N_3794);
xnor U4233 (N_4233,N_3823,N_3930);
nor U4234 (N_4234,N_3997,N_3797);
nand U4235 (N_4235,N_3801,N_3133);
and U4236 (N_4236,N_3066,N_3364);
and U4237 (N_4237,N_3333,N_3624);
nand U4238 (N_4238,N_3141,N_3707);
or U4239 (N_4239,N_3083,N_3783);
nand U4240 (N_4240,N_3297,N_3177);
or U4241 (N_4241,N_3102,N_3987);
nand U4242 (N_4242,N_3607,N_3662);
xor U4243 (N_4243,N_3932,N_3125);
nand U4244 (N_4244,N_3020,N_3556);
nor U4245 (N_4245,N_3154,N_3039);
nand U4246 (N_4246,N_3837,N_3358);
nor U4247 (N_4247,N_3164,N_3737);
or U4248 (N_4248,N_3537,N_3391);
nand U4249 (N_4249,N_3735,N_3887);
xnor U4250 (N_4250,N_3541,N_3202);
and U4251 (N_4251,N_3496,N_3760);
or U4252 (N_4252,N_3024,N_3809);
and U4253 (N_4253,N_3263,N_3922);
xor U4254 (N_4254,N_3952,N_3211);
nand U4255 (N_4255,N_3602,N_3558);
nor U4256 (N_4256,N_3866,N_3194);
xor U4257 (N_4257,N_3139,N_3679);
nand U4258 (N_4258,N_3788,N_3110);
nor U4259 (N_4259,N_3438,N_3500);
xor U4260 (N_4260,N_3401,N_3336);
nor U4261 (N_4261,N_3339,N_3804);
or U4262 (N_4262,N_3914,N_3542);
nor U4263 (N_4263,N_3224,N_3226);
nor U4264 (N_4264,N_3120,N_3750);
or U4265 (N_4265,N_3097,N_3863);
nor U4266 (N_4266,N_3460,N_3293);
nor U4267 (N_4267,N_3658,N_3960);
and U4268 (N_4268,N_3021,N_3523);
and U4269 (N_4269,N_3709,N_3957);
and U4270 (N_4270,N_3582,N_3507);
nand U4271 (N_4271,N_3425,N_3475);
and U4272 (N_4272,N_3815,N_3995);
nor U4273 (N_4273,N_3162,N_3062);
and U4274 (N_4274,N_3546,N_3389);
or U4275 (N_4275,N_3306,N_3061);
xor U4276 (N_4276,N_3479,N_3397);
xor U4277 (N_4277,N_3768,N_3596);
nand U4278 (N_4278,N_3480,N_3035);
xnor U4279 (N_4279,N_3776,N_3583);
or U4280 (N_4280,N_3331,N_3220);
nor U4281 (N_4281,N_3821,N_3335);
nor U4282 (N_4282,N_3726,N_3580);
xor U4283 (N_4283,N_3074,N_3135);
nand U4284 (N_4284,N_3227,N_3811);
or U4285 (N_4285,N_3562,N_3623);
nand U4286 (N_4286,N_3070,N_3468);
xor U4287 (N_4287,N_3257,N_3345);
nor U4288 (N_4288,N_3667,N_3182);
and U4289 (N_4289,N_3589,N_3555);
and U4290 (N_4290,N_3936,N_3808);
nand U4291 (N_4291,N_3412,N_3774);
nand U4292 (N_4292,N_3630,N_3545);
nor U4293 (N_4293,N_3751,N_3762);
xnor U4294 (N_4294,N_3080,N_3714);
or U4295 (N_4295,N_3640,N_3563);
nor U4296 (N_4296,N_3031,N_3395);
nand U4297 (N_4297,N_3529,N_3449);
nor U4298 (N_4298,N_3354,N_3575);
xnor U4299 (N_4299,N_3843,N_3147);
nand U4300 (N_4300,N_3965,N_3320);
nor U4301 (N_4301,N_3516,N_3214);
nand U4302 (N_4302,N_3900,N_3482);
or U4303 (N_4303,N_3037,N_3159);
nand U4304 (N_4304,N_3568,N_3802);
or U4305 (N_4305,N_3442,N_3892);
nand U4306 (N_4306,N_3341,N_3308);
and U4307 (N_4307,N_3947,N_3486);
or U4308 (N_4308,N_3708,N_3249);
nor U4309 (N_4309,N_3927,N_3436);
nand U4310 (N_4310,N_3663,N_3281);
nand U4311 (N_4311,N_3096,N_3969);
and U4312 (N_4312,N_3034,N_3906);
xor U4313 (N_4313,N_3234,N_3767);
nand U4314 (N_4314,N_3271,N_3659);
nand U4315 (N_4315,N_3520,N_3505);
nor U4316 (N_4316,N_3825,N_3359);
nor U4317 (N_4317,N_3665,N_3235);
xnor U4318 (N_4318,N_3343,N_3611);
xor U4319 (N_4319,N_3514,N_3572);
nor U4320 (N_4320,N_3576,N_3165);
nand U4321 (N_4321,N_3526,N_3810);
or U4322 (N_4322,N_3089,N_3118);
nand U4323 (N_4323,N_3521,N_3294);
nand U4324 (N_4324,N_3761,N_3538);
nor U4325 (N_4325,N_3270,N_3218);
nand U4326 (N_4326,N_3157,N_3047);
nor U4327 (N_4327,N_3385,N_3941);
nor U4328 (N_4328,N_3055,N_3244);
or U4329 (N_4329,N_3286,N_3416);
or U4330 (N_4330,N_3675,N_3778);
xor U4331 (N_4331,N_3260,N_3251);
and U4332 (N_4332,N_3685,N_3999);
and U4333 (N_4333,N_3179,N_3253);
and U4334 (N_4334,N_3571,N_3487);
or U4335 (N_4335,N_3880,N_3961);
nor U4336 (N_4336,N_3280,N_3241);
and U4337 (N_4337,N_3790,N_3420);
nor U4338 (N_4338,N_3528,N_3883);
xor U4339 (N_4339,N_3827,N_3835);
nand U4340 (N_4340,N_3923,N_3678);
and U4341 (N_4341,N_3369,N_3057);
nor U4342 (N_4342,N_3968,N_3413);
or U4343 (N_4343,N_3240,N_3363);
and U4344 (N_4344,N_3642,N_3042);
nor U4345 (N_4345,N_3830,N_3124);
or U4346 (N_4346,N_3258,N_3186);
xor U4347 (N_4347,N_3742,N_3248);
nor U4348 (N_4348,N_3759,N_3873);
nor U4349 (N_4349,N_3045,N_3009);
or U4350 (N_4350,N_3142,N_3011);
and U4351 (N_4351,N_3030,N_3954);
nand U4352 (N_4352,N_3325,N_3005);
xor U4353 (N_4353,N_3876,N_3166);
and U4354 (N_4354,N_3899,N_3451);
xnor U4355 (N_4355,N_3847,N_3498);
nand U4356 (N_4356,N_3893,N_3896);
nand U4357 (N_4357,N_3366,N_3497);
xnor U4358 (N_4358,N_3481,N_3149);
or U4359 (N_4359,N_3398,N_3477);
nand U4360 (N_4360,N_3908,N_3806);
nand U4361 (N_4361,N_3405,N_3765);
nand U4362 (N_4362,N_3299,N_3950);
xor U4363 (N_4363,N_3881,N_3181);
nor U4364 (N_4364,N_3474,N_3188);
nand U4365 (N_4365,N_3891,N_3715);
nand U4366 (N_4366,N_3004,N_3848);
nand U4367 (N_4367,N_3694,N_3939);
nor U4368 (N_4368,N_3427,N_3619);
and U4369 (N_4369,N_3744,N_3785);
nand U4370 (N_4370,N_3422,N_3012);
xnor U4371 (N_4371,N_3458,N_3828);
nor U4372 (N_4372,N_3901,N_3885);
nor U4373 (N_4373,N_3993,N_3860);
xnor U4374 (N_4374,N_3237,N_3079);
xnor U4375 (N_4375,N_3711,N_3116);
nor U4376 (N_4376,N_3419,N_3245);
nand U4377 (N_4377,N_3023,N_3015);
xnor U4378 (N_4378,N_3755,N_3434);
xor U4379 (N_4379,N_3829,N_3895);
nor U4380 (N_4380,N_3151,N_3637);
and U4381 (N_4381,N_3189,N_3134);
or U4382 (N_4382,N_3609,N_3612);
and U4383 (N_4383,N_3680,N_3532);
xor U4384 (N_4384,N_3647,N_3372);
and U4385 (N_4385,N_3668,N_3028);
nor U4386 (N_4386,N_3749,N_3200);
nand U4387 (N_4387,N_3739,N_3410);
or U4388 (N_4388,N_3087,N_3600);
or U4389 (N_4389,N_3447,N_3958);
or U4390 (N_4390,N_3365,N_3695);
nand U4391 (N_4391,N_3547,N_3510);
nor U4392 (N_4392,N_3782,N_3353);
xor U4393 (N_4393,N_3929,N_3228);
xor U4394 (N_4394,N_3841,N_3137);
nand U4395 (N_4395,N_3878,N_3674);
xor U4396 (N_4396,N_3136,N_3085);
and U4397 (N_4397,N_3666,N_3025);
or U4398 (N_4398,N_3266,N_3787);
nand U4399 (N_4399,N_3702,N_3996);
xor U4400 (N_4400,N_3738,N_3077);
or U4401 (N_4401,N_3178,N_3191);
nor U4402 (N_4402,N_3494,N_3803);
nand U4403 (N_4403,N_3195,N_3530);
xnor U4404 (N_4404,N_3400,N_3867);
or U4405 (N_4405,N_3003,N_3027);
nor U4406 (N_4406,N_3799,N_3290);
or U4407 (N_4407,N_3515,N_3409);
nand U4408 (N_4408,N_3615,N_3452);
and U4409 (N_4409,N_3832,N_3910);
and U4410 (N_4410,N_3557,N_3511);
and U4411 (N_4411,N_3805,N_3535);
or U4412 (N_4412,N_3403,N_3585);
xnor U4413 (N_4413,N_3898,N_3256);
or U4414 (N_4414,N_3155,N_3879);
and U4415 (N_4415,N_3380,N_3246);
nand U4416 (N_4416,N_3672,N_3661);
nor U4417 (N_4417,N_3086,N_3851);
nand U4418 (N_4418,N_3622,N_3038);
xnor U4419 (N_4419,N_3357,N_3924);
nor U4420 (N_4420,N_3326,N_3373);
and U4421 (N_4421,N_3721,N_3350);
and U4422 (N_4422,N_3127,N_3978);
xnor U4423 (N_4423,N_3081,N_3994);
or U4424 (N_4424,N_3356,N_3276);
xnor U4425 (N_4425,N_3644,N_3461);
and U4426 (N_4426,N_3402,N_3687);
or U4427 (N_4427,N_3942,N_3569);
nor U4428 (N_4428,N_3690,N_3903);
or U4429 (N_4429,N_3842,N_3371);
nand U4430 (N_4430,N_3277,N_3717);
nor U4431 (N_4431,N_3379,N_3230);
nor U4432 (N_4432,N_3223,N_3183);
xnor U4433 (N_4433,N_3512,N_3018);
xnor U4434 (N_4434,N_3238,N_3100);
xnor U4435 (N_4435,N_3724,N_3980);
nand U4436 (N_4436,N_3747,N_3536);
xor U4437 (N_4437,N_3549,N_3889);
nor U4438 (N_4438,N_3056,N_3008);
nand U4439 (N_4439,N_3059,N_3051);
or U4440 (N_4440,N_3631,N_3573);
nand U4441 (N_4441,N_3636,N_3504);
xnor U4442 (N_4442,N_3907,N_3106);
or U4443 (N_4443,N_3592,N_3033);
xnor U4444 (N_4444,N_3272,N_3818);
and U4445 (N_4445,N_3471,N_3780);
nor U4446 (N_4446,N_3453,N_3072);
and U4447 (N_4447,N_3651,N_3869);
and U4448 (N_4448,N_3145,N_3565);
nor U4449 (N_4449,N_3598,N_3108);
or U4450 (N_4450,N_3613,N_3606);
or U4451 (N_4451,N_3586,N_3951);
xor U4452 (N_4452,N_3983,N_3488);
xor U4453 (N_4453,N_3374,N_3953);
nand U4454 (N_4454,N_3152,N_3688);
nand U4455 (N_4455,N_3772,N_3463);
and U4456 (N_4456,N_3963,N_3304);
nor U4457 (N_4457,N_3524,N_3199);
or U4458 (N_4458,N_3543,N_3000);
nor U4459 (N_4459,N_3608,N_3981);
and U4460 (N_4460,N_3657,N_3119);
nor U4461 (N_4461,N_3641,N_3550);
or U4462 (N_4462,N_3485,N_3683);
nand U4463 (N_4463,N_3853,N_3756);
xor U4464 (N_4464,N_3495,N_3650);
xor U4465 (N_4465,N_3180,N_3275);
xnor U4466 (N_4466,N_3527,N_3421);
xnor U4467 (N_4467,N_3664,N_3437);
nor U4468 (N_4468,N_3013,N_3703);
xor U4469 (N_4469,N_3698,N_3604);
nand U4470 (N_4470,N_3130,N_3067);
and U4471 (N_4471,N_3292,N_3064);
nor U4472 (N_4472,N_3691,N_3763);
nand U4473 (N_4473,N_3689,N_3368);
and U4474 (N_4474,N_3729,N_3036);
or U4475 (N_4475,N_3444,N_3816);
nor U4476 (N_4476,N_3126,N_3752);
and U4477 (N_4477,N_3491,N_3103);
nand U4478 (N_4478,N_3769,N_3201);
nand U4479 (N_4479,N_3991,N_3614);
or U4480 (N_4480,N_3340,N_3148);
nand U4481 (N_4481,N_3210,N_3273);
or U4482 (N_4482,N_3831,N_3254);
and U4483 (N_4483,N_3423,N_3192);
xnor U4484 (N_4484,N_3913,N_3839);
and U4485 (N_4485,N_3259,N_3082);
or U4486 (N_4486,N_3284,N_3646);
nor U4487 (N_4487,N_3998,N_3784);
nand U4488 (N_4488,N_3605,N_3635);
nand U4489 (N_4489,N_3387,N_3383);
nand U4490 (N_4490,N_3868,N_3473);
or U4491 (N_4491,N_3730,N_3105);
and U4492 (N_4492,N_3001,N_3022);
nor U4493 (N_4493,N_3010,N_3736);
and U4494 (N_4494,N_3696,N_3626);
nor U4495 (N_4495,N_3633,N_3713);
xor U4496 (N_4496,N_3329,N_3533);
and U4497 (N_4497,N_3587,N_3173);
and U4498 (N_4498,N_3348,N_3727);
xor U4499 (N_4499,N_3455,N_3564);
nor U4500 (N_4500,N_3107,N_3266);
xor U4501 (N_4501,N_3582,N_3493);
nand U4502 (N_4502,N_3369,N_3581);
or U4503 (N_4503,N_3908,N_3549);
and U4504 (N_4504,N_3941,N_3485);
nand U4505 (N_4505,N_3077,N_3252);
xor U4506 (N_4506,N_3153,N_3840);
nand U4507 (N_4507,N_3732,N_3917);
or U4508 (N_4508,N_3525,N_3612);
nand U4509 (N_4509,N_3033,N_3243);
nor U4510 (N_4510,N_3032,N_3172);
nor U4511 (N_4511,N_3621,N_3715);
nand U4512 (N_4512,N_3102,N_3048);
and U4513 (N_4513,N_3524,N_3846);
and U4514 (N_4514,N_3549,N_3594);
or U4515 (N_4515,N_3743,N_3654);
nor U4516 (N_4516,N_3824,N_3295);
and U4517 (N_4517,N_3079,N_3199);
nor U4518 (N_4518,N_3281,N_3589);
xor U4519 (N_4519,N_3489,N_3824);
and U4520 (N_4520,N_3184,N_3386);
nor U4521 (N_4521,N_3221,N_3993);
or U4522 (N_4522,N_3477,N_3375);
xnor U4523 (N_4523,N_3700,N_3408);
or U4524 (N_4524,N_3290,N_3311);
xnor U4525 (N_4525,N_3382,N_3666);
or U4526 (N_4526,N_3440,N_3073);
nand U4527 (N_4527,N_3992,N_3710);
or U4528 (N_4528,N_3666,N_3437);
xor U4529 (N_4529,N_3209,N_3213);
and U4530 (N_4530,N_3774,N_3852);
or U4531 (N_4531,N_3713,N_3238);
or U4532 (N_4532,N_3330,N_3353);
nor U4533 (N_4533,N_3290,N_3796);
nor U4534 (N_4534,N_3983,N_3914);
or U4535 (N_4535,N_3683,N_3990);
or U4536 (N_4536,N_3444,N_3615);
nand U4537 (N_4537,N_3116,N_3243);
nor U4538 (N_4538,N_3070,N_3205);
xor U4539 (N_4539,N_3300,N_3036);
nand U4540 (N_4540,N_3914,N_3271);
nand U4541 (N_4541,N_3074,N_3408);
xnor U4542 (N_4542,N_3711,N_3644);
xor U4543 (N_4543,N_3133,N_3917);
xor U4544 (N_4544,N_3094,N_3776);
xnor U4545 (N_4545,N_3581,N_3848);
nor U4546 (N_4546,N_3824,N_3672);
nand U4547 (N_4547,N_3594,N_3174);
and U4548 (N_4548,N_3325,N_3804);
nor U4549 (N_4549,N_3184,N_3852);
nand U4550 (N_4550,N_3878,N_3469);
or U4551 (N_4551,N_3877,N_3765);
xor U4552 (N_4552,N_3563,N_3432);
and U4553 (N_4553,N_3995,N_3689);
and U4554 (N_4554,N_3844,N_3412);
and U4555 (N_4555,N_3775,N_3813);
xor U4556 (N_4556,N_3567,N_3473);
nand U4557 (N_4557,N_3538,N_3167);
or U4558 (N_4558,N_3907,N_3867);
or U4559 (N_4559,N_3740,N_3752);
nand U4560 (N_4560,N_3439,N_3588);
nand U4561 (N_4561,N_3453,N_3987);
and U4562 (N_4562,N_3714,N_3973);
and U4563 (N_4563,N_3449,N_3870);
or U4564 (N_4564,N_3716,N_3922);
and U4565 (N_4565,N_3269,N_3910);
nor U4566 (N_4566,N_3639,N_3875);
xnor U4567 (N_4567,N_3134,N_3769);
xnor U4568 (N_4568,N_3190,N_3603);
xor U4569 (N_4569,N_3240,N_3794);
nor U4570 (N_4570,N_3406,N_3682);
nor U4571 (N_4571,N_3567,N_3041);
nand U4572 (N_4572,N_3813,N_3245);
or U4573 (N_4573,N_3832,N_3875);
or U4574 (N_4574,N_3396,N_3579);
nand U4575 (N_4575,N_3004,N_3226);
and U4576 (N_4576,N_3601,N_3693);
or U4577 (N_4577,N_3497,N_3077);
and U4578 (N_4578,N_3589,N_3244);
nor U4579 (N_4579,N_3070,N_3190);
nor U4580 (N_4580,N_3842,N_3376);
nor U4581 (N_4581,N_3606,N_3966);
nor U4582 (N_4582,N_3295,N_3982);
xnor U4583 (N_4583,N_3292,N_3132);
nand U4584 (N_4584,N_3284,N_3702);
or U4585 (N_4585,N_3153,N_3902);
or U4586 (N_4586,N_3976,N_3856);
nand U4587 (N_4587,N_3238,N_3533);
xnor U4588 (N_4588,N_3457,N_3261);
nand U4589 (N_4589,N_3997,N_3734);
and U4590 (N_4590,N_3050,N_3501);
xnor U4591 (N_4591,N_3034,N_3863);
or U4592 (N_4592,N_3379,N_3072);
nor U4593 (N_4593,N_3760,N_3157);
nand U4594 (N_4594,N_3150,N_3514);
xnor U4595 (N_4595,N_3060,N_3733);
nor U4596 (N_4596,N_3259,N_3423);
nor U4597 (N_4597,N_3013,N_3745);
nor U4598 (N_4598,N_3564,N_3947);
nand U4599 (N_4599,N_3209,N_3265);
or U4600 (N_4600,N_3352,N_3313);
nor U4601 (N_4601,N_3726,N_3416);
nor U4602 (N_4602,N_3552,N_3398);
and U4603 (N_4603,N_3641,N_3486);
or U4604 (N_4604,N_3541,N_3890);
xor U4605 (N_4605,N_3285,N_3790);
xor U4606 (N_4606,N_3527,N_3314);
xnor U4607 (N_4607,N_3742,N_3962);
xnor U4608 (N_4608,N_3277,N_3544);
nand U4609 (N_4609,N_3095,N_3799);
and U4610 (N_4610,N_3137,N_3919);
nand U4611 (N_4611,N_3767,N_3290);
xnor U4612 (N_4612,N_3929,N_3687);
xnor U4613 (N_4613,N_3723,N_3471);
or U4614 (N_4614,N_3138,N_3385);
or U4615 (N_4615,N_3467,N_3975);
and U4616 (N_4616,N_3761,N_3027);
and U4617 (N_4617,N_3665,N_3205);
and U4618 (N_4618,N_3431,N_3840);
xnor U4619 (N_4619,N_3548,N_3565);
nor U4620 (N_4620,N_3999,N_3092);
or U4621 (N_4621,N_3093,N_3841);
nand U4622 (N_4622,N_3422,N_3621);
or U4623 (N_4623,N_3282,N_3560);
or U4624 (N_4624,N_3393,N_3333);
or U4625 (N_4625,N_3294,N_3168);
and U4626 (N_4626,N_3390,N_3587);
nand U4627 (N_4627,N_3320,N_3114);
and U4628 (N_4628,N_3204,N_3998);
nor U4629 (N_4629,N_3434,N_3885);
xor U4630 (N_4630,N_3749,N_3881);
and U4631 (N_4631,N_3773,N_3740);
nor U4632 (N_4632,N_3652,N_3184);
xnor U4633 (N_4633,N_3190,N_3314);
xnor U4634 (N_4634,N_3101,N_3316);
xnor U4635 (N_4635,N_3349,N_3567);
nor U4636 (N_4636,N_3554,N_3639);
xnor U4637 (N_4637,N_3024,N_3006);
nor U4638 (N_4638,N_3173,N_3984);
nor U4639 (N_4639,N_3516,N_3401);
and U4640 (N_4640,N_3408,N_3297);
xor U4641 (N_4641,N_3151,N_3118);
xnor U4642 (N_4642,N_3225,N_3694);
and U4643 (N_4643,N_3146,N_3211);
or U4644 (N_4644,N_3563,N_3046);
xnor U4645 (N_4645,N_3775,N_3143);
nand U4646 (N_4646,N_3686,N_3605);
and U4647 (N_4647,N_3251,N_3722);
and U4648 (N_4648,N_3919,N_3547);
xor U4649 (N_4649,N_3151,N_3000);
or U4650 (N_4650,N_3135,N_3150);
and U4651 (N_4651,N_3526,N_3226);
nand U4652 (N_4652,N_3980,N_3452);
nand U4653 (N_4653,N_3903,N_3990);
xnor U4654 (N_4654,N_3555,N_3238);
nor U4655 (N_4655,N_3927,N_3464);
and U4656 (N_4656,N_3929,N_3530);
nor U4657 (N_4657,N_3022,N_3824);
and U4658 (N_4658,N_3425,N_3481);
nand U4659 (N_4659,N_3903,N_3864);
and U4660 (N_4660,N_3696,N_3865);
or U4661 (N_4661,N_3985,N_3922);
xor U4662 (N_4662,N_3897,N_3833);
nand U4663 (N_4663,N_3659,N_3523);
and U4664 (N_4664,N_3256,N_3080);
and U4665 (N_4665,N_3883,N_3842);
nor U4666 (N_4666,N_3575,N_3953);
or U4667 (N_4667,N_3956,N_3240);
or U4668 (N_4668,N_3664,N_3847);
nand U4669 (N_4669,N_3404,N_3159);
or U4670 (N_4670,N_3361,N_3045);
nor U4671 (N_4671,N_3327,N_3510);
and U4672 (N_4672,N_3818,N_3891);
or U4673 (N_4673,N_3515,N_3063);
or U4674 (N_4674,N_3984,N_3587);
or U4675 (N_4675,N_3296,N_3177);
or U4676 (N_4676,N_3057,N_3775);
nor U4677 (N_4677,N_3414,N_3042);
xor U4678 (N_4678,N_3587,N_3460);
nand U4679 (N_4679,N_3632,N_3527);
nor U4680 (N_4680,N_3644,N_3822);
nor U4681 (N_4681,N_3960,N_3123);
nand U4682 (N_4682,N_3472,N_3707);
nor U4683 (N_4683,N_3022,N_3723);
xor U4684 (N_4684,N_3471,N_3133);
and U4685 (N_4685,N_3602,N_3136);
or U4686 (N_4686,N_3030,N_3984);
or U4687 (N_4687,N_3841,N_3148);
xnor U4688 (N_4688,N_3280,N_3338);
nor U4689 (N_4689,N_3026,N_3048);
nand U4690 (N_4690,N_3607,N_3469);
and U4691 (N_4691,N_3300,N_3436);
or U4692 (N_4692,N_3158,N_3525);
nor U4693 (N_4693,N_3766,N_3654);
nor U4694 (N_4694,N_3951,N_3008);
or U4695 (N_4695,N_3634,N_3261);
and U4696 (N_4696,N_3077,N_3650);
nand U4697 (N_4697,N_3305,N_3862);
nand U4698 (N_4698,N_3703,N_3488);
xor U4699 (N_4699,N_3474,N_3370);
xnor U4700 (N_4700,N_3102,N_3635);
nand U4701 (N_4701,N_3555,N_3250);
nor U4702 (N_4702,N_3582,N_3292);
nand U4703 (N_4703,N_3170,N_3676);
or U4704 (N_4704,N_3358,N_3552);
and U4705 (N_4705,N_3953,N_3873);
xor U4706 (N_4706,N_3058,N_3786);
nand U4707 (N_4707,N_3185,N_3103);
nor U4708 (N_4708,N_3457,N_3313);
or U4709 (N_4709,N_3589,N_3225);
and U4710 (N_4710,N_3109,N_3152);
xor U4711 (N_4711,N_3982,N_3539);
nand U4712 (N_4712,N_3556,N_3338);
and U4713 (N_4713,N_3297,N_3146);
or U4714 (N_4714,N_3922,N_3797);
nor U4715 (N_4715,N_3672,N_3567);
or U4716 (N_4716,N_3735,N_3290);
and U4717 (N_4717,N_3898,N_3502);
and U4718 (N_4718,N_3202,N_3329);
nand U4719 (N_4719,N_3987,N_3581);
nand U4720 (N_4720,N_3708,N_3847);
xor U4721 (N_4721,N_3281,N_3217);
nor U4722 (N_4722,N_3871,N_3906);
nor U4723 (N_4723,N_3335,N_3596);
and U4724 (N_4724,N_3199,N_3911);
nand U4725 (N_4725,N_3678,N_3384);
xor U4726 (N_4726,N_3360,N_3667);
and U4727 (N_4727,N_3869,N_3805);
nor U4728 (N_4728,N_3771,N_3502);
and U4729 (N_4729,N_3637,N_3322);
xnor U4730 (N_4730,N_3275,N_3737);
nand U4731 (N_4731,N_3980,N_3036);
nor U4732 (N_4732,N_3365,N_3261);
and U4733 (N_4733,N_3587,N_3915);
nor U4734 (N_4734,N_3813,N_3706);
nor U4735 (N_4735,N_3142,N_3098);
or U4736 (N_4736,N_3482,N_3161);
nand U4737 (N_4737,N_3350,N_3526);
nand U4738 (N_4738,N_3857,N_3965);
nor U4739 (N_4739,N_3546,N_3250);
and U4740 (N_4740,N_3077,N_3679);
xnor U4741 (N_4741,N_3381,N_3225);
or U4742 (N_4742,N_3260,N_3732);
or U4743 (N_4743,N_3763,N_3525);
xor U4744 (N_4744,N_3855,N_3811);
nor U4745 (N_4745,N_3791,N_3922);
nor U4746 (N_4746,N_3780,N_3397);
nand U4747 (N_4747,N_3424,N_3828);
or U4748 (N_4748,N_3257,N_3187);
or U4749 (N_4749,N_3346,N_3309);
nor U4750 (N_4750,N_3527,N_3235);
or U4751 (N_4751,N_3796,N_3555);
nor U4752 (N_4752,N_3183,N_3385);
and U4753 (N_4753,N_3819,N_3315);
nand U4754 (N_4754,N_3320,N_3545);
or U4755 (N_4755,N_3225,N_3519);
or U4756 (N_4756,N_3257,N_3062);
xor U4757 (N_4757,N_3968,N_3088);
nand U4758 (N_4758,N_3891,N_3100);
xor U4759 (N_4759,N_3189,N_3613);
nor U4760 (N_4760,N_3740,N_3097);
or U4761 (N_4761,N_3818,N_3128);
nand U4762 (N_4762,N_3640,N_3818);
nor U4763 (N_4763,N_3077,N_3779);
nor U4764 (N_4764,N_3137,N_3134);
nand U4765 (N_4765,N_3892,N_3969);
or U4766 (N_4766,N_3551,N_3200);
nand U4767 (N_4767,N_3256,N_3941);
nand U4768 (N_4768,N_3531,N_3758);
nor U4769 (N_4769,N_3802,N_3254);
nand U4770 (N_4770,N_3216,N_3974);
xnor U4771 (N_4771,N_3265,N_3117);
or U4772 (N_4772,N_3589,N_3510);
nand U4773 (N_4773,N_3416,N_3804);
or U4774 (N_4774,N_3316,N_3392);
xor U4775 (N_4775,N_3330,N_3901);
xnor U4776 (N_4776,N_3033,N_3956);
and U4777 (N_4777,N_3243,N_3289);
or U4778 (N_4778,N_3458,N_3714);
nor U4779 (N_4779,N_3667,N_3197);
xnor U4780 (N_4780,N_3634,N_3911);
nand U4781 (N_4781,N_3469,N_3348);
and U4782 (N_4782,N_3282,N_3685);
nand U4783 (N_4783,N_3105,N_3467);
nor U4784 (N_4784,N_3164,N_3178);
and U4785 (N_4785,N_3336,N_3513);
or U4786 (N_4786,N_3638,N_3744);
nand U4787 (N_4787,N_3718,N_3067);
and U4788 (N_4788,N_3003,N_3925);
xor U4789 (N_4789,N_3853,N_3006);
nor U4790 (N_4790,N_3070,N_3472);
nor U4791 (N_4791,N_3495,N_3496);
xnor U4792 (N_4792,N_3064,N_3881);
xor U4793 (N_4793,N_3989,N_3983);
or U4794 (N_4794,N_3103,N_3478);
or U4795 (N_4795,N_3208,N_3063);
nor U4796 (N_4796,N_3772,N_3217);
and U4797 (N_4797,N_3293,N_3800);
nor U4798 (N_4798,N_3584,N_3938);
nor U4799 (N_4799,N_3182,N_3216);
xor U4800 (N_4800,N_3754,N_3667);
nor U4801 (N_4801,N_3885,N_3339);
nor U4802 (N_4802,N_3359,N_3795);
or U4803 (N_4803,N_3802,N_3426);
or U4804 (N_4804,N_3215,N_3530);
and U4805 (N_4805,N_3355,N_3046);
nand U4806 (N_4806,N_3375,N_3851);
xnor U4807 (N_4807,N_3631,N_3280);
nor U4808 (N_4808,N_3244,N_3202);
xnor U4809 (N_4809,N_3840,N_3579);
nand U4810 (N_4810,N_3459,N_3288);
or U4811 (N_4811,N_3104,N_3843);
and U4812 (N_4812,N_3539,N_3435);
nor U4813 (N_4813,N_3148,N_3745);
or U4814 (N_4814,N_3909,N_3539);
and U4815 (N_4815,N_3401,N_3561);
nand U4816 (N_4816,N_3105,N_3817);
or U4817 (N_4817,N_3779,N_3944);
xnor U4818 (N_4818,N_3165,N_3664);
and U4819 (N_4819,N_3650,N_3838);
and U4820 (N_4820,N_3557,N_3705);
nor U4821 (N_4821,N_3250,N_3990);
nor U4822 (N_4822,N_3882,N_3709);
or U4823 (N_4823,N_3115,N_3195);
nand U4824 (N_4824,N_3596,N_3561);
and U4825 (N_4825,N_3211,N_3535);
nand U4826 (N_4826,N_3946,N_3252);
xor U4827 (N_4827,N_3082,N_3527);
xor U4828 (N_4828,N_3213,N_3793);
xor U4829 (N_4829,N_3866,N_3820);
nor U4830 (N_4830,N_3103,N_3923);
xnor U4831 (N_4831,N_3058,N_3744);
xor U4832 (N_4832,N_3318,N_3039);
and U4833 (N_4833,N_3355,N_3567);
nor U4834 (N_4834,N_3499,N_3433);
xor U4835 (N_4835,N_3833,N_3246);
nand U4836 (N_4836,N_3842,N_3714);
xnor U4837 (N_4837,N_3115,N_3658);
nor U4838 (N_4838,N_3539,N_3434);
and U4839 (N_4839,N_3298,N_3982);
nand U4840 (N_4840,N_3778,N_3038);
or U4841 (N_4841,N_3667,N_3912);
nor U4842 (N_4842,N_3846,N_3460);
nand U4843 (N_4843,N_3355,N_3734);
or U4844 (N_4844,N_3746,N_3813);
or U4845 (N_4845,N_3904,N_3694);
xnor U4846 (N_4846,N_3375,N_3010);
nor U4847 (N_4847,N_3382,N_3767);
xnor U4848 (N_4848,N_3252,N_3856);
nor U4849 (N_4849,N_3138,N_3340);
or U4850 (N_4850,N_3751,N_3363);
nor U4851 (N_4851,N_3479,N_3658);
or U4852 (N_4852,N_3902,N_3151);
nor U4853 (N_4853,N_3166,N_3796);
nor U4854 (N_4854,N_3463,N_3525);
or U4855 (N_4855,N_3790,N_3373);
or U4856 (N_4856,N_3791,N_3899);
or U4857 (N_4857,N_3717,N_3908);
or U4858 (N_4858,N_3785,N_3810);
nor U4859 (N_4859,N_3452,N_3955);
nand U4860 (N_4860,N_3521,N_3237);
or U4861 (N_4861,N_3730,N_3944);
nand U4862 (N_4862,N_3527,N_3240);
and U4863 (N_4863,N_3580,N_3407);
or U4864 (N_4864,N_3705,N_3370);
xor U4865 (N_4865,N_3885,N_3359);
xnor U4866 (N_4866,N_3258,N_3042);
nand U4867 (N_4867,N_3188,N_3835);
or U4868 (N_4868,N_3184,N_3294);
nand U4869 (N_4869,N_3782,N_3380);
or U4870 (N_4870,N_3221,N_3692);
xor U4871 (N_4871,N_3806,N_3788);
nand U4872 (N_4872,N_3825,N_3162);
or U4873 (N_4873,N_3483,N_3463);
or U4874 (N_4874,N_3449,N_3952);
and U4875 (N_4875,N_3464,N_3561);
nand U4876 (N_4876,N_3401,N_3279);
nor U4877 (N_4877,N_3571,N_3614);
xnor U4878 (N_4878,N_3495,N_3195);
or U4879 (N_4879,N_3006,N_3664);
nand U4880 (N_4880,N_3088,N_3367);
nor U4881 (N_4881,N_3143,N_3798);
or U4882 (N_4882,N_3382,N_3528);
or U4883 (N_4883,N_3970,N_3575);
or U4884 (N_4884,N_3471,N_3510);
and U4885 (N_4885,N_3925,N_3780);
nor U4886 (N_4886,N_3593,N_3194);
nor U4887 (N_4887,N_3065,N_3299);
nor U4888 (N_4888,N_3344,N_3627);
xnor U4889 (N_4889,N_3042,N_3196);
and U4890 (N_4890,N_3129,N_3150);
nor U4891 (N_4891,N_3414,N_3205);
and U4892 (N_4892,N_3692,N_3146);
or U4893 (N_4893,N_3485,N_3636);
nor U4894 (N_4894,N_3973,N_3870);
or U4895 (N_4895,N_3253,N_3758);
or U4896 (N_4896,N_3847,N_3051);
nand U4897 (N_4897,N_3033,N_3934);
nand U4898 (N_4898,N_3806,N_3141);
and U4899 (N_4899,N_3888,N_3980);
xor U4900 (N_4900,N_3308,N_3946);
xnor U4901 (N_4901,N_3398,N_3214);
nor U4902 (N_4902,N_3694,N_3367);
nor U4903 (N_4903,N_3310,N_3224);
xor U4904 (N_4904,N_3391,N_3982);
and U4905 (N_4905,N_3221,N_3872);
nor U4906 (N_4906,N_3880,N_3510);
nand U4907 (N_4907,N_3240,N_3505);
nand U4908 (N_4908,N_3272,N_3155);
nand U4909 (N_4909,N_3364,N_3401);
xor U4910 (N_4910,N_3525,N_3952);
or U4911 (N_4911,N_3924,N_3657);
nor U4912 (N_4912,N_3509,N_3241);
or U4913 (N_4913,N_3897,N_3296);
xor U4914 (N_4914,N_3113,N_3509);
nand U4915 (N_4915,N_3051,N_3260);
nor U4916 (N_4916,N_3111,N_3524);
nor U4917 (N_4917,N_3488,N_3731);
nand U4918 (N_4918,N_3253,N_3633);
xor U4919 (N_4919,N_3724,N_3138);
nand U4920 (N_4920,N_3573,N_3223);
or U4921 (N_4921,N_3685,N_3519);
or U4922 (N_4922,N_3611,N_3577);
xnor U4923 (N_4923,N_3904,N_3006);
nand U4924 (N_4924,N_3446,N_3537);
xnor U4925 (N_4925,N_3206,N_3192);
xor U4926 (N_4926,N_3164,N_3965);
or U4927 (N_4927,N_3278,N_3428);
xnor U4928 (N_4928,N_3156,N_3914);
and U4929 (N_4929,N_3205,N_3267);
xnor U4930 (N_4930,N_3790,N_3460);
and U4931 (N_4931,N_3848,N_3662);
or U4932 (N_4932,N_3741,N_3823);
and U4933 (N_4933,N_3604,N_3988);
and U4934 (N_4934,N_3207,N_3167);
or U4935 (N_4935,N_3789,N_3280);
nand U4936 (N_4936,N_3902,N_3364);
nor U4937 (N_4937,N_3128,N_3875);
nand U4938 (N_4938,N_3087,N_3785);
nor U4939 (N_4939,N_3344,N_3676);
nor U4940 (N_4940,N_3802,N_3880);
nand U4941 (N_4941,N_3013,N_3868);
nor U4942 (N_4942,N_3466,N_3584);
and U4943 (N_4943,N_3234,N_3959);
nand U4944 (N_4944,N_3750,N_3032);
or U4945 (N_4945,N_3273,N_3562);
and U4946 (N_4946,N_3696,N_3803);
and U4947 (N_4947,N_3227,N_3429);
nand U4948 (N_4948,N_3177,N_3168);
or U4949 (N_4949,N_3447,N_3159);
nand U4950 (N_4950,N_3921,N_3114);
nand U4951 (N_4951,N_3354,N_3162);
or U4952 (N_4952,N_3740,N_3760);
nand U4953 (N_4953,N_3308,N_3847);
nand U4954 (N_4954,N_3014,N_3103);
and U4955 (N_4955,N_3451,N_3648);
nand U4956 (N_4956,N_3485,N_3040);
or U4957 (N_4957,N_3656,N_3918);
nand U4958 (N_4958,N_3501,N_3315);
xnor U4959 (N_4959,N_3858,N_3989);
nor U4960 (N_4960,N_3266,N_3709);
or U4961 (N_4961,N_3162,N_3498);
nor U4962 (N_4962,N_3346,N_3885);
nand U4963 (N_4963,N_3560,N_3696);
xnor U4964 (N_4964,N_3145,N_3886);
xor U4965 (N_4965,N_3527,N_3307);
nand U4966 (N_4966,N_3415,N_3468);
nor U4967 (N_4967,N_3788,N_3493);
and U4968 (N_4968,N_3480,N_3080);
or U4969 (N_4969,N_3685,N_3053);
nand U4970 (N_4970,N_3844,N_3566);
and U4971 (N_4971,N_3473,N_3082);
and U4972 (N_4972,N_3171,N_3265);
nand U4973 (N_4973,N_3133,N_3848);
or U4974 (N_4974,N_3803,N_3921);
nor U4975 (N_4975,N_3979,N_3243);
nand U4976 (N_4976,N_3847,N_3852);
xnor U4977 (N_4977,N_3064,N_3459);
or U4978 (N_4978,N_3219,N_3140);
xor U4979 (N_4979,N_3620,N_3922);
xor U4980 (N_4980,N_3239,N_3211);
or U4981 (N_4981,N_3394,N_3059);
or U4982 (N_4982,N_3474,N_3569);
xor U4983 (N_4983,N_3650,N_3614);
xnor U4984 (N_4984,N_3605,N_3330);
or U4985 (N_4985,N_3392,N_3047);
nand U4986 (N_4986,N_3369,N_3188);
or U4987 (N_4987,N_3929,N_3677);
or U4988 (N_4988,N_3524,N_3906);
xnor U4989 (N_4989,N_3604,N_3535);
xnor U4990 (N_4990,N_3439,N_3713);
or U4991 (N_4991,N_3466,N_3742);
xnor U4992 (N_4992,N_3851,N_3239);
or U4993 (N_4993,N_3104,N_3543);
nand U4994 (N_4994,N_3996,N_3291);
and U4995 (N_4995,N_3217,N_3725);
and U4996 (N_4996,N_3760,N_3175);
and U4997 (N_4997,N_3001,N_3777);
and U4998 (N_4998,N_3776,N_3746);
or U4999 (N_4999,N_3380,N_3129);
nand U5000 (N_5000,N_4090,N_4544);
nor U5001 (N_5001,N_4583,N_4380);
and U5002 (N_5002,N_4297,N_4860);
nor U5003 (N_5003,N_4892,N_4674);
xor U5004 (N_5004,N_4741,N_4283);
nand U5005 (N_5005,N_4321,N_4653);
or U5006 (N_5006,N_4087,N_4398);
nor U5007 (N_5007,N_4926,N_4349);
xor U5008 (N_5008,N_4091,N_4346);
nor U5009 (N_5009,N_4226,N_4996);
nor U5010 (N_5010,N_4292,N_4818);
nor U5011 (N_5011,N_4855,N_4467);
or U5012 (N_5012,N_4964,N_4357);
xnor U5013 (N_5013,N_4714,N_4065);
xor U5014 (N_5014,N_4538,N_4883);
and U5015 (N_5015,N_4819,N_4061);
or U5016 (N_5016,N_4096,N_4602);
nor U5017 (N_5017,N_4198,N_4491);
and U5018 (N_5018,N_4811,N_4037);
or U5019 (N_5019,N_4638,N_4794);
or U5020 (N_5020,N_4401,N_4956);
or U5021 (N_5021,N_4399,N_4842);
nor U5022 (N_5022,N_4146,N_4421);
and U5023 (N_5023,N_4826,N_4940);
nor U5024 (N_5024,N_4931,N_4129);
or U5025 (N_5025,N_4231,N_4806);
nor U5026 (N_5026,N_4269,N_4325);
nand U5027 (N_5027,N_4577,N_4907);
nand U5028 (N_5028,N_4856,N_4782);
nor U5029 (N_5029,N_4257,N_4954);
nand U5030 (N_5030,N_4541,N_4063);
xnor U5031 (N_5031,N_4086,N_4507);
and U5032 (N_5032,N_4518,N_4685);
and U5033 (N_5033,N_4650,N_4625);
and U5034 (N_5034,N_4145,N_4698);
nand U5035 (N_5035,N_4252,N_4902);
nand U5036 (N_5036,N_4254,N_4118);
nand U5037 (N_5037,N_4026,N_4447);
nor U5038 (N_5038,N_4081,N_4578);
nor U5039 (N_5039,N_4052,N_4924);
nand U5040 (N_5040,N_4953,N_4114);
xor U5041 (N_5041,N_4763,N_4950);
xor U5042 (N_5042,N_4792,N_4474);
and U5043 (N_5043,N_4732,N_4360);
nand U5044 (N_5044,N_4497,N_4138);
and U5045 (N_5045,N_4862,N_4298);
xnor U5046 (N_5046,N_4895,N_4143);
or U5047 (N_5047,N_4024,N_4215);
nand U5048 (N_5048,N_4958,N_4821);
or U5049 (N_5049,N_4783,N_4069);
xnor U5050 (N_5050,N_4880,N_4475);
nand U5051 (N_5051,N_4457,N_4050);
nor U5052 (N_5052,N_4400,N_4709);
nor U5053 (N_5053,N_4974,N_4540);
nor U5054 (N_5054,N_4224,N_4847);
and U5055 (N_5055,N_4896,N_4435);
nand U5056 (N_5056,N_4867,N_4798);
or U5057 (N_5057,N_4678,N_4567);
nor U5058 (N_5058,N_4897,N_4730);
nand U5059 (N_5059,N_4075,N_4780);
nand U5060 (N_5060,N_4209,N_4484);
xnor U5061 (N_5061,N_4085,N_4303);
nand U5062 (N_5062,N_4828,N_4428);
or U5063 (N_5063,N_4839,N_4412);
nor U5064 (N_5064,N_4968,N_4492);
xnor U5065 (N_5065,N_4424,N_4749);
or U5066 (N_5066,N_4948,N_4604);
and U5067 (N_5067,N_4535,N_4468);
nor U5068 (N_5068,N_4162,N_4785);
nor U5069 (N_5069,N_4553,N_4773);
and U5070 (N_5070,N_4888,N_4779);
nand U5071 (N_5071,N_4098,N_4857);
xnor U5072 (N_5072,N_4853,N_4003);
nor U5073 (N_5073,N_4356,N_4432);
xnor U5074 (N_5074,N_4493,N_4980);
nand U5075 (N_5075,N_4646,N_4368);
or U5076 (N_5076,N_4726,N_4791);
and U5077 (N_5077,N_4595,N_4848);
nand U5078 (N_5078,N_4758,N_4031);
nand U5079 (N_5079,N_4654,N_4295);
nand U5080 (N_5080,N_4177,N_4530);
or U5081 (N_5081,N_4433,N_4438);
or U5082 (N_5082,N_4757,N_4374);
nand U5083 (N_5083,N_4988,N_4232);
nor U5084 (N_5084,N_4223,N_4505);
or U5085 (N_5085,N_4942,N_4205);
nor U5086 (N_5086,N_4967,N_4367);
and U5087 (N_5087,N_4584,N_4999);
nor U5088 (N_5088,N_4861,N_4289);
xnor U5089 (N_5089,N_4594,N_4469);
nand U5090 (N_5090,N_4204,N_4528);
or U5091 (N_5091,N_4719,N_4248);
xnor U5092 (N_5092,N_4846,N_4586);
nor U5093 (N_5093,N_4918,N_4001);
nor U5094 (N_5094,N_4312,N_4249);
xnor U5095 (N_5095,N_4179,N_4748);
and U5096 (N_5096,N_4620,N_4803);
and U5097 (N_5097,N_4489,N_4745);
and U5098 (N_5098,N_4152,N_4273);
nand U5099 (N_5099,N_4957,N_4739);
nor U5100 (N_5100,N_4488,N_4127);
xor U5101 (N_5101,N_4603,N_4669);
or U5102 (N_5102,N_4550,N_4606);
nand U5103 (N_5103,N_4291,N_4652);
and U5104 (N_5104,N_4245,N_4559);
nor U5105 (N_5105,N_4103,N_4120);
xor U5106 (N_5106,N_4724,N_4621);
nor U5107 (N_5107,N_4680,N_4569);
and U5108 (N_5108,N_4824,N_4391);
or U5109 (N_5109,N_4004,N_4115);
nor U5110 (N_5110,N_4056,N_4738);
nand U5111 (N_5111,N_4694,N_4985);
xnor U5112 (N_5112,N_4173,N_4994);
or U5113 (N_5113,N_4376,N_4844);
xor U5114 (N_5114,N_4728,N_4139);
nand U5115 (N_5115,N_4986,N_4126);
xnor U5116 (N_5116,N_4328,N_4419);
and U5117 (N_5117,N_4919,N_4845);
or U5118 (N_5118,N_4703,N_4000);
or U5119 (N_5119,N_4079,N_4626);
and U5120 (N_5120,N_4175,N_4765);
nand U5121 (N_5121,N_4210,N_4350);
or U5122 (N_5122,N_4201,N_4352);
nand U5123 (N_5123,N_4264,N_4941);
and U5124 (N_5124,N_4643,N_4082);
xor U5125 (N_5125,N_4080,N_4045);
and U5126 (N_5126,N_4333,N_4387);
nand U5127 (N_5127,N_4440,N_4416);
nor U5128 (N_5128,N_4556,N_4827);
nand U5129 (N_5129,N_4099,N_4822);
xor U5130 (N_5130,N_4723,N_4668);
and U5131 (N_5131,N_4989,N_4624);
nor U5132 (N_5132,N_4239,N_4908);
nor U5133 (N_5133,N_4351,N_4422);
and U5134 (N_5134,N_4263,N_4814);
nand U5135 (N_5135,N_4673,N_4778);
nor U5136 (N_5136,N_4453,N_4925);
xnor U5137 (N_5137,N_4557,N_4163);
or U5138 (N_5138,N_4952,N_4025);
and U5139 (N_5139,N_4051,N_4256);
nand U5140 (N_5140,N_4397,N_4459);
and U5141 (N_5141,N_4898,N_4364);
nand U5142 (N_5142,N_4211,N_4221);
nand U5143 (N_5143,N_4027,N_4700);
and U5144 (N_5144,N_4150,N_4002);
nand U5145 (N_5145,N_4601,N_4969);
nor U5146 (N_5146,N_4884,N_4377);
and U5147 (N_5147,N_4057,N_4049);
xnor U5148 (N_5148,N_4384,N_4890);
nor U5149 (N_5149,N_4006,N_4921);
nand U5150 (N_5150,N_4287,N_4716);
xor U5151 (N_5151,N_4308,N_4928);
nor U5152 (N_5152,N_4022,N_4517);
nor U5153 (N_5153,N_4592,N_4191);
xor U5154 (N_5154,N_4927,N_4587);
or U5155 (N_5155,N_4236,N_4717);
and U5156 (N_5156,N_4111,N_4032);
xor U5157 (N_5157,N_4310,N_4666);
and U5158 (N_5158,N_4914,N_4463);
xor U5159 (N_5159,N_4555,N_4410);
and U5160 (N_5160,N_4913,N_4119);
nand U5161 (N_5161,N_4326,N_4562);
xnor U5162 (N_5162,N_4502,N_4406);
and U5163 (N_5163,N_4202,N_4702);
nor U5164 (N_5164,N_4864,N_4677);
or U5165 (N_5165,N_4059,N_4268);
xnor U5166 (N_5166,N_4704,N_4481);
nand U5167 (N_5167,N_4414,N_4670);
xor U5168 (N_5168,N_4392,N_4966);
nand U5169 (N_5169,N_4279,N_4010);
xor U5170 (N_5170,N_4789,N_4165);
or U5171 (N_5171,N_4509,N_4110);
and U5172 (N_5172,N_4722,N_4740);
and U5173 (N_5173,N_4551,N_4452);
xnor U5174 (N_5174,N_4100,N_4200);
nor U5175 (N_5175,N_4238,N_4105);
nand U5176 (N_5176,N_4318,N_4690);
nor U5177 (N_5177,N_4344,N_4571);
xor U5178 (N_5178,N_4990,N_4074);
nor U5179 (N_5179,N_4686,N_4005);
and U5180 (N_5180,N_4471,N_4949);
nand U5181 (N_5181,N_4532,N_4102);
nor U5182 (N_5182,N_4870,N_4799);
and U5183 (N_5183,N_4007,N_4131);
and U5184 (N_5184,N_4598,N_4446);
xnor U5185 (N_5185,N_4886,N_4186);
and U5186 (N_5186,N_4930,N_4899);
xnor U5187 (N_5187,N_4564,N_4213);
and U5188 (N_5188,N_4802,N_4676);
and U5189 (N_5189,N_4539,N_4476);
nor U5190 (N_5190,N_4011,N_4154);
nand U5191 (N_5191,N_4906,N_4515);
and U5192 (N_5192,N_4813,N_4834);
nor U5193 (N_5193,N_4575,N_4465);
xnor U5194 (N_5194,N_4012,N_4720);
or U5195 (N_5195,N_4991,N_4448);
or U5196 (N_5196,N_4649,N_4591);
nand U5197 (N_5197,N_4938,N_4565);
or U5198 (N_5198,N_4640,N_4036);
or U5199 (N_5199,N_4237,N_4288);
or U5200 (N_5200,N_4379,N_4657);
and U5201 (N_5201,N_4825,N_4317);
xnor U5202 (N_5202,N_4997,N_4570);
and U5203 (N_5203,N_4258,N_4527);
xor U5204 (N_5204,N_4889,N_4337);
xor U5205 (N_5205,N_4608,N_4373);
nor U5206 (N_5206,N_4281,N_4441);
nor U5207 (N_5207,N_4929,N_4563);
xor U5208 (N_5208,N_4746,N_4240);
nor U5209 (N_5209,N_4663,N_4342);
and U5210 (N_5210,N_4250,N_4167);
nor U5211 (N_5211,N_4188,N_4083);
and U5212 (N_5212,N_4797,N_4836);
xor U5213 (N_5213,N_4104,N_4199);
and U5214 (N_5214,N_4151,N_4869);
nor U5215 (N_5215,N_4766,N_4504);
nor U5216 (N_5216,N_4547,N_4656);
or U5217 (N_5217,N_4498,N_4113);
nand U5218 (N_5218,N_4284,N_4731);
xnor U5219 (N_5219,N_4585,N_4434);
nand U5220 (N_5220,N_4180,N_4658);
nand U5221 (N_5221,N_4615,N_4235);
or U5222 (N_5222,N_4692,N_4920);
or U5223 (N_5223,N_4496,N_4993);
nand U5224 (N_5224,N_4275,N_4753);
nor U5225 (N_5225,N_4194,N_4047);
and U5226 (N_5226,N_4411,N_4353);
nor U5227 (N_5227,N_4420,N_4216);
nand U5228 (N_5228,N_4536,N_4361);
or U5229 (N_5229,N_4128,N_4568);
and U5230 (N_5230,N_4922,N_4381);
xnor U5231 (N_5231,N_4259,N_4939);
and U5232 (N_5232,N_4599,N_4593);
or U5233 (N_5233,N_4750,N_4072);
or U5234 (N_5234,N_4230,N_4286);
nand U5235 (N_5235,N_4451,N_4158);
xor U5236 (N_5236,N_4648,N_4442);
and U5237 (N_5237,N_4659,N_4875);
or U5238 (N_5238,N_4516,N_4644);
nand U5239 (N_5239,N_4262,N_4519);
nand U5240 (N_5240,N_4106,N_4808);
nand U5241 (N_5241,N_4332,N_4871);
or U5242 (N_5242,N_4909,N_4514);
nor U5243 (N_5243,N_4088,N_4971);
xnor U5244 (N_5244,N_4294,N_4937);
nor U5245 (N_5245,N_4034,N_4636);
nor U5246 (N_5246,N_4833,N_4588);
nor U5247 (N_5247,N_4157,N_4960);
nand U5248 (N_5248,N_4382,N_4097);
and U5249 (N_5249,N_4545,N_4979);
and U5250 (N_5250,N_4891,N_4214);
nand U5251 (N_5251,N_4030,N_4632);
and U5252 (N_5252,N_4522,N_4962);
and U5253 (N_5253,N_4309,N_4133);
nor U5254 (N_5254,N_4521,N_4835);
nor U5255 (N_5255,N_4661,N_4271);
or U5256 (N_5256,N_4301,N_4580);
or U5257 (N_5257,N_4543,N_4529);
and U5258 (N_5258,N_4850,N_4729);
nor U5259 (N_5259,N_4747,N_4959);
nor U5260 (N_5260,N_4417,N_4267);
xnor U5261 (N_5261,N_4480,N_4721);
and U5262 (N_5262,N_4296,N_4572);
nand U5263 (N_5263,N_4616,N_4781);
and U5264 (N_5264,N_4334,N_4458);
or U5265 (N_5265,N_4241,N_4371);
xor U5266 (N_5266,N_4560,N_4718);
xnor U5267 (N_5267,N_4987,N_4184);
xor U5268 (N_5268,N_4174,N_4073);
or U5269 (N_5269,N_4117,N_4917);
nand U5270 (N_5270,N_4060,N_4637);
nand U5271 (N_5271,N_4067,N_4627);
and U5272 (N_5272,N_4218,N_4044);
xor U5273 (N_5273,N_4490,N_4708);
xnor U5274 (N_5274,N_4647,N_4109);
and U5275 (N_5275,N_4655,N_4816);
nor U5276 (N_5276,N_4423,N_4915);
nand U5277 (N_5277,N_4089,N_4378);
nor U5278 (N_5278,N_4715,N_4299);
or U5279 (N_5279,N_4878,N_4479);
nor U5280 (N_5280,N_4300,N_4372);
nand U5281 (N_5281,N_4623,N_4710);
xor U5282 (N_5282,N_4134,N_4068);
and U5283 (N_5283,N_4664,N_4450);
xnor U5284 (N_5284,N_4343,N_4195);
xor U5285 (N_5285,N_4837,N_4831);
and U5286 (N_5286,N_4338,N_4774);
nand U5287 (N_5287,N_4307,N_4478);
or U5288 (N_5288,N_4243,N_4176);
and U5289 (N_5289,N_4701,N_4156);
or U5290 (N_5290,N_4095,N_4339);
and U5291 (N_5291,N_4501,N_4590);
nor U5292 (N_5292,N_4169,N_4066);
and U5293 (N_5293,N_4358,N_4932);
and U5294 (N_5294,N_4893,N_4903);
xnor U5295 (N_5295,N_4613,N_4612);
or U5296 (N_5296,N_4153,N_4879);
or U5297 (N_5297,N_4018,N_4212);
nor U5298 (N_5298,N_4054,N_4040);
xor U5299 (N_5299,N_4092,N_4029);
and U5300 (N_5300,N_4123,N_4359);
nand U5301 (N_5301,N_4282,N_4520);
and U5302 (N_5302,N_4220,N_4172);
xor U5303 (N_5303,N_4689,N_4800);
xor U5304 (N_5304,N_4375,N_4038);
nor U5305 (N_5305,N_4125,N_4777);
or U5306 (N_5306,N_4976,N_4735);
nand U5307 (N_5307,N_4630,N_4511);
nand U5308 (N_5308,N_4019,N_4341);
and U5309 (N_5309,N_4865,N_4852);
and U5310 (N_5310,N_4208,N_4436);
nor U5311 (N_5311,N_4671,N_4619);
xnor U5312 (N_5312,N_4877,N_4963);
nor U5313 (N_5313,N_4354,N_4234);
xnor U5314 (N_5314,N_4526,N_4331);
or U5315 (N_5315,N_4265,N_4549);
xor U5316 (N_5316,N_4048,N_4181);
nand U5317 (N_5317,N_4854,N_4820);
or U5318 (N_5318,N_4764,N_4278);
xnor U5319 (N_5319,N_4266,N_4445);
or U5320 (N_5320,N_4874,N_4682);
nor U5321 (N_5321,N_4314,N_4322);
nor U5322 (N_5322,N_4166,N_4039);
nor U5323 (N_5323,N_4116,N_4193);
nor U5324 (N_5324,N_4840,N_4135);
nor U5325 (N_5325,N_4768,N_4829);
or U5326 (N_5326,N_4810,N_4992);
or U5327 (N_5327,N_4635,N_4759);
and U5328 (N_5328,N_4933,N_4508);
xor U5329 (N_5329,N_4093,N_4253);
and U5330 (N_5330,N_4662,N_4229);
nor U5331 (N_5331,N_4772,N_4946);
nor U5332 (N_5332,N_4071,N_4455);
or U5333 (N_5333,N_4429,N_4881);
nor U5334 (N_5334,N_4631,N_4155);
xor U5335 (N_5335,N_4013,N_4274);
xnor U5336 (N_5336,N_4693,N_4147);
nand U5337 (N_5337,N_4363,N_4628);
or U5338 (N_5338,N_4887,N_4751);
xnor U5339 (N_5339,N_4485,N_4470);
nand U5340 (N_5340,N_4769,N_4043);
and U5341 (N_5341,N_4622,N_4255);
and U5342 (N_5342,N_4244,N_4904);
nand U5343 (N_5343,N_4629,N_4943);
nor U5344 (N_5344,N_4524,N_4639);
nand U5345 (N_5345,N_4542,N_4149);
or U5346 (N_5346,N_4576,N_4984);
or U5347 (N_5347,N_4160,N_4805);
or U5348 (N_5348,N_4923,N_4672);
nand U5349 (N_5349,N_4605,N_4159);
nand U5350 (N_5350,N_4633,N_4078);
nor U5351 (N_5351,N_4355,N_4832);
nor U5352 (N_5352,N_4033,N_4407);
nor U5353 (N_5353,N_4734,N_4276);
and U5354 (N_5354,N_4130,N_4998);
xor U5355 (N_5355,N_4665,N_4634);
nand U5356 (N_5356,N_4660,N_4849);
nand U5357 (N_5357,N_4062,N_4807);
nor U5358 (N_5358,N_4132,N_4965);
nor U5359 (N_5359,N_4449,N_4841);
nor U5360 (N_5360,N_4472,N_4064);
nand U5361 (N_5361,N_4260,N_4020);
nor U5362 (N_5362,N_4280,N_4618);
xor U5363 (N_5363,N_4916,N_4675);
nand U5364 (N_5364,N_4936,N_4456);
or U5365 (N_5365,N_4396,N_4512);
or U5366 (N_5366,N_4596,N_4461);
xnor U5367 (N_5367,N_4614,N_4046);
and U5368 (N_5368,N_4743,N_4561);
nor U5369 (N_5369,N_4144,N_4246);
or U5370 (N_5370,N_4369,N_4403);
nor U5371 (N_5371,N_4136,N_4684);
nor U5372 (N_5372,N_4405,N_4972);
and U5373 (N_5373,N_4737,N_4454);
nor U5374 (N_5374,N_4983,N_4219);
nand U5375 (N_5375,N_4513,N_4319);
nor U5376 (N_5376,N_4609,N_4466);
nand U5377 (N_5377,N_4679,N_4021);
nor U5378 (N_5378,N_4207,N_4164);
nand U5379 (N_5379,N_4304,N_4365);
xor U5380 (N_5380,N_4311,N_4336);
or U5381 (N_5381,N_4222,N_4141);
nand U5382 (N_5382,N_4531,N_4911);
nand U5383 (N_5383,N_4028,N_4537);
or U5384 (N_5384,N_4431,N_4305);
nand U5385 (N_5385,N_4823,N_4947);
or U5386 (N_5386,N_4077,N_4042);
nor U5387 (N_5387,N_4611,N_4945);
xor U5388 (N_5388,N_4770,N_4444);
or U5389 (N_5389,N_4389,N_4329);
nor U5390 (N_5390,N_4752,N_4885);
nor U5391 (N_5391,N_4793,N_4124);
xnor U5392 (N_5392,N_4755,N_4418);
nor U5393 (N_5393,N_4610,N_4784);
nand U5394 (N_5394,N_4699,N_4761);
nand U5395 (N_5395,N_4394,N_4206);
and U5396 (N_5396,N_4838,N_4320);
or U5397 (N_5397,N_4094,N_4788);
or U5398 (N_5398,N_4487,N_4995);
nand U5399 (N_5399,N_4754,N_4651);
or U5400 (N_5400,N_4863,N_4787);
or U5401 (N_5401,N_4041,N_4712);
nand U5402 (N_5402,N_4285,N_4951);
nand U5403 (N_5403,N_4443,N_4121);
nor U5404 (N_5404,N_4617,N_4168);
xnor U5405 (N_5405,N_4137,N_4302);
nand U5406 (N_5406,N_4771,N_4227);
nand U5407 (N_5407,N_4696,N_4462);
xnor U5408 (N_5408,N_4189,N_4786);
xnor U5409 (N_5409,N_4801,N_4776);
or U5410 (N_5410,N_4101,N_4477);
and U5411 (N_5411,N_4760,N_4395);
and U5412 (N_5412,N_4313,N_4736);
and U5413 (N_5413,N_4548,N_4713);
and U5414 (N_5414,N_4574,N_4706);
xor U5415 (N_5415,N_4641,N_4733);
and U5416 (N_5416,N_4324,N_4464);
or U5417 (N_5417,N_4579,N_4796);
or U5418 (N_5418,N_4247,N_4185);
nand U5419 (N_5419,N_4430,N_4261);
nand U5420 (N_5420,N_4830,N_4843);
nor U5421 (N_5421,N_4582,N_4494);
and U5422 (N_5422,N_4348,N_4055);
xor U5423 (N_5423,N_4725,N_4170);
and U5424 (N_5424,N_4683,N_4330);
or U5425 (N_5425,N_4882,N_4795);
nor U5426 (N_5426,N_4607,N_4015);
nor U5427 (N_5427,N_4345,N_4695);
and U5428 (N_5428,N_4552,N_4977);
xor U5429 (N_5429,N_4499,N_4554);
nor U5430 (N_5430,N_4973,N_4390);
nor U5431 (N_5431,N_4335,N_4014);
or U5432 (N_5432,N_4866,N_4386);
nor U5433 (N_5433,N_4762,N_4182);
nand U5434 (N_5434,N_4009,N_4197);
nand U5435 (N_5435,N_4727,N_4233);
nor U5436 (N_5436,N_4366,N_4851);
xnor U5437 (N_5437,N_4961,N_4894);
or U5438 (N_5438,N_4293,N_4868);
and U5439 (N_5439,N_4171,N_4597);
nor U5440 (N_5440,N_4272,N_4427);
xor U5441 (N_5441,N_4196,N_4402);
xor U5442 (N_5442,N_4362,N_4183);
nand U5443 (N_5443,N_4978,N_4905);
nand U5444 (N_5444,N_4053,N_4642);
nor U5445 (N_5445,N_4858,N_4142);
nand U5446 (N_5446,N_4122,N_4645);
or U5447 (N_5447,N_4935,N_4008);
xor U5448 (N_5448,N_4228,N_4178);
xor U5449 (N_5449,N_4681,N_4016);
nor U5450 (N_5450,N_4790,N_4534);
and U5451 (N_5451,N_4190,N_4315);
nand U5452 (N_5452,N_4711,N_4667);
xnor U5453 (N_5453,N_4691,N_4900);
nand U5454 (N_5454,N_4187,N_4503);
nor U5455 (N_5455,N_4910,N_4944);
or U5456 (N_5456,N_4327,N_4775);
or U5457 (N_5457,N_4161,N_4873);
xor U5458 (N_5458,N_4510,N_4388);
xor U5459 (N_5459,N_4408,N_4473);
or U5460 (N_5460,N_4756,N_4558);
xor U5461 (N_5461,N_4108,N_4705);
or U5462 (N_5462,N_4409,N_4306);
xnor U5463 (N_5463,N_4385,N_4934);
nor U5464 (N_5464,N_4566,N_4076);
nor U5465 (N_5465,N_4483,N_4573);
xnor U5466 (N_5466,N_4546,N_4217);
and U5467 (N_5467,N_4316,N_4437);
nor U5468 (N_5468,N_4697,N_4859);
nor U5469 (N_5469,N_4817,N_4525);
or U5470 (N_5470,N_4383,N_4815);
nor U5471 (N_5471,N_4404,N_4533);
nand U5472 (N_5472,N_4581,N_4148);
xor U5473 (N_5473,N_4370,N_4707);
and U5474 (N_5474,N_4460,N_4975);
and U5475 (N_5475,N_4688,N_4486);
or U5476 (N_5476,N_4140,N_4901);
nand U5477 (N_5477,N_4912,N_4290);
nand U5478 (N_5478,N_4482,N_4523);
nor U5479 (N_5479,N_4500,N_4084);
and U5480 (N_5480,N_4812,N_4340);
or U5481 (N_5481,N_4251,N_4225);
xor U5482 (N_5482,N_4981,N_4955);
nor U5483 (N_5483,N_4742,N_4242);
nand U5484 (N_5484,N_4023,N_4347);
nand U5485 (N_5485,N_4876,N_4277);
and U5486 (N_5486,N_4017,N_4426);
and U5487 (N_5487,N_4804,N_4600);
or U5488 (N_5488,N_4393,N_4982);
nor U5489 (N_5489,N_4323,N_4495);
and U5490 (N_5490,N_4107,N_4872);
nand U5491 (N_5491,N_4744,N_4425);
or U5492 (N_5492,N_4687,N_4035);
nand U5493 (N_5493,N_4413,N_4809);
nor U5494 (N_5494,N_4415,N_4767);
or U5495 (N_5495,N_4589,N_4070);
or U5496 (N_5496,N_4192,N_4439);
nand U5497 (N_5497,N_4970,N_4506);
or U5498 (N_5498,N_4112,N_4270);
and U5499 (N_5499,N_4058,N_4203);
nor U5500 (N_5500,N_4156,N_4050);
nor U5501 (N_5501,N_4682,N_4227);
nand U5502 (N_5502,N_4165,N_4712);
nor U5503 (N_5503,N_4164,N_4548);
or U5504 (N_5504,N_4859,N_4337);
xnor U5505 (N_5505,N_4112,N_4141);
nor U5506 (N_5506,N_4631,N_4021);
nor U5507 (N_5507,N_4283,N_4963);
nand U5508 (N_5508,N_4865,N_4300);
xnor U5509 (N_5509,N_4910,N_4644);
or U5510 (N_5510,N_4136,N_4671);
nor U5511 (N_5511,N_4344,N_4194);
nor U5512 (N_5512,N_4645,N_4129);
nor U5513 (N_5513,N_4847,N_4030);
xor U5514 (N_5514,N_4382,N_4790);
and U5515 (N_5515,N_4935,N_4937);
nand U5516 (N_5516,N_4961,N_4788);
and U5517 (N_5517,N_4613,N_4701);
and U5518 (N_5518,N_4021,N_4979);
and U5519 (N_5519,N_4801,N_4388);
nand U5520 (N_5520,N_4721,N_4007);
xor U5521 (N_5521,N_4864,N_4723);
xnor U5522 (N_5522,N_4731,N_4968);
or U5523 (N_5523,N_4370,N_4770);
or U5524 (N_5524,N_4210,N_4277);
or U5525 (N_5525,N_4159,N_4962);
xor U5526 (N_5526,N_4059,N_4815);
nor U5527 (N_5527,N_4858,N_4045);
nand U5528 (N_5528,N_4833,N_4874);
or U5529 (N_5529,N_4877,N_4412);
xor U5530 (N_5530,N_4175,N_4598);
or U5531 (N_5531,N_4491,N_4283);
nor U5532 (N_5532,N_4387,N_4325);
nand U5533 (N_5533,N_4158,N_4095);
xnor U5534 (N_5534,N_4273,N_4591);
nand U5535 (N_5535,N_4108,N_4202);
nand U5536 (N_5536,N_4777,N_4280);
xor U5537 (N_5537,N_4496,N_4468);
nor U5538 (N_5538,N_4603,N_4475);
xor U5539 (N_5539,N_4484,N_4544);
or U5540 (N_5540,N_4447,N_4944);
nand U5541 (N_5541,N_4734,N_4307);
xnor U5542 (N_5542,N_4912,N_4543);
nor U5543 (N_5543,N_4644,N_4451);
nand U5544 (N_5544,N_4216,N_4458);
and U5545 (N_5545,N_4372,N_4506);
nor U5546 (N_5546,N_4845,N_4544);
or U5547 (N_5547,N_4954,N_4246);
xnor U5548 (N_5548,N_4616,N_4946);
or U5549 (N_5549,N_4117,N_4249);
or U5550 (N_5550,N_4301,N_4669);
and U5551 (N_5551,N_4734,N_4858);
or U5552 (N_5552,N_4032,N_4669);
or U5553 (N_5553,N_4694,N_4418);
nor U5554 (N_5554,N_4466,N_4594);
and U5555 (N_5555,N_4170,N_4556);
or U5556 (N_5556,N_4118,N_4140);
or U5557 (N_5557,N_4616,N_4563);
xor U5558 (N_5558,N_4971,N_4449);
and U5559 (N_5559,N_4343,N_4059);
nand U5560 (N_5560,N_4552,N_4652);
xor U5561 (N_5561,N_4093,N_4388);
or U5562 (N_5562,N_4059,N_4307);
nand U5563 (N_5563,N_4529,N_4732);
nor U5564 (N_5564,N_4627,N_4670);
nand U5565 (N_5565,N_4596,N_4585);
or U5566 (N_5566,N_4260,N_4937);
or U5567 (N_5567,N_4863,N_4235);
or U5568 (N_5568,N_4185,N_4345);
or U5569 (N_5569,N_4459,N_4711);
xor U5570 (N_5570,N_4649,N_4494);
xor U5571 (N_5571,N_4183,N_4494);
nand U5572 (N_5572,N_4494,N_4218);
nor U5573 (N_5573,N_4515,N_4274);
and U5574 (N_5574,N_4418,N_4333);
or U5575 (N_5575,N_4900,N_4302);
xor U5576 (N_5576,N_4473,N_4752);
nand U5577 (N_5577,N_4458,N_4852);
or U5578 (N_5578,N_4917,N_4822);
xor U5579 (N_5579,N_4306,N_4089);
and U5580 (N_5580,N_4945,N_4121);
xnor U5581 (N_5581,N_4051,N_4614);
or U5582 (N_5582,N_4972,N_4019);
nor U5583 (N_5583,N_4250,N_4598);
and U5584 (N_5584,N_4095,N_4645);
nor U5585 (N_5585,N_4886,N_4667);
nor U5586 (N_5586,N_4270,N_4038);
and U5587 (N_5587,N_4278,N_4554);
or U5588 (N_5588,N_4457,N_4889);
and U5589 (N_5589,N_4726,N_4847);
and U5590 (N_5590,N_4164,N_4892);
or U5591 (N_5591,N_4021,N_4359);
or U5592 (N_5592,N_4025,N_4253);
xnor U5593 (N_5593,N_4214,N_4967);
nand U5594 (N_5594,N_4317,N_4501);
and U5595 (N_5595,N_4669,N_4684);
nor U5596 (N_5596,N_4854,N_4005);
and U5597 (N_5597,N_4290,N_4306);
nor U5598 (N_5598,N_4122,N_4673);
nor U5599 (N_5599,N_4729,N_4342);
xor U5600 (N_5600,N_4813,N_4879);
and U5601 (N_5601,N_4523,N_4255);
nor U5602 (N_5602,N_4658,N_4748);
and U5603 (N_5603,N_4263,N_4706);
or U5604 (N_5604,N_4448,N_4321);
or U5605 (N_5605,N_4790,N_4578);
or U5606 (N_5606,N_4396,N_4943);
or U5607 (N_5607,N_4619,N_4099);
nor U5608 (N_5608,N_4571,N_4058);
nand U5609 (N_5609,N_4571,N_4622);
or U5610 (N_5610,N_4413,N_4172);
or U5611 (N_5611,N_4287,N_4212);
nand U5612 (N_5612,N_4102,N_4379);
and U5613 (N_5613,N_4818,N_4670);
nor U5614 (N_5614,N_4509,N_4784);
xor U5615 (N_5615,N_4964,N_4191);
nand U5616 (N_5616,N_4622,N_4371);
or U5617 (N_5617,N_4340,N_4157);
and U5618 (N_5618,N_4598,N_4004);
nor U5619 (N_5619,N_4302,N_4148);
or U5620 (N_5620,N_4719,N_4226);
and U5621 (N_5621,N_4486,N_4852);
and U5622 (N_5622,N_4921,N_4866);
xnor U5623 (N_5623,N_4682,N_4977);
nor U5624 (N_5624,N_4653,N_4528);
and U5625 (N_5625,N_4935,N_4382);
xor U5626 (N_5626,N_4172,N_4840);
and U5627 (N_5627,N_4043,N_4549);
xor U5628 (N_5628,N_4792,N_4655);
or U5629 (N_5629,N_4382,N_4000);
and U5630 (N_5630,N_4241,N_4103);
nand U5631 (N_5631,N_4952,N_4605);
xor U5632 (N_5632,N_4292,N_4637);
xnor U5633 (N_5633,N_4086,N_4481);
xnor U5634 (N_5634,N_4958,N_4881);
nand U5635 (N_5635,N_4098,N_4961);
or U5636 (N_5636,N_4469,N_4737);
xor U5637 (N_5637,N_4083,N_4681);
nand U5638 (N_5638,N_4957,N_4511);
or U5639 (N_5639,N_4678,N_4488);
and U5640 (N_5640,N_4105,N_4183);
or U5641 (N_5641,N_4302,N_4051);
or U5642 (N_5642,N_4508,N_4282);
nand U5643 (N_5643,N_4526,N_4451);
xnor U5644 (N_5644,N_4026,N_4898);
nand U5645 (N_5645,N_4743,N_4386);
and U5646 (N_5646,N_4454,N_4732);
xnor U5647 (N_5647,N_4101,N_4702);
nor U5648 (N_5648,N_4811,N_4777);
xnor U5649 (N_5649,N_4518,N_4120);
and U5650 (N_5650,N_4039,N_4630);
or U5651 (N_5651,N_4056,N_4259);
or U5652 (N_5652,N_4106,N_4434);
nor U5653 (N_5653,N_4138,N_4197);
nor U5654 (N_5654,N_4078,N_4031);
xor U5655 (N_5655,N_4684,N_4545);
and U5656 (N_5656,N_4442,N_4209);
xor U5657 (N_5657,N_4040,N_4371);
nand U5658 (N_5658,N_4441,N_4804);
nand U5659 (N_5659,N_4310,N_4024);
or U5660 (N_5660,N_4666,N_4016);
or U5661 (N_5661,N_4974,N_4350);
nor U5662 (N_5662,N_4384,N_4316);
nand U5663 (N_5663,N_4958,N_4312);
nand U5664 (N_5664,N_4208,N_4391);
nand U5665 (N_5665,N_4543,N_4223);
or U5666 (N_5666,N_4528,N_4546);
nand U5667 (N_5667,N_4329,N_4904);
xnor U5668 (N_5668,N_4820,N_4798);
xor U5669 (N_5669,N_4873,N_4241);
or U5670 (N_5670,N_4675,N_4461);
or U5671 (N_5671,N_4458,N_4497);
nand U5672 (N_5672,N_4492,N_4484);
xnor U5673 (N_5673,N_4424,N_4606);
xor U5674 (N_5674,N_4056,N_4053);
xnor U5675 (N_5675,N_4877,N_4332);
or U5676 (N_5676,N_4163,N_4062);
xnor U5677 (N_5677,N_4635,N_4240);
or U5678 (N_5678,N_4480,N_4411);
nand U5679 (N_5679,N_4081,N_4855);
xnor U5680 (N_5680,N_4570,N_4415);
nand U5681 (N_5681,N_4052,N_4173);
xnor U5682 (N_5682,N_4412,N_4955);
nor U5683 (N_5683,N_4134,N_4882);
and U5684 (N_5684,N_4256,N_4304);
or U5685 (N_5685,N_4549,N_4576);
nor U5686 (N_5686,N_4001,N_4084);
and U5687 (N_5687,N_4846,N_4937);
or U5688 (N_5688,N_4853,N_4395);
and U5689 (N_5689,N_4836,N_4134);
nand U5690 (N_5690,N_4676,N_4674);
nor U5691 (N_5691,N_4239,N_4107);
and U5692 (N_5692,N_4434,N_4219);
nor U5693 (N_5693,N_4241,N_4332);
or U5694 (N_5694,N_4006,N_4219);
xnor U5695 (N_5695,N_4949,N_4718);
or U5696 (N_5696,N_4545,N_4535);
and U5697 (N_5697,N_4125,N_4657);
nor U5698 (N_5698,N_4019,N_4414);
xnor U5699 (N_5699,N_4153,N_4644);
nand U5700 (N_5700,N_4964,N_4842);
xnor U5701 (N_5701,N_4820,N_4746);
or U5702 (N_5702,N_4688,N_4990);
nor U5703 (N_5703,N_4283,N_4002);
nor U5704 (N_5704,N_4283,N_4261);
nand U5705 (N_5705,N_4562,N_4654);
or U5706 (N_5706,N_4456,N_4252);
or U5707 (N_5707,N_4302,N_4594);
nand U5708 (N_5708,N_4649,N_4293);
nor U5709 (N_5709,N_4839,N_4530);
and U5710 (N_5710,N_4132,N_4368);
nor U5711 (N_5711,N_4412,N_4419);
nand U5712 (N_5712,N_4071,N_4510);
nor U5713 (N_5713,N_4803,N_4832);
xnor U5714 (N_5714,N_4727,N_4817);
and U5715 (N_5715,N_4103,N_4391);
and U5716 (N_5716,N_4037,N_4455);
xor U5717 (N_5717,N_4935,N_4196);
nand U5718 (N_5718,N_4982,N_4456);
nand U5719 (N_5719,N_4292,N_4481);
or U5720 (N_5720,N_4840,N_4232);
nor U5721 (N_5721,N_4303,N_4156);
nand U5722 (N_5722,N_4630,N_4210);
nor U5723 (N_5723,N_4692,N_4091);
or U5724 (N_5724,N_4970,N_4137);
or U5725 (N_5725,N_4407,N_4097);
nor U5726 (N_5726,N_4183,N_4078);
nand U5727 (N_5727,N_4664,N_4454);
nand U5728 (N_5728,N_4666,N_4701);
and U5729 (N_5729,N_4974,N_4340);
or U5730 (N_5730,N_4143,N_4740);
and U5731 (N_5731,N_4859,N_4981);
or U5732 (N_5732,N_4940,N_4698);
and U5733 (N_5733,N_4458,N_4416);
xor U5734 (N_5734,N_4686,N_4538);
and U5735 (N_5735,N_4143,N_4529);
and U5736 (N_5736,N_4466,N_4425);
nor U5737 (N_5737,N_4745,N_4211);
or U5738 (N_5738,N_4821,N_4527);
xor U5739 (N_5739,N_4277,N_4030);
xor U5740 (N_5740,N_4248,N_4515);
xnor U5741 (N_5741,N_4667,N_4632);
nor U5742 (N_5742,N_4003,N_4831);
xnor U5743 (N_5743,N_4676,N_4781);
nor U5744 (N_5744,N_4918,N_4718);
or U5745 (N_5745,N_4674,N_4743);
nor U5746 (N_5746,N_4427,N_4172);
xnor U5747 (N_5747,N_4710,N_4844);
nand U5748 (N_5748,N_4768,N_4258);
xnor U5749 (N_5749,N_4222,N_4420);
nor U5750 (N_5750,N_4900,N_4478);
and U5751 (N_5751,N_4770,N_4769);
nor U5752 (N_5752,N_4267,N_4004);
and U5753 (N_5753,N_4400,N_4423);
xor U5754 (N_5754,N_4775,N_4420);
nand U5755 (N_5755,N_4086,N_4951);
and U5756 (N_5756,N_4289,N_4387);
or U5757 (N_5757,N_4538,N_4839);
nor U5758 (N_5758,N_4034,N_4011);
nand U5759 (N_5759,N_4269,N_4092);
nor U5760 (N_5760,N_4460,N_4953);
nor U5761 (N_5761,N_4383,N_4210);
nand U5762 (N_5762,N_4089,N_4123);
or U5763 (N_5763,N_4400,N_4861);
and U5764 (N_5764,N_4682,N_4181);
xnor U5765 (N_5765,N_4315,N_4856);
or U5766 (N_5766,N_4018,N_4614);
xnor U5767 (N_5767,N_4060,N_4229);
nand U5768 (N_5768,N_4489,N_4929);
xnor U5769 (N_5769,N_4164,N_4085);
and U5770 (N_5770,N_4067,N_4715);
and U5771 (N_5771,N_4636,N_4419);
nor U5772 (N_5772,N_4440,N_4246);
or U5773 (N_5773,N_4393,N_4860);
nor U5774 (N_5774,N_4682,N_4463);
or U5775 (N_5775,N_4052,N_4645);
and U5776 (N_5776,N_4538,N_4698);
nand U5777 (N_5777,N_4204,N_4610);
xnor U5778 (N_5778,N_4833,N_4943);
nand U5779 (N_5779,N_4498,N_4711);
xnor U5780 (N_5780,N_4292,N_4238);
or U5781 (N_5781,N_4304,N_4706);
or U5782 (N_5782,N_4758,N_4127);
nor U5783 (N_5783,N_4271,N_4938);
or U5784 (N_5784,N_4118,N_4921);
or U5785 (N_5785,N_4914,N_4453);
nor U5786 (N_5786,N_4049,N_4240);
nor U5787 (N_5787,N_4428,N_4398);
and U5788 (N_5788,N_4072,N_4300);
nand U5789 (N_5789,N_4382,N_4117);
nand U5790 (N_5790,N_4395,N_4344);
nand U5791 (N_5791,N_4211,N_4343);
and U5792 (N_5792,N_4791,N_4638);
xor U5793 (N_5793,N_4246,N_4861);
or U5794 (N_5794,N_4269,N_4798);
nor U5795 (N_5795,N_4338,N_4900);
nor U5796 (N_5796,N_4719,N_4599);
and U5797 (N_5797,N_4150,N_4957);
and U5798 (N_5798,N_4051,N_4104);
and U5799 (N_5799,N_4854,N_4573);
and U5800 (N_5800,N_4089,N_4589);
and U5801 (N_5801,N_4592,N_4578);
or U5802 (N_5802,N_4540,N_4042);
or U5803 (N_5803,N_4172,N_4589);
nand U5804 (N_5804,N_4940,N_4765);
nand U5805 (N_5805,N_4441,N_4812);
xor U5806 (N_5806,N_4785,N_4632);
xnor U5807 (N_5807,N_4247,N_4464);
xor U5808 (N_5808,N_4009,N_4846);
or U5809 (N_5809,N_4566,N_4088);
xor U5810 (N_5810,N_4892,N_4125);
or U5811 (N_5811,N_4104,N_4599);
nor U5812 (N_5812,N_4902,N_4724);
nor U5813 (N_5813,N_4913,N_4835);
and U5814 (N_5814,N_4663,N_4223);
and U5815 (N_5815,N_4721,N_4165);
and U5816 (N_5816,N_4306,N_4758);
xor U5817 (N_5817,N_4639,N_4721);
and U5818 (N_5818,N_4524,N_4545);
xnor U5819 (N_5819,N_4756,N_4475);
nor U5820 (N_5820,N_4060,N_4350);
or U5821 (N_5821,N_4532,N_4962);
nor U5822 (N_5822,N_4231,N_4127);
nand U5823 (N_5823,N_4452,N_4054);
and U5824 (N_5824,N_4229,N_4408);
or U5825 (N_5825,N_4224,N_4994);
nor U5826 (N_5826,N_4342,N_4497);
or U5827 (N_5827,N_4511,N_4063);
xor U5828 (N_5828,N_4887,N_4768);
nor U5829 (N_5829,N_4505,N_4022);
and U5830 (N_5830,N_4767,N_4307);
and U5831 (N_5831,N_4027,N_4061);
nor U5832 (N_5832,N_4106,N_4185);
and U5833 (N_5833,N_4761,N_4504);
and U5834 (N_5834,N_4301,N_4151);
nor U5835 (N_5835,N_4871,N_4975);
or U5836 (N_5836,N_4434,N_4129);
nor U5837 (N_5837,N_4562,N_4126);
and U5838 (N_5838,N_4727,N_4528);
and U5839 (N_5839,N_4451,N_4345);
or U5840 (N_5840,N_4884,N_4609);
and U5841 (N_5841,N_4320,N_4674);
xnor U5842 (N_5842,N_4334,N_4483);
nand U5843 (N_5843,N_4671,N_4127);
or U5844 (N_5844,N_4199,N_4015);
or U5845 (N_5845,N_4469,N_4691);
xor U5846 (N_5846,N_4581,N_4025);
nand U5847 (N_5847,N_4252,N_4692);
and U5848 (N_5848,N_4517,N_4882);
nor U5849 (N_5849,N_4334,N_4919);
and U5850 (N_5850,N_4361,N_4704);
and U5851 (N_5851,N_4258,N_4368);
nor U5852 (N_5852,N_4817,N_4679);
or U5853 (N_5853,N_4897,N_4638);
and U5854 (N_5854,N_4586,N_4112);
or U5855 (N_5855,N_4589,N_4757);
or U5856 (N_5856,N_4526,N_4900);
or U5857 (N_5857,N_4591,N_4157);
and U5858 (N_5858,N_4242,N_4236);
xnor U5859 (N_5859,N_4475,N_4155);
nor U5860 (N_5860,N_4698,N_4474);
xor U5861 (N_5861,N_4311,N_4595);
nand U5862 (N_5862,N_4377,N_4827);
nand U5863 (N_5863,N_4032,N_4829);
nand U5864 (N_5864,N_4929,N_4278);
xnor U5865 (N_5865,N_4344,N_4729);
xor U5866 (N_5866,N_4234,N_4888);
xnor U5867 (N_5867,N_4671,N_4332);
nand U5868 (N_5868,N_4544,N_4576);
nand U5869 (N_5869,N_4007,N_4160);
and U5870 (N_5870,N_4227,N_4867);
nor U5871 (N_5871,N_4613,N_4075);
and U5872 (N_5872,N_4455,N_4872);
xnor U5873 (N_5873,N_4218,N_4312);
nor U5874 (N_5874,N_4019,N_4891);
nor U5875 (N_5875,N_4567,N_4137);
nor U5876 (N_5876,N_4517,N_4262);
nor U5877 (N_5877,N_4581,N_4141);
and U5878 (N_5878,N_4682,N_4582);
and U5879 (N_5879,N_4396,N_4409);
and U5880 (N_5880,N_4870,N_4925);
or U5881 (N_5881,N_4829,N_4541);
nand U5882 (N_5882,N_4821,N_4675);
nor U5883 (N_5883,N_4880,N_4370);
nand U5884 (N_5884,N_4264,N_4343);
nand U5885 (N_5885,N_4827,N_4083);
nand U5886 (N_5886,N_4820,N_4243);
or U5887 (N_5887,N_4812,N_4970);
and U5888 (N_5888,N_4012,N_4257);
nand U5889 (N_5889,N_4674,N_4787);
nand U5890 (N_5890,N_4351,N_4113);
and U5891 (N_5891,N_4959,N_4577);
nand U5892 (N_5892,N_4553,N_4378);
xnor U5893 (N_5893,N_4723,N_4926);
nor U5894 (N_5894,N_4877,N_4520);
nand U5895 (N_5895,N_4961,N_4183);
xnor U5896 (N_5896,N_4693,N_4343);
nor U5897 (N_5897,N_4581,N_4279);
and U5898 (N_5898,N_4937,N_4010);
and U5899 (N_5899,N_4617,N_4206);
xnor U5900 (N_5900,N_4966,N_4920);
nor U5901 (N_5901,N_4942,N_4995);
nand U5902 (N_5902,N_4390,N_4118);
and U5903 (N_5903,N_4885,N_4065);
xnor U5904 (N_5904,N_4868,N_4134);
xnor U5905 (N_5905,N_4983,N_4198);
or U5906 (N_5906,N_4735,N_4012);
or U5907 (N_5907,N_4200,N_4146);
nor U5908 (N_5908,N_4560,N_4508);
nand U5909 (N_5909,N_4762,N_4846);
or U5910 (N_5910,N_4743,N_4402);
xor U5911 (N_5911,N_4625,N_4991);
nor U5912 (N_5912,N_4908,N_4726);
nor U5913 (N_5913,N_4571,N_4946);
xnor U5914 (N_5914,N_4074,N_4018);
or U5915 (N_5915,N_4488,N_4789);
or U5916 (N_5916,N_4196,N_4725);
nor U5917 (N_5917,N_4946,N_4766);
xor U5918 (N_5918,N_4004,N_4941);
xor U5919 (N_5919,N_4346,N_4542);
nand U5920 (N_5920,N_4911,N_4813);
and U5921 (N_5921,N_4200,N_4022);
or U5922 (N_5922,N_4579,N_4749);
xnor U5923 (N_5923,N_4604,N_4001);
or U5924 (N_5924,N_4097,N_4211);
or U5925 (N_5925,N_4877,N_4795);
nand U5926 (N_5926,N_4544,N_4223);
nor U5927 (N_5927,N_4892,N_4670);
nand U5928 (N_5928,N_4456,N_4640);
nand U5929 (N_5929,N_4222,N_4338);
or U5930 (N_5930,N_4020,N_4863);
or U5931 (N_5931,N_4573,N_4394);
or U5932 (N_5932,N_4881,N_4647);
nor U5933 (N_5933,N_4035,N_4658);
nor U5934 (N_5934,N_4566,N_4114);
nor U5935 (N_5935,N_4424,N_4664);
nand U5936 (N_5936,N_4422,N_4991);
and U5937 (N_5937,N_4143,N_4469);
and U5938 (N_5938,N_4720,N_4255);
xnor U5939 (N_5939,N_4839,N_4758);
and U5940 (N_5940,N_4733,N_4170);
nand U5941 (N_5941,N_4419,N_4714);
nor U5942 (N_5942,N_4984,N_4888);
nor U5943 (N_5943,N_4390,N_4116);
and U5944 (N_5944,N_4409,N_4341);
xor U5945 (N_5945,N_4873,N_4207);
or U5946 (N_5946,N_4617,N_4009);
or U5947 (N_5947,N_4752,N_4534);
xor U5948 (N_5948,N_4725,N_4114);
nor U5949 (N_5949,N_4016,N_4259);
xnor U5950 (N_5950,N_4785,N_4049);
or U5951 (N_5951,N_4036,N_4235);
nand U5952 (N_5952,N_4544,N_4652);
nand U5953 (N_5953,N_4558,N_4752);
nand U5954 (N_5954,N_4247,N_4434);
and U5955 (N_5955,N_4543,N_4813);
nand U5956 (N_5956,N_4808,N_4752);
xor U5957 (N_5957,N_4048,N_4339);
or U5958 (N_5958,N_4191,N_4912);
xor U5959 (N_5959,N_4857,N_4493);
or U5960 (N_5960,N_4474,N_4360);
or U5961 (N_5961,N_4217,N_4489);
nand U5962 (N_5962,N_4876,N_4371);
nand U5963 (N_5963,N_4622,N_4480);
nand U5964 (N_5964,N_4426,N_4332);
nor U5965 (N_5965,N_4949,N_4643);
and U5966 (N_5966,N_4190,N_4304);
or U5967 (N_5967,N_4568,N_4797);
and U5968 (N_5968,N_4679,N_4309);
nor U5969 (N_5969,N_4994,N_4506);
or U5970 (N_5970,N_4704,N_4454);
xor U5971 (N_5971,N_4434,N_4642);
xnor U5972 (N_5972,N_4049,N_4137);
nand U5973 (N_5973,N_4062,N_4965);
and U5974 (N_5974,N_4422,N_4252);
xor U5975 (N_5975,N_4626,N_4705);
xor U5976 (N_5976,N_4867,N_4364);
xor U5977 (N_5977,N_4281,N_4935);
or U5978 (N_5978,N_4767,N_4396);
or U5979 (N_5979,N_4303,N_4504);
nor U5980 (N_5980,N_4432,N_4570);
xor U5981 (N_5981,N_4705,N_4942);
or U5982 (N_5982,N_4187,N_4559);
xnor U5983 (N_5983,N_4037,N_4342);
xnor U5984 (N_5984,N_4961,N_4261);
nand U5985 (N_5985,N_4646,N_4167);
and U5986 (N_5986,N_4711,N_4977);
or U5987 (N_5987,N_4200,N_4452);
and U5988 (N_5988,N_4653,N_4802);
nor U5989 (N_5989,N_4934,N_4291);
and U5990 (N_5990,N_4632,N_4946);
nand U5991 (N_5991,N_4829,N_4483);
xor U5992 (N_5992,N_4066,N_4365);
nand U5993 (N_5993,N_4614,N_4015);
or U5994 (N_5994,N_4238,N_4342);
or U5995 (N_5995,N_4580,N_4212);
and U5996 (N_5996,N_4318,N_4575);
or U5997 (N_5997,N_4040,N_4964);
xor U5998 (N_5998,N_4830,N_4631);
and U5999 (N_5999,N_4795,N_4411);
xnor U6000 (N_6000,N_5667,N_5593);
or U6001 (N_6001,N_5163,N_5158);
and U6002 (N_6002,N_5495,N_5128);
xnor U6003 (N_6003,N_5179,N_5229);
or U6004 (N_6004,N_5866,N_5571);
or U6005 (N_6005,N_5724,N_5132);
and U6006 (N_6006,N_5883,N_5517);
and U6007 (N_6007,N_5116,N_5404);
xnor U6008 (N_6008,N_5335,N_5074);
and U6009 (N_6009,N_5527,N_5695);
and U6010 (N_6010,N_5015,N_5046);
or U6011 (N_6011,N_5783,N_5341);
xor U6012 (N_6012,N_5706,N_5945);
nand U6013 (N_6013,N_5786,N_5481);
nor U6014 (N_6014,N_5981,N_5394);
nand U6015 (N_6015,N_5955,N_5329);
nand U6016 (N_6016,N_5137,N_5662);
xor U6017 (N_6017,N_5871,N_5845);
nor U6018 (N_6018,N_5714,N_5071);
or U6019 (N_6019,N_5192,N_5644);
or U6020 (N_6020,N_5946,N_5185);
and U6021 (N_6021,N_5318,N_5916);
nand U6022 (N_6022,N_5687,N_5609);
and U6023 (N_6023,N_5770,N_5181);
nand U6024 (N_6024,N_5247,N_5225);
or U6025 (N_6025,N_5020,N_5756);
xor U6026 (N_6026,N_5001,N_5099);
nand U6027 (N_6027,N_5872,N_5171);
nand U6028 (N_6028,N_5103,N_5746);
nand U6029 (N_6029,N_5285,N_5196);
or U6030 (N_6030,N_5886,N_5450);
xor U6031 (N_6031,N_5135,N_5183);
nand U6032 (N_6032,N_5288,N_5791);
nand U6033 (N_6033,N_5009,N_5034);
xnor U6034 (N_6034,N_5856,N_5321);
nor U6035 (N_6035,N_5064,N_5650);
and U6036 (N_6036,N_5567,N_5283);
xnor U6037 (N_6037,N_5528,N_5828);
nand U6038 (N_6038,N_5852,N_5787);
nor U6039 (N_6039,N_5386,N_5210);
xnor U6040 (N_6040,N_5251,N_5459);
nor U6041 (N_6041,N_5173,N_5489);
or U6042 (N_6042,N_5053,N_5281);
nand U6043 (N_6043,N_5490,N_5387);
nand U6044 (N_6044,N_5168,N_5566);
xor U6045 (N_6045,N_5322,N_5758);
nand U6046 (N_6046,N_5118,N_5734);
nor U6047 (N_6047,N_5703,N_5606);
nand U6048 (N_6048,N_5529,N_5066);
xor U6049 (N_6049,N_5313,N_5747);
nor U6050 (N_6050,N_5563,N_5971);
and U6051 (N_6051,N_5487,N_5025);
or U6052 (N_6052,N_5467,N_5647);
nand U6053 (N_6053,N_5236,N_5078);
or U6054 (N_6054,N_5346,N_5767);
and U6055 (N_6055,N_5612,N_5337);
nand U6056 (N_6056,N_5095,N_5217);
and U6057 (N_6057,N_5154,N_5268);
nor U6058 (N_6058,N_5121,N_5351);
nor U6059 (N_6059,N_5499,N_5259);
xor U6060 (N_6060,N_5655,N_5514);
and U6061 (N_6061,N_5353,N_5441);
xnor U6062 (N_6062,N_5569,N_5968);
nand U6063 (N_6063,N_5545,N_5080);
or U6064 (N_6064,N_5142,N_5550);
nand U6065 (N_6065,N_5677,N_5083);
xnor U6066 (N_6066,N_5548,N_5925);
and U6067 (N_6067,N_5082,N_5839);
nand U6068 (N_6068,N_5426,N_5951);
nor U6069 (N_6069,N_5709,N_5397);
nor U6070 (N_6070,N_5508,N_5660);
nor U6071 (N_6071,N_5388,N_5543);
xor U6072 (N_6072,N_5933,N_5365);
xnor U6073 (N_6073,N_5019,N_5111);
nand U6074 (N_6074,N_5940,N_5881);
xnor U6075 (N_6075,N_5605,N_5950);
and U6076 (N_6076,N_5028,N_5223);
xor U6077 (N_6077,N_5284,N_5896);
or U6078 (N_6078,N_5598,N_5085);
nand U6079 (N_6079,N_5616,N_5840);
or U6080 (N_6080,N_5613,N_5357);
xnor U6081 (N_6081,N_5378,N_5350);
xnor U6082 (N_6082,N_5073,N_5018);
xor U6083 (N_6083,N_5802,N_5693);
nor U6084 (N_6084,N_5393,N_5782);
or U6085 (N_6085,N_5833,N_5238);
and U6086 (N_6086,N_5076,N_5013);
nor U6087 (N_6087,N_5948,N_5796);
nor U6088 (N_6088,N_5823,N_5043);
and U6089 (N_6089,N_5704,N_5162);
nand U6090 (N_6090,N_5184,N_5024);
nor U6091 (N_6091,N_5090,N_5546);
xor U6092 (N_6092,N_5474,N_5169);
nor U6093 (N_6093,N_5516,N_5800);
xor U6094 (N_6094,N_5718,N_5716);
xor U6095 (N_6095,N_5243,N_5539);
nand U6096 (N_6096,N_5822,N_5402);
nand U6097 (N_6097,N_5876,N_5141);
xor U6098 (N_6098,N_5319,N_5376);
or U6099 (N_6099,N_5072,N_5114);
nand U6100 (N_6100,N_5713,N_5698);
nor U6101 (N_6101,N_5045,N_5909);
nand U6102 (N_6102,N_5249,N_5984);
nor U6103 (N_6103,N_5148,N_5177);
and U6104 (N_6104,N_5811,N_5478);
nor U6105 (N_6105,N_5130,N_5765);
xnor U6106 (N_6106,N_5831,N_5577);
nand U6107 (N_6107,N_5873,N_5098);
nand U6108 (N_6108,N_5472,N_5809);
and U6109 (N_6109,N_5987,N_5501);
or U6110 (N_6110,N_5101,N_5728);
nor U6111 (N_6111,N_5875,N_5145);
xnor U6112 (N_6112,N_5473,N_5834);
xnor U6113 (N_6113,N_5070,N_5870);
xor U6114 (N_6114,N_5500,N_5776);
nand U6115 (N_6115,N_5937,N_5817);
xnor U6116 (N_6116,N_5764,N_5959);
and U6117 (N_6117,N_5956,N_5692);
or U6118 (N_6118,N_5115,N_5276);
nor U6119 (N_6119,N_5496,N_5794);
or U6120 (N_6120,N_5789,N_5637);
nor U6121 (N_6121,N_5576,N_5272);
xor U6122 (N_6122,N_5193,N_5112);
xor U6123 (N_6123,N_5861,N_5760);
nor U6124 (N_6124,N_5753,N_5970);
xnor U6125 (N_6125,N_5859,N_5869);
xor U6126 (N_6126,N_5000,N_5632);
nand U6127 (N_6127,N_5884,N_5924);
and U6128 (N_6128,N_5077,N_5614);
or U6129 (N_6129,N_5827,N_5656);
nor U6130 (N_6130,N_5907,N_5298);
nand U6131 (N_6131,N_5294,N_5156);
and U6132 (N_6132,N_5359,N_5688);
xor U6133 (N_6133,N_5301,N_5027);
nor U6134 (N_6134,N_5663,N_5425);
or U6135 (N_6135,N_5729,N_5842);
or U6136 (N_6136,N_5666,N_5668);
or U6137 (N_6137,N_5039,N_5400);
or U6138 (N_6138,N_5590,N_5140);
or U6139 (N_6139,N_5358,N_5736);
nor U6140 (N_6140,N_5458,N_5428);
nor U6141 (N_6141,N_5488,N_5067);
or U6142 (N_6142,N_5578,N_5557);
nand U6143 (N_6143,N_5362,N_5810);
nor U6144 (N_6144,N_5494,N_5645);
nor U6145 (N_6145,N_5580,N_5999);
nor U6146 (N_6146,N_5138,N_5235);
nor U6147 (N_6147,N_5819,N_5503);
xnor U6148 (N_6148,N_5248,N_5554);
nand U6149 (N_6149,N_5311,N_5586);
xnor U6150 (N_6150,N_5684,N_5306);
xor U6151 (N_6151,N_5913,N_5544);
or U6152 (N_6152,N_5844,N_5801);
nand U6153 (N_6153,N_5149,N_5087);
nor U6154 (N_6154,N_5038,N_5134);
or U6155 (N_6155,N_5370,N_5445);
xor U6156 (N_6156,N_5993,N_5058);
nand U6157 (N_6157,N_5265,N_5296);
and U6158 (N_6158,N_5424,N_5941);
nand U6159 (N_6159,N_5206,N_5929);
and U6160 (N_6160,N_5892,N_5300);
nor U6161 (N_6161,N_5205,N_5850);
or U6162 (N_6162,N_5750,N_5558);
nor U6163 (N_6163,N_5497,N_5126);
nand U6164 (N_6164,N_5146,N_5385);
and U6165 (N_6165,N_5965,N_5161);
and U6166 (N_6166,N_5914,N_5129);
nand U6167 (N_6167,N_5537,N_5615);
xnor U6168 (N_6168,N_5832,N_5017);
nand U6169 (N_6169,N_5390,N_5178);
xnor U6170 (N_6170,N_5412,N_5730);
and U6171 (N_6171,N_5690,N_5841);
nor U6172 (N_6172,N_5403,N_5150);
or U6173 (N_6173,N_5047,N_5254);
xnor U6174 (N_6174,N_5986,N_5224);
nand U6175 (N_6175,N_5199,N_5939);
or U6176 (N_6176,N_5702,N_5990);
nor U6177 (N_6177,N_5255,N_5621);
nand U6178 (N_6178,N_5638,N_5451);
and U6179 (N_6179,N_5799,N_5815);
and U6180 (N_6180,N_5784,N_5044);
nor U6181 (N_6181,N_5938,N_5919);
nor U6182 (N_6182,N_5752,N_5669);
nor U6183 (N_6183,N_5356,N_5820);
nor U6184 (N_6184,N_5538,N_5379);
nand U6185 (N_6185,N_5519,N_5816);
nor U6186 (N_6186,N_5777,N_5627);
nand U6187 (N_6187,N_5918,N_5654);
nor U6188 (N_6188,N_5417,N_5882);
nand U6189 (N_6189,N_5065,N_5050);
xnor U6190 (N_6190,N_5530,N_5194);
or U6191 (N_6191,N_5848,N_5700);
or U6192 (N_6192,N_5125,N_5769);
nor U6193 (N_6193,N_5710,N_5504);
nor U6194 (N_6194,N_5853,N_5635);
nor U6195 (N_6195,N_5587,N_5333);
nand U6196 (N_6196,N_5057,N_5512);
xnor U6197 (N_6197,N_5723,N_5160);
or U6198 (N_6198,N_5405,N_5464);
and U6199 (N_6199,N_5905,N_5542);
nor U6200 (N_6200,N_5106,N_5340);
nand U6201 (N_6201,N_5060,N_5282);
xor U6202 (N_6202,N_5680,N_5336);
nand U6203 (N_6203,N_5779,N_5269);
nand U6204 (N_6204,N_5409,N_5360);
and U6205 (N_6205,N_5485,N_5751);
or U6206 (N_6206,N_5222,N_5200);
xor U6207 (N_6207,N_5920,N_5596);
and U6208 (N_6208,N_5286,N_5936);
or U6209 (N_6209,N_5022,N_5204);
nand U6210 (N_6210,N_5665,N_5415);
or U6211 (N_6211,N_5055,N_5903);
nor U6212 (N_6212,N_5302,N_5910);
nor U6213 (N_6213,N_5643,N_5438);
nand U6214 (N_6214,N_5731,N_5960);
nand U6215 (N_6215,N_5541,N_5825);
xor U6216 (N_6216,N_5420,N_5442);
or U6217 (N_6217,N_5582,N_5030);
nand U6218 (N_6218,N_5182,N_5594);
xnor U6219 (N_6219,N_5785,N_5565);
nand U6220 (N_6220,N_5628,N_5476);
or U6221 (N_6221,N_5626,N_5392);
or U6222 (N_6222,N_5143,N_5293);
and U6223 (N_6223,N_5398,N_5682);
xnor U6224 (N_6224,N_5326,N_5380);
nand U6225 (N_6225,N_5317,N_5835);
or U6226 (N_6226,N_5649,N_5620);
xnor U6227 (N_6227,N_5423,N_5898);
xor U6228 (N_6228,N_5401,N_5513);
xnor U6229 (N_6229,N_5049,N_5868);
nor U6230 (N_6230,N_5717,N_5007);
or U6231 (N_6231,N_5836,N_5911);
and U6232 (N_6232,N_5893,N_5465);
nand U6233 (N_6233,N_5585,N_5763);
xor U6234 (N_6234,N_5051,N_5091);
xor U6235 (N_6235,N_5562,N_5005);
xnor U6236 (N_6236,N_5610,N_5089);
nor U6237 (N_6237,N_5821,N_5479);
xor U6238 (N_6238,N_5625,N_5954);
xnor U6239 (N_6239,N_5408,N_5372);
nor U6240 (N_6240,N_5958,N_5540);
nor U6241 (N_6241,N_5446,N_5737);
nor U6242 (N_6242,N_5081,N_5659);
xor U6243 (N_6243,N_5202,N_5855);
or U6244 (N_6244,N_5227,N_5452);
or U6245 (N_6245,N_5382,N_5773);
and U6246 (N_6246,N_5712,N_5310);
nand U6247 (N_6247,N_5579,N_5052);
nand U6248 (N_6248,N_5602,N_5040);
nor U6249 (N_6249,N_5444,N_5862);
xnor U6250 (N_6250,N_5768,N_5331);
xnor U6251 (N_6251,N_5124,N_5026);
and U6252 (N_6252,N_5917,N_5031);
nand U6253 (N_6253,N_5147,N_5309);
nand U6254 (N_6254,N_5953,N_5167);
xnor U6255 (N_6255,N_5744,N_5165);
nor U6256 (N_6256,N_5630,N_5691);
nor U6257 (N_6257,N_5701,N_5011);
and U6258 (N_6258,N_5983,N_5355);
or U6259 (N_6259,N_5498,N_5857);
xnor U6260 (N_6260,N_5526,N_5430);
and U6261 (N_6261,N_5292,N_5215);
xnor U6262 (N_6262,N_5486,N_5096);
and U6263 (N_6263,N_5339,N_5589);
or U6264 (N_6264,N_5988,N_5934);
or U6265 (N_6265,N_5699,N_5837);
xnor U6266 (N_6266,N_5119,N_5257);
nand U6267 (N_6267,N_5048,N_5727);
or U6268 (N_6268,N_5600,N_5639);
xor U6269 (N_6269,N_5029,N_5108);
or U6270 (N_6270,N_5922,N_5696);
nor U6271 (N_6271,N_5136,N_5509);
or U6272 (N_6272,N_5421,N_5399);
or U6273 (N_6273,N_5375,N_5766);
xor U6274 (N_6274,N_5814,N_5685);
and U6275 (N_6275,N_5812,N_5012);
and U6276 (N_6276,N_5641,N_5942);
xor U6277 (N_6277,N_5406,N_5931);
nand U6278 (N_6278,N_5757,N_5505);
or U6279 (N_6279,N_5260,N_5511);
xor U6280 (N_6280,N_5961,N_5962);
or U6281 (N_6281,N_5188,N_5172);
xnor U6282 (N_6282,N_5732,N_5493);
nor U6283 (N_6283,N_5761,N_5440);
or U6284 (N_6284,N_5720,N_5407);
nor U6285 (N_6285,N_5228,N_5510);
nor U6286 (N_6286,N_5633,N_5996);
xnor U6287 (N_6287,N_5413,N_5422);
nor U6288 (N_6288,N_5595,N_5435);
xnor U6289 (N_6289,N_5664,N_5573);
or U6290 (N_6290,N_5245,N_5369);
or U6291 (N_6291,N_5155,N_5477);
xnor U6292 (N_6292,N_5952,N_5622);
and U6293 (N_6293,N_5036,N_5016);
and U6294 (N_6294,N_5743,N_5471);
and U6295 (N_6295,N_5267,N_5711);
or U6296 (N_6296,N_5297,N_5256);
xnor U6297 (N_6297,N_5033,N_5439);
nand U6298 (N_6298,N_5583,N_5847);
nand U6299 (N_6299,N_5470,N_5570);
nand U6300 (N_6300,N_5396,N_5266);
nor U6301 (N_6301,N_5325,N_5127);
xor U6302 (N_6302,N_5042,N_5623);
nand U6303 (N_6303,N_5998,N_5246);
and U6304 (N_6304,N_5521,N_5880);
or U6305 (N_6305,N_5679,N_5271);
and U6306 (N_6306,N_5455,N_5793);
and U6307 (N_6307,N_5564,N_5790);
nand U6308 (N_6308,N_5233,N_5584);
nor U6309 (N_6309,N_5874,N_5806);
and U6310 (N_6310,N_5715,N_5234);
xnor U6311 (N_6311,N_5877,N_5109);
nand U6312 (N_6312,N_5289,N_5492);
and U6313 (N_6313,N_5930,N_5175);
nor U6314 (N_6314,N_5006,N_5556);
and U6315 (N_6315,N_5061,N_5902);
or U6316 (N_6316,N_5308,N_5969);
xnor U6317 (N_6317,N_5002,N_5642);
or U6318 (N_6318,N_5383,N_5277);
and U6319 (N_6319,N_5197,N_5588);
nor U6320 (N_6320,N_5159,N_5021);
nand U6321 (N_6321,N_5522,N_5239);
or U6322 (N_6322,N_5927,N_5186);
nor U6323 (N_6323,N_5591,N_5389);
and U6324 (N_6324,N_5547,N_5648);
or U6325 (N_6325,N_5220,N_5772);
nand U6326 (N_6326,N_5462,N_5434);
and U6327 (N_6327,N_5858,N_5536);
or U6328 (N_6328,N_5332,N_5552);
and U6329 (N_6329,N_5232,N_5176);
and U6330 (N_6330,N_5252,N_5218);
xnor U6331 (N_6331,N_5797,N_5304);
xor U6332 (N_6332,N_5807,N_5629);
or U6333 (N_6333,N_5480,N_5117);
nor U6334 (N_6334,N_5363,N_5972);
nand U6335 (N_6335,N_5974,N_5740);
and U6336 (N_6336,N_5231,N_5448);
and U6337 (N_6337,N_5944,N_5323);
nor U6338 (N_6338,N_5263,N_5592);
xnor U6339 (N_6339,N_5100,N_5475);
or U6340 (N_6340,N_5461,N_5781);
xnor U6341 (N_6341,N_5299,N_5418);
or U6342 (N_6342,N_5991,N_5104);
or U6343 (N_6343,N_5195,N_5980);
xor U6344 (N_6344,N_5830,N_5719);
or U6345 (N_6345,N_5994,N_5123);
nor U6346 (N_6346,N_5646,N_5603);
xor U6347 (N_6347,N_5997,N_5068);
or U6348 (N_6348,N_5771,N_5352);
nand U6349 (N_6349,N_5004,N_5805);
nand U6350 (N_6350,N_5273,N_5110);
or U6351 (N_6351,N_5242,N_5617);
and U6352 (N_6352,N_5608,N_5755);
nor U6353 (N_6353,N_5599,N_5581);
and U6354 (N_6354,N_5979,N_5678);
nor U6355 (N_6355,N_5240,N_5560);
nor U6356 (N_6356,N_5561,N_5967);
or U6357 (N_6357,N_5604,N_5675);
or U6358 (N_6358,N_5469,N_5894);
nor U6359 (N_6359,N_5804,N_5921);
or U6360 (N_6360,N_5741,N_5468);
or U6361 (N_6361,N_5555,N_5391);
nand U6362 (N_6362,N_5144,N_5084);
xor U6363 (N_6363,N_5947,N_5483);
and U6364 (N_6364,N_5964,N_5164);
nand U6365 (N_6365,N_5774,N_5201);
or U6366 (N_6366,N_5244,N_5694);
and U6367 (N_6367,N_5384,N_5525);
xnor U6368 (N_6368,N_5749,N_5673);
or U6369 (N_6369,N_5926,N_5611);
nand U6370 (N_6370,N_5287,N_5631);
or U6371 (N_6371,N_5433,N_5374);
nand U6372 (N_6372,N_5443,N_5535);
xor U6373 (N_6373,N_5216,N_5312);
xor U6374 (N_6374,N_5891,N_5803);
nand U6375 (N_6375,N_5726,N_5551);
xnor U6376 (N_6376,N_5533,N_5037);
and U6377 (N_6377,N_5102,N_5686);
and U6378 (N_6378,N_5963,N_5278);
nor U6379 (N_6379,N_5976,N_5191);
or U6380 (N_6380,N_5212,N_5985);
or U6381 (N_6381,N_5733,N_5657);
nand U6382 (N_6382,N_5754,N_5854);
xnor U6383 (N_6383,N_5069,N_5088);
nand U6384 (N_6384,N_5214,N_5906);
nand U6385 (N_6385,N_5345,N_5279);
and U6386 (N_6386,N_5867,N_5314);
nand U6387 (N_6387,N_5447,N_5054);
nor U6388 (N_6388,N_5411,N_5338);
nor U6389 (N_6389,N_5008,N_5105);
and U6390 (N_6390,N_5887,N_5762);
nor U6391 (N_6391,N_5334,N_5303);
nor U6392 (N_6392,N_5966,N_5658);
nand U6393 (N_6393,N_5895,N_5977);
xor U6394 (N_6394,N_5328,N_5863);
nand U6395 (N_6395,N_5721,N_5207);
nand U6396 (N_6396,N_5253,N_5568);
and U6397 (N_6397,N_5775,N_5932);
and U6398 (N_6398,N_5463,N_5315);
nand U6399 (N_6399,N_5506,N_5671);
or U6400 (N_6400,N_5366,N_5572);
and U6401 (N_6401,N_5739,N_5575);
xor U6402 (N_6402,N_5349,N_5824);
nor U6403 (N_6403,N_5532,N_5923);
xor U6404 (N_6404,N_5189,N_5466);
nand U6405 (N_6405,N_5707,N_5416);
and U6406 (N_6406,N_5305,N_5187);
nand U6407 (N_6407,N_5992,N_5838);
nor U6408 (N_6408,N_5410,N_5949);
xor U6409 (N_6409,N_5888,N_5460);
xor U6410 (N_6410,N_5262,N_5371);
nand U6411 (N_6411,N_5209,N_5957);
xor U6412 (N_6412,N_5221,N_5899);
and U6413 (N_6413,N_5208,N_5075);
or U6414 (N_6414,N_5131,N_5975);
xnor U6415 (N_6415,N_5414,N_5618);
nand U6416 (N_6416,N_5324,N_5274);
nor U6417 (N_6417,N_5377,N_5062);
xnor U6418 (N_6418,N_5735,N_5203);
and U6419 (N_6419,N_5327,N_5995);
xor U6420 (N_6420,N_5748,N_5361);
nand U6421 (N_6421,N_5901,N_5978);
xnor U6422 (N_6422,N_5436,N_5652);
xnor U6423 (N_6423,N_5818,N_5056);
xnor U6424 (N_6424,N_5190,N_5041);
or U6425 (N_6425,N_5381,N_5093);
or U6426 (N_6426,N_5674,N_5014);
and U6427 (N_6427,N_5122,N_5373);
and U6428 (N_6428,N_5482,N_5086);
nor U6429 (N_6429,N_5226,N_5943);
nand U6430 (N_6430,N_5549,N_5502);
and U6431 (N_6431,N_5230,N_5063);
nor U6432 (N_6432,N_5531,N_5250);
or U6433 (N_6433,N_5454,N_5559);
xor U6434 (N_6434,N_5097,N_5270);
nand U6435 (N_6435,N_5291,N_5010);
nor U6436 (N_6436,N_5973,N_5798);
or U6437 (N_6437,N_5860,N_5431);
or U6438 (N_6438,N_5885,N_5574);
nand U6439 (N_6439,N_5864,N_5170);
and U6440 (N_6440,N_5427,N_5237);
and U6441 (N_6441,N_5808,N_5367);
xnor U6442 (N_6442,N_5368,N_5553);
xor U6443 (N_6443,N_5534,N_5795);
nor U6444 (N_6444,N_5681,N_5219);
xnor U6445 (N_6445,N_5059,N_5879);
xnor U6446 (N_6446,N_5788,N_5343);
and U6447 (N_6447,N_5738,N_5989);
and U6448 (N_6448,N_5395,N_5107);
or U6449 (N_6449,N_5636,N_5619);
nor U6450 (N_6450,N_5023,N_5697);
or U6451 (N_6451,N_5601,N_5035);
or U6452 (N_6452,N_5151,N_5889);
nand U6453 (N_6453,N_5851,N_5829);
and U6454 (N_6454,N_5912,N_5928);
nand U6455 (N_6455,N_5597,N_5344);
nor U6456 (N_6456,N_5354,N_5742);
and U6457 (N_6457,N_5213,N_5676);
xnor U6458 (N_6458,N_5826,N_5153);
or U6459 (N_6459,N_5507,N_5518);
or U6460 (N_6460,N_5520,N_5330);
nand U6461 (N_6461,N_5429,N_5113);
and U6462 (N_6462,N_5180,N_5152);
or U6463 (N_6463,N_5897,N_5491);
xor U6464 (N_6464,N_5032,N_5419);
or U6465 (N_6465,N_5935,N_5515);
and U6466 (N_6466,N_5157,N_5780);
nand U6467 (N_6467,N_5258,N_5843);
nor U6468 (N_6468,N_5900,N_5449);
nor U6469 (N_6469,N_5722,N_5275);
or U6470 (N_6470,N_5437,N_5280);
or U6471 (N_6471,N_5348,N_5725);
or U6472 (N_6472,N_5264,N_5261);
xor U6473 (N_6473,N_5890,N_5290);
or U6474 (N_6474,N_5689,N_5670);
nand U6475 (N_6475,N_5982,N_5320);
nand U6476 (N_6476,N_5166,N_5661);
or U6477 (N_6477,N_5484,N_5456);
or U6478 (N_6478,N_5432,N_5705);
nand U6479 (N_6479,N_5342,N_5457);
xnor U6480 (N_6480,N_5092,N_5120);
nand U6481 (N_6481,N_5878,N_5865);
nor U6482 (N_6482,N_5524,N_5792);
nand U6483 (N_6483,N_5778,N_5849);
xnor U6484 (N_6484,N_5003,N_5094);
nand U6485 (N_6485,N_5634,N_5813);
nand U6486 (N_6486,N_5523,N_5453);
or U6487 (N_6487,N_5607,N_5174);
or U6488 (N_6488,N_5651,N_5624);
nor U6489 (N_6489,N_5079,N_5295);
nand U6490 (N_6490,N_5347,N_5683);
xor U6491 (N_6491,N_5139,N_5307);
and U6492 (N_6492,N_5904,N_5708);
and U6493 (N_6493,N_5915,N_5653);
and U6494 (N_6494,N_5759,N_5241);
nand U6495 (N_6495,N_5364,N_5908);
xor U6496 (N_6496,N_5745,N_5133);
nor U6497 (N_6497,N_5846,N_5316);
and U6498 (N_6498,N_5198,N_5211);
nor U6499 (N_6499,N_5672,N_5640);
xnor U6500 (N_6500,N_5308,N_5083);
or U6501 (N_6501,N_5087,N_5958);
or U6502 (N_6502,N_5130,N_5613);
xor U6503 (N_6503,N_5177,N_5678);
xor U6504 (N_6504,N_5974,N_5860);
nand U6505 (N_6505,N_5495,N_5182);
and U6506 (N_6506,N_5534,N_5098);
nand U6507 (N_6507,N_5718,N_5263);
xnor U6508 (N_6508,N_5150,N_5081);
nand U6509 (N_6509,N_5158,N_5120);
or U6510 (N_6510,N_5718,N_5192);
or U6511 (N_6511,N_5628,N_5104);
and U6512 (N_6512,N_5890,N_5316);
or U6513 (N_6513,N_5148,N_5275);
xnor U6514 (N_6514,N_5850,N_5902);
nor U6515 (N_6515,N_5371,N_5422);
or U6516 (N_6516,N_5050,N_5120);
nor U6517 (N_6517,N_5381,N_5034);
nor U6518 (N_6518,N_5929,N_5885);
xor U6519 (N_6519,N_5238,N_5204);
or U6520 (N_6520,N_5931,N_5567);
and U6521 (N_6521,N_5427,N_5101);
nand U6522 (N_6522,N_5019,N_5713);
or U6523 (N_6523,N_5624,N_5799);
xnor U6524 (N_6524,N_5039,N_5940);
nand U6525 (N_6525,N_5601,N_5534);
nand U6526 (N_6526,N_5065,N_5302);
xor U6527 (N_6527,N_5134,N_5293);
or U6528 (N_6528,N_5639,N_5748);
or U6529 (N_6529,N_5362,N_5496);
or U6530 (N_6530,N_5668,N_5286);
nand U6531 (N_6531,N_5980,N_5148);
xor U6532 (N_6532,N_5994,N_5536);
and U6533 (N_6533,N_5091,N_5744);
xnor U6534 (N_6534,N_5235,N_5432);
or U6535 (N_6535,N_5846,N_5272);
nand U6536 (N_6536,N_5120,N_5400);
nor U6537 (N_6537,N_5531,N_5657);
and U6538 (N_6538,N_5978,N_5923);
xor U6539 (N_6539,N_5894,N_5144);
xnor U6540 (N_6540,N_5499,N_5887);
and U6541 (N_6541,N_5670,N_5930);
nand U6542 (N_6542,N_5338,N_5073);
xor U6543 (N_6543,N_5606,N_5563);
and U6544 (N_6544,N_5486,N_5767);
nor U6545 (N_6545,N_5423,N_5310);
xor U6546 (N_6546,N_5171,N_5198);
xor U6547 (N_6547,N_5642,N_5244);
nor U6548 (N_6548,N_5100,N_5072);
and U6549 (N_6549,N_5868,N_5705);
and U6550 (N_6550,N_5227,N_5133);
xor U6551 (N_6551,N_5091,N_5965);
nand U6552 (N_6552,N_5753,N_5181);
and U6553 (N_6553,N_5936,N_5932);
xnor U6554 (N_6554,N_5148,N_5006);
xnor U6555 (N_6555,N_5394,N_5127);
or U6556 (N_6556,N_5889,N_5672);
nor U6557 (N_6557,N_5853,N_5375);
nor U6558 (N_6558,N_5647,N_5817);
and U6559 (N_6559,N_5873,N_5042);
nand U6560 (N_6560,N_5274,N_5086);
nor U6561 (N_6561,N_5850,N_5271);
nand U6562 (N_6562,N_5409,N_5946);
xor U6563 (N_6563,N_5191,N_5658);
or U6564 (N_6564,N_5508,N_5000);
nand U6565 (N_6565,N_5269,N_5735);
nor U6566 (N_6566,N_5636,N_5478);
or U6567 (N_6567,N_5210,N_5486);
and U6568 (N_6568,N_5133,N_5678);
nor U6569 (N_6569,N_5049,N_5407);
nor U6570 (N_6570,N_5967,N_5265);
or U6571 (N_6571,N_5494,N_5614);
nor U6572 (N_6572,N_5831,N_5152);
and U6573 (N_6573,N_5933,N_5037);
or U6574 (N_6574,N_5020,N_5152);
and U6575 (N_6575,N_5370,N_5839);
xnor U6576 (N_6576,N_5825,N_5535);
xnor U6577 (N_6577,N_5546,N_5821);
and U6578 (N_6578,N_5579,N_5110);
or U6579 (N_6579,N_5691,N_5684);
or U6580 (N_6580,N_5581,N_5694);
nand U6581 (N_6581,N_5759,N_5991);
and U6582 (N_6582,N_5276,N_5153);
and U6583 (N_6583,N_5187,N_5189);
xor U6584 (N_6584,N_5514,N_5935);
or U6585 (N_6585,N_5225,N_5407);
xor U6586 (N_6586,N_5627,N_5071);
nand U6587 (N_6587,N_5176,N_5677);
or U6588 (N_6588,N_5855,N_5119);
and U6589 (N_6589,N_5904,N_5966);
and U6590 (N_6590,N_5882,N_5068);
nor U6591 (N_6591,N_5968,N_5536);
or U6592 (N_6592,N_5849,N_5418);
nand U6593 (N_6593,N_5480,N_5050);
nor U6594 (N_6594,N_5885,N_5740);
nor U6595 (N_6595,N_5421,N_5422);
and U6596 (N_6596,N_5662,N_5116);
xor U6597 (N_6597,N_5557,N_5918);
nand U6598 (N_6598,N_5300,N_5574);
xnor U6599 (N_6599,N_5246,N_5745);
nor U6600 (N_6600,N_5764,N_5534);
nor U6601 (N_6601,N_5370,N_5451);
or U6602 (N_6602,N_5473,N_5359);
nand U6603 (N_6603,N_5888,N_5635);
xnor U6604 (N_6604,N_5559,N_5172);
nand U6605 (N_6605,N_5853,N_5446);
nand U6606 (N_6606,N_5283,N_5653);
xor U6607 (N_6607,N_5400,N_5460);
nand U6608 (N_6608,N_5048,N_5887);
or U6609 (N_6609,N_5017,N_5526);
nor U6610 (N_6610,N_5467,N_5040);
xnor U6611 (N_6611,N_5852,N_5310);
or U6612 (N_6612,N_5720,N_5580);
or U6613 (N_6613,N_5981,N_5504);
nor U6614 (N_6614,N_5306,N_5633);
xnor U6615 (N_6615,N_5427,N_5587);
nand U6616 (N_6616,N_5950,N_5806);
nand U6617 (N_6617,N_5482,N_5796);
nand U6618 (N_6618,N_5957,N_5533);
nor U6619 (N_6619,N_5556,N_5313);
and U6620 (N_6620,N_5029,N_5618);
or U6621 (N_6621,N_5667,N_5072);
and U6622 (N_6622,N_5124,N_5817);
nand U6623 (N_6623,N_5549,N_5320);
and U6624 (N_6624,N_5802,N_5342);
and U6625 (N_6625,N_5392,N_5636);
nand U6626 (N_6626,N_5382,N_5133);
nand U6627 (N_6627,N_5616,N_5807);
nand U6628 (N_6628,N_5372,N_5963);
xnor U6629 (N_6629,N_5533,N_5833);
and U6630 (N_6630,N_5731,N_5573);
nand U6631 (N_6631,N_5916,N_5602);
and U6632 (N_6632,N_5460,N_5896);
nand U6633 (N_6633,N_5185,N_5134);
nand U6634 (N_6634,N_5480,N_5593);
or U6635 (N_6635,N_5259,N_5849);
and U6636 (N_6636,N_5574,N_5426);
and U6637 (N_6637,N_5687,N_5863);
xnor U6638 (N_6638,N_5370,N_5000);
or U6639 (N_6639,N_5484,N_5412);
xor U6640 (N_6640,N_5465,N_5117);
or U6641 (N_6641,N_5904,N_5003);
or U6642 (N_6642,N_5091,N_5793);
nor U6643 (N_6643,N_5316,N_5712);
xor U6644 (N_6644,N_5452,N_5556);
nand U6645 (N_6645,N_5039,N_5683);
or U6646 (N_6646,N_5660,N_5639);
nor U6647 (N_6647,N_5598,N_5727);
nor U6648 (N_6648,N_5367,N_5829);
nand U6649 (N_6649,N_5629,N_5030);
xor U6650 (N_6650,N_5225,N_5766);
nand U6651 (N_6651,N_5716,N_5708);
nor U6652 (N_6652,N_5093,N_5505);
and U6653 (N_6653,N_5721,N_5205);
or U6654 (N_6654,N_5163,N_5625);
nor U6655 (N_6655,N_5710,N_5304);
and U6656 (N_6656,N_5187,N_5310);
and U6657 (N_6657,N_5233,N_5087);
and U6658 (N_6658,N_5342,N_5960);
and U6659 (N_6659,N_5448,N_5759);
xnor U6660 (N_6660,N_5210,N_5563);
nor U6661 (N_6661,N_5902,N_5220);
xor U6662 (N_6662,N_5978,N_5200);
and U6663 (N_6663,N_5370,N_5662);
and U6664 (N_6664,N_5216,N_5092);
and U6665 (N_6665,N_5173,N_5046);
xnor U6666 (N_6666,N_5452,N_5116);
and U6667 (N_6667,N_5519,N_5135);
nor U6668 (N_6668,N_5368,N_5092);
xor U6669 (N_6669,N_5884,N_5911);
nor U6670 (N_6670,N_5458,N_5133);
nand U6671 (N_6671,N_5532,N_5336);
or U6672 (N_6672,N_5269,N_5086);
xor U6673 (N_6673,N_5030,N_5945);
xnor U6674 (N_6674,N_5617,N_5676);
and U6675 (N_6675,N_5382,N_5801);
and U6676 (N_6676,N_5926,N_5638);
xnor U6677 (N_6677,N_5890,N_5142);
and U6678 (N_6678,N_5585,N_5941);
and U6679 (N_6679,N_5836,N_5326);
nor U6680 (N_6680,N_5569,N_5119);
or U6681 (N_6681,N_5242,N_5208);
xnor U6682 (N_6682,N_5595,N_5305);
nand U6683 (N_6683,N_5216,N_5808);
nor U6684 (N_6684,N_5153,N_5849);
xnor U6685 (N_6685,N_5531,N_5016);
and U6686 (N_6686,N_5227,N_5484);
nor U6687 (N_6687,N_5988,N_5625);
nor U6688 (N_6688,N_5291,N_5053);
xnor U6689 (N_6689,N_5877,N_5667);
nand U6690 (N_6690,N_5384,N_5625);
nor U6691 (N_6691,N_5401,N_5018);
nor U6692 (N_6692,N_5169,N_5945);
nor U6693 (N_6693,N_5155,N_5168);
xor U6694 (N_6694,N_5266,N_5879);
nor U6695 (N_6695,N_5400,N_5713);
nor U6696 (N_6696,N_5357,N_5652);
xnor U6697 (N_6697,N_5229,N_5942);
nand U6698 (N_6698,N_5844,N_5247);
xor U6699 (N_6699,N_5089,N_5414);
or U6700 (N_6700,N_5536,N_5956);
xor U6701 (N_6701,N_5213,N_5211);
or U6702 (N_6702,N_5103,N_5017);
nor U6703 (N_6703,N_5523,N_5497);
or U6704 (N_6704,N_5596,N_5533);
or U6705 (N_6705,N_5924,N_5262);
nor U6706 (N_6706,N_5790,N_5450);
nand U6707 (N_6707,N_5614,N_5504);
xnor U6708 (N_6708,N_5805,N_5659);
nor U6709 (N_6709,N_5112,N_5063);
or U6710 (N_6710,N_5249,N_5967);
or U6711 (N_6711,N_5906,N_5604);
and U6712 (N_6712,N_5620,N_5194);
or U6713 (N_6713,N_5288,N_5043);
nand U6714 (N_6714,N_5218,N_5729);
xor U6715 (N_6715,N_5972,N_5973);
xor U6716 (N_6716,N_5112,N_5350);
xnor U6717 (N_6717,N_5923,N_5549);
or U6718 (N_6718,N_5654,N_5292);
nand U6719 (N_6719,N_5795,N_5013);
nand U6720 (N_6720,N_5523,N_5787);
nand U6721 (N_6721,N_5656,N_5398);
nor U6722 (N_6722,N_5079,N_5085);
nor U6723 (N_6723,N_5593,N_5529);
xor U6724 (N_6724,N_5602,N_5064);
nor U6725 (N_6725,N_5294,N_5384);
nand U6726 (N_6726,N_5848,N_5353);
xnor U6727 (N_6727,N_5760,N_5463);
xor U6728 (N_6728,N_5695,N_5276);
nor U6729 (N_6729,N_5762,N_5655);
and U6730 (N_6730,N_5032,N_5099);
nand U6731 (N_6731,N_5381,N_5595);
or U6732 (N_6732,N_5653,N_5450);
and U6733 (N_6733,N_5902,N_5458);
xor U6734 (N_6734,N_5071,N_5128);
xnor U6735 (N_6735,N_5542,N_5710);
and U6736 (N_6736,N_5229,N_5364);
and U6737 (N_6737,N_5228,N_5069);
and U6738 (N_6738,N_5011,N_5704);
xnor U6739 (N_6739,N_5491,N_5218);
nor U6740 (N_6740,N_5925,N_5942);
nor U6741 (N_6741,N_5798,N_5189);
or U6742 (N_6742,N_5012,N_5906);
nand U6743 (N_6743,N_5209,N_5861);
xor U6744 (N_6744,N_5637,N_5435);
nor U6745 (N_6745,N_5567,N_5642);
or U6746 (N_6746,N_5452,N_5925);
xnor U6747 (N_6747,N_5102,N_5141);
or U6748 (N_6748,N_5542,N_5643);
nor U6749 (N_6749,N_5701,N_5081);
xnor U6750 (N_6750,N_5690,N_5360);
and U6751 (N_6751,N_5440,N_5452);
nand U6752 (N_6752,N_5786,N_5128);
and U6753 (N_6753,N_5953,N_5484);
and U6754 (N_6754,N_5818,N_5148);
xor U6755 (N_6755,N_5990,N_5003);
nor U6756 (N_6756,N_5233,N_5351);
nor U6757 (N_6757,N_5851,N_5701);
or U6758 (N_6758,N_5113,N_5092);
nor U6759 (N_6759,N_5760,N_5302);
xor U6760 (N_6760,N_5238,N_5397);
xnor U6761 (N_6761,N_5706,N_5309);
nor U6762 (N_6762,N_5469,N_5604);
xnor U6763 (N_6763,N_5850,N_5954);
xor U6764 (N_6764,N_5744,N_5611);
and U6765 (N_6765,N_5836,N_5270);
and U6766 (N_6766,N_5774,N_5547);
and U6767 (N_6767,N_5035,N_5596);
and U6768 (N_6768,N_5631,N_5693);
nand U6769 (N_6769,N_5629,N_5736);
or U6770 (N_6770,N_5090,N_5778);
nor U6771 (N_6771,N_5238,N_5393);
nor U6772 (N_6772,N_5889,N_5784);
or U6773 (N_6773,N_5635,N_5056);
and U6774 (N_6774,N_5250,N_5246);
nand U6775 (N_6775,N_5885,N_5874);
nand U6776 (N_6776,N_5384,N_5690);
or U6777 (N_6777,N_5966,N_5892);
nor U6778 (N_6778,N_5629,N_5007);
nor U6779 (N_6779,N_5290,N_5221);
nor U6780 (N_6780,N_5347,N_5745);
nor U6781 (N_6781,N_5030,N_5250);
or U6782 (N_6782,N_5616,N_5466);
and U6783 (N_6783,N_5852,N_5515);
nand U6784 (N_6784,N_5218,N_5998);
or U6785 (N_6785,N_5047,N_5074);
or U6786 (N_6786,N_5906,N_5423);
nand U6787 (N_6787,N_5852,N_5844);
and U6788 (N_6788,N_5828,N_5433);
nand U6789 (N_6789,N_5416,N_5486);
nor U6790 (N_6790,N_5779,N_5861);
or U6791 (N_6791,N_5249,N_5166);
and U6792 (N_6792,N_5984,N_5725);
nor U6793 (N_6793,N_5593,N_5264);
or U6794 (N_6794,N_5840,N_5240);
nand U6795 (N_6795,N_5887,N_5996);
nor U6796 (N_6796,N_5646,N_5848);
xor U6797 (N_6797,N_5909,N_5930);
or U6798 (N_6798,N_5603,N_5573);
or U6799 (N_6799,N_5926,N_5454);
nand U6800 (N_6800,N_5644,N_5806);
nor U6801 (N_6801,N_5102,N_5305);
nand U6802 (N_6802,N_5398,N_5239);
or U6803 (N_6803,N_5928,N_5397);
or U6804 (N_6804,N_5239,N_5902);
nor U6805 (N_6805,N_5218,N_5346);
or U6806 (N_6806,N_5165,N_5683);
or U6807 (N_6807,N_5639,N_5152);
xnor U6808 (N_6808,N_5391,N_5199);
and U6809 (N_6809,N_5748,N_5436);
and U6810 (N_6810,N_5557,N_5739);
or U6811 (N_6811,N_5160,N_5172);
and U6812 (N_6812,N_5791,N_5053);
xnor U6813 (N_6813,N_5195,N_5522);
nor U6814 (N_6814,N_5124,N_5927);
or U6815 (N_6815,N_5578,N_5841);
and U6816 (N_6816,N_5201,N_5068);
xor U6817 (N_6817,N_5060,N_5938);
and U6818 (N_6818,N_5281,N_5627);
nor U6819 (N_6819,N_5819,N_5034);
nand U6820 (N_6820,N_5146,N_5604);
and U6821 (N_6821,N_5043,N_5667);
and U6822 (N_6822,N_5068,N_5166);
and U6823 (N_6823,N_5110,N_5905);
nor U6824 (N_6824,N_5767,N_5558);
xnor U6825 (N_6825,N_5313,N_5944);
nand U6826 (N_6826,N_5012,N_5557);
nand U6827 (N_6827,N_5750,N_5946);
nand U6828 (N_6828,N_5322,N_5605);
and U6829 (N_6829,N_5424,N_5161);
xor U6830 (N_6830,N_5361,N_5066);
or U6831 (N_6831,N_5615,N_5168);
and U6832 (N_6832,N_5453,N_5216);
or U6833 (N_6833,N_5760,N_5453);
nand U6834 (N_6834,N_5694,N_5274);
or U6835 (N_6835,N_5680,N_5906);
nor U6836 (N_6836,N_5095,N_5858);
or U6837 (N_6837,N_5139,N_5706);
and U6838 (N_6838,N_5875,N_5131);
xor U6839 (N_6839,N_5826,N_5079);
xnor U6840 (N_6840,N_5147,N_5632);
nand U6841 (N_6841,N_5682,N_5357);
or U6842 (N_6842,N_5316,N_5658);
nor U6843 (N_6843,N_5722,N_5615);
or U6844 (N_6844,N_5099,N_5186);
and U6845 (N_6845,N_5058,N_5899);
nand U6846 (N_6846,N_5444,N_5402);
or U6847 (N_6847,N_5370,N_5734);
nor U6848 (N_6848,N_5040,N_5134);
or U6849 (N_6849,N_5208,N_5897);
or U6850 (N_6850,N_5822,N_5216);
xnor U6851 (N_6851,N_5783,N_5716);
and U6852 (N_6852,N_5872,N_5551);
nor U6853 (N_6853,N_5894,N_5142);
or U6854 (N_6854,N_5279,N_5739);
xor U6855 (N_6855,N_5431,N_5001);
xnor U6856 (N_6856,N_5129,N_5436);
and U6857 (N_6857,N_5022,N_5490);
xor U6858 (N_6858,N_5609,N_5803);
and U6859 (N_6859,N_5422,N_5367);
nand U6860 (N_6860,N_5097,N_5526);
nor U6861 (N_6861,N_5628,N_5783);
or U6862 (N_6862,N_5026,N_5353);
nand U6863 (N_6863,N_5146,N_5720);
or U6864 (N_6864,N_5313,N_5653);
nor U6865 (N_6865,N_5759,N_5600);
nor U6866 (N_6866,N_5147,N_5017);
xnor U6867 (N_6867,N_5888,N_5577);
xor U6868 (N_6868,N_5466,N_5630);
xor U6869 (N_6869,N_5798,N_5815);
xor U6870 (N_6870,N_5300,N_5980);
nor U6871 (N_6871,N_5503,N_5639);
nand U6872 (N_6872,N_5799,N_5136);
nor U6873 (N_6873,N_5131,N_5482);
and U6874 (N_6874,N_5267,N_5117);
nor U6875 (N_6875,N_5646,N_5447);
and U6876 (N_6876,N_5881,N_5446);
nand U6877 (N_6877,N_5616,N_5050);
and U6878 (N_6878,N_5458,N_5333);
and U6879 (N_6879,N_5200,N_5905);
and U6880 (N_6880,N_5629,N_5285);
nand U6881 (N_6881,N_5578,N_5761);
or U6882 (N_6882,N_5042,N_5164);
or U6883 (N_6883,N_5744,N_5615);
nor U6884 (N_6884,N_5286,N_5448);
xor U6885 (N_6885,N_5787,N_5148);
or U6886 (N_6886,N_5714,N_5539);
nand U6887 (N_6887,N_5302,N_5811);
nand U6888 (N_6888,N_5586,N_5345);
and U6889 (N_6889,N_5303,N_5826);
or U6890 (N_6890,N_5206,N_5885);
nor U6891 (N_6891,N_5413,N_5446);
nand U6892 (N_6892,N_5212,N_5566);
xnor U6893 (N_6893,N_5659,N_5186);
or U6894 (N_6894,N_5734,N_5049);
or U6895 (N_6895,N_5649,N_5892);
nor U6896 (N_6896,N_5672,N_5506);
xor U6897 (N_6897,N_5863,N_5918);
or U6898 (N_6898,N_5131,N_5807);
nor U6899 (N_6899,N_5443,N_5783);
nand U6900 (N_6900,N_5990,N_5323);
and U6901 (N_6901,N_5061,N_5295);
xnor U6902 (N_6902,N_5010,N_5801);
or U6903 (N_6903,N_5478,N_5933);
nor U6904 (N_6904,N_5604,N_5592);
nor U6905 (N_6905,N_5820,N_5449);
nand U6906 (N_6906,N_5620,N_5088);
xnor U6907 (N_6907,N_5847,N_5638);
xor U6908 (N_6908,N_5928,N_5334);
and U6909 (N_6909,N_5470,N_5769);
and U6910 (N_6910,N_5968,N_5459);
xor U6911 (N_6911,N_5838,N_5553);
nor U6912 (N_6912,N_5334,N_5092);
and U6913 (N_6913,N_5588,N_5268);
nand U6914 (N_6914,N_5806,N_5681);
nor U6915 (N_6915,N_5169,N_5351);
nor U6916 (N_6916,N_5762,N_5286);
xnor U6917 (N_6917,N_5602,N_5310);
xor U6918 (N_6918,N_5943,N_5314);
nand U6919 (N_6919,N_5025,N_5579);
or U6920 (N_6920,N_5480,N_5829);
and U6921 (N_6921,N_5575,N_5294);
and U6922 (N_6922,N_5934,N_5985);
nand U6923 (N_6923,N_5161,N_5252);
or U6924 (N_6924,N_5551,N_5236);
xnor U6925 (N_6925,N_5239,N_5119);
nand U6926 (N_6926,N_5318,N_5615);
or U6927 (N_6927,N_5932,N_5978);
nor U6928 (N_6928,N_5057,N_5847);
or U6929 (N_6929,N_5329,N_5000);
nand U6930 (N_6930,N_5186,N_5166);
and U6931 (N_6931,N_5032,N_5539);
nand U6932 (N_6932,N_5655,N_5642);
nand U6933 (N_6933,N_5842,N_5695);
xor U6934 (N_6934,N_5468,N_5478);
nor U6935 (N_6935,N_5739,N_5336);
and U6936 (N_6936,N_5154,N_5262);
or U6937 (N_6937,N_5058,N_5374);
and U6938 (N_6938,N_5079,N_5251);
nand U6939 (N_6939,N_5760,N_5378);
nor U6940 (N_6940,N_5632,N_5979);
nor U6941 (N_6941,N_5750,N_5176);
or U6942 (N_6942,N_5137,N_5211);
and U6943 (N_6943,N_5058,N_5558);
nor U6944 (N_6944,N_5650,N_5106);
and U6945 (N_6945,N_5463,N_5206);
or U6946 (N_6946,N_5201,N_5768);
nor U6947 (N_6947,N_5932,N_5391);
xor U6948 (N_6948,N_5587,N_5223);
nor U6949 (N_6949,N_5978,N_5750);
nand U6950 (N_6950,N_5557,N_5685);
xnor U6951 (N_6951,N_5069,N_5631);
or U6952 (N_6952,N_5609,N_5876);
or U6953 (N_6953,N_5339,N_5693);
and U6954 (N_6954,N_5624,N_5771);
or U6955 (N_6955,N_5105,N_5924);
or U6956 (N_6956,N_5670,N_5634);
nand U6957 (N_6957,N_5686,N_5745);
and U6958 (N_6958,N_5802,N_5817);
xor U6959 (N_6959,N_5006,N_5064);
xnor U6960 (N_6960,N_5107,N_5292);
xor U6961 (N_6961,N_5168,N_5862);
and U6962 (N_6962,N_5903,N_5425);
nor U6963 (N_6963,N_5992,N_5911);
nand U6964 (N_6964,N_5053,N_5764);
nor U6965 (N_6965,N_5249,N_5042);
and U6966 (N_6966,N_5429,N_5831);
xor U6967 (N_6967,N_5523,N_5783);
or U6968 (N_6968,N_5148,N_5595);
and U6969 (N_6969,N_5776,N_5509);
xnor U6970 (N_6970,N_5149,N_5081);
or U6971 (N_6971,N_5881,N_5155);
nand U6972 (N_6972,N_5150,N_5742);
xnor U6973 (N_6973,N_5266,N_5905);
or U6974 (N_6974,N_5469,N_5058);
nand U6975 (N_6975,N_5072,N_5912);
nand U6976 (N_6976,N_5382,N_5738);
and U6977 (N_6977,N_5522,N_5049);
and U6978 (N_6978,N_5873,N_5930);
and U6979 (N_6979,N_5200,N_5365);
and U6980 (N_6980,N_5541,N_5577);
nor U6981 (N_6981,N_5589,N_5561);
xnor U6982 (N_6982,N_5355,N_5917);
and U6983 (N_6983,N_5495,N_5098);
and U6984 (N_6984,N_5752,N_5948);
xor U6985 (N_6985,N_5597,N_5902);
nor U6986 (N_6986,N_5470,N_5340);
nand U6987 (N_6987,N_5124,N_5101);
and U6988 (N_6988,N_5928,N_5947);
xor U6989 (N_6989,N_5552,N_5710);
and U6990 (N_6990,N_5628,N_5838);
xor U6991 (N_6991,N_5739,N_5510);
nand U6992 (N_6992,N_5087,N_5388);
nand U6993 (N_6993,N_5813,N_5256);
xor U6994 (N_6994,N_5290,N_5618);
nor U6995 (N_6995,N_5396,N_5282);
nor U6996 (N_6996,N_5198,N_5463);
xnor U6997 (N_6997,N_5603,N_5910);
or U6998 (N_6998,N_5346,N_5092);
nor U6999 (N_6999,N_5296,N_5503);
or U7000 (N_7000,N_6335,N_6188);
xor U7001 (N_7001,N_6765,N_6763);
xor U7002 (N_7002,N_6899,N_6028);
nor U7003 (N_7003,N_6803,N_6439);
xor U7004 (N_7004,N_6777,N_6648);
or U7005 (N_7005,N_6527,N_6396);
and U7006 (N_7006,N_6161,N_6878);
xnor U7007 (N_7007,N_6271,N_6566);
or U7008 (N_7008,N_6965,N_6636);
nand U7009 (N_7009,N_6924,N_6992);
nor U7010 (N_7010,N_6302,N_6366);
nor U7011 (N_7011,N_6189,N_6886);
nor U7012 (N_7012,N_6283,N_6670);
or U7013 (N_7013,N_6157,N_6855);
and U7014 (N_7014,N_6957,N_6860);
xnor U7015 (N_7015,N_6608,N_6953);
or U7016 (N_7016,N_6251,N_6498);
xor U7017 (N_7017,N_6696,N_6693);
xnor U7018 (N_7018,N_6208,N_6340);
and U7019 (N_7019,N_6902,N_6871);
or U7020 (N_7020,N_6404,N_6213);
nor U7021 (N_7021,N_6543,N_6460);
or U7022 (N_7022,N_6916,N_6958);
nor U7023 (N_7023,N_6782,N_6625);
nand U7024 (N_7024,N_6417,N_6114);
or U7025 (N_7025,N_6504,N_6268);
nor U7026 (N_7026,N_6424,N_6526);
xor U7027 (N_7027,N_6416,N_6699);
or U7028 (N_7028,N_6657,N_6661);
nand U7029 (N_7029,N_6132,N_6808);
xnor U7030 (N_7030,N_6863,N_6063);
nand U7031 (N_7031,N_6178,N_6914);
and U7032 (N_7032,N_6621,N_6182);
xor U7033 (N_7033,N_6509,N_6180);
and U7034 (N_7034,N_6336,N_6284);
nor U7035 (N_7035,N_6787,N_6331);
nor U7036 (N_7036,N_6123,N_6736);
nand U7037 (N_7037,N_6394,N_6111);
nor U7038 (N_7038,N_6956,N_6370);
or U7039 (N_7039,N_6497,N_6294);
xor U7040 (N_7040,N_6053,N_6843);
xnor U7041 (N_7041,N_6649,N_6673);
and U7042 (N_7042,N_6514,N_6406);
nor U7043 (N_7043,N_6805,N_6982);
nand U7044 (N_7044,N_6952,N_6116);
and U7045 (N_7045,N_6589,N_6119);
and U7046 (N_7046,N_6606,N_6741);
or U7047 (N_7047,N_6609,N_6092);
xnor U7048 (N_7048,N_6304,N_6254);
nand U7049 (N_7049,N_6219,N_6493);
nor U7050 (N_7050,N_6379,N_6517);
xnor U7051 (N_7051,N_6584,N_6017);
nor U7052 (N_7052,N_6462,N_6272);
or U7053 (N_7053,N_6140,N_6541);
or U7054 (N_7054,N_6716,N_6840);
nand U7055 (N_7055,N_6906,N_6922);
nor U7056 (N_7056,N_6680,N_6296);
and U7057 (N_7057,N_6666,N_6635);
xor U7058 (N_7058,N_6739,N_6731);
nand U7059 (N_7059,N_6263,N_6454);
and U7060 (N_7060,N_6230,N_6050);
nor U7061 (N_7061,N_6072,N_6455);
or U7062 (N_7062,N_6653,N_6133);
xnor U7063 (N_7063,N_6773,N_6276);
or U7064 (N_7064,N_6764,N_6233);
or U7065 (N_7065,N_6298,N_6849);
or U7066 (N_7066,N_6890,N_6784);
nand U7067 (N_7067,N_6904,N_6908);
and U7068 (N_7068,N_6684,N_6138);
nand U7069 (N_7069,N_6110,N_6875);
nor U7070 (N_7070,N_6386,N_6991);
nand U7071 (N_7071,N_6576,N_6872);
xor U7072 (N_7072,N_6437,N_6196);
xor U7073 (N_7073,N_6442,N_6175);
nand U7074 (N_7074,N_6363,N_6715);
nand U7075 (N_7075,N_6828,N_6647);
nor U7076 (N_7076,N_6832,N_6382);
nor U7077 (N_7077,N_6099,N_6478);
and U7078 (N_7078,N_6996,N_6000);
or U7079 (N_7079,N_6241,N_6246);
xnor U7080 (N_7080,N_6620,N_6681);
nand U7081 (N_7081,N_6227,N_6311);
and U7082 (N_7082,N_6411,N_6546);
nor U7083 (N_7083,N_6788,N_6614);
nand U7084 (N_7084,N_6937,N_6744);
or U7085 (N_7085,N_6658,N_6995);
nand U7086 (N_7086,N_6717,N_6101);
or U7087 (N_7087,N_6853,N_6148);
xnor U7088 (N_7088,N_6426,N_6469);
or U7089 (N_7089,N_6791,N_6652);
nand U7090 (N_7090,N_6868,N_6605);
or U7091 (N_7091,N_6950,N_6122);
nor U7092 (N_7092,N_6361,N_6238);
nor U7093 (N_7093,N_6139,N_6578);
nor U7094 (N_7094,N_6405,N_6934);
xor U7095 (N_7095,N_6740,N_6326);
nand U7096 (N_7096,N_6938,N_6389);
or U7097 (N_7097,N_6894,N_6195);
xnor U7098 (N_7098,N_6983,N_6295);
and U7099 (N_7099,N_6553,N_6354);
or U7100 (N_7100,N_6051,N_6003);
nand U7101 (N_7101,N_6796,N_6240);
or U7102 (N_7102,N_6203,N_6702);
xnor U7103 (N_7103,N_6436,N_6206);
nand U7104 (N_7104,N_6435,N_6976);
nor U7105 (N_7105,N_6274,N_6323);
xor U7106 (N_7106,N_6960,N_6260);
nand U7107 (N_7107,N_6282,N_6714);
or U7108 (N_7108,N_6951,N_6646);
nor U7109 (N_7109,N_6984,N_6826);
nand U7110 (N_7110,N_6107,N_6806);
and U7111 (N_7111,N_6809,N_6540);
nor U7112 (N_7112,N_6719,N_6743);
or U7113 (N_7113,N_6535,N_6380);
nand U7114 (N_7114,N_6852,N_6367);
nand U7115 (N_7115,N_6727,N_6624);
and U7116 (N_7116,N_6306,N_6496);
and U7117 (N_7117,N_6501,N_6262);
and U7118 (N_7118,N_6359,N_6758);
or U7119 (N_7119,N_6876,N_6309);
or U7120 (N_7120,N_6040,N_6930);
xor U7121 (N_7121,N_6597,N_6163);
or U7122 (N_7122,N_6135,N_6619);
and U7123 (N_7123,N_6468,N_6602);
or U7124 (N_7124,N_6165,N_6559);
xnor U7125 (N_7125,N_6117,N_6001);
nand U7126 (N_7126,N_6058,N_6007);
xor U7127 (N_7127,N_6793,N_6754);
nor U7128 (N_7128,N_6009,N_6185);
or U7129 (N_7129,N_6324,N_6850);
xnor U7130 (N_7130,N_6722,N_6836);
nand U7131 (N_7131,N_6459,N_6156);
nor U7132 (N_7132,N_6569,N_6512);
nand U7133 (N_7133,N_6476,N_6697);
nor U7134 (N_7134,N_6325,N_6289);
and U7135 (N_7135,N_6672,N_6954);
nor U7136 (N_7136,N_6688,N_6328);
or U7137 (N_7137,N_6037,N_6008);
and U7138 (N_7138,N_6663,N_6356);
or U7139 (N_7139,N_6834,N_6373);
xor U7140 (N_7140,N_6089,N_6239);
nor U7141 (N_7141,N_6923,N_6994);
nor U7142 (N_7142,N_6898,N_6748);
or U7143 (N_7143,N_6821,N_6634);
xnor U7144 (N_7144,N_6495,N_6989);
or U7145 (N_7145,N_6068,N_6160);
nand U7146 (N_7146,N_6980,N_6330);
and U7147 (N_7147,N_6143,N_6313);
and U7148 (N_7148,N_6613,N_6461);
nor U7149 (N_7149,N_6884,N_6529);
nor U7150 (N_7150,N_6745,N_6757);
nor U7151 (N_7151,N_6870,N_6244);
and U7152 (N_7152,N_6145,N_6835);
nand U7153 (N_7153,N_6299,N_6491);
and U7154 (N_7154,N_6901,N_6480);
and U7155 (N_7155,N_6665,N_6257);
xor U7156 (N_7156,N_6993,N_6974);
xor U7157 (N_7157,N_6785,N_6959);
or U7158 (N_7158,N_6686,N_6617);
and U7159 (N_7159,N_6287,N_6291);
nand U7160 (N_7160,N_6747,N_6293);
xnor U7161 (N_7161,N_6059,N_6275);
nor U7162 (N_7162,N_6909,N_6467);
or U7163 (N_7163,N_6709,N_6544);
and U7164 (N_7164,N_6795,N_6664);
and U7165 (N_7165,N_6388,N_6968);
or U7166 (N_7166,N_6481,N_6432);
xor U7167 (N_7167,N_6494,N_6513);
and U7168 (N_7168,N_6199,N_6761);
and U7169 (N_7169,N_6510,N_6940);
and U7170 (N_7170,N_6842,N_6637);
nand U7171 (N_7171,N_6060,N_6557);
or U7172 (N_7172,N_6485,N_6593);
nand U7173 (N_7173,N_6942,N_6016);
and U7174 (N_7174,N_6452,N_6713);
nand U7175 (N_7175,N_6204,N_6162);
xor U7176 (N_7176,N_6499,N_6742);
nand U7177 (N_7177,N_6470,N_6750);
nand U7178 (N_7178,N_6242,N_6874);
and U7179 (N_7179,N_6466,N_6997);
and U7180 (N_7180,N_6112,N_6025);
nand U7181 (N_7181,N_6895,N_6611);
nor U7182 (N_7182,N_6746,N_6098);
or U7183 (N_7183,N_6216,N_6171);
nor U7184 (N_7184,N_6538,N_6897);
and U7185 (N_7185,N_6560,N_6641);
xnor U7186 (N_7186,N_6026,N_6749);
nand U7187 (N_7187,N_6177,N_6319);
xnor U7188 (N_7188,N_6679,N_6408);
nand U7189 (N_7189,N_6457,N_6712);
xor U7190 (N_7190,N_6586,N_6622);
or U7191 (N_7191,N_6228,N_6151);
nor U7192 (N_7192,N_6015,N_6700);
nor U7193 (N_7193,N_6285,N_6243);
nand U7194 (N_7194,N_6660,N_6103);
xnor U7195 (N_7195,N_6728,N_6531);
or U7196 (N_7196,N_6292,N_6255);
xnor U7197 (N_7197,N_6817,N_6558);
nand U7198 (N_7198,N_6091,N_6447);
xnor U7199 (N_7199,N_6610,N_6489);
or U7200 (N_7200,N_6214,N_6031);
or U7201 (N_7201,N_6288,N_6598);
nor U7202 (N_7202,N_6236,N_6550);
nor U7203 (N_7203,N_6572,N_6223);
or U7204 (N_7204,N_6054,N_6887);
nand U7205 (N_7205,N_6174,N_6004);
nor U7206 (N_7206,N_6453,N_6445);
nand U7207 (N_7207,N_6618,N_6039);
nor U7208 (N_7208,N_6858,N_6390);
xor U7209 (N_7209,N_6418,N_6153);
and U7210 (N_7210,N_6802,N_6705);
nor U7211 (N_7211,N_6385,N_6534);
nand U7212 (N_7212,N_6594,N_6192);
or U7213 (N_7213,N_6250,N_6628);
xnor U7214 (N_7214,N_6674,N_6905);
nor U7215 (N_7215,N_6656,N_6603);
nand U7216 (N_7216,N_6524,N_6183);
or U7217 (N_7217,N_6536,N_6378);
and U7218 (N_7218,N_6915,N_6813);
nand U7219 (N_7219,N_6322,N_6772);
and U7220 (N_7220,N_6252,N_6108);
nand U7221 (N_7221,N_6095,N_6044);
xnor U7222 (N_7222,N_6479,N_6794);
xor U7223 (N_7223,N_6824,N_6917);
or U7224 (N_7224,N_6662,N_6176);
xor U7225 (N_7225,N_6869,N_6212);
or U7226 (N_7226,N_6281,N_6321);
xnor U7227 (N_7227,N_6781,N_6574);
xor U7228 (N_7228,N_6303,N_6318);
xor U7229 (N_7229,N_6925,N_6018);
nand U7230 (N_7230,N_6730,N_6790);
nor U7231 (N_7231,N_6383,N_6846);
xor U7232 (N_7232,N_6259,N_6172);
nand U7233 (N_7233,N_6990,N_6070);
nor U7234 (N_7234,N_6082,N_6429);
nand U7235 (N_7235,N_6775,N_6170);
nand U7236 (N_7236,N_6399,N_6011);
xor U7237 (N_7237,N_6542,N_6677);
or U7238 (N_7238,N_6987,N_6643);
or U7239 (N_7239,N_6630,N_6768);
nor U7240 (N_7240,N_6364,N_6570);
nand U7241 (N_7241,N_6207,N_6533);
or U7242 (N_7242,N_6197,N_6723);
nor U7243 (N_7243,N_6823,N_6409);
nand U7244 (N_7244,N_6353,N_6220);
nor U7245 (N_7245,N_6694,N_6305);
nand U7246 (N_7246,N_6555,N_6537);
nand U7247 (N_7247,N_6804,N_6839);
and U7248 (N_7248,N_6725,N_6487);
xor U7249 (N_7249,N_6086,N_6087);
or U7250 (N_7250,N_6695,N_6807);
or U7251 (N_7251,N_6316,N_6315);
nand U7252 (N_7252,N_6631,N_6726);
or U7253 (N_7253,N_6339,N_6030);
xor U7254 (N_7254,N_6301,N_6933);
xor U7255 (N_7255,N_6946,N_6438);
nand U7256 (N_7256,N_6341,N_6261);
or U7257 (N_7257,N_6596,N_6488);
and U7258 (N_7258,N_6645,N_6430);
xnor U7259 (N_7259,N_6027,N_6190);
xor U7260 (N_7260,N_6819,N_6484);
nand U7261 (N_7261,N_6019,N_6845);
or U7262 (N_7262,N_6751,N_6343);
nand U7263 (N_7263,N_6146,N_6774);
and U7264 (N_7264,N_6351,N_6651);
xnor U7265 (N_7265,N_6888,N_6191);
or U7266 (N_7266,N_6346,N_6671);
nor U7267 (N_7267,N_6626,N_6423);
or U7268 (N_7268,N_6522,N_6482);
or U7269 (N_7269,N_6347,N_6978);
nand U7270 (N_7270,N_6607,N_6848);
and U7271 (N_7271,N_6421,N_6032);
nand U7272 (N_7272,N_6381,N_6711);
or U7273 (N_7273,N_6473,N_6080);
nand U7274 (N_7274,N_6800,N_6943);
or U7275 (N_7275,N_6226,N_6913);
nor U7276 (N_7276,N_6412,N_6097);
and U7277 (N_7277,N_6720,N_6124);
xnor U7278 (N_7278,N_6981,N_6279);
or U7279 (N_7279,N_6278,N_6256);
or U7280 (N_7280,N_6397,N_6320);
and U7281 (N_7281,N_6444,N_6615);
nand U7282 (N_7282,N_6939,N_6910);
or U7283 (N_7283,N_6629,N_6414);
nand U7284 (N_7284,N_6141,N_6471);
and U7285 (N_7285,N_6024,N_6766);
or U7286 (N_7286,N_6838,N_6822);
nor U7287 (N_7287,N_6737,N_6779);
nor U7288 (N_7288,N_6049,N_6595);
nor U7289 (N_7289,N_6857,N_6732);
nor U7290 (N_7290,N_6955,N_6277);
nor U7291 (N_7291,N_6721,N_6164);
xor U7292 (N_7292,N_6879,N_6120);
xnor U7293 (N_7293,N_6300,N_6961);
and U7294 (N_7294,N_6734,N_6883);
nand U7295 (N_7295,N_6882,N_6094);
and U7296 (N_7296,N_6682,N_6801);
nor U7297 (N_7297,N_6985,N_6451);
and U7298 (N_7298,N_6523,N_6685);
and U7299 (N_7299,N_6374,N_6358);
xnor U7300 (N_7300,N_6312,N_6573);
xnor U7301 (N_7301,N_6014,N_6820);
nor U7302 (N_7302,N_6193,N_6733);
nand U7303 (N_7303,N_6632,N_6556);
xor U7304 (N_7304,N_6102,N_6975);
nand U7305 (N_7305,N_6210,N_6759);
or U7306 (N_7306,N_6113,N_6355);
and U7307 (N_7307,N_6181,N_6456);
nand U7308 (N_7308,N_6200,N_6237);
nor U7309 (N_7309,N_6783,N_6859);
nand U7310 (N_7310,N_6064,N_6528);
or U7311 (N_7311,N_6873,N_6267);
nor U7312 (N_7312,N_6041,N_6892);
nor U7313 (N_7313,N_6448,N_6912);
and U7314 (N_7314,N_6604,N_6074);
and U7315 (N_7315,N_6592,N_6856);
nand U7316 (N_7316,N_6971,N_6128);
nand U7317 (N_7317,N_6770,N_6738);
nor U7318 (N_7318,N_6577,N_6034);
and U7319 (N_7319,N_6472,N_6575);
xnor U7320 (N_7320,N_6413,N_6167);
or U7321 (N_7321,N_6490,N_6169);
or U7322 (N_7322,N_6159,N_6446);
nand U7323 (N_7323,N_6581,N_6568);
xnor U7324 (N_7324,N_6235,N_6704);
nand U7325 (N_7325,N_6701,N_6047);
xnor U7326 (N_7326,N_6391,N_6465);
nor U7327 (N_7327,N_6753,N_6225);
xnor U7328 (N_7328,N_6265,N_6075);
and U7329 (N_7329,N_6639,N_6023);
nand U7330 (N_7330,N_6941,N_6329);
nor U7331 (N_7331,N_6392,N_6580);
nor U7332 (N_7332,N_6066,N_6010);
nand U7333 (N_7333,N_6231,N_6689);
and U7334 (N_7334,N_6187,N_6972);
nor U7335 (N_7335,N_6136,N_6038);
nand U7336 (N_7336,N_6198,N_6929);
nor U7337 (N_7337,N_6642,N_6350);
or U7338 (N_7338,N_6571,N_6247);
and U7339 (N_7339,N_6362,N_6797);
and U7340 (N_7340,N_6090,N_6623);
nand U7341 (N_7341,N_6376,N_6920);
and U7342 (N_7342,N_6458,N_6073);
or U7343 (N_7343,N_6118,N_6927);
xnor U7344 (N_7344,N_6121,N_6654);
nor U7345 (N_7345,N_6724,N_6932);
and U7346 (N_7346,N_6209,N_6503);
and U7347 (N_7347,N_6627,N_6729);
and U7348 (N_7348,N_6154,N_6563);
and U7349 (N_7349,N_6515,N_6708);
nor U7350 (N_7350,N_6109,N_6062);
nor U7351 (N_7351,N_6264,N_6889);
and U7352 (N_7352,N_6348,N_6310);
nand U7353 (N_7353,N_6562,N_6425);
nor U7354 (N_7354,N_6085,N_6477);
and U7355 (N_7355,N_6368,N_6464);
xnor U7356 (N_7356,N_6683,N_6078);
nor U7357 (N_7357,N_6218,N_6600);
nand U7358 (N_7358,N_6035,N_6530);
nor U7359 (N_7359,N_6431,N_6520);
nor U7360 (N_7360,N_6449,N_6434);
or U7361 (N_7361,N_6964,N_6061);
nor U7362 (N_7362,N_6640,N_6337);
or U7363 (N_7363,N_6475,N_6829);
or U7364 (N_7364,N_6907,N_6767);
nor U7365 (N_7365,N_6644,N_6201);
nor U7366 (N_7366,N_6345,N_6786);
xnor U7367 (N_7367,N_6043,N_6422);
or U7368 (N_7368,N_6048,N_6847);
nor U7369 (N_7369,N_6825,N_6150);
and U7370 (N_7370,N_6830,N_6771);
nor U7371 (N_7371,N_6710,N_6332);
nor U7372 (N_7372,N_6827,N_6104);
nor U7373 (N_7373,N_6258,N_6342);
xor U7374 (N_7374,N_6194,N_6893);
xnor U7375 (N_7375,N_6552,N_6137);
and U7376 (N_7376,N_6988,N_6401);
or U7377 (N_7377,N_6548,N_6881);
nand U7378 (N_7378,N_6678,N_6234);
or U7379 (N_7379,N_6862,N_6308);
nor U7380 (N_7380,N_6492,N_6221);
and U7381 (N_7381,N_6900,N_6168);
and U7382 (N_7382,N_6273,N_6129);
xor U7383 (N_7383,N_6149,N_6327);
xor U7384 (N_7384,N_6756,N_6880);
and U7385 (N_7385,N_6516,N_6142);
and U7386 (N_7386,N_6998,N_6735);
nand U7387 (N_7387,N_6186,N_6921);
nand U7388 (N_7388,N_6083,N_6387);
xor U7389 (N_7389,N_6071,N_6591);
and U7390 (N_7390,N_6105,N_6115);
and U7391 (N_7391,N_6703,N_6076);
xnor U7392 (N_7392,N_6410,N_6266);
and U7393 (N_7393,N_6052,N_6590);
xor U7394 (N_7394,N_6205,N_6081);
and U7395 (N_7395,N_6601,N_6999);
nor U7396 (N_7396,N_6587,N_6511);
and U7397 (N_7397,N_6963,N_6069);
nand U7398 (N_7398,N_6065,N_6903);
xor U7399 (N_7399,N_6349,N_6760);
or U7400 (N_7400,N_6067,N_6055);
nor U7401 (N_7401,N_6926,N_6928);
xnor U7402 (N_7402,N_6463,N_6502);
nor U7403 (N_7403,N_6357,N_6215);
and U7404 (N_7404,N_6861,N_6211);
xor U7405 (N_7405,N_6935,N_6002);
nor U7406 (N_7406,N_6224,N_6131);
nor U7407 (N_7407,N_6815,N_6518);
and U7408 (N_7408,N_6249,N_6833);
nor U7409 (N_7409,N_6811,N_6633);
xnor U7410 (N_7410,N_6769,N_6778);
nand U7411 (N_7411,N_6564,N_6179);
or U7412 (N_7412,N_6949,N_6655);
xnor U7413 (N_7413,N_6021,N_6706);
and U7414 (N_7414,N_6551,N_6042);
or U7415 (N_7415,N_6029,N_6565);
nor U7416 (N_7416,N_6166,N_6232);
nand U7417 (N_7417,N_6420,N_6789);
nand U7418 (N_7418,N_6100,N_6384);
and U7419 (N_7419,N_6338,N_6134);
nor U7420 (N_7420,N_6317,N_6588);
or U7421 (N_7421,N_6918,N_6173);
and U7422 (N_7422,N_6440,N_6896);
nand U7423 (N_7423,N_6507,N_6307);
xnor U7424 (N_7424,N_6885,N_6864);
and U7425 (N_7425,N_6752,N_6486);
or U7426 (N_7426,N_6152,N_6433);
xor U7427 (N_7427,N_6415,N_6579);
nor U7428 (N_7428,N_6377,N_6547);
nand U7429 (N_7429,N_6269,N_6127);
nand U7430 (N_7430,N_6508,N_6290);
and U7431 (N_7431,N_6612,N_6334);
xor U7432 (N_7432,N_6297,N_6532);
or U7433 (N_7433,N_6931,N_6812);
and U7434 (N_7434,N_6369,N_6599);
and U7435 (N_7435,N_6854,N_6690);
nor U7436 (N_7436,N_6184,N_6911);
xor U7437 (N_7437,N_6393,N_6762);
xnor U7438 (N_7438,N_6799,N_6539);
or U7439 (N_7439,N_6096,N_6837);
nand U7440 (N_7440,N_6500,N_6554);
and U7441 (N_7441,N_6687,N_6036);
and U7442 (N_7442,N_6969,N_6755);
or U7443 (N_7443,N_6202,N_6020);
or U7444 (N_7444,N_6945,N_6561);
and U7445 (N_7445,N_6400,N_6314);
nand U7446 (N_7446,N_6372,N_6816);
xnor U7447 (N_7447,N_6698,N_6398);
nand U7448 (N_7448,N_6005,N_6077);
and U7449 (N_7449,N_6814,N_6253);
nor U7450 (N_7450,N_6944,N_6013);
and U7451 (N_7451,N_6549,N_6147);
nand U7452 (N_7452,N_6093,N_6427);
and U7453 (N_7453,N_6371,N_6865);
and U7454 (N_7454,N_6375,N_6659);
nor U7455 (N_7455,N_6582,N_6443);
or U7456 (N_7456,N_6245,N_6891);
and U7457 (N_7457,N_6585,N_6667);
nor U7458 (N_7458,N_6365,N_6810);
nand U7459 (N_7459,N_6780,N_6676);
nand U7460 (N_7460,N_6718,N_6428);
or U7461 (N_7461,N_6056,N_6545);
and U7462 (N_7462,N_6217,N_6776);
nand U7463 (N_7463,N_6525,N_6877);
and U7464 (N_7464,N_6919,N_6521);
xnor U7465 (N_7465,N_6947,N_6125);
or U7466 (N_7466,N_6851,N_6792);
or U7467 (N_7467,N_6403,N_6650);
or U7468 (N_7468,N_6844,N_6866);
and U7469 (N_7469,N_6668,N_6691);
and U7470 (N_7470,N_6841,N_6979);
nand U7471 (N_7471,N_6033,N_6519);
nor U7472 (N_7472,N_6130,N_6126);
or U7473 (N_7473,N_6948,N_6222);
or U7474 (N_7474,N_6158,N_6280);
nand U7475 (N_7475,N_6986,N_6395);
and U7476 (N_7476,N_6106,N_6079);
or U7477 (N_7477,N_6286,N_6144);
and U7478 (N_7478,N_6818,N_6669);
xnor U7479 (N_7479,N_6419,N_6506);
and U7480 (N_7480,N_6474,N_6407);
nor U7481 (N_7481,N_6088,N_6616);
nor U7482 (N_7482,N_6966,N_6967);
xnor U7483 (N_7483,N_6973,N_6270);
nor U7484 (N_7484,N_6692,N_6022);
and U7485 (N_7485,N_6483,N_6936);
or U7486 (N_7486,N_6970,N_6977);
or U7487 (N_7487,N_6012,N_6229);
and U7488 (N_7488,N_6352,N_6707);
nand U7489 (N_7489,N_6344,N_6248);
nand U7490 (N_7490,N_6831,N_6450);
xnor U7491 (N_7491,N_6057,N_6638);
or U7492 (N_7492,N_6867,N_6402);
and U7493 (N_7493,N_6505,N_6045);
xnor U7494 (N_7494,N_6798,N_6084);
xor U7495 (N_7495,N_6583,N_6155);
nor U7496 (N_7496,N_6962,N_6333);
xnor U7497 (N_7497,N_6675,N_6360);
or U7498 (N_7498,N_6006,N_6567);
and U7499 (N_7499,N_6046,N_6441);
nor U7500 (N_7500,N_6094,N_6138);
xnor U7501 (N_7501,N_6070,N_6027);
nand U7502 (N_7502,N_6461,N_6135);
or U7503 (N_7503,N_6670,N_6294);
or U7504 (N_7504,N_6537,N_6467);
or U7505 (N_7505,N_6167,N_6668);
and U7506 (N_7506,N_6015,N_6399);
nor U7507 (N_7507,N_6797,N_6437);
nor U7508 (N_7508,N_6846,N_6212);
xor U7509 (N_7509,N_6633,N_6238);
and U7510 (N_7510,N_6025,N_6564);
xnor U7511 (N_7511,N_6979,N_6723);
xnor U7512 (N_7512,N_6685,N_6090);
and U7513 (N_7513,N_6786,N_6748);
or U7514 (N_7514,N_6320,N_6473);
xor U7515 (N_7515,N_6172,N_6098);
or U7516 (N_7516,N_6175,N_6786);
or U7517 (N_7517,N_6836,N_6560);
or U7518 (N_7518,N_6713,N_6176);
nor U7519 (N_7519,N_6599,N_6932);
xnor U7520 (N_7520,N_6649,N_6498);
or U7521 (N_7521,N_6087,N_6523);
or U7522 (N_7522,N_6785,N_6383);
xnor U7523 (N_7523,N_6378,N_6816);
nor U7524 (N_7524,N_6596,N_6105);
nor U7525 (N_7525,N_6341,N_6237);
or U7526 (N_7526,N_6781,N_6903);
and U7527 (N_7527,N_6985,N_6869);
or U7528 (N_7528,N_6985,N_6614);
xnor U7529 (N_7529,N_6816,N_6546);
nor U7530 (N_7530,N_6418,N_6119);
nor U7531 (N_7531,N_6292,N_6703);
xnor U7532 (N_7532,N_6398,N_6259);
xnor U7533 (N_7533,N_6079,N_6927);
nand U7534 (N_7534,N_6680,N_6349);
nor U7535 (N_7535,N_6554,N_6302);
xnor U7536 (N_7536,N_6086,N_6197);
nor U7537 (N_7537,N_6331,N_6247);
nor U7538 (N_7538,N_6269,N_6342);
nand U7539 (N_7539,N_6949,N_6960);
and U7540 (N_7540,N_6650,N_6644);
nor U7541 (N_7541,N_6319,N_6087);
or U7542 (N_7542,N_6212,N_6399);
nor U7543 (N_7543,N_6954,N_6354);
xor U7544 (N_7544,N_6481,N_6442);
xor U7545 (N_7545,N_6796,N_6039);
nand U7546 (N_7546,N_6513,N_6274);
and U7547 (N_7547,N_6961,N_6905);
nor U7548 (N_7548,N_6753,N_6376);
and U7549 (N_7549,N_6553,N_6695);
xnor U7550 (N_7550,N_6624,N_6233);
nand U7551 (N_7551,N_6892,N_6406);
or U7552 (N_7552,N_6942,N_6149);
nand U7553 (N_7553,N_6104,N_6953);
nor U7554 (N_7554,N_6902,N_6346);
xnor U7555 (N_7555,N_6008,N_6518);
nor U7556 (N_7556,N_6723,N_6676);
nand U7557 (N_7557,N_6739,N_6307);
nor U7558 (N_7558,N_6326,N_6440);
nor U7559 (N_7559,N_6835,N_6035);
nor U7560 (N_7560,N_6437,N_6220);
and U7561 (N_7561,N_6072,N_6168);
and U7562 (N_7562,N_6759,N_6001);
xor U7563 (N_7563,N_6537,N_6898);
xnor U7564 (N_7564,N_6636,N_6358);
nand U7565 (N_7565,N_6539,N_6184);
or U7566 (N_7566,N_6488,N_6207);
or U7567 (N_7567,N_6922,N_6455);
xor U7568 (N_7568,N_6198,N_6806);
nor U7569 (N_7569,N_6898,N_6356);
nand U7570 (N_7570,N_6995,N_6547);
or U7571 (N_7571,N_6001,N_6748);
nor U7572 (N_7572,N_6117,N_6884);
and U7573 (N_7573,N_6759,N_6280);
nor U7574 (N_7574,N_6424,N_6692);
xnor U7575 (N_7575,N_6892,N_6427);
or U7576 (N_7576,N_6590,N_6575);
nand U7577 (N_7577,N_6431,N_6754);
xor U7578 (N_7578,N_6184,N_6989);
and U7579 (N_7579,N_6491,N_6242);
nand U7580 (N_7580,N_6560,N_6482);
nand U7581 (N_7581,N_6728,N_6628);
or U7582 (N_7582,N_6946,N_6872);
nor U7583 (N_7583,N_6593,N_6060);
and U7584 (N_7584,N_6602,N_6259);
nor U7585 (N_7585,N_6261,N_6138);
nor U7586 (N_7586,N_6382,N_6214);
and U7587 (N_7587,N_6629,N_6707);
and U7588 (N_7588,N_6111,N_6419);
and U7589 (N_7589,N_6364,N_6591);
nor U7590 (N_7590,N_6503,N_6004);
xor U7591 (N_7591,N_6776,N_6623);
nand U7592 (N_7592,N_6712,N_6202);
xor U7593 (N_7593,N_6912,N_6271);
nand U7594 (N_7594,N_6031,N_6490);
or U7595 (N_7595,N_6555,N_6437);
xnor U7596 (N_7596,N_6723,N_6841);
nor U7597 (N_7597,N_6845,N_6740);
nand U7598 (N_7598,N_6252,N_6096);
or U7599 (N_7599,N_6855,N_6411);
or U7600 (N_7600,N_6276,N_6469);
xor U7601 (N_7601,N_6670,N_6181);
and U7602 (N_7602,N_6422,N_6619);
nor U7603 (N_7603,N_6975,N_6751);
xor U7604 (N_7604,N_6541,N_6785);
nand U7605 (N_7605,N_6532,N_6907);
nand U7606 (N_7606,N_6324,N_6826);
and U7607 (N_7607,N_6115,N_6932);
and U7608 (N_7608,N_6287,N_6481);
or U7609 (N_7609,N_6080,N_6077);
xnor U7610 (N_7610,N_6512,N_6510);
nand U7611 (N_7611,N_6558,N_6027);
nand U7612 (N_7612,N_6050,N_6191);
nand U7613 (N_7613,N_6107,N_6966);
nand U7614 (N_7614,N_6913,N_6171);
and U7615 (N_7615,N_6761,N_6422);
xnor U7616 (N_7616,N_6416,N_6246);
xnor U7617 (N_7617,N_6018,N_6516);
xor U7618 (N_7618,N_6821,N_6917);
and U7619 (N_7619,N_6293,N_6122);
nor U7620 (N_7620,N_6930,N_6416);
and U7621 (N_7621,N_6176,N_6380);
xor U7622 (N_7622,N_6743,N_6892);
and U7623 (N_7623,N_6909,N_6266);
xnor U7624 (N_7624,N_6102,N_6990);
and U7625 (N_7625,N_6369,N_6210);
or U7626 (N_7626,N_6922,N_6388);
nand U7627 (N_7627,N_6696,N_6559);
or U7628 (N_7628,N_6376,N_6349);
or U7629 (N_7629,N_6839,N_6961);
or U7630 (N_7630,N_6422,N_6190);
nor U7631 (N_7631,N_6073,N_6837);
and U7632 (N_7632,N_6621,N_6848);
and U7633 (N_7633,N_6420,N_6676);
or U7634 (N_7634,N_6624,N_6215);
or U7635 (N_7635,N_6776,N_6226);
nand U7636 (N_7636,N_6928,N_6265);
xnor U7637 (N_7637,N_6287,N_6303);
or U7638 (N_7638,N_6299,N_6807);
nand U7639 (N_7639,N_6993,N_6558);
and U7640 (N_7640,N_6128,N_6236);
and U7641 (N_7641,N_6894,N_6899);
nand U7642 (N_7642,N_6768,N_6364);
nor U7643 (N_7643,N_6266,N_6478);
nor U7644 (N_7644,N_6674,N_6549);
nor U7645 (N_7645,N_6784,N_6258);
or U7646 (N_7646,N_6796,N_6594);
xnor U7647 (N_7647,N_6450,N_6879);
nand U7648 (N_7648,N_6143,N_6604);
xor U7649 (N_7649,N_6093,N_6334);
nand U7650 (N_7650,N_6498,N_6773);
nand U7651 (N_7651,N_6949,N_6304);
nand U7652 (N_7652,N_6314,N_6137);
and U7653 (N_7653,N_6089,N_6577);
nor U7654 (N_7654,N_6803,N_6881);
or U7655 (N_7655,N_6586,N_6757);
xor U7656 (N_7656,N_6806,N_6931);
nor U7657 (N_7657,N_6555,N_6702);
nand U7658 (N_7658,N_6603,N_6273);
and U7659 (N_7659,N_6850,N_6277);
nor U7660 (N_7660,N_6316,N_6042);
and U7661 (N_7661,N_6146,N_6439);
xnor U7662 (N_7662,N_6364,N_6859);
or U7663 (N_7663,N_6282,N_6823);
nand U7664 (N_7664,N_6159,N_6921);
nand U7665 (N_7665,N_6482,N_6887);
nand U7666 (N_7666,N_6435,N_6985);
and U7667 (N_7667,N_6311,N_6285);
or U7668 (N_7668,N_6899,N_6271);
nand U7669 (N_7669,N_6695,N_6897);
and U7670 (N_7670,N_6932,N_6997);
nor U7671 (N_7671,N_6815,N_6425);
or U7672 (N_7672,N_6057,N_6552);
xnor U7673 (N_7673,N_6991,N_6264);
xnor U7674 (N_7674,N_6700,N_6218);
xnor U7675 (N_7675,N_6950,N_6850);
and U7676 (N_7676,N_6368,N_6068);
and U7677 (N_7677,N_6907,N_6698);
nand U7678 (N_7678,N_6339,N_6517);
xnor U7679 (N_7679,N_6164,N_6942);
or U7680 (N_7680,N_6727,N_6615);
and U7681 (N_7681,N_6174,N_6025);
nand U7682 (N_7682,N_6085,N_6545);
and U7683 (N_7683,N_6137,N_6661);
xor U7684 (N_7684,N_6072,N_6601);
xor U7685 (N_7685,N_6049,N_6014);
nor U7686 (N_7686,N_6448,N_6798);
and U7687 (N_7687,N_6796,N_6900);
and U7688 (N_7688,N_6593,N_6036);
xnor U7689 (N_7689,N_6426,N_6578);
nand U7690 (N_7690,N_6227,N_6587);
xnor U7691 (N_7691,N_6689,N_6808);
and U7692 (N_7692,N_6270,N_6169);
and U7693 (N_7693,N_6600,N_6669);
xor U7694 (N_7694,N_6571,N_6808);
nand U7695 (N_7695,N_6981,N_6839);
xnor U7696 (N_7696,N_6765,N_6985);
xor U7697 (N_7697,N_6713,N_6716);
and U7698 (N_7698,N_6674,N_6379);
and U7699 (N_7699,N_6425,N_6801);
xnor U7700 (N_7700,N_6718,N_6244);
or U7701 (N_7701,N_6507,N_6709);
and U7702 (N_7702,N_6047,N_6750);
nor U7703 (N_7703,N_6814,N_6184);
nor U7704 (N_7704,N_6613,N_6789);
nand U7705 (N_7705,N_6660,N_6506);
or U7706 (N_7706,N_6982,N_6088);
or U7707 (N_7707,N_6399,N_6952);
nor U7708 (N_7708,N_6270,N_6353);
xor U7709 (N_7709,N_6769,N_6080);
or U7710 (N_7710,N_6100,N_6559);
xor U7711 (N_7711,N_6396,N_6782);
xnor U7712 (N_7712,N_6579,N_6300);
nand U7713 (N_7713,N_6936,N_6110);
xor U7714 (N_7714,N_6380,N_6056);
nand U7715 (N_7715,N_6512,N_6715);
nor U7716 (N_7716,N_6505,N_6273);
and U7717 (N_7717,N_6801,N_6217);
or U7718 (N_7718,N_6546,N_6034);
xnor U7719 (N_7719,N_6409,N_6243);
xor U7720 (N_7720,N_6816,N_6121);
xor U7721 (N_7721,N_6260,N_6877);
or U7722 (N_7722,N_6772,N_6516);
nand U7723 (N_7723,N_6540,N_6533);
xnor U7724 (N_7724,N_6245,N_6641);
nand U7725 (N_7725,N_6436,N_6406);
nor U7726 (N_7726,N_6150,N_6675);
or U7727 (N_7727,N_6606,N_6668);
nand U7728 (N_7728,N_6786,N_6055);
and U7729 (N_7729,N_6332,N_6729);
nand U7730 (N_7730,N_6030,N_6459);
and U7731 (N_7731,N_6318,N_6435);
or U7732 (N_7732,N_6927,N_6919);
nor U7733 (N_7733,N_6731,N_6527);
or U7734 (N_7734,N_6033,N_6593);
nor U7735 (N_7735,N_6263,N_6779);
nor U7736 (N_7736,N_6864,N_6707);
nand U7737 (N_7737,N_6252,N_6301);
nand U7738 (N_7738,N_6157,N_6074);
nor U7739 (N_7739,N_6323,N_6042);
and U7740 (N_7740,N_6987,N_6253);
and U7741 (N_7741,N_6351,N_6557);
xnor U7742 (N_7742,N_6095,N_6733);
nor U7743 (N_7743,N_6075,N_6034);
or U7744 (N_7744,N_6167,N_6117);
xnor U7745 (N_7745,N_6538,N_6404);
nor U7746 (N_7746,N_6051,N_6004);
nor U7747 (N_7747,N_6744,N_6434);
nor U7748 (N_7748,N_6344,N_6507);
nand U7749 (N_7749,N_6688,N_6074);
and U7750 (N_7750,N_6635,N_6826);
nor U7751 (N_7751,N_6262,N_6283);
nor U7752 (N_7752,N_6265,N_6827);
and U7753 (N_7753,N_6845,N_6024);
nand U7754 (N_7754,N_6925,N_6009);
nor U7755 (N_7755,N_6699,N_6129);
nand U7756 (N_7756,N_6194,N_6107);
xor U7757 (N_7757,N_6992,N_6003);
nand U7758 (N_7758,N_6777,N_6845);
nor U7759 (N_7759,N_6317,N_6849);
and U7760 (N_7760,N_6521,N_6406);
and U7761 (N_7761,N_6373,N_6992);
xor U7762 (N_7762,N_6370,N_6137);
nor U7763 (N_7763,N_6551,N_6813);
or U7764 (N_7764,N_6219,N_6077);
xnor U7765 (N_7765,N_6754,N_6024);
xor U7766 (N_7766,N_6549,N_6024);
nand U7767 (N_7767,N_6050,N_6786);
nand U7768 (N_7768,N_6217,N_6652);
nor U7769 (N_7769,N_6717,N_6358);
nand U7770 (N_7770,N_6486,N_6201);
or U7771 (N_7771,N_6240,N_6329);
nor U7772 (N_7772,N_6037,N_6406);
nor U7773 (N_7773,N_6838,N_6707);
nor U7774 (N_7774,N_6787,N_6827);
nand U7775 (N_7775,N_6683,N_6816);
nor U7776 (N_7776,N_6318,N_6239);
or U7777 (N_7777,N_6364,N_6105);
xnor U7778 (N_7778,N_6828,N_6589);
nand U7779 (N_7779,N_6670,N_6932);
or U7780 (N_7780,N_6662,N_6423);
xor U7781 (N_7781,N_6486,N_6063);
nor U7782 (N_7782,N_6618,N_6438);
nor U7783 (N_7783,N_6143,N_6114);
and U7784 (N_7784,N_6965,N_6421);
nor U7785 (N_7785,N_6824,N_6386);
or U7786 (N_7786,N_6697,N_6555);
xnor U7787 (N_7787,N_6097,N_6975);
nor U7788 (N_7788,N_6253,N_6147);
xor U7789 (N_7789,N_6099,N_6485);
nand U7790 (N_7790,N_6784,N_6419);
and U7791 (N_7791,N_6070,N_6442);
nand U7792 (N_7792,N_6720,N_6240);
nand U7793 (N_7793,N_6198,N_6458);
or U7794 (N_7794,N_6864,N_6754);
nor U7795 (N_7795,N_6509,N_6483);
nor U7796 (N_7796,N_6002,N_6989);
or U7797 (N_7797,N_6107,N_6817);
nand U7798 (N_7798,N_6169,N_6410);
nor U7799 (N_7799,N_6738,N_6150);
or U7800 (N_7800,N_6337,N_6771);
nor U7801 (N_7801,N_6443,N_6114);
nor U7802 (N_7802,N_6574,N_6306);
nand U7803 (N_7803,N_6890,N_6075);
nor U7804 (N_7804,N_6271,N_6120);
and U7805 (N_7805,N_6519,N_6990);
or U7806 (N_7806,N_6182,N_6170);
and U7807 (N_7807,N_6615,N_6245);
xnor U7808 (N_7808,N_6741,N_6582);
and U7809 (N_7809,N_6696,N_6361);
xnor U7810 (N_7810,N_6595,N_6754);
and U7811 (N_7811,N_6934,N_6916);
nand U7812 (N_7812,N_6104,N_6632);
or U7813 (N_7813,N_6347,N_6713);
nand U7814 (N_7814,N_6399,N_6553);
and U7815 (N_7815,N_6986,N_6389);
and U7816 (N_7816,N_6424,N_6517);
nor U7817 (N_7817,N_6230,N_6888);
and U7818 (N_7818,N_6049,N_6589);
nor U7819 (N_7819,N_6084,N_6533);
nand U7820 (N_7820,N_6195,N_6131);
xnor U7821 (N_7821,N_6470,N_6334);
xor U7822 (N_7822,N_6010,N_6461);
and U7823 (N_7823,N_6520,N_6828);
or U7824 (N_7824,N_6120,N_6109);
or U7825 (N_7825,N_6747,N_6183);
nor U7826 (N_7826,N_6542,N_6259);
xnor U7827 (N_7827,N_6240,N_6931);
xnor U7828 (N_7828,N_6154,N_6161);
nor U7829 (N_7829,N_6048,N_6928);
and U7830 (N_7830,N_6245,N_6917);
or U7831 (N_7831,N_6849,N_6944);
and U7832 (N_7832,N_6027,N_6938);
xnor U7833 (N_7833,N_6780,N_6048);
nor U7834 (N_7834,N_6692,N_6042);
nor U7835 (N_7835,N_6280,N_6734);
nand U7836 (N_7836,N_6357,N_6185);
and U7837 (N_7837,N_6306,N_6732);
nor U7838 (N_7838,N_6469,N_6958);
or U7839 (N_7839,N_6387,N_6312);
or U7840 (N_7840,N_6049,N_6797);
or U7841 (N_7841,N_6825,N_6554);
and U7842 (N_7842,N_6521,N_6508);
nor U7843 (N_7843,N_6968,N_6770);
xnor U7844 (N_7844,N_6061,N_6277);
nor U7845 (N_7845,N_6152,N_6101);
and U7846 (N_7846,N_6643,N_6269);
nand U7847 (N_7847,N_6008,N_6307);
and U7848 (N_7848,N_6204,N_6867);
xnor U7849 (N_7849,N_6784,N_6065);
nand U7850 (N_7850,N_6110,N_6787);
xor U7851 (N_7851,N_6251,N_6168);
nor U7852 (N_7852,N_6533,N_6019);
nor U7853 (N_7853,N_6327,N_6022);
xnor U7854 (N_7854,N_6002,N_6696);
nand U7855 (N_7855,N_6614,N_6741);
nor U7856 (N_7856,N_6976,N_6613);
nor U7857 (N_7857,N_6472,N_6862);
nand U7858 (N_7858,N_6861,N_6002);
nor U7859 (N_7859,N_6149,N_6777);
xor U7860 (N_7860,N_6310,N_6500);
or U7861 (N_7861,N_6025,N_6341);
nor U7862 (N_7862,N_6814,N_6678);
or U7863 (N_7863,N_6022,N_6440);
nor U7864 (N_7864,N_6498,N_6797);
or U7865 (N_7865,N_6834,N_6623);
or U7866 (N_7866,N_6736,N_6231);
or U7867 (N_7867,N_6787,N_6905);
and U7868 (N_7868,N_6608,N_6724);
and U7869 (N_7869,N_6448,N_6044);
nor U7870 (N_7870,N_6903,N_6570);
and U7871 (N_7871,N_6783,N_6140);
nor U7872 (N_7872,N_6977,N_6079);
or U7873 (N_7873,N_6261,N_6791);
xnor U7874 (N_7874,N_6087,N_6557);
xor U7875 (N_7875,N_6188,N_6579);
xor U7876 (N_7876,N_6758,N_6588);
nor U7877 (N_7877,N_6352,N_6128);
xor U7878 (N_7878,N_6782,N_6912);
or U7879 (N_7879,N_6153,N_6966);
nor U7880 (N_7880,N_6863,N_6456);
and U7881 (N_7881,N_6907,N_6195);
or U7882 (N_7882,N_6013,N_6113);
nand U7883 (N_7883,N_6760,N_6917);
nand U7884 (N_7884,N_6490,N_6211);
xnor U7885 (N_7885,N_6182,N_6932);
nor U7886 (N_7886,N_6269,N_6514);
or U7887 (N_7887,N_6401,N_6137);
nor U7888 (N_7888,N_6289,N_6082);
nor U7889 (N_7889,N_6591,N_6010);
xnor U7890 (N_7890,N_6642,N_6236);
nor U7891 (N_7891,N_6186,N_6544);
and U7892 (N_7892,N_6301,N_6064);
nand U7893 (N_7893,N_6951,N_6662);
xnor U7894 (N_7894,N_6853,N_6919);
xnor U7895 (N_7895,N_6153,N_6470);
or U7896 (N_7896,N_6510,N_6793);
nand U7897 (N_7897,N_6518,N_6918);
xnor U7898 (N_7898,N_6801,N_6469);
nor U7899 (N_7899,N_6447,N_6054);
nor U7900 (N_7900,N_6615,N_6297);
or U7901 (N_7901,N_6575,N_6599);
nor U7902 (N_7902,N_6693,N_6906);
and U7903 (N_7903,N_6828,N_6167);
nand U7904 (N_7904,N_6764,N_6377);
nand U7905 (N_7905,N_6517,N_6340);
or U7906 (N_7906,N_6916,N_6471);
and U7907 (N_7907,N_6989,N_6503);
and U7908 (N_7908,N_6736,N_6216);
nand U7909 (N_7909,N_6014,N_6841);
and U7910 (N_7910,N_6673,N_6092);
nand U7911 (N_7911,N_6080,N_6240);
and U7912 (N_7912,N_6011,N_6588);
or U7913 (N_7913,N_6325,N_6464);
or U7914 (N_7914,N_6886,N_6823);
nor U7915 (N_7915,N_6387,N_6131);
nor U7916 (N_7916,N_6232,N_6605);
nand U7917 (N_7917,N_6507,N_6001);
xnor U7918 (N_7918,N_6812,N_6316);
and U7919 (N_7919,N_6557,N_6161);
and U7920 (N_7920,N_6180,N_6658);
xnor U7921 (N_7921,N_6476,N_6586);
nand U7922 (N_7922,N_6669,N_6228);
xor U7923 (N_7923,N_6081,N_6418);
or U7924 (N_7924,N_6179,N_6609);
and U7925 (N_7925,N_6862,N_6606);
nand U7926 (N_7926,N_6381,N_6082);
or U7927 (N_7927,N_6944,N_6144);
xnor U7928 (N_7928,N_6868,N_6609);
or U7929 (N_7929,N_6341,N_6644);
xor U7930 (N_7930,N_6731,N_6351);
and U7931 (N_7931,N_6342,N_6193);
nor U7932 (N_7932,N_6357,N_6166);
nand U7933 (N_7933,N_6460,N_6993);
and U7934 (N_7934,N_6863,N_6265);
nor U7935 (N_7935,N_6998,N_6607);
nand U7936 (N_7936,N_6427,N_6773);
and U7937 (N_7937,N_6745,N_6908);
xor U7938 (N_7938,N_6542,N_6574);
or U7939 (N_7939,N_6664,N_6907);
nor U7940 (N_7940,N_6056,N_6066);
nor U7941 (N_7941,N_6298,N_6730);
and U7942 (N_7942,N_6933,N_6830);
nor U7943 (N_7943,N_6711,N_6301);
or U7944 (N_7944,N_6060,N_6828);
nand U7945 (N_7945,N_6543,N_6740);
xnor U7946 (N_7946,N_6787,N_6121);
nand U7947 (N_7947,N_6586,N_6059);
nand U7948 (N_7948,N_6890,N_6884);
nor U7949 (N_7949,N_6148,N_6050);
and U7950 (N_7950,N_6117,N_6760);
xnor U7951 (N_7951,N_6685,N_6651);
nor U7952 (N_7952,N_6556,N_6852);
nor U7953 (N_7953,N_6714,N_6109);
and U7954 (N_7954,N_6129,N_6790);
or U7955 (N_7955,N_6097,N_6441);
and U7956 (N_7956,N_6972,N_6819);
and U7957 (N_7957,N_6785,N_6972);
or U7958 (N_7958,N_6689,N_6880);
nor U7959 (N_7959,N_6040,N_6780);
or U7960 (N_7960,N_6662,N_6664);
or U7961 (N_7961,N_6696,N_6013);
xnor U7962 (N_7962,N_6373,N_6494);
and U7963 (N_7963,N_6741,N_6389);
nor U7964 (N_7964,N_6097,N_6095);
xor U7965 (N_7965,N_6264,N_6915);
nand U7966 (N_7966,N_6778,N_6689);
nor U7967 (N_7967,N_6474,N_6996);
nand U7968 (N_7968,N_6214,N_6430);
nand U7969 (N_7969,N_6411,N_6174);
xnor U7970 (N_7970,N_6711,N_6607);
nand U7971 (N_7971,N_6099,N_6959);
and U7972 (N_7972,N_6439,N_6547);
nor U7973 (N_7973,N_6616,N_6090);
xnor U7974 (N_7974,N_6553,N_6656);
and U7975 (N_7975,N_6549,N_6428);
nand U7976 (N_7976,N_6837,N_6303);
nor U7977 (N_7977,N_6889,N_6762);
and U7978 (N_7978,N_6714,N_6363);
nor U7979 (N_7979,N_6401,N_6447);
or U7980 (N_7980,N_6393,N_6073);
and U7981 (N_7981,N_6451,N_6094);
and U7982 (N_7982,N_6662,N_6670);
nor U7983 (N_7983,N_6345,N_6378);
nor U7984 (N_7984,N_6950,N_6797);
or U7985 (N_7985,N_6254,N_6008);
xnor U7986 (N_7986,N_6948,N_6899);
nand U7987 (N_7987,N_6119,N_6262);
or U7988 (N_7988,N_6882,N_6402);
or U7989 (N_7989,N_6620,N_6170);
nand U7990 (N_7990,N_6647,N_6785);
and U7991 (N_7991,N_6913,N_6102);
or U7992 (N_7992,N_6098,N_6629);
and U7993 (N_7993,N_6500,N_6365);
and U7994 (N_7994,N_6288,N_6490);
xnor U7995 (N_7995,N_6207,N_6698);
nand U7996 (N_7996,N_6052,N_6602);
nor U7997 (N_7997,N_6389,N_6001);
or U7998 (N_7998,N_6541,N_6962);
and U7999 (N_7999,N_6604,N_6520);
nand U8000 (N_8000,N_7728,N_7770);
nand U8001 (N_8001,N_7972,N_7699);
xor U8002 (N_8002,N_7226,N_7193);
nand U8003 (N_8003,N_7706,N_7351);
xor U8004 (N_8004,N_7129,N_7067);
nor U8005 (N_8005,N_7813,N_7059);
nor U8006 (N_8006,N_7923,N_7230);
nand U8007 (N_8007,N_7619,N_7611);
nor U8008 (N_8008,N_7063,N_7383);
or U8009 (N_8009,N_7371,N_7055);
nor U8010 (N_8010,N_7103,N_7707);
xor U8011 (N_8011,N_7773,N_7431);
xnor U8012 (N_8012,N_7427,N_7280);
and U8013 (N_8013,N_7057,N_7519);
xnor U8014 (N_8014,N_7962,N_7062);
or U8015 (N_8015,N_7152,N_7325);
nor U8016 (N_8016,N_7704,N_7856);
and U8017 (N_8017,N_7549,N_7612);
or U8018 (N_8018,N_7092,N_7889);
or U8019 (N_8019,N_7981,N_7645);
nand U8020 (N_8020,N_7228,N_7281);
nor U8021 (N_8021,N_7698,N_7974);
and U8022 (N_8022,N_7732,N_7462);
nor U8023 (N_8023,N_7410,N_7158);
nand U8024 (N_8024,N_7591,N_7545);
nor U8025 (N_8025,N_7454,N_7581);
and U8026 (N_8026,N_7747,N_7742);
nand U8027 (N_8027,N_7763,N_7366);
or U8028 (N_8028,N_7328,N_7276);
and U8029 (N_8029,N_7234,N_7621);
or U8030 (N_8030,N_7093,N_7458);
or U8031 (N_8031,N_7133,N_7620);
nor U8032 (N_8032,N_7583,N_7385);
and U8033 (N_8033,N_7177,N_7329);
xor U8034 (N_8034,N_7102,N_7758);
and U8035 (N_8035,N_7888,N_7041);
or U8036 (N_8036,N_7484,N_7195);
xnor U8037 (N_8037,N_7561,N_7126);
or U8038 (N_8038,N_7210,N_7712);
xor U8039 (N_8039,N_7899,N_7941);
nor U8040 (N_8040,N_7687,N_7378);
or U8041 (N_8041,N_7927,N_7904);
xor U8042 (N_8042,N_7364,N_7594);
and U8043 (N_8043,N_7844,N_7425);
or U8044 (N_8044,N_7944,N_7933);
and U8045 (N_8045,N_7413,N_7219);
nand U8046 (N_8046,N_7926,N_7155);
nor U8047 (N_8047,N_7039,N_7402);
or U8048 (N_8048,N_7022,N_7843);
xor U8049 (N_8049,N_7789,N_7816);
nand U8050 (N_8050,N_7984,N_7331);
and U8051 (N_8051,N_7876,N_7991);
nand U8052 (N_8052,N_7377,N_7068);
nand U8053 (N_8053,N_7223,N_7100);
nand U8054 (N_8054,N_7287,N_7541);
nand U8055 (N_8055,N_7029,N_7358);
and U8056 (N_8056,N_7426,N_7250);
nor U8057 (N_8057,N_7920,N_7942);
nand U8058 (N_8058,N_7081,N_7394);
xnor U8059 (N_8059,N_7001,N_7298);
nand U8060 (N_8060,N_7428,N_7143);
nand U8061 (N_8061,N_7389,N_7162);
or U8062 (N_8062,N_7064,N_7811);
and U8063 (N_8063,N_7714,N_7603);
and U8064 (N_8064,N_7648,N_7930);
nand U8065 (N_8065,N_7472,N_7890);
nand U8066 (N_8066,N_7205,N_7750);
or U8067 (N_8067,N_7830,N_7047);
nor U8068 (N_8068,N_7360,N_7967);
and U8069 (N_8069,N_7312,N_7913);
xor U8070 (N_8070,N_7640,N_7797);
or U8071 (N_8071,N_7236,N_7467);
nand U8072 (N_8072,N_7679,N_7649);
nand U8073 (N_8073,N_7352,N_7632);
nor U8074 (N_8074,N_7660,N_7282);
nor U8075 (N_8075,N_7496,N_7490);
or U8076 (N_8076,N_7900,N_7852);
nor U8077 (N_8077,N_7015,N_7662);
or U8078 (N_8078,N_7993,N_7269);
xor U8079 (N_8079,N_7979,N_7782);
or U8080 (N_8080,N_7863,N_7183);
or U8081 (N_8081,N_7909,N_7414);
nor U8082 (N_8082,N_7809,N_7300);
nand U8083 (N_8083,N_7301,N_7424);
xnor U8084 (N_8084,N_7864,N_7135);
or U8085 (N_8085,N_7638,N_7585);
or U8086 (N_8086,N_7992,N_7453);
xnor U8087 (N_8087,N_7723,N_7566);
xor U8088 (N_8088,N_7990,N_7589);
xnor U8089 (N_8089,N_7542,N_7370);
nand U8090 (N_8090,N_7161,N_7829);
or U8091 (N_8091,N_7036,N_7422);
and U8092 (N_8092,N_7895,N_7249);
or U8093 (N_8093,N_7340,N_7266);
xnor U8094 (N_8094,N_7186,N_7051);
xor U8095 (N_8095,N_7500,N_7988);
nor U8096 (N_8096,N_7008,N_7290);
and U8097 (N_8097,N_7049,N_7615);
or U8098 (N_8098,N_7802,N_7908);
or U8099 (N_8099,N_7762,N_7602);
or U8100 (N_8100,N_7845,N_7697);
nor U8101 (N_8101,N_7609,N_7271);
nand U8102 (N_8102,N_7877,N_7673);
nand U8103 (N_8103,N_7518,N_7606);
and U8104 (N_8104,N_7480,N_7634);
nor U8105 (N_8105,N_7828,N_7626);
nor U8106 (N_8106,N_7316,N_7091);
and U8107 (N_8107,N_7191,N_7918);
nor U8108 (N_8108,N_7213,N_7775);
or U8109 (N_8109,N_7009,N_7246);
nand U8110 (N_8110,N_7071,N_7175);
xnor U8111 (N_8111,N_7463,N_7465);
xor U8112 (N_8112,N_7898,N_7344);
nand U8113 (N_8113,N_7817,N_7263);
or U8114 (N_8114,N_7995,N_7444);
or U8115 (N_8115,N_7089,N_7869);
nor U8116 (N_8116,N_7169,N_7952);
nand U8117 (N_8117,N_7715,N_7043);
or U8118 (N_8118,N_7517,N_7503);
or U8119 (N_8119,N_7450,N_7885);
nand U8120 (N_8120,N_7491,N_7087);
xnor U8121 (N_8121,N_7224,N_7790);
xor U8122 (N_8122,N_7363,N_7504);
nand U8123 (N_8123,N_7215,N_7556);
nand U8124 (N_8124,N_7243,N_7073);
xnor U8125 (N_8125,N_7421,N_7973);
or U8126 (N_8126,N_7105,N_7115);
and U8127 (N_8127,N_7806,N_7744);
and U8128 (N_8128,N_7357,N_7456);
xnor U8129 (N_8129,N_7189,N_7310);
or U8130 (N_8130,N_7268,N_7074);
nand U8131 (N_8131,N_7576,N_7145);
nand U8132 (N_8132,N_7875,N_7292);
and U8133 (N_8133,N_7661,N_7146);
nor U8134 (N_8134,N_7674,N_7185);
and U8135 (N_8135,N_7006,N_7823);
and U8136 (N_8136,N_7408,N_7940);
nor U8137 (N_8137,N_7886,N_7586);
or U8138 (N_8138,N_7842,N_7018);
or U8139 (N_8139,N_7231,N_7168);
or U8140 (N_8140,N_7173,N_7451);
xor U8141 (N_8141,N_7359,N_7880);
xnor U8142 (N_8142,N_7655,N_7297);
and U8143 (N_8143,N_7957,N_7977);
xor U8144 (N_8144,N_7682,N_7666);
and U8145 (N_8145,N_7767,N_7148);
xor U8146 (N_8146,N_7535,N_7031);
nor U8147 (N_8147,N_7954,N_7857);
xor U8148 (N_8148,N_7324,N_7999);
and U8149 (N_8149,N_7724,N_7562);
and U8150 (N_8150,N_7070,N_7590);
nor U8151 (N_8151,N_7733,N_7283);
or U8152 (N_8152,N_7379,N_7931);
xnor U8153 (N_8153,N_7532,N_7505);
xor U8154 (N_8154,N_7752,N_7274);
xnor U8155 (N_8155,N_7194,N_7448);
xor U8156 (N_8156,N_7212,N_7819);
xor U8157 (N_8157,N_7065,N_7851);
nand U8158 (N_8158,N_7664,N_7207);
or U8159 (N_8159,N_7859,N_7313);
and U8160 (N_8160,N_7582,N_7232);
or U8161 (N_8161,N_7172,N_7607);
or U8162 (N_8162,N_7044,N_7179);
and U8163 (N_8163,N_7771,N_7601);
xnor U8164 (N_8164,N_7635,N_7220);
or U8165 (N_8165,N_7110,N_7007);
or U8166 (N_8166,N_7537,N_7291);
nor U8167 (N_8167,N_7711,N_7253);
or U8168 (N_8168,N_7305,N_7384);
or U8169 (N_8169,N_7214,N_7306);
nand U8170 (N_8170,N_7761,N_7021);
nand U8171 (N_8171,N_7037,N_7111);
or U8172 (N_8172,N_7373,N_7987);
or U8173 (N_8173,N_7746,N_7641);
and U8174 (N_8174,N_7457,N_7112);
nor U8175 (N_8175,N_7256,N_7109);
and U8176 (N_8176,N_7947,N_7150);
xnor U8177 (N_8177,N_7137,N_7080);
and U8178 (N_8178,N_7552,N_7240);
nand U8179 (N_8179,N_7964,N_7865);
nor U8180 (N_8180,N_7748,N_7053);
nor U8181 (N_8181,N_7182,N_7437);
nor U8182 (N_8182,N_7891,N_7798);
and U8183 (N_8183,N_7989,N_7337);
and U8184 (N_8184,N_7369,N_7754);
nor U8185 (N_8185,N_7099,N_7709);
nor U8186 (N_8186,N_7855,N_7795);
and U8187 (N_8187,N_7116,N_7046);
and U8188 (N_8188,N_7343,N_7393);
and U8189 (N_8189,N_7184,N_7722);
nand U8190 (N_8190,N_7630,N_7409);
and U8191 (N_8191,N_7639,N_7882);
xnor U8192 (N_8192,N_7095,N_7285);
xnor U8193 (N_8193,N_7710,N_7976);
nor U8194 (N_8194,N_7516,N_7834);
nand U8195 (N_8195,N_7739,N_7468);
or U8196 (N_8196,N_7494,N_7951);
and U8197 (N_8197,N_7027,N_7959);
or U8198 (N_8198,N_7289,N_7832);
and U8199 (N_8199,N_7629,N_7368);
or U8200 (N_8200,N_7440,N_7356);
or U8201 (N_8201,N_7814,N_7163);
or U8202 (N_8202,N_7555,N_7314);
and U8203 (N_8203,N_7956,N_7235);
nand U8204 (N_8204,N_7076,N_7793);
and U8205 (N_8205,N_7060,N_7523);
nand U8206 (N_8206,N_7592,N_7040);
xnor U8207 (N_8207,N_7983,N_7906);
nor U8208 (N_8208,N_7320,N_7005);
nand U8209 (N_8209,N_7689,N_7716);
nor U8210 (N_8210,N_7106,N_7831);
nor U8211 (N_8211,N_7125,N_7361);
nand U8212 (N_8212,N_7565,N_7692);
xor U8213 (N_8213,N_7200,N_7245);
nand U8214 (N_8214,N_7769,N_7050);
nor U8215 (N_8215,N_7508,N_7872);
nand U8216 (N_8216,N_7078,N_7753);
or U8217 (N_8217,N_7244,N_7669);
xnor U8218 (N_8218,N_7934,N_7209);
xnor U8219 (N_8219,N_7618,N_7493);
or U8220 (N_8220,N_7760,N_7558);
nand U8221 (N_8221,N_7738,N_7052);
and U8222 (N_8222,N_7391,N_7252);
or U8223 (N_8223,N_7751,N_7731);
nand U8224 (N_8224,N_7788,N_7960);
nor U8225 (N_8225,N_7735,N_7072);
or U8226 (N_8226,N_7084,N_7905);
and U8227 (N_8227,N_7211,N_7570);
nor U8228 (N_8228,N_7997,N_7097);
and U8229 (N_8229,N_7094,N_7154);
xnor U8230 (N_8230,N_7435,N_7013);
and U8231 (N_8231,N_7251,N_7725);
nor U8232 (N_8232,N_7141,N_7568);
nor U8233 (N_8233,N_7935,N_7002);
nor U8234 (N_8234,N_7376,N_7800);
nand U8235 (N_8235,N_7943,N_7878);
nand U8236 (N_8236,N_7395,N_7339);
and U8237 (N_8237,N_7239,N_7515);
and U8238 (N_8238,N_7330,N_7970);
xor U8239 (N_8239,N_7447,N_7955);
nand U8240 (N_8240,N_7659,N_7190);
or U8241 (N_8241,N_7308,N_7557);
nor U8242 (N_8242,N_7347,N_7432);
nor U8243 (N_8243,N_7799,N_7196);
and U8244 (N_8244,N_7489,N_7833);
nand U8245 (N_8245,N_7916,N_7117);
nor U8246 (N_8246,N_7866,N_7780);
xnor U8247 (N_8247,N_7374,N_7077);
or U8248 (N_8248,N_7466,N_7350);
nand U8249 (N_8249,N_7333,N_7783);
nor U8250 (N_8250,N_7971,N_7255);
and U8251 (N_8251,N_7726,N_7404);
xor U8252 (N_8252,N_7528,N_7538);
xor U8253 (N_8253,N_7501,N_7694);
nor U8254 (N_8254,N_7530,N_7805);
xor U8255 (N_8255,N_7014,N_7151);
xor U8256 (N_8256,N_7627,N_7729);
nor U8257 (N_8257,N_7965,N_7939);
nor U8258 (N_8258,N_7020,N_7569);
or U8259 (N_8259,N_7691,N_7871);
or U8260 (N_8260,N_7262,N_7108);
and U8261 (N_8261,N_7654,N_7187);
and U8262 (N_8262,N_7381,N_7642);
nand U8263 (N_8263,N_7804,N_7142);
or U8264 (N_8264,N_7417,N_7225);
and U8265 (N_8265,N_7375,N_7085);
nor U8266 (N_8266,N_7838,N_7327);
xor U8267 (N_8267,N_7884,N_7550);
and U8268 (N_8268,N_7840,N_7610);
xor U8269 (N_8269,N_7901,N_7958);
nand U8270 (N_8270,N_7846,N_7120);
xnor U8271 (N_8271,N_7636,N_7968);
and U8272 (N_8272,N_7524,N_7708);
or U8273 (N_8273,N_7123,N_7577);
and U8274 (N_8274,N_7171,N_7925);
or U8275 (N_8275,N_7267,N_7304);
and U8276 (N_8276,N_7801,N_7907);
xor U8277 (N_8277,N_7665,N_7676);
or U8278 (N_8278,N_7513,N_7443);
and U8279 (N_8279,N_7222,N_7403);
and U8280 (N_8280,N_7392,N_7030);
or U8281 (N_8281,N_7719,N_7862);
nor U8282 (N_8282,N_7588,N_7487);
or U8283 (N_8283,N_7396,N_7406);
xor U8284 (N_8284,N_7631,N_7218);
nor U8285 (N_8285,N_7915,N_7743);
nand U8286 (N_8286,N_7338,N_7362);
nand U8287 (N_8287,N_7273,N_7946);
and U8288 (N_8288,N_7703,N_7953);
nand U8289 (N_8289,N_7867,N_7288);
nand U8290 (N_8290,N_7257,N_7647);
nor U8291 (N_8291,N_7580,N_7779);
nand U8292 (N_8292,N_7045,N_7159);
nor U8293 (N_8293,N_7420,N_7003);
or U8294 (N_8294,N_7756,N_7605);
or U8295 (N_8295,N_7121,N_7663);
xnor U8296 (N_8296,N_7309,N_7341);
or U8297 (N_8297,N_7579,N_7336);
or U8298 (N_8298,N_7405,N_7319);
xor U8299 (N_8299,N_7140,N_7028);
nor U8300 (N_8300,N_7452,N_7157);
xnor U8301 (N_8301,N_7459,N_7994);
or U8302 (N_8302,N_7672,N_7502);
nand U8303 (N_8303,N_7737,N_7894);
xnor U8304 (N_8304,N_7668,N_7104);
nand U8305 (N_8305,N_7278,N_7181);
xnor U8306 (N_8306,N_7734,N_7938);
nor U8307 (N_8307,N_7345,N_7492);
nand U8308 (N_8308,N_7980,N_7717);
nor U8309 (N_8309,N_7048,N_7054);
xnor U8310 (N_8310,N_7386,N_7471);
nand U8311 (N_8311,N_7026,N_7096);
or U8312 (N_8312,N_7688,N_7657);
nor U8313 (N_8313,N_7841,N_7460);
or U8314 (N_8314,N_7353,N_7613);
and U8315 (N_8315,N_7066,N_7924);
or U8316 (N_8316,N_7132,N_7033);
nor U8317 (N_8317,N_7608,N_7765);
xor U8318 (N_8318,N_7397,N_7367);
nand U8319 (N_8319,N_7398,N_7810);
and U8320 (N_8320,N_7893,N_7826);
nor U8321 (N_8321,N_7348,N_7265);
nand U8322 (N_8322,N_7985,N_7270);
xor U8323 (N_8323,N_7670,N_7461);
nor U8324 (N_8324,N_7896,N_7936);
or U8325 (N_8325,N_7578,N_7587);
nor U8326 (N_8326,N_7966,N_7778);
nor U8327 (N_8327,N_7149,N_7527);
xnor U8328 (N_8328,N_7416,N_7260);
nand U8329 (N_8329,N_7540,N_7922);
xnor U8330 (N_8330,N_7533,N_7593);
xnor U8331 (N_8331,N_7208,N_7777);
xnor U8332 (N_8332,N_7643,N_7418);
or U8333 (N_8333,N_7791,N_7019);
nand U8334 (N_8334,N_7919,N_7766);
nor U8335 (N_8335,N_7727,N_7702);
nand U8336 (N_8336,N_7010,N_7004);
and U8337 (N_8337,N_7180,N_7623);
xnor U8338 (N_8338,N_7914,N_7476);
nor U8339 (N_8339,N_7101,N_7982);
xnor U8340 (N_8340,N_7512,N_7658);
xnor U8341 (N_8341,N_7883,N_7430);
xor U8342 (N_8342,N_7713,N_7318);
and U8343 (N_8343,N_7488,N_7616);
nand U8344 (N_8344,N_7881,N_7796);
xor U8345 (N_8345,N_7238,N_7061);
nand U8346 (N_8346,N_7812,N_7975);
or U8347 (N_8347,N_7848,N_7677);
xor U8348 (N_8348,N_7012,N_7614);
nor U8349 (N_8349,N_7241,N_7628);
nand U8350 (N_8350,N_7365,N_7521);
and U8351 (N_8351,N_7113,N_7911);
or U8352 (N_8352,N_7701,N_7474);
xor U8353 (N_8353,N_7441,N_7445);
and U8354 (N_8354,N_7204,N_7617);
and U8355 (N_8355,N_7407,N_7870);
or U8356 (N_8356,N_7794,N_7134);
nand U8357 (N_8357,N_7575,N_7622);
or U8358 (N_8358,N_7025,N_7399);
and U8359 (N_8359,N_7509,N_7595);
or U8360 (N_8360,N_7573,N_7653);
and U8361 (N_8361,N_7625,N_7455);
or U8362 (N_8362,N_7317,N_7860);
or U8363 (N_8363,N_7247,N_7144);
xnor U8364 (N_8364,N_7963,N_7695);
xnor U8365 (N_8365,N_7434,N_7685);
xnor U8366 (N_8366,N_7229,N_7335);
or U8367 (N_8367,N_7948,N_7429);
xnor U8368 (N_8368,N_7671,N_7449);
nor U8369 (N_8369,N_7740,N_7165);
or U8370 (N_8370,N_7174,N_7887);
or U8371 (N_8371,N_7294,N_7721);
nor U8372 (N_8372,N_7675,N_7536);
nand U8373 (N_8373,N_7083,N_7107);
nor U8374 (N_8374,N_7127,N_7478);
or U8375 (N_8375,N_7700,N_7510);
nand U8376 (N_8376,N_7481,N_7693);
xor U8377 (N_8377,N_7929,N_7815);
or U8378 (N_8378,N_7600,N_7529);
xnor U8379 (N_8379,N_7824,N_7201);
and U8380 (N_8380,N_7526,N_7138);
nand U8381 (N_8381,N_7683,N_7854);
or U8382 (N_8382,N_7950,N_7818);
and U8383 (N_8383,N_7439,N_7130);
or U8384 (N_8384,N_7650,N_7254);
and U8385 (N_8385,N_7539,N_7741);
or U8386 (N_8386,N_7903,N_7604);
xnor U8387 (N_8387,N_7075,N_7221);
and U8388 (N_8388,N_7264,N_7868);
nand U8389 (N_8389,N_7119,N_7544);
nor U8390 (N_8390,N_7961,N_7299);
nor U8391 (N_8391,N_7122,N_7902);
or U8392 (N_8392,N_7118,N_7412);
and U8393 (N_8393,N_7035,N_7598);
xor U8394 (N_8394,N_7419,N_7438);
xnor U8395 (N_8395,N_7216,N_7757);
nand U8396 (N_8396,N_7825,N_7563);
or U8397 (N_8397,N_7446,N_7473);
nor U8398 (N_8398,N_7258,N_7346);
xnor U8399 (N_8399,N_7322,N_7293);
nor U8400 (N_8400,N_7038,N_7202);
nand U8401 (N_8401,N_7560,N_7433);
nand U8402 (N_8402,N_7522,N_7633);
or U8403 (N_8403,N_7442,N_7114);
nand U8404 (N_8404,N_7978,N_7786);
xor U8405 (N_8405,N_7482,N_7032);
xor U8406 (N_8406,N_7917,N_7355);
nand U8407 (N_8407,N_7277,N_7847);
and U8408 (N_8408,N_7525,N_7197);
or U8409 (N_8409,N_7511,N_7090);
nor U8410 (N_8410,N_7497,N_7764);
or U8411 (N_8411,N_7259,N_7928);
and U8412 (N_8412,N_7275,N_7772);
nor U8413 (N_8413,N_7949,N_7514);
nor U8414 (N_8414,N_7332,N_7464);
nor U8415 (N_8415,N_7969,N_7506);
or U8416 (N_8416,N_7996,N_7837);
nor U8417 (N_8417,N_7380,N_7910);
nand U8418 (N_8418,N_7861,N_7156);
or U8419 (N_8419,N_7774,N_7166);
xor U8420 (N_8420,N_7567,N_7646);
nand U8421 (N_8421,N_7088,N_7198);
nand U8422 (N_8422,N_7387,N_7534);
or U8423 (N_8423,N_7768,N_7597);
xor U8424 (N_8424,N_7932,N_7543);
and U8425 (N_8425,N_7897,N_7034);
nor U8426 (N_8426,N_7736,N_7787);
or U8427 (N_8427,N_7199,N_7827);
and U8428 (N_8428,N_7718,N_7307);
nand U8429 (N_8429,N_7921,N_7164);
and U8430 (N_8430,N_7296,N_7176);
nor U8431 (N_8431,N_7551,N_7242);
nor U8432 (N_8432,N_7520,N_7781);
and U8433 (N_8433,N_7599,N_7853);
nand U8434 (N_8434,N_7874,N_7637);
or U8435 (N_8435,N_7153,N_7667);
or U8436 (N_8436,N_7696,N_7279);
or U8437 (N_8437,N_7261,N_7056);
xnor U8438 (N_8438,N_7124,N_7086);
or U8439 (N_8439,N_7286,N_7479);
nor U8440 (N_8440,N_7401,N_7192);
xor U8441 (N_8441,N_7303,N_7098);
or U8442 (N_8442,N_7839,N_7058);
or U8443 (N_8443,N_7720,N_7507);
nor U8444 (N_8444,N_7690,N_7559);
nand U8445 (N_8445,N_7564,N_7820);
nand U8446 (N_8446,N_7656,N_7469);
nand U8447 (N_8447,N_7553,N_7400);
xnor U8448 (N_8448,N_7749,N_7167);
nand U8449 (N_8449,N_7785,N_7024);
nor U8450 (N_8450,N_7349,N_7548);
and U8451 (N_8451,N_7016,N_7069);
and U8452 (N_8452,N_7571,N_7188);
xor U8453 (N_8453,N_7784,N_7485);
nor U8454 (N_8454,N_7334,N_7079);
xnor U8455 (N_8455,N_7372,N_7326);
nand U8456 (N_8456,N_7596,N_7237);
and U8457 (N_8457,N_7082,N_7477);
nand U8458 (N_8458,N_7295,N_7531);
and U8459 (N_8459,N_7284,N_7705);
nand U8460 (N_8460,N_7745,N_7986);
nor U8461 (N_8461,N_7546,N_7217);
nand U8462 (N_8462,N_7354,N_7233);
or U8463 (N_8463,N_7792,N_7203);
nand U8464 (N_8464,N_7776,N_7547);
nor U8465 (N_8465,N_7011,N_7342);
nor U8466 (N_8466,N_7835,N_7390);
xnor U8467 (N_8467,N_7821,N_7486);
nor U8468 (N_8468,N_7170,N_7023);
nand U8469 (N_8469,N_7302,N_7498);
or U8470 (N_8470,N_7998,N_7136);
xor U8471 (N_8471,N_7206,N_7139);
nand U8472 (N_8472,N_7808,N_7945);
and U8473 (N_8473,N_7873,N_7272);
xor U8474 (N_8474,N_7730,N_7686);
xor U8475 (N_8475,N_7892,N_7311);
nor U8476 (N_8476,N_7131,N_7554);
nand U8477 (N_8477,N_7572,N_7836);
nor U8478 (N_8478,N_7803,N_7912);
nor U8479 (N_8479,N_7584,N_7017);
nor U8480 (N_8480,N_7680,N_7644);
nor U8481 (N_8481,N_7624,N_7000);
xor U8482 (N_8482,N_7755,N_7495);
nor U8483 (N_8483,N_7411,N_7475);
nor U8484 (N_8484,N_7128,N_7499);
and U8485 (N_8485,N_7415,N_7807);
or U8486 (N_8486,N_7483,N_7849);
and U8487 (N_8487,N_7248,N_7042);
and U8488 (N_8488,N_7759,N_7423);
nand U8489 (N_8489,N_7227,N_7681);
or U8490 (N_8490,N_7388,N_7937);
xnor U8491 (N_8491,N_7678,N_7850);
nand U8492 (N_8492,N_7652,N_7147);
or U8493 (N_8493,N_7879,N_7684);
or U8494 (N_8494,N_7321,N_7315);
nand U8495 (N_8495,N_7323,N_7858);
nor U8496 (N_8496,N_7160,N_7574);
and U8497 (N_8497,N_7178,N_7651);
nor U8498 (N_8498,N_7436,N_7822);
xnor U8499 (N_8499,N_7470,N_7382);
nor U8500 (N_8500,N_7954,N_7036);
nor U8501 (N_8501,N_7340,N_7739);
nand U8502 (N_8502,N_7045,N_7788);
nand U8503 (N_8503,N_7355,N_7175);
and U8504 (N_8504,N_7786,N_7135);
nand U8505 (N_8505,N_7412,N_7686);
or U8506 (N_8506,N_7381,N_7003);
nand U8507 (N_8507,N_7271,N_7424);
and U8508 (N_8508,N_7881,N_7527);
and U8509 (N_8509,N_7238,N_7113);
and U8510 (N_8510,N_7556,N_7115);
nand U8511 (N_8511,N_7115,N_7810);
xor U8512 (N_8512,N_7307,N_7143);
nor U8513 (N_8513,N_7433,N_7272);
nand U8514 (N_8514,N_7570,N_7004);
xor U8515 (N_8515,N_7733,N_7621);
and U8516 (N_8516,N_7375,N_7358);
and U8517 (N_8517,N_7670,N_7414);
nor U8518 (N_8518,N_7831,N_7723);
nor U8519 (N_8519,N_7235,N_7714);
nor U8520 (N_8520,N_7730,N_7751);
and U8521 (N_8521,N_7379,N_7770);
and U8522 (N_8522,N_7166,N_7547);
or U8523 (N_8523,N_7390,N_7576);
nor U8524 (N_8524,N_7138,N_7073);
nor U8525 (N_8525,N_7348,N_7454);
xnor U8526 (N_8526,N_7730,N_7066);
nand U8527 (N_8527,N_7672,N_7676);
and U8528 (N_8528,N_7199,N_7668);
nand U8529 (N_8529,N_7255,N_7167);
nor U8530 (N_8530,N_7807,N_7643);
xor U8531 (N_8531,N_7381,N_7301);
nor U8532 (N_8532,N_7228,N_7313);
nand U8533 (N_8533,N_7479,N_7809);
nand U8534 (N_8534,N_7102,N_7465);
nand U8535 (N_8535,N_7470,N_7496);
and U8536 (N_8536,N_7468,N_7011);
or U8537 (N_8537,N_7609,N_7760);
nor U8538 (N_8538,N_7219,N_7629);
xor U8539 (N_8539,N_7059,N_7065);
xor U8540 (N_8540,N_7095,N_7920);
nand U8541 (N_8541,N_7391,N_7928);
and U8542 (N_8542,N_7418,N_7783);
or U8543 (N_8543,N_7275,N_7277);
nand U8544 (N_8544,N_7814,N_7221);
and U8545 (N_8545,N_7727,N_7118);
or U8546 (N_8546,N_7078,N_7756);
or U8547 (N_8547,N_7301,N_7595);
or U8548 (N_8548,N_7272,N_7369);
nor U8549 (N_8549,N_7126,N_7803);
and U8550 (N_8550,N_7471,N_7720);
nand U8551 (N_8551,N_7660,N_7526);
xnor U8552 (N_8552,N_7601,N_7197);
nor U8553 (N_8553,N_7654,N_7210);
and U8554 (N_8554,N_7485,N_7200);
and U8555 (N_8555,N_7958,N_7306);
or U8556 (N_8556,N_7465,N_7333);
and U8557 (N_8557,N_7135,N_7512);
xor U8558 (N_8558,N_7805,N_7307);
nand U8559 (N_8559,N_7142,N_7248);
or U8560 (N_8560,N_7172,N_7133);
or U8561 (N_8561,N_7370,N_7195);
xnor U8562 (N_8562,N_7631,N_7191);
nand U8563 (N_8563,N_7981,N_7589);
or U8564 (N_8564,N_7153,N_7726);
or U8565 (N_8565,N_7832,N_7660);
or U8566 (N_8566,N_7614,N_7651);
and U8567 (N_8567,N_7042,N_7023);
and U8568 (N_8568,N_7358,N_7946);
nor U8569 (N_8569,N_7459,N_7021);
or U8570 (N_8570,N_7028,N_7888);
xor U8571 (N_8571,N_7079,N_7792);
or U8572 (N_8572,N_7634,N_7895);
and U8573 (N_8573,N_7570,N_7772);
or U8574 (N_8574,N_7567,N_7570);
and U8575 (N_8575,N_7239,N_7839);
xnor U8576 (N_8576,N_7599,N_7954);
nand U8577 (N_8577,N_7774,N_7300);
nor U8578 (N_8578,N_7008,N_7090);
and U8579 (N_8579,N_7058,N_7984);
or U8580 (N_8580,N_7975,N_7725);
nor U8581 (N_8581,N_7539,N_7106);
nor U8582 (N_8582,N_7561,N_7951);
or U8583 (N_8583,N_7463,N_7839);
and U8584 (N_8584,N_7271,N_7159);
or U8585 (N_8585,N_7728,N_7236);
xnor U8586 (N_8586,N_7746,N_7223);
or U8587 (N_8587,N_7563,N_7722);
xnor U8588 (N_8588,N_7824,N_7617);
nand U8589 (N_8589,N_7455,N_7557);
and U8590 (N_8590,N_7946,N_7204);
nand U8591 (N_8591,N_7320,N_7774);
xor U8592 (N_8592,N_7092,N_7886);
nor U8593 (N_8593,N_7027,N_7593);
and U8594 (N_8594,N_7615,N_7291);
and U8595 (N_8595,N_7544,N_7150);
and U8596 (N_8596,N_7261,N_7263);
nor U8597 (N_8597,N_7742,N_7618);
and U8598 (N_8598,N_7072,N_7157);
nand U8599 (N_8599,N_7444,N_7265);
nand U8600 (N_8600,N_7450,N_7087);
nor U8601 (N_8601,N_7303,N_7685);
xor U8602 (N_8602,N_7012,N_7051);
nand U8603 (N_8603,N_7642,N_7267);
nor U8604 (N_8604,N_7176,N_7129);
xor U8605 (N_8605,N_7517,N_7605);
nand U8606 (N_8606,N_7418,N_7954);
or U8607 (N_8607,N_7062,N_7349);
nand U8608 (N_8608,N_7837,N_7278);
nor U8609 (N_8609,N_7574,N_7539);
or U8610 (N_8610,N_7413,N_7918);
xor U8611 (N_8611,N_7177,N_7333);
or U8612 (N_8612,N_7649,N_7085);
nand U8613 (N_8613,N_7205,N_7611);
or U8614 (N_8614,N_7713,N_7993);
nand U8615 (N_8615,N_7533,N_7172);
or U8616 (N_8616,N_7668,N_7750);
and U8617 (N_8617,N_7040,N_7427);
xnor U8618 (N_8618,N_7805,N_7336);
or U8619 (N_8619,N_7870,N_7711);
or U8620 (N_8620,N_7631,N_7246);
nor U8621 (N_8621,N_7647,N_7644);
or U8622 (N_8622,N_7012,N_7372);
xor U8623 (N_8623,N_7121,N_7399);
nand U8624 (N_8624,N_7797,N_7433);
or U8625 (N_8625,N_7259,N_7884);
nand U8626 (N_8626,N_7339,N_7024);
xnor U8627 (N_8627,N_7450,N_7553);
nand U8628 (N_8628,N_7742,N_7481);
nand U8629 (N_8629,N_7547,N_7908);
xnor U8630 (N_8630,N_7037,N_7040);
or U8631 (N_8631,N_7348,N_7351);
nand U8632 (N_8632,N_7631,N_7411);
nand U8633 (N_8633,N_7643,N_7591);
nor U8634 (N_8634,N_7311,N_7564);
and U8635 (N_8635,N_7672,N_7213);
xnor U8636 (N_8636,N_7051,N_7262);
xnor U8637 (N_8637,N_7933,N_7561);
xor U8638 (N_8638,N_7178,N_7084);
or U8639 (N_8639,N_7225,N_7438);
or U8640 (N_8640,N_7694,N_7078);
or U8641 (N_8641,N_7802,N_7626);
xnor U8642 (N_8642,N_7960,N_7666);
and U8643 (N_8643,N_7982,N_7184);
nand U8644 (N_8644,N_7941,N_7107);
nor U8645 (N_8645,N_7856,N_7144);
nor U8646 (N_8646,N_7434,N_7004);
nor U8647 (N_8647,N_7045,N_7210);
xnor U8648 (N_8648,N_7648,N_7021);
nand U8649 (N_8649,N_7160,N_7923);
and U8650 (N_8650,N_7239,N_7430);
nor U8651 (N_8651,N_7101,N_7837);
nand U8652 (N_8652,N_7884,N_7895);
xor U8653 (N_8653,N_7781,N_7012);
nor U8654 (N_8654,N_7733,N_7086);
nand U8655 (N_8655,N_7529,N_7104);
nand U8656 (N_8656,N_7295,N_7346);
nand U8657 (N_8657,N_7757,N_7742);
or U8658 (N_8658,N_7696,N_7776);
or U8659 (N_8659,N_7545,N_7061);
nor U8660 (N_8660,N_7893,N_7937);
or U8661 (N_8661,N_7126,N_7331);
nor U8662 (N_8662,N_7467,N_7775);
or U8663 (N_8663,N_7212,N_7355);
nor U8664 (N_8664,N_7769,N_7855);
xor U8665 (N_8665,N_7765,N_7454);
or U8666 (N_8666,N_7297,N_7159);
or U8667 (N_8667,N_7397,N_7647);
or U8668 (N_8668,N_7208,N_7794);
nor U8669 (N_8669,N_7704,N_7288);
nand U8670 (N_8670,N_7484,N_7420);
xnor U8671 (N_8671,N_7885,N_7193);
or U8672 (N_8672,N_7278,N_7474);
nand U8673 (N_8673,N_7496,N_7789);
and U8674 (N_8674,N_7116,N_7061);
xnor U8675 (N_8675,N_7144,N_7373);
nor U8676 (N_8676,N_7690,N_7317);
or U8677 (N_8677,N_7545,N_7700);
nand U8678 (N_8678,N_7971,N_7475);
xor U8679 (N_8679,N_7596,N_7300);
nor U8680 (N_8680,N_7334,N_7350);
xnor U8681 (N_8681,N_7524,N_7481);
nand U8682 (N_8682,N_7254,N_7181);
nand U8683 (N_8683,N_7994,N_7191);
nand U8684 (N_8684,N_7254,N_7124);
or U8685 (N_8685,N_7548,N_7395);
or U8686 (N_8686,N_7471,N_7559);
and U8687 (N_8687,N_7342,N_7716);
xor U8688 (N_8688,N_7656,N_7059);
nor U8689 (N_8689,N_7784,N_7491);
or U8690 (N_8690,N_7038,N_7175);
and U8691 (N_8691,N_7031,N_7461);
nand U8692 (N_8692,N_7950,N_7683);
nand U8693 (N_8693,N_7939,N_7245);
nor U8694 (N_8694,N_7180,N_7881);
and U8695 (N_8695,N_7618,N_7915);
or U8696 (N_8696,N_7460,N_7484);
or U8697 (N_8697,N_7816,N_7834);
nand U8698 (N_8698,N_7533,N_7423);
or U8699 (N_8699,N_7710,N_7330);
xnor U8700 (N_8700,N_7549,N_7865);
nand U8701 (N_8701,N_7025,N_7867);
nor U8702 (N_8702,N_7717,N_7419);
or U8703 (N_8703,N_7506,N_7321);
or U8704 (N_8704,N_7270,N_7956);
nand U8705 (N_8705,N_7489,N_7352);
xor U8706 (N_8706,N_7625,N_7714);
or U8707 (N_8707,N_7728,N_7388);
xnor U8708 (N_8708,N_7066,N_7237);
or U8709 (N_8709,N_7545,N_7687);
xor U8710 (N_8710,N_7777,N_7412);
xnor U8711 (N_8711,N_7163,N_7860);
nor U8712 (N_8712,N_7182,N_7770);
or U8713 (N_8713,N_7733,N_7540);
nor U8714 (N_8714,N_7726,N_7640);
or U8715 (N_8715,N_7464,N_7098);
xnor U8716 (N_8716,N_7551,N_7899);
nand U8717 (N_8717,N_7934,N_7125);
nand U8718 (N_8718,N_7741,N_7579);
nor U8719 (N_8719,N_7070,N_7883);
and U8720 (N_8720,N_7356,N_7361);
nor U8721 (N_8721,N_7484,N_7669);
or U8722 (N_8722,N_7545,N_7624);
nand U8723 (N_8723,N_7113,N_7143);
xor U8724 (N_8724,N_7990,N_7069);
nor U8725 (N_8725,N_7010,N_7319);
nand U8726 (N_8726,N_7662,N_7981);
nor U8727 (N_8727,N_7670,N_7109);
nand U8728 (N_8728,N_7787,N_7588);
nand U8729 (N_8729,N_7320,N_7533);
xor U8730 (N_8730,N_7915,N_7052);
xnor U8731 (N_8731,N_7466,N_7433);
nor U8732 (N_8732,N_7198,N_7683);
or U8733 (N_8733,N_7435,N_7547);
and U8734 (N_8734,N_7152,N_7839);
nor U8735 (N_8735,N_7670,N_7848);
nand U8736 (N_8736,N_7864,N_7717);
nand U8737 (N_8737,N_7921,N_7811);
nor U8738 (N_8738,N_7105,N_7175);
nor U8739 (N_8739,N_7875,N_7038);
or U8740 (N_8740,N_7042,N_7511);
xor U8741 (N_8741,N_7596,N_7395);
nand U8742 (N_8742,N_7388,N_7978);
nand U8743 (N_8743,N_7418,N_7284);
nand U8744 (N_8744,N_7958,N_7411);
nor U8745 (N_8745,N_7212,N_7433);
nand U8746 (N_8746,N_7515,N_7273);
nand U8747 (N_8747,N_7575,N_7920);
and U8748 (N_8748,N_7196,N_7180);
or U8749 (N_8749,N_7325,N_7773);
or U8750 (N_8750,N_7829,N_7758);
nor U8751 (N_8751,N_7869,N_7176);
nand U8752 (N_8752,N_7606,N_7072);
or U8753 (N_8753,N_7922,N_7891);
nor U8754 (N_8754,N_7736,N_7131);
or U8755 (N_8755,N_7495,N_7627);
nand U8756 (N_8756,N_7038,N_7110);
nand U8757 (N_8757,N_7941,N_7163);
or U8758 (N_8758,N_7935,N_7605);
and U8759 (N_8759,N_7883,N_7439);
nor U8760 (N_8760,N_7976,N_7453);
or U8761 (N_8761,N_7068,N_7062);
nand U8762 (N_8762,N_7042,N_7270);
and U8763 (N_8763,N_7866,N_7538);
nand U8764 (N_8764,N_7147,N_7385);
or U8765 (N_8765,N_7338,N_7361);
and U8766 (N_8766,N_7023,N_7802);
or U8767 (N_8767,N_7922,N_7545);
or U8768 (N_8768,N_7234,N_7690);
xnor U8769 (N_8769,N_7156,N_7173);
nor U8770 (N_8770,N_7021,N_7908);
or U8771 (N_8771,N_7990,N_7092);
nor U8772 (N_8772,N_7117,N_7084);
nor U8773 (N_8773,N_7660,N_7643);
xor U8774 (N_8774,N_7596,N_7462);
nor U8775 (N_8775,N_7066,N_7928);
xnor U8776 (N_8776,N_7380,N_7113);
nand U8777 (N_8777,N_7317,N_7668);
xnor U8778 (N_8778,N_7070,N_7375);
xor U8779 (N_8779,N_7790,N_7152);
and U8780 (N_8780,N_7717,N_7004);
or U8781 (N_8781,N_7757,N_7476);
nand U8782 (N_8782,N_7828,N_7417);
or U8783 (N_8783,N_7357,N_7530);
and U8784 (N_8784,N_7525,N_7719);
nor U8785 (N_8785,N_7925,N_7727);
xor U8786 (N_8786,N_7573,N_7650);
nor U8787 (N_8787,N_7709,N_7227);
or U8788 (N_8788,N_7384,N_7484);
nor U8789 (N_8789,N_7007,N_7471);
xor U8790 (N_8790,N_7547,N_7718);
nand U8791 (N_8791,N_7930,N_7203);
or U8792 (N_8792,N_7094,N_7513);
or U8793 (N_8793,N_7022,N_7944);
nand U8794 (N_8794,N_7855,N_7518);
xnor U8795 (N_8795,N_7982,N_7324);
and U8796 (N_8796,N_7812,N_7000);
xnor U8797 (N_8797,N_7826,N_7700);
nor U8798 (N_8798,N_7895,N_7863);
xor U8799 (N_8799,N_7560,N_7370);
or U8800 (N_8800,N_7474,N_7040);
nor U8801 (N_8801,N_7701,N_7597);
nor U8802 (N_8802,N_7249,N_7923);
and U8803 (N_8803,N_7352,N_7172);
and U8804 (N_8804,N_7184,N_7191);
nor U8805 (N_8805,N_7465,N_7864);
nor U8806 (N_8806,N_7048,N_7180);
or U8807 (N_8807,N_7230,N_7008);
or U8808 (N_8808,N_7543,N_7915);
and U8809 (N_8809,N_7549,N_7407);
xnor U8810 (N_8810,N_7741,N_7250);
xnor U8811 (N_8811,N_7596,N_7071);
or U8812 (N_8812,N_7499,N_7816);
or U8813 (N_8813,N_7299,N_7059);
or U8814 (N_8814,N_7959,N_7005);
nand U8815 (N_8815,N_7710,N_7961);
or U8816 (N_8816,N_7645,N_7920);
xor U8817 (N_8817,N_7289,N_7451);
nand U8818 (N_8818,N_7715,N_7826);
or U8819 (N_8819,N_7751,N_7915);
nor U8820 (N_8820,N_7102,N_7270);
and U8821 (N_8821,N_7571,N_7106);
or U8822 (N_8822,N_7556,N_7816);
or U8823 (N_8823,N_7712,N_7693);
or U8824 (N_8824,N_7024,N_7641);
xor U8825 (N_8825,N_7044,N_7194);
and U8826 (N_8826,N_7220,N_7068);
nor U8827 (N_8827,N_7528,N_7133);
nand U8828 (N_8828,N_7929,N_7816);
nor U8829 (N_8829,N_7536,N_7178);
and U8830 (N_8830,N_7046,N_7088);
or U8831 (N_8831,N_7017,N_7606);
xnor U8832 (N_8832,N_7824,N_7207);
and U8833 (N_8833,N_7911,N_7788);
nand U8834 (N_8834,N_7266,N_7747);
or U8835 (N_8835,N_7487,N_7099);
nand U8836 (N_8836,N_7612,N_7501);
nand U8837 (N_8837,N_7925,N_7659);
or U8838 (N_8838,N_7576,N_7839);
or U8839 (N_8839,N_7643,N_7506);
nand U8840 (N_8840,N_7215,N_7860);
or U8841 (N_8841,N_7463,N_7044);
and U8842 (N_8842,N_7215,N_7407);
or U8843 (N_8843,N_7431,N_7728);
nor U8844 (N_8844,N_7747,N_7678);
xor U8845 (N_8845,N_7623,N_7774);
nor U8846 (N_8846,N_7201,N_7909);
nand U8847 (N_8847,N_7713,N_7129);
or U8848 (N_8848,N_7843,N_7285);
nor U8849 (N_8849,N_7276,N_7052);
xor U8850 (N_8850,N_7387,N_7589);
or U8851 (N_8851,N_7611,N_7659);
or U8852 (N_8852,N_7714,N_7076);
nor U8853 (N_8853,N_7055,N_7480);
xor U8854 (N_8854,N_7494,N_7386);
or U8855 (N_8855,N_7318,N_7388);
nand U8856 (N_8856,N_7053,N_7471);
and U8857 (N_8857,N_7222,N_7323);
or U8858 (N_8858,N_7980,N_7312);
or U8859 (N_8859,N_7164,N_7584);
nand U8860 (N_8860,N_7418,N_7699);
and U8861 (N_8861,N_7548,N_7259);
xor U8862 (N_8862,N_7022,N_7340);
nand U8863 (N_8863,N_7454,N_7247);
and U8864 (N_8864,N_7531,N_7329);
and U8865 (N_8865,N_7979,N_7937);
nor U8866 (N_8866,N_7341,N_7673);
or U8867 (N_8867,N_7352,N_7328);
xnor U8868 (N_8868,N_7615,N_7453);
xor U8869 (N_8869,N_7451,N_7814);
xnor U8870 (N_8870,N_7208,N_7683);
nand U8871 (N_8871,N_7872,N_7494);
xor U8872 (N_8872,N_7978,N_7490);
nand U8873 (N_8873,N_7792,N_7076);
nor U8874 (N_8874,N_7371,N_7661);
and U8875 (N_8875,N_7086,N_7118);
xnor U8876 (N_8876,N_7771,N_7677);
nor U8877 (N_8877,N_7598,N_7727);
nand U8878 (N_8878,N_7954,N_7570);
xor U8879 (N_8879,N_7146,N_7623);
and U8880 (N_8880,N_7461,N_7214);
or U8881 (N_8881,N_7030,N_7621);
xor U8882 (N_8882,N_7178,N_7969);
and U8883 (N_8883,N_7202,N_7225);
and U8884 (N_8884,N_7944,N_7967);
or U8885 (N_8885,N_7087,N_7051);
and U8886 (N_8886,N_7326,N_7381);
nand U8887 (N_8887,N_7132,N_7417);
xnor U8888 (N_8888,N_7427,N_7685);
nor U8889 (N_8889,N_7695,N_7261);
xnor U8890 (N_8890,N_7901,N_7507);
xnor U8891 (N_8891,N_7931,N_7340);
nor U8892 (N_8892,N_7382,N_7502);
nor U8893 (N_8893,N_7462,N_7887);
nand U8894 (N_8894,N_7090,N_7400);
and U8895 (N_8895,N_7306,N_7663);
and U8896 (N_8896,N_7859,N_7484);
nand U8897 (N_8897,N_7040,N_7850);
xnor U8898 (N_8898,N_7624,N_7837);
nand U8899 (N_8899,N_7535,N_7042);
nand U8900 (N_8900,N_7276,N_7101);
xnor U8901 (N_8901,N_7546,N_7006);
and U8902 (N_8902,N_7859,N_7222);
xor U8903 (N_8903,N_7701,N_7128);
nor U8904 (N_8904,N_7811,N_7430);
nand U8905 (N_8905,N_7513,N_7257);
and U8906 (N_8906,N_7735,N_7757);
and U8907 (N_8907,N_7082,N_7985);
nand U8908 (N_8908,N_7753,N_7051);
or U8909 (N_8909,N_7842,N_7175);
xnor U8910 (N_8910,N_7310,N_7858);
or U8911 (N_8911,N_7456,N_7365);
and U8912 (N_8912,N_7045,N_7560);
or U8913 (N_8913,N_7904,N_7801);
or U8914 (N_8914,N_7734,N_7496);
or U8915 (N_8915,N_7183,N_7680);
or U8916 (N_8916,N_7110,N_7274);
xnor U8917 (N_8917,N_7040,N_7845);
and U8918 (N_8918,N_7332,N_7063);
nand U8919 (N_8919,N_7413,N_7890);
and U8920 (N_8920,N_7208,N_7291);
nand U8921 (N_8921,N_7735,N_7508);
nor U8922 (N_8922,N_7224,N_7448);
nand U8923 (N_8923,N_7451,N_7327);
nor U8924 (N_8924,N_7863,N_7502);
nor U8925 (N_8925,N_7308,N_7684);
xor U8926 (N_8926,N_7559,N_7894);
nor U8927 (N_8927,N_7497,N_7552);
or U8928 (N_8928,N_7702,N_7742);
xnor U8929 (N_8929,N_7855,N_7585);
or U8930 (N_8930,N_7606,N_7063);
nand U8931 (N_8931,N_7908,N_7730);
xor U8932 (N_8932,N_7926,N_7051);
or U8933 (N_8933,N_7574,N_7755);
xnor U8934 (N_8934,N_7122,N_7662);
or U8935 (N_8935,N_7461,N_7250);
nor U8936 (N_8936,N_7411,N_7035);
xor U8937 (N_8937,N_7351,N_7680);
nor U8938 (N_8938,N_7162,N_7169);
nor U8939 (N_8939,N_7668,N_7442);
xnor U8940 (N_8940,N_7098,N_7404);
nor U8941 (N_8941,N_7516,N_7711);
or U8942 (N_8942,N_7869,N_7347);
and U8943 (N_8943,N_7859,N_7263);
nand U8944 (N_8944,N_7021,N_7980);
or U8945 (N_8945,N_7324,N_7477);
xnor U8946 (N_8946,N_7734,N_7047);
or U8947 (N_8947,N_7309,N_7196);
and U8948 (N_8948,N_7267,N_7777);
xnor U8949 (N_8949,N_7253,N_7009);
xnor U8950 (N_8950,N_7102,N_7355);
xnor U8951 (N_8951,N_7759,N_7697);
nand U8952 (N_8952,N_7250,N_7282);
or U8953 (N_8953,N_7981,N_7456);
nor U8954 (N_8954,N_7276,N_7971);
nand U8955 (N_8955,N_7295,N_7677);
nor U8956 (N_8956,N_7829,N_7374);
and U8957 (N_8957,N_7170,N_7326);
and U8958 (N_8958,N_7790,N_7751);
nand U8959 (N_8959,N_7232,N_7413);
and U8960 (N_8960,N_7744,N_7439);
and U8961 (N_8961,N_7589,N_7193);
xor U8962 (N_8962,N_7475,N_7402);
or U8963 (N_8963,N_7988,N_7117);
nor U8964 (N_8964,N_7834,N_7843);
nand U8965 (N_8965,N_7813,N_7357);
or U8966 (N_8966,N_7369,N_7797);
nand U8967 (N_8967,N_7160,N_7835);
nand U8968 (N_8968,N_7552,N_7612);
and U8969 (N_8969,N_7034,N_7370);
nor U8970 (N_8970,N_7574,N_7670);
nor U8971 (N_8971,N_7295,N_7305);
and U8972 (N_8972,N_7177,N_7290);
and U8973 (N_8973,N_7731,N_7685);
nand U8974 (N_8974,N_7991,N_7272);
nor U8975 (N_8975,N_7507,N_7669);
nor U8976 (N_8976,N_7847,N_7356);
xor U8977 (N_8977,N_7610,N_7670);
nor U8978 (N_8978,N_7691,N_7942);
nor U8979 (N_8979,N_7219,N_7110);
xor U8980 (N_8980,N_7247,N_7112);
or U8981 (N_8981,N_7271,N_7052);
xor U8982 (N_8982,N_7481,N_7034);
and U8983 (N_8983,N_7565,N_7388);
nand U8984 (N_8984,N_7052,N_7167);
xor U8985 (N_8985,N_7724,N_7768);
or U8986 (N_8986,N_7189,N_7263);
xnor U8987 (N_8987,N_7927,N_7455);
xor U8988 (N_8988,N_7524,N_7573);
xor U8989 (N_8989,N_7137,N_7856);
and U8990 (N_8990,N_7248,N_7512);
xor U8991 (N_8991,N_7292,N_7658);
and U8992 (N_8992,N_7465,N_7578);
or U8993 (N_8993,N_7918,N_7061);
nor U8994 (N_8994,N_7961,N_7865);
and U8995 (N_8995,N_7663,N_7436);
nor U8996 (N_8996,N_7587,N_7634);
xnor U8997 (N_8997,N_7401,N_7162);
and U8998 (N_8998,N_7266,N_7278);
xnor U8999 (N_8999,N_7635,N_7767);
or U9000 (N_9000,N_8427,N_8611);
xor U9001 (N_9001,N_8226,N_8652);
xor U9002 (N_9002,N_8367,N_8359);
nand U9003 (N_9003,N_8428,N_8979);
nand U9004 (N_9004,N_8866,N_8386);
xnor U9005 (N_9005,N_8331,N_8655);
and U9006 (N_9006,N_8351,N_8038);
xor U9007 (N_9007,N_8911,N_8947);
nor U9008 (N_9008,N_8784,N_8348);
xor U9009 (N_9009,N_8678,N_8174);
or U9010 (N_9010,N_8531,N_8244);
and U9011 (N_9011,N_8294,N_8301);
xnor U9012 (N_9012,N_8801,N_8315);
nand U9013 (N_9013,N_8568,N_8023);
nand U9014 (N_9014,N_8218,N_8882);
nand U9015 (N_9015,N_8300,N_8070);
nand U9016 (N_9016,N_8977,N_8164);
and U9017 (N_9017,N_8747,N_8610);
and U9018 (N_9018,N_8625,N_8551);
and U9019 (N_9019,N_8021,N_8389);
nor U9020 (N_9020,N_8724,N_8480);
nor U9021 (N_9021,N_8227,N_8131);
nand U9022 (N_9022,N_8970,N_8103);
or U9023 (N_9023,N_8897,N_8371);
and U9024 (N_9024,N_8879,N_8697);
nor U9025 (N_9025,N_8715,N_8566);
nand U9026 (N_9026,N_8250,N_8529);
nand U9027 (N_9027,N_8769,N_8317);
and U9028 (N_9028,N_8790,N_8939);
and U9029 (N_9029,N_8604,N_8425);
nand U9030 (N_9030,N_8653,N_8245);
nor U9031 (N_9031,N_8717,N_8414);
nor U9032 (N_9032,N_8749,N_8114);
and U9033 (N_9033,N_8839,N_8843);
or U9034 (N_9034,N_8100,N_8046);
nand U9035 (N_9035,N_8908,N_8775);
xnor U9036 (N_9036,N_8085,N_8334);
nor U9037 (N_9037,N_8042,N_8436);
xor U9038 (N_9038,N_8370,N_8483);
and U9039 (N_9039,N_8401,N_8881);
xor U9040 (N_9040,N_8829,N_8206);
nor U9041 (N_9041,N_8337,N_8382);
xor U9042 (N_9042,N_8640,N_8745);
xnor U9043 (N_9043,N_8659,N_8589);
nand U9044 (N_9044,N_8274,N_8516);
xnor U9045 (N_9045,N_8402,N_8471);
nor U9046 (N_9046,N_8253,N_8285);
xnor U9047 (N_9047,N_8701,N_8230);
or U9048 (N_9048,N_8209,N_8918);
and U9049 (N_9049,N_8508,N_8913);
xnor U9050 (N_9050,N_8054,N_8433);
xnor U9051 (N_9051,N_8669,N_8109);
or U9052 (N_9052,N_8963,N_8110);
or U9053 (N_9053,N_8132,N_8810);
and U9054 (N_9054,N_8763,N_8290);
and U9055 (N_9055,N_8362,N_8614);
xnor U9056 (N_9056,N_8646,N_8395);
and U9057 (N_9057,N_8107,N_8656);
or U9058 (N_9058,N_8426,N_8242);
nand U9059 (N_9059,N_8251,N_8058);
xor U9060 (N_9060,N_8826,N_8276);
and U9061 (N_9061,N_8437,N_8994);
xnor U9062 (N_9062,N_8845,N_8836);
xor U9063 (N_9063,N_8733,N_8819);
nor U9064 (N_9064,N_8104,N_8378);
nand U9065 (N_9065,N_8357,N_8316);
nor U9066 (N_9066,N_8392,N_8528);
or U9067 (N_9067,N_8720,N_8406);
xor U9068 (N_9068,N_8986,N_8906);
and U9069 (N_9069,N_8592,N_8466);
nand U9070 (N_9070,N_8214,N_8506);
xnor U9071 (N_9071,N_8022,N_8848);
nand U9072 (N_9072,N_8917,N_8945);
and U9073 (N_9073,N_8481,N_8312);
or U9074 (N_9074,N_8014,N_8795);
or U9075 (N_9075,N_8078,N_8309);
xnor U9076 (N_9076,N_8375,N_8598);
nand U9077 (N_9077,N_8940,N_8243);
and U9078 (N_9078,N_8044,N_8187);
xor U9079 (N_9079,N_8412,N_8456);
xnor U9080 (N_9080,N_8034,N_8252);
nor U9081 (N_9081,N_8565,N_8702);
nor U9082 (N_9082,N_8629,N_8522);
nand U9083 (N_9083,N_8295,N_8239);
nor U9084 (N_9084,N_8990,N_8853);
xnor U9085 (N_9085,N_8575,N_8624);
xnor U9086 (N_9086,N_8686,N_8995);
nand U9087 (N_9087,N_8943,N_8518);
nor U9088 (N_9088,N_8479,N_8171);
nand U9089 (N_9089,N_8783,N_8658);
nand U9090 (N_9090,N_8444,N_8088);
xor U9091 (N_9091,N_8605,N_8129);
nor U9092 (N_9092,N_8050,N_8003);
xor U9093 (N_9093,N_8996,N_8883);
or U9094 (N_9094,N_8207,N_8045);
nand U9095 (N_9095,N_8356,N_8649);
or U9096 (N_9096,N_8229,N_8837);
nor U9097 (N_9097,N_8086,N_8677);
and U9098 (N_9098,N_8800,N_8205);
nor U9099 (N_9099,N_8419,N_8993);
and U9100 (N_9100,N_8695,N_8390);
nand U9101 (N_9101,N_8163,N_8318);
and U9102 (N_9102,N_8681,N_8458);
or U9103 (N_9103,N_8024,N_8854);
and U9104 (N_9104,N_8791,N_8139);
nand U9105 (N_9105,N_8018,N_8825);
nor U9106 (N_9106,N_8327,N_8124);
or U9107 (N_9107,N_8588,N_8916);
nor U9108 (N_9108,N_8319,N_8329);
or U9109 (N_9109,N_8519,N_8344);
and U9110 (N_9110,N_8645,N_8012);
or U9111 (N_9111,N_8867,N_8169);
xnor U9112 (N_9112,N_8053,N_8289);
and U9113 (N_9113,N_8496,N_8676);
xor U9114 (N_9114,N_8435,N_8474);
nor U9115 (N_9115,N_8446,N_8929);
and U9116 (N_9116,N_8778,N_8484);
nor U9117 (N_9117,N_8926,N_8950);
nand U9118 (N_9118,N_8079,N_8786);
xnor U9119 (N_9119,N_8280,N_8136);
nand U9120 (N_9120,N_8478,N_8620);
nand U9121 (N_9121,N_8644,N_8776);
or U9122 (N_9122,N_8532,N_8602);
and U9123 (N_9123,N_8524,N_8584);
and U9124 (N_9124,N_8377,N_8748);
nor U9125 (N_9125,N_8912,N_8505);
and U9126 (N_9126,N_8521,N_8666);
nor U9127 (N_9127,N_8056,N_8095);
nand U9128 (N_9128,N_8762,N_8526);
nand U9129 (N_9129,N_8777,N_8254);
and U9130 (N_9130,N_8952,N_8236);
and U9131 (N_9131,N_8743,N_8111);
nor U9132 (N_9132,N_8539,N_8064);
nor U9133 (N_9133,N_8346,N_8661);
xor U9134 (N_9134,N_8320,N_8654);
xor U9135 (N_9135,N_8621,N_8641);
and U9136 (N_9136,N_8313,N_8472);
or U9137 (N_9137,N_8156,N_8262);
nor U9138 (N_9138,N_8513,N_8257);
xor U9139 (N_9139,N_8507,N_8706);
nand U9140 (N_9140,N_8992,N_8158);
nand U9141 (N_9141,N_8739,N_8036);
xnor U9142 (N_9142,N_8121,N_8721);
and U9143 (N_9143,N_8464,N_8974);
xnor U9144 (N_9144,N_8221,N_8647);
nor U9145 (N_9145,N_8544,N_8609);
or U9146 (N_9146,N_8333,N_8905);
nand U9147 (N_9147,N_8664,N_8942);
xnor U9148 (N_9148,N_8851,N_8821);
and U9149 (N_9149,N_8955,N_8190);
nand U9150 (N_9150,N_8219,N_8674);
and U9151 (N_9151,N_8071,N_8149);
xor U9152 (N_9152,N_8953,N_8418);
and U9153 (N_9153,N_8451,N_8092);
nand U9154 (N_9154,N_8284,N_8490);
nor U9155 (N_9155,N_8608,N_8048);
xnor U9156 (N_9156,N_8117,N_8183);
xnor U9157 (N_9157,N_8997,N_8314);
and U9158 (N_9158,N_8090,N_8440);
xnor U9159 (N_9159,N_8411,N_8286);
nand U9160 (N_9160,N_8051,N_8010);
xor U9161 (N_9161,N_8732,N_8693);
and U9162 (N_9162,N_8886,N_8449);
nand U9163 (N_9163,N_8525,N_8146);
and U9164 (N_9164,N_8040,N_8536);
nor U9165 (N_9165,N_8718,N_8765);
nor U9166 (N_9166,N_8865,N_8445);
or U9167 (N_9167,N_8757,N_8384);
and U9168 (N_9168,N_8618,N_8258);
nand U9169 (N_9169,N_8827,N_8511);
or U9170 (N_9170,N_8597,N_8985);
or U9171 (N_9171,N_8059,N_8298);
and U9172 (N_9172,N_8713,N_8862);
xnor U9173 (N_9173,N_8358,N_8961);
xor U9174 (N_9174,N_8751,N_8188);
and U9175 (N_9175,N_8461,N_8328);
or U9176 (N_9176,N_8157,N_8991);
nand U9177 (N_9177,N_8794,N_8208);
and U9178 (N_9178,N_8699,N_8880);
nor U9179 (N_9179,N_8830,N_8273);
and U9180 (N_9180,N_8630,N_8260);
nor U9181 (N_9181,N_8842,N_8944);
or U9182 (N_9182,N_8350,N_8073);
xnor U9183 (N_9183,N_8712,N_8308);
and U9184 (N_9184,N_8907,N_8166);
or U9185 (N_9185,N_8140,N_8971);
nor U9186 (N_9186,N_8075,N_8398);
nand U9187 (N_9187,N_8335,N_8857);
or U9188 (N_9188,N_8213,N_8781);
and U9189 (N_9189,N_8930,N_8583);
nand U9190 (N_9190,N_8416,N_8964);
and U9191 (N_9191,N_8360,N_8192);
or U9192 (N_9192,N_8491,N_8303);
nor U9193 (N_9193,N_8901,N_8723);
and U9194 (N_9194,N_8736,N_8394);
and U9195 (N_9195,N_8409,N_8266);
nor U9196 (N_9196,N_8302,N_8577);
nand U9197 (N_9197,N_8469,N_8694);
or U9198 (N_9198,N_8147,N_8859);
xnor U9199 (N_9199,N_8155,N_8636);
or U9200 (N_9200,N_8580,N_8197);
and U9201 (N_9201,N_8637,N_8138);
xnor U9202 (N_9202,N_8893,N_8161);
nand U9203 (N_9203,N_8980,N_8322);
or U9204 (N_9204,N_8962,N_8613);
and U9205 (N_9205,N_8020,N_8041);
and U9206 (N_9206,N_8601,N_8808);
nand U9207 (N_9207,N_8773,N_8144);
nor U9208 (N_9208,N_8931,N_8112);
nor U9209 (N_9209,N_8366,N_8201);
nand U9210 (N_9210,N_8872,N_8898);
xor U9211 (N_9211,N_8787,N_8987);
nand U9212 (N_9212,N_8581,N_8856);
or U9213 (N_9213,N_8441,N_8269);
nand U9214 (N_9214,N_8855,N_8231);
and U9215 (N_9215,N_8247,N_8607);
nor U9216 (N_9216,N_8307,N_8510);
or U9217 (N_9217,N_8310,N_8013);
nand U9218 (N_9218,N_8560,N_8707);
and U9219 (N_9219,N_8657,N_8049);
and U9220 (N_9220,N_8497,N_8729);
and U9221 (N_9221,N_8016,N_8969);
xor U9222 (N_9222,N_8672,N_8225);
and U9223 (N_9223,N_8332,N_8639);
and U9224 (N_9224,N_8442,N_8069);
or U9225 (N_9225,N_8460,N_8098);
and U9226 (N_9226,N_8126,N_8692);
xor U9227 (N_9227,N_8072,N_8635);
nor U9228 (N_9228,N_8615,N_8113);
and U9229 (N_9229,N_8453,N_8860);
nand U9230 (N_9230,N_8015,N_8871);
nand U9231 (N_9231,N_8582,N_8448);
or U9232 (N_9232,N_8934,N_8026);
and U9233 (N_9233,N_8477,N_8028);
nand U9234 (N_9234,N_8771,N_8336);
nand U9235 (N_9235,N_8503,N_8989);
or U9236 (N_9236,N_8922,N_8162);
and U9237 (N_9237,N_8354,N_8710);
nor U9238 (N_9238,N_8734,N_8740);
and U9239 (N_9239,N_8679,N_8324);
nand U9240 (N_9240,N_8788,N_8181);
nand U9241 (N_9241,N_8704,N_8423);
or U9242 (N_9242,N_8271,N_8530);
or U9243 (N_9243,N_8960,N_8108);
nand U9244 (N_9244,N_8550,N_8540);
nor U9245 (N_9245,N_8793,N_8632);
or U9246 (N_9246,N_8545,N_8616);
or U9247 (N_9247,N_8972,N_8822);
and U9248 (N_9248,N_8556,N_8383);
xor U9249 (N_9249,N_8864,N_8097);
nand U9250 (N_9250,N_8397,N_8204);
or U9251 (N_9251,N_8549,N_8792);
nor U9252 (N_9252,N_8047,N_8730);
nand U9253 (N_9253,N_8287,N_8080);
nor U9254 (N_9254,N_8805,N_8115);
nor U9255 (N_9255,N_8283,N_8339);
and U9256 (N_9256,N_8002,N_8714);
nand U9257 (N_9257,N_8341,N_8145);
nor U9258 (N_9258,N_8809,N_8282);
nor U9259 (N_9259,N_8372,N_8407);
xnor U9260 (N_9260,N_8574,N_8305);
nand U9261 (N_9261,N_8379,N_8415);
xnor U9262 (N_9262,N_8234,N_8703);
or U9263 (N_9263,N_8537,N_8052);
or U9264 (N_9264,N_8921,N_8141);
nor U9265 (N_9265,N_8571,N_8564);
and U9266 (N_9266,N_8746,N_8684);
and U9267 (N_9267,N_8459,N_8224);
xnor U9268 (N_9268,N_8288,N_8936);
xor U9269 (N_9269,N_8999,N_8680);
or U9270 (N_9270,N_8089,N_8179);
nor U9271 (N_9271,N_8489,N_8439);
nand U9272 (N_9272,N_8888,N_8202);
nand U9273 (N_9273,N_8925,N_8828);
nor U9274 (N_9274,N_8265,N_8467);
or U9275 (N_9275,N_8754,N_8199);
nor U9276 (N_9276,N_8281,N_8772);
nor U9277 (N_9277,N_8849,N_8399);
and U9278 (N_9278,N_8454,N_8587);
or U9279 (N_9279,N_8951,N_8761);
and U9280 (N_9280,N_8306,N_8981);
xor U9281 (N_9281,N_8403,N_8626);
nand U9282 (N_9282,N_8420,N_8689);
or U9283 (N_9283,N_8958,N_8065);
nand U9284 (N_9284,N_8178,N_8173);
nor U9285 (N_9285,N_8186,N_8292);
and U9286 (N_9286,N_8259,N_8998);
and U9287 (N_9287,N_8172,N_8846);
and U9288 (N_9288,N_8326,N_8373);
xor U9289 (N_9289,N_8920,N_8184);
and U9290 (N_9290,N_8457,N_8535);
nand U9291 (N_9291,N_8957,N_8685);
and U9292 (N_9292,N_8708,N_8768);
nor U9293 (N_9293,N_8264,N_8009);
nand U9294 (N_9294,N_8812,N_8120);
xor U9295 (N_9295,N_8063,N_8485);
nor U9296 (N_9296,N_8450,N_8128);
or U9297 (N_9297,N_8735,N_8404);
nand U9298 (N_9298,N_8452,N_8083);
or U9299 (N_9299,N_8482,N_8475);
nor U9300 (N_9300,N_8062,N_8594);
xnor U9301 (N_9301,N_8858,N_8542);
nand U9302 (N_9302,N_8638,N_8633);
nor U9303 (N_9303,N_8220,N_8391);
xor U9304 (N_9304,N_8767,N_8758);
nand U9305 (N_9305,N_8180,N_8408);
and U9306 (N_9306,N_8623,N_8538);
or U9307 (N_9307,N_8567,N_8744);
nor U9308 (N_9308,N_8151,N_8068);
or U9309 (N_9309,N_8919,N_8330);
nor U9310 (N_9310,N_8004,N_8241);
nor U9311 (N_9311,N_8338,N_8831);
xnor U9312 (N_9312,N_8727,N_8494);
nand U9313 (N_9313,N_8668,N_8430);
and U9314 (N_9314,N_8385,N_8501);
and U9315 (N_9315,N_8975,N_8554);
and U9316 (N_9316,N_8099,N_8650);
nor U9317 (N_9317,N_8563,N_8593);
or U9318 (N_9318,N_8504,N_8737);
or U9319 (N_9319,N_8820,N_8956);
and U9320 (N_9320,N_8363,N_8082);
and U9321 (N_9321,N_8275,N_8572);
and U9322 (N_9322,N_8585,N_8818);
nor U9323 (N_9323,N_8914,N_8870);
or U9324 (N_9324,N_8473,N_8067);
nor U9325 (N_9325,N_8968,N_8811);
or U9326 (N_9326,N_8782,N_8096);
or U9327 (N_9327,N_8492,N_8802);
xor U9328 (N_9328,N_8691,N_8612);
xor U9329 (N_9329,N_8852,N_8562);
or U9330 (N_9330,N_8586,N_8590);
or U9331 (N_9331,N_8393,N_8033);
xor U9332 (N_9332,N_8682,N_8847);
or U9333 (N_9333,N_8705,N_8248);
and U9334 (N_9334,N_8816,N_8222);
nand U9335 (N_9335,N_8533,N_8591);
or U9336 (N_9336,N_8966,N_8076);
nand U9337 (N_9337,N_8035,N_8277);
and U9338 (N_9338,N_8011,N_8462);
xnor U9339 (N_9339,N_8470,N_8675);
or U9340 (N_9340,N_8698,N_8122);
nand U9341 (N_9341,N_8299,N_8514);
and U9342 (N_9342,N_8885,N_8954);
and U9343 (N_9343,N_8495,N_8753);
xor U9344 (N_9344,N_8025,N_8774);
and U9345 (N_9345,N_8973,N_8487);
and U9346 (N_9346,N_8619,N_8168);
or U9347 (N_9347,N_8892,N_8160);
and U9348 (N_9348,N_8716,N_8832);
and U9349 (N_9349,N_8722,N_8463);
or U9350 (N_9350,N_8493,N_8561);
or U9351 (N_9351,N_8381,N_8130);
and U9352 (N_9352,N_8928,N_8084);
nand U9353 (N_9353,N_8127,N_8240);
nand U9354 (N_9354,N_8750,N_8541);
and U9355 (N_9355,N_8868,N_8291);
and U9356 (N_9356,N_8438,N_8850);
or U9357 (N_9357,N_8643,N_8797);
and U9358 (N_9358,N_8548,N_8387);
xnor U9359 (N_9359,N_8660,N_8364);
nor U9360 (N_9360,N_8833,N_8237);
nand U9361 (N_9361,N_8631,N_8134);
nor U9362 (N_9362,N_8417,N_8671);
xor U9363 (N_9363,N_8352,N_8223);
nor U9364 (N_9364,N_8817,N_8915);
or U9365 (N_9365,N_8941,N_8434);
and U9366 (N_9366,N_8877,N_8967);
and U9367 (N_9367,N_8520,N_8311);
xnor U9368 (N_9368,N_8878,N_8932);
xnor U9369 (N_9369,N_8648,N_8891);
nand U9370 (N_9370,N_8884,N_8909);
nand U9371 (N_9371,N_8074,N_8000);
nor U9372 (N_9372,N_8345,N_8578);
or U9373 (N_9373,N_8861,N_8217);
nor U9374 (N_9374,N_8101,N_8512);
nor U9375 (N_9375,N_8037,N_8876);
nand U9376 (N_9376,N_8509,N_8443);
nor U9377 (N_9377,N_8904,N_8910);
xor U9378 (N_9378,N_8167,N_8796);
nand U9379 (N_9379,N_8628,N_8725);
xor U9380 (N_9380,N_8200,N_8486);
nor U9381 (N_9381,N_8923,N_8106);
or U9382 (N_9382,N_8353,N_8374);
nand U9383 (N_9383,N_8413,N_8185);
and U9384 (N_9384,N_8844,N_8342);
nand U9385 (N_9385,N_8663,N_8978);
xor U9386 (N_9386,N_8949,N_8983);
nor U9387 (N_9387,N_8488,N_8203);
nor U9388 (N_9388,N_8043,N_8573);
nor U9389 (N_9389,N_8742,N_8102);
nand U9390 (N_9390,N_8665,N_8455);
or U9391 (N_9391,N_8424,N_8270);
and U9392 (N_9392,N_8840,N_8400);
or U9393 (N_9393,N_8304,N_8001);
and U9394 (N_9394,N_8600,N_8447);
nor U9395 (N_9395,N_8396,N_8687);
and U9396 (N_9396,N_8150,N_8709);
xor U9397 (N_9397,N_8651,N_8534);
and U9398 (N_9398,N_8125,N_8347);
or U9399 (N_9399,N_8690,N_8711);
or U9400 (N_9400,N_8815,N_8177);
xnor U9401 (N_9401,N_8595,N_8297);
nor U9402 (N_9402,N_8216,N_8933);
and U9403 (N_9403,N_8196,N_8195);
nor U9404 (N_9404,N_8008,N_8133);
nand U9405 (N_9405,N_8803,N_8603);
and U9406 (N_9406,N_8935,N_8365);
and U9407 (N_9407,N_8869,N_8228);
xnor U9408 (N_9408,N_8232,N_8982);
xor U9409 (N_9409,N_8093,N_8077);
and U9410 (N_9410,N_8764,N_8029);
or U9411 (N_9411,N_8546,N_8135);
or U9412 (N_9412,N_8527,N_8343);
and U9413 (N_9413,N_8670,N_8060);
and U9414 (N_9414,N_8938,N_8175);
or U9415 (N_9415,N_8557,N_8116);
or U9416 (N_9416,N_8965,N_8361);
nor U9417 (N_9417,N_8838,N_8642);
and U9418 (N_9418,N_8142,N_8874);
and U9419 (N_9419,N_8606,N_8760);
nand U9420 (N_9420,N_8789,N_8515);
or U9421 (N_9421,N_8355,N_8210);
or U9422 (N_9422,N_8756,N_8006);
nand U9423 (N_9423,N_8032,N_8726);
nand U9424 (N_9424,N_8576,N_8268);
nand U9425 (N_9425,N_8959,N_8321);
xnor U9426 (N_9426,N_8559,N_8895);
xnor U9427 (N_9427,N_8159,N_8176);
and U9428 (N_9428,N_8903,N_8278);
xor U9429 (N_9429,N_8055,N_8017);
nor U9430 (N_9430,N_8799,N_8759);
or U9431 (N_9431,N_8731,N_8081);
nor U9432 (N_9432,N_8937,N_8137);
nor U9433 (N_9433,N_8667,N_8900);
and U9434 (N_9434,N_8215,N_8517);
or U9435 (N_9435,N_8946,N_8388);
nor U9436 (N_9436,N_8779,N_8770);
nor U9437 (N_9437,N_8570,N_8165);
nand U9438 (N_9438,N_8323,N_8766);
or U9439 (N_9439,N_8738,N_8780);
xnor U9440 (N_9440,N_8984,N_8087);
nor U9441 (N_9441,N_8579,N_8523);
or U9442 (N_9442,N_8105,N_8152);
and U9443 (N_9443,N_8804,N_8976);
xnor U9444 (N_9444,N_8118,N_8019);
xor U9445 (N_9445,N_8255,N_8263);
nor U9446 (N_9446,N_8432,N_8148);
xor U9447 (N_9447,N_8182,N_8476);
and U9448 (N_9448,N_8212,N_8368);
nor U9449 (N_9449,N_8189,N_8369);
xnor U9450 (N_9450,N_8823,N_8552);
and U9451 (N_9451,N_8405,N_8547);
nor U9452 (N_9452,N_8700,N_8170);
nand U9453 (N_9453,N_8039,N_8031);
nand U9454 (N_9454,N_8153,N_8814);
xor U9455 (N_9455,N_8755,N_8057);
nand U9456 (N_9456,N_8261,N_8249);
nand U9457 (N_9457,N_8875,N_8785);
nand U9458 (N_9458,N_8143,N_8325);
nand U9459 (N_9459,N_8500,N_8376);
xnor U9460 (N_9460,N_8841,N_8340);
nor U9461 (N_9461,N_8553,N_8431);
nand U9462 (N_9462,N_8027,N_8696);
nand U9463 (N_9463,N_8429,N_8899);
nor U9464 (N_9464,N_8061,N_8465);
nor U9465 (N_9465,N_8617,N_8902);
and U9466 (N_9466,N_8256,N_8627);
nand U9467 (N_9467,N_8502,N_8030);
xnor U9468 (N_9468,N_8296,N_8688);
nand U9469 (N_9469,N_8924,N_8835);
xor U9470 (N_9470,N_8662,N_8123);
xor U9471 (N_9471,N_8555,N_8410);
nor U9472 (N_9472,N_8198,N_8119);
nand U9473 (N_9473,N_8246,N_8728);
or U9474 (N_9474,N_8890,N_8272);
nand U9475 (N_9475,N_8622,N_8896);
nor U9476 (N_9476,N_8558,N_8091);
nor U9477 (N_9477,N_8673,N_8752);
and U9478 (N_9478,N_8235,N_8498);
or U9479 (N_9479,N_8380,N_8741);
xor U9480 (N_9480,N_8233,N_8889);
nor U9481 (N_9481,N_8596,N_8066);
or U9482 (N_9482,N_8421,N_8927);
xor U9483 (N_9483,N_8569,N_8873);
and U9484 (N_9484,N_8293,N_8194);
and U9485 (N_9485,N_8094,N_8887);
or U9486 (N_9486,N_8422,N_8834);
and U9487 (N_9487,N_8634,N_8349);
and U9488 (N_9488,N_8211,N_8279);
and U9489 (N_9489,N_8988,N_8894);
nor U9490 (N_9490,N_8599,N_8807);
and U9491 (N_9491,N_8468,N_8005);
xnor U9492 (N_9492,N_8719,N_8813);
xnor U9493 (N_9493,N_8543,N_8683);
and U9494 (N_9494,N_8007,N_8824);
and U9495 (N_9495,N_8238,N_8798);
nor U9496 (N_9496,N_8193,N_8267);
or U9497 (N_9497,N_8191,N_8154);
or U9498 (N_9498,N_8948,N_8806);
and U9499 (N_9499,N_8499,N_8863);
nor U9500 (N_9500,N_8789,N_8749);
and U9501 (N_9501,N_8544,N_8041);
and U9502 (N_9502,N_8698,N_8433);
nor U9503 (N_9503,N_8000,N_8795);
nor U9504 (N_9504,N_8095,N_8226);
and U9505 (N_9505,N_8301,N_8085);
nand U9506 (N_9506,N_8464,N_8656);
or U9507 (N_9507,N_8454,N_8317);
nand U9508 (N_9508,N_8619,N_8276);
and U9509 (N_9509,N_8558,N_8746);
and U9510 (N_9510,N_8370,N_8108);
or U9511 (N_9511,N_8964,N_8968);
or U9512 (N_9512,N_8997,N_8434);
nor U9513 (N_9513,N_8638,N_8234);
and U9514 (N_9514,N_8040,N_8063);
or U9515 (N_9515,N_8540,N_8891);
or U9516 (N_9516,N_8540,N_8467);
nor U9517 (N_9517,N_8111,N_8278);
or U9518 (N_9518,N_8854,N_8744);
nand U9519 (N_9519,N_8751,N_8785);
or U9520 (N_9520,N_8784,N_8810);
nand U9521 (N_9521,N_8067,N_8528);
or U9522 (N_9522,N_8481,N_8273);
nand U9523 (N_9523,N_8287,N_8735);
xnor U9524 (N_9524,N_8263,N_8940);
nor U9525 (N_9525,N_8911,N_8553);
nand U9526 (N_9526,N_8847,N_8114);
and U9527 (N_9527,N_8321,N_8646);
nand U9528 (N_9528,N_8368,N_8757);
xor U9529 (N_9529,N_8984,N_8377);
xor U9530 (N_9530,N_8362,N_8951);
or U9531 (N_9531,N_8572,N_8217);
or U9532 (N_9532,N_8232,N_8576);
nor U9533 (N_9533,N_8925,N_8263);
nand U9534 (N_9534,N_8278,N_8011);
and U9535 (N_9535,N_8948,N_8367);
xor U9536 (N_9536,N_8285,N_8114);
xor U9537 (N_9537,N_8303,N_8409);
or U9538 (N_9538,N_8249,N_8380);
and U9539 (N_9539,N_8563,N_8191);
nor U9540 (N_9540,N_8138,N_8062);
xnor U9541 (N_9541,N_8574,N_8762);
or U9542 (N_9542,N_8099,N_8199);
and U9543 (N_9543,N_8080,N_8942);
or U9544 (N_9544,N_8286,N_8646);
and U9545 (N_9545,N_8988,N_8258);
nand U9546 (N_9546,N_8719,N_8835);
nand U9547 (N_9547,N_8131,N_8064);
and U9548 (N_9548,N_8624,N_8060);
xnor U9549 (N_9549,N_8153,N_8211);
or U9550 (N_9550,N_8819,N_8535);
and U9551 (N_9551,N_8757,N_8480);
and U9552 (N_9552,N_8818,N_8656);
nand U9553 (N_9553,N_8231,N_8145);
nand U9554 (N_9554,N_8627,N_8284);
nand U9555 (N_9555,N_8643,N_8397);
and U9556 (N_9556,N_8859,N_8259);
xnor U9557 (N_9557,N_8412,N_8158);
nand U9558 (N_9558,N_8790,N_8409);
or U9559 (N_9559,N_8094,N_8774);
xnor U9560 (N_9560,N_8302,N_8118);
nand U9561 (N_9561,N_8430,N_8333);
xnor U9562 (N_9562,N_8526,N_8340);
and U9563 (N_9563,N_8519,N_8704);
nand U9564 (N_9564,N_8818,N_8282);
and U9565 (N_9565,N_8754,N_8186);
and U9566 (N_9566,N_8350,N_8776);
or U9567 (N_9567,N_8629,N_8217);
or U9568 (N_9568,N_8816,N_8618);
nor U9569 (N_9569,N_8103,N_8862);
or U9570 (N_9570,N_8015,N_8031);
and U9571 (N_9571,N_8674,N_8959);
and U9572 (N_9572,N_8381,N_8551);
or U9573 (N_9573,N_8351,N_8770);
or U9574 (N_9574,N_8248,N_8442);
nand U9575 (N_9575,N_8557,N_8228);
and U9576 (N_9576,N_8705,N_8647);
and U9577 (N_9577,N_8082,N_8634);
xnor U9578 (N_9578,N_8114,N_8514);
or U9579 (N_9579,N_8713,N_8333);
nand U9580 (N_9580,N_8066,N_8625);
nor U9581 (N_9581,N_8342,N_8885);
nor U9582 (N_9582,N_8288,N_8762);
and U9583 (N_9583,N_8503,N_8215);
and U9584 (N_9584,N_8048,N_8322);
nand U9585 (N_9585,N_8350,N_8670);
nand U9586 (N_9586,N_8992,N_8255);
and U9587 (N_9587,N_8233,N_8763);
nor U9588 (N_9588,N_8674,N_8664);
nand U9589 (N_9589,N_8586,N_8797);
nand U9590 (N_9590,N_8240,N_8957);
nor U9591 (N_9591,N_8290,N_8289);
xnor U9592 (N_9592,N_8718,N_8921);
and U9593 (N_9593,N_8394,N_8002);
or U9594 (N_9594,N_8705,N_8341);
or U9595 (N_9595,N_8873,N_8047);
nand U9596 (N_9596,N_8660,N_8064);
nand U9597 (N_9597,N_8645,N_8304);
nand U9598 (N_9598,N_8685,N_8673);
nand U9599 (N_9599,N_8368,N_8392);
nor U9600 (N_9600,N_8742,N_8493);
nand U9601 (N_9601,N_8081,N_8699);
or U9602 (N_9602,N_8327,N_8147);
nor U9603 (N_9603,N_8058,N_8011);
or U9604 (N_9604,N_8457,N_8684);
nor U9605 (N_9605,N_8289,N_8293);
or U9606 (N_9606,N_8101,N_8745);
nor U9607 (N_9607,N_8564,N_8968);
nor U9608 (N_9608,N_8379,N_8486);
or U9609 (N_9609,N_8600,N_8560);
and U9610 (N_9610,N_8923,N_8790);
and U9611 (N_9611,N_8371,N_8846);
xnor U9612 (N_9612,N_8583,N_8897);
nand U9613 (N_9613,N_8167,N_8590);
or U9614 (N_9614,N_8274,N_8982);
nand U9615 (N_9615,N_8919,N_8499);
nand U9616 (N_9616,N_8151,N_8993);
or U9617 (N_9617,N_8227,N_8637);
xnor U9618 (N_9618,N_8090,N_8190);
xor U9619 (N_9619,N_8935,N_8511);
xnor U9620 (N_9620,N_8808,N_8582);
or U9621 (N_9621,N_8510,N_8962);
nand U9622 (N_9622,N_8590,N_8465);
and U9623 (N_9623,N_8935,N_8495);
nor U9624 (N_9624,N_8351,N_8613);
or U9625 (N_9625,N_8612,N_8155);
xor U9626 (N_9626,N_8603,N_8325);
nor U9627 (N_9627,N_8405,N_8199);
or U9628 (N_9628,N_8671,N_8897);
or U9629 (N_9629,N_8390,N_8467);
nand U9630 (N_9630,N_8422,N_8355);
nor U9631 (N_9631,N_8773,N_8114);
nand U9632 (N_9632,N_8865,N_8882);
nand U9633 (N_9633,N_8308,N_8283);
nor U9634 (N_9634,N_8851,N_8586);
and U9635 (N_9635,N_8852,N_8999);
xnor U9636 (N_9636,N_8147,N_8606);
and U9637 (N_9637,N_8727,N_8953);
xor U9638 (N_9638,N_8319,N_8043);
and U9639 (N_9639,N_8964,N_8975);
and U9640 (N_9640,N_8619,N_8220);
nand U9641 (N_9641,N_8534,N_8871);
and U9642 (N_9642,N_8903,N_8260);
nor U9643 (N_9643,N_8150,N_8545);
and U9644 (N_9644,N_8811,N_8382);
or U9645 (N_9645,N_8423,N_8733);
or U9646 (N_9646,N_8974,N_8524);
nand U9647 (N_9647,N_8699,N_8449);
and U9648 (N_9648,N_8445,N_8677);
nor U9649 (N_9649,N_8798,N_8979);
nor U9650 (N_9650,N_8022,N_8099);
xnor U9651 (N_9651,N_8248,N_8111);
and U9652 (N_9652,N_8820,N_8196);
and U9653 (N_9653,N_8741,N_8105);
and U9654 (N_9654,N_8625,N_8218);
xor U9655 (N_9655,N_8926,N_8443);
or U9656 (N_9656,N_8879,N_8590);
and U9657 (N_9657,N_8293,N_8379);
or U9658 (N_9658,N_8302,N_8053);
xnor U9659 (N_9659,N_8664,N_8732);
nor U9660 (N_9660,N_8444,N_8113);
and U9661 (N_9661,N_8415,N_8690);
or U9662 (N_9662,N_8942,N_8999);
and U9663 (N_9663,N_8708,N_8069);
nor U9664 (N_9664,N_8009,N_8334);
xnor U9665 (N_9665,N_8426,N_8934);
and U9666 (N_9666,N_8197,N_8538);
nand U9667 (N_9667,N_8558,N_8505);
nor U9668 (N_9668,N_8470,N_8248);
or U9669 (N_9669,N_8668,N_8455);
or U9670 (N_9670,N_8360,N_8824);
xor U9671 (N_9671,N_8882,N_8019);
nand U9672 (N_9672,N_8179,N_8449);
or U9673 (N_9673,N_8387,N_8002);
xnor U9674 (N_9674,N_8904,N_8855);
or U9675 (N_9675,N_8354,N_8056);
xnor U9676 (N_9676,N_8623,N_8404);
xor U9677 (N_9677,N_8282,N_8091);
nand U9678 (N_9678,N_8279,N_8596);
xor U9679 (N_9679,N_8629,N_8234);
nand U9680 (N_9680,N_8105,N_8693);
and U9681 (N_9681,N_8604,N_8347);
and U9682 (N_9682,N_8395,N_8368);
or U9683 (N_9683,N_8546,N_8041);
xor U9684 (N_9684,N_8746,N_8580);
and U9685 (N_9685,N_8750,N_8893);
or U9686 (N_9686,N_8268,N_8767);
xnor U9687 (N_9687,N_8090,N_8781);
xor U9688 (N_9688,N_8125,N_8367);
xor U9689 (N_9689,N_8899,N_8888);
or U9690 (N_9690,N_8551,N_8928);
and U9691 (N_9691,N_8368,N_8230);
xnor U9692 (N_9692,N_8196,N_8512);
and U9693 (N_9693,N_8171,N_8089);
nand U9694 (N_9694,N_8644,N_8892);
nand U9695 (N_9695,N_8215,N_8945);
or U9696 (N_9696,N_8382,N_8226);
and U9697 (N_9697,N_8216,N_8678);
xnor U9698 (N_9698,N_8926,N_8710);
xnor U9699 (N_9699,N_8838,N_8530);
nor U9700 (N_9700,N_8703,N_8815);
xor U9701 (N_9701,N_8062,N_8154);
nand U9702 (N_9702,N_8339,N_8783);
and U9703 (N_9703,N_8799,N_8084);
nand U9704 (N_9704,N_8214,N_8394);
nor U9705 (N_9705,N_8208,N_8913);
or U9706 (N_9706,N_8485,N_8017);
nor U9707 (N_9707,N_8441,N_8446);
nor U9708 (N_9708,N_8262,N_8186);
nor U9709 (N_9709,N_8228,N_8173);
xor U9710 (N_9710,N_8272,N_8412);
nand U9711 (N_9711,N_8662,N_8950);
nor U9712 (N_9712,N_8520,N_8633);
and U9713 (N_9713,N_8837,N_8124);
or U9714 (N_9714,N_8631,N_8202);
and U9715 (N_9715,N_8887,N_8491);
xnor U9716 (N_9716,N_8815,N_8067);
or U9717 (N_9717,N_8827,N_8478);
and U9718 (N_9718,N_8944,N_8139);
xor U9719 (N_9719,N_8334,N_8546);
nor U9720 (N_9720,N_8342,N_8394);
or U9721 (N_9721,N_8060,N_8847);
nor U9722 (N_9722,N_8331,N_8171);
and U9723 (N_9723,N_8640,N_8193);
and U9724 (N_9724,N_8984,N_8615);
nand U9725 (N_9725,N_8966,N_8846);
and U9726 (N_9726,N_8155,N_8531);
nor U9727 (N_9727,N_8312,N_8212);
nor U9728 (N_9728,N_8726,N_8180);
and U9729 (N_9729,N_8795,N_8612);
or U9730 (N_9730,N_8176,N_8867);
or U9731 (N_9731,N_8176,N_8979);
nand U9732 (N_9732,N_8166,N_8388);
nand U9733 (N_9733,N_8924,N_8070);
and U9734 (N_9734,N_8508,N_8158);
xor U9735 (N_9735,N_8657,N_8950);
xor U9736 (N_9736,N_8719,N_8641);
nand U9737 (N_9737,N_8923,N_8383);
xor U9738 (N_9738,N_8802,N_8662);
nand U9739 (N_9739,N_8753,N_8264);
nand U9740 (N_9740,N_8210,N_8393);
nor U9741 (N_9741,N_8725,N_8365);
and U9742 (N_9742,N_8171,N_8571);
nor U9743 (N_9743,N_8234,N_8242);
and U9744 (N_9744,N_8062,N_8026);
nor U9745 (N_9745,N_8255,N_8216);
xnor U9746 (N_9746,N_8896,N_8006);
xor U9747 (N_9747,N_8623,N_8503);
or U9748 (N_9748,N_8885,N_8669);
nand U9749 (N_9749,N_8805,N_8092);
and U9750 (N_9750,N_8236,N_8564);
nand U9751 (N_9751,N_8771,N_8899);
nand U9752 (N_9752,N_8383,N_8637);
nand U9753 (N_9753,N_8233,N_8695);
or U9754 (N_9754,N_8809,N_8351);
or U9755 (N_9755,N_8683,N_8317);
or U9756 (N_9756,N_8446,N_8702);
nor U9757 (N_9757,N_8776,N_8939);
nor U9758 (N_9758,N_8039,N_8487);
nand U9759 (N_9759,N_8413,N_8268);
xor U9760 (N_9760,N_8154,N_8164);
and U9761 (N_9761,N_8710,N_8168);
or U9762 (N_9762,N_8616,N_8281);
or U9763 (N_9763,N_8260,N_8604);
and U9764 (N_9764,N_8492,N_8004);
or U9765 (N_9765,N_8969,N_8226);
xnor U9766 (N_9766,N_8187,N_8590);
and U9767 (N_9767,N_8624,N_8754);
xnor U9768 (N_9768,N_8039,N_8566);
nor U9769 (N_9769,N_8860,N_8271);
xnor U9770 (N_9770,N_8266,N_8708);
nor U9771 (N_9771,N_8490,N_8853);
and U9772 (N_9772,N_8511,N_8419);
and U9773 (N_9773,N_8006,N_8321);
xnor U9774 (N_9774,N_8849,N_8539);
or U9775 (N_9775,N_8619,N_8628);
and U9776 (N_9776,N_8994,N_8220);
nand U9777 (N_9777,N_8678,N_8179);
nand U9778 (N_9778,N_8962,N_8423);
or U9779 (N_9779,N_8859,N_8271);
nor U9780 (N_9780,N_8018,N_8636);
nor U9781 (N_9781,N_8634,N_8501);
or U9782 (N_9782,N_8885,N_8141);
nand U9783 (N_9783,N_8186,N_8725);
nor U9784 (N_9784,N_8683,N_8965);
nor U9785 (N_9785,N_8288,N_8626);
or U9786 (N_9786,N_8071,N_8629);
nand U9787 (N_9787,N_8439,N_8124);
and U9788 (N_9788,N_8555,N_8284);
nand U9789 (N_9789,N_8739,N_8045);
xor U9790 (N_9790,N_8123,N_8954);
nand U9791 (N_9791,N_8040,N_8818);
and U9792 (N_9792,N_8629,N_8379);
nand U9793 (N_9793,N_8800,N_8923);
nor U9794 (N_9794,N_8303,N_8488);
and U9795 (N_9795,N_8780,N_8377);
and U9796 (N_9796,N_8036,N_8127);
nand U9797 (N_9797,N_8807,N_8585);
nor U9798 (N_9798,N_8052,N_8234);
nand U9799 (N_9799,N_8816,N_8142);
or U9800 (N_9800,N_8230,N_8675);
or U9801 (N_9801,N_8047,N_8719);
xor U9802 (N_9802,N_8360,N_8335);
and U9803 (N_9803,N_8763,N_8115);
and U9804 (N_9804,N_8500,N_8454);
or U9805 (N_9805,N_8471,N_8389);
and U9806 (N_9806,N_8481,N_8774);
nand U9807 (N_9807,N_8689,N_8478);
nor U9808 (N_9808,N_8022,N_8460);
xnor U9809 (N_9809,N_8988,N_8673);
or U9810 (N_9810,N_8923,N_8601);
nand U9811 (N_9811,N_8545,N_8290);
xnor U9812 (N_9812,N_8243,N_8734);
xor U9813 (N_9813,N_8108,N_8065);
nand U9814 (N_9814,N_8577,N_8186);
xnor U9815 (N_9815,N_8244,N_8297);
and U9816 (N_9816,N_8033,N_8554);
nor U9817 (N_9817,N_8283,N_8690);
and U9818 (N_9818,N_8519,N_8750);
or U9819 (N_9819,N_8451,N_8766);
and U9820 (N_9820,N_8666,N_8851);
nand U9821 (N_9821,N_8976,N_8364);
and U9822 (N_9822,N_8792,N_8888);
nand U9823 (N_9823,N_8679,N_8459);
nand U9824 (N_9824,N_8124,N_8772);
xnor U9825 (N_9825,N_8950,N_8713);
and U9826 (N_9826,N_8534,N_8366);
nand U9827 (N_9827,N_8052,N_8507);
and U9828 (N_9828,N_8711,N_8257);
nor U9829 (N_9829,N_8669,N_8355);
and U9830 (N_9830,N_8636,N_8729);
and U9831 (N_9831,N_8910,N_8702);
nand U9832 (N_9832,N_8393,N_8208);
nor U9833 (N_9833,N_8664,N_8439);
nand U9834 (N_9834,N_8013,N_8187);
xor U9835 (N_9835,N_8460,N_8632);
nor U9836 (N_9836,N_8253,N_8696);
nor U9837 (N_9837,N_8896,N_8717);
or U9838 (N_9838,N_8434,N_8201);
and U9839 (N_9839,N_8653,N_8201);
xnor U9840 (N_9840,N_8511,N_8995);
nand U9841 (N_9841,N_8669,N_8229);
or U9842 (N_9842,N_8212,N_8477);
nand U9843 (N_9843,N_8274,N_8892);
or U9844 (N_9844,N_8651,N_8964);
nor U9845 (N_9845,N_8677,N_8986);
or U9846 (N_9846,N_8874,N_8646);
and U9847 (N_9847,N_8103,N_8455);
or U9848 (N_9848,N_8579,N_8324);
xnor U9849 (N_9849,N_8451,N_8238);
nor U9850 (N_9850,N_8929,N_8169);
nor U9851 (N_9851,N_8686,N_8413);
nand U9852 (N_9852,N_8093,N_8946);
nand U9853 (N_9853,N_8217,N_8020);
nor U9854 (N_9854,N_8292,N_8698);
nand U9855 (N_9855,N_8715,N_8760);
nand U9856 (N_9856,N_8657,N_8106);
xor U9857 (N_9857,N_8133,N_8804);
xor U9858 (N_9858,N_8293,N_8992);
or U9859 (N_9859,N_8467,N_8684);
xnor U9860 (N_9860,N_8214,N_8461);
nor U9861 (N_9861,N_8501,N_8677);
or U9862 (N_9862,N_8901,N_8084);
xor U9863 (N_9863,N_8444,N_8644);
and U9864 (N_9864,N_8289,N_8201);
nand U9865 (N_9865,N_8779,N_8911);
nor U9866 (N_9866,N_8711,N_8210);
nor U9867 (N_9867,N_8315,N_8080);
xor U9868 (N_9868,N_8115,N_8939);
or U9869 (N_9869,N_8022,N_8016);
and U9870 (N_9870,N_8407,N_8445);
or U9871 (N_9871,N_8062,N_8633);
and U9872 (N_9872,N_8649,N_8582);
or U9873 (N_9873,N_8193,N_8717);
and U9874 (N_9874,N_8088,N_8369);
xnor U9875 (N_9875,N_8193,N_8653);
nor U9876 (N_9876,N_8712,N_8992);
nand U9877 (N_9877,N_8652,N_8598);
or U9878 (N_9878,N_8749,N_8216);
nor U9879 (N_9879,N_8362,N_8813);
or U9880 (N_9880,N_8587,N_8659);
nor U9881 (N_9881,N_8397,N_8637);
and U9882 (N_9882,N_8193,N_8148);
or U9883 (N_9883,N_8996,N_8317);
nor U9884 (N_9884,N_8071,N_8639);
nand U9885 (N_9885,N_8270,N_8832);
xor U9886 (N_9886,N_8002,N_8599);
or U9887 (N_9887,N_8599,N_8451);
nor U9888 (N_9888,N_8422,N_8152);
xor U9889 (N_9889,N_8419,N_8182);
and U9890 (N_9890,N_8905,N_8416);
or U9891 (N_9891,N_8712,N_8698);
nand U9892 (N_9892,N_8526,N_8513);
nand U9893 (N_9893,N_8148,N_8492);
nand U9894 (N_9894,N_8522,N_8168);
and U9895 (N_9895,N_8015,N_8908);
or U9896 (N_9896,N_8634,N_8585);
nand U9897 (N_9897,N_8011,N_8204);
nand U9898 (N_9898,N_8473,N_8979);
nor U9899 (N_9899,N_8824,N_8886);
and U9900 (N_9900,N_8031,N_8330);
nand U9901 (N_9901,N_8173,N_8184);
or U9902 (N_9902,N_8352,N_8553);
nor U9903 (N_9903,N_8316,N_8986);
and U9904 (N_9904,N_8681,N_8705);
or U9905 (N_9905,N_8524,N_8518);
nor U9906 (N_9906,N_8289,N_8114);
and U9907 (N_9907,N_8464,N_8088);
and U9908 (N_9908,N_8454,N_8090);
and U9909 (N_9909,N_8699,N_8877);
nor U9910 (N_9910,N_8629,N_8850);
nor U9911 (N_9911,N_8511,N_8806);
and U9912 (N_9912,N_8041,N_8774);
and U9913 (N_9913,N_8064,N_8220);
xnor U9914 (N_9914,N_8680,N_8115);
xor U9915 (N_9915,N_8109,N_8604);
or U9916 (N_9916,N_8047,N_8071);
nor U9917 (N_9917,N_8264,N_8341);
nand U9918 (N_9918,N_8734,N_8611);
nand U9919 (N_9919,N_8578,N_8347);
xor U9920 (N_9920,N_8914,N_8581);
and U9921 (N_9921,N_8571,N_8678);
nand U9922 (N_9922,N_8742,N_8804);
or U9923 (N_9923,N_8624,N_8704);
or U9924 (N_9924,N_8750,N_8259);
nand U9925 (N_9925,N_8908,N_8622);
xor U9926 (N_9926,N_8196,N_8935);
and U9927 (N_9927,N_8407,N_8373);
or U9928 (N_9928,N_8866,N_8453);
nand U9929 (N_9929,N_8430,N_8432);
and U9930 (N_9930,N_8455,N_8269);
or U9931 (N_9931,N_8820,N_8589);
or U9932 (N_9932,N_8152,N_8707);
or U9933 (N_9933,N_8626,N_8121);
and U9934 (N_9934,N_8695,N_8073);
xor U9935 (N_9935,N_8675,N_8212);
or U9936 (N_9936,N_8155,N_8800);
xor U9937 (N_9937,N_8304,N_8049);
or U9938 (N_9938,N_8532,N_8196);
nand U9939 (N_9939,N_8621,N_8871);
or U9940 (N_9940,N_8374,N_8666);
xor U9941 (N_9941,N_8045,N_8368);
nor U9942 (N_9942,N_8934,N_8021);
or U9943 (N_9943,N_8567,N_8254);
and U9944 (N_9944,N_8947,N_8312);
nor U9945 (N_9945,N_8940,N_8135);
or U9946 (N_9946,N_8878,N_8450);
and U9947 (N_9947,N_8131,N_8123);
and U9948 (N_9948,N_8324,N_8155);
nand U9949 (N_9949,N_8839,N_8895);
or U9950 (N_9950,N_8667,N_8257);
or U9951 (N_9951,N_8198,N_8403);
and U9952 (N_9952,N_8711,N_8536);
nand U9953 (N_9953,N_8674,N_8461);
nor U9954 (N_9954,N_8992,N_8109);
xnor U9955 (N_9955,N_8951,N_8458);
nor U9956 (N_9956,N_8894,N_8232);
xnor U9957 (N_9957,N_8197,N_8296);
xor U9958 (N_9958,N_8704,N_8840);
nand U9959 (N_9959,N_8567,N_8252);
xnor U9960 (N_9960,N_8366,N_8313);
and U9961 (N_9961,N_8100,N_8843);
nand U9962 (N_9962,N_8654,N_8592);
or U9963 (N_9963,N_8104,N_8428);
and U9964 (N_9964,N_8609,N_8681);
and U9965 (N_9965,N_8871,N_8474);
and U9966 (N_9966,N_8547,N_8926);
xnor U9967 (N_9967,N_8082,N_8281);
or U9968 (N_9968,N_8444,N_8819);
or U9969 (N_9969,N_8994,N_8340);
nor U9970 (N_9970,N_8872,N_8572);
nor U9971 (N_9971,N_8798,N_8082);
and U9972 (N_9972,N_8524,N_8713);
nor U9973 (N_9973,N_8233,N_8642);
nor U9974 (N_9974,N_8087,N_8644);
or U9975 (N_9975,N_8902,N_8455);
or U9976 (N_9976,N_8297,N_8934);
nand U9977 (N_9977,N_8086,N_8970);
or U9978 (N_9978,N_8804,N_8598);
nand U9979 (N_9979,N_8558,N_8894);
nor U9980 (N_9980,N_8337,N_8706);
nand U9981 (N_9981,N_8728,N_8666);
and U9982 (N_9982,N_8475,N_8323);
xnor U9983 (N_9983,N_8642,N_8124);
xnor U9984 (N_9984,N_8359,N_8941);
or U9985 (N_9985,N_8456,N_8082);
nor U9986 (N_9986,N_8952,N_8680);
nand U9987 (N_9987,N_8275,N_8166);
or U9988 (N_9988,N_8650,N_8063);
and U9989 (N_9989,N_8846,N_8209);
nand U9990 (N_9990,N_8040,N_8948);
and U9991 (N_9991,N_8223,N_8290);
nand U9992 (N_9992,N_8381,N_8048);
nor U9993 (N_9993,N_8921,N_8168);
xnor U9994 (N_9994,N_8381,N_8545);
nand U9995 (N_9995,N_8730,N_8806);
xor U9996 (N_9996,N_8540,N_8051);
or U9997 (N_9997,N_8553,N_8700);
and U9998 (N_9998,N_8758,N_8539);
and U9999 (N_9999,N_8497,N_8598);
xnor UO_0 (O_0,N_9585,N_9478);
or UO_1 (O_1,N_9964,N_9457);
or UO_2 (O_2,N_9292,N_9367);
nand UO_3 (O_3,N_9064,N_9032);
nand UO_4 (O_4,N_9284,N_9142);
nand UO_5 (O_5,N_9613,N_9118);
xor UO_6 (O_6,N_9098,N_9130);
or UO_7 (O_7,N_9249,N_9742);
and UO_8 (O_8,N_9406,N_9180);
and UO_9 (O_9,N_9340,N_9391);
nand UO_10 (O_10,N_9820,N_9814);
or UO_11 (O_11,N_9153,N_9554);
and UO_12 (O_12,N_9815,N_9945);
nor UO_13 (O_13,N_9464,N_9777);
and UO_14 (O_14,N_9233,N_9159);
and UO_15 (O_15,N_9986,N_9677);
nor UO_16 (O_16,N_9879,N_9960);
and UO_17 (O_17,N_9418,N_9397);
or UO_18 (O_18,N_9358,N_9845);
and UO_19 (O_19,N_9607,N_9876);
or UO_20 (O_20,N_9447,N_9303);
nand UO_21 (O_21,N_9229,N_9014);
and UO_22 (O_22,N_9254,N_9881);
xnor UO_23 (O_23,N_9663,N_9051);
nor UO_24 (O_24,N_9054,N_9207);
or UO_25 (O_25,N_9047,N_9530);
and UO_26 (O_26,N_9381,N_9966);
nand UO_27 (O_27,N_9730,N_9536);
or UO_28 (O_28,N_9754,N_9955);
or UO_29 (O_29,N_9701,N_9917);
and UO_30 (O_30,N_9366,N_9022);
xor UO_31 (O_31,N_9011,N_9204);
and UO_32 (O_32,N_9526,N_9949);
nand UO_33 (O_33,N_9532,N_9557);
xor UO_34 (O_34,N_9637,N_9185);
xor UO_35 (O_35,N_9178,N_9334);
nor UO_36 (O_36,N_9594,N_9856);
or UO_37 (O_37,N_9596,N_9188);
xnor UO_38 (O_38,N_9831,N_9546);
xnor UO_39 (O_39,N_9737,N_9595);
xor UO_40 (O_40,N_9529,N_9643);
nand UO_41 (O_41,N_9039,N_9860);
nand UO_42 (O_42,N_9665,N_9518);
nand UO_43 (O_43,N_9510,N_9893);
nor UO_44 (O_44,N_9283,N_9538);
and UO_45 (O_45,N_9902,N_9310);
or UO_46 (O_46,N_9693,N_9706);
or UO_47 (O_47,N_9985,N_9555);
nor UO_48 (O_48,N_9650,N_9989);
and UO_49 (O_49,N_9355,N_9658);
nand UO_50 (O_50,N_9921,N_9847);
xnor UO_51 (O_51,N_9439,N_9980);
xnor UO_52 (O_52,N_9275,N_9928);
xor UO_53 (O_53,N_9041,N_9822);
and UO_54 (O_54,N_9516,N_9450);
or UO_55 (O_55,N_9676,N_9660);
nand UO_56 (O_56,N_9190,N_9357);
nor UO_57 (O_57,N_9774,N_9463);
and UO_58 (O_58,N_9056,N_9927);
xnor UO_59 (O_59,N_9487,N_9779);
or UO_60 (O_60,N_9436,N_9217);
or UO_61 (O_61,N_9316,N_9992);
or UO_62 (O_62,N_9537,N_9084);
and UO_63 (O_63,N_9887,N_9168);
or UO_64 (O_64,N_9388,N_9498);
and UO_65 (O_65,N_9884,N_9946);
nand UO_66 (O_66,N_9030,N_9135);
nor UO_67 (O_67,N_9053,N_9776);
and UO_68 (O_68,N_9709,N_9323);
and UO_69 (O_69,N_9788,N_9052);
nor UO_70 (O_70,N_9850,N_9019);
and UO_71 (O_71,N_9844,N_9352);
and UO_72 (O_72,N_9095,N_9790);
xnor UO_73 (O_73,N_9187,N_9266);
and UO_74 (O_74,N_9553,N_9308);
xnor UO_75 (O_75,N_9981,N_9453);
xor UO_76 (O_76,N_9026,N_9751);
or UO_77 (O_77,N_9348,N_9760);
and UO_78 (O_78,N_9091,N_9008);
nor UO_79 (O_79,N_9525,N_9664);
nand UO_80 (O_80,N_9561,N_9396);
or UO_81 (O_81,N_9200,N_9382);
xnor UO_82 (O_82,N_9191,N_9655);
or UO_83 (O_83,N_9269,N_9503);
nor UO_84 (O_84,N_9891,N_9816);
and UO_85 (O_85,N_9982,N_9652);
nand UO_86 (O_86,N_9489,N_9152);
or UO_87 (O_87,N_9624,N_9231);
nor UO_88 (O_88,N_9714,N_9076);
xor UO_89 (O_89,N_9507,N_9282);
nor UO_90 (O_90,N_9990,N_9398);
nor UO_91 (O_91,N_9719,N_9160);
xnor UO_92 (O_92,N_9248,N_9186);
xnor UO_93 (O_93,N_9110,N_9771);
and UO_94 (O_94,N_9710,N_9281);
nand UO_95 (O_95,N_9659,N_9021);
nor UO_96 (O_96,N_9865,N_9297);
xor UO_97 (O_97,N_9608,N_9247);
xor UO_98 (O_98,N_9048,N_9695);
and UO_99 (O_99,N_9027,N_9471);
and UO_100 (O_100,N_9020,N_9127);
and UO_101 (O_101,N_9101,N_9519);
xnor UO_102 (O_102,N_9818,N_9792);
and UO_103 (O_103,N_9924,N_9544);
nor UO_104 (O_104,N_9100,N_9678);
xnor UO_105 (O_105,N_9642,N_9549);
xor UO_106 (O_106,N_9430,N_9956);
xor UO_107 (O_107,N_9023,N_9745);
xor UO_108 (O_108,N_9307,N_9370);
and UO_109 (O_109,N_9647,N_9145);
nand UO_110 (O_110,N_9550,N_9028);
and UO_111 (O_111,N_9469,N_9531);
nor UO_112 (O_112,N_9733,N_9113);
xor UO_113 (O_113,N_9081,N_9885);
and UO_114 (O_114,N_9798,N_9267);
xor UO_115 (O_115,N_9409,N_9134);
and UO_116 (O_116,N_9983,N_9506);
or UO_117 (O_117,N_9309,N_9727);
nand UO_118 (O_118,N_9963,N_9304);
nor UO_119 (O_119,N_9944,N_9648);
nand UO_120 (O_120,N_9897,N_9910);
or UO_121 (O_121,N_9832,N_9606);
xnor UO_122 (O_122,N_9230,N_9038);
nor UO_123 (O_123,N_9387,N_9636);
xor UO_124 (O_124,N_9634,N_9684);
nand UO_125 (O_125,N_9619,N_9795);
xnor UO_126 (O_126,N_9468,N_9029);
nand UO_127 (O_127,N_9424,N_9566);
nor UO_128 (O_128,N_9791,N_9003);
nand UO_129 (O_129,N_9728,N_9286);
or UO_130 (O_130,N_9768,N_9006);
or UO_131 (O_131,N_9569,N_9895);
xor UO_132 (O_132,N_9128,N_9973);
nand UO_133 (O_133,N_9103,N_9732);
nor UO_134 (O_134,N_9122,N_9037);
or UO_135 (O_135,N_9163,N_9681);
nor UO_136 (O_136,N_9589,N_9155);
nor UO_137 (O_137,N_9700,N_9718);
or UO_138 (O_138,N_9414,N_9962);
xor UO_139 (O_139,N_9456,N_9562);
nand UO_140 (O_140,N_9074,N_9939);
or UO_141 (O_141,N_9942,N_9215);
xnor UO_142 (O_142,N_9715,N_9344);
nand UO_143 (O_143,N_9720,N_9036);
or UO_144 (O_144,N_9654,N_9328);
or UO_145 (O_145,N_9901,N_9558);
nor UO_146 (O_146,N_9431,N_9579);
nand UO_147 (O_147,N_9488,N_9184);
nand UO_148 (O_148,N_9116,N_9260);
nor UO_149 (O_149,N_9043,N_9123);
nor UO_150 (O_150,N_9067,N_9094);
xor UO_151 (O_151,N_9373,N_9392);
and UO_152 (O_152,N_9143,N_9697);
xnor UO_153 (O_153,N_9961,N_9476);
or UO_154 (O_154,N_9285,N_9057);
or UO_155 (O_155,N_9671,N_9623);
and UO_156 (O_156,N_9482,N_9769);
or UO_157 (O_157,N_9126,N_9222);
and UO_158 (O_158,N_9408,N_9954);
nor UO_159 (O_159,N_9124,N_9073);
or UO_160 (O_160,N_9375,N_9333);
or UO_161 (O_161,N_9686,N_9915);
or UO_162 (O_162,N_9616,N_9545);
nor UO_163 (O_163,N_9683,N_9315);
nor UO_164 (O_164,N_9484,N_9878);
nor UO_165 (O_165,N_9661,N_9138);
nand UO_166 (O_166,N_9179,N_9739);
nor UO_167 (O_167,N_9383,N_9242);
nor UO_168 (O_168,N_9801,N_9426);
and UO_169 (O_169,N_9459,N_9514);
nand UO_170 (O_170,N_9347,N_9889);
xnor UO_171 (O_171,N_9725,N_9451);
nor UO_172 (O_172,N_9106,N_9206);
nor UO_173 (O_173,N_9587,N_9762);
or UO_174 (O_174,N_9552,N_9610);
xnor UO_175 (O_175,N_9108,N_9428);
xor UO_176 (O_176,N_9353,N_9794);
nor UO_177 (O_177,N_9764,N_9121);
nand UO_178 (O_178,N_9778,N_9724);
or UO_179 (O_179,N_9688,N_9953);
nand UO_180 (O_180,N_9827,N_9287);
xnor UO_181 (O_181,N_9626,N_9470);
and UO_182 (O_182,N_9970,N_9258);
and UO_183 (O_183,N_9322,N_9735);
or UO_184 (O_184,N_9541,N_9240);
nand UO_185 (O_185,N_9598,N_9314);
or UO_186 (O_186,N_9120,N_9148);
and UO_187 (O_187,N_9189,N_9062);
and UO_188 (O_188,N_9882,N_9176);
and UO_189 (O_189,N_9063,N_9279);
nand UO_190 (O_190,N_9363,N_9079);
xnor UO_191 (O_191,N_9351,N_9505);
or UO_192 (O_192,N_9389,N_9851);
and UO_193 (O_193,N_9289,N_9004);
nand UO_194 (O_194,N_9295,N_9293);
nor UO_195 (O_195,N_9477,N_9035);
or UO_196 (O_196,N_9244,N_9691);
nand UO_197 (O_197,N_9040,N_9016);
and UO_198 (O_198,N_9548,N_9994);
or UO_199 (O_199,N_9326,N_9903);
nand UO_200 (O_200,N_9114,N_9046);
xor UO_201 (O_201,N_9227,N_9574);
nor UO_202 (O_202,N_9501,N_9429);
or UO_203 (O_203,N_9717,N_9861);
or UO_204 (O_204,N_9508,N_9354);
or UO_205 (O_205,N_9919,N_9490);
xnor UO_206 (O_206,N_9385,N_9926);
or UO_207 (O_207,N_9854,N_9483);
xnor UO_208 (O_208,N_9540,N_9789);
xor UO_209 (O_209,N_9465,N_9369);
xor UO_210 (O_210,N_9165,N_9628);
xnor UO_211 (O_211,N_9433,N_9455);
or UO_212 (O_212,N_9937,N_9183);
nor UO_213 (O_213,N_9149,N_9330);
and UO_214 (O_214,N_9515,N_9797);
or UO_215 (O_215,N_9810,N_9427);
and UO_216 (O_216,N_9611,N_9298);
xnor UO_217 (O_217,N_9495,N_9662);
or UO_218 (O_218,N_9524,N_9723);
and UO_219 (O_219,N_9205,N_9072);
nor UO_220 (O_220,N_9133,N_9086);
and UO_221 (O_221,N_9338,N_9259);
nand UO_222 (O_222,N_9971,N_9068);
or UO_223 (O_223,N_9950,N_9241);
nor UO_224 (O_224,N_9336,N_9007);
xnor UO_225 (O_225,N_9571,N_9911);
nand UO_226 (O_226,N_9609,N_9687);
or UO_227 (O_227,N_9443,N_9807);
or UO_228 (O_228,N_9274,N_9224);
nand UO_229 (O_229,N_9957,N_9842);
nor UO_230 (O_230,N_9460,N_9422);
nor UO_231 (O_231,N_9033,N_9726);
nor UO_232 (O_232,N_9087,N_9932);
nand UO_233 (O_233,N_9226,N_9836);
nor UO_234 (O_234,N_9834,N_9045);
nand UO_235 (O_235,N_9781,N_9622);
nor UO_236 (O_236,N_9502,N_9934);
xnor UO_237 (O_237,N_9864,N_9584);
and UO_238 (O_238,N_9920,N_9632);
and UO_239 (O_239,N_9232,N_9402);
xnor UO_240 (O_240,N_9306,N_9829);
xnor UO_241 (O_241,N_9682,N_9320);
nor UO_242 (O_242,N_9245,N_9150);
or UO_243 (O_243,N_9166,N_9952);
and UO_244 (O_244,N_9401,N_9042);
xnor UO_245 (O_245,N_9621,N_9689);
nor UO_246 (O_246,N_9547,N_9784);
and UO_247 (O_247,N_9657,N_9640);
or UO_248 (O_248,N_9025,N_9753);
xor UO_249 (O_249,N_9452,N_9496);
and UO_250 (O_250,N_9638,N_9757);
and UO_251 (O_251,N_9883,N_9602);
xnor UO_252 (O_252,N_9243,N_9093);
nor UO_253 (O_253,N_9194,N_9835);
nor UO_254 (O_254,N_9192,N_9786);
or UO_255 (O_255,N_9914,N_9238);
xnor UO_256 (O_256,N_9830,N_9500);
nand UO_257 (O_257,N_9603,N_9362);
and UO_258 (O_258,N_9480,N_9823);
nand UO_259 (O_259,N_9301,N_9995);
nand UO_260 (O_260,N_9372,N_9617);
nor UO_261 (O_261,N_9291,N_9975);
and UO_262 (O_262,N_9273,N_9132);
and UO_263 (O_263,N_9290,N_9565);
and UO_264 (O_264,N_9112,N_9704);
nand UO_265 (O_265,N_9649,N_9533);
and UO_266 (O_266,N_9886,N_9441);
nand UO_267 (O_267,N_9808,N_9800);
xor UO_268 (O_268,N_9085,N_9568);
or UO_269 (O_269,N_9872,N_9393);
xnor UO_270 (O_270,N_9486,N_9690);
nor UO_271 (O_271,N_9858,N_9253);
xnor UO_272 (O_272,N_9846,N_9935);
or UO_273 (O_273,N_9862,N_9350);
nand UO_274 (O_274,N_9341,N_9237);
or UO_275 (O_275,N_9641,N_9627);
or UO_276 (O_276,N_9839,N_9824);
nor UO_277 (O_277,N_9923,N_9219);
nand UO_278 (O_278,N_9305,N_9843);
nand UO_279 (O_279,N_9175,N_9984);
or UO_280 (O_280,N_9473,N_9412);
nor UO_281 (O_281,N_9193,N_9013);
and UO_282 (O_282,N_9821,N_9413);
and UO_283 (O_283,N_9890,N_9109);
xor UO_284 (O_284,N_9645,N_9535);
and UO_285 (O_285,N_9346,N_9070);
or UO_286 (O_286,N_9813,N_9894);
xnor UO_287 (O_287,N_9685,N_9674);
or UO_288 (O_288,N_9875,N_9140);
and UO_289 (O_289,N_9395,N_9913);
and UO_290 (O_290,N_9772,N_9947);
nor UO_291 (O_291,N_9218,N_9467);
or UO_292 (O_292,N_9672,N_9157);
nor UO_293 (O_293,N_9511,N_9692);
and UO_294 (O_294,N_9870,N_9716);
xor UO_295 (O_295,N_9379,N_9411);
xnor UO_296 (O_296,N_9221,N_9837);
and UO_297 (O_297,N_9899,N_9630);
xor UO_298 (O_298,N_9588,N_9146);
nor UO_299 (O_299,N_9104,N_9485);
nor UO_300 (O_300,N_9793,N_9520);
or UO_301 (O_301,N_9527,N_9590);
nand UO_302 (O_302,N_9089,N_9852);
nand UO_303 (O_303,N_9578,N_9252);
nor UO_304 (O_304,N_9107,N_9102);
or UO_305 (O_305,N_9817,N_9223);
nor UO_306 (O_306,N_9580,N_9376);
nand UO_307 (O_307,N_9147,N_9492);
nor UO_308 (O_308,N_9105,N_9169);
nand UO_309 (O_309,N_9417,N_9208);
and UO_310 (O_310,N_9698,N_9472);
nor UO_311 (O_311,N_9805,N_9906);
nor UO_312 (O_312,N_9335,N_9542);
xnor UO_313 (O_313,N_9201,N_9216);
nor UO_314 (O_314,N_9088,N_9421);
or UO_315 (O_315,N_9318,N_9246);
nand UO_316 (O_316,N_9078,N_9479);
and UO_317 (O_317,N_9390,N_9877);
or UO_318 (O_318,N_9448,N_9171);
xnor UO_319 (O_319,N_9129,N_9577);
xnor UO_320 (O_320,N_9423,N_9907);
or UO_321 (O_321,N_9410,N_9667);
nor UO_322 (O_322,N_9857,N_9024);
and UO_323 (O_323,N_9696,N_9804);
and UO_324 (O_324,N_9071,N_9010);
or UO_325 (O_325,N_9629,N_9898);
and UO_326 (O_326,N_9212,N_9528);
nand UO_327 (O_327,N_9722,N_9400);
nor UO_328 (O_328,N_9420,N_9059);
xor UO_329 (O_329,N_9251,N_9614);
nor UO_330 (O_330,N_9517,N_9405);
xnor UO_331 (O_331,N_9838,N_9466);
xnor UO_332 (O_332,N_9618,N_9702);
or UO_333 (O_333,N_9151,N_9278);
or UO_334 (O_334,N_9065,N_9741);
and UO_335 (O_335,N_9270,N_9077);
nand UO_336 (O_336,N_9356,N_9058);
nor UO_337 (O_337,N_9239,N_9263);
xnor UO_338 (O_338,N_9438,N_9250);
or UO_339 (O_339,N_9181,N_9977);
or UO_340 (O_340,N_9987,N_9563);
xnor UO_341 (O_341,N_9539,N_9705);
and UO_342 (O_342,N_9359,N_9481);
nor UO_343 (O_343,N_9137,N_9203);
or UO_344 (O_344,N_9866,N_9600);
xnor UO_345 (O_345,N_9440,N_9512);
xnor UO_346 (O_346,N_9434,N_9271);
nor UO_347 (O_347,N_9329,N_9656);
xnor UO_348 (O_348,N_9900,N_9294);
or UO_349 (O_349,N_9633,N_9841);
or UO_350 (O_350,N_9435,N_9491);
xnor UO_351 (O_351,N_9651,N_9930);
nor UO_352 (O_352,N_9001,N_9680);
and UO_353 (O_353,N_9969,N_9182);
nor UO_354 (O_354,N_9748,N_9668);
nor UO_355 (O_355,N_9556,N_9236);
xor UO_356 (O_356,N_9755,N_9597);
nor UO_357 (O_357,N_9097,N_9625);
xor UO_358 (O_358,N_9277,N_9604);
nor UO_359 (O_359,N_9750,N_9965);
nand UO_360 (O_360,N_9075,N_9871);
xnor UO_361 (O_361,N_9276,N_9374);
nand UO_362 (O_362,N_9378,N_9069);
nor UO_363 (O_363,N_9922,N_9111);
and UO_364 (O_364,N_9812,N_9721);
and UO_365 (O_365,N_9738,N_9752);
nand UO_366 (O_366,N_9765,N_9999);
nand UO_367 (O_367,N_9474,N_9261);
nor UO_368 (O_368,N_9031,N_9734);
and UO_369 (O_369,N_9386,N_9321);
or UO_370 (O_370,N_9080,N_9703);
nor UO_371 (O_371,N_9908,N_9740);
or UO_372 (O_372,N_9343,N_9324);
and UO_373 (O_373,N_9896,N_9131);
and UO_374 (O_374,N_9399,N_9445);
and UO_375 (O_375,N_9669,N_9044);
xnor UO_376 (O_376,N_9736,N_9912);
nor UO_377 (O_377,N_9174,N_9666);
and UO_378 (O_378,N_9234,N_9806);
and UO_379 (O_379,N_9712,N_9228);
nor UO_380 (O_380,N_9012,N_9675);
or UO_381 (O_381,N_9639,N_9312);
nand UO_382 (O_382,N_9933,N_9437);
and UO_383 (O_383,N_9302,N_9005);
nor UO_384 (O_384,N_9017,N_9235);
and UO_385 (O_385,N_9567,N_9199);
nand UO_386 (O_386,N_9782,N_9050);
and UO_387 (O_387,N_9198,N_9117);
xor UO_388 (O_388,N_9635,N_9559);
and UO_389 (O_389,N_9317,N_9493);
and UO_390 (O_390,N_9670,N_9202);
nand UO_391 (O_391,N_9853,N_9331);
xor UO_392 (O_392,N_9313,N_9729);
xnor UO_393 (O_393,N_9268,N_9197);
or UO_394 (O_394,N_9711,N_9593);
and UO_395 (O_395,N_9384,N_9494);
and UO_396 (O_396,N_9599,N_9136);
xor UO_397 (O_397,N_9744,N_9646);
nand UO_398 (O_398,N_9694,N_9766);
and UO_399 (O_399,N_9407,N_9958);
and UO_400 (O_400,N_9560,N_9775);
nor UO_401 (O_401,N_9015,N_9060);
and UO_402 (O_402,N_9158,N_9360);
and UO_403 (O_403,N_9581,N_9377);
and UO_404 (O_404,N_9849,N_9394);
nor UO_405 (O_405,N_9523,N_9264);
or UO_406 (O_406,N_9009,N_9257);
nand UO_407 (O_407,N_9936,N_9941);
xor UO_408 (O_408,N_9615,N_9918);
nand UO_409 (O_409,N_9773,N_9991);
nand UO_410 (O_410,N_9840,N_9172);
nor UO_411 (O_411,N_9213,N_9499);
nand UO_412 (O_412,N_9167,N_9763);
and UO_413 (O_413,N_9415,N_9534);
and UO_414 (O_414,N_9096,N_9002);
or UO_415 (O_415,N_9564,N_9214);
or UO_416 (O_416,N_9967,N_9458);
xnor UO_417 (O_417,N_9968,N_9880);
and UO_418 (O_418,N_9997,N_9925);
nor UO_419 (O_419,N_9707,N_9868);
nor UO_420 (O_420,N_9272,N_9988);
or UO_421 (O_421,N_9938,N_9731);
xnor UO_422 (O_422,N_9948,N_9713);
xor UO_423 (O_423,N_9959,N_9888);
xnor UO_424 (O_424,N_9342,N_9115);
nand UO_425 (O_425,N_9299,N_9170);
xnor UO_426 (O_426,N_9905,N_9404);
nor UO_427 (O_427,N_9653,N_9591);
xnor UO_428 (O_428,N_9161,N_9859);
nor UO_429 (O_429,N_9867,N_9572);
or UO_430 (O_430,N_9758,N_9280);
nand UO_431 (O_431,N_9586,N_9220);
and UO_432 (O_432,N_9940,N_9177);
or UO_433 (O_433,N_9543,N_9000);
nand UO_434 (O_434,N_9475,N_9432);
nor UO_435 (O_435,N_9825,N_9454);
nor UO_436 (O_436,N_9673,N_9582);
and UO_437 (O_437,N_9743,N_9034);
and UO_438 (O_438,N_9605,N_9265);
and UO_439 (O_439,N_9380,N_9979);
or UO_440 (O_440,N_9371,N_9442);
or UO_441 (O_441,N_9592,N_9497);
xor UO_442 (O_442,N_9262,N_9300);
nor UO_443 (O_443,N_9049,N_9869);
or UO_444 (O_444,N_9972,N_9337);
nor UO_445 (O_445,N_9679,N_9996);
nand UO_446 (O_446,N_9349,N_9092);
nand UO_447 (O_447,N_9787,N_9747);
nand UO_448 (O_448,N_9819,N_9978);
xor UO_449 (O_449,N_9620,N_9916);
or UO_450 (O_450,N_9931,N_9570);
xor UO_451 (O_451,N_9327,N_9099);
and UO_452 (O_452,N_9785,N_9892);
nand UO_453 (O_453,N_9770,N_9210);
and UO_454 (O_454,N_9018,N_9461);
or UO_455 (O_455,N_9909,N_9576);
xor UO_456 (O_456,N_9416,N_9425);
and UO_457 (O_457,N_9365,N_9332);
or UO_458 (O_458,N_9904,N_9976);
and UO_459 (O_459,N_9783,N_9767);
nand UO_460 (O_460,N_9513,N_9256);
and UO_461 (O_461,N_9855,N_9951);
or UO_462 (O_462,N_9066,N_9125);
nor UO_463 (O_463,N_9631,N_9288);
xor UO_464 (O_464,N_9255,N_9446);
and UO_465 (O_465,N_9863,N_9826);
and UO_466 (O_466,N_9154,N_9296);
nand UO_467 (O_467,N_9090,N_9345);
xor UO_468 (O_468,N_9708,N_9943);
xnor UO_469 (O_469,N_9583,N_9055);
and UO_470 (O_470,N_9156,N_9211);
nand UO_471 (O_471,N_9522,N_9874);
or UO_472 (O_472,N_9575,N_9796);
nand UO_473 (O_473,N_9164,N_9196);
or UO_474 (O_474,N_9462,N_9811);
or UO_475 (O_475,N_9509,N_9195);
nor UO_476 (O_476,N_9551,N_9780);
xnor UO_477 (O_477,N_9974,N_9612);
or UO_478 (O_478,N_9803,N_9756);
xor UO_479 (O_479,N_9833,N_9083);
or UO_480 (O_480,N_9449,N_9141);
and UO_481 (O_481,N_9809,N_9802);
or UO_482 (O_482,N_9368,N_9311);
nor UO_483 (O_483,N_9119,N_9873);
nor UO_484 (O_484,N_9828,N_9746);
and UO_485 (O_485,N_9061,N_9521);
xor UO_486 (O_486,N_9209,N_9082);
or UO_487 (O_487,N_9325,N_9225);
nand UO_488 (O_488,N_9848,N_9361);
or UO_489 (O_489,N_9139,N_9403);
nor UO_490 (O_490,N_9419,N_9929);
xor UO_491 (O_491,N_9162,N_9761);
nor UO_492 (O_492,N_9601,N_9319);
nand UO_493 (O_493,N_9699,N_9339);
or UO_494 (O_494,N_9749,N_9799);
and UO_495 (O_495,N_9759,N_9144);
or UO_496 (O_496,N_9573,N_9173);
nand UO_497 (O_497,N_9993,N_9444);
nand UO_498 (O_498,N_9364,N_9504);
nor UO_499 (O_499,N_9998,N_9644);
nor UO_500 (O_500,N_9692,N_9075);
or UO_501 (O_501,N_9101,N_9643);
and UO_502 (O_502,N_9204,N_9546);
and UO_503 (O_503,N_9472,N_9566);
and UO_504 (O_504,N_9976,N_9930);
nand UO_505 (O_505,N_9093,N_9663);
or UO_506 (O_506,N_9857,N_9886);
nand UO_507 (O_507,N_9248,N_9986);
nand UO_508 (O_508,N_9045,N_9643);
and UO_509 (O_509,N_9169,N_9264);
nor UO_510 (O_510,N_9283,N_9035);
nand UO_511 (O_511,N_9670,N_9442);
or UO_512 (O_512,N_9840,N_9429);
and UO_513 (O_513,N_9999,N_9853);
or UO_514 (O_514,N_9909,N_9194);
nor UO_515 (O_515,N_9316,N_9840);
xnor UO_516 (O_516,N_9120,N_9088);
or UO_517 (O_517,N_9036,N_9290);
nand UO_518 (O_518,N_9806,N_9249);
or UO_519 (O_519,N_9978,N_9672);
or UO_520 (O_520,N_9725,N_9965);
nor UO_521 (O_521,N_9019,N_9790);
nor UO_522 (O_522,N_9413,N_9282);
xor UO_523 (O_523,N_9022,N_9563);
xnor UO_524 (O_524,N_9193,N_9406);
nor UO_525 (O_525,N_9241,N_9031);
xnor UO_526 (O_526,N_9344,N_9769);
nor UO_527 (O_527,N_9745,N_9952);
or UO_528 (O_528,N_9164,N_9187);
nand UO_529 (O_529,N_9638,N_9810);
xnor UO_530 (O_530,N_9903,N_9336);
xnor UO_531 (O_531,N_9852,N_9585);
xnor UO_532 (O_532,N_9124,N_9585);
nor UO_533 (O_533,N_9025,N_9683);
nand UO_534 (O_534,N_9577,N_9045);
nand UO_535 (O_535,N_9186,N_9808);
xor UO_536 (O_536,N_9646,N_9999);
or UO_537 (O_537,N_9653,N_9394);
and UO_538 (O_538,N_9269,N_9216);
xnor UO_539 (O_539,N_9806,N_9332);
xor UO_540 (O_540,N_9069,N_9962);
nand UO_541 (O_541,N_9042,N_9674);
and UO_542 (O_542,N_9310,N_9292);
and UO_543 (O_543,N_9479,N_9110);
or UO_544 (O_544,N_9594,N_9246);
xnor UO_545 (O_545,N_9781,N_9962);
xnor UO_546 (O_546,N_9597,N_9179);
xor UO_547 (O_547,N_9472,N_9492);
nor UO_548 (O_548,N_9066,N_9504);
or UO_549 (O_549,N_9445,N_9015);
nor UO_550 (O_550,N_9523,N_9191);
or UO_551 (O_551,N_9664,N_9150);
nor UO_552 (O_552,N_9725,N_9342);
nand UO_553 (O_553,N_9555,N_9152);
and UO_554 (O_554,N_9054,N_9618);
and UO_555 (O_555,N_9624,N_9174);
xnor UO_556 (O_556,N_9708,N_9337);
xnor UO_557 (O_557,N_9599,N_9039);
and UO_558 (O_558,N_9815,N_9193);
xor UO_559 (O_559,N_9179,N_9704);
nor UO_560 (O_560,N_9578,N_9560);
nor UO_561 (O_561,N_9050,N_9478);
or UO_562 (O_562,N_9547,N_9524);
or UO_563 (O_563,N_9870,N_9751);
xnor UO_564 (O_564,N_9079,N_9238);
nand UO_565 (O_565,N_9610,N_9489);
or UO_566 (O_566,N_9155,N_9900);
and UO_567 (O_567,N_9557,N_9914);
nand UO_568 (O_568,N_9345,N_9413);
or UO_569 (O_569,N_9509,N_9147);
nand UO_570 (O_570,N_9307,N_9409);
or UO_571 (O_571,N_9006,N_9477);
nand UO_572 (O_572,N_9709,N_9119);
or UO_573 (O_573,N_9198,N_9262);
nor UO_574 (O_574,N_9624,N_9725);
or UO_575 (O_575,N_9225,N_9446);
nor UO_576 (O_576,N_9942,N_9451);
xor UO_577 (O_577,N_9096,N_9727);
nand UO_578 (O_578,N_9951,N_9939);
xnor UO_579 (O_579,N_9885,N_9019);
and UO_580 (O_580,N_9108,N_9767);
or UO_581 (O_581,N_9760,N_9465);
or UO_582 (O_582,N_9542,N_9214);
nand UO_583 (O_583,N_9420,N_9241);
or UO_584 (O_584,N_9419,N_9011);
xnor UO_585 (O_585,N_9212,N_9279);
xor UO_586 (O_586,N_9211,N_9051);
nor UO_587 (O_587,N_9751,N_9951);
nor UO_588 (O_588,N_9999,N_9747);
nand UO_589 (O_589,N_9993,N_9720);
and UO_590 (O_590,N_9884,N_9803);
xnor UO_591 (O_591,N_9930,N_9540);
or UO_592 (O_592,N_9781,N_9682);
or UO_593 (O_593,N_9479,N_9641);
nand UO_594 (O_594,N_9493,N_9049);
or UO_595 (O_595,N_9485,N_9344);
nand UO_596 (O_596,N_9645,N_9266);
or UO_597 (O_597,N_9471,N_9709);
xnor UO_598 (O_598,N_9941,N_9272);
and UO_599 (O_599,N_9868,N_9317);
xor UO_600 (O_600,N_9724,N_9412);
or UO_601 (O_601,N_9409,N_9432);
and UO_602 (O_602,N_9698,N_9944);
nand UO_603 (O_603,N_9442,N_9063);
nand UO_604 (O_604,N_9448,N_9017);
xor UO_605 (O_605,N_9473,N_9042);
nand UO_606 (O_606,N_9075,N_9681);
xnor UO_607 (O_607,N_9344,N_9609);
and UO_608 (O_608,N_9704,N_9153);
xnor UO_609 (O_609,N_9903,N_9602);
and UO_610 (O_610,N_9891,N_9282);
and UO_611 (O_611,N_9389,N_9759);
xor UO_612 (O_612,N_9972,N_9136);
xor UO_613 (O_613,N_9004,N_9873);
xnor UO_614 (O_614,N_9036,N_9323);
xnor UO_615 (O_615,N_9305,N_9433);
and UO_616 (O_616,N_9269,N_9679);
and UO_617 (O_617,N_9656,N_9947);
nor UO_618 (O_618,N_9829,N_9696);
nand UO_619 (O_619,N_9358,N_9144);
or UO_620 (O_620,N_9515,N_9029);
or UO_621 (O_621,N_9476,N_9661);
xor UO_622 (O_622,N_9864,N_9904);
or UO_623 (O_623,N_9451,N_9176);
and UO_624 (O_624,N_9685,N_9665);
xor UO_625 (O_625,N_9030,N_9533);
and UO_626 (O_626,N_9349,N_9196);
xnor UO_627 (O_627,N_9482,N_9112);
or UO_628 (O_628,N_9531,N_9278);
nor UO_629 (O_629,N_9464,N_9662);
xnor UO_630 (O_630,N_9775,N_9022);
or UO_631 (O_631,N_9127,N_9344);
and UO_632 (O_632,N_9050,N_9591);
xor UO_633 (O_633,N_9337,N_9541);
nor UO_634 (O_634,N_9349,N_9973);
xor UO_635 (O_635,N_9142,N_9811);
nor UO_636 (O_636,N_9124,N_9912);
nor UO_637 (O_637,N_9334,N_9568);
nor UO_638 (O_638,N_9170,N_9505);
nor UO_639 (O_639,N_9963,N_9180);
nor UO_640 (O_640,N_9008,N_9214);
nor UO_641 (O_641,N_9471,N_9206);
nand UO_642 (O_642,N_9997,N_9524);
xnor UO_643 (O_643,N_9076,N_9339);
and UO_644 (O_644,N_9567,N_9671);
nand UO_645 (O_645,N_9109,N_9190);
nand UO_646 (O_646,N_9922,N_9624);
xnor UO_647 (O_647,N_9532,N_9380);
nor UO_648 (O_648,N_9101,N_9629);
and UO_649 (O_649,N_9544,N_9875);
nand UO_650 (O_650,N_9379,N_9270);
or UO_651 (O_651,N_9356,N_9814);
xor UO_652 (O_652,N_9275,N_9643);
nand UO_653 (O_653,N_9796,N_9834);
nor UO_654 (O_654,N_9724,N_9118);
and UO_655 (O_655,N_9918,N_9243);
nand UO_656 (O_656,N_9197,N_9567);
and UO_657 (O_657,N_9438,N_9636);
nor UO_658 (O_658,N_9585,N_9907);
and UO_659 (O_659,N_9425,N_9434);
nand UO_660 (O_660,N_9385,N_9354);
and UO_661 (O_661,N_9363,N_9404);
nand UO_662 (O_662,N_9826,N_9473);
nor UO_663 (O_663,N_9315,N_9837);
nand UO_664 (O_664,N_9014,N_9420);
nand UO_665 (O_665,N_9843,N_9377);
or UO_666 (O_666,N_9222,N_9271);
nor UO_667 (O_667,N_9025,N_9603);
and UO_668 (O_668,N_9845,N_9878);
and UO_669 (O_669,N_9583,N_9658);
xnor UO_670 (O_670,N_9590,N_9752);
nand UO_671 (O_671,N_9917,N_9970);
or UO_672 (O_672,N_9734,N_9377);
nand UO_673 (O_673,N_9194,N_9897);
nor UO_674 (O_674,N_9011,N_9752);
or UO_675 (O_675,N_9088,N_9478);
and UO_676 (O_676,N_9843,N_9173);
and UO_677 (O_677,N_9787,N_9371);
xor UO_678 (O_678,N_9513,N_9820);
or UO_679 (O_679,N_9616,N_9640);
nor UO_680 (O_680,N_9177,N_9497);
or UO_681 (O_681,N_9531,N_9849);
nor UO_682 (O_682,N_9369,N_9651);
or UO_683 (O_683,N_9212,N_9379);
nand UO_684 (O_684,N_9454,N_9059);
nand UO_685 (O_685,N_9256,N_9713);
or UO_686 (O_686,N_9095,N_9061);
xor UO_687 (O_687,N_9668,N_9787);
and UO_688 (O_688,N_9781,N_9848);
xnor UO_689 (O_689,N_9719,N_9985);
or UO_690 (O_690,N_9963,N_9179);
nand UO_691 (O_691,N_9443,N_9128);
or UO_692 (O_692,N_9842,N_9470);
and UO_693 (O_693,N_9678,N_9568);
nor UO_694 (O_694,N_9095,N_9351);
and UO_695 (O_695,N_9299,N_9640);
nand UO_696 (O_696,N_9376,N_9246);
xor UO_697 (O_697,N_9847,N_9561);
or UO_698 (O_698,N_9961,N_9437);
nor UO_699 (O_699,N_9320,N_9993);
xnor UO_700 (O_700,N_9229,N_9333);
nor UO_701 (O_701,N_9906,N_9591);
nor UO_702 (O_702,N_9427,N_9613);
nand UO_703 (O_703,N_9623,N_9110);
nand UO_704 (O_704,N_9378,N_9185);
or UO_705 (O_705,N_9917,N_9736);
and UO_706 (O_706,N_9913,N_9823);
nor UO_707 (O_707,N_9052,N_9237);
nand UO_708 (O_708,N_9623,N_9217);
or UO_709 (O_709,N_9307,N_9148);
or UO_710 (O_710,N_9647,N_9473);
xor UO_711 (O_711,N_9264,N_9746);
nor UO_712 (O_712,N_9188,N_9082);
and UO_713 (O_713,N_9023,N_9015);
and UO_714 (O_714,N_9066,N_9137);
nor UO_715 (O_715,N_9403,N_9973);
or UO_716 (O_716,N_9734,N_9691);
xnor UO_717 (O_717,N_9439,N_9694);
and UO_718 (O_718,N_9264,N_9818);
or UO_719 (O_719,N_9836,N_9849);
nor UO_720 (O_720,N_9706,N_9247);
and UO_721 (O_721,N_9002,N_9288);
and UO_722 (O_722,N_9381,N_9784);
or UO_723 (O_723,N_9343,N_9548);
nand UO_724 (O_724,N_9523,N_9692);
and UO_725 (O_725,N_9965,N_9807);
xor UO_726 (O_726,N_9526,N_9918);
or UO_727 (O_727,N_9133,N_9572);
xnor UO_728 (O_728,N_9406,N_9379);
xnor UO_729 (O_729,N_9810,N_9821);
nor UO_730 (O_730,N_9987,N_9511);
xnor UO_731 (O_731,N_9673,N_9414);
and UO_732 (O_732,N_9637,N_9042);
xnor UO_733 (O_733,N_9783,N_9754);
or UO_734 (O_734,N_9069,N_9227);
nor UO_735 (O_735,N_9080,N_9815);
nand UO_736 (O_736,N_9838,N_9012);
and UO_737 (O_737,N_9688,N_9265);
nor UO_738 (O_738,N_9903,N_9724);
nand UO_739 (O_739,N_9275,N_9114);
nor UO_740 (O_740,N_9300,N_9427);
or UO_741 (O_741,N_9467,N_9846);
nor UO_742 (O_742,N_9849,N_9015);
xor UO_743 (O_743,N_9958,N_9552);
and UO_744 (O_744,N_9757,N_9259);
nand UO_745 (O_745,N_9666,N_9954);
or UO_746 (O_746,N_9986,N_9393);
xor UO_747 (O_747,N_9267,N_9326);
or UO_748 (O_748,N_9114,N_9051);
or UO_749 (O_749,N_9998,N_9836);
nor UO_750 (O_750,N_9450,N_9010);
nand UO_751 (O_751,N_9766,N_9036);
nor UO_752 (O_752,N_9120,N_9209);
nand UO_753 (O_753,N_9168,N_9216);
nor UO_754 (O_754,N_9533,N_9415);
xor UO_755 (O_755,N_9540,N_9210);
or UO_756 (O_756,N_9738,N_9021);
or UO_757 (O_757,N_9728,N_9457);
xor UO_758 (O_758,N_9734,N_9309);
and UO_759 (O_759,N_9231,N_9435);
or UO_760 (O_760,N_9561,N_9589);
or UO_761 (O_761,N_9817,N_9531);
and UO_762 (O_762,N_9839,N_9195);
and UO_763 (O_763,N_9548,N_9015);
nand UO_764 (O_764,N_9529,N_9339);
or UO_765 (O_765,N_9412,N_9887);
or UO_766 (O_766,N_9932,N_9080);
nand UO_767 (O_767,N_9100,N_9216);
nand UO_768 (O_768,N_9513,N_9778);
xnor UO_769 (O_769,N_9443,N_9173);
or UO_770 (O_770,N_9371,N_9113);
xor UO_771 (O_771,N_9224,N_9476);
nand UO_772 (O_772,N_9348,N_9127);
or UO_773 (O_773,N_9666,N_9310);
nor UO_774 (O_774,N_9134,N_9730);
or UO_775 (O_775,N_9670,N_9179);
or UO_776 (O_776,N_9090,N_9317);
nand UO_777 (O_777,N_9656,N_9904);
xnor UO_778 (O_778,N_9599,N_9943);
and UO_779 (O_779,N_9521,N_9303);
nor UO_780 (O_780,N_9076,N_9002);
nand UO_781 (O_781,N_9850,N_9243);
xnor UO_782 (O_782,N_9169,N_9069);
or UO_783 (O_783,N_9544,N_9511);
and UO_784 (O_784,N_9365,N_9582);
nor UO_785 (O_785,N_9990,N_9406);
or UO_786 (O_786,N_9085,N_9331);
nor UO_787 (O_787,N_9046,N_9320);
nor UO_788 (O_788,N_9951,N_9668);
and UO_789 (O_789,N_9080,N_9220);
and UO_790 (O_790,N_9311,N_9540);
nand UO_791 (O_791,N_9941,N_9513);
nand UO_792 (O_792,N_9275,N_9208);
nand UO_793 (O_793,N_9150,N_9052);
xnor UO_794 (O_794,N_9800,N_9946);
xor UO_795 (O_795,N_9079,N_9214);
or UO_796 (O_796,N_9554,N_9928);
nor UO_797 (O_797,N_9473,N_9009);
and UO_798 (O_798,N_9143,N_9804);
nor UO_799 (O_799,N_9375,N_9197);
nand UO_800 (O_800,N_9716,N_9426);
or UO_801 (O_801,N_9310,N_9446);
nand UO_802 (O_802,N_9789,N_9195);
or UO_803 (O_803,N_9046,N_9040);
nand UO_804 (O_804,N_9293,N_9746);
and UO_805 (O_805,N_9828,N_9460);
and UO_806 (O_806,N_9411,N_9516);
or UO_807 (O_807,N_9525,N_9193);
nand UO_808 (O_808,N_9783,N_9490);
xor UO_809 (O_809,N_9650,N_9601);
and UO_810 (O_810,N_9274,N_9152);
xnor UO_811 (O_811,N_9831,N_9256);
and UO_812 (O_812,N_9655,N_9743);
or UO_813 (O_813,N_9688,N_9434);
or UO_814 (O_814,N_9945,N_9128);
xor UO_815 (O_815,N_9829,N_9810);
nor UO_816 (O_816,N_9457,N_9606);
and UO_817 (O_817,N_9882,N_9184);
nor UO_818 (O_818,N_9118,N_9487);
nand UO_819 (O_819,N_9226,N_9856);
nand UO_820 (O_820,N_9831,N_9674);
and UO_821 (O_821,N_9764,N_9857);
nand UO_822 (O_822,N_9510,N_9414);
nor UO_823 (O_823,N_9169,N_9710);
and UO_824 (O_824,N_9886,N_9767);
xnor UO_825 (O_825,N_9017,N_9190);
or UO_826 (O_826,N_9642,N_9068);
xor UO_827 (O_827,N_9793,N_9259);
xor UO_828 (O_828,N_9169,N_9306);
nor UO_829 (O_829,N_9413,N_9472);
and UO_830 (O_830,N_9931,N_9106);
and UO_831 (O_831,N_9814,N_9852);
and UO_832 (O_832,N_9818,N_9725);
or UO_833 (O_833,N_9682,N_9628);
nand UO_834 (O_834,N_9250,N_9024);
nor UO_835 (O_835,N_9435,N_9767);
or UO_836 (O_836,N_9845,N_9315);
nand UO_837 (O_837,N_9520,N_9476);
nor UO_838 (O_838,N_9573,N_9592);
or UO_839 (O_839,N_9530,N_9409);
nor UO_840 (O_840,N_9050,N_9951);
nand UO_841 (O_841,N_9066,N_9371);
and UO_842 (O_842,N_9314,N_9629);
xnor UO_843 (O_843,N_9759,N_9364);
nor UO_844 (O_844,N_9523,N_9913);
and UO_845 (O_845,N_9972,N_9816);
and UO_846 (O_846,N_9057,N_9706);
or UO_847 (O_847,N_9415,N_9984);
xnor UO_848 (O_848,N_9767,N_9586);
nand UO_849 (O_849,N_9290,N_9270);
nand UO_850 (O_850,N_9910,N_9540);
nand UO_851 (O_851,N_9149,N_9989);
or UO_852 (O_852,N_9503,N_9558);
nand UO_853 (O_853,N_9121,N_9605);
and UO_854 (O_854,N_9719,N_9074);
nand UO_855 (O_855,N_9775,N_9386);
nand UO_856 (O_856,N_9083,N_9471);
nand UO_857 (O_857,N_9637,N_9661);
nor UO_858 (O_858,N_9779,N_9488);
nand UO_859 (O_859,N_9634,N_9770);
xor UO_860 (O_860,N_9884,N_9887);
and UO_861 (O_861,N_9183,N_9807);
nand UO_862 (O_862,N_9026,N_9201);
and UO_863 (O_863,N_9146,N_9756);
and UO_864 (O_864,N_9927,N_9528);
nor UO_865 (O_865,N_9889,N_9822);
and UO_866 (O_866,N_9201,N_9039);
nand UO_867 (O_867,N_9907,N_9769);
and UO_868 (O_868,N_9214,N_9703);
xor UO_869 (O_869,N_9636,N_9807);
nor UO_870 (O_870,N_9466,N_9705);
nor UO_871 (O_871,N_9208,N_9465);
xor UO_872 (O_872,N_9952,N_9422);
nor UO_873 (O_873,N_9239,N_9840);
nand UO_874 (O_874,N_9864,N_9756);
or UO_875 (O_875,N_9390,N_9554);
nor UO_876 (O_876,N_9166,N_9161);
or UO_877 (O_877,N_9680,N_9148);
or UO_878 (O_878,N_9539,N_9208);
or UO_879 (O_879,N_9306,N_9855);
xnor UO_880 (O_880,N_9415,N_9206);
or UO_881 (O_881,N_9750,N_9515);
xor UO_882 (O_882,N_9356,N_9000);
xor UO_883 (O_883,N_9558,N_9816);
nand UO_884 (O_884,N_9413,N_9017);
and UO_885 (O_885,N_9269,N_9684);
xor UO_886 (O_886,N_9906,N_9111);
xor UO_887 (O_887,N_9371,N_9547);
nand UO_888 (O_888,N_9647,N_9406);
nand UO_889 (O_889,N_9102,N_9249);
nand UO_890 (O_890,N_9867,N_9406);
nor UO_891 (O_891,N_9595,N_9192);
and UO_892 (O_892,N_9507,N_9321);
xor UO_893 (O_893,N_9337,N_9328);
nor UO_894 (O_894,N_9402,N_9170);
xor UO_895 (O_895,N_9145,N_9610);
nor UO_896 (O_896,N_9946,N_9040);
xor UO_897 (O_897,N_9732,N_9024);
nand UO_898 (O_898,N_9386,N_9179);
or UO_899 (O_899,N_9276,N_9092);
or UO_900 (O_900,N_9308,N_9185);
xnor UO_901 (O_901,N_9923,N_9621);
nand UO_902 (O_902,N_9685,N_9175);
and UO_903 (O_903,N_9662,N_9727);
and UO_904 (O_904,N_9828,N_9379);
and UO_905 (O_905,N_9705,N_9963);
nand UO_906 (O_906,N_9658,N_9520);
nand UO_907 (O_907,N_9656,N_9010);
nor UO_908 (O_908,N_9189,N_9328);
nor UO_909 (O_909,N_9423,N_9197);
xor UO_910 (O_910,N_9999,N_9841);
nand UO_911 (O_911,N_9118,N_9213);
or UO_912 (O_912,N_9254,N_9371);
xnor UO_913 (O_913,N_9590,N_9055);
xor UO_914 (O_914,N_9482,N_9714);
nand UO_915 (O_915,N_9111,N_9694);
nand UO_916 (O_916,N_9441,N_9254);
xor UO_917 (O_917,N_9574,N_9495);
nor UO_918 (O_918,N_9023,N_9817);
or UO_919 (O_919,N_9316,N_9632);
nand UO_920 (O_920,N_9761,N_9251);
or UO_921 (O_921,N_9414,N_9360);
nor UO_922 (O_922,N_9146,N_9729);
nor UO_923 (O_923,N_9808,N_9989);
and UO_924 (O_924,N_9553,N_9360);
xor UO_925 (O_925,N_9716,N_9906);
xnor UO_926 (O_926,N_9984,N_9233);
or UO_927 (O_927,N_9376,N_9628);
nor UO_928 (O_928,N_9689,N_9334);
and UO_929 (O_929,N_9980,N_9894);
and UO_930 (O_930,N_9159,N_9331);
xor UO_931 (O_931,N_9311,N_9191);
xor UO_932 (O_932,N_9709,N_9320);
or UO_933 (O_933,N_9290,N_9055);
and UO_934 (O_934,N_9097,N_9063);
and UO_935 (O_935,N_9046,N_9533);
nor UO_936 (O_936,N_9762,N_9111);
and UO_937 (O_937,N_9749,N_9716);
and UO_938 (O_938,N_9884,N_9743);
xor UO_939 (O_939,N_9085,N_9872);
and UO_940 (O_940,N_9646,N_9274);
or UO_941 (O_941,N_9269,N_9135);
or UO_942 (O_942,N_9976,N_9068);
or UO_943 (O_943,N_9533,N_9605);
xnor UO_944 (O_944,N_9479,N_9092);
and UO_945 (O_945,N_9507,N_9374);
xnor UO_946 (O_946,N_9350,N_9984);
nand UO_947 (O_947,N_9161,N_9164);
or UO_948 (O_948,N_9036,N_9981);
or UO_949 (O_949,N_9121,N_9014);
and UO_950 (O_950,N_9982,N_9333);
nor UO_951 (O_951,N_9427,N_9202);
nand UO_952 (O_952,N_9429,N_9175);
xor UO_953 (O_953,N_9316,N_9130);
xor UO_954 (O_954,N_9694,N_9332);
xor UO_955 (O_955,N_9230,N_9303);
and UO_956 (O_956,N_9106,N_9454);
nand UO_957 (O_957,N_9526,N_9015);
xnor UO_958 (O_958,N_9149,N_9002);
or UO_959 (O_959,N_9361,N_9078);
and UO_960 (O_960,N_9042,N_9588);
nand UO_961 (O_961,N_9896,N_9163);
xor UO_962 (O_962,N_9514,N_9233);
nor UO_963 (O_963,N_9181,N_9114);
nor UO_964 (O_964,N_9059,N_9372);
xor UO_965 (O_965,N_9197,N_9531);
or UO_966 (O_966,N_9647,N_9316);
and UO_967 (O_967,N_9501,N_9450);
xor UO_968 (O_968,N_9467,N_9400);
nor UO_969 (O_969,N_9767,N_9637);
and UO_970 (O_970,N_9721,N_9384);
and UO_971 (O_971,N_9068,N_9780);
or UO_972 (O_972,N_9800,N_9522);
nand UO_973 (O_973,N_9411,N_9718);
nor UO_974 (O_974,N_9683,N_9162);
nor UO_975 (O_975,N_9092,N_9107);
xnor UO_976 (O_976,N_9821,N_9886);
or UO_977 (O_977,N_9812,N_9571);
xnor UO_978 (O_978,N_9604,N_9539);
and UO_979 (O_979,N_9203,N_9454);
and UO_980 (O_980,N_9672,N_9675);
or UO_981 (O_981,N_9766,N_9631);
and UO_982 (O_982,N_9994,N_9760);
nand UO_983 (O_983,N_9403,N_9148);
xnor UO_984 (O_984,N_9024,N_9507);
nand UO_985 (O_985,N_9807,N_9604);
or UO_986 (O_986,N_9158,N_9184);
nand UO_987 (O_987,N_9171,N_9302);
or UO_988 (O_988,N_9873,N_9394);
nand UO_989 (O_989,N_9215,N_9670);
xor UO_990 (O_990,N_9498,N_9442);
xor UO_991 (O_991,N_9532,N_9895);
nand UO_992 (O_992,N_9230,N_9222);
xor UO_993 (O_993,N_9890,N_9028);
xor UO_994 (O_994,N_9982,N_9920);
nand UO_995 (O_995,N_9399,N_9751);
or UO_996 (O_996,N_9720,N_9018);
or UO_997 (O_997,N_9323,N_9356);
or UO_998 (O_998,N_9961,N_9146);
xor UO_999 (O_999,N_9180,N_9802);
xor UO_1000 (O_1000,N_9077,N_9566);
xnor UO_1001 (O_1001,N_9791,N_9678);
nand UO_1002 (O_1002,N_9479,N_9770);
or UO_1003 (O_1003,N_9553,N_9000);
nor UO_1004 (O_1004,N_9071,N_9451);
xnor UO_1005 (O_1005,N_9470,N_9047);
xnor UO_1006 (O_1006,N_9540,N_9467);
and UO_1007 (O_1007,N_9080,N_9162);
nand UO_1008 (O_1008,N_9649,N_9662);
or UO_1009 (O_1009,N_9750,N_9615);
xor UO_1010 (O_1010,N_9777,N_9343);
or UO_1011 (O_1011,N_9360,N_9895);
nor UO_1012 (O_1012,N_9687,N_9569);
and UO_1013 (O_1013,N_9306,N_9809);
or UO_1014 (O_1014,N_9272,N_9742);
nand UO_1015 (O_1015,N_9718,N_9602);
xnor UO_1016 (O_1016,N_9324,N_9102);
xor UO_1017 (O_1017,N_9793,N_9680);
nor UO_1018 (O_1018,N_9922,N_9253);
and UO_1019 (O_1019,N_9597,N_9826);
or UO_1020 (O_1020,N_9617,N_9446);
or UO_1021 (O_1021,N_9715,N_9730);
xor UO_1022 (O_1022,N_9546,N_9524);
or UO_1023 (O_1023,N_9187,N_9644);
nor UO_1024 (O_1024,N_9041,N_9689);
and UO_1025 (O_1025,N_9632,N_9988);
or UO_1026 (O_1026,N_9250,N_9408);
and UO_1027 (O_1027,N_9988,N_9330);
xor UO_1028 (O_1028,N_9556,N_9860);
nor UO_1029 (O_1029,N_9901,N_9181);
and UO_1030 (O_1030,N_9911,N_9095);
and UO_1031 (O_1031,N_9340,N_9408);
nor UO_1032 (O_1032,N_9487,N_9560);
nand UO_1033 (O_1033,N_9284,N_9480);
xnor UO_1034 (O_1034,N_9324,N_9980);
and UO_1035 (O_1035,N_9944,N_9826);
and UO_1036 (O_1036,N_9918,N_9633);
xnor UO_1037 (O_1037,N_9939,N_9955);
and UO_1038 (O_1038,N_9791,N_9815);
nand UO_1039 (O_1039,N_9181,N_9587);
and UO_1040 (O_1040,N_9160,N_9006);
xor UO_1041 (O_1041,N_9906,N_9174);
and UO_1042 (O_1042,N_9986,N_9595);
nand UO_1043 (O_1043,N_9081,N_9228);
nand UO_1044 (O_1044,N_9499,N_9928);
xnor UO_1045 (O_1045,N_9571,N_9274);
or UO_1046 (O_1046,N_9847,N_9611);
nor UO_1047 (O_1047,N_9433,N_9063);
nand UO_1048 (O_1048,N_9361,N_9161);
or UO_1049 (O_1049,N_9739,N_9565);
and UO_1050 (O_1050,N_9375,N_9171);
and UO_1051 (O_1051,N_9341,N_9083);
or UO_1052 (O_1052,N_9314,N_9274);
or UO_1053 (O_1053,N_9813,N_9855);
xor UO_1054 (O_1054,N_9779,N_9234);
nor UO_1055 (O_1055,N_9958,N_9754);
or UO_1056 (O_1056,N_9778,N_9071);
or UO_1057 (O_1057,N_9419,N_9638);
nor UO_1058 (O_1058,N_9770,N_9219);
and UO_1059 (O_1059,N_9966,N_9492);
nand UO_1060 (O_1060,N_9521,N_9110);
nand UO_1061 (O_1061,N_9110,N_9295);
and UO_1062 (O_1062,N_9838,N_9228);
and UO_1063 (O_1063,N_9456,N_9310);
or UO_1064 (O_1064,N_9965,N_9720);
nor UO_1065 (O_1065,N_9304,N_9069);
nor UO_1066 (O_1066,N_9253,N_9109);
nand UO_1067 (O_1067,N_9063,N_9240);
nor UO_1068 (O_1068,N_9879,N_9806);
xnor UO_1069 (O_1069,N_9281,N_9857);
nor UO_1070 (O_1070,N_9710,N_9926);
and UO_1071 (O_1071,N_9860,N_9968);
or UO_1072 (O_1072,N_9215,N_9065);
nor UO_1073 (O_1073,N_9546,N_9632);
xor UO_1074 (O_1074,N_9175,N_9171);
xnor UO_1075 (O_1075,N_9918,N_9256);
or UO_1076 (O_1076,N_9015,N_9405);
or UO_1077 (O_1077,N_9058,N_9790);
or UO_1078 (O_1078,N_9669,N_9855);
nand UO_1079 (O_1079,N_9057,N_9210);
nor UO_1080 (O_1080,N_9965,N_9094);
and UO_1081 (O_1081,N_9163,N_9834);
nor UO_1082 (O_1082,N_9117,N_9851);
or UO_1083 (O_1083,N_9187,N_9288);
or UO_1084 (O_1084,N_9372,N_9195);
nor UO_1085 (O_1085,N_9959,N_9756);
and UO_1086 (O_1086,N_9332,N_9235);
or UO_1087 (O_1087,N_9444,N_9903);
or UO_1088 (O_1088,N_9150,N_9633);
xnor UO_1089 (O_1089,N_9982,N_9246);
or UO_1090 (O_1090,N_9767,N_9820);
nand UO_1091 (O_1091,N_9641,N_9913);
or UO_1092 (O_1092,N_9533,N_9967);
nand UO_1093 (O_1093,N_9941,N_9729);
nand UO_1094 (O_1094,N_9062,N_9261);
xnor UO_1095 (O_1095,N_9687,N_9577);
and UO_1096 (O_1096,N_9511,N_9366);
or UO_1097 (O_1097,N_9587,N_9114);
or UO_1098 (O_1098,N_9120,N_9900);
or UO_1099 (O_1099,N_9569,N_9132);
nor UO_1100 (O_1100,N_9125,N_9487);
and UO_1101 (O_1101,N_9293,N_9127);
nor UO_1102 (O_1102,N_9953,N_9272);
xnor UO_1103 (O_1103,N_9161,N_9903);
or UO_1104 (O_1104,N_9280,N_9601);
or UO_1105 (O_1105,N_9371,N_9309);
xnor UO_1106 (O_1106,N_9693,N_9308);
nor UO_1107 (O_1107,N_9046,N_9157);
nand UO_1108 (O_1108,N_9682,N_9904);
and UO_1109 (O_1109,N_9872,N_9258);
and UO_1110 (O_1110,N_9303,N_9789);
nand UO_1111 (O_1111,N_9703,N_9456);
nand UO_1112 (O_1112,N_9454,N_9735);
and UO_1113 (O_1113,N_9864,N_9757);
xor UO_1114 (O_1114,N_9880,N_9350);
and UO_1115 (O_1115,N_9619,N_9735);
nor UO_1116 (O_1116,N_9318,N_9620);
nand UO_1117 (O_1117,N_9964,N_9085);
nor UO_1118 (O_1118,N_9730,N_9773);
and UO_1119 (O_1119,N_9810,N_9341);
nand UO_1120 (O_1120,N_9729,N_9583);
or UO_1121 (O_1121,N_9208,N_9202);
xnor UO_1122 (O_1122,N_9776,N_9741);
xnor UO_1123 (O_1123,N_9060,N_9313);
xnor UO_1124 (O_1124,N_9131,N_9763);
and UO_1125 (O_1125,N_9623,N_9261);
xor UO_1126 (O_1126,N_9112,N_9723);
xnor UO_1127 (O_1127,N_9871,N_9604);
nand UO_1128 (O_1128,N_9826,N_9883);
nand UO_1129 (O_1129,N_9773,N_9705);
nor UO_1130 (O_1130,N_9676,N_9383);
nor UO_1131 (O_1131,N_9665,N_9508);
and UO_1132 (O_1132,N_9551,N_9614);
xor UO_1133 (O_1133,N_9839,N_9996);
or UO_1134 (O_1134,N_9757,N_9838);
xnor UO_1135 (O_1135,N_9443,N_9582);
and UO_1136 (O_1136,N_9623,N_9306);
and UO_1137 (O_1137,N_9825,N_9126);
or UO_1138 (O_1138,N_9326,N_9252);
nor UO_1139 (O_1139,N_9429,N_9652);
nand UO_1140 (O_1140,N_9542,N_9225);
and UO_1141 (O_1141,N_9317,N_9459);
and UO_1142 (O_1142,N_9918,N_9641);
nand UO_1143 (O_1143,N_9694,N_9907);
nor UO_1144 (O_1144,N_9969,N_9201);
xnor UO_1145 (O_1145,N_9522,N_9377);
nand UO_1146 (O_1146,N_9775,N_9896);
nand UO_1147 (O_1147,N_9822,N_9863);
nor UO_1148 (O_1148,N_9441,N_9524);
or UO_1149 (O_1149,N_9377,N_9057);
nand UO_1150 (O_1150,N_9197,N_9414);
or UO_1151 (O_1151,N_9207,N_9434);
nor UO_1152 (O_1152,N_9149,N_9750);
nor UO_1153 (O_1153,N_9567,N_9833);
or UO_1154 (O_1154,N_9107,N_9312);
nand UO_1155 (O_1155,N_9044,N_9096);
xor UO_1156 (O_1156,N_9836,N_9186);
nor UO_1157 (O_1157,N_9378,N_9793);
and UO_1158 (O_1158,N_9653,N_9375);
or UO_1159 (O_1159,N_9381,N_9839);
and UO_1160 (O_1160,N_9855,N_9955);
or UO_1161 (O_1161,N_9712,N_9838);
xor UO_1162 (O_1162,N_9432,N_9477);
nor UO_1163 (O_1163,N_9488,N_9210);
or UO_1164 (O_1164,N_9467,N_9506);
nor UO_1165 (O_1165,N_9030,N_9425);
nor UO_1166 (O_1166,N_9158,N_9853);
nor UO_1167 (O_1167,N_9294,N_9382);
or UO_1168 (O_1168,N_9707,N_9938);
nor UO_1169 (O_1169,N_9902,N_9755);
nand UO_1170 (O_1170,N_9056,N_9847);
or UO_1171 (O_1171,N_9642,N_9964);
and UO_1172 (O_1172,N_9185,N_9144);
and UO_1173 (O_1173,N_9368,N_9188);
nor UO_1174 (O_1174,N_9090,N_9947);
or UO_1175 (O_1175,N_9435,N_9587);
xnor UO_1176 (O_1176,N_9262,N_9211);
or UO_1177 (O_1177,N_9348,N_9998);
nor UO_1178 (O_1178,N_9691,N_9005);
xnor UO_1179 (O_1179,N_9876,N_9761);
nand UO_1180 (O_1180,N_9536,N_9153);
nor UO_1181 (O_1181,N_9002,N_9023);
and UO_1182 (O_1182,N_9611,N_9834);
nand UO_1183 (O_1183,N_9186,N_9224);
nor UO_1184 (O_1184,N_9852,N_9395);
nor UO_1185 (O_1185,N_9643,N_9985);
and UO_1186 (O_1186,N_9127,N_9935);
nand UO_1187 (O_1187,N_9428,N_9064);
or UO_1188 (O_1188,N_9818,N_9483);
or UO_1189 (O_1189,N_9435,N_9136);
nand UO_1190 (O_1190,N_9211,N_9155);
nor UO_1191 (O_1191,N_9388,N_9728);
and UO_1192 (O_1192,N_9257,N_9939);
xor UO_1193 (O_1193,N_9090,N_9303);
nor UO_1194 (O_1194,N_9374,N_9693);
and UO_1195 (O_1195,N_9964,N_9989);
nand UO_1196 (O_1196,N_9063,N_9781);
nor UO_1197 (O_1197,N_9907,N_9032);
or UO_1198 (O_1198,N_9297,N_9571);
nor UO_1199 (O_1199,N_9158,N_9602);
and UO_1200 (O_1200,N_9253,N_9202);
and UO_1201 (O_1201,N_9257,N_9146);
and UO_1202 (O_1202,N_9044,N_9992);
or UO_1203 (O_1203,N_9789,N_9761);
xnor UO_1204 (O_1204,N_9488,N_9219);
or UO_1205 (O_1205,N_9408,N_9419);
or UO_1206 (O_1206,N_9933,N_9471);
nor UO_1207 (O_1207,N_9617,N_9068);
nor UO_1208 (O_1208,N_9673,N_9094);
nor UO_1209 (O_1209,N_9611,N_9189);
xnor UO_1210 (O_1210,N_9909,N_9669);
or UO_1211 (O_1211,N_9828,N_9651);
nor UO_1212 (O_1212,N_9324,N_9442);
nand UO_1213 (O_1213,N_9168,N_9222);
nand UO_1214 (O_1214,N_9645,N_9028);
nand UO_1215 (O_1215,N_9512,N_9592);
xnor UO_1216 (O_1216,N_9644,N_9135);
and UO_1217 (O_1217,N_9024,N_9365);
or UO_1218 (O_1218,N_9561,N_9954);
nand UO_1219 (O_1219,N_9363,N_9377);
nor UO_1220 (O_1220,N_9551,N_9825);
xor UO_1221 (O_1221,N_9219,N_9265);
nand UO_1222 (O_1222,N_9665,N_9805);
and UO_1223 (O_1223,N_9569,N_9740);
or UO_1224 (O_1224,N_9681,N_9056);
xor UO_1225 (O_1225,N_9257,N_9274);
xnor UO_1226 (O_1226,N_9510,N_9587);
xnor UO_1227 (O_1227,N_9956,N_9772);
xnor UO_1228 (O_1228,N_9844,N_9654);
and UO_1229 (O_1229,N_9216,N_9139);
nor UO_1230 (O_1230,N_9722,N_9079);
xor UO_1231 (O_1231,N_9071,N_9568);
and UO_1232 (O_1232,N_9803,N_9391);
nor UO_1233 (O_1233,N_9312,N_9361);
and UO_1234 (O_1234,N_9610,N_9890);
and UO_1235 (O_1235,N_9136,N_9848);
or UO_1236 (O_1236,N_9731,N_9465);
nand UO_1237 (O_1237,N_9739,N_9473);
or UO_1238 (O_1238,N_9642,N_9254);
nand UO_1239 (O_1239,N_9868,N_9796);
or UO_1240 (O_1240,N_9450,N_9386);
xor UO_1241 (O_1241,N_9319,N_9262);
or UO_1242 (O_1242,N_9410,N_9210);
or UO_1243 (O_1243,N_9831,N_9561);
and UO_1244 (O_1244,N_9852,N_9042);
nor UO_1245 (O_1245,N_9929,N_9201);
and UO_1246 (O_1246,N_9383,N_9428);
nand UO_1247 (O_1247,N_9126,N_9799);
xor UO_1248 (O_1248,N_9657,N_9601);
nand UO_1249 (O_1249,N_9217,N_9076);
nand UO_1250 (O_1250,N_9672,N_9080);
xnor UO_1251 (O_1251,N_9926,N_9649);
and UO_1252 (O_1252,N_9876,N_9693);
nor UO_1253 (O_1253,N_9016,N_9582);
or UO_1254 (O_1254,N_9209,N_9589);
nand UO_1255 (O_1255,N_9030,N_9069);
and UO_1256 (O_1256,N_9085,N_9461);
nand UO_1257 (O_1257,N_9070,N_9422);
xor UO_1258 (O_1258,N_9274,N_9003);
or UO_1259 (O_1259,N_9528,N_9818);
nand UO_1260 (O_1260,N_9363,N_9528);
xor UO_1261 (O_1261,N_9014,N_9421);
or UO_1262 (O_1262,N_9152,N_9591);
and UO_1263 (O_1263,N_9637,N_9187);
or UO_1264 (O_1264,N_9829,N_9228);
and UO_1265 (O_1265,N_9811,N_9792);
xor UO_1266 (O_1266,N_9273,N_9180);
or UO_1267 (O_1267,N_9741,N_9981);
nor UO_1268 (O_1268,N_9765,N_9088);
nor UO_1269 (O_1269,N_9684,N_9369);
nor UO_1270 (O_1270,N_9601,N_9690);
nor UO_1271 (O_1271,N_9910,N_9614);
nand UO_1272 (O_1272,N_9875,N_9441);
nand UO_1273 (O_1273,N_9014,N_9472);
and UO_1274 (O_1274,N_9979,N_9151);
xor UO_1275 (O_1275,N_9729,N_9539);
xor UO_1276 (O_1276,N_9920,N_9187);
or UO_1277 (O_1277,N_9945,N_9625);
or UO_1278 (O_1278,N_9533,N_9520);
and UO_1279 (O_1279,N_9647,N_9838);
and UO_1280 (O_1280,N_9388,N_9691);
nand UO_1281 (O_1281,N_9204,N_9422);
nor UO_1282 (O_1282,N_9705,N_9825);
xor UO_1283 (O_1283,N_9566,N_9749);
nand UO_1284 (O_1284,N_9868,N_9606);
nor UO_1285 (O_1285,N_9199,N_9859);
nand UO_1286 (O_1286,N_9148,N_9247);
and UO_1287 (O_1287,N_9023,N_9368);
and UO_1288 (O_1288,N_9563,N_9175);
xor UO_1289 (O_1289,N_9448,N_9258);
and UO_1290 (O_1290,N_9822,N_9203);
nand UO_1291 (O_1291,N_9134,N_9280);
or UO_1292 (O_1292,N_9282,N_9990);
nand UO_1293 (O_1293,N_9250,N_9934);
or UO_1294 (O_1294,N_9810,N_9748);
xnor UO_1295 (O_1295,N_9532,N_9171);
nand UO_1296 (O_1296,N_9384,N_9244);
nand UO_1297 (O_1297,N_9761,N_9662);
xnor UO_1298 (O_1298,N_9998,N_9924);
xnor UO_1299 (O_1299,N_9886,N_9579);
nand UO_1300 (O_1300,N_9164,N_9405);
and UO_1301 (O_1301,N_9990,N_9886);
xnor UO_1302 (O_1302,N_9358,N_9149);
nand UO_1303 (O_1303,N_9365,N_9683);
and UO_1304 (O_1304,N_9158,N_9908);
xnor UO_1305 (O_1305,N_9702,N_9848);
and UO_1306 (O_1306,N_9626,N_9386);
xnor UO_1307 (O_1307,N_9452,N_9922);
nand UO_1308 (O_1308,N_9029,N_9709);
nor UO_1309 (O_1309,N_9569,N_9581);
nor UO_1310 (O_1310,N_9946,N_9653);
xnor UO_1311 (O_1311,N_9182,N_9748);
nor UO_1312 (O_1312,N_9247,N_9466);
and UO_1313 (O_1313,N_9957,N_9618);
or UO_1314 (O_1314,N_9052,N_9663);
or UO_1315 (O_1315,N_9813,N_9940);
nor UO_1316 (O_1316,N_9028,N_9101);
nor UO_1317 (O_1317,N_9228,N_9703);
xor UO_1318 (O_1318,N_9498,N_9454);
and UO_1319 (O_1319,N_9264,N_9384);
nor UO_1320 (O_1320,N_9651,N_9776);
xnor UO_1321 (O_1321,N_9289,N_9082);
and UO_1322 (O_1322,N_9785,N_9417);
and UO_1323 (O_1323,N_9414,N_9910);
or UO_1324 (O_1324,N_9560,N_9064);
nor UO_1325 (O_1325,N_9598,N_9950);
or UO_1326 (O_1326,N_9611,N_9147);
nor UO_1327 (O_1327,N_9126,N_9484);
and UO_1328 (O_1328,N_9274,N_9909);
and UO_1329 (O_1329,N_9969,N_9481);
nor UO_1330 (O_1330,N_9543,N_9291);
nor UO_1331 (O_1331,N_9709,N_9925);
or UO_1332 (O_1332,N_9445,N_9419);
xor UO_1333 (O_1333,N_9058,N_9728);
or UO_1334 (O_1334,N_9964,N_9679);
xnor UO_1335 (O_1335,N_9806,N_9158);
nor UO_1336 (O_1336,N_9084,N_9654);
nand UO_1337 (O_1337,N_9970,N_9350);
nor UO_1338 (O_1338,N_9474,N_9298);
nand UO_1339 (O_1339,N_9929,N_9040);
and UO_1340 (O_1340,N_9112,N_9980);
or UO_1341 (O_1341,N_9166,N_9193);
or UO_1342 (O_1342,N_9401,N_9641);
and UO_1343 (O_1343,N_9200,N_9039);
xor UO_1344 (O_1344,N_9349,N_9932);
nor UO_1345 (O_1345,N_9567,N_9556);
xnor UO_1346 (O_1346,N_9174,N_9386);
xor UO_1347 (O_1347,N_9309,N_9350);
xor UO_1348 (O_1348,N_9665,N_9528);
and UO_1349 (O_1349,N_9337,N_9476);
nand UO_1350 (O_1350,N_9853,N_9800);
and UO_1351 (O_1351,N_9250,N_9068);
xnor UO_1352 (O_1352,N_9216,N_9399);
xor UO_1353 (O_1353,N_9685,N_9616);
or UO_1354 (O_1354,N_9250,N_9280);
and UO_1355 (O_1355,N_9133,N_9625);
nor UO_1356 (O_1356,N_9981,N_9779);
and UO_1357 (O_1357,N_9787,N_9779);
nand UO_1358 (O_1358,N_9854,N_9966);
nand UO_1359 (O_1359,N_9091,N_9251);
nand UO_1360 (O_1360,N_9045,N_9129);
nor UO_1361 (O_1361,N_9460,N_9613);
or UO_1362 (O_1362,N_9079,N_9690);
nand UO_1363 (O_1363,N_9833,N_9389);
nand UO_1364 (O_1364,N_9815,N_9033);
nand UO_1365 (O_1365,N_9599,N_9317);
or UO_1366 (O_1366,N_9999,N_9424);
xnor UO_1367 (O_1367,N_9841,N_9258);
or UO_1368 (O_1368,N_9422,N_9629);
xor UO_1369 (O_1369,N_9305,N_9467);
nand UO_1370 (O_1370,N_9901,N_9161);
and UO_1371 (O_1371,N_9083,N_9789);
or UO_1372 (O_1372,N_9006,N_9686);
nor UO_1373 (O_1373,N_9621,N_9217);
and UO_1374 (O_1374,N_9824,N_9528);
xor UO_1375 (O_1375,N_9570,N_9419);
nand UO_1376 (O_1376,N_9458,N_9307);
and UO_1377 (O_1377,N_9185,N_9075);
xnor UO_1378 (O_1378,N_9756,N_9835);
and UO_1379 (O_1379,N_9073,N_9495);
or UO_1380 (O_1380,N_9486,N_9463);
nand UO_1381 (O_1381,N_9542,N_9652);
or UO_1382 (O_1382,N_9235,N_9496);
nand UO_1383 (O_1383,N_9476,N_9480);
nor UO_1384 (O_1384,N_9154,N_9176);
xnor UO_1385 (O_1385,N_9619,N_9229);
or UO_1386 (O_1386,N_9794,N_9051);
and UO_1387 (O_1387,N_9457,N_9463);
and UO_1388 (O_1388,N_9236,N_9581);
nand UO_1389 (O_1389,N_9815,N_9856);
and UO_1390 (O_1390,N_9253,N_9640);
xnor UO_1391 (O_1391,N_9380,N_9000);
or UO_1392 (O_1392,N_9815,N_9908);
nand UO_1393 (O_1393,N_9578,N_9695);
nor UO_1394 (O_1394,N_9071,N_9927);
nor UO_1395 (O_1395,N_9064,N_9982);
or UO_1396 (O_1396,N_9183,N_9044);
xor UO_1397 (O_1397,N_9035,N_9552);
nand UO_1398 (O_1398,N_9321,N_9701);
or UO_1399 (O_1399,N_9730,N_9652);
and UO_1400 (O_1400,N_9964,N_9550);
and UO_1401 (O_1401,N_9591,N_9871);
xor UO_1402 (O_1402,N_9916,N_9651);
or UO_1403 (O_1403,N_9668,N_9064);
and UO_1404 (O_1404,N_9510,N_9072);
nand UO_1405 (O_1405,N_9115,N_9617);
xnor UO_1406 (O_1406,N_9515,N_9085);
xor UO_1407 (O_1407,N_9174,N_9370);
and UO_1408 (O_1408,N_9724,N_9495);
and UO_1409 (O_1409,N_9816,N_9999);
and UO_1410 (O_1410,N_9288,N_9274);
nor UO_1411 (O_1411,N_9765,N_9724);
or UO_1412 (O_1412,N_9127,N_9805);
nand UO_1413 (O_1413,N_9474,N_9625);
nor UO_1414 (O_1414,N_9648,N_9770);
and UO_1415 (O_1415,N_9145,N_9685);
xnor UO_1416 (O_1416,N_9501,N_9992);
and UO_1417 (O_1417,N_9155,N_9521);
and UO_1418 (O_1418,N_9073,N_9294);
nand UO_1419 (O_1419,N_9930,N_9750);
and UO_1420 (O_1420,N_9359,N_9874);
and UO_1421 (O_1421,N_9636,N_9329);
xnor UO_1422 (O_1422,N_9407,N_9427);
nor UO_1423 (O_1423,N_9694,N_9044);
nor UO_1424 (O_1424,N_9325,N_9637);
xnor UO_1425 (O_1425,N_9805,N_9342);
nand UO_1426 (O_1426,N_9230,N_9061);
or UO_1427 (O_1427,N_9567,N_9764);
nor UO_1428 (O_1428,N_9360,N_9218);
nor UO_1429 (O_1429,N_9752,N_9174);
nand UO_1430 (O_1430,N_9758,N_9912);
and UO_1431 (O_1431,N_9478,N_9566);
or UO_1432 (O_1432,N_9306,N_9176);
nand UO_1433 (O_1433,N_9627,N_9588);
or UO_1434 (O_1434,N_9720,N_9774);
or UO_1435 (O_1435,N_9683,N_9054);
or UO_1436 (O_1436,N_9468,N_9067);
nand UO_1437 (O_1437,N_9855,N_9988);
xor UO_1438 (O_1438,N_9471,N_9494);
nor UO_1439 (O_1439,N_9171,N_9547);
nor UO_1440 (O_1440,N_9115,N_9798);
nand UO_1441 (O_1441,N_9175,N_9954);
or UO_1442 (O_1442,N_9296,N_9122);
and UO_1443 (O_1443,N_9331,N_9982);
or UO_1444 (O_1444,N_9557,N_9811);
xor UO_1445 (O_1445,N_9705,N_9428);
nor UO_1446 (O_1446,N_9791,N_9729);
or UO_1447 (O_1447,N_9951,N_9918);
and UO_1448 (O_1448,N_9303,N_9950);
or UO_1449 (O_1449,N_9572,N_9186);
nor UO_1450 (O_1450,N_9325,N_9674);
nand UO_1451 (O_1451,N_9517,N_9269);
nand UO_1452 (O_1452,N_9083,N_9342);
nor UO_1453 (O_1453,N_9726,N_9446);
nor UO_1454 (O_1454,N_9551,N_9405);
or UO_1455 (O_1455,N_9240,N_9059);
nand UO_1456 (O_1456,N_9966,N_9791);
or UO_1457 (O_1457,N_9836,N_9796);
xor UO_1458 (O_1458,N_9747,N_9702);
and UO_1459 (O_1459,N_9707,N_9287);
nand UO_1460 (O_1460,N_9029,N_9563);
nor UO_1461 (O_1461,N_9741,N_9983);
nand UO_1462 (O_1462,N_9956,N_9404);
or UO_1463 (O_1463,N_9681,N_9819);
nor UO_1464 (O_1464,N_9399,N_9385);
nor UO_1465 (O_1465,N_9521,N_9268);
nor UO_1466 (O_1466,N_9917,N_9805);
nor UO_1467 (O_1467,N_9009,N_9869);
and UO_1468 (O_1468,N_9204,N_9746);
or UO_1469 (O_1469,N_9705,N_9736);
and UO_1470 (O_1470,N_9074,N_9016);
and UO_1471 (O_1471,N_9099,N_9106);
xnor UO_1472 (O_1472,N_9417,N_9510);
nand UO_1473 (O_1473,N_9860,N_9441);
or UO_1474 (O_1474,N_9988,N_9926);
and UO_1475 (O_1475,N_9244,N_9751);
and UO_1476 (O_1476,N_9059,N_9842);
nand UO_1477 (O_1477,N_9384,N_9745);
xnor UO_1478 (O_1478,N_9507,N_9935);
nor UO_1479 (O_1479,N_9705,N_9922);
nand UO_1480 (O_1480,N_9524,N_9951);
and UO_1481 (O_1481,N_9223,N_9913);
xor UO_1482 (O_1482,N_9595,N_9362);
or UO_1483 (O_1483,N_9752,N_9213);
or UO_1484 (O_1484,N_9306,N_9191);
and UO_1485 (O_1485,N_9900,N_9271);
xnor UO_1486 (O_1486,N_9101,N_9828);
and UO_1487 (O_1487,N_9091,N_9223);
or UO_1488 (O_1488,N_9391,N_9053);
xor UO_1489 (O_1489,N_9714,N_9445);
nand UO_1490 (O_1490,N_9010,N_9314);
xor UO_1491 (O_1491,N_9813,N_9458);
nand UO_1492 (O_1492,N_9698,N_9473);
nand UO_1493 (O_1493,N_9178,N_9198);
or UO_1494 (O_1494,N_9522,N_9074);
or UO_1495 (O_1495,N_9797,N_9762);
nor UO_1496 (O_1496,N_9200,N_9793);
xor UO_1497 (O_1497,N_9852,N_9966);
nand UO_1498 (O_1498,N_9669,N_9437);
nor UO_1499 (O_1499,N_9344,N_9828);
endmodule