module basic_500_3000_500_6_levels_1xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_114,In_323);
or U1 (N_1,In_60,In_126);
nand U2 (N_2,In_62,In_395);
nand U3 (N_3,In_47,In_91);
nand U4 (N_4,In_473,In_454);
xnor U5 (N_5,In_362,In_210);
or U6 (N_6,In_41,In_327);
and U7 (N_7,In_484,In_198);
or U8 (N_8,In_200,In_292);
nor U9 (N_9,In_445,In_279);
nand U10 (N_10,In_178,In_312);
nor U11 (N_11,In_69,In_70);
and U12 (N_12,In_162,In_427);
nor U13 (N_13,In_9,In_486);
or U14 (N_14,In_461,In_274);
nor U15 (N_15,In_185,In_104);
nor U16 (N_16,In_251,In_230);
or U17 (N_17,In_197,In_453);
nand U18 (N_18,In_346,In_189);
nand U19 (N_19,In_388,In_144);
nand U20 (N_20,In_316,In_287);
and U21 (N_21,In_363,In_223);
nand U22 (N_22,In_171,In_353);
and U23 (N_23,In_406,In_478);
nor U24 (N_24,In_66,In_333);
nand U25 (N_25,In_277,In_293);
nor U26 (N_26,In_377,In_263);
or U27 (N_27,In_23,In_122);
and U28 (N_28,In_101,In_42);
nand U29 (N_29,In_494,In_205);
nor U30 (N_30,In_372,In_160);
nor U31 (N_31,In_402,In_225);
and U32 (N_32,In_100,In_102);
nor U33 (N_33,In_493,In_381);
or U34 (N_34,In_467,In_95);
nand U35 (N_35,In_89,In_439);
or U36 (N_36,In_284,In_375);
nand U37 (N_37,In_370,In_421);
nand U38 (N_38,In_246,In_79);
nand U39 (N_39,In_474,In_182);
and U40 (N_40,In_186,In_432);
and U41 (N_41,In_280,In_25);
nand U42 (N_42,In_255,In_350);
nor U43 (N_43,In_286,In_224);
nand U44 (N_44,In_368,In_465);
or U45 (N_45,In_308,In_7);
nand U46 (N_46,In_228,In_184);
nand U47 (N_47,In_499,In_260);
nand U48 (N_48,In_158,In_67);
and U49 (N_49,In_151,In_482);
and U50 (N_50,In_26,In_222);
nand U51 (N_51,In_218,In_455);
nand U52 (N_52,In_103,In_302);
nor U53 (N_53,In_27,In_12);
and U54 (N_54,In_65,In_366);
and U55 (N_55,In_249,In_40);
and U56 (N_56,In_492,In_305);
and U57 (N_57,In_146,In_397);
nand U58 (N_58,In_418,In_391);
nor U59 (N_59,In_342,In_219);
or U60 (N_60,In_19,In_409);
and U61 (N_61,In_275,In_108);
nor U62 (N_62,In_11,In_121);
xnor U63 (N_63,In_301,In_264);
xnor U64 (N_64,In_129,In_119);
nor U65 (N_65,In_125,In_63);
and U66 (N_66,In_30,In_360);
and U67 (N_67,In_242,In_426);
and U68 (N_68,In_236,In_425);
and U69 (N_69,In_221,In_152);
and U70 (N_70,In_481,In_206);
nor U71 (N_71,In_383,In_442);
or U72 (N_72,In_97,In_194);
nor U73 (N_73,In_64,In_38);
nor U74 (N_74,In_124,In_468);
and U75 (N_75,In_56,In_247);
nor U76 (N_76,In_78,In_273);
nor U77 (N_77,In_477,In_84);
nor U78 (N_78,In_299,In_32);
or U79 (N_79,In_334,In_6);
or U80 (N_80,In_433,In_234);
nand U81 (N_81,In_498,In_376);
and U82 (N_82,In_470,In_85);
or U83 (N_83,In_90,In_207);
nor U84 (N_84,In_39,In_357);
nand U85 (N_85,In_335,In_451);
or U86 (N_86,In_45,In_139);
and U87 (N_87,In_110,In_106);
nor U88 (N_88,In_488,In_438);
nor U89 (N_89,In_213,In_109);
nand U90 (N_90,In_52,In_138);
or U91 (N_91,In_303,In_460);
and U92 (N_92,In_289,In_140);
nand U93 (N_93,In_320,In_349);
nand U94 (N_94,In_183,In_414);
or U95 (N_95,In_319,In_233);
and U96 (N_96,In_44,In_252);
nor U97 (N_97,In_177,In_257);
nor U98 (N_98,In_94,In_336);
nand U99 (N_99,In_87,In_456);
or U100 (N_100,In_471,In_115);
or U101 (N_101,In_417,In_20);
nand U102 (N_102,In_459,In_322);
nor U103 (N_103,In_387,In_365);
and U104 (N_104,In_373,In_83);
nor U105 (N_105,In_338,In_36);
nor U106 (N_106,In_389,In_29);
nand U107 (N_107,In_49,In_297);
nand U108 (N_108,In_462,In_154);
nor U109 (N_109,In_440,In_169);
and U110 (N_110,In_295,In_328);
nor U111 (N_111,In_364,In_400);
nor U112 (N_112,In_396,In_340);
and U113 (N_113,In_410,In_201);
nand U114 (N_114,In_384,In_380);
and U115 (N_115,In_248,In_332);
nor U116 (N_116,In_398,In_86);
and U117 (N_117,In_261,In_485);
and U118 (N_118,In_361,In_192);
nor U119 (N_119,In_2,In_98);
and U120 (N_120,In_476,In_72);
nand U121 (N_121,In_188,In_120);
and U122 (N_122,In_318,In_16);
and U123 (N_123,In_428,In_155);
nor U124 (N_124,In_345,In_479);
nor U125 (N_125,In_475,In_325);
and U126 (N_126,In_176,In_227);
or U127 (N_127,In_276,In_163);
nor U128 (N_128,In_283,In_133);
nor U129 (N_129,In_130,In_422);
and U130 (N_130,In_281,In_168);
or U131 (N_131,In_76,In_212);
or U132 (N_132,In_226,In_173);
nor U133 (N_133,In_447,In_164);
and U134 (N_134,In_93,In_148);
and U135 (N_135,In_54,In_132);
and U136 (N_136,In_229,In_369);
or U137 (N_137,In_497,In_306);
and U138 (N_138,In_231,In_244);
or U139 (N_139,In_430,In_354);
and U140 (N_140,In_37,In_304);
nand U141 (N_141,In_43,In_238);
or U142 (N_142,In_250,In_240);
or U143 (N_143,In_167,In_436);
nand U144 (N_144,In_270,In_393);
and U145 (N_145,In_190,In_142);
and U146 (N_146,In_127,In_203);
nor U147 (N_147,In_495,In_339);
or U148 (N_148,In_416,In_408);
or U149 (N_149,In_399,In_131);
nand U150 (N_150,In_166,In_296);
or U151 (N_151,In_321,In_150);
and U152 (N_152,In_0,In_483);
nand U153 (N_153,In_385,In_143);
or U154 (N_154,In_187,In_256);
nor U155 (N_155,In_392,In_35);
or U156 (N_156,In_153,In_394);
or U157 (N_157,In_170,In_241);
and U158 (N_158,In_258,In_431);
xnor U159 (N_159,In_267,In_450);
nor U160 (N_160,In_435,In_282);
nor U161 (N_161,In_415,In_271);
nand U162 (N_162,In_31,In_217);
nand U163 (N_163,In_112,In_75);
or U164 (N_164,In_118,In_268);
or U165 (N_165,In_55,In_21);
or U166 (N_166,In_420,In_390);
or U167 (N_167,In_269,In_358);
nand U168 (N_168,In_294,In_337);
nand U169 (N_169,In_82,In_324);
and U170 (N_170,In_235,In_135);
nor U171 (N_171,In_330,In_208);
nand U172 (N_172,In_161,In_3);
and U173 (N_173,In_113,In_15);
nor U174 (N_174,In_180,In_480);
or U175 (N_175,In_266,In_172);
nor U176 (N_176,In_452,In_191);
or U177 (N_177,In_466,In_359);
nand U178 (N_178,In_204,In_272);
nor U179 (N_179,In_1,In_443);
nand U180 (N_180,In_331,In_179);
nor U181 (N_181,In_313,In_489);
nand U182 (N_182,In_117,In_457);
or U183 (N_183,In_254,In_10);
or U184 (N_184,In_134,In_50);
nor U185 (N_185,In_159,In_374);
nor U186 (N_186,In_449,In_199);
and U187 (N_187,In_278,In_496);
nand U188 (N_188,In_413,In_444);
nor U189 (N_189,In_472,In_237);
and U190 (N_190,In_28,In_193);
or U191 (N_191,In_259,In_53);
nor U192 (N_192,In_220,In_285);
or U193 (N_193,In_314,In_33);
nor U194 (N_194,In_352,In_262);
and U195 (N_195,In_215,In_51);
or U196 (N_196,In_92,In_5);
and U197 (N_197,In_73,In_348);
nor U198 (N_198,In_77,In_356);
or U199 (N_199,In_136,In_490);
or U200 (N_200,In_309,In_347);
nor U201 (N_201,In_423,In_446);
nand U202 (N_202,In_401,In_105);
nand U203 (N_203,In_96,In_441);
nor U204 (N_204,In_81,In_8);
or U205 (N_205,In_434,In_57);
or U206 (N_206,In_14,In_329);
nand U207 (N_207,In_24,In_59);
nor U208 (N_208,In_341,In_367);
nor U209 (N_209,In_239,In_165);
or U210 (N_210,In_379,In_403);
nand U211 (N_211,In_469,In_487);
or U212 (N_212,In_310,In_141);
nand U213 (N_213,In_174,In_371);
nand U214 (N_214,In_58,In_448);
nor U215 (N_215,In_147,In_46);
nand U216 (N_216,In_88,In_407);
or U217 (N_217,In_17,In_288);
and U218 (N_218,In_245,In_405);
nor U219 (N_219,In_68,In_343);
nand U220 (N_220,In_464,In_61);
or U221 (N_221,In_326,In_253);
or U222 (N_222,In_419,In_344);
and U223 (N_223,In_491,In_216);
and U224 (N_224,In_156,In_355);
and U225 (N_225,In_34,In_404);
nand U226 (N_226,In_214,In_137);
nand U227 (N_227,In_300,In_307);
nand U228 (N_228,In_458,In_424);
nand U229 (N_229,In_80,In_123);
and U230 (N_230,In_128,In_437);
nor U231 (N_231,In_411,In_22);
and U232 (N_232,In_13,In_317);
nor U233 (N_233,In_74,In_175);
nor U234 (N_234,In_290,In_386);
nor U235 (N_235,In_429,In_111);
and U236 (N_236,In_71,In_157);
or U237 (N_237,In_145,In_291);
and U238 (N_238,In_265,In_232);
nor U239 (N_239,In_382,In_149);
and U240 (N_240,In_48,In_463);
or U241 (N_241,In_4,In_196);
nand U242 (N_242,In_211,In_202);
or U243 (N_243,In_116,In_18);
nand U244 (N_244,In_412,In_243);
nor U245 (N_245,In_209,In_298);
nor U246 (N_246,In_99,In_315);
nand U247 (N_247,In_378,In_351);
and U248 (N_248,In_311,In_181);
nor U249 (N_249,In_107,In_195);
nand U250 (N_250,In_470,In_236);
nor U251 (N_251,In_13,In_44);
and U252 (N_252,In_155,In_173);
nor U253 (N_253,In_450,In_219);
or U254 (N_254,In_398,In_131);
nand U255 (N_255,In_220,In_379);
nor U256 (N_256,In_402,In_312);
or U257 (N_257,In_102,In_147);
and U258 (N_258,In_318,In_158);
nor U259 (N_259,In_3,In_153);
or U260 (N_260,In_23,In_52);
and U261 (N_261,In_24,In_155);
and U262 (N_262,In_135,In_129);
nor U263 (N_263,In_209,In_361);
or U264 (N_264,In_224,In_146);
or U265 (N_265,In_221,In_202);
and U266 (N_266,In_353,In_386);
nor U267 (N_267,In_414,In_195);
or U268 (N_268,In_268,In_354);
or U269 (N_269,In_225,In_339);
nor U270 (N_270,In_105,In_227);
and U271 (N_271,In_331,In_29);
nor U272 (N_272,In_125,In_212);
and U273 (N_273,In_136,In_187);
nand U274 (N_274,In_459,In_254);
or U275 (N_275,In_150,In_35);
nand U276 (N_276,In_143,In_283);
or U277 (N_277,In_169,In_256);
nor U278 (N_278,In_484,In_208);
nor U279 (N_279,In_263,In_368);
or U280 (N_280,In_359,In_106);
and U281 (N_281,In_199,In_122);
nor U282 (N_282,In_436,In_280);
nand U283 (N_283,In_312,In_69);
and U284 (N_284,In_281,In_27);
nor U285 (N_285,In_413,In_342);
nor U286 (N_286,In_171,In_333);
and U287 (N_287,In_44,In_177);
or U288 (N_288,In_359,In_490);
and U289 (N_289,In_255,In_66);
nor U290 (N_290,In_470,In_96);
or U291 (N_291,In_361,In_419);
or U292 (N_292,In_302,In_260);
and U293 (N_293,In_256,In_67);
nand U294 (N_294,In_18,In_430);
and U295 (N_295,In_165,In_472);
nor U296 (N_296,In_298,In_113);
or U297 (N_297,In_499,In_487);
or U298 (N_298,In_416,In_435);
nor U299 (N_299,In_229,In_433);
or U300 (N_300,In_420,In_212);
nor U301 (N_301,In_287,In_60);
nor U302 (N_302,In_108,In_72);
nor U303 (N_303,In_99,In_195);
or U304 (N_304,In_229,In_272);
or U305 (N_305,In_340,In_343);
nor U306 (N_306,In_40,In_112);
and U307 (N_307,In_466,In_298);
and U308 (N_308,In_319,In_164);
and U309 (N_309,In_37,In_419);
and U310 (N_310,In_122,In_298);
nor U311 (N_311,In_458,In_44);
nor U312 (N_312,In_231,In_65);
nand U313 (N_313,In_396,In_382);
or U314 (N_314,In_111,In_326);
nand U315 (N_315,In_359,In_208);
or U316 (N_316,In_124,In_108);
nand U317 (N_317,In_227,In_330);
or U318 (N_318,In_360,In_266);
or U319 (N_319,In_19,In_314);
nand U320 (N_320,In_260,In_61);
and U321 (N_321,In_34,In_187);
or U322 (N_322,In_222,In_427);
nor U323 (N_323,In_402,In_318);
and U324 (N_324,In_308,In_315);
or U325 (N_325,In_225,In_360);
or U326 (N_326,In_366,In_479);
and U327 (N_327,In_328,In_149);
and U328 (N_328,In_328,In_479);
nand U329 (N_329,In_387,In_109);
and U330 (N_330,In_421,In_227);
nand U331 (N_331,In_246,In_93);
and U332 (N_332,In_454,In_176);
nand U333 (N_333,In_474,In_267);
or U334 (N_334,In_341,In_59);
nand U335 (N_335,In_65,In_395);
nor U336 (N_336,In_74,In_249);
nand U337 (N_337,In_320,In_213);
or U338 (N_338,In_277,In_136);
or U339 (N_339,In_382,In_62);
or U340 (N_340,In_73,In_375);
nand U341 (N_341,In_199,In_437);
or U342 (N_342,In_221,In_109);
and U343 (N_343,In_180,In_243);
and U344 (N_344,In_200,In_308);
and U345 (N_345,In_487,In_411);
nand U346 (N_346,In_461,In_275);
nand U347 (N_347,In_315,In_14);
nand U348 (N_348,In_317,In_130);
or U349 (N_349,In_407,In_155);
or U350 (N_350,In_165,In_304);
and U351 (N_351,In_218,In_315);
nand U352 (N_352,In_385,In_453);
and U353 (N_353,In_154,In_394);
nand U354 (N_354,In_332,In_87);
nor U355 (N_355,In_398,In_207);
nor U356 (N_356,In_265,In_484);
nor U357 (N_357,In_34,In_88);
nor U358 (N_358,In_217,In_34);
or U359 (N_359,In_393,In_461);
and U360 (N_360,In_54,In_75);
or U361 (N_361,In_367,In_41);
nand U362 (N_362,In_154,In_425);
and U363 (N_363,In_12,In_137);
nand U364 (N_364,In_204,In_176);
and U365 (N_365,In_118,In_425);
and U366 (N_366,In_303,In_112);
nor U367 (N_367,In_10,In_358);
nor U368 (N_368,In_334,In_437);
or U369 (N_369,In_417,In_271);
nor U370 (N_370,In_93,In_12);
nand U371 (N_371,In_103,In_183);
nand U372 (N_372,In_151,In_94);
nor U373 (N_373,In_192,In_319);
nand U374 (N_374,In_144,In_422);
or U375 (N_375,In_180,In_23);
nor U376 (N_376,In_471,In_146);
and U377 (N_377,In_248,In_438);
nand U378 (N_378,In_453,In_227);
nor U379 (N_379,In_69,In_459);
nand U380 (N_380,In_293,In_4);
and U381 (N_381,In_489,In_347);
or U382 (N_382,In_154,In_153);
nor U383 (N_383,In_421,In_479);
nand U384 (N_384,In_481,In_385);
and U385 (N_385,In_336,In_129);
nor U386 (N_386,In_371,In_486);
nor U387 (N_387,In_253,In_175);
nor U388 (N_388,In_313,In_76);
nor U389 (N_389,In_320,In_371);
nor U390 (N_390,In_484,In_1);
and U391 (N_391,In_350,In_301);
and U392 (N_392,In_50,In_56);
and U393 (N_393,In_74,In_248);
nor U394 (N_394,In_405,In_203);
nor U395 (N_395,In_408,In_475);
nand U396 (N_396,In_102,In_1);
nand U397 (N_397,In_439,In_486);
and U398 (N_398,In_99,In_408);
and U399 (N_399,In_309,In_441);
nand U400 (N_400,In_405,In_427);
nor U401 (N_401,In_116,In_372);
nand U402 (N_402,In_125,In_218);
nand U403 (N_403,In_300,In_228);
or U404 (N_404,In_149,In_73);
and U405 (N_405,In_464,In_319);
nor U406 (N_406,In_135,In_295);
nor U407 (N_407,In_82,In_240);
nor U408 (N_408,In_137,In_89);
nor U409 (N_409,In_291,In_364);
nand U410 (N_410,In_286,In_193);
nand U411 (N_411,In_331,In_153);
nand U412 (N_412,In_373,In_143);
nand U413 (N_413,In_169,In_332);
or U414 (N_414,In_436,In_7);
and U415 (N_415,In_85,In_309);
nor U416 (N_416,In_194,In_49);
nor U417 (N_417,In_176,In_464);
nand U418 (N_418,In_52,In_113);
nor U419 (N_419,In_368,In_482);
and U420 (N_420,In_425,In_471);
nor U421 (N_421,In_32,In_381);
and U422 (N_422,In_387,In_355);
nand U423 (N_423,In_62,In_185);
nor U424 (N_424,In_350,In_382);
nor U425 (N_425,In_215,In_209);
or U426 (N_426,In_6,In_189);
nand U427 (N_427,In_212,In_195);
and U428 (N_428,In_312,In_281);
nor U429 (N_429,In_313,In_249);
and U430 (N_430,In_51,In_361);
nor U431 (N_431,In_27,In_180);
nand U432 (N_432,In_462,In_51);
nor U433 (N_433,In_107,In_301);
nand U434 (N_434,In_180,In_71);
nor U435 (N_435,In_483,In_254);
nand U436 (N_436,In_60,In_76);
nand U437 (N_437,In_263,In_91);
and U438 (N_438,In_4,In_86);
or U439 (N_439,In_134,In_125);
or U440 (N_440,In_208,In_498);
nand U441 (N_441,In_349,In_287);
nand U442 (N_442,In_468,In_453);
or U443 (N_443,In_56,In_15);
nor U444 (N_444,In_184,In_69);
nor U445 (N_445,In_482,In_44);
or U446 (N_446,In_432,In_41);
or U447 (N_447,In_456,In_39);
or U448 (N_448,In_0,In_130);
nand U449 (N_449,In_92,In_22);
nor U450 (N_450,In_305,In_347);
or U451 (N_451,In_426,In_7);
or U452 (N_452,In_485,In_284);
and U453 (N_453,In_316,In_40);
nand U454 (N_454,In_260,In_33);
or U455 (N_455,In_214,In_356);
or U456 (N_456,In_403,In_11);
and U457 (N_457,In_270,In_132);
and U458 (N_458,In_208,In_430);
or U459 (N_459,In_358,In_168);
nand U460 (N_460,In_228,In_461);
and U461 (N_461,In_244,In_391);
and U462 (N_462,In_298,In_431);
nor U463 (N_463,In_433,In_446);
and U464 (N_464,In_180,In_149);
nand U465 (N_465,In_156,In_398);
or U466 (N_466,In_268,In_186);
or U467 (N_467,In_209,In_49);
nand U468 (N_468,In_494,In_343);
nand U469 (N_469,In_333,In_323);
and U470 (N_470,In_419,In_467);
nor U471 (N_471,In_244,In_350);
and U472 (N_472,In_301,In_390);
nor U473 (N_473,In_302,In_140);
nor U474 (N_474,In_29,In_373);
or U475 (N_475,In_176,In_122);
or U476 (N_476,In_360,In_85);
nor U477 (N_477,In_370,In_114);
nor U478 (N_478,In_121,In_164);
nor U479 (N_479,In_309,In_92);
nand U480 (N_480,In_207,In_404);
or U481 (N_481,In_195,In_149);
and U482 (N_482,In_141,In_436);
nand U483 (N_483,In_223,In_163);
and U484 (N_484,In_332,In_403);
nand U485 (N_485,In_150,In_238);
nand U486 (N_486,In_356,In_0);
and U487 (N_487,In_249,In_305);
nand U488 (N_488,In_442,In_385);
or U489 (N_489,In_399,In_224);
nor U490 (N_490,In_327,In_200);
nand U491 (N_491,In_394,In_131);
nand U492 (N_492,In_169,In_469);
and U493 (N_493,In_402,In_37);
nand U494 (N_494,In_25,In_343);
or U495 (N_495,In_193,In_95);
nor U496 (N_496,In_378,In_392);
nand U497 (N_497,In_40,In_332);
and U498 (N_498,In_120,In_315);
xor U499 (N_499,In_340,In_411);
nand U500 (N_500,N_131,N_376);
nor U501 (N_501,N_264,N_234);
nand U502 (N_502,N_298,N_228);
nand U503 (N_503,N_107,N_144);
nand U504 (N_504,N_472,N_322);
nor U505 (N_505,N_72,N_377);
nand U506 (N_506,N_186,N_291);
nand U507 (N_507,N_270,N_450);
and U508 (N_508,N_118,N_425);
or U509 (N_509,N_256,N_277);
and U510 (N_510,N_61,N_143);
or U511 (N_511,N_310,N_76);
nor U512 (N_512,N_400,N_329);
or U513 (N_513,N_0,N_417);
or U514 (N_514,N_299,N_482);
nand U515 (N_515,N_427,N_140);
and U516 (N_516,N_134,N_338);
xnor U517 (N_517,N_240,N_94);
and U518 (N_518,N_163,N_415);
or U519 (N_519,N_261,N_403);
nand U520 (N_520,N_448,N_369);
nor U521 (N_521,N_60,N_89);
or U522 (N_522,N_31,N_388);
or U523 (N_523,N_458,N_405);
and U524 (N_524,N_193,N_386);
nand U525 (N_525,N_8,N_153);
nor U526 (N_526,N_232,N_187);
nor U527 (N_527,N_346,N_460);
or U528 (N_528,N_190,N_481);
or U529 (N_529,N_241,N_343);
nor U530 (N_530,N_429,N_10);
and U531 (N_531,N_81,N_401);
nand U532 (N_532,N_181,N_217);
nand U533 (N_533,N_274,N_29);
and U534 (N_534,N_473,N_244);
nor U535 (N_535,N_145,N_32);
or U536 (N_536,N_324,N_236);
and U537 (N_537,N_229,N_230);
xnor U538 (N_538,N_96,N_127);
and U539 (N_539,N_476,N_423);
or U540 (N_540,N_142,N_149);
nand U541 (N_541,N_320,N_119);
nand U542 (N_542,N_114,N_408);
nor U543 (N_543,N_286,N_316);
nand U544 (N_544,N_156,N_252);
and U545 (N_545,N_339,N_254);
or U546 (N_546,N_479,N_125);
or U547 (N_547,N_133,N_441);
and U548 (N_548,N_58,N_411);
nor U549 (N_549,N_260,N_311);
nor U550 (N_550,N_287,N_67);
nand U551 (N_551,N_20,N_259);
nor U552 (N_552,N_392,N_344);
and U553 (N_553,N_161,N_215);
nor U554 (N_554,N_273,N_21);
and U555 (N_555,N_88,N_359);
or U556 (N_556,N_211,N_435);
and U557 (N_557,N_51,N_253);
and U558 (N_558,N_50,N_185);
nand U559 (N_559,N_56,N_135);
nor U560 (N_560,N_440,N_251);
and U561 (N_561,N_182,N_381);
or U562 (N_562,N_166,N_465);
nand U563 (N_563,N_462,N_295);
and U564 (N_564,N_115,N_227);
and U565 (N_565,N_348,N_318);
nand U566 (N_566,N_70,N_188);
and U567 (N_567,N_98,N_255);
or U568 (N_568,N_378,N_396);
or U569 (N_569,N_432,N_213);
or U570 (N_570,N_453,N_148);
and U571 (N_571,N_41,N_113);
nor U572 (N_572,N_304,N_406);
nand U573 (N_573,N_24,N_2);
nand U574 (N_574,N_300,N_196);
or U575 (N_575,N_219,N_395);
nor U576 (N_576,N_34,N_201);
and U577 (N_577,N_293,N_202);
nand U578 (N_578,N_466,N_342);
or U579 (N_579,N_49,N_87);
and U580 (N_580,N_375,N_200);
nand U581 (N_581,N_99,N_484);
nor U582 (N_582,N_57,N_490);
nor U583 (N_583,N_111,N_266);
or U584 (N_584,N_86,N_282);
and U585 (N_585,N_357,N_223);
nor U586 (N_586,N_136,N_333);
nand U587 (N_587,N_120,N_55);
or U588 (N_588,N_416,N_75);
or U589 (N_589,N_306,N_433);
or U590 (N_590,N_170,N_38);
nor U591 (N_591,N_289,N_404);
or U592 (N_592,N_454,N_288);
or U593 (N_593,N_257,N_455);
nor U594 (N_594,N_319,N_474);
nand U595 (N_595,N_459,N_480);
nor U596 (N_596,N_285,N_48);
and U597 (N_597,N_340,N_13);
nor U598 (N_598,N_250,N_497);
and U599 (N_599,N_110,N_206);
nand U600 (N_600,N_297,N_189);
nor U601 (N_601,N_485,N_1);
or U602 (N_602,N_283,N_325);
nand U603 (N_603,N_45,N_390);
or U604 (N_604,N_457,N_197);
xnor U605 (N_605,N_27,N_362);
nand U606 (N_606,N_301,N_160);
nor U607 (N_607,N_470,N_246);
nand U608 (N_608,N_467,N_290);
nor U609 (N_609,N_93,N_90);
nand U610 (N_610,N_267,N_471);
or U611 (N_611,N_436,N_216);
or U612 (N_612,N_336,N_276);
nand U613 (N_613,N_245,N_428);
or U614 (N_614,N_430,N_350);
nand U615 (N_615,N_22,N_451);
or U616 (N_616,N_68,N_159);
or U617 (N_617,N_265,N_437);
nand U618 (N_618,N_494,N_103);
and U619 (N_619,N_370,N_317);
or U620 (N_620,N_360,N_397);
nand U621 (N_621,N_421,N_409);
nand U622 (N_622,N_139,N_272);
nand U623 (N_623,N_203,N_85);
nand U624 (N_624,N_207,N_194);
nor U625 (N_625,N_361,N_308);
nand U626 (N_626,N_43,N_180);
or U627 (N_627,N_199,N_468);
or U628 (N_628,N_422,N_358);
nor U629 (N_629,N_64,N_487);
nor U630 (N_630,N_78,N_19);
nor U631 (N_631,N_221,N_469);
nand U632 (N_632,N_493,N_249);
nor U633 (N_633,N_419,N_323);
nand U634 (N_634,N_198,N_205);
nor U635 (N_635,N_35,N_239);
and U636 (N_636,N_141,N_92);
xnor U637 (N_637,N_36,N_231);
nand U638 (N_638,N_373,N_498);
nand U639 (N_639,N_184,N_168);
and U640 (N_640,N_347,N_4);
or U641 (N_641,N_62,N_73);
or U642 (N_642,N_439,N_238);
and U643 (N_643,N_281,N_26);
nor U644 (N_644,N_157,N_69);
nand U645 (N_645,N_214,N_130);
nor U646 (N_646,N_52,N_183);
nor U647 (N_647,N_351,N_413);
or U648 (N_648,N_491,N_384);
nand U649 (N_649,N_258,N_383);
nor U650 (N_650,N_146,N_393);
and U651 (N_651,N_321,N_391);
nand U652 (N_652,N_109,N_30);
nor U653 (N_653,N_162,N_224);
nor U654 (N_654,N_444,N_6);
nand U655 (N_655,N_235,N_208);
nor U656 (N_656,N_334,N_164);
or U657 (N_657,N_499,N_464);
or U658 (N_658,N_363,N_175);
and U659 (N_659,N_284,N_495);
nor U660 (N_660,N_177,N_486);
nor U661 (N_661,N_488,N_121);
nand U662 (N_662,N_477,N_438);
or U663 (N_663,N_46,N_275);
nand U664 (N_664,N_65,N_167);
or U665 (N_665,N_332,N_105);
or U666 (N_666,N_366,N_151);
nand U667 (N_667,N_95,N_326);
xor U668 (N_668,N_442,N_3);
nor U669 (N_669,N_9,N_204);
or U670 (N_670,N_132,N_434);
nand U671 (N_671,N_101,N_44);
nor U672 (N_672,N_195,N_218);
or U673 (N_673,N_128,N_176);
nand U674 (N_674,N_302,N_47);
nor U675 (N_675,N_102,N_147);
and U676 (N_676,N_420,N_492);
or U677 (N_677,N_353,N_279);
and U678 (N_678,N_209,N_312);
nand U679 (N_679,N_226,N_305);
and U680 (N_680,N_337,N_233);
and U681 (N_681,N_398,N_372);
and U682 (N_682,N_445,N_16);
nor U683 (N_683,N_17,N_368);
nand U684 (N_684,N_100,N_155);
and U685 (N_685,N_210,N_414);
and U686 (N_686,N_174,N_379);
or U687 (N_687,N_447,N_475);
nor U688 (N_688,N_327,N_117);
nor U689 (N_689,N_278,N_399);
nor U690 (N_690,N_83,N_374);
nor U691 (N_691,N_303,N_394);
or U692 (N_692,N_426,N_39);
and U693 (N_693,N_313,N_371);
or U694 (N_694,N_489,N_382);
and U695 (N_695,N_63,N_367);
nand U696 (N_696,N_496,N_222);
or U697 (N_697,N_104,N_247);
or U698 (N_698,N_331,N_122);
nor U699 (N_699,N_463,N_106);
nor U700 (N_700,N_91,N_171);
and U701 (N_701,N_355,N_280);
nand U702 (N_702,N_315,N_356);
nor U703 (N_703,N_191,N_84);
or U704 (N_704,N_263,N_59);
nor U705 (N_705,N_28,N_33);
nand U706 (N_706,N_192,N_7);
nand U707 (N_707,N_40,N_354);
nor U708 (N_708,N_269,N_341);
nand U709 (N_709,N_23,N_179);
nor U710 (N_710,N_126,N_410);
nand U711 (N_711,N_54,N_129);
nand U712 (N_712,N_330,N_407);
and U713 (N_713,N_178,N_365);
and U714 (N_714,N_108,N_380);
nor U715 (N_715,N_173,N_387);
and U716 (N_716,N_412,N_74);
nor U717 (N_717,N_25,N_80);
nand U718 (N_718,N_150,N_15);
nand U719 (N_719,N_456,N_385);
nor U720 (N_720,N_237,N_82);
or U721 (N_721,N_123,N_53);
and U722 (N_722,N_165,N_116);
and U723 (N_723,N_66,N_328);
and U724 (N_724,N_307,N_225);
or U725 (N_725,N_172,N_483);
and U726 (N_726,N_268,N_77);
nand U727 (N_727,N_443,N_296);
or U728 (N_728,N_112,N_71);
and U729 (N_729,N_262,N_37);
or U730 (N_730,N_169,N_79);
nor U731 (N_731,N_212,N_452);
nor U732 (N_732,N_42,N_418);
nand U733 (N_733,N_124,N_11);
and U734 (N_734,N_294,N_138);
xor U735 (N_735,N_424,N_152);
and U736 (N_736,N_242,N_352);
or U737 (N_737,N_345,N_158);
or U738 (N_738,N_314,N_154);
or U739 (N_739,N_402,N_461);
and U740 (N_740,N_271,N_335);
nand U741 (N_741,N_220,N_431);
or U742 (N_742,N_349,N_5);
nor U743 (N_743,N_14,N_309);
and U744 (N_744,N_248,N_12);
or U745 (N_745,N_292,N_137);
or U746 (N_746,N_446,N_97);
and U747 (N_747,N_364,N_389);
nor U748 (N_748,N_478,N_18);
and U749 (N_749,N_449,N_243);
and U750 (N_750,N_246,N_24);
nand U751 (N_751,N_10,N_1);
or U752 (N_752,N_363,N_166);
nand U753 (N_753,N_155,N_421);
nand U754 (N_754,N_462,N_123);
nand U755 (N_755,N_330,N_221);
nand U756 (N_756,N_91,N_246);
or U757 (N_757,N_285,N_389);
nor U758 (N_758,N_220,N_472);
nor U759 (N_759,N_112,N_283);
nor U760 (N_760,N_337,N_48);
nor U761 (N_761,N_233,N_5);
and U762 (N_762,N_350,N_460);
or U763 (N_763,N_241,N_0);
or U764 (N_764,N_54,N_55);
nand U765 (N_765,N_34,N_204);
and U766 (N_766,N_373,N_371);
nor U767 (N_767,N_48,N_243);
and U768 (N_768,N_339,N_99);
nor U769 (N_769,N_134,N_387);
or U770 (N_770,N_151,N_144);
nor U771 (N_771,N_493,N_52);
or U772 (N_772,N_112,N_371);
nor U773 (N_773,N_28,N_286);
or U774 (N_774,N_316,N_242);
and U775 (N_775,N_424,N_435);
nor U776 (N_776,N_127,N_237);
or U777 (N_777,N_189,N_360);
and U778 (N_778,N_464,N_250);
and U779 (N_779,N_133,N_213);
or U780 (N_780,N_388,N_192);
nor U781 (N_781,N_277,N_65);
or U782 (N_782,N_74,N_35);
nor U783 (N_783,N_491,N_194);
or U784 (N_784,N_361,N_12);
nand U785 (N_785,N_334,N_29);
nand U786 (N_786,N_437,N_453);
or U787 (N_787,N_245,N_15);
nor U788 (N_788,N_170,N_489);
nand U789 (N_789,N_93,N_278);
nor U790 (N_790,N_465,N_134);
nand U791 (N_791,N_3,N_222);
nor U792 (N_792,N_321,N_236);
and U793 (N_793,N_86,N_197);
and U794 (N_794,N_285,N_61);
and U795 (N_795,N_324,N_279);
and U796 (N_796,N_164,N_230);
and U797 (N_797,N_61,N_457);
or U798 (N_798,N_443,N_391);
nor U799 (N_799,N_460,N_73);
nor U800 (N_800,N_185,N_61);
or U801 (N_801,N_405,N_480);
and U802 (N_802,N_438,N_379);
nand U803 (N_803,N_10,N_200);
or U804 (N_804,N_265,N_130);
nor U805 (N_805,N_51,N_41);
nor U806 (N_806,N_488,N_436);
nor U807 (N_807,N_437,N_242);
nand U808 (N_808,N_97,N_421);
and U809 (N_809,N_278,N_397);
or U810 (N_810,N_295,N_30);
nor U811 (N_811,N_193,N_107);
and U812 (N_812,N_160,N_451);
or U813 (N_813,N_161,N_373);
or U814 (N_814,N_121,N_435);
or U815 (N_815,N_185,N_192);
nor U816 (N_816,N_46,N_177);
and U817 (N_817,N_154,N_168);
or U818 (N_818,N_282,N_272);
and U819 (N_819,N_84,N_223);
nor U820 (N_820,N_9,N_386);
nor U821 (N_821,N_170,N_362);
and U822 (N_822,N_88,N_453);
nand U823 (N_823,N_328,N_59);
and U824 (N_824,N_443,N_466);
nor U825 (N_825,N_369,N_2);
nor U826 (N_826,N_416,N_173);
nor U827 (N_827,N_441,N_357);
and U828 (N_828,N_88,N_185);
nor U829 (N_829,N_108,N_344);
xnor U830 (N_830,N_370,N_295);
and U831 (N_831,N_260,N_65);
nor U832 (N_832,N_344,N_174);
nor U833 (N_833,N_317,N_166);
and U834 (N_834,N_315,N_185);
and U835 (N_835,N_291,N_39);
and U836 (N_836,N_59,N_273);
nand U837 (N_837,N_449,N_492);
and U838 (N_838,N_332,N_169);
nor U839 (N_839,N_129,N_378);
or U840 (N_840,N_412,N_123);
and U841 (N_841,N_448,N_267);
and U842 (N_842,N_98,N_403);
and U843 (N_843,N_252,N_29);
nor U844 (N_844,N_1,N_160);
or U845 (N_845,N_418,N_255);
nor U846 (N_846,N_418,N_50);
nor U847 (N_847,N_74,N_215);
and U848 (N_848,N_20,N_367);
xor U849 (N_849,N_422,N_266);
and U850 (N_850,N_304,N_147);
nand U851 (N_851,N_200,N_336);
nand U852 (N_852,N_219,N_280);
and U853 (N_853,N_380,N_8);
nor U854 (N_854,N_9,N_362);
or U855 (N_855,N_107,N_285);
or U856 (N_856,N_21,N_403);
or U857 (N_857,N_2,N_494);
nor U858 (N_858,N_231,N_457);
xnor U859 (N_859,N_88,N_105);
nor U860 (N_860,N_118,N_332);
nand U861 (N_861,N_89,N_355);
nand U862 (N_862,N_241,N_269);
nor U863 (N_863,N_174,N_374);
or U864 (N_864,N_322,N_140);
nor U865 (N_865,N_80,N_223);
and U866 (N_866,N_497,N_0);
nor U867 (N_867,N_292,N_134);
and U868 (N_868,N_498,N_44);
nor U869 (N_869,N_251,N_52);
and U870 (N_870,N_130,N_298);
nor U871 (N_871,N_34,N_296);
and U872 (N_872,N_364,N_37);
nor U873 (N_873,N_463,N_126);
or U874 (N_874,N_369,N_10);
nor U875 (N_875,N_416,N_54);
nor U876 (N_876,N_355,N_183);
nand U877 (N_877,N_286,N_438);
and U878 (N_878,N_489,N_93);
nor U879 (N_879,N_485,N_337);
and U880 (N_880,N_485,N_291);
and U881 (N_881,N_310,N_239);
nor U882 (N_882,N_114,N_262);
nor U883 (N_883,N_120,N_436);
or U884 (N_884,N_372,N_244);
nand U885 (N_885,N_334,N_489);
nor U886 (N_886,N_474,N_454);
nand U887 (N_887,N_263,N_256);
or U888 (N_888,N_118,N_373);
or U889 (N_889,N_461,N_40);
or U890 (N_890,N_74,N_184);
nor U891 (N_891,N_345,N_371);
nor U892 (N_892,N_385,N_186);
nor U893 (N_893,N_285,N_88);
nand U894 (N_894,N_218,N_43);
nor U895 (N_895,N_353,N_40);
nor U896 (N_896,N_424,N_280);
nor U897 (N_897,N_363,N_20);
and U898 (N_898,N_340,N_198);
and U899 (N_899,N_131,N_130);
or U900 (N_900,N_204,N_458);
and U901 (N_901,N_306,N_98);
and U902 (N_902,N_434,N_242);
and U903 (N_903,N_187,N_475);
and U904 (N_904,N_472,N_131);
or U905 (N_905,N_297,N_187);
nand U906 (N_906,N_421,N_338);
and U907 (N_907,N_257,N_202);
nor U908 (N_908,N_494,N_41);
nor U909 (N_909,N_17,N_196);
nor U910 (N_910,N_339,N_157);
nand U911 (N_911,N_229,N_311);
and U912 (N_912,N_290,N_279);
xnor U913 (N_913,N_393,N_406);
nand U914 (N_914,N_407,N_134);
and U915 (N_915,N_481,N_467);
nor U916 (N_916,N_92,N_229);
or U917 (N_917,N_89,N_292);
and U918 (N_918,N_405,N_164);
or U919 (N_919,N_60,N_225);
nor U920 (N_920,N_71,N_346);
nand U921 (N_921,N_101,N_150);
nand U922 (N_922,N_215,N_44);
nor U923 (N_923,N_247,N_432);
and U924 (N_924,N_336,N_410);
and U925 (N_925,N_266,N_325);
and U926 (N_926,N_303,N_7);
nand U927 (N_927,N_429,N_200);
and U928 (N_928,N_455,N_113);
nor U929 (N_929,N_70,N_391);
nand U930 (N_930,N_38,N_380);
nand U931 (N_931,N_457,N_79);
nand U932 (N_932,N_97,N_416);
and U933 (N_933,N_124,N_329);
nand U934 (N_934,N_141,N_245);
or U935 (N_935,N_164,N_489);
nor U936 (N_936,N_488,N_45);
and U937 (N_937,N_6,N_399);
nand U938 (N_938,N_45,N_146);
or U939 (N_939,N_386,N_237);
nor U940 (N_940,N_277,N_247);
nor U941 (N_941,N_69,N_119);
or U942 (N_942,N_428,N_465);
nand U943 (N_943,N_469,N_392);
nor U944 (N_944,N_238,N_437);
nor U945 (N_945,N_376,N_170);
or U946 (N_946,N_80,N_247);
nand U947 (N_947,N_433,N_357);
and U948 (N_948,N_482,N_81);
nand U949 (N_949,N_153,N_377);
and U950 (N_950,N_381,N_118);
xor U951 (N_951,N_300,N_123);
nor U952 (N_952,N_408,N_25);
nor U953 (N_953,N_16,N_17);
nand U954 (N_954,N_131,N_241);
nor U955 (N_955,N_26,N_122);
and U956 (N_956,N_230,N_109);
and U957 (N_957,N_254,N_226);
nor U958 (N_958,N_196,N_187);
nor U959 (N_959,N_10,N_301);
nand U960 (N_960,N_262,N_221);
nand U961 (N_961,N_238,N_216);
or U962 (N_962,N_197,N_118);
and U963 (N_963,N_173,N_191);
nor U964 (N_964,N_499,N_23);
or U965 (N_965,N_129,N_165);
and U966 (N_966,N_240,N_370);
nor U967 (N_967,N_292,N_400);
nand U968 (N_968,N_242,N_492);
nor U969 (N_969,N_287,N_459);
nand U970 (N_970,N_408,N_368);
or U971 (N_971,N_118,N_292);
nor U972 (N_972,N_413,N_312);
nand U973 (N_973,N_339,N_126);
nor U974 (N_974,N_345,N_327);
nor U975 (N_975,N_407,N_423);
and U976 (N_976,N_228,N_361);
and U977 (N_977,N_102,N_104);
nand U978 (N_978,N_76,N_184);
or U979 (N_979,N_42,N_282);
or U980 (N_980,N_105,N_452);
and U981 (N_981,N_370,N_285);
and U982 (N_982,N_232,N_220);
nand U983 (N_983,N_254,N_362);
nor U984 (N_984,N_428,N_19);
or U985 (N_985,N_378,N_437);
or U986 (N_986,N_221,N_184);
nand U987 (N_987,N_276,N_337);
or U988 (N_988,N_366,N_68);
nor U989 (N_989,N_415,N_38);
or U990 (N_990,N_253,N_159);
or U991 (N_991,N_87,N_466);
nor U992 (N_992,N_392,N_84);
nand U993 (N_993,N_127,N_87);
nand U994 (N_994,N_425,N_267);
or U995 (N_995,N_236,N_397);
nand U996 (N_996,N_25,N_425);
nor U997 (N_997,N_190,N_322);
or U998 (N_998,N_39,N_232);
or U999 (N_999,N_156,N_279);
nand U1000 (N_1000,N_801,N_505);
or U1001 (N_1001,N_639,N_675);
nand U1002 (N_1002,N_694,N_573);
nand U1003 (N_1003,N_773,N_654);
or U1004 (N_1004,N_670,N_788);
or U1005 (N_1005,N_542,N_893);
nor U1006 (N_1006,N_723,N_725);
or U1007 (N_1007,N_916,N_998);
and U1008 (N_1008,N_722,N_557);
nor U1009 (N_1009,N_648,N_881);
and U1010 (N_1010,N_958,N_930);
or U1011 (N_1011,N_949,N_671);
nor U1012 (N_1012,N_932,N_574);
nand U1013 (N_1013,N_592,N_527);
nand U1014 (N_1014,N_611,N_710);
nor U1015 (N_1015,N_552,N_892);
nand U1016 (N_1016,N_595,N_660);
nor U1017 (N_1017,N_735,N_709);
nor U1018 (N_1018,N_996,N_622);
nand U1019 (N_1019,N_524,N_697);
nor U1020 (N_1020,N_942,N_823);
nor U1021 (N_1021,N_793,N_685);
nor U1022 (N_1022,N_640,N_791);
nor U1023 (N_1023,N_668,N_577);
nand U1024 (N_1024,N_764,N_630);
nand U1025 (N_1025,N_575,N_727);
and U1026 (N_1026,N_978,N_604);
and U1027 (N_1027,N_845,N_726);
and U1028 (N_1028,N_976,N_692);
and U1029 (N_1029,N_812,N_681);
or U1030 (N_1030,N_646,N_861);
and U1031 (N_1031,N_866,N_927);
or U1032 (N_1032,N_848,N_761);
and U1033 (N_1033,N_997,N_880);
nand U1034 (N_1034,N_917,N_599);
or U1035 (N_1035,N_736,N_947);
nor U1036 (N_1036,N_840,N_663);
nand U1037 (N_1037,N_982,N_829);
nand U1038 (N_1038,N_642,N_683);
and U1039 (N_1039,N_855,N_854);
nand U1040 (N_1040,N_706,N_810);
nand U1041 (N_1041,N_826,N_730);
nor U1042 (N_1042,N_538,N_512);
nand U1043 (N_1043,N_568,N_924);
and U1044 (N_1044,N_547,N_655);
or U1045 (N_1045,N_563,N_669);
and U1046 (N_1046,N_621,N_689);
xor U1047 (N_1047,N_526,N_863);
nand U1048 (N_1048,N_853,N_939);
or U1049 (N_1049,N_799,N_545);
nor U1050 (N_1050,N_502,N_860);
or U1051 (N_1051,N_822,N_561);
nand U1052 (N_1052,N_914,N_973);
nor U1053 (N_1053,N_515,N_827);
or U1054 (N_1054,N_590,N_833);
and U1055 (N_1055,N_509,N_875);
or U1056 (N_1056,N_907,N_757);
or U1057 (N_1057,N_865,N_816);
or U1058 (N_1058,N_740,N_531);
nand U1059 (N_1059,N_532,N_904);
or U1060 (N_1060,N_558,N_748);
nand U1061 (N_1061,N_772,N_528);
or U1062 (N_1062,N_955,N_883);
xnor U1063 (N_1063,N_818,N_613);
or U1064 (N_1064,N_782,N_923);
and U1065 (N_1065,N_915,N_921);
or U1066 (N_1066,N_603,N_696);
and U1067 (N_1067,N_713,N_500);
and U1068 (N_1068,N_662,N_755);
nand U1069 (N_1069,N_790,N_898);
and U1070 (N_1070,N_806,N_828);
and U1071 (N_1071,N_744,N_800);
nor U1072 (N_1072,N_682,N_627);
nand U1073 (N_1073,N_597,N_733);
and U1074 (N_1074,N_843,N_503);
and U1075 (N_1075,N_677,N_514);
and U1076 (N_1076,N_536,N_644);
nor U1077 (N_1077,N_809,N_795);
nand U1078 (N_1078,N_605,N_580);
nor U1079 (N_1079,N_572,N_749);
or U1080 (N_1080,N_615,N_578);
and U1081 (N_1081,N_732,N_819);
nor U1082 (N_1082,N_541,N_925);
and U1083 (N_1083,N_598,N_811);
and U1084 (N_1084,N_762,N_581);
or U1085 (N_1085,N_956,N_784);
and U1086 (N_1086,N_564,N_868);
nand U1087 (N_1087,N_824,N_929);
and U1088 (N_1088,N_889,N_544);
nor U1089 (N_1089,N_678,N_873);
and U1090 (N_1090,N_775,N_712);
nand U1091 (N_1091,N_789,N_896);
or U1092 (N_1092,N_649,N_901);
nor U1093 (N_1093,N_551,N_647);
and U1094 (N_1094,N_959,N_624);
and U1095 (N_1095,N_543,N_767);
nor U1096 (N_1096,N_742,N_571);
or U1097 (N_1097,N_933,N_900);
nand U1098 (N_1098,N_862,N_588);
or U1099 (N_1099,N_867,N_886);
nand U1100 (N_1100,N_969,N_618);
nor U1101 (N_1101,N_659,N_807);
and U1102 (N_1102,N_501,N_815);
and U1103 (N_1103,N_708,N_535);
and U1104 (N_1104,N_747,N_817);
nor U1105 (N_1105,N_787,N_674);
nor U1106 (N_1106,N_842,N_877);
and U1107 (N_1107,N_928,N_641);
nand U1108 (N_1108,N_752,N_769);
nand U1109 (N_1109,N_596,N_802);
and U1110 (N_1110,N_879,N_852);
or U1111 (N_1111,N_995,N_768);
and U1112 (N_1112,N_651,N_684);
and U1113 (N_1113,N_513,N_583);
and U1114 (N_1114,N_984,N_794);
and U1115 (N_1115,N_688,N_864);
or U1116 (N_1116,N_779,N_946);
and U1117 (N_1117,N_602,N_922);
nand U1118 (N_1118,N_632,N_741);
nor U1119 (N_1119,N_972,N_834);
nand U1120 (N_1120,N_780,N_835);
or U1121 (N_1121,N_533,N_550);
nand U1122 (N_1122,N_693,N_771);
or U1123 (N_1123,N_715,N_970);
and U1124 (N_1124,N_620,N_954);
nor U1125 (N_1125,N_664,N_737);
nor U1126 (N_1126,N_600,N_638);
and U1127 (N_1127,N_971,N_560);
and U1128 (N_1128,N_555,N_792);
and U1129 (N_1129,N_980,N_825);
or U1130 (N_1130,N_738,N_576);
and U1131 (N_1131,N_776,N_656);
and U1132 (N_1132,N_781,N_556);
or U1133 (N_1133,N_909,N_628);
nor U1134 (N_1134,N_548,N_891);
nor U1135 (N_1135,N_546,N_520);
nand U1136 (N_1136,N_798,N_634);
and U1137 (N_1137,N_720,N_690);
nor U1138 (N_1138,N_832,N_841);
and U1139 (N_1139,N_945,N_756);
or U1140 (N_1140,N_797,N_814);
nand U1141 (N_1141,N_657,N_965);
nor U1142 (N_1142,N_607,N_619);
or U1143 (N_1143,N_510,N_871);
and U1144 (N_1144,N_585,N_796);
nand U1145 (N_1145,N_623,N_724);
and U1146 (N_1146,N_729,N_992);
or U1147 (N_1147,N_844,N_702);
and U1148 (N_1148,N_631,N_813);
nor U1149 (N_1149,N_918,N_616);
xnor U1150 (N_1150,N_988,N_948);
nor U1151 (N_1151,N_746,N_521);
and U1152 (N_1152,N_629,N_537);
and U1153 (N_1153,N_765,N_745);
or U1154 (N_1154,N_850,N_963);
nor U1155 (N_1155,N_858,N_643);
or U1156 (N_1156,N_977,N_601);
and U1157 (N_1157,N_872,N_687);
nor U1158 (N_1158,N_989,N_549);
and U1159 (N_1159,N_887,N_587);
nor U1160 (N_1160,N_523,N_808);
nor U1161 (N_1161,N_570,N_936);
and U1162 (N_1162,N_897,N_878);
and U1163 (N_1163,N_593,N_903);
or U1164 (N_1164,N_507,N_836);
or U1165 (N_1165,N_941,N_519);
and U1166 (N_1166,N_704,N_635);
nor U1167 (N_1167,N_987,N_703);
nor U1168 (N_1168,N_562,N_952);
or U1169 (N_1169,N_743,N_966);
nand U1170 (N_1170,N_721,N_940);
or U1171 (N_1171,N_803,N_985);
and U1172 (N_1172,N_511,N_837);
or U1173 (N_1173,N_739,N_758);
and U1174 (N_1174,N_943,N_874);
nand U1175 (N_1175,N_981,N_626);
nor U1176 (N_1176,N_934,N_565);
nor U1177 (N_1177,N_777,N_870);
and U1178 (N_1178,N_579,N_584);
nor U1179 (N_1179,N_633,N_888);
or U1180 (N_1180,N_979,N_516);
and U1181 (N_1181,N_964,N_680);
and U1182 (N_1182,N_957,N_566);
and U1183 (N_1183,N_691,N_983);
nand U1184 (N_1184,N_529,N_951);
or U1185 (N_1185,N_665,N_522);
and U1186 (N_1186,N_920,N_766);
nor U1187 (N_1187,N_778,N_658);
or U1188 (N_1188,N_695,N_763);
nand U1189 (N_1189,N_609,N_559);
nor U1190 (N_1190,N_913,N_999);
nor U1191 (N_1191,N_717,N_582);
nor U1192 (N_1192,N_770,N_591);
or U1193 (N_1193,N_567,N_719);
nor U1194 (N_1194,N_912,N_974);
and U1195 (N_1195,N_990,N_968);
nor U1196 (N_1196,N_991,N_760);
or U1197 (N_1197,N_851,N_950);
and U1198 (N_1198,N_540,N_589);
and U1199 (N_1199,N_650,N_857);
and U1200 (N_1200,N_938,N_919);
nor U1201 (N_1201,N_707,N_820);
nor U1202 (N_1202,N_849,N_884);
or U1203 (N_1203,N_653,N_847);
or U1204 (N_1204,N_804,N_839);
nor U1205 (N_1205,N_911,N_993);
nor U1206 (N_1206,N_508,N_783);
nor U1207 (N_1207,N_679,N_705);
and U1208 (N_1208,N_944,N_902);
and U1209 (N_1209,N_960,N_539);
nand U1210 (N_1210,N_869,N_805);
or U1211 (N_1211,N_753,N_935);
or U1212 (N_1212,N_838,N_554);
nor U1213 (N_1213,N_906,N_926);
nor U1214 (N_1214,N_899,N_625);
or U1215 (N_1215,N_734,N_885);
nand U1216 (N_1216,N_608,N_525);
nand U1217 (N_1217,N_645,N_910);
nor U1218 (N_1218,N_714,N_517);
nor U1219 (N_1219,N_931,N_937);
nand U1220 (N_1220,N_534,N_700);
nand U1221 (N_1221,N_594,N_672);
or U1222 (N_1222,N_967,N_831);
and U1223 (N_1223,N_986,N_711);
and U1224 (N_1224,N_859,N_673);
nand U1225 (N_1225,N_754,N_612);
and U1226 (N_1226,N_774,N_610);
nand U1227 (N_1227,N_504,N_882);
and U1228 (N_1228,N_718,N_894);
nand U1229 (N_1229,N_701,N_785);
nor U1230 (N_1230,N_606,N_750);
nor U1231 (N_1231,N_876,N_751);
nor U1232 (N_1232,N_716,N_905);
nand U1233 (N_1233,N_994,N_518);
and U1234 (N_1234,N_553,N_530);
nand U1235 (N_1235,N_652,N_759);
nand U1236 (N_1236,N_699,N_908);
nand U1237 (N_1237,N_961,N_661);
nand U1238 (N_1238,N_830,N_617);
nor U1239 (N_1239,N_953,N_637);
nor U1240 (N_1240,N_506,N_821);
and U1241 (N_1241,N_962,N_569);
or U1242 (N_1242,N_667,N_786);
nand U1243 (N_1243,N_676,N_698);
and U1244 (N_1244,N_666,N_895);
nor U1245 (N_1245,N_975,N_890);
and U1246 (N_1246,N_586,N_636);
nand U1247 (N_1247,N_731,N_614);
nor U1248 (N_1248,N_846,N_686);
or U1249 (N_1249,N_728,N_856);
and U1250 (N_1250,N_530,N_810);
nor U1251 (N_1251,N_851,N_616);
nor U1252 (N_1252,N_886,N_818);
or U1253 (N_1253,N_894,N_631);
or U1254 (N_1254,N_612,N_693);
nand U1255 (N_1255,N_835,N_555);
or U1256 (N_1256,N_814,N_687);
nor U1257 (N_1257,N_959,N_659);
or U1258 (N_1258,N_785,N_894);
nor U1259 (N_1259,N_721,N_973);
nand U1260 (N_1260,N_994,N_563);
nor U1261 (N_1261,N_580,N_810);
nand U1262 (N_1262,N_707,N_616);
or U1263 (N_1263,N_944,N_530);
nand U1264 (N_1264,N_993,N_598);
nor U1265 (N_1265,N_923,N_568);
nand U1266 (N_1266,N_522,N_583);
and U1267 (N_1267,N_927,N_873);
nor U1268 (N_1268,N_899,N_586);
nand U1269 (N_1269,N_627,N_707);
or U1270 (N_1270,N_855,N_823);
nand U1271 (N_1271,N_819,N_972);
nand U1272 (N_1272,N_976,N_956);
and U1273 (N_1273,N_964,N_589);
and U1274 (N_1274,N_961,N_680);
nand U1275 (N_1275,N_962,N_717);
or U1276 (N_1276,N_824,N_519);
nand U1277 (N_1277,N_999,N_767);
nor U1278 (N_1278,N_570,N_985);
or U1279 (N_1279,N_535,N_981);
and U1280 (N_1280,N_987,N_990);
nor U1281 (N_1281,N_650,N_511);
nor U1282 (N_1282,N_744,N_809);
nand U1283 (N_1283,N_857,N_965);
nand U1284 (N_1284,N_871,N_583);
nand U1285 (N_1285,N_890,N_737);
or U1286 (N_1286,N_529,N_669);
or U1287 (N_1287,N_977,N_695);
and U1288 (N_1288,N_804,N_815);
and U1289 (N_1289,N_531,N_937);
and U1290 (N_1290,N_939,N_696);
nand U1291 (N_1291,N_533,N_690);
nand U1292 (N_1292,N_908,N_953);
nand U1293 (N_1293,N_690,N_529);
nand U1294 (N_1294,N_550,N_597);
nand U1295 (N_1295,N_767,N_608);
and U1296 (N_1296,N_508,N_772);
nor U1297 (N_1297,N_520,N_600);
or U1298 (N_1298,N_697,N_825);
and U1299 (N_1299,N_542,N_935);
or U1300 (N_1300,N_503,N_942);
and U1301 (N_1301,N_888,N_897);
nand U1302 (N_1302,N_950,N_744);
nand U1303 (N_1303,N_954,N_818);
nand U1304 (N_1304,N_915,N_975);
or U1305 (N_1305,N_512,N_733);
nand U1306 (N_1306,N_816,N_570);
or U1307 (N_1307,N_524,N_889);
and U1308 (N_1308,N_602,N_675);
or U1309 (N_1309,N_943,N_528);
nand U1310 (N_1310,N_501,N_788);
and U1311 (N_1311,N_672,N_559);
and U1312 (N_1312,N_614,N_755);
nand U1313 (N_1313,N_699,N_745);
or U1314 (N_1314,N_523,N_724);
or U1315 (N_1315,N_604,N_983);
nor U1316 (N_1316,N_812,N_654);
or U1317 (N_1317,N_613,N_721);
and U1318 (N_1318,N_854,N_687);
nand U1319 (N_1319,N_855,N_501);
and U1320 (N_1320,N_777,N_924);
and U1321 (N_1321,N_910,N_695);
nor U1322 (N_1322,N_618,N_562);
or U1323 (N_1323,N_976,N_909);
nand U1324 (N_1324,N_976,N_997);
or U1325 (N_1325,N_567,N_809);
and U1326 (N_1326,N_897,N_993);
and U1327 (N_1327,N_993,N_510);
nor U1328 (N_1328,N_856,N_589);
nor U1329 (N_1329,N_803,N_761);
and U1330 (N_1330,N_958,N_859);
nor U1331 (N_1331,N_995,N_912);
nor U1332 (N_1332,N_712,N_530);
nor U1333 (N_1333,N_830,N_740);
nand U1334 (N_1334,N_597,N_559);
nand U1335 (N_1335,N_668,N_911);
nand U1336 (N_1336,N_518,N_575);
and U1337 (N_1337,N_811,N_658);
nand U1338 (N_1338,N_526,N_500);
and U1339 (N_1339,N_598,N_589);
or U1340 (N_1340,N_870,N_527);
or U1341 (N_1341,N_832,N_753);
nor U1342 (N_1342,N_864,N_595);
or U1343 (N_1343,N_721,N_816);
nor U1344 (N_1344,N_823,N_575);
nand U1345 (N_1345,N_576,N_530);
and U1346 (N_1346,N_838,N_692);
or U1347 (N_1347,N_662,N_632);
nor U1348 (N_1348,N_799,N_632);
nor U1349 (N_1349,N_854,N_540);
or U1350 (N_1350,N_736,N_677);
nand U1351 (N_1351,N_916,N_612);
and U1352 (N_1352,N_887,N_938);
nand U1353 (N_1353,N_520,N_706);
and U1354 (N_1354,N_831,N_575);
nand U1355 (N_1355,N_579,N_604);
nor U1356 (N_1356,N_765,N_818);
or U1357 (N_1357,N_726,N_968);
nand U1358 (N_1358,N_823,N_520);
nor U1359 (N_1359,N_565,N_562);
nand U1360 (N_1360,N_768,N_907);
or U1361 (N_1361,N_810,N_612);
nor U1362 (N_1362,N_861,N_609);
or U1363 (N_1363,N_740,N_913);
or U1364 (N_1364,N_964,N_950);
nor U1365 (N_1365,N_993,N_536);
nor U1366 (N_1366,N_687,N_684);
or U1367 (N_1367,N_599,N_597);
or U1368 (N_1368,N_830,N_744);
nand U1369 (N_1369,N_758,N_574);
nand U1370 (N_1370,N_726,N_508);
nor U1371 (N_1371,N_915,N_704);
nand U1372 (N_1372,N_934,N_571);
or U1373 (N_1373,N_893,N_936);
and U1374 (N_1374,N_913,N_969);
nor U1375 (N_1375,N_721,N_978);
and U1376 (N_1376,N_546,N_782);
nor U1377 (N_1377,N_862,N_558);
nand U1378 (N_1378,N_968,N_742);
nor U1379 (N_1379,N_674,N_549);
and U1380 (N_1380,N_592,N_743);
nor U1381 (N_1381,N_718,N_564);
and U1382 (N_1382,N_930,N_533);
and U1383 (N_1383,N_680,N_895);
and U1384 (N_1384,N_516,N_930);
or U1385 (N_1385,N_936,N_664);
or U1386 (N_1386,N_522,N_878);
and U1387 (N_1387,N_717,N_877);
nor U1388 (N_1388,N_743,N_792);
or U1389 (N_1389,N_745,N_951);
or U1390 (N_1390,N_987,N_698);
nand U1391 (N_1391,N_621,N_643);
nor U1392 (N_1392,N_723,N_702);
nand U1393 (N_1393,N_945,N_621);
nor U1394 (N_1394,N_699,N_569);
nor U1395 (N_1395,N_998,N_562);
and U1396 (N_1396,N_519,N_514);
or U1397 (N_1397,N_813,N_948);
nand U1398 (N_1398,N_685,N_544);
nand U1399 (N_1399,N_725,N_938);
or U1400 (N_1400,N_787,N_518);
and U1401 (N_1401,N_853,N_767);
and U1402 (N_1402,N_886,N_705);
or U1403 (N_1403,N_779,N_960);
nor U1404 (N_1404,N_820,N_733);
nand U1405 (N_1405,N_672,N_851);
nor U1406 (N_1406,N_936,N_600);
and U1407 (N_1407,N_688,N_570);
and U1408 (N_1408,N_778,N_645);
nand U1409 (N_1409,N_568,N_598);
nor U1410 (N_1410,N_909,N_533);
nand U1411 (N_1411,N_650,N_844);
nor U1412 (N_1412,N_817,N_610);
nand U1413 (N_1413,N_549,N_542);
and U1414 (N_1414,N_594,N_844);
or U1415 (N_1415,N_705,N_593);
or U1416 (N_1416,N_750,N_754);
nand U1417 (N_1417,N_599,N_989);
nor U1418 (N_1418,N_865,N_800);
and U1419 (N_1419,N_800,N_628);
nand U1420 (N_1420,N_891,N_786);
or U1421 (N_1421,N_696,N_953);
or U1422 (N_1422,N_800,N_670);
nand U1423 (N_1423,N_673,N_988);
and U1424 (N_1424,N_730,N_609);
xnor U1425 (N_1425,N_505,N_552);
nor U1426 (N_1426,N_995,N_696);
nand U1427 (N_1427,N_976,N_792);
and U1428 (N_1428,N_803,N_665);
and U1429 (N_1429,N_913,N_885);
nand U1430 (N_1430,N_571,N_999);
nand U1431 (N_1431,N_922,N_981);
nand U1432 (N_1432,N_522,N_835);
xnor U1433 (N_1433,N_999,N_852);
and U1434 (N_1434,N_695,N_729);
nor U1435 (N_1435,N_996,N_551);
nand U1436 (N_1436,N_638,N_879);
or U1437 (N_1437,N_881,N_508);
nor U1438 (N_1438,N_925,N_784);
nor U1439 (N_1439,N_891,N_689);
nand U1440 (N_1440,N_891,N_751);
nor U1441 (N_1441,N_978,N_638);
or U1442 (N_1442,N_935,N_659);
nand U1443 (N_1443,N_625,N_845);
nand U1444 (N_1444,N_652,N_819);
nor U1445 (N_1445,N_774,N_781);
or U1446 (N_1446,N_541,N_814);
or U1447 (N_1447,N_857,N_568);
and U1448 (N_1448,N_832,N_721);
nand U1449 (N_1449,N_556,N_627);
and U1450 (N_1450,N_878,N_654);
nand U1451 (N_1451,N_918,N_961);
nand U1452 (N_1452,N_669,N_681);
and U1453 (N_1453,N_656,N_577);
nor U1454 (N_1454,N_557,N_776);
or U1455 (N_1455,N_858,N_661);
or U1456 (N_1456,N_680,N_852);
nand U1457 (N_1457,N_732,N_886);
nand U1458 (N_1458,N_530,N_517);
and U1459 (N_1459,N_892,N_561);
or U1460 (N_1460,N_624,N_584);
nand U1461 (N_1461,N_557,N_658);
nand U1462 (N_1462,N_901,N_766);
nor U1463 (N_1463,N_869,N_924);
and U1464 (N_1464,N_987,N_523);
or U1465 (N_1465,N_941,N_836);
or U1466 (N_1466,N_560,N_673);
or U1467 (N_1467,N_819,N_763);
xor U1468 (N_1468,N_905,N_876);
nand U1469 (N_1469,N_775,N_629);
and U1470 (N_1470,N_948,N_535);
and U1471 (N_1471,N_940,N_908);
nand U1472 (N_1472,N_779,N_931);
nor U1473 (N_1473,N_751,N_954);
nand U1474 (N_1474,N_752,N_525);
nand U1475 (N_1475,N_670,N_993);
nand U1476 (N_1476,N_783,N_665);
nand U1477 (N_1477,N_570,N_738);
nand U1478 (N_1478,N_665,N_874);
nand U1479 (N_1479,N_611,N_683);
or U1480 (N_1480,N_552,N_610);
nand U1481 (N_1481,N_899,N_667);
nor U1482 (N_1482,N_762,N_619);
or U1483 (N_1483,N_572,N_927);
nor U1484 (N_1484,N_744,N_856);
or U1485 (N_1485,N_793,N_533);
nor U1486 (N_1486,N_508,N_612);
nor U1487 (N_1487,N_837,N_822);
nor U1488 (N_1488,N_893,N_876);
nor U1489 (N_1489,N_823,N_798);
nand U1490 (N_1490,N_705,N_507);
or U1491 (N_1491,N_845,N_541);
nand U1492 (N_1492,N_651,N_863);
nand U1493 (N_1493,N_816,N_943);
nor U1494 (N_1494,N_820,N_663);
and U1495 (N_1495,N_708,N_794);
or U1496 (N_1496,N_879,N_741);
nor U1497 (N_1497,N_931,N_578);
and U1498 (N_1498,N_944,N_517);
nor U1499 (N_1499,N_756,N_599);
nor U1500 (N_1500,N_1324,N_1011);
nand U1501 (N_1501,N_1079,N_1026);
and U1502 (N_1502,N_1498,N_1341);
nand U1503 (N_1503,N_1226,N_1097);
nand U1504 (N_1504,N_1189,N_1092);
nor U1505 (N_1505,N_1423,N_1383);
or U1506 (N_1506,N_1493,N_1233);
nor U1507 (N_1507,N_1147,N_1497);
nor U1508 (N_1508,N_1457,N_1081);
and U1509 (N_1509,N_1474,N_1204);
nand U1510 (N_1510,N_1289,N_1365);
nand U1511 (N_1511,N_1452,N_1330);
nand U1512 (N_1512,N_1184,N_1394);
and U1513 (N_1513,N_1308,N_1279);
nand U1514 (N_1514,N_1076,N_1054);
nor U1515 (N_1515,N_1294,N_1481);
and U1516 (N_1516,N_1491,N_1486);
or U1517 (N_1517,N_1302,N_1379);
xnor U1518 (N_1518,N_1166,N_1133);
nand U1519 (N_1519,N_1215,N_1203);
and U1520 (N_1520,N_1047,N_1187);
or U1521 (N_1521,N_1409,N_1216);
nand U1522 (N_1522,N_1313,N_1051);
or U1523 (N_1523,N_1311,N_1208);
and U1524 (N_1524,N_1415,N_1299);
and U1525 (N_1525,N_1209,N_1471);
nor U1526 (N_1526,N_1362,N_1263);
nand U1527 (N_1527,N_1321,N_1101);
or U1528 (N_1528,N_1250,N_1327);
nand U1529 (N_1529,N_1165,N_1141);
nor U1530 (N_1530,N_1041,N_1361);
nor U1531 (N_1531,N_1462,N_1314);
and U1532 (N_1532,N_1085,N_1373);
nand U1533 (N_1533,N_1036,N_1134);
or U1534 (N_1534,N_1420,N_1170);
or U1535 (N_1535,N_1459,N_1048);
and U1536 (N_1536,N_1214,N_1149);
and U1537 (N_1537,N_1103,N_1439);
or U1538 (N_1538,N_1364,N_1091);
and U1539 (N_1539,N_1089,N_1447);
and U1540 (N_1540,N_1344,N_1372);
or U1541 (N_1541,N_1159,N_1231);
and U1542 (N_1542,N_1205,N_1237);
nand U1543 (N_1543,N_1405,N_1354);
nand U1544 (N_1544,N_1242,N_1432);
nand U1545 (N_1545,N_1375,N_1006);
nor U1546 (N_1546,N_1320,N_1297);
or U1547 (N_1547,N_1228,N_1106);
or U1548 (N_1548,N_1012,N_1470);
or U1549 (N_1549,N_1254,N_1136);
or U1550 (N_1550,N_1014,N_1118);
nand U1551 (N_1551,N_1368,N_1438);
and U1552 (N_1552,N_1400,N_1013);
nand U1553 (N_1553,N_1169,N_1171);
nor U1554 (N_1554,N_1355,N_1251);
nand U1555 (N_1555,N_1393,N_1199);
or U1556 (N_1556,N_1333,N_1010);
or U1557 (N_1557,N_1062,N_1325);
and U1558 (N_1558,N_1061,N_1290);
nor U1559 (N_1559,N_1413,N_1306);
and U1560 (N_1560,N_1175,N_1040);
nand U1561 (N_1561,N_1119,N_1286);
or U1562 (N_1562,N_1059,N_1315);
nor U1563 (N_1563,N_1109,N_1283);
nand U1564 (N_1564,N_1449,N_1053);
and U1565 (N_1565,N_1016,N_1145);
or U1566 (N_1566,N_1454,N_1069);
or U1567 (N_1567,N_1024,N_1173);
or U1568 (N_1568,N_1261,N_1066);
or U1569 (N_1569,N_1367,N_1282);
nor U1570 (N_1570,N_1125,N_1273);
nand U1571 (N_1571,N_1213,N_1406);
nor U1572 (N_1572,N_1156,N_1262);
or U1573 (N_1573,N_1358,N_1023);
nand U1574 (N_1574,N_1494,N_1356);
and U1575 (N_1575,N_1220,N_1412);
nor U1576 (N_1576,N_1198,N_1331);
nor U1577 (N_1577,N_1402,N_1437);
nor U1578 (N_1578,N_1359,N_1377);
nor U1579 (N_1579,N_1063,N_1143);
or U1580 (N_1580,N_1392,N_1129);
or U1581 (N_1581,N_1241,N_1150);
and U1582 (N_1582,N_1426,N_1046);
and U1583 (N_1583,N_1245,N_1458);
nand U1584 (N_1584,N_1374,N_1223);
nor U1585 (N_1585,N_1234,N_1080);
nor U1586 (N_1586,N_1366,N_1138);
and U1587 (N_1587,N_1192,N_1293);
and U1588 (N_1588,N_1280,N_1335);
nand U1589 (N_1589,N_1148,N_1068);
and U1590 (N_1590,N_1422,N_1492);
nor U1591 (N_1591,N_1489,N_1072);
and U1592 (N_1592,N_1487,N_1064);
and U1593 (N_1593,N_1132,N_1248);
nand U1594 (N_1594,N_1028,N_1116);
or U1595 (N_1595,N_1408,N_1135);
or U1596 (N_1596,N_1466,N_1395);
xor U1597 (N_1597,N_1269,N_1194);
nand U1598 (N_1598,N_1317,N_1312);
nor U1599 (N_1599,N_1259,N_1021);
or U1600 (N_1600,N_1476,N_1083);
and U1601 (N_1601,N_1146,N_1099);
xor U1602 (N_1602,N_1300,N_1182);
nand U1603 (N_1603,N_1378,N_1418);
or U1604 (N_1604,N_1456,N_1433);
or U1605 (N_1605,N_1117,N_1084);
and U1606 (N_1606,N_1285,N_1446);
nand U1607 (N_1607,N_1104,N_1403);
nor U1608 (N_1608,N_1045,N_1060);
and U1609 (N_1609,N_1202,N_1472);
xnor U1610 (N_1610,N_1167,N_1464);
nand U1611 (N_1611,N_1448,N_1020);
nand U1612 (N_1612,N_1193,N_1275);
nand U1613 (N_1613,N_1332,N_1381);
and U1614 (N_1614,N_1292,N_1496);
and U1615 (N_1615,N_1347,N_1086);
nand U1616 (N_1616,N_1266,N_1111);
nor U1617 (N_1617,N_1094,N_1218);
nand U1618 (N_1618,N_1391,N_1130);
nor U1619 (N_1619,N_1239,N_1281);
nor U1620 (N_1620,N_1307,N_1442);
and U1621 (N_1621,N_1077,N_1428);
xnor U1622 (N_1622,N_1087,N_1318);
or U1623 (N_1623,N_1178,N_1288);
or U1624 (N_1624,N_1495,N_1398);
nand U1625 (N_1625,N_1009,N_1386);
nor U1626 (N_1626,N_1272,N_1304);
nand U1627 (N_1627,N_1396,N_1485);
and U1628 (N_1628,N_1219,N_1029);
nor U1629 (N_1629,N_1181,N_1253);
and U1630 (N_1630,N_1033,N_1336);
nor U1631 (N_1631,N_1258,N_1227);
and U1632 (N_1632,N_1276,N_1058);
nand U1633 (N_1633,N_1157,N_1278);
and U1634 (N_1634,N_1477,N_1206);
or U1635 (N_1635,N_1034,N_1343);
or U1636 (N_1636,N_1360,N_1049);
nor U1637 (N_1637,N_1349,N_1287);
and U1638 (N_1638,N_1455,N_1351);
and U1639 (N_1639,N_1108,N_1031);
nor U1640 (N_1640,N_1211,N_1329);
nand U1641 (N_1641,N_1430,N_1007);
nor U1642 (N_1642,N_1404,N_1088);
nor U1643 (N_1643,N_1107,N_1399);
or U1644 (N_1644,N_1376,N_1389);
or U1645 (N_1645,N_1483,N_1144);
xor U1646 (N_1646,N_1110,N_1093);
and U1647 (N_1647,N_1003,N_1467);
or U1648 (N_1648,N_1124,N_1270);
nand U1649 (N_1649,N_1480,N_1340);
nor U1650 (N_1650,N_1015,N_1431);
nand U1651 (N_1651,N_1073,N_1411);
or U1652 (N_1652,N_1112,N_1390);
nand U1653 (N_1653,N_1309,N_1421);
or U1654 (N_1654,N_1388,N_1161);
nand U1655 (N_1655,N_1095,N_1443);
or U1656 (N_1656,N_1338,N_1139);
nand U1657 (N_1657,N_1291,N_1074);
nor U1658 (N_1658,N_1055,N_1441);
and U1659 (N_1659,N_1328,N_1256);
nand U1660 (N_1660,N_1191,N_1429);
and U1661 (N_1661,N_1098,N_1078);
nor U1662 (N_1662,N_1222,N_1350);
nand U1663 (N_1663,N_1484,N_1043);
nand U1664 (N_1664,N_1005,N_1252);
or U1665 (N_1665,N_1353,N_1018);
and U1666 (N_1666,N_1255,N_1153);
or U1667 (N_1667,N_1468,N_1035);
nor U1668 (N_1668,N_1186,N_1337);
and U1669 (N_1669,N_1499,N_1444);
and U1670 (N_1670,N_1339,N_1382);
and U1671 (N_1671,N_1075,N_1195);
nand U1672 (N_1672,N_1052,N_1001);
nor U1673 (N_1673,N_1478,N_1152);
nand U1674 (N_1674,N_1039,N_1142);
or U1675 (N_1675,N_1128,N_1475);
nor U1676 (N_1676,N_1316,N_1229);
nand U1677 (N_1677,N_1345,N_1235);
and U1678 (N_1678,N_1200,N_1380);
nand U1679 (N_1679,N_1407,N_1419);
or U1680 (N_1680,N_1310,N_1154);
nor U1681 (N_1681,N_1174,N_1185);
and U1682 (N_1682,N_1436,N_1158);
nand U1683 (N_1683,N_1162,N_1196);
and U1684 (N_1684,N_1183,N_1131);
and U1685 (N_1685,N_1440,N_1461);
nor U1686 (N_1686,N_1180,N_1303);
nor U1687 (N_1687,N_1071,N_1115);
nor U1688 (N_1688,N_1277,N_1424);
nor U1689 (N_1689,N_1022,N_1151);
nand U1690 (N_1690,N_1473,N_1267);
or U1691 (N_1691,N_1463,N_1322);
and U1692 (N_1692,N_1232,N_1264);
nand U1693 (N_1693,N_1168,N_1105);
and U1694 (N_1694,N_1257,N_1244);
and U1695 (N_1695,N_1469,N_1247);
or U1696 (N_1696,N_1217,N_1102);
nand U1697 (N_1697,N_1387,N_1295);
or U1698 (N_1698,N_1427,N_1038);
nand U1699 (N_1699,N_1070,N_1008);
or U1700 (N_1700,N_1246,N_1271);
nor U1701 (N_1701,N_1027,N_1460);
nor U1702 (N_1702,N_1342,N_1201);
nand U1703 (N_1703,N_1348,N_1369);
xor U1704 (N_1704,N_1179,N_1163);
nand U1705 (N_1705,N_1030,N_1090);
nor U1706 (N_1706,N_1249,N_1450);
nor U1707 (N_1707,N_1260,N_1114);
nor U1708 (N_1708,N_1384,N_1044);
nand U1709 (N_1709,N_1298,N_1479);
or U1710 (N_1710,N_1453,N_1268);
and U1711 (N_1711,N_1434,N_1352);
nor U1712 (N_1712,N_1296,N_1056);
nand U1713 (N_1713,N_1000,N_1207);
nor U1714 (N_1714,N_1140,N_1451);
or U1715 (N_1715,N_1127,N_1197);
nand U1716 (N_1716,N_1224,N_1371);
nor U1717 (N_1717,N_1490,N_1172);
nor U1718 (N_1718,N_1274,N_1236);
nand U1719 (N_1719,N_1401,N_1160);
and U1720 (N_1720,N_1319,N_1212);
and U1721 (N_1721,N_1017,N_1037);
nor U1722 (N_1722,N_1177,N_1370);
and U1723 (N_1723,N_1334,N_1155);
or U1724 (N_1724,N_1425,N_1410);
and U1725 (N_1725,N_1230,N_1238);
nor U1726 (N_1726,N_1385,N_1284);
nor U1727 (N_1727,N_1445,N_1465);
nand U1728 (N_1728,N_1397,N_1096);
nor U1729 (N_1729,N_1100,N_1210);
nand U1730 (N_1730,N_1126,N_1488);
and U1731 (N_1731,N_1057,N_1363);
nand U1732 (N_1732,N_1225,N_1221);
nor U1733 (N_1733,N_1042,N_1032);
nor U1734 (N_1734,N_1326,N_1305);
and U1735 (N_1735,N_1082,N_1414);
or U1736 (N_1736,N_1019,N_1482);
or U1737 (N_1737,N_1164,N_1121);
nand U1738 (N_1738,N_1190,N_1065);
nand U1739 (N_1739,N_1357,N_1323);
and U1740 (N_1740,N_1435,N_1002);
and U1741 (N_1741,N_1050,N_1265);
and U1742 (N_1742,N_1067,N_1137);
and U1743 (N_1743,N_1123,N_1113);
nand U1744 (N_1744,N_1004,N_1025);
nand U1745 (N_1745,N_1301,N_1416);
nor U1746 (N_1746,N_1176,N_1188);
and U1747 (N_1747,N_1417,N_1240);
or U1748 (N_1748,N_1346,N_1120);
or U1749 (N_1749,N_1122,N_1243);
nand U1750 (N_1750,N_1359,N_1179);
and U1751 (N_1751,N_1481,N_1352);
or U1752 (N_1752,N_1488,N_1204);
nor U1753 (N_1753,N_1047,N_1366);
or U1754 (N_1754,N_1330,N_1010);
nor U1755 (N_1755,N_1280,N_1167);
and U1756 (N_1756,N_1192,N_1099);
nand U1757 (N_1757,N_1416,N_1264);
and U1758 (N_1758,N_1282,N_1193);
and U1759 (N_1759,N_1094,N_1204);
nor U1760 (N_1760,N_1111,N_1497);
and U1761 (N_1761,N_1245,N_1252);
and U1762 (N_1762,N_1387,N_1089);
and U1763 (N_1763,N_1039,N_1224);
or U1764 (N_1764,N_1253,N_1411);
nand U1765 (N_1765,N_1366,N_1349);
and U1766 (N_1766,N_1091,N_1411);
and U1767 (N_1767,N_1080,N_1438);
nor U1768 (N_1768,N_1487,N_1499);
nor U1769 (N_1769,N_1137,N_1454);
or U1770 (N_1770,N_1325,N_1117);
or U1771 (N_1771,N_1126,N_1193);
or U1772 (N_1772,N_1401,N_1225);
nand U1773 (N_1773,N_1476,N_1123);
and U1774 (N_1774,N_1088,N_1097);
nand U1775 (N_1775,N_1079,N_1261);
nand U1776 (N_1776,N_1282,N_1085);
or U1777 (N_1777,N_1177,N_1110);
and U1778 (N_1778,N_1418,N_1231);
and U1779 (N_1779,N_1179,N_1263);
and U1780 (N_1780,N_1334,N_1183);
and U1781 (N_1781,N_1193,N_1380);
or U1782 (N_1782,N_1138,N_1106);
or U1783 (N_1783,N_1401,N_1366);
nor U1784 (N_1784,N_1496,N_1296);
nand U1785 (N_1785,N_1022,N_1003);
and U1786 (N_1786,N_1459,N_1120);
or U1787 (N_1787,N_1139,N_1275);
nand U1788 (N_1788,N_1276,N_1454);
and U1789 (N_1789,N_1186,N_1220);
nor U1790 (N_1790,N_1491,N_1110);
or U1791 (N_1791,N_1224,N_1466);
or U1792 (N_1792,N_1274,N_1207);
nand U1793 (N_1793,N_1414,N_1353);
or U1794 (N_1794,N_1440,N_1251);
or U1795 (N_1795,N_1173,N_1373);
nor U1796 (N_1796,N_1172,N_1124);
and U1797 (N_1797,N_1352,N_1424);
and U1798 (N_1798,N_1287,N_1175);
nor U1799 (N_1799,N_1306,N_1137);
nand U1800 (N_1800,N_1017,N_1173);
or U1801 (N_1801,N_1064,N_1375);
or U1802 (N_1802,N_1219,N_1308);
and U1803 (N_1803,N_1070,N_1195);
nor U1804 (N_1804,N_1492,N_1057);
and U1805 (N_1805,N_1092,N_1016);
nand U1806 (N_1806,N_1054,N_1079);
and U1807 (N_1807,N_1486,N_1384);
or U1808 (N_1808,N_1300,N_1228);
nand U1809 (N_1809,N_1232,N_1251);
nand U1810 (N_1810,N_1473,N_1356);
and U1811 (N_1811,N_1022,N_1158);
or U1812 (N_1812,N_1365,N_1267);
or U1813 (N_1813,N_1410,N_1336);
and U1814 (N_1814,N_1439,N_1493);
nand U1815 (N_1815,N_1078,N_1158);
nor U1816 (N_1816,N_1479,N_1263);
nor U1817 (N_1817,N_1379,N_1234);
nand U1818 (N_1818,N_1148,N_1446);
nor U1819 (N_1819,N_1457,N_1253);
and U1820 (N_1820,N_1120,N_1172);
nor U1821 (N_1821,N_1295,N_1489);
nand U1822 (N_1822,N_1305,N_1422);
nor U1823 (N_1823,N_1490,N_1275);
or U1824 (N_1824,N_1044,N_1434);
nor U1825 (N_1825,N_1100,N_1339);
nand U1826 (N_1826,N_1436,N_1267);
and U1827 (N_1827,N_1225,N_1108);
and U1828 (N_1828,N_1460,N_1190);
nand U1829 (N_1829,N_1448,N_1470);
nor U1830 (N_1830,N_1044,N_1168);
nor U1831 (N_1831,N_1358,N_1011);
or U1832 (N_1832,N_1294,N_1118);
nand U1833 (N_1833,N_1289,N_1277);
and U1834 (N_1834,N_1263,N_1406);
and U1835 (N_1835,N_1429,N_1384);
or U1836 (N_1836,N_1412,N_1073);
and U1837 (N_1837,N_1168,N_1137);
or U1838 (N_1838,N_1149,N_1221);
xor U1839 (N_1839,N_1227,N_1179);
nand U1840 (N_1840,N_1102,N_1174);
nor U1841 (N_1841,N_1353,N_1331);
nand U1842 (N_1842,N_1210,N_1156);
and U1843 (N_1843,N_1314,N_1060);
nor U1844 (N_1844,N_1131,N_1008);
nor U1845 (N_1845,N_1186,N_1322);
or U1846 (N_1846,N_1141,N_1059);
nand U1847 (N_1847,N_1426,N_1215);
nor U1848 (N_1848,N_1219,N_1422);
or U1849 (N_1849,N_1148,N_1338);
nor U1850 (N_1850,N_1016,N_1380);
and U1851 (N_1851,N_1348,N_1233);
nor U1852 (N_1852,N_1378,N_1399);
or U1853 (N_1853,N_1228,N_1254);
and U1854 (N_1854,N_1326,N_1020);
and U1855 (N_1855,N_1120,N_1355);
and U1856 (N_1856,N_1001,N_1012);
and U1857 (N_1857,N_1378,N_1483);
nor U1858 (N_1858,N_1226,N_1092);
or U1859 (N_1859,N_1007,N_1407);
or U1860 (N_1860,N_1397,N_1245);
nor U1861 (N_1861,N_1372,N_1158);
nor U1862 (N_1862,N_1022,N_1469);
or U1863 (N_1863,N_1360,N_1034);
nor U1864 (N_1864,N_1298,N_1339);
or U1865 (N_1865,N_1290,N_1404);
or U1866 (N_1866,N_1324,N_1419);
xor U1867 (N_1867,N_1277,N_1335);
or U1868 (N_1868,N_1194,N_1264);
nand U1869 (N_1869,N_1429,N_1055);
nor U1870 (N_1870,N_1012,N_1302);
nor U1871 (N_1871,N_1015,N_1254);
or U1872 (N_1872,N_1399,N_1270);
or U1873 (N_1873,N_1054,N_1300);
nor U1874 (N_1874,N_1098,N_1290);
nand U1875 (N_1875,N_1269,N_1399);
nand U1876 (N_1876,N_1170,N_1202);
nand U1877 (N_1877,N_1485,N_1132);
or U1878 (N_1878,N_1333,N_1167);
and U1879 (N_1879,N_1008,N_1071);
nor U1880 (N_1880,N_1384,N_1382);
nand U1881 (N_1881,N_1100,N_1466);
and U1882 (N_1882,N_1091,N_1398);
nand U1883 (N_1883,N_1280,N_1131);
or U1884 (N_1884,N_1209,N_1412);
nor U1885 (N_1885,N_1494,N_1297);
nor U1886 (N_1886,N_1323,N_1215);
nor U1887 (N_1887,N_1358,N_1436);
nand U1888 (N_1888,N_1108,N_1006);
nor U1889 (N_1889,N_1438,N_1482);
xnor U1890 (N_1890,N_1466,N_1139);
nor U1891 (N_1891,N_1361,N_1349);
and U1892 (N_1892,N_1023,N_1105);
or U1893 (N_1893,N_1373,N_1349);
or U1894 (N_1894,N_1488,N_1290);
or U1895 (N_1895,N_1307,N_1363);
nor U1896 (N_1896,N_1184,N_1191);
nor U1897 (N_1897,N_1051,N_1237);
nand U1898 (N_1898,N_1349,N_1089);
xnor U1899 (N_1899,N_1369,N_1210);
and U1900 (N_1900,N_1352,N_1201);
or U1901 (N_1901,N_1396,N_1117);
nand U1902 (N_1902,N_1193,N_1175);
nand U1903 (N_1903,N_1318,N_1089);
and U1904 (N_1904,N_1189,N_1167);
nand U1905 (N_1905,N_1365,N_1410);
nor U1906 (N_1906,N_1462,N_1476);
nand U1907 (N_1907,N_1378,N_1459);
and U1908 (N_1908,N_1101,N_1232);
or U1909 (N_1909,N_1389,N_1232);
and U1910 (N_1910,N_1233,N_1246);
or U1911 (N_1911,N_1101,N_1465);
and U1912 (N_1912,N_1399,N_1384);
nand U1913 (N_1913,N_1434,N_1423);
or U1914 (N_1914,N_1387,N_1175);
nor U1915 (N_1915,N_1200,N_1154);
nor U1916 (N_1916,N_1223,N_1022);
and U1917 (N_1917,N_1498,N_1400);
nand U1918 (N_1918,N_1289,N_1191);
nor U1919 (N_1919,N_1200,N_1241);
nor U1920 (N_1920,N_1068,N_1287);
nor U1921 (N_1921,N_1173,N_1041);
and U1922 (N_1922,N_1272,N_1375);
nand U1923 (N_1923,N_1462,N_1008);
or U1924 (N_1924,N_1449,N_1041);
or U1925 (N_1925,N_1499,N_1408);
nand U1926 (N_1926,N_1026,N_1090);
and U1927 (N_1927,N_1160,N_1395);
nor U1928 (N_1928,N_1304,N_1396);
or U1929 (N_1929,N_1152,N_1482);
and U1930 (N_1930,N_1352,N_1195);
or U1931 (N_1931,N_1293,N_1226);
nand U1932 (N_1932,N_1216,N_1339);
or U1933 (N_1933,N_1181,N_1143);
nor U1934 (N_1934,N_1083,N_1071);
nor U1935 (N_1935,N_1125,N_1167);
and U1936 (N_1936,N_1021,N_1404);
nand U1937 (N_1937,N_1453,N_1155);
and U1938 (N_1938,N_1176,N_1061);
nor U1939 (N_1939,N_1254,N_1482);
and U1940 (N_1940,N_1495,N_1347);
nand U1941 (N_1941,N_1280,N_1139);
nor U1942 (N_1942,N_1282,N_1299);
or U1943 (N_1943,N_1025,N_1267);
nand U1944 (N_1944,N_1081,N_1033);
and U1945 (N_1945,N_1093,N_1165);
and U1946 (N_1946,N_1387,N_1346);
nor U1947 (N_1947,N_1158,N_1288);
and U1948 (N_1948,N_1341,N_1391);
nor U1949 (N_1949,N_1190,N_1011);
and U1950 (N_1950,N_1284,N_1369);
nand U1951 (N_1951,N_1352,N_1381);
or U1952 (N_1952,N_1116,N_1403);
or U1953 (N_1953,N_1478,N_1452);
or U1954 (N_1954,N_1281,N_1053);
or U1955 (N_1955,N_1343,N_1144);
and U1956 (N_1956,N_1304,N_1352);
and U1957 (N_1957,N_1407,N_1210);
and U1958 (N_1958,N_1485,N_1138);
and U1959 (N_1959,N_1265,N_1349);
and U1960 (N_1960,N_1311,N_1293);
and U1961 (N_1961,N_1030,N_1053);
nand U1962 (N_1962,N_1309,N_1142);
or U1963 (N_1963,N_1453,N_1475);
or U1964 (N_1964,N_1065,N_1251);
nand U1965 (N_1965,N_1395,N_1271);
nor U1966 (N_1966,N_1017,N_1440);
or U1967 (N_1967,N_1036,N_1185);
and U1968 (N_1968,N_1167,N_1325);
xnor U1969 (N_1969,N_1476,N_1207);
nor U1970 (N_1970,N_1060,N_1453);
and U1971 (N_1971,N_1433,N_1073);
nor U1972 (N_1972,N_1121,N_1411);
or U1973 (N_1973,N_1046,N_1366);
or U1974 (N_1974,N_1000,N_1026);
and U1975 (N_1975,N_1406,N_1438);
nand U1976 (N_1976,N_1230,N_1222);
and U1977 (N_1977,N_1302,N_1289);
or U1978 (N_1978,N_1456,N_1354);
nand U1979 (N_1979,N_1086,N_1309);
and U1980 (N_1980,N_1103,N_1154);
or U1981 (N_1981,N_1215,N_1080);
nand U1982 (N_1982,N_1073,N_1238);
or U1983 (N_1983,N_1317,N_1192);
nand U1984 (N_1984,N_1356,N_1089);
and U1985 (N_1985,N_1034,N_1465);
nand U1986 (N_1986,N_1476,N_1010);
nor U1987 (N_1987,N_1358,N_1217);
and U1988 (N_1988,N_1372,N_1118);
nand U1989 (N_1989,N_1244,N_1462);
nor U1990 (N_1990,N_1433,N_1358);
or U1991 (N_1991,N_1407,N_1163);
nor U1992 (N_1992,N_1179,N_1157);
and U1993 (N_1993,N_1288,N_1066);
or U1994 (N_1994,N_1227,N_1184);
nand U1995 (N_1995,N_1294,N_1077);
nand U1996 (N_1996,N_1441,N_1451);
nand U1997 (N_1997,N_1492,N_1168);
and U1998 (N_1998,N_1183,N_1056);
nor U1999 (N_1999,N_1333,N_1016);
and U2000 (N_2000,N_1764,N_1646);
or U2001 (N_2001,N_1977,N_1962);
nor U2002 (N_2002,N_1789,N_1701);
and U2003 (N_2003,N_1557,N_1520);
nor U2004 (N_2004,N_1842,N_1569);
nor U2005 (N_2005,N_1617,N_1503);
and U2006 (N_2006,N_1758,N_1887);
and U2007 (N_2007,N_1637,N_1865);
or U2008 (N_2008,N_1753,N_1636);
and U2009 (N_2009,N_1559,N_1814);
nand U2010 (N_2010,N_1872,N_1524);
or U2011 (N_2011,N_1800,N_1951);
or U2012 (N_2012,N_1712,N_1914);
nand U2013 (N_2013,N_1711,N_1666);
nor U2014 (N_2014,N_1660,N_1526);
and U2015 (N_2015,N_1974,N_1732);
nor U2016 (N_2016,N_1669,N_1912);
nor U2017 (N_2017,N_1766,N_1851);
xnor U2018 (N_2018,N_1863,N_1548);
or U2019 (N_2019,N_1762,N_1978);
nand U2020 (N_2020,N_1692,N_1835);
nand U2021 (N_2021,N_1932,N_1791);
nor U2022 (N_2022,N_1650,N_1558);
and U2023 (N_2023,N_1573,N_1964);
and U2024 (N_2024,N_1609,N_1828);
nand U2025 (N_2025,N_1723,N_1922);
nand U2026 (N_2026,N_1936,N_1952);
and U2027 (N_2027,N_1947,N_1570);
and U2028 (N_2028,N_1769,N_1605);
and U2029 (N_2029,N_1856,N_1787);
nand U2030 (N_2030,N_1598,N_1901);
nand U2031 (N_2031,N_1981,N_1755);
or U2032 (N_2032,N_1907,N_1565);
or U2033 (N_2033,N_1987,N_1906);
nand U2034 (N_2034,N_1674,N_1709);
and U2035 (N_2035,N_1943,N_1999);
nand U2036 (N_2036,N_1904,N_1895);
or U2037 (N_2037,N_1748,N_1546);
and U2038 (N_2038,N_1514,N_1919);
or U2039 (N_2039,N_1774,N_1556);
nor U2040 (N_2040,N_1809,N_1903);
and U2041 (N_2041,N_1622,N_1626);
and U2042 (N_2042,N_1663,N_1632);
and U2043 (N_2043,N_1505,N_1840);
or U2044 (N_2044,N_1536,N_1765);
and U2045 (N_2045,N_1855,N_1533);
nand U2046 (N_2046,N_1615,N_1795);
and U2047 (N_2047,N_1593,N_1928);
nand U2048 (N_2048,N_1591,N_1985);
or U2049 (N_2049,N_1600,N_1816);
nor U2050 (N_2050,N_1576,N_1584);
or U2051 (N_2051,N_1727,N_1850);
and U2052 (N_2052,N_1799,N_1881);
and U2053 (N_2053,N_1549,N_1721);
nor U2054 (N_2054,N_1679,N_1956);
and U2055 (N_2055,N_1635,N_1624);
or U2056 (N_2056,N_1511,N_1859);
and U2057 (N_2057,N_1619,N_1934);
nor U2058 (N_2058,N_1807,N_1633);
nor U2059 (N_2059,N_1797,N_1757);
and U2060 (N_2060,N_1921,N_1606);
nor U2061 (N_2061,N_1671,N_1992);
or U2062 (N_2062,N_1740,N_1927);
nand U2063 (N_2063,N_1829,N_1942);
or U2064 (N_2064,N_1501,N_1811);
nor U2065 (N_2065,N_1984,N_1849);
or U2066 (N_2066,N_1862,N_1661);
nand U2067 (N_2067,N_1995,N_1880);
or U2068 (N_2068,N_1886,N_1720);
nor U2069 (N_2069,N_1547,N_1518);
nor U2070 (N_2070,N_1885,N_1819);
or U2071 (N_2071,N_1909,N_1568);
nor U2072 (N_2072,N_1954,N_1513);
nor U2073 (N_2073,N_1715,N_1967);
nor U2074 (N_2074,N_1644,N_1935);
and U2075 (N_2075,N_1640,N_1852);
nand U2076 (N_2076,N_1698,N_1733);
or U2077 (N_2077,N_1993,N_1686);
nand U2078 (N_2078,N_1543,N_1877);
and U2079 (N_2079,N_1542,N_1902);
and U2080 (N_2080,N_1680,N_1878);
nor U2081 (N_2081,N_1986,N_1836);
or U2082 (N_2082,N_1890,N_1752);
nor U2083 (N_2083,N_1823,N_1554);
and U2084 (N_2084,N_1508,N_1714);
nor U2085 (N_2085,N_1776,N_1638);
or U2086 (N_2086,N_1868,N_1794);
nor U2087 (N_2087,N_1920,N_1681);
nor U2088 (N_2088,N_1938,N_1695);
nor U2089 (N_2089,N_1631,N_1704);
and U2090 (N_2090,N_1911,N_1824);
or U2091 (N_2091,N_1676,N_1623);
nand U2092 (N_2092,N_1893,N_1832);
or U2093 (N_2093,N_1930,N_1580);
and U2094 (N_2094,N_1519,N_1566);
and U2095 (N_2095,N_1949,N_1678);
or U2096 (N_2096,N_1759,N_1627);
nor U2097 (N_2097,N_1529,N_1905);
or U2098 (N_2098,N_1792,N_1899);
and U2099 (N_2099,N_1785,N_1687);
and U2100 (N_2100,N_1782,N_1694);
nor U2101 (N_2101,N_1725,N_1804);
or U2102 (N_2102,N_1882,N_1929);
or U2103 (N_2103,N_1971,N_1892);
nor U2104 (N_2104,N_1729,N_1708);
and U2105 (N_2105,N_1801,N_1963);
nand U2106 (N_2106,N_1634,N_1983);
nor U2107 (N_2107,N_1749,N_1768);
and U2108 (N_2108,N_1628,N_1970);
nand U2109 (N_2109,N_1817,N_1608);
nand U2110 (N_2110,N_1530,N_1771);
and U2111 (N_2111,N_1826,N_1846);
nor U2112 (N_2112,N_1891,N_1563);
or U2113 (N_2113,N_1810,N_1702);
or U2114 (N_2114,N_1586,N_1916);
or U2115 (N_2115,N_1577,N_1643);
and U2116 (N_2116,N_1923,N_1652);
nor U2117 (N_2117,N_1958,N_1957);
and U2118 (N_2118,N_1675,N_1838);
or U2119 (N_2119,N_1837,N_1629);
and U2120 (N_2120,N_1754,N_1802);
nor U2121 (N_2121,N_1502,N_1839);
or U2122 (N_2122,N_1739,N_1788);
and U2123 (N_2123,N_1790,N_1841);
or U2124 (N_2124,N_1888,N_1761);
nor U2125 (N_2125,N_1825,N_1815);
or U2126 (N_2126,N_1763,N_1560);
nor U2127 (N_2127,N_1588,N_1614);
nor U2128 (N_2128,N_1553,N_1610);
or U2129 (N_2129,N_1976,N_1690);
nand U2130 (N_2130,N_1592,N_1706);
nor U2131 (N_2131,N_1621,N_1875);
or U2132 (N_2132,N_1900,N_1994);
or U2133 (N_2133,N_1726,N_1741);
nand U2134 (N_2134,N_1528,N_1781);
nand U2135 (N_2135,N_1572,N_1717);
nand U2136 (N_2136,N_1866,N_1604);
or U2137 (N_2137,N_1939,N_1784);
nand U2138 (N_2138,N_1767,N_1630);
and U2139 (N_2139,N_1688,N_1668);
nor U2140 (N_2140,N_1858,N_1673);
nor U2141 (N_2141,N_1517,N_1579);
nand U2142 (N_2142,N_1818,N_1522);
nor U2143 (N_2143,N_1988,N_1778);
or U2144 (N_2144,N_1898,N_1830);
and U2145 (N_2145,N_1889,N_1843);
and U2146 (N_2146,N_1979,N_1793);
nor U2147 (N_2147,N_1589,N_1571);
nand U2148 (N_2148,N_1750,N_1657);
or U2149 (N_2149,N_1595,N_1662);
and U2150 (N_2150,N_1504,N_1998);
or U2151 (N_2151,N_1870,N_1500);
nand U2152 (N_2152,N_1770,N_1854);
and U2153 (N_2153,N_1742,N_1532);
nor U2154 (N_2154,N_1587,N_1990);
and U2155 (N_2155,N_1596,N_1651);
nand U2156 (N_2156,N_1777,N_1869);
or U2157 (N_2157,N_1747,N_1691);
nor U2158 (N_2158,N_1871,N_1808);
and U2159 (N_2159,N_1989,N_1744);
xnor U2160 (N_2160,N_1917,N_1509);
and U2161 (N_2161,N_1915,N_1924);
nand U2162 (N_2162,N_1857,N_1734);
or U2163 (N_2163,N_1751,N_1796);
nor U2164 (N_2164,N_1894,N_1773);
and U2165 (N_2165,N_1876,N_1506);
and U2166 (N_2166,N_1555,N_1937);
or U2167 (N_2167,N_1848,N_1980);
nor U2168 (N_2168,N_1718,N_1525);
and U2169 (N_2169,N_1590,N_1966);
nor U2170 (N_2170,N_1521,N_1918);
and U2171 (N_2171,N_1705,N_1940);
and U2172 (N_2172,N_1585,N_1834);
nand U2173 (N_2173,N_1813,N_1670);
and U2174 (N_2174,N_1516,N_1719);
nand U2175 (N_2175,N_1672,N_1689);
or U2176 (N_2176,N_1515,N_1655);
or U2177 (N_2177,N_1746,N_1625);
and U2178 (N_2178,N_1659,N_1973);
and U2179 (N_2179,N_1710,N_1745);
and U2180 (N_2180,N_1561,N_1541);
and U2181 (N_2181,N_1982,N_1845);
or U2182 (N_2182,N_1847,N_1735);
or U2183 (N_2183,N_1601,N_1738);
nand U2184 (N_2184,N_1583,N_1578);
and U2185 (N_2185,N_1879,N_1731);
nand U2186 (N_2186,N_1693,N_1884);
and U2187 (N_2187,N_1944,N_1616);
nor U2188 (N_2188,N_1953,N_1961);
or U2189 (N_2189,N_1827,N_1550);
and U2190 (N_2190,N_1562,N_1933);
nor U2191 (N_2191,N_1775,N_1665);
nor U2192 (N_2192,N_1664,N_1743);
or U2193 (N_2193,N_1613,N_1703);
and U2194 (N_2194,N_1716,N_1684);
and U2195 (N_2195,N_1696,N_1772);
and U2196 (N_2196,N_1975,N_1965);
nor U2197 (N_2197,N_1853,N_1540);
and U2198 (N_2198,N_1594,N_1645);
or U2199 (N_2199,N_1867,N_1786);
and U2200 (N_2200,N_1677,N_1897);
nand U2201 (N_2201,N_1783,N_1683);
nor U2202 (N_2202,N_1948,N_1582);
nor U2203 (N_2203,N_1658,N_1607);
nor U2204 (N_2204,N_1822,N_1535);
nand U2205 (N_2205,N_1737,N_1896);
nor U2206 (N_2206,N_1697,N_1779);
or U2207 (N_2207,N_1642,N_1527);
nand U2208 (N_2208,N_1883,N_1972);
or U2209 (N_2209,N_1567,N_1581);
or U2210 (N_2210,N_1861,N_1656);
and U2211 (N_2211,N_1946,N_1959);
nand U2212 (N_2212,N_1945,N_1537);
nand U2213 (N_2213,N_1682,N_1507);
nand U2214 (N_2214,N_1812,N_1602);
and U2215 (N_2215,N_1736,N_1925);
or U2216 (N_2216,N_1538,N_1926);
and U2217 (N_2217,N_1564,N_1510);
nand U2218 (N_2218,N_1798,N_1864);
or U2219 (N_2219,N_1603,N_1831);
nor U2220 (N_2220,N_1969,N_1873);
or U2221 (N_2221,N_1599,N_1968);
or U2222 (N_2222,N_1539,N_1654);
nand U2223 (N_2223,N_1618,N_1667);
nand U2224 (N_2224,N_1707,N_1728);
and U2225 (N_2225,N_1833,N_1724);
nand U2226 (N_2226,N_1648,N_1760);
nor U2227 (N_2227,N_1551,N_1941);
and U2228 (N_2228,N_1820,N_1780);
nor U2229 (N_2229,N_1641,N_1722);
nor U2230 (N_2230,N_1685,N_1806);
and U2231 (N_2231,N_1991,N_1713);
nand U2232 (N_2232,N_1574,N_1803);
nand U2233 (N_2233,N_1534,N_1910);
and U2234 (N_2234,N_1647,N_1612);
and U2235 (N_2235,N_1545,N_1996);
nor U2236 (N_2236,N_1805,N_1997);
or U2237 (N_2237,N_1931,N_1950);
nor U2238 (N_2238,N_1844,N_1700);
nand U2239 (N_2239,N_1531,N_1860);
nor U2240 (N_2240,N_1955,N_1960);
nor U2241 (N_2241,N_1611,N_1649);
or U2242 (N_2242,N_1620,N_1699);
and U2243 (N_2243,N_1874,N_1544);
or U2244 (N_2244,N_1597,N_1908);
and U2245 (N_2245,N_1913,N_1653);
or U2246 (N_2246,N_1552,N_1523);
or U2247 (N_2247,N_1575,N_1756);
nand U2248 (N_2248,N_1821,N_1512);
nor U2249 (N_2249,N_1730,N_1639);
and U2250 (N_2250,N_1754,N_1852);
or U2251 (N_2251,N_1678,N_1659);
nor U2252 (N_2252,N_1636,N_1551);
or U2253 (N_2253,N_1837,N_1651);
or U2254 (N_2254,N_1939,N_1607);
nor U2255 (N_2255,N_1852,N_1563);
and U2256 (N_2256,N_1833,N_1524);
or U2257 (N_2257,N_1958,N_1795);
and U2258 (N_2258,N_1546,N_1593);
nor U2259 (N_2259,N_1574,N_1504);
nor U2260 (N_2260,N_1691,N_1865);
nand U2261 (N_2261,N_1687,N_1972);
or U2262 (N_2262,N_1842,N_1814);
nor U2263 (N_2263,N_1932,N_1944);
nor U2264 (N_2264,N_1707,N_1561);
or U2265 (N_2265,N_1688,N_1926);
nand U2266 (N_2266,N_1953,N_1754);
nand U2267 (N_2267,N_1879,N_1726);
nand U2268 (N_2268,N_1547,N_1947);
or U2269 (N_2269,N_1803,N_1767);
nand U2270 (N_2270,N_1765,N_1645);
and U2271 (N_2271,N_1584,N_1766);
nor U2272 (N_2272,N_1581,N_1989);
nand U2273 (N_2273,N_1504,N_1792);
or U2274 (N_2274,N_1699,N_1512);
nor U2275 (N_2275,N_1512,N_1958);
or U2276 (N_2276,N_1695,N_1831);
or U2277 (N_2277,N_1541,N_1864);
nor U2278 (N_2278,N_1921,N_1614);
nor U2279 (N_2279,N_1792,N_1601);
or U2280 (N_2280,N_1534,N_1823);
nor U2281 (N_2281,N_1646,N_1953);
and U2282 (N_2282,N_1993,N_1802);
or U2283 (N_2283,N_1631,N_1731);
nand U2284 (N_2284,N_1696,N_1654);
nand U2285 (N_2285,N_1574,N_1770);
or U2286 (N_2286,N_1607,N_1951);
and U2287 (N_2287,N_1629,N_1800);
and U2288 (N_2288,N_1960,N_1655);
and U2289 (N_2289,N_1748,N_1644);
or U2290 (N_2290,N_1652,N_1955);
and U2291 (N_2291,N_1844,N_1596);
and U2292 (N_2292,N_1605,N_1578);
nor U2293 (N_2293,N_1606,N_1791);
nor U2294 (N_2294,N_1748,N_1849);
nand U2295 (N_2295,N_1990,N_1656);
or U2296 (N_2296,N_1842,N_1896);
or U2297 (N_2297,N_1856,N_1601);
or U2298 (N_2298,N_1794,N_1838);
xor U2299 (N_2299,N_1829,N_1511);
nand U2300 (N_2300,N_1838,N_1780);
nor U2301 (N_2301,N_1556,N_1763);
nand U2302 (N_2302,N_1650,N_1583);
nand U2303 (N_2303,N_1566,N_1855);
or U2304 (N_2304,N_1629,N_1788);
nor U2305 (N_2305,N_1718,N_1918);
nor U2306 (N_2306,N_1891,N_1532);
nand U2307 (N_2307,N_1689,N_1812);
nor U2308 (N_2308,N_1559,N_1772);
nand U2309 (N_2309,N_1980,N_1930);
or U2310 (N_2310,N_1940,N_1701);
or U2311 (N_2311,N_1546,N_1747);
or U2312 (N_2312,N_1587,N_1920);
nor U2313 (N_2313,N_1768,N_1980);
nand U2314 (N_2314,N_1633,N_1947);
and U2315 (N_2315,N_1899,N_1920);
nand U2316 (N_2316,N_1784,N_1710);
nor U2317 (N_2317,N_1758,N_1845);
nand U2318 (N_2318,N_1671,N_1912);
nor U2319 (N_2319,N_1726,N_1865);
and U2320 (N_2320,N_1560,N_1959);
or U2321 (N_2321,N_1906,N_1965);
nand U2322 (N_2322,N_1664,N_1518);
nor U2323 (N_2323,N_1854,N_1723);
and U2324 (N_2324,N_1872,N_1772);
nand U2325 (N_2325,N_1777,N_1724);
nor U2326 (N_2326,N_1731,N_1642);
and U2327 (N_2327,N_1586,N_1873);
or U2328 (N_2328,N_1718,N_1823);
or U2329 (N_2329,N_1943,N_1510);
and U2330 (N_2330,N_1872,N_1806);
nor U2331 (N_2331,N_1565,N_1704);
nand U2332 (N_2332,N_1840,N_1600);
and U2333 (N_2333,N_1665,N_1805);
nor U2334 (N_2334,N_1913,N_1515);
and U2335 (N_2335,N_1687,N_1569);
nor U2336 (N_2336,N_1776,N_1855);
or U2337 (N_2337,N_1648,N_1646);
nand U2338 (N_2338,N_1867,N_1534);
nor U2339 (N_2339,N_1753,N_1871);
and U2340 (N_2340,N_1801,N_1914);
or U2341 (N_2341,N_1720,N_1585);
or U2342 (N_2342,N_1626,N_1901);
or U2343 (N_2343,N_1955,N_1815);
nand U2344 (N_2344,N_1609,N_1606);
and U2345 (N_2345,N_1904,N_1897);
or U2346 (N_2346,N_1808,N_1623);
or U2347 (N_2347,N_1693,N_1847);
and U2348 (N_2348,N_1874,N_1863);
and U2349 (N_2349,N_1679,N_1606);
or U2350 (N_2350,N_1722,N_1693);
or U2351 (N_2351,N_1927,N_1741);
nor U2352 (N_2352,N_1910,N_1557);
or U2353 (N_2353,N_1510,N_1593);
or U2354 (N_2354,N_1534,N_1631);
and U2355 (N_2355,N_1588,N_1894);
or U2356 (N_2356,N_1614,N_1742);
nor U2357 (N_2357,N_1599,N_1884);
nor U2358 (N_2358,N_1745,N_1510);
and U2359 (N_2359,N_1756,N_1722);
and U2360 (N_2360,N_1707,N_1649);
and U2361 (N_2361,N_1633,N_1643);
and U2362 (N_2362,N_1673,N_1733);
or U2363 (N_2363,N_1560,N_1984);
nand U2364 (N_2364,N_1775,N_1574);
or U2365 (N_2365,N_1886,N_1858);
nor U2366 (N_2366,N_1695,N_1533);
nand U2367 (N_2367,N_1836,N_1961);
or U2368 (N_2368,N_1997,N_1984);
nor U2369 (N_2369,N_1805,N_1675);
xnor U2370 (N_2370,N_1816,N_1599);
nor U2371 (N_2371,N_1820,N_1988);
nand U2372 (N_2372,N_1526,N_1661);
or U2373 (N_2373,N_1504,N_1859);
nand U2374 (N_2374,N_1540,N_1934);
nor U2375 (N_2375,N_1991,N_1883);
nand U2376 (N_2376,N_1610,N_1929);
nor U2377 (N_2377,N_1860,N_1614);
nand U2378 (N_2378,N_1530,N_1794);
nor U2379 (N_2379,N_1735,N_1932);
nand U2380 (N_2380,N_1860,N_1520);
or U2381 (N_2381,N_1779,N_1920);
nand U2382 (N_2382,N_1927,N_1615);
nor U2383 (N_2383,N_1917,N_1734);
nand U2384 (N_2384,N_1765,N_1608);
and U2385 (N_2385,N_1928,N_1910);
nor U2386 (N_2386,N_1518,N_1729);
and U2387 (N_2387,N_1875,N_1552);
nand U2388 (N_2388,N_1903,N_1981);
and U2389 (N_2389,N_1710,N_1783);
and U2390 (N_2390,N_1697,N_1947);
nor U2391 (N_2391,N_1537,N_1841);
nor U2392 (N_2392,N_1818,N_1952);
nor U2393 (N_2393,N_1610,N_1557);
nand U2394 (N_2394,N_1762,N_1859);
nor U2395 (N_2395,N_1803,N_1757);
or U2396 (N_2396,N_1666,N_1632);
and U2397 (N_2397,N_1830,N_1755);
and U2398 (N_2398,N_1517,N_1537);
nor U2399 (N_2399,N_1927,N_1919);
or U2400 (N_2400,N_1703,N_1916);
and U2401 (N_2401,N_1929,N_1542);
nor U2402 (N_2402,N_1687,N_1811);
nand U2403 (N_2403,N_1570,N_1805);
and U2404 (N_2404,N_1841,N_1934);
nor U2405 (N_2405,N_1767,N_1859);
nor U2406 (N_2406,N_1537,N_1934);
and U2407 (N_2407,N_1965,N_1898);
or U2408 (N_2408,N_1866,N_1770);
or U2409 (N_2409,N_1823,N_1500);
or U2410 (N_2410,N_1936,N_1833);
or U2411 (N_2411,N_1751,N_1820);
nor U2412 (N_2412,N_1791,N_1523);
nor U2413 (N_2413,N_1589,N_1753);
or U2414 (N_2414,N_1578,N_1952);
and U2415 (N_2415,N_1787,N_1586);
nor U2416 (N_2416,N_1700,N_1706);
or U2417 (N_2417,N_1983,N_1547);
or U2418 (N_2418,N_1593,N_1792);
nor U2419 (N_2419,N_1694,N_1631);
or U2420 (N_2420,N_1989,N_1901);
or U2421 (N_2421,N_1909,N_1860);
or U2422 (N_2422,N_1535,N_1930);
or U2423 (N_2423,N_1632,N_1642);
or U2424 (N_2424,N_1865,N_1666);
nand U2425 (N_2425,N_1895,N_1818);
nand U2426 (N_2426,N_1606,N_1862);
nand U2427 (N_2427,N_1782,N_1701);
nand U2428 (N_2428,N_1882,N_1674);
nand U2429 (N_2429,N_1951,N_1641);
nor U2430 (N_2430,N_1803,N_1809);
and U2431 (N_2431,N_1801,N_1725);
and U2432 (N_2432,N_1700,N_1712);
and U2433 (N_2433,N_1900,N_1609);
and U2434 (N_2434,N_1750,N_1588);
xor U2435 (N_2435,N_1981,N_1718);
nand U2436 (N_2436,N_1742,N_1786);
nand U2437 (N_2437,N_1964,N_1634);
nand U2438 (N_2438,N_1835,N_1715);
nand U2439 (N_2439,N_1937,N_1778);
or U2440 (N_2440,N_1832,N_1640);
and U2441 (N_2441,N_1999,N_1989);
nand U2442 (N_2442,N_1682,N_1815);
nor U2443 (N_2443,N_1869,N_1929);
nor U2444 (N_2444,N_1615,N_1778);
or U2445 (N_2445,N_1568,N_1908);
or U2446 (N_2446,N_1946,N_1783);
or U2447 (N_2447,N_1833,N_1742);
and U2448 (N_2448,N_1575,N_1615);
and U2449 (N_2449,N_1944,N_1806);
and U2450 (N_2450,N_1956,N_1751);
and U2451 (N_2451,N_1847,N_1632);
and U2452 (N_2452,N_1710,N_1962);
nor U2453 (N_2453,N_1658,N_1608);
and U2454 (N_2454,N_1965,N_1875);
or U2455 (N_2455,N_1632,N_1745);
nor U2456 (N_2456,N_1692,N_1999);
or U2457 (N_2457,N_1550,N_1723);
nand U2458 (N_2458,N_1621,N_1961);
nor U2459 (N_2459,N_1782,N_1998);
nand U2460 (N_2460,N_1525,N_1967);
or U2461 (N_2461,N_1839,N_1816);
nand U2462 (N_2462,N_1665,N_1693);
and U2463 (N_2463,N_1526,N_1902);
nor U2464 (N_2464,N_1967,N_1776);
or U2465 (N_2465,N_1820,N_1783);
nand U2466 (N_2466,N_1843,N_1833);
nor U2467 (N_2467,N_1590,N_1546);
or U2468 (N_2468,N_1745,N_1821);
or U2469 (N_2469,N_1740,N_1566);
nand U2470 (N_2470,N_1734,N_1728);
and U2471 (N_2471,N_1804,N_1906);
nand U2472 (N_2472,N_1538,N_1694);
and U2473 (N_2473,N_1986,N_1969);
or U2474 (N_2474,N_1529,N_1769);
or U2475 (N_2475,N_1829,N_1727);
or U2476 (N_2476,N_1964,N_1563);
nand U2477 (N_2477,N_1551,N_1741);
and U2478 (N_2478,N_1753,N_1639);
nand U2479 (N_2479,N_1981,N_1662);
and U2480 (N_2480,N_1833,N_1510);
nand U2481 (N_2481,N_1509,N_1862);
nand U2482 (N_2482,N_1882,N_1979);
nor U2483 (N_2483,N_1596,N_1924);
nand U2484 (N_2484,N_1900,N_1561);
or U2485 (N_2485,N_1551,N_1833);
or U2486 (N_2486,N_1538,N_1876);
and U2487 (N_2487,N_1930,N_1892);
and U2488 (N_2488,N_1615,N_1819);
nand U2489 (N_2489,N_1635,N_1728);
or U2490 (N_2490,N_1895,N_1759);
nand U2491 (N_2491,N_1590,N_1750);
nand U2492 (N_2492,N_1502,N_1872);
nor U2493 (N_2493,N_1590,N_1632);
nor U2494 (N_2494,N_1889,N_1721);
nand U2495 (N_2495,N_1539,N_1563);
and U2496 (N_2496,N_1868,N_1550);
or U2497 (N_2497,N_1943,N_1843);
nor U2498 (N_2498,N_1882,N_1521);
or U2499 (N_2499,N_1976,N_1678);
nor U2500 (N_2500,N_2282,N_2317);
nor U2501 (N_2501,N_2321,N_2355);
nor U2502 (N_2502,N_2346,N_2224);
nor U2503 (N_2503,N_2125,N_2376);
nor U2504 (N_2504,N_2336,N_2203);
or U2505 (N_2505,N_2131,N_2001);
and U2506 (N_2506,N_2470,N_2169);
nor U2507 (N_2507,N_2495,N_2497);
nor U2508 (N_2508,N_2366,N_2049);
nand U2509 (N_2509,N_2303,N_2420);
nand U2510 (N_2510,N_2273,N_2426);
nand U2511 (N_2511,N_2486,N_2374);
or U2512 (N_2512,N_2348,N_2188);
or U2513 (N_2513,N_2124,N_2425);
nor U2514 (N_2514,N_2380,N_2270);
nor U2515 (N_2515,N_2170,N_2084);
or U2516 (N_2516,N_2061,N_2266);
nand U2517 (N_2517,N_2329,N_2216);
nor U2518 (N_2518,N_2221,N_2096);
or U2519 (N_2519,N_2372,N_2387);
nor U2520 (N_2520,N_2293,N_2173);
nor U2521 (N_2521,N_2073,N_2043);
or U2522 (N_2522,N_2256,N_2069);
nand U2523 (N_2523,N_2441,N_2236);
nand U2524 (N_2524,N_2166,N_2119);
nand U2525 (N_2525,N_2085,N_2029);
or U2526 (N_2526,N_2167,N_2245);
or U2527 (N_2527,N_2455,N_2337);
or U2528 (N_2528,N_2250,N_2064);
nor U2529 (N_2529,N_2395,N_2031);
or U2530 (N_2530,N_2295,N_2392);
nor U2531 (N_2531,N_2230,N_2396);
nor U2532 (N_2532,N_2060,N_2363);
or U2533 (N_2533,N_2429,N_2254);
or U2534 (N_2534,N_2118,N_2264);
or U2535 (N_2535,N_2228,N_2488);
or U2536 (N_2536,N_2445,N_2422);
or U2537 (N_2537,N_2176,N_2491);
or U2538 (N_2538,N_2186,N_2474);
and U2539 (N_2539,N_2121,N_2241);
or U2540 (N_2540,N_2105,N_2283);
or U2541 (N_2541,N_2385,N_2034);
nand U2542 (N_2542,N_2150,N_2180);
xor U2543 (N_2543,N_2259,N_2021);
nand U2544 (N_2544,N_2443,N_2432);
or U2545 (N_2545,N_2151,N_2223);
or U2546 (N_2546,N_2431,N_2171);
or U2547 (N_2547,N_2292,N_2407);
nand U2548 (N_2548,N_2162,N_2101);
and U2549 (N_2549,N_2020,N_2490);
and U2550 (N_2550,N_2314,N_2319);
nor U2551 (N_2551,N_2251,N_2320);
nand U2552 (N_2552,N_2227,N_2424);
nor U2553 (N_2553,N_2377,N_2435);
or U2554 (N_2554,N_2439,N_2214);
nor U2555 (N_2555,N_2480,N_2217);
or U2556 (N_2556,N_2107,N_2233);
or U2557 (N_2557,N_2145,N_2464);
or U2558 (N_2558,N_2129,N_2433);
or U2559 (N_2559,N_2370,N_2094);
nor U2560 (N_2560,N_2209,N_2326);
or U2561 (N_2561,N_2324,N_2197);
or U2562 (N_2562,N_2100,N_2479);
or U2563 (N_2563,N_2017,N_2436);
xnor U2564 (N_2564,N_2083,N_2373);
nand U2565 (N_2565,N_2413,N_2123);
or U2566 (N_2566,N_2262,N_2072);
nand U2567 (N_2567,N_2446,N_2165);
nand U2568 (N_2568,N_2218,N_2331);
nand U2569 (N_2569,N_2114,N_2229);
nor U2570 (N_2570,N_2352,N_2386);
nand U2571 (N_2571,N_2014,N_2341);
and U2572 (N_2572,N_2322,N_2333);
and U2573 (N_2573,N_2112,N_2378);
nand U2574 (N_2574,N_2304,N_2057);
or U2575 (N_2575,N_2133,N_2406);
or U2576 (N_2576,N_2247,N_2260);
or U2577 (N_2577,N_2279,N_2063);
and U2578 (N_2578,N_2198,N_2409);
xor U2579 (N_2579,N_2397,N_2185);
nor U2580 (N_2580,N_2059,N_2301);
nand U2581 (N_2581,N_2065,N_2110);
and U2582 (N_2582,N_2115,N_2332);
or U2583 (N_2583,N_2290,N_2234);
nand U2584 (N_2584,N_2484,N_2312);
or U2585 (N_2585,N_2210,N_2277);
and U2586 (N_2586,N_2461,N_2405);
nor U2587 (N_2587,N_2257,N_2485);
nand U2588 (N_2588,N_2196,N_2310);
nand U2589 (N_2589,N_2062,N_2442);
or U2590 (N_2590,N_2371,N_2369);
nand U2591 (N_2591,N_2242,N_2481);
nor U2592 (N_2592,N_2074,N_2010);
nor U2593 (N_2593,N_2231,N_2201);
nand U2594 (N_2594,N_2309,N_2478);
or U2595 (N_2595,N_2476,N_2106);
or U2596 (N_2596,N_2416,N_2238);
and U2597 (N_2597,N_2161,N_2421);
and U2598 (N_2598,N_2291,N_2354);
nor U2599 (N_2599,N_2012,N_2349);
nand U2600 (N_2600,N_2274,N_2297);
or U2601 (N_2601,N_2148,N_2360);
nand U2602 (N_2602,N_2097,N_2434);
or U2603 (N_2603,N_2459,N_2206);
nor U2604 (N_2604,N_2207,N_2302);
nor U2605 (N_2605,N_2335,N_2306);
and U2606 (N_2606,N_2286,N_2456);
or U2607 (N_2607,N_2122,N_2163);
nor U2608 (N_2608,N_2184,N_2313);
xnor U2609 (N_2609,N_2200,N_2258);
nand U2610 (N_2610,N_2268,N_2038);
nor U2611 (N_2611,N_2368,N_2089);
and U2612 (N_2612,N_2493,N_2095);
nor U2613 (N_2613,N_2299,N_2158);
nand U2614 (N_2614,N_2391,N_2437);
nand U2615 (N_2615,N_2452,N_2454);
nand U2616 (N_2616,N_2127,N_2111);
and U2617 (N_2617,N_2356,N_2120);
or U2618 (N_2618,N_2382,N_2323);
and U2619 (N_2619,N_2492,N_2342);
nor U2620 (N_2620,N_2311,N_2460);
and U2621 (N_2621,N_2149,N_2152);
or U2622 (N_2622,N_2006,N_2237);
or U2623 (N_2623,N_2141,N_2033);
nand U2624 (N_2624,N_2081,N_2272);
nor U2625 (N_2625,N_2410,N_2157);
nand U2626 (N_2626,N_2213,N_2082);
nand U2627 (N_2627,N_2450,N_2086);
and U2628 (N_2628,N_2343,N_2136);
nor U2629 (N_2629,N_2202,N_2177);
nand U2630 (N_2630,N_2199,N_2281);
nor U2631 (N_2631,N_2155,N_2467);
nor U2632 (N_2632,N_2246,N_2267);
or U2633 (N_2633,N_2076,N_2253);
nand U2634 (N_2634,N_2179,N_2330);
or U2635 (N_2635,N_2019,N_2305);
nor U2636 (N_2636,N_2025,N_2427);
nand U2637 (N_2637,N_2411,N_2004);
nor U2638 (N_2638,N_2013,N_2002);
nor U2639 (N_2639,N_2191,N_2130);
nand U2640 (N_2640,N_2448,N_2102);
nor U2641 (N_2641,N_2142,N_2359);
nand U2642 (N_2642,N_2007,N_2126);
and U2643 (N_2643,N_2023,N_2402);
xor U2644 (N_2644,N_2249,N_2092);
nor U2645 (N_2645,N_2219,N_2022);
nor U2646 (N_2646,N_2164,N_2389);
or U2647 (N_2647,N_2080,N_2153);
and U2648 (N_2648,N_2350,N_2071);
nand U2649 (N_2649,N_2175,N_2364);
nand U2650 (N_2650,N_2487,N_2362);
or U2651 (N_2651,N_2016,N_2318);
and U2652 (N_2652,N_2339,N_2090);
nor U2653 (N_2653,N_2208,N_2394);
or U2654 (N_2654,N_2139,N_2466);
nor U2655 (N_2655,N_2398,N_2052);
or U2656 (N_2656,N_2183,N_2357);
or U2657 (N_2657,N_2172,N_2271);
or U2658 (N_2658,N_2269,N_2109);
and U2659 (N_2659,N_2296,N_2401);
nand U2660 (N_2660,N_2030,N_2381);
and U2661 (N_2661,N_2168,N_2351);
or U2662 (N_2662,N_2462,N_2367);
nor U2663 (N_2663,N_2220,N_2103);
nor U2664 (N_2664,N_2032,N_2104);
nand U2665 (N_2665,N_2015,N_2027);
or U2666 (N_2666,N_2018,N_2138);
nand U2667 (N_2667,N_2154,N_2423);
or U2668 (N_2668,N_2046,N_2365);
nand U2669 (N_2669,N_2316,N_2066);
and U2670 (N_2670,N_2211,N_2419);
nand U2671 (N_2671,N_2428,N_2040);
or U2672 (N_2672,N_2050,N_2047);
nand U2673 (N_2673,N_2134,N_2128);
and U2674 (N_2674,N_2132,N_2300);
nand U2675 (N_2675,N_2334,N_2340);
or U2676 (N_2676,N_2144,N_2280);
nand U2677 (N_2677,N_2353,N_2026);
or U2678 (N_2678,N_2189,N_2137);
and U2679 (N_2679,N_2388,N_2054);
nor U2680 (N_2680,N_2393,N_2225);
nand U2681 (N_2681,N_2327,N_2159);
or U2682 (N_2682,N_2099,N_2463);
or U2683 (N_2683,N_2325,N_2068);
or U2684 (N_2684,N_2451,N_2117);
or U2685 (N_2685,N_2156,N_2498);
and U2686 (N_2686,N_2265,N_2414);
or U2687 (N_2687,N_2344,N_2496);
nand U2688 (N_2688,N_2289,N_2041);
or U2689 (N_2689,N_2375,N_2244);
or U2690 (N_2690,N_2240,N_2070);
and U2691 (N_2691,N_2193,N_2383);
or U2692 (N_2692,N_2499,N_2028);
and U2693 (N_2693,N_2307,N_2178);
nor U2694 (N_2694,N_2205,N_2473);
or U2695 (N_2695,N_2252,N_2358);
nand U2696 (N_2696,N_2048,N_2039);
and U2697 (N_2697,N_2143,N_2475);
or U2698 (N_2698,N_2042,N_2024);
or U2699 (N_2699,N_2494,N_2035);
and U2700 (N_2700,N_2078,N_2438);
nor U2701 (N_2701,N_2000,N_2255);
or U2702 (N_2702,N_2472,N_2408);
nand U2703 (N_2703,N_2449,N_2384);
nor U2704 (N_2704,N_2285,N_2412);
or U2705 (N_2705,N_2404,N_2093);
nand U2706 (N_2706,N_2204,N_2051);
and U2707 (N_2707,N_2056,N_2075);
or U2708 (N_2708,N_2284,N_2160);
and U2709 (N_2709,N_2308,N_2036);
nor U2710 (N_2710,N_2403,N_2079);
and U2711 (N_2711,N_2471,N_2108);
nand U2712 (N_2712,N_2288,N_2328);
and U2713 (N_2713,N_2418,N_2465);
and U2714 (N_2714,N_2190,N_2037);
and U2715 (N_2715,N_2055,N_2468);
nor U2716 (N_2716,N_2009,N_2187);
nand U2717 (N_2717,N_2399,N_2003);
or U2718 (N_2718,N_2058,N_2011);
nor U2719 (N_2719,N_2215,N_2345);
and U2720 (N_2720,N_2379,N_2005);
or U2721 (N_2721,N_2116,N_2181);
or U2722 (N_2722,N_2430,N_2239);
nor U2723 (N_2723,N_2243,N_2261);
and U2724 (N_2724,N_2444,N_2192);
and U2725 (N_2725,N_2469,N_2477);
and U2726 (N_2726,N_2457,N_2417);
or U2727 (N_2727,N_2489,N_2222);
nand U2728 (N_2728,N_2453,N_2482);
and U2729 (N_2729,N_2113,N_2400);
and U2730 (N_2730,N_2087,N_2338);
nand U2731 (N_2731,N_2212,N_2182);
or U2732 (N_2732,N_2053,N_2278);
nand U2733 (N_2733,N_2483,N_2390);
and U2734 (N_2734,N_2088,N_2091);
nor U2735 (N_2735,N_2235,N_2226);
or U2736 (N_2736,N_2447,N_2077);
nand U2737 (N_2737,N_2045,N_2440);
nor U2738 (N_2738,N_2415,N_2458);
or U2739 (N_2739,N_2194,N_2294);
or U2740 (N_2740,N_2195,N_2298);
nor U2741 (N_2741,N_2287,N_2315);
nor U2742 (N_2742,N_2098,N_2174);
and U2743 (N_2743,N_2275,N_2140);
nand U2744 (N_2744,N_2147,N_2146);
or U2745 (N_2745,N_2347,N_2067);
or U2746 (N_2746,N_2135,N_2361);
nor U2747 (N_2747,N_2232,N_2008);
or U2748 (N_2748,N_2248,N_2263);
and U2749 (N_2749,N_2276,N_2044);
nor U2750 (N_2750,N_2263,N_2063);
or U2751 (N_2751,N_2406,N_2424);
nor U2752 (N_2752,N_2141,N_2229);
nand U2753 (N_2753,N_2091,N_2403);
or U2754 (N_2754,N_2489,N_2104);
or U2755 (N_2755,N_2080,N_2492);
nor U2756 (N_2756,N_2034,N_2406);
nor U2757 (N_2757,N_2285,N_2024);
or U2758 (N_2758,N_2416,N_2333);
or U2759 (N_2759,N_2340,N_2127);
and U2760 (N_2760,N_2254,N_2203);
nand U2761 (N_2761,N_2132,N_2435);
nor U2762 (N_2762,N_2455,N_2300);
or U2763 (N_2763,N_2287,N_2280);
nand U2764 (N_2764,N_2310,N_2323);
nor U2765 (N_2765,N_2056,N_2449);
and U2766 (N_2766,N_2181,N_2489);
and U2767 (N_2767,N_2230,N_2132);
or U2768 (N_2768,N_2428,N_2325);
nand U2769 (N_2769,N_2219,N_2054);
nand U2770 (N_2770,N_2004,N_2088);
or U2771 (N_2771,N_2122,N_2240);
nand U2772 (N_2772,N_2386,N_2093);
and U2773 (N_2773,N_2343,N_2295);
nand U2774 (N_2774,N_2463,N_2283);
and U2775 (N_2775,N_2497,N_2444);
and U2776 (N_2776,N_2283,N_2334);
and U2777 (N_2777,N_2158,N_2386);
or U2778 (N_2778,N_2258,N_2261);
or U2779 (N_2779,N_2013,N_2112);
nand U2780 (N_2780,N_2031,N_2336);
or U2781 (N_2781,N_2212,N_2031);
nor U2782 (N_2782,N_2224,N_2349);
nor U2783 (N_2783,N_2052,N_2486);
and U2784 (N_2784,N_2408,N_2038);
nand U2785 (N_2785,N_2389,N_2407);
or U2786 (N_2786,N_2167,N_2429);
or U2787 (N_2787,N_2293,N_2366);
and U2788 (N_2788,N_2418,N_2493);
nand U2789 (N_2789,N_2274,N_2219);
nand U2790 (N_2790,N_2206,N_2118);
and U2791 (N_2791,N_2446,N_2399);
and U2792 (N_2792,N_2439,N_2092);
or U2793 (N_2793,N_2163,N_2258);
or U2794 (N_2794,N_2298,N_2225);
or U2795 (N_2795,N_2117,N_2239);
nand U2796 (N_2796,N_2055,N_2080);
or U2797 (N_2797,N_2463,N_2142);
and U2798 (N_2798,N_2443,N_2302);
nand U2799 (N_2799,N_2123,N_2460);
nand U2800 (N_2800,N_2077,N_2277);
nand U2801 (N_2801,N_2418,N_2442);
nor U2802 (N_2802,N_2390,N_2067);
and U2803 (N_2803,N_2309,N_2370);
nor U2804 (N_2804,N_2065,N_2055);
nor U2805 (N_2805,N_2087,N_2169);
xor U2806 (N_2806,N_2309,N_2158);
nand U2807 (N_2807,N_2003,N_2406);
nand U2808 (N_2808,N_2384,N_2043);
nor U2809 (N_2809,N_2409,N_2067);
nor U2810 (N_2810,N_2123,N_2045);
or U2811 (N_2811,N_2263,N_2082);
nor U2812 (N_2812,N_2113,N_2477);
and U2813 (N_2813,N_2225,N_2231);
or U2814 (N_2814,N_2460,N_2432);
nand U2815 (N_2815,N_2473,N_2307);
nand U2816 (N_2816,N_2045,N_2048);
nor U2817 (N_2817,N_2410,N_2029);
nor U2818 (N_2818,N_2485,N_2068);
nor U2819 (N_2819,N_2415,N_2360);
or U2820 (N_2820,N_2256,N_2252);
nor U2821 (N_2821,N_2308,N_2027);
and U2822 (N_2822,N_2299,N_2061);
nor U2823 (N_2823,N_2197,N_2354);
and U2824 (N_2824,N_2149,N_2090);
nor U2825 (N_2825,N_2003,N_2361);
xor U2826 (N_2826,N_2393,N_2475);
or U2827 (N_2827,N_2391,N_2248);
nor U2828 (N_2828,N_2218,N_2285);
and U2829 (N_2829,N_2005,N_2377);
or U2830 (N_2830,N_2413,N_2369);
and U2831 (N_2831,N_2381,N_2348);
nand U2832 (N_2832,N_2033,N_2136);
and U2833 (N_2833,N_2279,N_2201);
nor U2834 (N_2834,N_2161,N_2021);
nand U2835 (N_2835,N_2225,N_2040);
nor U2836 (N_2836,N_2444,N_2181);
and U2837 (N_2837,N_2328,N_2254);
nand U2838 (N_2838,N_2411,N_2397);
and U2839 (N_2839,N_2285,N_2102);
nand U2840 (N_2840,N_2171,N_2120);
nor U2841 (N_2841,N_2079,N_2103);
or U2842 (N_2842,N_2276,N_2185);
and U2843 (N_2843,N_2272,N_2456);
nand U2844 (N_2844,N_2331,N_2189);
nor U2845 (N_2845,N_2135,N_2143);
or U2846 (N_2846,N_2249,N_2370);
and U2847 (N_2847,N_2345,N_2162);
nor U2848 (N_2848,N_2175,N_2248);
and U2849 (N_2849,N_2102,N_2271);
nand U2850 (N_2850,N_2441,N_2065);
or U2851 (N_2851,N_2156,N_2395);
nor U2852 (N_2852,N_2486,N_2138);
and U2853 (N_2853,N_2168,N_2366);
nor U2854 (N_2854,N_2386,N_2249);
nand U2855 (N_2855,N_2006,N_2266);
or U2856 (N_2856,N_2248,N_2481);
nor U2857 (N_2857,N_2325,N_2473);
nand U2858 (N_2858,N_2226,N_2112);
nor U2859 (N_2859,N_2252,N_2081);
or U2860 (N_2860,N_2130,N_2034);
or U2861 (N_2861,N_2042,N_2298);
and U2862 (N_2862,N_2485,N_2237);
nor U2863 (N_2863,N_2385,N_2210);
or U2864 (N_2864,N_2137,N_2293);
nor U2865 (N_2865,N_2058,N_2452);
nand U2866 (N_2866,N_2115,N_2497);
and U2867 (N_2867,N_2048,N_2259);
or U2868 (N_2868,N_2013,N_2241);
and U2869 (N_2869,N_2054,N_2251);
nor U2870 (N_2870,N_2358,N_2030);
and U2871 (N_2871,N_2381,N_2366);
nand U2872 (N_2872,N_2175,N_2413);
nand U2873 (N_2873,N_2136,N_2248);
and U2874 (N_2874,N_2241,N_2200);
or U2875 (N_2875,N_2373,N_2118);
nand U2876 (N_2876,N_2044,N_2429);
nor U2877 (N_2877,N_2049,N_2178);
nand U2878 (N_2878,N_2152,N_2432);
or U2879 (N_2879,N_2405,N_2345);
or U2880 (N_2880,N_2492,N_2392);
nor U2881 (N_2881,N_2039,N_2105);
nor U2882 (N_2882,N_2049,N_2374);
or U2883 (N_2883,N_2435,N_2498);
and U2884 (N_2884,N_2065,N_2403);
nor U2885 (N_2885,N_2499,N_2281);
and U2886 (N_2886,N_2437,N_2077);
nand U2887 (N_2887,N_2198,N_2208);
and U2888 (N_2888,N_2007,N_2292);
or U2889 (N_2889,N_2461,N_2264);
or U2890 (N_2890,N_2493,N_2032);
nor U2891 (N_2891,N_2469,N_2175);
nand U2892 (N_2892,N_2496,N_2339);
or U2893 (N_2893,N_2419,N_2109);
or U2894 (N_2894,N_2119,N_2340);
nor U2895 (N_2895,N_2033,N_2182);
nor U2896 (N_2896,N_2427,N_2238);
nand U2897 (N_2897,N_2243,N_2231);
and U2898 (N_2898,N_2024,N_2118);
nand U2899 (N_2899,N_2258,N_2427);
or U2900 (N_2900,N_2330,N_2398);
or U2901 (N_2901,N_2295,N_2440);
nor U2902 (N_2902,N_2061,N_2445);
nand U2903 (N_2903,N_2332,N_2325);
nor U2904 (N_2904,N_2194,N_2291);
or U2905 (N_2905,N_2284,N_2301);
or U2906 (N_2906,N_2223,N_2297);
or U2907 (N_2907,N_2438,N_2272);
or U2908 (N_2908,N_2433,N_2408);
nand U2909 (N_2909,N_2224,N_2075);
nor U2910 (N_2910,N_2047,N_2139);
nor U2911 (N_2911,N_2118,N_2490);
nand U2912 (N_2912,N_2217,N_2180);
nor U2913 (N_2913,N_2381,N_2321);
and U2914 (N_2914,N_2136,N_2121);
nand U2915 (N_2915,N_2431,N_2315);
and U2916 (N_2916,N_2067,N_2025);
nor U2917 (N_2917,N_2399,N_2327);
and U2918 (N_2918,N_2465,N_2073);
nand U2919 (N_2919,N_2100,N_2355);
and U2920 (N_2920,N_2001,N_2305);
or U2921 (N_2921,N_2254,N_2379);
or U2922 (N_2922,N_2154,N_2409);
nor U2923 (N_2923,N_2346,N_2402);
and U2924 (N_2924,N_2181,N_2169);
and U2925 (N_2925,N_2178,N_2251);
nor U2926 (N_2926,N_2394,N_2431);
nand U2927 (N_2927,N_2485,N_2271);
nor U2928 (N_2928,N_2318,N_2422);
nand U2929 (N_2929,N_2099,N_2032);
and U2930 (N_2930,N_2260,N_2353);
nand U2931 (N_2931,N_2015,N_2487);
nand U2932 (N_2932,N_2331,N_2034);
and U2933 (N_2933,N_2079,N_2327);
and U2934 (N_2934,N_2010,N_2107);
or U2935 (N_2935,N_2422,N_2487);
or U2936 (N_2936,N_2167,N_2023);
and U2937 (N_2937,N_2468,N_2156);
or U2938 (N_2938,N_2141,N_2375);
and U2939 (N_2939,N_2102,N_2288);
and U2940 (N_2940,N_2224,N_2378);
nand U2941 (N_2941,N_2180,N_2107);
and U2942 (N_2942,N_2393,N_2366);
or U2943 (N_2943,N_2157,N_2083);
and U2944 (N_2944,N_2070,N_2075);
or U2945 (N_2945,N_2110,N_2148);
nand U2946 (N_2946,N_2464,N_2408);
and U2947 (N_2947,N_2457,N_2199);
and U2948 (N_2948,N_2237,N_2196);
and U2949 (N_2949,N_2311,N_2009);
nand U2950 (N_2950,N_2152,N_2178);
and U2951 (N_2951,N_2471,N_2035);
nand U2952 (N_2952,N_2256,N_2379);
and U2953 (N_2953,N_2436,N_2182);
or U2954 (N_2954,N_2231,N_2353);
xnor U2955 (N_2955,N_2101,N_2411);
nor U2956 (N_2956,N_2145,N_2137);
and U2957 (N_2957,N_2196,N_2002);
or U2958 (N_2958,N_2149,N_2378);
or U2959 (N_2959,N_2169,N_2211);
or U2960 (N_2960,N_2477,N_2144);
nor U2961 (N_2961,N_2086,N_2481);
and U2962 (N_2962,N_2294,N_2125);
xor U2963 (N_2963,N_2402,N_2327);
or U2964 (N_2964,N_2387,N_2334);
or U2965 (N_2965,N_2071,N_2238);
nor U2966 (N_2966,N_2412,N_2311);
nor U2967 (N_2967,N_2339,N_2347);
nor U2968 (N_2968,N_2341,N_2275);
and U2969 (N_2969,N_2161,N_2470);
or U2970 (N_2970,N_2383,N_2473);
nand U2971 (N_2971,N_2046,N_2241);
or U2972 (N_2972,N_2210,N_2363);
and U2973 (N_2973,N_2082,N_2122);
and U2974 (N_2974,N_2482,N_2442);
and U2975 (N_2975,N_2054,N_2376);
nor U2976 (N_2976,N_2479,N_2163);
and U2977 (N_2977,N_2015,N_2140);
nor U2978 (N_2978,N_2440,N_2086);
nor U2979 (N_2979,N_2436,N_2263);
nor U2980 (N_2980,N_2250,N_2139);
nand U2981 (N_2981,N_2371,N_2283);
nand U2982 (N_2982,N_2150,N_2100);
and U2983 (N_2983,N_2374,N_2067);
nand U2984 (N_2984,N_2238,N_2111);
and U2985 (N_2985,N_2132,N_2448);
nand U2986 (N_2986,N_2061,N_2218);
nand U2987 (N_2987,N_2211,N_2386);
nand U2988 (N_2988,N_2168,N_2494);
and U2989 (N_2989,N_2111,N_2279);
and U2990 (N_2990,N_2179,N_2394);
nor U2991 (N_2991,N_2239,N_2398);
nand U2992 (N_2992,N_2033,N_2408);
or U2993 (N_2993,N_2210,N_2075);
nand U2994 (N_2994,N_2014,N_2253);
or U2995 (N_2995,N_2025,N_2352);
or U2996 (N_2996,N_2084,N_2007);
nand U2997 (N_2997,N_2425,N_2332);
and U2998 (N_2998,N_2196,N_2070);
and U2999 (N_2999,N_2219,N_2013);
or UO_0 (O_0,N_2766,N_2945);
and UO_1 (O_1,N_2750,N_2730);
nor UO_2 (O_2,N_2725,N_2623);
or UO_3 (O_3,N_2701,N_2600);
or UO_4 (O_4,N_2811,N_2867);
nand UO_5 (O_5,N_2972,N_2924);
nor UO_6 (O_6,N_2598,N_2506);
or UO_7 (O_7,N_2836,N_2514);
nor UO_8 (O_8,N_2943,N_2685);
and UO_9 (O_9,N_2752,N_2930);
or UO_10 (O_10,N_2736,N_2641);
or UO_11 (O_11,N_2553,N_2923);
or UO_12 (O_12,N_2662,N_2852);
nand UO_13 (O_13,N_2941,N_2773);
nand UO_14 (O_14,N_2997,N_2619);
nand UO_15 (O_15,N_2861,N_2952);
or UO_16 (O_16,N_2721,N_2599);
and UO_17 (O_17,N_2983,N_2783);
nor UO_18 (O_18,N_2743,N_2869);
nand UO_19 (O_19,N_2785,N_2853);
nand UO_20 (O_20,N_2905,N_2760);
nand UO_21 (O_21,N_2964,N_2695);
and UO_22 (O_22,N_2893,N_2603);
nor UO_23 (O_23,N_2890,N_2799);
or UO_24 (O_24,N_2871,N_2570);
nand UO_25 (O_25,N_2769,N_2966);
nor UO_26 (O_26,N_2948,N_2712);
or UO_27 (O_27,N_2607,N_2805);
and UO_28 (O_28,N_2899,N_2857);
or UO_29 (O_29,N_2779,N_2927);
nand UO_30 (O_30,N_2904,N_2802);
or UO_31 (O_31,N_2568,N_2894);
nor UO_32 (O_32,N_2956,N_2963);
nand UO_33 (O_33,N_2660,N_2593);
and UO_34 (O_34,N_2788,N_2771);
and UO_35 (O_35,N_2957,N_2666);
and UO_36 (O_36,N_2960,N_2965);
nand UO_37 (O_37,N_2870,N_2675);
nor UO_38 (O_38,N_2513,N_2551);
nor UO_39 (O_39,N_2678,N_2765);
or UO_40 (O_40,N_2700,N_2801);
nand UO_41 (O_41,N_2592,N_2579);
nand UO_42 (O_42,N_2648,N_2746);
nor UO_43 (O_43,N_2544,N_2990);
and UO_44 (O_44,N_2611,N_2804);
and UO_45 (O_45,N_2994,N_2714);
or UO_46 (O_46,N_2794,N_2724);
or UO_47 (O_47,N_2552,N_2504);
or UO_48 (O_48,N_2708,N_2680);
nand UO_49 (O_49,N_2572,N_2606);
or UO_50 (O_50,N_2643,N_2699);
nor UO_51 (O_51,N_2885,N_2880);
or UO_52 (O_52,N_2974,N_2989);
nand UO_53 (O_53,N_2955,N_2646);
or UO_54 (O_54,N_2792,N_2732);
nor UO_55 (O_55,N_2764,N_2912);
nand UO_56 (O_56,N_2958,N_2667);
or UO_57 (O_57,N_2873,N_2649);
nand UO_58 (O_58,N_2795,N_2538);
or UO_59 (O_59,N_2531,N_2523);
nand UO_60 (O_60,N_2854,N_2991);
nor UO_61 (O_61,N_2696,N_2775);
or UO_62 (O_62,N_2577,N_2816);
or UO_63 (O_63,N_2718,N_2671);
or UO_64 (O_64,N_2686,N_2637);
or UO_65 (O_65,N_2796,N_2817);
or UO_66 (O_66,N_2605,N_2874);
nand UO_67 (O_67,N_2889,N_2781);
nor UO_68 (O_68,N_2673,N_2876);
nor UO_69 (O_69,N_2507,N_2534);
nor UO_70 (O_70,N_2705,N_2782);
nand UO_71 (O_71,N_2967,N_2809);
and UO_72 (O_72,N_2753,N_2800);
nand UO_73 (O_73,N_2588,N_2501);
nor UO_74 (O_74,N_2982,N_2831);
nor UO_75 (O_75,N_2868,N_2668);
nor UO_76 (O_76,N_2840,N_2936);
nor UO_77 (O_77,N_2672,N_2825);
nand UO_78 (O_78,N_2527,N_2888);
or UO_79 (O_79,N_2689,N_2502);
or UO_80 (O_80,N_2558,N_2741);
or UO_81 (O_81,N_2716,N_2803);
and UO_82 (O_82,N_2535,N_2629);
nor UO_83 (O_83,N_2855,N_2713);
or UO_84 (O_84,N_2729,N_2787);
or UO_85 (O_85,N_2832,N_2995);
and UO_86 (O_86,N_2872,N_2954);
nor UO_87 (O_87,N_2797,N_2949);
nor UO_88 (O_88,N_2862,N_2946);
nor UO_89 (O_89,N_2711,N_2702);
nand UO_90 (O_90,N_2674,N_2710);
nand UO_91 (O_91,N_2933,N_2925);
and UO_92 (O_92,N_2833,N_2758);
or UO_93 (O_93,N_2968,N_2510);
nand UO_94 (O_94,N_2537,N_2574);
and UO_95 (O_95,N_2582,N_2882);
and UO_96 (O_96,N_2772,N_2953);
nand UO_97 (O_97,N_2683,N_2541);
nand UO_98 (O_98,N_2986,N_2652);
nand UO_99 (O_99,N_2661,N_2934);
nor UO_100 (O_100,N_2704,N_2642);
nand UO_101 (O_101,N_2992,N_2812);
or UO_102 (O_102,N_2707,N_2737);
nor UO_103 (O_103,N_2658,N_2546);
nor UO_104 (O_104,N_2891,N_2814);
or UO_105 (O_105,N_2877,N_2723);
and UO_106 (O_106,N_2500,N_2590);
or UO_107 (O_107,N_2980,N_2935);
or UO_108 (O_108,N_2973,N_2848);
and UO_109 (O_109,N_2516,N_2818);
and UO_110 (O_110,N_2971,N_2536);
nand UO_111 (O_111,N_2850,N_2609);
nand UO_112 (O_112,N_2665,N_2914);
xnor UO_113 (O_113,N_2720,N_2977);
nand UO_114 (O_114,N_2647,N_2621);
or UO_115 (O_115,N_2613,N_2910);
and UO_116 (O_116,N_2639,N_2520);
nand UO_117 (O_117,N_2524,N_2521);
nor UO_118 (O_118,N_2940,N_2916);
and UO_119 (O_119,N_2719,N_2896);
nor UO_120 (O_120,N_2778,N_2906);
nor UO_121 (O_121,N_2624,N_2561);
or UO_122 (O_122,N_2847,N_2944);
nor UO_123 (O_123,N_2951,N_2628);
and UO_124 (O_124,N_2728,N_2808);
and UO_125 (O_125,N_2676,N_2790);
nor UO_126 (O_126,N_2756,N_2898);
and UO_127 (O_127,N_2851,N_2557);
or UO_128 (O_128,N_2726,N_2519);
or UO_129 (O_129,N_2841,N_2875);
or UO_130 (O_130,N_2970,N_2822);
and UO_131 (O_131,N_2902,N_2543);
nand UO_132 (O_132,N_2824,N_2597);
or UO_133 (O_133,N_2633,N_2845);
or UO_134 (O_134,N_2610,N_2614);
nor UO_135 (O_135,N_2587,N_2540);
nor UO_136 (O_136,N_2975,N_2566);
nor UO_137 (O_137,N_2921,N_2865);
or UO_138 (O_138,N_2763,N_2976);
and UO_139 (O_139,N_2884,N_2807);
or UO_140 (O_140,N_2657,N_2616);
and UO_141 (O_141,N_2886,N_2757);
or UO_142 (O_142,N_2709,N_2601);
and UO_143 (O_143,N_2767,N_2595);
and UO_144 (O_144,N_2586,N_2813);
xnor UO_145 (O_145,N_2512,N_2669);
nor UO_146 (O_146,N_2937,N_2950);
nand UO_147 (O_147,N_2591,N_2985);
and UO_148 (O_148,N_2670,N_2681);
and UO_149 (O_149,N_2897,N_2585);
nor UO_150 (O_150,N_2618,N_2717);
and UO_151 (O_151,N_2820,N_2735);
nor UO_152 (O_152,N_2694,N_2734);
nand UO_153 (O_153,N_2731,N_2564);
and UO_154 (O_154,N_2858,N_2554);
or UO_155 (O_155,N_2749,N_2575);
nand UO_156 (O_156,N_2917,N_2528);
nand UO_157 (O_157,N_2580,N_2835);
nand UO_158 (O_158,N_2645,N_2838);
nand UO_159 (O_159,N_2703,N_2962);
nor UO_160 (O_160,N_2739,N_2849);
and UO_161 (O_161,N_2644,N_2693);
nand UO_162 (O_162,N_2602,N_2996);
or UO_163 (O_163,N_2526,N_2632);
or UO_164 (O_164,N_2837,N_2761);
nor UO_165 (O_165,N_2748,N_2684);
and UO_166 (O_166,N_2697,N_2786);
nand UO_167 (O_167,N_2987,N_2583);
or UO_168 (O_168,N_2744,N_2682);
nand UO_169 (O_169,N_2550,N_2690);
nor UO_170 (O_170,N_2895,N_2505);
or UO_171 (O_171,N_2545,N_2698);
nand UO_172 (O_172,N_2908,N_2863);
or UO_173 (O_173,N_2830,N_2692);
or UO_174 (O_174,N_2548,N_2784);
nand UO_175 (O_175,N_2573,N_2920);
nor UO_176 (O_176,N_2777,N_2834);
and UO_177 (O_177,N_2864,N_2636);
and UO_178 (O_178,N_2608,N_2856);
and UO_179 (O_179,N_2612,N_2768);
nor UO_180 (O_180,N_2878,N_2843);
nor UO_181 (O_181,N_2620,N_2659);
or UO_182 (O_182,N_2939,N_2740);
and UO_183 (O_183,N_2776,N_2615);
nor UO_184 (O_184,N_2525,N_2511);
or UO_185 (O_185,N_2542,N_2979);
nor UO_186 (O_186,N_2774,N_2576);
or UO_187 (O_187,N_2687,N_2745);
or UO_188 (O_188,N_2518,N_2581);
and UO_189 (O_189,N_2981,N_2823);
nor UO_190 (O_190,N_2655,N_2562);
or UO_191 (O_191,N_2931,N_2663);
nor UO_192 (O_192,N_2998,N_2547);
nor UO_193 (O_193,N_2625,N_2738);
or UO_194 (O_194,N_2630,N_2900);
nand UO_195 (O_195,N_2529,N_2829);
nor UO_196 (O_196,N_2650,N_2879);
or UO_197 (O_197,N_2715,N_2656);
nor UO_198 (O_198,N_2622,N_2881);
and UO_199 (O_199,N_2815,N_2751);
or UO_200 (O_200,N_2789,N_2922);
nand UO_201 (O_201,N_2634,N_2806);
xor UO_202 (O_202,N_2942,N_2887);
nor UO_203 (O_203,N_2827,N_2727);
and UO_204 (O_204,N_2503,N_2780);
nor UO_205 (O_205,N_2993,N_2560);
nand UO_206 (O_206,N_2919,N_2584);
nand UO_207 (O_207,N_2604,N_2640);
or UO_208 (O_208,N_2754,N_2509);
nand UO_209 (O_209,N_2999,N_2928);
nand UO_210 (O_210,N_2932,N_2688);
or UO_211 (O_211,N_2569,N_2762);
and UO_212 (O_212,N_2571,N_2839);
or UO_213 (O_213,N_2860,N_2892);
and UO_214 (O_214,N_2929,N_2901);
nor UO_215 (O_215,N_2617,N_2810);
or UO_216 (O_216,N_2664,N_2508);
nor UO_217 (O_217,N_2926,N_2755);
or UO_218 (O_218,N_2578,N_2747);
nand UO_219 (O_219,N_2915,N_2677);
and UO_220 (O_220,N_2883,N_2742);
nand UO_221 (O_221,N_2626,N_2959);
and UO_222 (O_222,N_2793,N_2907);
nand UO_223 (O_223,N_2631,N_2589);
and UO_224 (O_224,N_2969,N_2826);
and UO_225 (O_225,N_2654,N_2961);
and UO_226 (O_226,N_2828,N_2635);
nor UO_227 (O_227,N_2653,N_2563);
nand UO_228 (O_228,N_2549,N_2791);
and UO_229 (O_229,N_2866,N_2798);
nor UO_230 (O_230,N_2559,N_2532);
nor UO_231 (O_231,N_2567,N_2596);
nor UO_232 (O_232,N_2938,N_2722);
and UO_233 (O_233,N_2842,N_2947);
or UO_234 (O_234,N_2555,N_2903);
and UO_235 (O_235,N_2821,N_2691);
and UO_236 (O_236,N_2988,N_2522);
nand UO_237 (O_237,N_2517,N_2539);
and UO_238 (O_238,N_2556,N_2759);
nand UO_239 (O_239,N_2911,N_2733);
or UO_240 (O_240,N_2770,N_2565);
nand UO_241 (O_241,N_2594,N_2638);
or UO_242 (O_242,N_2844,N_2627);
or UO_243 (O_243,N_2918,N_2533);
and UO_244 (O_244,N_2859,N_2984);
or UO_245 (O_245,N_2846,N_2978);
or UO_246 (O_246,N_2515,N_2651);
nand UO_247 (O_247,N_2913,N_2706);
and UO_248 (O_248,N_2909,N_2530);
or UO_249 (O_249,N_2819,N_2679);
or UO_250 (O_250,N_2723,N_2953);
and UO_251 (O_251,N_2984,N_2585);
nor UO_252 (O_252,N_2647,N_2534);
nand UO_253 (O_253,N_2585,N_2987);
nor UO_254 (O_254,N_2712,N_2676);
and UO_255 (O_255,N_2891,N_2785);
nor UO_256 (O_256,N_2834,N_2952);
or UO_257 (O_257,N_2546,N_2780);
nor UO_258 (O_258,N_2510,N_2508);
and UO_259 (O_259,N_2708,N_2918);
nor UO_260 (O_260,N_2668,N_2638);
nand UO_261 (O_261,N_2936,N_2503);
and UO_262 (O_262,N_2905,N_2606);
nor UO_263 (O_263,N_2791,N_2723);
nand UO_264 (O_264,N_2708,N_2663);
and UO_265 (O_265,N_2806,N_2857);
nand UO_266 (O_266,N_2832,N_2698);
nand UO_267 (O_267,N_2805,N_2803);
nor UO_268 (O_268,N_2511,N_2567);
and UO_269 (O_269,N_2880,N_2665);
nand UO_270 (O_270,N_2742,N_2682);
nand UO_271 (O_271,N_2679,N_2873);
or UO_272 (O_272,N_2533,N_2632);
or UO_273 (O_273,N_2991,N_2897);
or UO_274 (O_274,N_2880,N_2836);
nand UO_275 (O_275,N_2635,N_2554);
or UO_276 (O_276,N_2587,N_2837);
and UO_277 (O_277,N_2755,N_2659);
nand UO_278 (O_278,N_2926,N_2898);
or UO_279 (O_279,N_2880,N_2573);
nor UO_280 (O_280,N_2818,N_2677);
or UO_281 (O_281,N_2930,N_2524);
nor UO_282 (O_282,N_2644,N_2529);
nand UO_283 (O_283,N_2501,N_2656);
nor UO_284 (O_284,N_2899,N_2535);
and UO_285 (O_285,N_2784,N_2568);
or UO_286 (O_286,N_2509,N_2849);
nand UO_287 (O_287,N_2987,N_2855);
xnor UO_288 (O_288,N_2669,N_2636);
nand UO_289 (O_289,N_2943,N_2927);
or UO_290 (O_290,N_2799,N_2885);
or UO_291 (O_291,N_2533,N_2932);
and UO_292 (O_292,N_2589,N_2789);
or UO_293 (O_293,N_2947,N_2702);
or UO_294 (O_294,N_2789,N_2988);
or UO_295 (O_295,N_2560,N_2860);
and UO_296 (O_296,N_2747,N_2518);
or UO_297 (O_297,N_2827,N_2567);
nor UO_298 (O_298,N_2581,N_2966);
nand UO_299 (O_299,N_2926,N_2749);
and UO_300 (O_300,N_2920,N_2965);
nand UO_301 (O_301,N_2583,N_2985);
nand UO_302 (O_302,N_2613,N_2733);
or UO_303 (O_303,N_2917,N_2701);
nand UO_304 (O_304,N_2951,N_2708);
nand UO_305 (O_305,N_2766,N_2841);
and UO_306 (O_306,N_2889,N_2722);
and UO_307 (O_307,N_2591,N_2710);
or UO_308 (O_308,N_2612,N_2605);
nor UO_309 (O_309,N_2505,N_2856);
and UO_310 (O_310,N_2967,N_2555);
and UO_311 (O_311,N_2965,N_2528);
and UO_312 (O_312,N_2849,N_2588);
nor UO_313 (O_313,N_2779,N_2784);
or UO_314 (O_314,N_2981,N_2523);
and UO_315 (O_315,N_2898,N_2630);
nor UO_316 (O_316,N_2974,N_2616);
or UO_317 (O_317,N_2775,N_2818);
and UO_318 (O_318,N_2683,N_2791);
nor UO_319 (O_319,N_2985,N_2945);
nand UO_320 (O_320,N_2855,N_2743);
or UO_321 (O_321,N_2898,N_2533);
nand UO_322 (O_322,N_2584,N_2764);
and UO_323 (O_323,N_2968,N_2819);
nor UO_324 (O_324,N_2700,N_2711);
and UO_325 (O_325,N_2841,N_2550);
nand UO_326 (O_326,N_2727,N_2868);
nor UO_327 (O_327,N_2553,N_2824);
or UO_328 (O_328,N_2747,N_2828);
and UO_329 (O_329,N_2884,N_2914);
or UO_330 (O_330,N_2529,N_2970);
nand UO_331 (O_331,N_2796,N_2843);
or UO_332 (O_332,N_2822,N_2567);
or UO_333 (O_333,N_2772,N_2879);
nand UO_334 (O_334,N_2895,N_2917);
and UO_335 (O_335,N_2817,N_2626);
or UO_336 (O_336,N_2525,N_2829);
nand UO_337 (O_337,N_2562,N_2539);
nand UO_338 (O_338,N_2862,N_2552);
or UO_339 (O_339,N_2830,N_2570);
xor UO_340 (O_340,N_2538,N_2851);
nor UO_341 (O_341,N_2580,N_2542);
nand UO_342 (O_342,N_2643,N_2626);
or UO_343 (O_343,N_2775,N_2568);
nand UO_344 (O_344,N_2649,N_2656);
or UO_345 (O_345,N_2599,N_2924);
nor UO_346 (O_346,N_2529,N_2609);
nor UO_347 (O_347,N_2852,N_2982);
or UO_348 (O_348,N_2595,N_2838);
nor UO_349 (O_349,N_2699,N_2587);
nor UO_350 (O_350,N_2733,N_2698);
nor UO_351 (O_351,N_2830,N_2920);
nand UO_352 (O_352,N_2857,N_2902);
nor UO_353 (O_353,N_2660,N_2813);
nor UO_354 (O_354,N_2856,N_2889);
and UO_355 (O_355,N_2804,N_2733);
nor UO_356 (O_356,N_2564,N_2645);
or UO_357 (O_357,N_2716,N_2507);
nor UO_358 (O_358,N_2779,N_2614);
nand UO_359 (O_359,N_2583,N_2709);
and UO_360 (O_360,N_2952,N_2758);
or UO_361 (O_361,N_2865,N_2922);
and UO_362 (O_362,N_2722,N_2566);
nand UO_363 (O_363,N_2672,N_2878);
or UO_364 (O_364,N_2597,N_2780);
or UO_365 (O_365,N_2652,N_2857);
nor UO_366 (O_366,N_2759,N_2911);
nor UO_367 (O_367,N_2613,N_2622);
and UO_368 (O_368,N_2934,N_2833);
nor UO_369 (O_369,N_2716,N_2714);
and UO_370 (O_370,N_2522,N_2893);
and UO_371 (O_371,N_2703,N_2780);
or UO_372 (O_372,N_2792,N_2523);
and UO_373 (O_373,N_2675,N_2970);
and UO_374 (O_374,N_2870,N_2637);
nand UO_375 (O_375,N_2632,N_2977);
nand UO_376 (O_376,N_2686,N_2820);
or UO_377 (O_377,N_2524,N_2963);
and UO_378 (O_378,N_2631,N_2533);
or UO_379 (O_379,N_2963,N_2941);
and UO_380 (O_380,N_2960,N_2850);
or UO_381 (O_381,N_2951,N_2952);
nor UO_382 (O_382,N_2720,N_2539);
and UO_383 (O_383,N_2862,N_2539);
and UO_384 (O_384,N_2665,N_2989);
and UO_385 (O_385,N_2911,N_2632);
nand UO_386 (O_386,N_2650,N_2682);
nor UO_387 (O_387,N_2746,N_2722);
nand UO_388 (O_388,N_2620,N_2928);
nand UO_389 (O_389,N_2800,N_2524);
or UO_390 (O_390,N_2970,N_2636);
nor UO_391 (O_391,N_2802,N_2647);
or UO_392 (O_392,N_2901,N_2840);
nor UO_393 (O_393,N_2663,N_2991);
and UO_394 (O_394,N_2878,N_2569);
nor UO_395 (O_395,N_2834,N_2790);
nor UO_396 (O_396,N_2670,N_2544);
nor UO_397 (O_397,N_2807,N_2990);
and UO_398 (O_398,N_2739,N_2636);
or UO_399 (O_399,N_2919,N_2897);
and UO_400 (O_400,N_2530,N_2991);
nor UO_401 (O_401,N_2964,N_2811);
nand UO_402 (O_402,N_2764,N_2629);
nand UO_403 (O_403,N_2889,N_2635);
nand UO_404 (O_404,N_2574,N_2669);
and UO_405 (O_405,N_2871,N_2588);
nor UO_406 (O_406,N_2666,N_2862);
and UO_407 (O_407,N_2627,N_2886);
and UO_408 (O_408,N_2607,N_2511);
nand UO_409 (O_409,N_2694,N_2810);
nand UO_410 (O_410,N_2986,N_2852);
and UO_411 (O_411,N_2841,N_2914);
and UO_412 (O_412,N_2713,N_2678);
or UO_413 (O_413,N_2874,N_2765);
and UO_414 (O_414,N_2738,N_2631);
and UO_415 (O_415,N_2679,N_2848);
nand UO_416 (O_416,N_2968,N_2767);
or UO_417 (O_417,N_2645,N_2959);
nor UO_418 (O_418,N_2638,N_2659);
or UO_419 (O_419,N_2587,N_2801);
and UO_420 (O_420,N_2622,N_2905);
nor UO_421 (O_421,N_2871,N_2730);
and UO_422 (O_422,N_2807,N_2613);
nand UO_423 (O_423,N_2777,N_2626);
nor UO_424 (O_424,N_2791,N_2697);
or UO_425 (O_425,N_2827,N_2735);
nand UO_426 (O_426,N_2684,N_2810);
xnor UO_427 (O_427,N_2668,N_2667);
or UO_428 (O_428,N_2665,N_2904);
nand UO_429 (O_429,N_2584,N_2724);
nor UO_430 (O_430,N_2536,N_2610);
nand UO_431 (O_431,N_2844,N_2737);
or UO_432 (O_432,N_2872,N_2699);
nor UO_433 (O_433,N_2772,N_2848);
nand UO_434 (O_434,N_2505,N_2745);
nor UO_435 (O_435,N_2525,N_2893);
and UO_436 (O_436,N_2582,N_2866);
and UO_437 (O_437,N_2639,N_2551);
nor UO_438 (O_438,N_2934,N_2818);
nand UO_439 (O_439,N_2933,N_2941);
nand UO_440 (O_440,N_2515,N_2852);
and UO_441 (O_441,N_2554,N_2895);
and UO_442 (O_442,N_2953,N_2846);
nor UO_443 (O_443,N_2766,N_2985);
and UO_444 (O_444,N_2650,N_2721);
or UO_445 (O_445,N_2549,N_2912);
nand UO_446 (O_446,N_2859,N_2980);
nand UO_447 (O_447,N_2675,N_2974);
nand UO_448 (O_448,N_2813,N_2564);
nand UO_449 (O_449,N_2882,N_2962);
nand UO_450 (O_450,N_2576,N_2772);
nand UO_451 (O_451,N_2603,N_2963);
nand UO_452 (O_452,N_2593,N_2883);
or UO_453 (O_453,N_2640,N_2986);
or UO_454 (O_454,N_2716,N_2912);
nor UO_455 (O_455,N_2915,N_2990);
nor UO_456 (O_456,N_2782,N_2656);
nor UO_457 (O_457,N_2832,N_2983);
and UO_458 (O_458,N_2990,N_2621);
nand UO_459 (O_459,N_2746,N_2643);
and UO_460 (O_460,N_2977,N_2589);
or UO_461 (O_461,N_2545,N_2743);
and UO_462 (O_462,N_2748,N_2772);
and UO_463 (O_463,N_2720,N_2749);
and UO_464 (O_464,N_2871,N_2924);
or UO_465 (O_465,N_2712,N_2706);
xnor UO_466 (O_466,N_2641,N_2874);
or UO_467 (O_467,N_2556,N_2613);
or UO_468 (O_468,N_2816,N_2639);
and UO_469 (O_469,N_2592,N_2899);
nand UO_470 (O_470,N_2766,N_2948);
xor UO_471 (O_471,N_2507,N_2912);
nand UO_472 (O_472,N_2543,N_2923);
or UO_473 (O_473,N_2741,N_2511);
nand UO_474 (O_474,N_2933,N_2529);
nor UO_475 (O_475,N_2660,N_2800);
nand UO_476 (O_476,N_2505,N_2527);
nand UO_477 (O_477,N_2937,N_2903);
nor UO_478 (O_478,N_2625,N_2926);
or UO_479 (O_479,N_2704,N_2699);
nor UO_480 (O_480,N_2775,N_2628);
or UO_481 (O_481,N_2982,N_2954);
nor UO_482 (O_482,N_2739,N_2592);
or UO_483 (O_483,N_2705,N_2807);
nor UO_484 (O_484,N_2731,N_2544);
nand UO_485 (O_485,N_2887,N_2899);
nor UO_486 (O_486,N_2959,N_2594);
and UO_487 (O_487,N_2597,N_2857);
nand UO_488 (O_488,N_2606,N_2854);
or UO_489 (O_489,N_2602,N_2895);
and UO_490 (O_490,N_2665,N_2734);
nor UO_491 (O_491,N_2856,N_2663);
or UO_492 (O_492,N_2708,N_2619);
or UO_493 (O_493,N_2753,N_2739);
and UO_494 (O_494,N_2677,N_2953);
and UO_495 (O_495,N_2629,N_2680);
or UO_496 (O_496,N_2786,N_2912);
xnor UO_497 (O_497,N_2988,N_2670);
nor UO_498 (O_498,N_2717,N_2791);
nor UO_499 (O_499,N_2906,N_2706);
endmodule