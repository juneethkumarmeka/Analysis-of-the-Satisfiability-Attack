module basic_1000_10000_1500_2_levels_2xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5006,N_5007,N_5013,N_5014,N_5016,N_5017,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5033,N_5040,N_5041,N_5043,N_5046,N_5047,N_5048,N_5049,N_5051,N_5052,N_5053,N_5057,N_5058,N_5060,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5070,N_5074,N_5082,N_5083,N_5086,N_5087,N_5090,N_5092,N_5094,N_5095,N_5096,N_5097,N_5098,N_5101,N_5102,N_5106,N_5107,N_5108,N_5110,N_5111,N_5112,N_5113,N_5116,N_5117,N_5118,N_5119,N_5121,N_5124,N_5125,N_5126,N_5127,N_5129,N_5131,N_5135,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5149,N_5150,N_5151,N_5152,N_5153,N_5155,N_5158,N_5160,N_5161,N_5164,N_5166,N_5170,N_5172,N_5173,N_5176,N_5177,N_5179,N_5181,N_5182,N_5184,N_5185,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5196,N_5199,N_5200,N_5202,N_5206,N_5208,N_5209,N_5213,N_5215,N_5217,N_5219,N_5220,N_5222,N_5224,N_5227,N_5229,N_5230,N_5231,N_5232,N_5234,N_5236,N_5237,N_5238,N_5239,N_5240,N_5244,N_5246,N_5248,N_5250,N_5251,N_5252,N_5253,N_5255,N_5256,N_5257,N_5259,N_5260,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5274,N_5277,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5287,N_5288,N_5290,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5301,N_5303,N_5304,N_5305,N_5307,N_5308,N_5310,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5322,N_5323,N_5326,N_5327,N_5329,N_5330,N_5334,N_5335,N_5336,N_5337,N_5338,N_5340,N_5342,N_5345,N_5346,N_5347,N_5348,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5358,N_5359,N_5361,N_5363,N_5364,N_5365,N_5366,N_5368,N_5369,N_5370,N_5373,N_5375,N_5377,N_5380,N_5381,N_5383,N_5384,N_5385,N_5387,N_5388,N_5389,N_5390,N_5394,N_5395,N_5396,N_5398,N_5399,N_5400,N_5402,N_5405,N_5406,N_5407,N_5409,N_5410,N_5414,N_5415,N_5420,N_5421,N_5423,N_5424,N_5427,N_5429,N_5431,N_5433,N_5435,N_5436,N_5440,N_5443,N_5444,N_5445,N_5447,N_5449,N_5450,N_5452,N_5453,N_5454,N_5456,N_5458,N_5459,N_5461,N_5462,N_5463,N_5464,N_5466,N_5467,N_5469,N_5472,N_5473,N_5474,N_5476,N_5479,N_5482,N_5485,N_5487,N_5488,N_5489,N_5490,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5501,N_5502,N_5504,N_5506,N_5508,N_5509,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5523,N_5524,N_5526,N_5527,N_5529,N_5531,N_5534,N_5535,N_5536,N_5537,N_5539,N_5541,N_5542,N_5546,N_5552,N_5554,N_5558,N_5559,N_5560,N_5561,N_5563,N_5564,N_5566,N_5568,N_5571,N_5572,N_5573,N_5574,N_5576,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5586,N_5587,N_5588,N_5590,N_5591,N_5592,N_5594,N_5595,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5606,N_5608,N_5609,N_5613,N_5614,N_5615,N_5616,N_5617,N_5622,N_5624,N_5625,N_5628,N_5629,N_5630,N_5631,N_5633,N_5634,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5645,N_5646,N_5647,N_5649,N_5651,N_5652,N_5653,N_5655,N_5656,N_5657,N_5660,N_5661,N_5663,N_5664,N_5666,N_5667,N_5668,N_5670,N_5671,N_5675,N_5676,N_5679,N_5680,N_5681,N_5682,N_5683,N_5686,N_5687,N_5688,N_5690,N_5691,N_5692,N_5693,N_5695,N_5699,N_5701,N_5702,N_5703,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5716,N_5719,N_5721,N_5722,N_5724,N_5725,N_5726,N_5727,N_5728,N_5731,N_5732,N_5733,N_5735,N_5736,N_5737,N_5739,N_5741,N_5742,N_5744,N_5749,N_5751,N_5753,N_5755,N_5756,N_5757,N_5759,N_5760,N_5761,N_5763,N_5766,N_5767,N_5768,N_5769,N_5770,N_5772,N_5773,N_5777,N_5778,N_5781,N_5783,N_5784,N_5785,N_5787,N_5788,N_5790,N_5791,N_5792,N_5797,N_5799,N_5801,N_5802,N_5804,N_5805,N_5806,N_5807,N_5810,N_5812,N_5813,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5824,N_5827,N_5830,N_5834,N_5838,N_5840,N_5841,N_5842,N_5843,N_5844,N_5848,N_5849,N_5851,N_5852,N_5853,N_5855,N_5857,N_5858,N_5859,N_5861,N_5862,N_5866,N_5867,N_5869,N_5870,N_5872,N_5875,N_5876,N_5877,N_5878,N_5880,N_5882,N_5886,N_5887,N_5889,N_5891,N_5892,N_5893,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5907,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5919,N_5920,N_5921,N_5922,N_5923,N_5925,N_5926,N_5927,N_5929,N_5930,N_5931,N_5932,N_5934,N_5935,N_5937,N_5938,N_5941,N_5942,N_5943,N_5945,N_5947,N_5948,N_5949,N_5951,N_5952,N_5954,N_5956,N_5957,N_5958,N_5959,N_5962,N_5963,N_5964,N_5965,N_5966,N_5969,N_5970,N_5975,N_5977,N_5978,N_5980,N_5981,N_5987,N_5988,N_5989,N_5990,N_5991,N_5993,N_5994,N_5996,N_5997,N_5998,N_6000,N_6001,N_6002,N_6003,N_6005,N_6007,N_6010,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6024,N_6029,N_6031,N_6032,N_6033,N_6035,N_6037,N_6038,N_6041,N_6042,N_6043,N_6045,N_6046,N_6047,N_6048,N_6049,N_6051,N_6052,N_6054,N_6056,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6068,N_6069,N_6071,N_6072,N_6073,N_6074,N_6075,N_6077,N_6079,N_6084,N_6086,N_6087,N_6088,N_6090,N_6091,N_6092,N_6094,N_6096,N_6097,N_6098,N_6102,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6115,N_6116,N_6118,N_6120,N_6121,N_6122,N_6123,N_6124,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6141,N_6142,N_6144,N_6146,N_6147,N_6148,N_6149,N_6151,N_6155,N_6157,N_6158,N_6159,N_6161,N_6162,N_6166,N_6167,N_6169,N_6170,N_6171,N_6173,N_6177,N_6181,N_6184,N_6186,N_6188,N_6189,N_6191,N_6195,N_6196,N_6198,N_6199,N_6200,N_6201,N_6202,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6213,N_6215,N_6216,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6229,N_6231,N_6232,N_6235,N_6236,N_6237,N_6238,N_6242,N_6243,N_6244,N_6246,N_6247,N_6248,N_6250,N_6251,N_6252,N_6256,N_6257,N_6258,N_6261,N_6262,N_6266,N_6267,N_6268,N_6270,N_6271,N_6274,N_6275,N_6276,N_6277,N_6279,N_6280,N_6281,N_6286,N_6290,N_6292,N_6293,N_6294,N_6295,N_6296,N_6298,N_6299,N_6302,N_6303,N_6305,N_6307,N_6310,N_6311,N_6313,N_6315,N_6318,N_6319,N_6320,N_6324,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6334,N_6335,N_6336,N_6337,N_6338,N_6345,N_6346,N_6347,N_6348,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6358,N_6359,N_6361,N_6362,N_6363,N_6366,N_6369,N_6370,N_6373,N_6374,N_6375,N_6376,N_6377,N_6379,N_6381,N_6382,N_6383,N_6384,N_6385,N_6388,N_6389,N_6390,N_6392,N_6394,N_6395,N_6397,N_6398,N_6399,N_6401,N_6404,N_6405,N_6406,N_6407,N_6410,N_6412,N_6415,N_6416,N_6417,N_6419,N_6420,N_6422,N_6423,N_6426,N_6429,N_6431,N_6434,N_6435,N_6438,N_6440,N_6441,N_6442,N_6444,N_6447,N_6449,N_6450,N_6453,N_6454,N_6456,N_6458,N_6460,N_6461,N_6462,N_6463,N_6466,N_6470,N_6471,N_6472,N_6477,N_6479,N_6481,N_6482,N_6485,N_6486,N_6487,N_6488,N_6490,N_6491,N_6492,N_6493,N_6496,N_6498,N_6499,N_6501,N_6505,N_6507,N_6508,N_6511,N_6512,N_6516,N_6517,N_6518,N_6523,N_6526,N_6528,N_6529,N_6530,N_6532,N_6534,N_6536,N_6537,N_6539,N_6541,N_6543,N_6545,N_6547,N_6548,N_6549,N_6550,N_6553,N_6554,N_6556,N_6557,N_6558,N_6559,N_6560,N_6562,N_6563,N_6565,N_6566,N_6568,N_6569,N_6572,N_6573,N_6574,N_6575,N_6577,N_6585,N_6586,N_6588,N_6590,N_6591,N_6593,N_6595,N_6596,N_6600,N_6601,N_6602,N_6604,N_6605,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6621,N_6622,N_6624,N_6625,N_6627,N_6628,N_6630,N_6632,N_6633,N_6634,N_6635,N_6637,N_6638,N_6641,N_6643,N_6644,N_6645,N_6646,N_6647,N_6650,N_6651,N_6652,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6662,N_6664,N_6669,N_6672,N_6673,N_6674,N_6677,N_6679,N_6683,N_6685,N_6686,N_6687,N_6689,N_6691,N_6692,N_6695,N_6697,N_6698,N_6699,N_6700,N_6703,N_6706,N_6707,N_6708,N_6709,N_6711,N_6713,N_6714,N_6716,N_6717,N_6718,N_6719,N_6721,N_6724,N_6725,N_6726,N_6727,N_6728,N_6733,N_6734,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6746,N_6747,N_6751,N_6752,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6773,N_6774,N_6777,N_6779,N_6780,N_6784,N_6787,N_6789,N_6790,N_6791,N_6792,N_6793,N_6795,N_6796,N_6797,N_6800,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6812,N_6814,N_6815,N_6816,N_6817,N_6818,N_6820,N_6821,N_6822,N_6825,N_6826,N_6829,N_6830,N_6831,N_6832,N_6833,N_6836,N_6838,N_6841,N_6842,N_6846,N_6848,N_6851,N_6852,N_6854,N_6855,N_6857,N_6858,N_6859,N_6860,N_6866,N_6868,N_6870,N_6871,N_6874,N_6877,N_6880,N_6884,N_6885,N_6886,N_6889,N_6891,N_6892,N_6895,N_6897,N_6901,N_6902,N_6907,N_6913,N_6915,N_6916,N_6917,N_6918,N_6921,N_6923,N_6926,N_6930,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6941,N_6942,N_6944,N_6945,N_6947,N_6949,N_6951,N_6952,N_6953,N_6954,N_6955,N_6958,N_6959,N_6962,N_6967,N_6968,N_6969,N_6970,N_6976,N_6978,N_6981,N_6982,N_6984,N_6987,N_6988,N_6989,N_6990,N_6991,N_6993,N_6994,N_6996,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7006,N_7009,N_7010,N_7011,N_7012,N_7015,N_7018,N_7019,N_7020,N_7021,N_7022,N_7025,N_7027,N_7028,N_7029,N_7031,N_7033,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7042,N_7045,N_7046,N_7049,N_7050,N_7052,N_7053,N_7055,N_7056,N_7060,N_7061,N_7063,N_7064,N_7067,N_7068,N_7069,N_7075,N_7076,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7086,N_7087,N_7088,N_7090,N_7091,N_7092,N_7093,N_7094,N_7096,N_7099,N_7101,N_7102,N_7103,N_7104,N_7107,N_7110,N_7113,N_7115,N_7116,N_7119,N_7120,N_7126,N_7127,N_7131,N_7133,N_7134,N_7136,N_7137,N_7140,N_7141,N_7142,N_7143,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7163,N_7164,N_7165,N_7166,N_7168,N_7169,N_7172,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7184,N_7185,N_7186,N_7187,N_7189,N_7190,N_7193,N_7194,N_7195,N_7196,N_7198,N_7199,N_7200,N_7203,N_7205,N_7207,N_7208,N_7209,N_7210,N_7213,N_7215,N_7216,N_7217,N_7219,N_7220,N_7222,N_7224,N_7225,N_7226,N_7227,N_7228,N_7230,N_7231,N_7235,N_7236,N_7240,N_7241,N_7243,N_7244,N_7246,N_7249,N_7251,N_7252,N_7253,N_7254,N_7257,N_7260,N_7262,N_7264,N_7265,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7276,N_7278,N_7280,N_7281,N_7282,N_7283,N_7284,N_7287,N_7288,N_7289,N_7292,N_7294,N_7295,N_7297,N_7298,N_7299,N_7301,N_7303,N_7305,N_7308,N_7309,N_7311,N_7313,N_7314,N_7315,N_7319,N_7320,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7329,N_7333,N_7334,N_7336,N_7337,N_7338,N_7341,N_7344,N_7346,N_7348,N_7351,N_7353,N_7354,N_7355,N_7356,N_7358,N_7360,N_7361,N_7363,N_7364,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7394,N_7395,N_7397,N_7398,N_7399,N_7400,N_7402,N_7403,N_7404,N_7407,N_7408,N_7411,N_7412,N_7414,N_7416,N_7419,N_7420,N_7421,N_7422,N_7424,N_7426,N_7429,N_7430,N_7431,N_7432,N_7433,N_7435,N_7436,N_7438,N_7440,N_7443,N_7445,N_7446,N_7448,N_7450,N_7451,N_7452,N_7454,N_7455,N_7456,N_7458,N_7459,N_7463,N_7464,N_7466,N_7468,N_7469,N_7474,N_7475,N_7478,N_7479,N_7480,N_7483,N_7487,N_7490,N_7491,N_7492,N_7495,N_7499,N_7500,N_7503,N_7504,N_7505,N_7508,N_7509,N_7513,N_7514,N_7515,N_7518,N_7520,N_7521,N_7524,N_7525,N_7527,N_7528,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7537,N_7541,N_7542,N_7544,N_7547,N_7552,N_7553,N_7556,N_7557,N_7560,N_7562,N_7564,N_7566,N_7567,N_7568,N_7569,N_7571,N_7577,N_7579,N_7580,N_7581,N_7582,N_7584,N_7586,N_7587,N_7591,N_7592,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7603,N_7606,N_7608,N_7609,N_7612,N_7615,N_7616,N_7621,N_7623,N_7624,N_7626,N_7627,N_7632,N_7633,N_7634,N_7635,N_7637,N_7638,N_7639,N_7640,N_7644,N_7647,N_7651,N_7652,N_7653,N_7654,N_7655,N_7659,N_7662,N_7663,N_7666,N_7667,N_7668,N_7669,N_7671,N_7672,N_7673,N_7676,N_7678,N_7679,N_7681,N_7682,N_7684,N_7685,N_7687,N_7694,N_7696,N_7698,N_7700,N_7702,N_7703,N_7706,N_7708,N_7710,N_7712,N_7719,N_7720,N_7722,N_7723,N_7724,N_7725,N_7729,N_7731,N_7735,N_7737,N_7739,N_7742,N_7743,N_7746,N_7748,N_7749,N_7750,N_7751,N_7752,N_7755,N_7756,N_7757,N_7758,N_7760,N_7764,N_7767,N_7768,N_7770,N_7771,N_7772,N_7774,N_7776,N_7778,N_7779,N_7780,N_7783,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7793,N_7794,N_7796,N_7797,N_7799,N_7800,N_7801,N_7803,N_7807,N_7808,N_7809,N_7810,N_7813,N_7815,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7824,N_7825,N_7828,N_7832,N_7833,N_7836,N_7837,N_7841,N_7842,N_7843,N_7845,N_7846,N_7847,N_7849,N_7851,N_7855,N_7858,N_7859,N_7860,N_7861,N_7862,N_7865,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7876,N_7877,N_7878,N_7880,N_7881,N_7882,N_7883,N_7885,N_7886,N_7888,N_7889,N_7893,N_7895,N_7897,N_7898,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7912,N_7913,N_7915,N_7917,N_7918,N_7919,N_7920,N_7921,N_7924,N_7925,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7937,N_7938,N_7940,N_7945,N_7946,N_7947,N_7948,N_7949,N_7951,N_7952,N_7953,N_7956,N_7957,N_7958,N_7959,N_7960,N_7962,N_7963,N_7964,N_7965,N_7968,N_7971,N_7975,N_7976,N_7977,N_7978,N_7980,N_7982,N_7984,N_7985,N_7987,N_7991,N_7995,N_7997,N_7999,N_8000,N_8001,N_8003,N_8004,N_8006,N_8008,N_8009,N_8011,N_8013,N_8014,N_8018,N_8020,N_8022,N_8024,N_8025,N_8027,N_8028,N_8032,N_8033,N_8034,N_8037,N_8039,N_8040,N_8041,N_8045,N_8046,N_8048,N_8049,N_8051,N_8054,N_8055,N_8056,N_8058,N_8059,N_8060,N_8064,N_8065,N_8070,N_8073,N_8074,N_8075,N_8076,N_8080,N_8081,N_8082,N_8084,N_8087,N_8088,N_8089,N_8090,N_8093,N_8094,N_8095,N_8096,N_8097,N_8099,N_8100,N_8101,N_8102,N_8103,N_8106,N_8107,N_8108,N_8110,N_8111,N_8115,N_8117,N_8119,N_8121,N_8122,N_8124,N_8125,N_8126,N_8128,N_8130,N_8131,N_8132,N_8134,N_8135,N_8136,N_8141,N_8142,N_8143,N_8144,N_8146,N_8147,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8156,N_8157,N_8158,N_8160,N_8161,N_8162,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8171,N_8172,N_8174,N_8175,N_8178,N_8179,N_8180,N_8181,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8190,N_8191,N_8192,N_8194,N_8196,N_8199,N_8201,N_8202,N_8204,N_8205,N_8206,N_8208,N_8209,N_8210,N_8211,N_8213,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8223,N_8224,N_8225,N_8227,N_8232,N_8234,N_8235,N_8236,N_8238,N_8239,N_8240,N_8242,N_8245,N_8246,N_8250,N_8251,N_8254,N_8256,N_8259,N_8261,N_8262,N_8263,N_8264,N_8267,N_8269,N_8270,N_8271,N_8272,N_8274,N_8275,N_8276,N_8283,N_8284,N_8285,N_8287,N_8292,N_8293,N_8294,N_8296,N_8297,N_8298,N_8300,N_8301,N_8302,N_8303,N_8304,N_8307,N_8314,N_8319,N_8320,N_8321,N_8322,N_8323,N_8328,N_8330,N_8333,N_8335,N_8338,N_8340,N_8342,N_8343,N_8344,N_8346,N_8347,N_8349,N_8351,N_8352,N_8353,N_8354,N_8356,N_8357,N_8358,N_8361,N_8363,N_8366,N_8367,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8376,N_8377,N_8378,N_8379,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8393,N_8394,N_8395,N_8397,N_8404,N_8405,N_8406,N_8415,N_8418,N_8421,N_8423,N_8424,N_8425,N_8426,N_8427,N_8430,N_8432,N_8433,N_8435,N_8436,N_8438,N_8441,N_8442,N_8443,N_8444,N_8446,N_8447,N_8448,N_8450,N_8451,N_8455,N_8457,N_8458,N_8459,N_8462,N_8464,N_8465,N_8466,N_8470,N_8471,N_8472,N_8474,N_8476,N_8477,N_8480,N_8482,N_8485,N_8488,N_8489,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8499,N_8500,N_8501,N_8504,N_8505,N_8506,N_8507,N_8508,N_8511,N_8512,N_8513,N_8515,N_8518,N_8519,N_8522,N_8524,N_8525,N_8527,N_8529,N_8531,N_8532,N_8533,N_8534,N_8535,N_8537,N_8539,N_8540,N_8541,N_8544,N_8545,N_8546,N_8548,N_8549,N_8552,N_8553,N_8554,N_8556,N_8557,N_8558,N_8561,N_8562,N_8563,N_8565,N_8566,N_8568,N_8569,N_8570,N_8573,N_8575,N_8576,N_8578,N_8579,N_8580,N_8581,N_8584,N_8587,N_8588,N_8589,N_8590,N_8593,N_8594,N_8598,N_8600,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8609,N_8610,N_8611,N_8612,N_8614,N_8616,N_8618,N_8620,N_8621,N_8623,N_8626,N_8628,N_8633,N_8635,N_8636,N_8638,N_8639,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8652,N_8653,N_8656,N_8659,N_8661,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8671,N_8672,N_8673,N_8674,N_8675,N_8679,N_8680,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8693,N_8697,N_8699,N_8700,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8719,N_8720,N_8721,N_8722,N_8723,N_8725,N_8726,N_8728,N_8730,N_8731,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8741,N_8744,N_8745,N_8747,N_8748,N_8750,N_8752,N_8754,N_8755,N_8757,N_8758,N_8761,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8773,N_8774,N_8775,N_8779,N_8781,N_8782,N_8785,N_8786,N_8787,N_8788,N_8793,N_8795,N_8796,N_8798,N_8799,N_8800,N_8802,N_8804,N_8805,N_8806,N_8808,N_8809,N_8816,N_8817,N_8820,N_8821,N_8822,N_8824,N_8825,N_8826,N_8831,N_8832,N_8835,N_8836,N_8837,N_8840,N_8842,N_8843,N_8844,N_8846,N_8847,N_8849,N_8850,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8861,N_8862,N_8866,N_8868,N_8869,N_8870,N_8871,N_8874,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8883,N_8885,N_8887,N_8889,N_8890,N_8892,N_8893,N_8895,N_8896,N_8897,N_8901,N_8902,N_8903,N_8906,N_8907,N_8908,N_8909,N_8911,N_8913,N_8914,N_8915,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8933,N_8934,N_8935,N_8936,N_8939,N_8940,N_8942,N_8945,N_8946,N_8947,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8958,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8975,N_8976,N_8978,N_8979,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8988,N_8990,N_8991,N_8993,N_8995,N_8996,N_9002,N_9004,N_9005,N_9006,N_9007,N_9012,N_9013,N_9014,N_9015,N_9017,N_9019,N_9022,N_9024,N_9025,N_9026,N_9030,N_9031,N_9035,N_9036,N_9039,N_9040,N_9041,N_9042,N_9043,N_9045,N_9047,N_9048,N_9050,N_9051,N_9053,N_9055,N_9056,N_9059,N_9060,N_9061,N_9065,N_9066,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9075,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9087,N_9088,N_9089,N_9090,N_9092,N_9093,N_9094,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9105,N_9108,N_9110,N_9113,N_9114,N_9116,N_9118,N_9123,N_9124,N_9125,N_9126,N_9128,N_9131,N_9133,N_9134,N_9137,N_9138,N_9139,N_9142,N_9146,N_9147,N_9151,N_9153,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9167,N_9168,N_9170,N_9172,N_9176,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9189,N_9191,N_9192,N_9195,N_9196,N_9197,N_9198,N_9200,N_9201,N_9203,N_9204,N_9205,N_9207,N_9209,N_9210,N_9214,N_9216,N_9217,N_9218,N_9220,N_9221,N_9223,N_9225,N_9226,N_9229,N_9230,N_9232,N_9233,N_9236,N_9240,N_9241,N_9242,N_9243,N_9245,N_9247,N_9250,N_9251,N_9252,N_9254,N_9255,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9269,N_9271,N_9272,N_9274,N_9276,N_9278,N_9280,N_9283,N_9284,N_9287,N_9288,N_9289,N_9290,N_9292,N_9293,N_9294,N_9295,N_9298,N_9301,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9313,N_9314,N_9319,N_9320,N_9323,N_9324,N_9325,N_9327,N_9329,N_9330,N_9333,N_9335,N_9336,N_9337,N_9339,N_9341,N_9342,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9360,N_9362,N_9363,N_9365,N_9368,N_9369,N_9370,N_9373,N_9374,N_9375,N_9376,N_9380,N_9383,N_9385,N_9386,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9398,N_9399,N_9400,N_9402,N_9405,N_9406,N_9407,N_9409,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9420,N_9421,N_9422,N_9424,N_9425,N_9427,N_9429,N_9430,N_9431,N_9432,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9443,N_9446,N_9447,N_9448,N_9450,N_9451,N_9453,N_9454,N_9456,N_9458,N_9459,N_9460,N_9461,N_9463,N_9467,N_9468,N_9472,N_9473,N_9474,N_9476,N_9477,N_9478,N_9479,N_9481,N_9482,N_9483,N_9484,N_9487,N_9489,N_9490,N_9491,N_9493,N_9494,N_9495,N_9496,N_9498,N_9499,N_9500,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9510,N_9511,N_9512,N_9514,N_9515,N_9516,N_9518,N_9519,N_9521,N_9522,N_9523,N_9524,N_9529,N_9530,N_9532,N_9533,N_9534,N_9536,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9557,N_9558,N_9560,N_9564,N_9566,N_9567,N_9568,N_9569,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9579,N_9582,N_9585,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9601,N_9602,N_9603,N_9605,N_9606,N_9607,N_9610,N_9611,N_9612,N_9614,N_9615,N_9617,N_9618,N_9619,N_9620,N_9623,N_9624,N_9626,N_9627,N_9629,N_9631,N_9633,N_9634,N_9635,N_9636,N_9639,N_9640,N_9642,N_9643,N_9646,N_9647,N_9649,N_9650,N_9651,N_9653,N_9655,N_9659,N_9662,N_9663,N_9664,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9674,N_9676,N_9677,N_9680,N_9682,N_9684,N_9685,N_9686,N_9687,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9699,N_9702,N_9705,N_9706,N_9707,N_9708,N_9709,N_9711,N_9713,N_9715,N_9716,N_9717,N_9718,N_9719,N_9721,N_9722,N_9725,N_9731,N_9732,N_9733,N_9734,N_9735,N_9738,N_9739,N_9740,N_9743,N_9745,N_9747,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9758,N_9759,N_9760,N_9762,N_9764,N_9765,N_9767,N_9769,N_9772,N_9778,N_9779,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9788,N_9790,N_9791,N_9793,N_9795,N_9800,N_9803,N_9805,N_9810,N_9813,N_9814,N_9816,N_9817,N_9819,N_9820,N_9821,N_9822,N_9824,N_9826,N_9829,N_9831,N_9835,N_9836,N_9838,N_9839,N_9840,N_9841,N_9843,N_9844,N_9845,N_9846,N_9848,N_9849,N_9851,N_9852,N_9853,N_9855,N_9856,N_9857,N_9858,N_9860,N_9862,N_9864,N_9867,N_9868,N_9869,N_9870,N_9871,N_9873,N_9874,N_9876,N_9878,N_9879,N_9882,N_9883,N_9884,N_9885,N_9886,N_9888,N_9889,N_9891,N_9894,N_9895,N_9896,N_9897,N_9898,N_9902,N_9903,N_9905,N_9906,N_9907,N_9908,N_9910,N_9911,N_9912,N_9913,N_9914,N_9917,N_9919,N_9921,N_9923,N_9925,N_9927,N_9928,N_9929,N_9930,N_9932,N_9933,N_9934,N_9935,N_9936,N_9939,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9984,N_9986,N_9989,N_9990,N_9991,N_9992,N_9993,N_9995,N_9996,N_9997,N_9999;
nor U0 (N_0,In_311,In_964);
nor U1 (N_1,In_116,In_809);
nor U2 (N_2,In_463,In_806);
nand U3 (N_3,In_803,In_589);
nand U4 (N_4,In_847,In_628);
nand U5 (N_5,In_716,In_15);
and U6 (N_6,In_679,In_118);
nor U7 (N_7,In_71,In_101);
nand U8 (N_8,In_310,In_102);
and U9 (N_9,In_551,In_884);
or U10 (N_10,In_352,In_117);
or U11 (N_11,In_170,In_487);
nor U12 (N_12,In_692,In_504);
and U13 (N_13,In_201,In_432);
or U14 (N_14,In_251,In_660);
or U15 (N_15,In_133,In_1);
or U16 (N_16,In_388,In_888);
nor U17 (N_17,In_217,In_435);
and U18 (N_18,In_603,In_528);
nor U19 (N_19,In_357,In_287);
and U20 (N_20,In_488,In_649);
or U21 (N_21,In_824,In_778);
nand U22 (N_22,In_976,In_663);
or U23 (N_23,In_265,In_212);
nand U24 (N_24,In_637,In_10);
nor U25 (N_25,In_210,In_490);
and U26 (N_26,In_986,In_796);
nor U27 (N_27,In_507,In_676);
nand U28 (N_28,In_655,In_50);
nand U29 (N_29,In_685,In_455);
or U30 (N_30,In_6,In_171);
and U31 (N_31,In_99,In_256);
and U32 (N_32,In_963,In_861);
nor U33 (N_33,In_169,In_669);
nor U34 (N_34,In_387,In_804);
and U35 (N_35,In_48,In_233);
nand U36 (N_36,In_565,In_893);
nor U37 (N_37,In_393,In_390);
or U38 (N_38,In_899,In_264);
nor U39 (N_39,In_304,In_181);
and U40 (N_40,In_200,In_776);
or U41 (N_41,In_404,In_242);
and U42 (N_42,In_829,In_911);
and U43 (N_43,In_25,In_120);
nand U44 (N_44,In_254,In_224);
nand U45 (N_45,In_524,In_834);
or U46 (N_46,In_672,In_623);
nand U47 (N_47,In_330,In_398);
nor U48 (N_48,In_46,In_703);
and U49 (N_49,In_510,In_682);
or U50 (N_50,In_0,In_444);
or U51 (N_51,In_837,In_990);
nor U52 (N_52,In_947,In_536);
and U53 (N_53,In_844,In_100);
or U54 (N_54,In_593,In_842);
and U55 (N_55,In_44,In_850);
or U56 (N_56,In_278,In_7);
or U57 (N_57,In_907,In_949);
or U58 (N_58,In_706,In_502);
and U59 (N_59,In_106,In_903);
xor U60 (N_60,In_744,In_552);
nor U61 (N_61,In_789,In_857);
nand U62 (N_62,In_443,In_710);
nand U63 (N_63,In_600,In_817);
and U64 (N_64,In_599,In_209);
and U65 (N_65,In_695,In_422);
nor U66 (N_66,In_496,In_508);
or U67 (N_67,In_895,In_621);
nor U68 (N_68,In_318,In_225);
nand U69 (N_69,In_157,In_972);
and U70 (N_70,In_82,In_61);
nor U71 (N_71,In_428,In_67);
or U72 (N_72,In_403,In_790);
and U73 (N_73,In_51,In_702);
nand U74 (N_74,In_522,In_671);
and U75 (N_75,In_968,In_701);
xnor U76 (N_76,In_627,In_841);
nand U77 (N_77,In_944,In_440);
or U78 (N_78,In_412,In_883);
and U79 (N_79,In_196,In_529);
nor U80 (N_80,In_312,In_831);
nor U81 (N_81,In_743,In_696);
nand U82 (N_82,In_275,In_182);
or U83 (N_83,In_250,In_408);
and U84 (N_84,In_900,In_202);
or U85 (N_85,In_854,In_784);
xor U86 (N_86,In_997,In_184);
or U87 (N_87,In_625,In_800);
nand U88 (N_88,In_786,In_173);
nand U89 (N_89,In_152,In_684);
or U90 (N_90,In_610,In_650);
nand U91 (N_91,In_713,In_582);
or U92 (N_92,In_535,In_550);
nand U93 (N_93,In_283,In_125);
nor U94 (N_94,In_140,In_475);
nor U95 (N_95,In_467,In_991);
or U96 (N_96,In_41,In_172);
and U97 (N_97,In_165,In_104);
nand U98 (N_98,In_189,In_291);
and U99 (N_99,In_161,In_820);
nand U100 (N_100,In_369,In_73);
nor U101 (N_101,In_305,In_92);
nor U102 (N_102,In_747,In_816);
or U103 (N_103,In_849,In_481);
and U104 (N_104,In_979,In_728);
nand U105 (N_105,In_114,In_176);
or U106 (N_106,In_795,In_731);
or U107 (N_107,In_186,In_109);
nand U108 (N_108,In_592,In_881);
nor U109 (N_109,In_436,In_754);
and U110 (N_110,In_29,In_775);
or U111 (N_111,In_699,In_909);
nor U112 (N_112,In_215,In_810);
and U113 (N_113,In_822,In_213);
nand U114 (N_114,In_420,In_447);
and U115 (N_115,In_503,In_424);
nor U116 (N_116,In_833,In_853);
nand U117 (N_117,In_675,In_768);
nor U118 (N_118,In_76,In_517);
nor U119 (N_119,In_765,In_647);
nor U120 (N_120,In_917,In_783);
nand U121 (N_121,In_838,In_864);
and U122 (N_122,In_68,In_164);
or U123 (N_123,In_557,In_180);
nand U124 (N_124,In_150,In_587);
or U125 (N_125,In_244,In_630);
nand U126 (N_126,In_260,In_129);
or U127 (N_127,In_954,In_58);
nor U128 (N_128,In_658,In_666);
nand U129 (N_129,In_770,In_323);
nand U130 (N_130,In_662,In_985);
nor U131 (N_131,In_43,In_574);
nor U132 (N_132,In_236,In_411);
or U133 (N_133,In_322,In_926);
and U134 (N_134,In_220,In_95);
and U135 (N_135,In_762,In_158);
or U136 (N_136,In_818,In_400);
xor U137 (N_137,In_920,In_518);
and U138 (N_138,In_472,In_544);
and U139 (N_139,In_945,In_742);
and U140 (N_140,In_492,In_232);
nand U141 (N_141,In_825,In_644);
xor U142 (N_142,In_119,In_23);
nand U143 (N_143,In_590,In_280);
or U144 (N_144,In_908,In_808);
nand U145 (N_145,In_286,In_755);
and U146 (N_146,In_384,In_103);
nand U147 (N_147,In_539,In_429);
nand U148 (N_148,In_878,In_77);
nand U149 (N_149,In_867,In_335);
nor U150 (N_150,In_559,In_933);
nand U151 (N_151,In_690,In_668);
or U152 (N_152,In_758,In_197);
nor U153 (N_153,In_358,In_511);
nor U154 (N_154,In_446,In_640);
nand U155 (N_155,In_179,In_154);
and U156 (N_156,In_49,In_868);
nand U157 (N_157,In_537,In_266);
and U158 (N_158,In_607,In_717);
and U159 (N_159,In_601,In_329);
xnor U160 (N_160,In_477,In_484);
nor U161 (N_161,In_892,In_268);
nor U162 (N_162,In_930,In_950);
nand U163 (N_163,In_230,In_723);
and U164 (N_164,In_110,In_22);
nor U165 (N_165,In_585,In_284);
nor U166 (N_166,In_313,In_781);
and U167 (N_167,In_724,In_319);
or U168 (N_168,In_395,In_708);
nand U169 (N_169,In_247,In_417);
and U170 (N_170,In_819,In_320);
and U171 (N_171,In_63,In_356);
nand U172 (N_172,In_427,In_901);
or U173 (N_173,In_894,In_188);
or U174 (N_174,In_545,In_392);
and U175 (N_175,In_707,In_293);
nand U176 (N_176,In_64,In_890);
or U177 (N_177,In_111,In_577);
and U178 (N_178,In_923,In_555);
and U179 (N_179,In_714,In_343);
or U180 (N_180,In_315,In_897);
nor U181 (N_181,In_56,In_681);
and U182 (N_182,In_938,In_228);
or U183 (N_183,In_107,In_361);
or U184 (N_184,In_556,In_693);
nor U185 (N_185,In_190,In_813);
and U186 (N_186,In_826,In_580);
nor U187 (N_187,In_85,In_961);
nand U188 (N_188,In_345,In_664);
xor U189 (N_189,In_360,In_97);
nand U190 (N_190,In_126,In_66);
and U191 (N_191,In_397,In_141);
nand U192 (N_192,In_843,In_439);
and U193 (N_193,In_880,In_547);
nor U194 (N_194,In_996,In_289);
nor U195 (N_195,In_90,In_223);
and U196 (N_196,In_20,In_147);
or U197 (N_197,In_136,In_348);
nand U198 (N_198,In_636,In_277);
nor U199 (N_199,In_174,In_252);
and U200 (N_200,In_870,In_983);
nor U201 (N_201,In_840,In_78);
xor U202 (N_202,In_460,In_626);
and U203 (N_203,In_777,In_469);
nand U204 (N_204,In_764,In_137);
and U205 (N_205,In_981,In_887);
xor U206 (N_206,In_47,In_350);
nand U207 (N_207,In_498,In_711);
nor U208 (N_208,In_726,In_325);
and U209 (N_209,In_643,In_321);
and U210 (N_210,In_269,In_60);
and U211 (N_211,In_121,In_858);
nand U212 (N_212,In_471,In_652);
nand U213 (N_213,In_379,In_752);
and U214 (N_214,In_36,In_769);
or U215 (N_215,In_175,In_937);
and U216 (N_216,In_382,In_211);
and U217 (N_217,In_377,In_386);
and U218 (N_218,In_814,In_124);
and U219 (N_219,In_499,In_418);
or U220 (N_220,In_573,In_543);
xnor U221 (N_221,In_656,In_457);
nand U222 (N_222,In_454,In_263);
or U223 (N_223,In_866,In_191);
nand U224 (N_224,In_569,In_328);
nor U225 (N_225,In_326,In_549);
nand U226 (N_226,In_351,In_598);
or U227 (N_227,In_402,In_689);
nand U228 (N_228,In_309,In_4);
and U229 (N_229,In_115,In_376);
xor U230 (N_230,In_494,In_2);
nor U231 (N_231,In_952,In_13);
nor U232 (N_232,In_542,In_339);
nand U233 (N_233,In_654,In_505);
or U234 (N_234,In_365,In_279);
or U235 (N_235,In_218,In_801);
and U236 (N_236,In_468,In_595);
nor U237 (N_237,In_146,In_896);
nor U238 (N_238,In_729,In_530);
or U239 (N_239,In_192,In_482);
or U240 (N_240,In_929,In_296);
nor U241 (N_241,In_648,In_787);
nand U242 (N_242,In_738,In_88);
and U243 (N_243,In_55,In_597);
nor U244 (N_244,In_353,In_239);
or U245 (N_245,In_670,In_94);
nor U246 (N_246,In_462,In_53);
nand U247 (N_247,In_486,In_958);
and U248 (N_248,In_812,In_383);
nand U249 (N_249,In_26,In_782);
or U250 (N_250,In_767,In_302);
and U251 (N_251,In_969,In_401);
nand U252 (N_252,In_521,In_928);
nor U253 (N_253,In_295,In_34);
nand U254 (N_254,In_229,In_359);
or U255 (N_255,In_259,In_619);
and U256 (N_256,In_425,In_875);
and U257 (N_257,In_583,In_736);
nand U258 (N_258,In_389,In_588);
nor U259 (N_259,In_285,In_281);
nand U260 (N_260,In_300,In_37);
nor U261 (N_261,In_445,In_288);
nand U262 (N_262,In_45,In_772);
nand U263 (N_263,In_862,In_354);
or U264 (N_264,In_303,In_391);
nor U265 (N_265,In_112,In_364);
nand U266 (N_266,In_779,In_130);
nand U267 (N_267,In_891,In_21);
nor U268 (N_268,In_591,In_608);
nor U269 (N_269,In_617,In_380);
and U270 (N_270,In_271,In_546);
nor U271 (N_271,In_344,In_378);
or U272 (N_272,In_461,In_28);
or U273 (N_273,In_629,In_553);
nor U274 (N_274,In_307,In_959);
nand U275 (N_275,In_931,In_519);
and U276 (N_276,In_665,In_915);
or U277 (N_277,In_451,In_459);
nand U278 (N_278,In_142,In_327);
or U279 (N_279,In_815,In_602);
nor U280 (N_280,In_774,In_240);
and U281 (N_281,In_415,In_992);
xor U282 (N_282,In_520,In_962);
or U283 (N_283,In_571,In_988);
or U284 (N_284,In_995,In_199);
and U285 (N_285,In_533,In_674);
nand U286 (N_286,In_128,In_661);
nand U287 (N_287,In_54,In_678);
nor U288 (N_288,In_127,In_677);
or U289 (N_289,In_32,In_38);
or U290 (N_290,In_253,In_470);
nand U291 (N_291,In_659,In_579);
and U292 (N_292,In_434,In_456);
nor U293 (N_293,In_299,In_410);
or U294 (N_294,In_187,In_262);
xor U295 (N_295,In_978,In_913);
or U296 (N_296,In_148,In_105);
and U297 (N_297,In_297,In_156);
and U298 (N_298,In_879,In_877);
nand U299 (N_299,In_832,In_616);
nor U300 (N_300,In_59,In_168);
nor U301 (N_301,In_749,In_122);
or U302 (N_302,In_821,In_430);
and U303 (N_303,In_618,In_414);
or U304 (N_304,In_596,In_480);
or U305 (N_305,In_856,In_802);
or U306 (N_306,In_791,In_999);
or U307 (N_307,In_513,In_491);
nor U308 (N_308,In_453,In_975);
or U309 (N_309,In_205,In_135);
nand U310 (N_310,In_123,In_509);
or U311 (N_311,In_340,In_394);
nand U312 (N_312,In_955,In_835);
or U313 (N_313,In_347,In_646);
and U314 (N_314,In_761,In_960);
nor U315 (N_315,In_575,In_438);
nand U316 (N_316,In_166,In_860);
and U317 (N_317,In_349,In_586);
nor U318 (N_318,In_612,In_741);
nor U319 (N_319,In_74,In_301);
nand U320 (N_320,In_567,In_902);
and U321 (N_321,In_96,In_686);
nor U322 (N_322,In_921,In_653);
or U323 (N_323,In_241,In_698);
and U324 (N_324,In_722,In_614);
nand U325 (N_325,In_993,In_14);
nand U326 (N_326,In_984,In_914);
nor U327 (N_327,In_423,In_785);
nor U328 (N_328,In_620,In_576);
and U329 (N_329,In_760,In_407);
or U330 (N_330,In_151,In_735);
and U331 (N_331,In_362,In_160);
nand U332 (N_332,In_381,In_194);
and U333 (N_333,In_771,In_516);
and U334 (N_334,In_317,In_437);
and U335 (N_335,In_756,In_906);
or U336 (N_336,In_87,In_965);
nand U337 (N_337,In_971,In_939);
or U338 (N_338,In_584,In_273);
and U339 (N_339,In_967,In_581);
nand U340 (N_340,In_966,In_144);
nand U341 (N_341,In_916,In_474);
nor U342 (N_342,In_534,In_846);
nor U343 (N_343,In_632,In_27);
or U344 (N_344,In_163,In_11);
and U345 (N_345,In_178,In_594);
or U346 (N_346,In_70,In_235);
nand U347 (N_347,In_237,In_807);
and U348 (N_348,In_561,In_84);
or U349 (N_349,In_385,In_442);
nand U350 (N_350,In_927,In_609);
nand U351 (N_351,In_905,In_255);
or U352 (N_352,In_977,In_341);
nor U353 (N_353,In_139,In_89);
nor U354 (N_354,In_998,In_57);
and U355 (N_355,In_538,In_645);
and U356 (N_356,In_162,In_290);
nor U357 (N_357,In_953,In_206);
or U358 (N_358,In_221,In_869);
nand U359 (N_359,In_207,In_697);
or U360 (N_360,In_872,In_134);
and U361 (N_361,In_132,In_375);
and U362 (N_362,In_919,In_336);
or U363 (N_363,In_874,In_40);
nor U364 (N_364,In_370,In_578);
nand U365 (N_365,In_799,In_149);
nand U366 (N_366,In_638,In_563);
nand U367 (N_367,In_924,In_372);
or U368 (N_368,In_257,In_396);
or U369 (N_369,In_982,In_267);
nand U370 (N_370,In_243,In_560);
nor U371 (N_371,In_974,In_548);
nand U372 (N_372,In_709,In_635);
nand U373 (N_373,In_848,In_721);
xor U374 (N_374,In_80,In_143);
or U375 (N_375,In_419,In_727);
and U376 (N_376,In_501,In_641);
nor U377 (N_377,In_33,In_934);
and U378 (N_378,In_355,In_421);
or U379 (N_379,In_332,In_465);
nor U380 (N_380,In_495,In_195);
and U381 (N_381,In_406,In_93);
nand U382 (N_382,In_483,In_409);
nor U383 (N_383,In_604,In_828);
nor U384 (N_384,In_918,In_153);
or U385 (N_385,In_852,In_86);
nor U386 (N_386,In_987,In_9);
or U387 (N_387,In_346,In_248);
or U388 (N_388,In_527,In_448);
or U389 (N_389,In_624,In_940);
nand U390 (N_390,In_298,In_970);
nor U391 (N_391,In_12,In_793);
and U392 (N_392,In_936,In_514);
nor U393 (N_393,In_338,In_306);
nand U394 (N_394,In_433,In_431);
nand U395 (N_395,In_942,In_526);
nor U396 (N_396,In_753,In_737);
or U397 (N_397,In_145,In_568);
nand U398 (N_398,In_532,In_798);
and U399 (N_399,In_688,In_91);
nor U400 (N_400,In_606,In_367);
nor U401 (N_401,In_131,In_155);
nor U402 (N_402,In_757,In_751);
nand U403 (N_403,In_35,In_30);
nand U404 (N_404,In_167,In_712);
or U405 (N_405,In_270,In_631);
and U406 (N_406,In_214,In_234);
and U407 (N_407,In_912,In_932);
and U408 (N_408,In_65,In_941);
nand U409 (N_409,In_566,In_374);
and U410 (N_410,In_855,In_994);
and U411 (N_411,In_622,In_845);
nand U412 (N_412,In_72,In_108);
nand U413 (N_413,In_525,In_540);
or U414 (N_414,In_863,In_732);
nand U415 (N_415,In_691,In_177);
and U416 (N_416,In_763,In_198);
and U417 (N_417,In_836,In_839);
and U418 (N_418,In_24,In_558);
nor U419 (N_419,In_75,In_368);
nand U420 (N_420,In_562,In_238);
nand U421 (N_421,In_450,In_740);
and U422 (N_422,In_426,In_113);
or U423 (N_423,In_337,In_464);
or U424 (N_424,In_792,In_773);
nand U425 (N_425,In_333,In_700);
and U426 (N_426,In_42,In_642);
nor U427 (N_427,In_687,In_739);
nand U428 (N_428,In_18,In_633);
or U429 (N_429,In_31,In_613);
nor U430 (N_430,In_851,In_203);
and U431 (N_431,In_657,In_683);
and U432 (N_432,In_16,In_925);
or U433 (N_433,In_493,In_980);
or U434 (N_434,In_943,In_231);
or U435 (N_435,In_957,In_720);
and U436 (N_436,In_441,In_497);
nor U437 (N_437,In_208,In_541);
and U438 (N_438,In_572,In_605);
or U439 (N_439,In_366,In_39);
nand U440 (N_440,In_951,In_485);
nor U441 (N_441,In_3,In_219);
nand U442 (N_442,In_730,In_399);
and U443 (N_443,In_805,In_859);
nand U444 (N_444,In_185,In_882);
or U445 (N_445,In_667,In_935);
or U446 (N_446,In_889,In_989);
or U447 (N_447,In_258,In_973);
nor U448 (N_448,In_363,In_811);
or U449 (N_449,In_748,In_371);
xor U450 (N_450,In_314,In_873);
or U451 (N_451,In_830,In_342);
nor U452 (N_452,In_797,In_458);
and U453 (N_453,In_17,In_245);
or U454 (N_454,In_704,In_413);
or U455 (N_455,In_138,In_885);
or U456 (N_456,In_733,In_261);
nand U457 (N_457,In_512,In_780);
xnor U458 (N_458,In_489,In_222);
or U459 (N_459,In_308,In_715);
or U460 (N_460,In_373,In_745);
nand U461 (N_461,In_705,In_718);
or U462 (N_462,In_272,In_292);
nor U463 (N_463,In_69,In_827);
nor U464 (N_464,In_956,In_865);
nor U465 (N_465,In_570,In_766);
nor U466 (N_466,In_193,In_216);
or U467 (N_467,In_81,In_794);
or U468 (N_468,In_500,In_746);
nor U469 (N_469,In_554,In_331);
or U470 (N_470,In_324,In_62);
or U471 (N_471,In_876,In_946);
nand U472 (N_472,In_904,In_466);
nor U473 (N_473,In_416,In_531);
or U474 (N_474,In_898,In_910);
nor U475 (N_475,In_5,In_871);
or U476 (N_476,In_476,In_226);
nor U477 (N_477,In_478,In_183);
nor U478 (N_478,In_276,In_734);
nand U479 (N_479,In_473,In_405);
and U480 (N_480,In_316,In_564);
nand U481 (N_481,In_79,In_719);
nor U482 (N_482,In_515,In_334);
and U483 (N_483,In_227,In_98);
and U484 (N_484,In_651,In_204);
xor U485 (N_485,In_823,In_922);
or U486 (N_486,In_19,In_479);
nor U487 (N_487,In_615,In_452);
nand U488 (N_488,In_282,In_680);
and U489 (N_489,In_694,In_886);
nor U490 (N_490,In_294,In_159);
or U491 (N_491,In_948,In_246);
or U492 (N_492,In_274,In_506);
or U493 (N_493,In_639,In_8);
or U494 (N_494,In_673,In_725);
and U495 (N_495,In_83,In_634);
or U496 (N_496,In_759,In_249);
and U497 (N_497,In_52,In_449);
or U498 (N_498,In_788,In_523);
nor U499 (N_499,In_750,In_611);
nor U500 (N_500,In_702,In_332);
or U501 (N_501,In_940,In_590);
or U502 (N_502,In_454,In_771);
nand U503 (N_503,In_77,In_688);
nand U504 (N_504,In_368,In_447);
nand U505 (N_505,In_75,In_386);
nand U506 (N_506,In_454,In_929);
or U507 (N_507,In_683,In_201);
and U508 (N_508,In_224,In_545);
and U509 (N_509,In_27,In_163);
or U510 (N_510,In_325,In_191);
nor U511 (N_511,In_242,In_158);
and U512 (N_512,In_456,In_571);
nand U513 (N_513,In_100,In_380);
nand U514 (N_514,In_625,In_521);
nand U515 (N_515,In_280,In_197);
or U516 (N_516,In_390,In_384);
nor U517 (N_517,In_504,In_307);
or U518 (N_518,In_918,In_258);
or U519 (N_519,In_40,In_372);
and U520 (N_520,In_788,In_108);
nand U521 (N_521,In_914,In_648);
nand U522 (N_522,In_197,In_727);
and U523 (N_523,In_44,In_763);
nand U524 (N_524,In_59,In_794);
nor U525 (N_525,In_582,In_282);
and U526 (N_526,In_851,In_603);
and U527 (N_527,In_443,In_242);
or U528 (N_528,In_851,In_478);
and U529 (N_529,In_211,In_142);
nand U530 (N_530,In_468,In_228);
nor U531 (N_531,In_387,In_611);
nand U532 (N_532,In_138,In_608);
and U533 (N_533,In_745,In_983);
and U534 (N_534,In_818,In_412);
or U535 (N_535,In_137,In_407);
and U536 (N_536,In_156,In_870);
nor U537 (N_537,In_545,In_821);
nand U538 (N_538,In_99,In_593);
nand U539 (N_539,In_589,In_738);
nand U540 (N_540,In_935,In_988);
or U541 (N_541,In_352,In_187);
or U542 (N_542,In_813,In_375);
nor U543 (N_543,In_85,In_123);
or U544 (N_544,In_97,In_861);
and U545 (N_545,In_209,In_844);
and U546 (N_546,In_859,In_928);
or U547 (N_547,In_756,In_703);
nor U548 (N_548,In_691,In_391);
nand U549 (N_549,In_601,In_731);
or U550 (N_550,In_884,In_270);
and U551 (N_551,In_275,In_23);
or U552 (N_552,In_362,In_472);
nor U553 (N_553,In_848,In_945);
nor U554 (N_554,In_71,In_991);
and U555 (N_555,In_480,In_60);
nor U556 (N_556,In_267,In_433);
nand U557 (N_557,In_281,In_216);
and U558 (N_558,In_689,In_858);
and U559 (N_559,In_348,In_267);
nor U560 (N_560,In_671,In_375);
or U561 (N_561,In_332,In_8);
and U562 (N_562,In_489,In_358);
or U563 (N_563,In_513,In_790);
or U564 (N_564,In_918,In_243);
and U565 (N_565,In_150,In_82);
or U566 (N_566,In_463,In_219);
or U567 (N_567,In_979,In_11);
and U568 (N_568,In_679,In_82);
and U569 (N_569,In_960,In_621);
or U570 (N_570,In_910,In_31);
nand U571 (N_571,In_53,In_172);
and U572 (N_572,In_543,In_732);
nand U573 (N_573,In_697,In_529);
or U574 (N_574,In_270,In_637);
or U575 (N_575,In_309,In_506);
nand U576 (N_576,In_23,In_633);
and U577 (N_577,In_60,In_709);
or U578 (N_578,In_345,In_680);
or U579 (N_579,In_557,In_337);
and U580 (N_580,In_949,In_58);
and U581 (N_581,In_677,In_546);
nor U582 (N_582,In_833,In_376);
nor U583 (N_583,In_577,In_759);
nand U584 (N_584,In_784,In_489);
nor U585 (N_585,In_391,In_769);
nand U586 (N_586,In_672,In_283);
or U587 (N_587,In_441,In_953);
or U588 (N_588,In_170,In_490);
nor U589 (N_589,In_308,In_693);
or U590 (N_590,In_298,In_844);
and U591 (N_591,In_391,In_940);
or U592 (N_592,In_169,In_85);
xnor U593 (N_593,In_169,In_954);
and U594 (N_594,In_654,In_885);
nand U595 (N_595,In_730,In_134);
or U596 (N_596,In_311,In_710);
or U597 (N_597,In_797,In_916);
nor U598 (N_598,In_473,In_461);
nand U599 (N_599,In_775,In_139);
or U600 (N_600,In_760,In_859);
nand U601 (N_601,In_240,In_583);
nand U602 (N_602,In_780,In_770);
nand U603 (N_603,In_742,In_656);
and U604 (N_604,In_568,In_779);
nor U605 (N_605,In_668,In_181);
nor U606 (N_606,In_177,In_464);
or U607 (N_607,In_220,In_953);
xor U608 (N_608,In_278,In_251);
or U609 (N_609,In_846,In_670);
or U610 (N_610,In_754,In_946);
nand U611 (N_611,In_360,In_512);
nor U612 (N_612,In_380,In_400);
or U613 (N_613,In_193,In_252);
nor U614 (N_614,In_985,In_498);
nand U615 (N_615,In_666,In_115);
and U616 (N_616,In_210,In_962);
or U617 (N_617,In_0,In_342);
nor U618 (N_618,In_406,In_864);
or U619 (N_619,In_981,In_314);
nor U620 (N_620,In_31,In_45);
nand U621 (N_621,In_750,In_39);
nor U622 (N_622,In_759,In_909);
or U623 (N_623,In_53,In_883);
and U624 (N_624,In_63,In_607);
nand U625 (N_625,In_619,In_879);
nand U626 (N_626,In_8,In_235);
nand U627 (N_627,In_309,In_41);
and U628 (N_628,In_644,In_223);
and U629 (N_629,In_31,In_460);
or U630 (N_630,In_892,In_621);
nand U631 (N_631,In_998,In_357);
or U632 (N_632,In_562,In_479);
or U633 (N_633,In_634,In_483);
nand U634 (N_634,In_217,In_813);
nand U635 (N_635,In_913,In_378);
nor U636 (N_636,In_927,In_475);
nor U637 (N_637,In_701,In_987);
or U638 (N_638,In_162,In_464);
or U639 (N_639,In_874,In_917);
and U640 (N_640,In_976,In_944);
or U641 (N_641,In_69,In_846);
and U642 (N_642,In_11,In_338);
nor U643 (N_643,In_591,In_271);
nand U644 (N_644,In_121,In_639);
or U645 (N_645,In_201,In_141);
nand U646 (N_646,In_446,In_375);
nor U647 (N_647,In_200,In_831);
nor U648 (N_648,In_690,In_209);
and U649 (N_649,In_845,In_612);
or U650 (N_650,In_754,In_494);
and U651 (N_651,In_781,In_334);
nor U652 (N_652,In_158,In_440);
and U653 (N_653,In_126,In_177);
or U654 (N_654,In_821,In_198);
and U655 (N_655,In_403,In_923);
or U656 (N_656,In_823,In_670);
and U657 (N_657,In_534,In_337);
nand U658 (N_658,In_400,In_501);
or U659 (N_659,In_427,In_196);
nand U660 (N_660,In_245,In_914);
nand U661 (N_661,In_621,In_447);
xnor U662 (N_662,In_254,In_902);
or U663 (N_663,In_649,In_137);
and U664 (N_664,In_983,In_264);
nand U665 (N_665,In_687,In_768);
or U666 (N_666,In_630,In_627);
nand U667 (N_667,In_984,In_610);
and U668 (N_668,In_351,In_997);
nor U669 (N_669,In_144,In_373);
nand U670 (N_670,In_568,In_621);
nor U671 (N_671,In_235,In_617);
or U672 (N_672,In_59,In_188);
nand U673 (N_673,In_370,In_472);
or U674 (N_674,In_733,In_307);
and U675 (N_675,In_466,In_968);
nor U676 (N_676,In_654,In_453);
nand U677 (N_677,In_105,In_337);
nor U678 (N_678,In_755,In_628);
nor U679 (N_679,In_455,In_242);
xor U680 (N_680,In_924,In_890);
nand U681 (N_681,In_896,In_148);
nand U682 (N_682,In_801,In_877);
and U683 (N_683,In_733,In_582);
nand U684 (N_684,In_758,In_838);
nor U685 (N_685,In_120,In_241);
or U686 (N_686,In_827,In_299);
nor U687 (N_687,In_120,In_760);
and U688 (N_688,In_316,In_786);
and U689 (N_689,In_912,In_647);
and U690 (N_690,In_742,In_0);
and U691 (N_691,In_391,In_910);
nor U692 (N_692,In_377,In_188);
nand U693 (N_693,In_87,In_273);
nor U694 (N_694,In_547,In_396);
or U695 (N_695,In_482,In_772);
or U696 (N_696,In_463,In_527);
nand U697 (N_697,In_478,In_808);
nand U698 (N_698,In_289,In_267);
nor U699 (N_699,In_276,In_443);
xor U700 (N_700,In_156,In_460);
and U701 (N_701,In_781,In_133);
or U702 (N_702,In_694,In_217);
nand U703 (N_703,In_589,In_64);
nor U704 (N_704,In_955,In_163);
nor U705 (N_705,In_534,In_224);
and U706 (N_706,In_546,In_976);
and U707 (N_707,In_847,In_947);
nand U708 (N_708,In_365,In_747);
and U709 (N_709,In_318,In_307);
nor U710 (N_710,In_267,In_414);
and U711 (N_711,In_387,In_955);
nand U712 (N_712,In_407,In_583);
nor U713 (N_713,In_806,In_165);
nor U714 (N_714,In_290,In_95);
xor U715 (N_715,In_498,In_116);
and U716 (N_716,In_695,In_510);
nor U717 (N_717,In_597,In_603);
or U718 (N_718,In_788,In_340);
and U719 (N_719,In_371,In_470);
nand U720 (N_720,In_947,In_253);
or U721 (N_721,In_102,In_798);
nor U722 (N_722,In_377,In_704);
and U723 (N_723,In_75,In_494);
or U724 (N_724,In_498,In_234);
nor U725 (N_725,In_489,In_318);
nor U726 (N_726,In_623,In_374);
nand U727 (N_727,In_158,In_128);
or U728 (N_728,In_858,In_823);
and U729 (N_729,In_331,In_133);
nor U730 (N_730,In_5,In_533);
nand U731 (N_731,In_209,In_18);
nor U732 (N_732,In_91,In_504);
and U733 (N_733,In_397,In_798);
nand U734 (N_734,In_783,In_431);
and U735 (N_735,In_976,In_551);
and U736 (N_736,In_796,In_800);
xor U737 (N_737,In_136,In_262);
and U738 (N_738,In_863,In_771);
nor U739 (N_739,In_825,In_716);
or U740 (N_740,In_785,In_200);
or U741 (N_741,In_938,In_369);
or U742 (N_742,In_177,In_430);
and U743 (N_743,In_896,In_979);
and U744 (N_744,In_176,In_804);
nor U745 (N_745,In_629,In_849);
and U746 (N_746,In_957,In_190);
or U747 (N_747,In_180,In_630);
nor U748 (N_748,In_706,In_15);
nand U749 (N_749,In_571,In_185);
nor U750 (N_750,In_249,In_857);
or U751 (N_751,In_361,In_503);
nand U752 (N_752,In_621,In_869);
and U753 (N_753,In_82,In_253);
nand U754 (N_754,In_133,In_687);
and U755 (N_755,In_97,In_540);
and U756 (N_756,In_498,In_895);
nor U757 (N_757,In_595,In_966);
nor U758 (N_758,In_24,In_660);
nor U759 (N_759,In_11,In_968);
or U760 (N_760,In_171,In_376);
and U761 (N_761,In_794,In_993);
nor U762 (N_762,In_822,In_604);
nor U763 (N_763,In_154,In_277);
nand U764 (N_764,In_851,In_350);
and U765 (N_765,In_6,In_130);
and U766 (N_766,In_695,In_788);
or U767 (N_767,In_196,In_840);
nor U768 (N_768,In_100,In_43);
or U769 (N_769,In_967,In_355);
nor U770 (N_770,In_876,In_948);
nand U771 (N_771,In_872,In_587);
nand U772 (N_772,In_34,In_107);
and U773 (N_773,In_275,In_99);
nor U774 (N_774,In_676,In_150);
nand U775 (N_775,In_864,In_527);
nor U776 (N_776,In_220,In_908);
xor U777 (N_777,In_30,In_54);
and U778 (N_778,In_197,In_471);
and U779 (N_779,In_320,In_921);
nor U780 (N_780,In_108,In_588);
nor U781 (N_781,In_988,In_525);
or U782 (N_782,In_22,In_135);
nor U783 (N_783,In_986,In_49);
nor U784 (N_784,In_469,In_647);
and U785 (N_785,In_82,In_20);
and U786 (N_786,In_910,In_452);
nor U787 (N_787,In_578,In_179);
and U788 (N_788,In_508,In_871);
nor U789 (N_789,In_268,In_461);
nand U790 (N_790,In_632,In_870);
nor U791 (N_791,In_290,In_326);
nand U792 (N_792,In_711,In_869);
xnor U793 (N_793,In_549,In_601);
or U794 (N_794,In_271,In_324);
nor U795 (N_795,In_233,In_23);
nand U796 (N_796,In_628,In_306);
nor U797 (N_797,In_926,In_206);
nand U798 (N_798,In_91,In_781);
nor U799 (N_799,In_704,In_385);
or U800 (N_800,In_149,In_990);
or U801 (N_801,In_147,In_273);
nand U802 (N_802,In_861,In_447);
nand U803 (N_803,In_414,In_337);
and U804 (N_804,In_576,In_827);
nand U805 (N_805,In_761,In_590);
nand U806 (N_806,In_655,In_731);
nand U807 (N_807,In_217,In_803);
nor U808 (N_808,In_22,In_888);
xor U809 (N_809,In_894,In_701);
xor U810 (N_810,In_375,In_298);
nand U811 (N_811,In_319,In_704);
or U812 (N_812,In_162,In_715);
and U813 (N_813,In_713,In_696);
and U814 (N_814,In_113,In_447);
nor U815 (N_815,In_998,In_352);
or U816 (N_816,In_723,In_169);
or U817 (N_817,In_278,In_821);
and U818 (N_818,In_424,In_823);
nor U819 (N_819,In_921,In_472);
and U820 (N_820,In_643,In_12);
or U821 (N_821,In_230,In_373);
and U822 (N_822,In_432,In_549);
and U823 (N_823,In_398,In_110);
nand U824 (N_824,In_337,In_270);
nor U825 (N_825,In_187,In_770);
and U826 (N_826,In_730,In_99);
nor U827 (N_827,In_185,In_319);
nor U828 (N_828,In_464,In_600);
nand U829 (N_829,In_864,In_953);
and U830 (N_830,In_564,In_944);
or U831 (N_831,In_992,In_206);
or U832 (N_832,In_293,In_667);
or U833 (N_833,In_626,In_440);
or U834 (N_834,In_430,In_998);
and U835 (N_835,In_12,In_301);
and U836 (N_836,In_520,In_214);
nor U837 (N_837,In_377,In_383);
and U838 (N_838,In_614,In_180);
nand U839 (N_839,In_206,In_962);
nor U840 (N_840,In_134,In_313);
nand U841 (N_841,In_923,In_874);
nor U842 (N_842,In_274,In_367);
xor U843 (N_843,In_302,In_749);
nor U844 (N_844,In_502,In_283);
and U845 (N_845,In_491,In_345);
or U846 (N_846,In_171,In_648);
nand U847 (N_847,In_835,In_689);
nand U848 (N_848,In_783,In_7);
nand U849 (N_849,In_927,In_579);
or U850 (N_850,In_786,In_305);
or U851 (N_851,In_425,In_697);
nor U852 (N_852,In_37,In_265);
or U853 (N_853,In_828,In_679);
xor U854 (N_854,In_419,In_615);
and U855 (N_855,In_832,In_500);
and U856 (N_856,In_8,In_497);
and U857 (N_857,In_620,In_357);
xnor U858 (N_858,In_220,In_82);
and U859 (N_859,In_596,In_641);
or U860 (N_860,In_773,In_329);
and U861 (N_861,In_931,In_721);
or U862 (N_862,In_954,In_60);
nor U863 (N_863,In_291,In_391);
nand U864 (N_864,In_788,In_659);
and U865 (N_865,In_78,In_655);
and U866 (N_866,In_229,In_360);
and U867 (N_867,In_599,In_620);
or U868 (N_868,In_806,In_232);
or U869 (N_869,In_106,In_391);
xnor U870 (N_870,In_430,In_775);
xnor U871 (N_871,In_496,In_516);
nor U872 (N_872,In_722,In_156);
nand U873 (N_873,In_49,In_524);
or U874 (N_874,In_301,In_550);
and U875 (N_875,In_983,In_902);
nor U876 (N_876,In_281,In_481);
nand U877 (N_877,In_321,In_362);
nor U878 (N_878,In_333,In_552);
nor U879 (N_879,In_318,In_787);
nor U880 (N_880,In_966,In_505);
or U881 (N_881,In_384,In_598);
nor U882 (N_882,In_198,In_228);
or U883 (N_883,In_839,In_455);
nor U884 (N_884,In_416,In_86);
xor U885 (N_885,In_171,In_44);
nand U886 (N_886,In_294,In_291);
and U887 (N_887,In_519,In_150);
nand U888 (N_888,In_581,In_157);
nor U889 (N_889,In_571,In_353);
nand U890 (N_890,In_675,In_606);
or U891 (N_891,In_50,In_186);
and U892 (N_892,In_423,In_160);
nand U893 (N_893,In_39,In_791);
xor U894 (N_894,In_130,In_587);
or U895 (N_895,In_270,In_706);
or U896 (N_896,In_49,In_444);
nand U897 (N_897,In_29,In_22);
or U898 (N_898,In_696,In_771);
nand U899 (N_899,In_952,In_239);
nand U900 (N_900,In_438,In_296);
or U901 (N_901,In_374,In_106);
or U902 (N_902,In_300,In_453);
and U903 (N_903,In_196,In_566);
or U904 (N_904,In_161,In_677);
or U905 (N_905,In_260,In_496);
or U906 (N_906,In_579,In_901);
and U907 (N_907,In_994,In_379);
nor U908 (N_908,In_650,In_549);
or U909 (N_909,In_808,In_627);
nor U910 (N_910,In_557,In_421);
nand U911 (N_911,In_425,In_715);
or U912 (N_912,In_243,In_386);
nand U913 (N_913,In_610,In_550);
and U914 (N_914,In_869,In_257);
or U915 (N_915,In_278,In_14);
nand U916 (N_916,In_451,In_864);
nor U917 (N_917,In_695,In_406);
nand U918 (N_918,In_745,In_404);
nand U919 (N_919,In_181,In_104);
and U920 (N_920,In_377,In_567);
or U921 (N_921,In_3,In_393);
nor U922 (N_922,In_357,In_38);
nand U923 (N_923,In_141,In_780);
nor U924 (N_924,In_957,In_289);
nand U925 (N_925,In_993,In_528);
nand U926 (N_926,In_586,In_642);
nor U927 (N_927,In_214,In_451);
and U928 (N_928,In_936,In_430);
nor U929 (N_929,In_43,In_809);
and U930 (N_930,In_50,In_177);
or U931 (N_931,In_77,In_4);
nor U932 (N_932,In_453,In_920);
nand U933 (N_933,In_639,In_710);
or U934 (N_934,In_145,In_572);
or U935 (N_935,In_701,In_651);
nor U936 (N_936,In_317,In_791);
or U937 (N_937,In_902,In_501);
and U938 (N_938,In_700,In_88);
nand U939 (N_939,In_953,In_171);
and U940 (N_940,In_68,In_363);
or U941 (N_941,In_149,In_193);
or U942 (N_942,In_67,In_973);
nor U943 (N_943,In_347,In_968);
and U944 (N_944,In_484,In_525);
nor U945 (N_945,In_873,In_85);
xnor U946 (N_946,In_962,In_252);
nand U947 (N_947,In_845,In_292);
nor U948 (N_948,In_450,In_0);
or U949 (N_949,In_483,In_525);
nor U950 (N_950,In_645,In_560);
xnor U951 (N_951,In_863,In_802);
and U952 (N_952,In_563,In_707);
nor U953 (N_953,In_625,In_642);
and U954 (N_954,In_734,In_323);
and U955 (N_955,In_753,In_545);
nand U956 (N_956,In_365,In_505);
and U957 (N_957,In_298,In_377);
nor U958 (N_958,In_515,In_807);
nor U959 (N_959,In_451,In_170);
nor U960 (N_960,In_290,In_663);
and U961 (N_961,In_871,In_163);
nor U962 (N_962,In_887,In_8);
nand U963 (N_963,In_269,In_25);
and U964 (N_964,In_420,In_910);
or U965 (N_965,In_633,In_299);
nor U966 (N_966,In_650,In_727);
nor U967 (N_967,In_768,In_833);
and U968 (N_968,In_562,In_774);
or U969 (N_969,In_199,In_103);
nand U970 (N_970,In_471,In_863);
or U971 (N_971,In_142,In_368);
or U972 (N_972,In_140,In_544);
or U973 (N_973,In_883,In_603);
and U974 (N_974,In_770,In_470);
and U975 (N_975,In_562,In_678);
nor U976 (N_976,In_726,In_719);
nor U977 (N_977,In_780,In_830);
nor U978 (N_978,In_888,In_220);
nand U979 (N_979,In_208,In_617);
and U980 (N_980,In_863,In_581);
and U981 (N_981,In_467,In_930);
or U982 (N_982,In_46,In_212);
nand U983 (N_983,In_893,In_316);
or U984 (N_984,In_920,In_251);
or U985 (N_985,In_341,In_95);
or U986 (N_986,In_368,In_529);
and U987 (N_987,In_89,In_307);
nor U988 (N_988,In_528,In_165);
and U989 (N_989,In_87,In_416);
nor U990 (N_990,In_77,In_257);
nor U991 (N_991,In_683,In_402);
and U992 (N_992,In_20,In_837);
nand U993 (N_993,In_972,In_754);
nor U994 (N_994,In_95,In_533);
and U995 (N_995,In_224,In_291);
or U996 (N_996,In_885,In_906);
or U997 (N_997,In_556,In_588);
and U998 (N_998,In_826,In_962);
nor U999 (N_999,In_157,In_352);
nor U1000 (N_1000,In_81,In_457);
or U1001 (N_1001,In_292,In_178);
nand U1002 (N_1002,In_630,In_363);
or U1003 (N_1003,In_326,In_264);
nor U1004 (N_1004,In_463,In_714);
nor U1005 (N_1005,In_242,In_900);
and U1006 (N_1006,In_851,In_964);
and U1007 (N_1007,In_64,In_777);
and U1008 (N_1008,In_916,In_671);
nor U1009 (N_1009,In_599,In_39);
xor U1010 (N_1010,In_863,In_899);
or U1011 (N_1011,In_401,In_354);
and U1012 (N_1012,In_696,In_388);
nand U1013 (N_1013,In_696,In_5);
and U1014 (N_1014,In_48,In_77);
nor U1015 (N_1015,In_674,In_135);
and U1016 (N_1016,In_145,In_498);
nand U1017 (N_1017,In_409,In_837);
and U1018 (N_1018,In_590,In_0);
nor U1019 (N_1019,In_612,In_983);
nor U1020 (N_1020,In_718,In_115);
nor U1021 (N_1021,In_0,In_618);
and U1022 (N_1022,In_640,In_322);
nor U1023 (N_1023,In_433,In_642);
and U1024 (N_1024,In_710,In_256);
nand U1025 (N_1025,In_806,In_591);
or U1026 (N_1026,In_741,In_156);
nand U1027 (N_1027,In_489,In_270);
nand U1028 (N_1028,In_421,In_82);
and U1029 (N_1029,In_215,In_71);
or U1030 (N_1030,In_200,In_8);
nand U1031 (N_1031,In_996,In_419);
and U1032 (N_1032,In_507,In_408);
or U1033 (N_1033,In_375,In_803);
nand U1034 (N_1034,In_200,In_237);
nor U1035 (N_1035,In_374,In_840);
or U1036 (N_1036,In_689,In_367);
nor U1037 (N_1037,In_680,In_429);
or U1038 (N_1038,In_428,In_691);
xnor U1039 (N_1039,In_152,In_296);
nand U1040 (N_1040,In_669,In_532);
or U1041 (N_1041,In_50,In_6);
nor U1042 (N_1042,In_357,In_59);
nor U1043 (N_1043,In_832,In_153);
and U1044 (N_1044,In_347,In_266);
or U1045 (N_1045,In_282,In_815);
xnor U1046 (N_1046,In_698,In_959);
nor U1047 (N_1047,In_130,In_473);
nand U1048 (N_1048,In_473,In_428);
nor U1049 (N_1049,In_637,In_441);
nor U1050 (N_1050,In_529,In_589);
nand U1051 (N_1051,In_712,In_480);
xnor U1052 (N_1052,In_177,In_998);
nand U1053 (N_1053,In_838,In_682);
and U1054 (N_1054,In_620,In_832);
and U1055 (N_1055,In_492,In_900);
nand U1056 (N_1056,In_185,In_370);
xnor U1057 (N_1057,In_457,In_492);
or U1058 (N_1058,In_574,In_143);
and U1059 (N_1059,In_800,In_339);
xnor U1060 (N_1060,In_218,In_294);
nor U1061 (N_1061,In_219,In_538);
nor U1062 (N_1062,In_950,In_632);
or U1063 (N_1063,In_931,In_860);
nand U1064 (N_1064,In_692,In_586);
or U1065 (N_1065,In_353,In_802);
nor U1066 (N_1066,In_485,In_339);
nor U1067 (N_1067,In_251,In_766);
and U1068 (N_1068,In_607,In_777);
and U1069 (N_1069,In_685,In_769);
nand U1070 (N_1070,In_398,In_965);
nand U1071 (N_1071,In_895,In_584);
or U1072 (N_1072,In_666,In_911);
nand U1073 (N_1073,In_404,In_171);
nand U1074 (N_1074,In_278,In_880);
nor U1075 (N_1075,In_551,In_6);
nand U1076 (N_1076,In_21,In_793);
or U1077 (N_1077,In_588,In_609);
and U1078 (N_1078,In_951,In_987);
or U1079 (N_1079,In_857,In_738);
nor U1080 (N_1080,In_75,In_114);
nand U1081 (N_1081,In_356,In_384);
nor U1082 (N_1082,In_430,In_526);
and U1083 (N_1083,In_679,In_44);
or U1084 (N_1084,In_262,In_785);
nor U1085 (N_1085,In_908,In_603);
nand U1086 (N_1086,In_166,In_584);
nand U1087 (N_1087,In_490,In_751);
or U1088 (N_1088,In_410,In_162);
or U1089 (N_1089,In_840,In_215);
or U1090 (N_1090,In_411,In_61);
and U1091 (N_1091,In_140,In_734);
or U1092 (N_1092,In_195,In_594);
and U1093 (N_1093,In_641,In_21);
and U1094 (N_1094,In_511,In_993);
or U1095 (N_1095,In_388,In_157);
or U1096 (N_1096,In_862,In_741);
nand U1097 (N_1097,In_294,In_812);
and U1098 (N_1098,In_636,In_223);
nor U1099 (N_1099,In_368,In_477);
nand U1100 (N_1100,In_799,In_845);
or U1101 (N_1101,In_288,In_45);
nand U1102 (N_1102,In_550,In_492);
or U1103 (N_1103,In_231,In_786);
nand U1104 (N_1104,In_790,In_353);
nor U1105 (N_1105,In_205,In_741);
xor U1106 (N_1106,In_301,In_529);
nand U1107 (N_1107,In_952,In_282);
nand U1108 (N_1108,In_34,In_552);
nor U1109 (N_1109,In_642,In_86);
nand U1110 (N_1110,In_815,In_515);
and U1111 (N_1111,In_783,In_371);
nor U1112 (N_1112,In_220,In_479);
nand U1113 (N_1113,In_118,In_670);
nor U1114 (N_1114,In_77,In_422);
nor U1115 (N_1115,In_577,In_662);
or U1116 (N_1116,In_881,In_653);
or U1117 (N_1117,In_788,In_280);
and U1118 (N_1118,In_862,In_128);
or U1119 (N_1119,In_325,In_7);
nor U1120 (N_1120,In_859,In_429);
nor U1121 (N_1121,In_78,In_797);
nand U1122 (N_1122,In_311,In_110);
nand U1123 (N_1123,In_830,In_18);
nor U1124 (N_1124,In_980,In_840);
and U1125 (N_1125,In_284,In_907);
or U1126 (N_1126,In_953,In_248);
and U1127 (N_1127,In_710,In_188);
nand U1128 (N_1128,In_683,In_733);
and U1129 (N_1129,In_482,In_571);
or U1130 (N_1130,In_13,In_753);
or U1131 (N_1131,In_673,In_63);
or U1132 (N_1132,In_827,In_129);
or U1133 (N_1133,In_914,In_122);
and U1134 (N_1134,In_335,In_237);
nand U1135 (N_1135,In_897,In_580);
nor U1136 (N_1136,In_89,In_662);
and U1137 (N_1137,In_360,In_407);
and U1138 (N_1138,In_171,In_113);
nand U1139 (N_1139,In_486,In_66);
nand U1140 (N_1140,In_203,In_998);
xnor U1141 (N_1141,In_445,In_935);
nand U1142 (N_1142,In_659,In_703);
and U1143 (N_1143,In_130,In_918);
or U1144 (N_1144,In_753,In_130);
nor U1145 (N_1145,In_413,In_633);
nor U1146 (N_1146,In_930,In_456);
nand U1147 (N_1147,In_563,In_926);
nand U1148 (N_1148,In_775,In_321);
and U1149 (N_1149,In_463,In_791);
or U1150 (N_1150,In_278,In_907);
nand U1151 (N_1151,In_156,In_91);
and U1152 (N_1152,In_321,In_411);
nor U1153 (N_1153,In_889,In_797);
or U1154 (N_1154,In_378,In_306);
and U1155 (N_1155,In_726,In_776);
nor U1156 (N_1156,In_156,In_703);
xor U1157 (N_1157,In_576,In_64);
nand U1158 (N_1158,In_581,In_874);
nor U1159 (N_1159,In_416,In_438);
and U1160 (N_1160,In_995,In_813);
or U1161 (N_1161,In_148,In_560);
or U1162 (N_1162,In_249,In_993);
nor U1163 (N_1163,In_49,In_262);
nand U1164 (N_1164,In_518,In_874);
and U1165 (N_1165,In_659,In_228);
nor U1166 (N_1166,In_595,In_263);
nand U1167 (N_1167,In_955,In_633);
xnor U1168 (N_1168,In_70,In_386);
or U1169 (N_1169,In_381,In_584);
xor U1170 (N_1170,In_36,In_279);
xnor U1171 (N_1171,In_541,In_607);
or U1172 (N_1172,In_192,In_2);
and U1173 (N_1173,In_70,In_13);
or U1174 (N_1174,In_756,In_712);
nand U1175 (N_1175,In_777,In_209);
and U1176 (N_1176,In_90,In_931);
nor U1177 (N_1177,In_346,In_310);
and U1178 (N_1178,In_665,In_427);
xnor U1179 (N_1179,In_961,In_234);
nand U1180 (N_1180,In_685,In_421);
nand U1181 (N_1181,In_917,In_26);
and U1182 (N_1182,In_191,In_935);
nor U1183 (N_1183,In_932,In_799);
nand U1184 (N_1184,In_670,In_10);
and U1185 (N_1185,In_600,In_705);
and U1186 (N_1186,In_480,In_737);
or U1187 (N_1187,In_907,In_417);
or U1188 (N_1188,In_463,In_498);
or U1189 (N_1189,In_907,In_78);
and U1190 (N_1190,In_42,In_832);
and U1191 (N_1191,In_100,In_652);
or U1192 (N_1192,In_134,In_650);
and U1193 (N_1193,In_406,In_127);
nand U1194 (N_1194,In_648,In_658);
nor U1195 (N_1195,In_655,In_8);
nor U1196 (N_1196,In_122,In_317);
nand U1197 (N_1197,In_783,In_910);
nand U1198 (N_1198,In_933,In_578);
or U1199 (N_1199,In_958,In_394);
or U1200 (N_1200,In_990,In_428);
or U1201 (N_1201,In_146,In_103);
nor U1202 (N_1202,In_939,In_932);
and U1203 (N_1203,In_211,In_198);
and U1204 (N_1204,In_472,In_501);
nand U1205 (N_1205,In_104,In_481);
nor U1206 (N_1206,In_478,In_822);
nor U1207 (N_1207,In_90,In_217);
nor U1208 (N_1208,In_668,In_694);
and U1209 (N_1209,In_779,In_587);
and U1210 (N_1210,In_128,In_168);
nand U1211 (N_1211,In_40,In_988);
nand U1212 (N_1212,In_831,In_578);
and U1213 (N_1213,In_944,In_378);
and U1214 (N_1214,In_399,In_275);
nor U1215 (N_1215,In_748,In_167);
or U1216 (N_1216,In_31,In_766);
nand U1217 (N_1217,In_607,In_287);
nand U1218 (N_1218,In_986,In_687);
nand U1219 (N_1219,In_962,In_749);
nor U1220 (N_1220,In_562,In_287);
and U1221 (N_1221,In_933,In_182);
nor U1222 (N_1222,In_822,In_892);
xnor U1223 (N_1223,In_478,In_796);
nor U1224 (N_1224,In_194,In_176);
and U1225 (N_1225,In_728,In_153);
nor U1226 (N_1226,In_215,In_576);
nand U1227 (N_1227,In_639,In_503);
nor U1228 (N_1228,In_991,In_36);
nand U1229 (N_1229,In_572,In_211);
nor U1230 (N_1230,In_375,In_349);
nor U1231 (N_1231,In_833,In_556);
xor U1232 (N_1232,In_566,In_142);
nor U1233 (N_1233,In_859,In_763);
and U1234 (N_1234,In_177,In_165);
and U1235 (N_1235,In_653,In_0);
and U1236 (N_1236,In_510,In_623);
and U1237 (N_1237,In_519,In_29);
or U1238 (N_1238,In_411,In_266);
nand U1239 (N_1239,In_876,In_119);
nor U1240 (N_1240,In_388,In_985);
nand U1241 (N_1241,In_129,In_768);
and U1242 (N_1242,In_510,In_857);
nor U1243 (N_1243,In_482,In_210);
or U1244 (N_1244,In_467,In_414);
xnor U1245 (N_1245,In_284,In_858);
nand U1246 (N_1246,In_8,In_724);
nand U1247 (N_1247,In_711,In_580);
nor U1248 (N_1248,In_136,In_335);
nor U1249 (N_1249,In_614,In_487);
and U1250 (N_1250,In_911,In_389);
and U1251 (N_1251,In_828,In_926);
nor U1252 (N_1252,In_108,In_46);
nor U1253 (N_1253,In_977,In_80);
nand U1254 (N_1254,In_231,In_504);
nand U1255 (N_1255,In_641,In_32);
nand U1256 (N_1256,In_179,In_584);
nor U1257 (N_1257,In_472,In_317);
or U1258 (N_1258,In_948,In_313);
and U1259 (N_1259,In_638,In_652);
nor U1260 (N_1260,In_227,In_956);
nand U1261 (N_1261,In_212,In_187);
or U1262 (N_1262,In_513,In_228);
and U1263 (N_1263,In_105,In_346);
nor U1264 (N_1264,In_481,In_709);
and U1265 (N_1265,In_279,In_350);
and U1266 (N_1266,In_350,In_814);
nand U1267 (N_1267,In_552,In_829);
nor U1268 (N_1268,In_656,In_943);
nand U1269 (N_1269,In_970,In_622);
or U1270 (N_1270,In_713,In_377);
nor U1271 (N_1271,In_639,In_65);
nand U1272 (N_1272,In_868,In_442);
and U1273 (N_1273,In_379,In_281);
or U1274 (N_1274,In_119,In_554);
or U1275 (N_1275,In_241,In_846);
and U1276 (N_1276,In_482,In_796);
nand U1277 (N_1277,In_647,In_455);
nand U1278 (N_1278,In_619,In_130);
and U1279 (N_1279,In_664,In_459);
and U1280 (N_1280,In_662,In_123);
and U1281 (N_1281,In_129,In_771);
nand U1282 (N_1282,In_691,In_57);
nand U1283 (N_1283,In_636,In_525);
nor U1284 (N_1284,In_696,In_973);
nor U1285 (N_1285,In_708,In_712);
nor U1286 (N_1286,In_35,In_987);
nor U1287 (N_1287,In_188,In_847);
or U1288 (N_1288,In_518,In_444);
and U1289 (N_1289,In_610,In_256);
nor U1290 (N_1290,In_912,In_117);
and U1291 (N_1291,In_815,In_417);
and U1292 (N_1292,In_969,In_364);
nor U1293 (N_1293,In_337,In_681);
and U1294 (N_1294,In_362,In_311);
or U1295 (N_1295,In_950,In_946);
nor U1296 (N_1296,In_654,In_356);
nor U1297 (N_1297,In_105,In_10);
nand U1298 (N_1298,In_673,In_60);
nor U1299 (N_1299,In_11,In_736);
or U1300 (N_1300,In_733,In_444);
and U1301 (N_1301,In_496,In_331);
xor U1302 (N_1302,In_127,In_303);
nand U1303 (N_1303,In_576,In_640);
or U1304 (N_1304,In_4,In_542);
nor U1305 (N_1305,In_333,In_182);
nor U1306 (N_1306,In_609,In_413);
nand U1307 (N_1307,In_163,In_495);
and U1308 (N_1308,In_328,In_212);
and U1309 (N_1309,In_683,In_299);
and U1310 (N_1310,In_468,In_180);
nand U1311 (N_1311,In_308,In_12);
nor U1312 (N_1312,In_188,In_73);
and U1313 (N_1313,In_621,In_552);
nand U1314 (N_1314,In_827,In_198);
or U1315 (N_1315,In_284,In_171);
and U1316 (N_1316,In_71,In_487);
and U1317 (N_1317,In_955,In_836);
nand U1318 (N_1318,In_630,In_331);
and U1319 (N_1319,In_739,In_833);
and U1320 (N_1320,In_131,In_747);
nor U1321 (N_1321,In_255,In_231);
nand U1322 (N_1322,In_813,In_439);
nand U1323 (N_1323,In_869,In_455);
or U1324 (N_1324,In_674,In_678);
nand U1325 (N_1325,In_684,In_776);
or U1326 (N_1326,In_760,In_964);
nand U1327 (N_1327,In_174,In_326);
or U1328 (N_1328,In_880,In_159);
nand U1329 (N_1329,In_521,In_797);
and U1330 (N_1330,In_650,In_342);
nand U1331 (N_1331,In_211,In_186);
and U1332 (N_1332,In_100,In_334);
or U1333 (N_1333,In_17,In_69);
nand U1334 (N_1334,In_44,In_808);
and U1335 (N_1335,In_730,In_622);
or U1336 (N_1336,In_127,In_394);
nor U1337 (N_1337,In_479,In_707);
nor U1338 (N_1338,In_289,In_217);
nand U1339 (N_1339,In_775,In_117);
nor U1340 (N_1340,In_504,In_841);
nand U1341 (N_1341,In_915,In_144);
or U1342 (N_1342,In_526,In_726);
nor U1343 (N_1343,In_444,In_907);
nand U1344 (N_1344,In_232,In_810);
and U1345 (N_1345,In_479,In_662);
and U1346 (N_1346,In_980,In_87);
and U1347 (N_1347,In_718,In_155);
or U1348 (N_1348,In_978,In_836);
or U1349 (N_1349,In_719,In_667);
xor U1350 (N_1350,In_297,In_857);
and U1351 (N_1351,In_770,In_683);
nand U1352 (N_1352,In_490,In_331);
nand U1353 (N_1353,In_756,In_954);
nor U1354 (N_1354,In_392,In_154);
nand U1355 (N_1355,In_267,In_545);
or U1356 (N_1356,In_886,In_65);
or U1357 (N_1357,In_527,In_932);
or U1358 (N_1358,In_406,In_409);
nor U1359 (N_1359,In_206,In_465);
and U1360 (N_1360,In_272,In_540);
xor U1361 (N_1361,In_85,In_43);
nand U1362 (N_1362,In_559,In_456);
and U1363 (N_1363,In_460,In_961);
nand U1364 (N_1364,In_615,In_820);
and U1365 (N_1365,In_379,In_726);
or U1366 (N_1366,In_262,In_17);
and U1367 (N_1367,In_331,In_907);
nand U1368 (N_1368,In_633,In_289);
or U1369 (N_1369,In_328,In_261);
or U1370 (N_1370,In_965,In_622);
nand U1371 (N_1371,In_464,In_42);
and U1372 (N_1372,In_497,In_603);
nand U1373 (N_1373,In_249,In_448);
nor U1374 (N_1374,In_394,In_53);
nand U1375 (N_1375,In_195,In_550);
nand U1376 (N_1376,In_547,In_281);
nor U1377 (N_1377,In_965,In_560);
or U1378 (N_1378,In_1,In_829);
nor U1379 (N_1379,In_70,In_786);
or U1380 (N_1380,In_164,In_53);
and U1381 (N_1381,In_160,In_419);
nand U1382 (N_1382,In_819,In_648);
nand U1383 (N_1383,In_940,In_448);
and U1384 (N_1384,In_292,In_216);
and U1385 (N_1385,In_311,In_498);
nor U1386 (N_1386,In_197,In_450);
nand U1387 (N_1387,In_808,In_167);
nor U1388 (N_1388,In_64,In_718);
and U1389 (N_1389,In_692,In_973);
nor U1390 (N_1390,In_173,In_418);
nand U1391 (N_1391,In_477,In_965);
nand U1392 (N_1392,In_692,In_200);
nand U1393 (N_1393,In_695,In_990);
nand U1394 (N_1394,In_416,In_145);
or U1395 (N_1395,In_821,In_558);
or U1396 (N_1396,In_32,In_474);
or U1397 (N_1397,In_905,In_151);
and U1398 (N_1398,In_529,In_432);
or U1399 (N_1399,In_390,In_911);
and U1400 (N_1400,In_864,In_229);
or U1401 (N_1401,In_179,In_714);
and U1402 (N_1402,In_164,In_969);
nand U1403 (N_1403,In_337,In_80);
and U1404 (N_1404,In_666,In_764);
or U1405 (N_1405,In_110,In_182);
and U1406 (N_1406,In_493,In_444);
or U1407 (N_1407,In_990,In_460);
and U1408 (N_1408,In_164,In_850);
xor U1409 (N_1409,In_413,In_919);
or U1410 (N_1410,In_284,In_971);
nand U1411 (N_1411,In_332,In_749);
or U1412 (N_1412,In_832,In_472);
nand U1413 (N_1413,In_350,In_320);
and U1414 (N_1414,In_616,In_322);
and U1415 (N_1415,In_178,In_184);
nor U1416 (N_1416,In_716,In_57);
nor U1417 (N_1417,In_924,In_975);
nor U1418 (N_1418,In_196,In_596);
or U1419 (N_1419,In_594,In_29);
nand U1420 (N_1420,In_18,In_329);
and U1421 (N_1421,In_457,In_897);
and U1422 (N_1422,In_431,In_256);
and U1423 (N_1423,In_939,In_97);
nand U1424 (N_1424,In_511,In_261);
nand U1425 (N_1425,In_140,In_485);
and U1426 (N_1426,In_300,In_245);
nand U1427 (N_1427,In_264,In_752);
or U1428 (N_1428,In_263,In_771);
or U1429 (N_1429,In_536,In_854);
nor U1430 (N_1430,In_556,In_497);
nand U1431 (N_1431,In_161,In_650);
or U1432 (N_1432,In_821,In_481);
nand U1433 (N_1433,In_852,In_103);
and U1434 (N_1434,In_214,In_668);
and U1435 (N_1435,In_317,In_231);
nand U1436 (N_1436,In_557,In_457);
and U1437 (N_1437,In_556,In_252);
or U1438 (N_1438,In_219,In_306);
nand U1439 (N_1439,In_632,In_726);
and U1440 (N_1440,In_150,In_493);
and U1441 (N_1441,In_652,In_579);
or U1442 (N_1442,In_815,In_956);
nor U1443 (N_1443,In_886,In_879);
nand U1444 (N_1444,In_890,In_610);
nand U1445 (N_1445,In_64,In_764);
and U1446 (N_1446,In_397,In_947);
nor U1447 (N_1447,In_575,In_950);
xnor U1448 (N_1448,In_77,In_721);
or U1449 (N_1449,In_678,In_433);
or U1450 (N_1450,In_574,In_4);
nor U1451 (N_1451,In_31,In_985);
nand U1452 (N_1452,In_563,In_785);
nor U1453 (N_1453,In_931,In_960);
or U1454 (N_1454,In_211,In_353);
and U1455 (N_1455,In_544,In_130);
nor U1456 (N_1456,In_785,In_231);
or U1457 (N_1457,In_197,In_489);
nand U1458 (N_1458,In_231,In_517);
and U1459 (N_1459,In_197,In_881);
nand U1460 (N_1460,In_919,In_272);
and U1461 (N_1461,In_610,In_90);
nor U1462 (N_1462,In_283,In_454);
or U1463 (N_1463,In_93,In_976);
and U1464 (N_1464,In_944,In_458);
or U1465 (N_1465,In_464,In_157);
and U1466 (N_1466,In_852,In_539);
or U1467 (N_1467,In_515,In_114);
or U1468 (N_1468,In_829,In_408);
or U1469 (N_1469,In_639,In_215);
nand U1470 (N_1470,In_133,In_703);
nand U1471 (N_1471,In_284,In_688);
and U1472 (N_1472,In_139,In_491);
nand U1473 (N_1473,In_373,In_936);
nor U1474 (N_1474,In_170,In_711);
and U1475 (N_1475,In_410,In_789);
nand U1476 (N_1476,In_816,In_825);
nand U1477 (N_1477,In_536,In_206);
or U1478 (N_1478,In_332,In_884);
nand U1479 (N_1479,In_419,In_755);
nand U1480 (N_1480,In_143,In_735);
nor U1481 (N_1481,In_295,In_149);
nor U1482 (N_1482,In_297,In_920);
or U1483 (N_1483,In_485,In_488);
or U1484 (N_1484,In_64,In_59);
nand U1485 (N_1485,In_128,In_288);
and U1486 (N_1486,In_563,In_191);
and U1487 (N_1487,In_712,In_135);
and U1488 (N_1488,In_531,In_270);
and U1489 (N_1489,In_171,In_126);
nand U1490 (N_1490,In_562,In_489);
xnor U1491 (N_1491,In_560,In_829);
nand U1492 (N_1492,In_230,In_919);
nand U1493 (N_1493,In_162,In_538);
and U1494 (N_1494,In_552,In_905);
and U1495 (N_1495,In_343,In_213);
xor U1496 (N_1496,In_956,In_606);
nor U1497 (N_1497,In_696,In_461);
nor U1498 (N_1498,In_680,In_128);
or U1499 (N_1499,In_682,In_120);
nor U1500 (N_1500,In_777,In_856);
or U1501 (N_1501,In_301,In_706);
and U1502 (N_1502,In_649,In_957);
nand U1503 (N_1503,In_237,In_8);
or U1504 (N_1504,In_635,In_923);
or U1505 (N_1505,In_594,In_622);
and U1506 (N_1506,In_985,In_435);
or U1507 (N_1507,In_672,In_975);
nand U1508 (N_1508,In_355,In_799);
nor U1509 (N_1509,In_288,In_198);
nor U1510 (N_1510,In_846,In_760);
nand U1511 (N_1511,In_864,In_669);
and U1512 (N_1512,In_307,In_297);
and U1513 (N_1513,In_712,In_729);
nor U1514 (N_1514,In_130,In_910);
nor U1515 (N_1515,In_952,In_349);
nor U1516 (N_1516,In_780,In_424);
xnor U1517 (N_1517,In_656,In_806);
or U1518 (N_1518,In_231,In_550);
nand U1519 (N_1519,In_835,In_738);
nand U1520 (N_1520,In_494,In_520);
or U1521 (N_1521,In_466,In_44);
and U1522 (N_1522,In_341,In_271);
nor U1523 (N_1523,In_147,In_724);
and U1524 (N_1524,In_108,In_57);
or U1525 (N_1525,In_555,In_553);
nor U1526 (N_1526,In_347,In_798);
or U1527 (N_1527,In_165,In_0);
or U1528 (N_1528,In_692,In_593);
nand U1529 (N_1529,In_433,In_858);
nor U1530 (N_1530,In_404,In_946);
or U1531 (N_1531,In_514,In_386);
and U1532 (N_1532,In_895,In_273);
and U1533 (N_1533,In_4,In_58);
or U1534 (N_1534,In_958,In_268);
or U1535 (N_1535,In_484,In_535);
and U1536 (N_1536,In_484,In_701);
or U1537 (N_1537,In_400,In_742);
and U1538 (N_1538,In_83,In_192);
nand U1539 (N_1539,In_448,In_32);
or U1540 (N_1540,In_653,In_295);
and U1541 (N_1541,In_862,In_642);
nor U1542 (N_1542,In_547,In_729);
or U1543 (N_1543,In_816,In_773);
xor U1544 (N_1544,In_413,In_93);
xor U1545 (N_1545,In_239,In_167);
and U1546 (N_1546,In_975,In_890);
or U1547 (N_1547,In_689,In_196);
or U1548 (N_1548,In_66,In_852);
nand U1549 (N_1549,In_639,In_795);
and U1550 (N_1550,In_674,In_235);
and U1551 (N_1551,In_565,In_80);
and U1552 (N_1552,In_790,In_185);
and U1553 (N_1553,In_141,In_914);
or U1554 (N_1554,In_842,In_896);
and U1555 (N_1555,In_29,In_809);
and U1556 (N_1556,In_996,In_166);
nor U1557 (N_1557,In_185,In_984);
and U1558 (N_1558,In_448,In_183);
or U1559 (N_1559,In_233,In_888);
or U1560 (N_1560,In_523,In_398);
nand U1561 (N_1561,In_908,In_616);
and U1562 (N_1562,In_997,In_968);
or U1563 (N_1563,In_740,In_410);
or U1564 (N_1564,In_835,In_799);
nand U1565 (N_1565,In_921,In_881);
and U1566 (N_1566,In_644,In_342);
nand U1567 (N_1567,In_497,In_6);
nand U1568 (N_1568,In_787,In_93);
or U1569 (N_1569,In_373,In_894);
nor U1570 (N_1570,In_627,In_861);
and U1571 (N_1571,In_477,In_541);
nor U1572 (N_1572,In_891,In_92);
nor U1573 (N_1573,In_470,In_482);
or U1574 (N_1574,In_405,In_925);
and U1575 (N_1575,In_539,In_991);
nand U1576 (N_1576,In_871,In_562);
nor U1577 (N_1577,In_756,In_440);
xnor U1578 (N_1578,In_517,In_640);
nor U1579 (N_1579,In_873,In_765);
xnor U1580 (N_1580,In_525,In_794);
nand U1581 (N_1581,In_804,In_909);
nand U1582 (N_1582,In_517,In_671);
or U1583 (N_1583,In_505,In_374);
and U1584 (N_1584,In_443,In_999);
or U1585 (N_1585,In_455,In_272);
nor U1586 (N_1586,In_941,In_192);
nor U1587 (N_1587,In_958,In_367);
nor U1588 (N_1588,In_474,In_231);
or U1589 (N_1589,In_440,In_449);
and U1590 (N_1590,In_311,In_682);
or U1591 (N_1591,In_513,In_395);
nor U1592 (N_1592,In_827,In_375);
nand U1593 (N_1593,In_663,In_941);
and U1594 (N_1594,In_78,In_801);
nor U1595 (N_1595,In_130,In_485);
nand U1596 (N_1596,In_351,In_18);
nand U1597 (N_1597,In_107,In_923);
and U1598 (N_1598,In_800,In_16);
nand U1599 (N_1599,In_769,In_811);
and U1600 (N_1600,In_214,In_8);
nand U1601 (N_1601,In_208,In_913);
and U1602 (N_1602,In_754,In_348);
nor U1603 (N_1603,In_230,In_422);
nor U1604 (N_1604,In_49,In_451);
nor U1605 (N_1605,In_303,In_448);
nor U1606 (N_1606,In_975,In_376);
nor U1607 (N_1607,In_830,In_82);
nand U1608 (N_1608,In_326,In_838);
and U1609 (N_1609,In_429,In_77);
or U1610 (N_1610,In_362,In_596);
nor U1611 (N_1611,In_773,In_152);
nor U1612 (N_1612,In_799,In_848);
nand U1613 (N_1613,In_891,In_570);
and U1614 (N_1614,In_115,In_653);
nor U1615 (N_1615,In_561,In_606);
nor U1616 (N_1616,In_448,In_653);
nor U1617 (N_1617,In_367,In_903);
xnor U1618 (N_1618,In_100,In_742);
nand U1619 (N_1619,In_495,In_855);
and U1620 (N_1620,In_469,In_301);
nor U1621 (N_1621,In_858,In_129);
nor U1622 (N_1622,In_293,In_696);
nand U1623 (N_1623,In_765,In_955);
and U1624 (N_1624,In_979,In_833);
nand U1625 (N_1625,In_302,In_19);
xnor U1626 (N_1626,In_798,In_897);
nand U1627 (N_1627,In_461,In_334);
nor U1628 (N_1628,In_448,In_928);
nor U1629 (N_1629,In_510,In_346);
nand U1630 (N_1630,In_937,In_999);
and U1631 (N_1631,In_107,In_548);
and U1632 (N_1632,In_444,In_552);
and U1633 (N_1633,In_722,In_990);
nand U1634 (N_1634,In_701,In_158);
or U1635 (N_1635,In_558,In_578);
or U1636 (N_1636,In_404,In_31);
nor U1637 (N_1637,In_158,In_850);
or U1638 (N_1638,In_429,In_706);
nor U1639 (N_1639,In_357,In_688);
nor U1640 (N_1640,In_148,In_916);
and U1641 (N_1641,In_959,In_884);
or U1642 (N_1642,In_468,In_421);
nor U1643 (N_1643,In_280,In_427);
nor U1644 (N_1644,In_988,In_345);
or U1645 (N_1645,In_615,In_689);
or U1646 (N_1646,In_490,In_240);
or U1647 (N_1647,In_950,In_966);
or U1648 (N_1648,In_684,In_405);
or U1649 (N_1649,In_946,In_957);
or U1650 (N_1650,In_230,In_784);
and U1651 (N_1651,In_262,In_745);
nor U1652 (N_1652,In_607,In_285);
nor U1653 (N_1653,In_359,In_389);
nor U1654 (N_1654,In_521,In_341);
and U1655 (N_1655,In_410,In_477);
nand U1656 (N_1656,In_707,In_732);
nand U1657 (N_1657,In_838,In_788);
nor U1658 (N_1658,In_173,In_627);
and U1659 (N_1659,In_281,In_705);
xnor U1660 (N_1660,In_521,In_598);
nor U1661 (N_1661,In_882,In_331);
nor U1662 (N_1662,In_640,In_151);
nand U1663 (N_1663,In_997,In_989);
nor U1664 (N_1664,In_170,In_846);
and U1665 (N_1665,In_566,In_332);
nor U1666 (N_1666,In_40,In_810);
or U1667 (N_1667,In_314,In_159);
or U1668 (N_1668,In_68,In_639);
or U1669 (N_1669,In_294,In_239);
or U1670 (N_1670,In_760,In_713);
and U1671 (N_1671,In_424,In_210);
nor U1672 (N_1672,In_382,In_330);
nor U1673 (N_1673,In_407,In_240);
and U1674 (N_1674,In_967,In_851);
or U1675 (N_1675,In_781,In_948);
and U1676 (N_1676,In_526,In_519);
nand U1677 (N_1677,In_766,In_227);
or U1678 (N_1678,In_495,In_607);
nand U1679 (N_1679,In_717,In_311);
and U1680 (N_1680,In_724,In_833);
or U1681 (N_1681,In_278,In_259);
and U1682 (N_1682,In_926,In_21);
nand U1683 (N_1683,In_192,In_916);
and U1684 (N_1684,In_712,In_447);
or U1685 (N_1685,In_12,In_790);
and U1686 (N_1686,In_988,In_597);
and U1687 (N_1687,In_940,In_838);
nand U1688 (N_1688,In_425,In_274);
or U1689 (N_1689,In_508,In_941);
and U1690 (N_1690,In_889,In_357);
nor U1691 (N_1691,In_532,In_813);
nor U1692 (N_1692,In_436,In_264);
nand U1693 (N_1693,In_347,In_613);
nand U1694 (N_1694,In_43,In_411);
and U1695 (N_1695,In_562,In_667);
or U1696 (N_1696,In_698,In_746);
and U1697 (N_1697,In_697,In_848);
or U1698 (N_1698,In_240,In_696);
and U1699 (N_1699,In_289,In_246);
and U1700 (N_1700,In_178,In_495);
nor U1701 (N_1701,In_424,In_341);
or U1702 (N_1702,In_453,In_63);
or U1703 (N_1703,In_458,In_763);
nor U1704 (N_1704,In_329,In_691);
and U1705 (N_1705,In_795,In_916);
or U1706 (N_1706,In_393,In_40);
nor U1707 (N_1707,In_357,In_232);
nor U1708 (N_1708,In_744,In_350);
or U1709 (N_1709,In_640,In_698);
or U1710 (N_1710,In_166,In_265);
or U1711 (N_1711,In_859,In_366);
or U1712 (N_1712,In_163,In_823);
nor U1713 (N_1713,In_420,In_743);
or U1714 (N_1714,In_33,In_399);
or U1715 (N_1715,In_276,In_343);
nand U1716 (N_1716,In_44,In_286);
and U1717 (N_1717,In_820,In_974);
nor U1718 (N_1718,In_993,In_113);
nor U1719 (N_1719,In_670,In_244);
nand U1720 (N_1720,In_720,In_497);
and U1721 (N_1721,In_425,In_493);
nor U1722 (N_1722,In_379,In_452);
or U1723 (N_1723,In_890,In_640);
nand U1724 (N_1724,In_697,In_822);
and U1725 (N_1725,In_796,In_648);
nor U1726 (N_1726,In_473,In_712);
or U1727 (N_1727,In_501,In_685);
or U1728 (N_1728,In_987,In_458);
nand U1729 (N_1729,In_33,In_412);
or U1730 (N_1730,In_309,In_901);
or U1731 (N_1731,In_230,In_356);
nand U1732 (N_1732,In_230,In_162);
nand U1733 (N_1733,In_682,In_844);
or U1734 (N_1734,In_642,In_224);
nor U1735 (N_1735,In_652,In_406);
nor U1736 (N_1736,In_600,In_780);
nand U1737 (N_1737,In_562,In_258);
nor U1738 (N_1738,In_950,In_912);
nor U1739 (N_1739,In_182,In_60);
nand U1740 (N_1740,In_896,In_332);
nand U1741 (N_1741,In_487,In_478);
or U1742 (N_1742,In_559,In_2);
nand U1743 (N_1743,In_115,In_344);
nor U1744 (N_1744,In_206,In_61);
and U1745 (N_1745,In_605,In_982);
or U1746 (N_1746,In_864,In_364);
or U1747 (N_1747,In_656,In_645);
nor U1748 (N_1748,In_873,In_37);
or U1749 (N_1749,In_905,In_162);
and U1750 (N_1750,In_245,In_121);
and U1751 (N_1751,In_971,In_54);
nor U1752 (N_1752,In_467,In_33);
nor U1753 (N_1753,In_545,In_385);
and U1754 (N_1754,In_274,In_830);
and U1755 (N_1755,In_223,In_468);
nand U1756 (N_1756,In_49,In_671);
or U1757 (N_1757,In_809,In_841);
or U1758 (N_1758,In_756,In_781);
or U1759 (N_1759,In_229,In_913);
or U1760 (N_1760,In_206,In_706);
nor U1761 (N_1761,In_796,In_475);
nand U1762 (N_1762,In_51,In_85);
or U1763 (N_1763,In_976,In_950);
and U1764 (N_1764,In_53,In_191);
nor U1765 (N_1765,In_919,In_627);
or U1766 (N_1766,In_284,In_341);
nor U1767 (N_1767,In_526,In_559);
nor U1768 (N_1768,In_869,In_689);
nand U1769 (N_1769,In_643,In_632);
and U1770 (N_1770,In_654,In_947);
and U1771 (N_1771,In_198,In_792);
or U1772 (N_1772,In_851,In_650);
nor U1773 (N_1773,In_672,In_411);
nor U1774 (N_1774,In_48,In_170);
nor U1775 (N_1775,In_795,In_285);
or U1776 (N_1776,In_576,In_47);
nand U1777 (N_1777,In_694,In_92);
nand U1778 (N_1778,In_291,In_484);
nand U1779 (N_1779,In_792,In_548);
nand U1780 (N_1780,In_413,In_977);
xor U1781 (N_1781,In_708,In_967);
or U1782 (N_1782,In_55,In_137);
nand U1783 (N_1783,In_16,In_775);
nor U1784 (N_1784,In_269,In_787);
nand U1785 (N_1785,In_224,In_758);
or U1786 (N_1786,In_608,In_757);
nor U1787 (N_1787,In_205,In_187);
nor U1788 (N_1788,In_633,In_332);
and U1789 (N_1789,In_85,In_912);
nor U1790 (N_1790,In_838,In_806);
nor U1791 (N_1791,In_83,In_977);
and U1792 (N_1792,In_628,In_577);
or U1793 (N_1793,In_874,In_855);
nand U1794 (N_1794,In_480,In_880);
and U1795 (N_1795,In_205,In_975);
nor U1796 (N_1796,In_542,In_128);
nand U1797 (N_1797,In_371,In_543);
and U1798 (N_1798,In_902,In_418);
nor U1799 (N_1799,In_72,In_226);
and U1800 (N_1800,In_482,In_373);
and U1801 (N_1801,In_838,In_567);
or U1802 (N_1802,In_860,In_756);
nand U1803 (N_1803,In_765,In_139);
or U1804 (N_1804,In_42,In_118);
and U1805 (N_1805,In_130,In_613);
nor U1806 (N_1806,In_997,In_252);
or U1807 (N_1807,In_822,In_674);
nor U1808 (N_1808,In_633,In_346);
and U1809 (N_1809,In_491,In_947);
or U1810 (N_1810,In_275,In_769);
nand U1811 (N_1811,In_479,In_568);
nor U1812 (N_1812,In_971,In_615);
nor U1813 (N_1813,In_383,In_547);
and U1814 (N_1814,In_799,In_881);
and U1815 (N_1815,In_983,In_827);
or U1816 (N_1816,In_475,In_107);
nor U1817 (N_1817,In_355,In_925);
or U1818 (N_1818,In_201,In_335);
and U1819 (N_1819,In_481,In_774);
or U1820 (N_1820,In_333,In_759);
nor U1821 (N_1821,In_307,In_181);
or U1822 (N_1822,In_189,In_466);
or U1823 (N_1823,In_571,In_612);
nor U1824 (N_1824,In_175,In_925);
and U1825 (N_1825,In_775,In_762);
nand U1826 (N_1826,In_214,In_783);
or U1827 (N_1827,In_227,In_728);
and U1828 (N_1828,In_82,In_696);
nor U1829 (N_1829,In_524,In_820);
or U1830 (N_1830,In_684,In_476);
nor U1831 (N_1831,In_464,In_223);
and U1832 (N_1832,In_141,In_190);
and U1833 (N_1833,In_153,In_858);
and U1834 (N_1834,In_79,In_972);
and U1835 (N_1835,In_104,In_812);
nor U1836 (N_1836,In_160,In_551);
or U1837 (N_1837,In_213,In_315);
nor U1838 (N_1838,In_693,In_775);
nand U1839 (N_1839,In_946,In_377);
or U1840 (N_1840,In_911,In_553);
and U1841 (N_1841,In_579,In_205);
nand U1842 (N_1842,In_999,In_468);
nor U1843 (N_1843,In_177,In_221);
nand U1844 (N_1844,In_213,In_846);
nor U1845 (N_1845,In_301,In_537);
nand U1846 (N_1846,In_190,In_611);
nand U1847 (N_1847,In_656,In_616);
nor U1848 (N_1848,In_451,In_54);
or U1849 (N_1849,In_190,In_564);
or U1850 (N_1850,In_596,In_437);
or U1851 (N_1851,In_545,In_7);
nand U1852 (N_1852,In_536,In_181);
or U1853 (N_1853,In_420,In_80);
or U1854 (N_1854,In_641,In_204);
nor U1855 (N_1855,In_926,In_840);
nor U1856 (N_1856,In_221,In_74);
nor U1857 (N_1857,In_530,In_224);
or U1858 (N_1858,In_448,In_834);
nor U1859 (N_1859,In_742,In_221);
nand U1860 (N_1860,In_531,In_543);
nor U1861 (N_1861,In_939,In_362);
nand U1862 (N_1862,In_322,In_586);
or U1863 (N_1863,In_155,In_559);
nor U1864 (N_1864,In_885,In_635);
nor U1865 (N_1865,In_325,In_763);
and U1866 (N_1866,In_544,In_26);
nor U1867 (N_1867,In_302,In_162);
or U1868 (N_1868,In_929,In_696);
and U1869 (N_1869,In_753,In_609);
nand U1870 (N_1870,In_922,In_995);
nor U1871 (N_1871,In_259,In_448);
nand U1872 (N_1872,In_756,In_585);
and U1873 (N_1873,In_369,In_926);
nor U1874 (N_1874,In_693,In_208);
or U1875 (N_1875,In_933,In_160);
and U1876 (N_1876,In_858,In_9);
or U1877 (N_1877,In_396,In_457);
nand U1878 (N_1878,In_667,In_852);
nor U1879 (N_1879,In_199,In_483);
nand U1880 (N_1880,In_776,In_26);
or U1881 (N_1881,In_819,In_724);
nor U1882 (N_1882,In_759,In_973);
nor U1883 (N_1883,In_70,In_329);
and U1884 (N_1884,In_533,In_587);
nor U1885 (N_1885,In_168,In_21);
or U1886 (N_1886,In_826,In_950);
or U1887 (N_1887,In_228,In_948);
nand U1888 (N_1888,In_62,In_661);
nand U1889 (N_1889,In_260,In_519);
nor U1890 (N_1890,In_417,In_376);
nor U1891 (N_1891,In_914,In_204);
nand U1892 (N_1892,In_203,In_93);
or U1893 (N_1893,In_570,In_145);
and U1894 (N_1894,In_176,In_834);
and U1895 (N_1895,In_517,In_143);
or U1896 (N_1896,In_846,In_909);
and U1897 (N_1897,In_946,In_656);
and U1898 (N_1898,In_134,In_757);
nand U1899 (N_1899,In_313,In_325);
or U1900 (N_1900,In_745,In_564);
nand U1901 (N_1901,In_604,In_917);
and U1902 (N_1902,In_191,In_26);
nand U1903 (N_1903,In_169,In_585);
and U1904 (N_1904,In_860,In_531);
nand U1905 (N_1905,In_379,In_676);
and U1906 (N_1906,In_266,In_226);
or U1907 (N_1907,In_48,In_540);
or U1908 (N_1908,In_183,In_764);
xor U1909 (N_1909,In_545,In_77);
nor U1910 (N_1910,In_400,In_309);
nor U1911 (N_1911,In_558,In_733);
nand U1912 (N_1912,In_60,In_541);
or U1913 (N_1913,In_670,In_536);
nand U1914 (N_1914,In_538,In_308);
and U1915 (N_1915,In_479,In_197);
xor U1916 (N_1916,In_32,In_213);
nor U1917 (N_1917,In_920,In_284);
nor U1918 (N_1918,In_431,In_673);
nand U1919 (N_1919,In_950,In_540);
nor U1920 (N_1920,In_668,In_795);
or U1921 (N_1921,In_998,In_322);
nand U1922 (N_1922,In_409,In_401);
and U1923 (N_1923,In_183,In_361);
or U1924 (N_1924,In_93,In_542);
nand U1925 (N_1925,In_503,In_919);
nor U1926 (N_1926,In_64,In_591);
or U1927 (N_1927,In_163,In_963);
or U1928 (N_1928,In_737,In_263);
or U1929 (N_1929,In_164,In_672);
nor U1930 (N_1930,In_502,In_948);
and U1931 (N_1931,In_997,In_504);
or U1932 (N_1932,In_166,In_461);
and U1933 (N_1933,In_759,In_144);
nor U1934 (N_1934,In_441,In_97);
nor U1935 (N_1935,In_859,In_124);
nor U1936 (N_1936,In_791,In_832);
nand U1937 (N_1937,In_801,In_921);
or U1938 (N_1938,In_982,In_135);
and U1939 (N_1939,In_866,In_460);
nand U1940 (N_1940,In_876,In_900);
nor U1941 (N_1941,In_207,In_177);
nor U1942 (N_1942,In_168,In_336);
nand U1943 (N_1943,In_747,In_32);
and U1944 (N_1944,In_844,In_470);
nor U1945 (N_1945,In_862,In_644);
nand U1946 (N_1946,In_75,In_955);
nor U1947 (N_1947,In_468,In_484);
or U1948 (N_1948,In_400,In_569);
nor U1949 (N_1949,In_75,In_268);
nand U1950 (N_1950,In_308,In_649);
nand U1951 (N_1951,In_139,In_826);
or U1952 (N_1952,In_755,In_816);
nor U1953 (N_1953,In_975,In_937);
or U1954 (N_1954,In_401,In_621);
nand U1955 (N_1955,In_340,In_468);
or U1956 (N_1956,In_631,In_524);
nor U1957 (N_1957,In_766,In_324);
or U1958 (N_1958,In_690,In_827);
and U1959 (N_1959,In_761,In_633);
or U1960 (N_1960,In_661,In_718);
and U1961 (N_1961,In_300,In_59);
nand U1962 (N_1962,In_425,In_737);
nand U1963 (N_1963,In_598,In_187);
nand U1964 (N_1964,In_468,In_29);
nand U1965 (N_1965,In_418,In_283);
nor U1966 (N_1966,In_41,In_372);
nand U1967 (N_1967,In_773,In_225);
nand U1968 (N_1968,In_373,In_912);
and U1969 (N_1969,In_660,In_348);
nor U1970 (N_1970,In_746,In_695);
xnor U1971 (N_1971,In_957,In_488);
and U1972 (N_1972,In_147,In_984);
nor U1973 (N_1973,In_337,In_167);
nand U1974 (N_1974,In_259,In_655);
nor U1975 (N_1975,In_363,In_920);
nand U1976 (N_1976,In_746,In_307);
and U1977 (N_1977,In_867,In_285);
nor U1978 (N_1978,In_91,In_60);
nor U1979 (N_1979,In_349,In_262);
nor U1980 (N_1980,In_22,In_88);
nand U1981 (N_1981,In_203,In_152);
xor U1982 (N_1982,In_998,In_726);
nand U1983 (N_1983,In_504,In_777);
nand U1984 (N_1984,In_140,In_852);
or U1985 (N_1985,In_802,In_871);
or U1986 (N_1986,In_690,In_991);
and U1987 (N_1987,In_773,In_969);
nand U1988 (N_1988,In_195,In_751);
and U1989 (N_1989,In_394,In_839);
nor U1990 (N_1990,In_603,In_294);
or U1991 (N_1991,In_410,In_67);
or U1992 (N_1992,In_125,In_853);
nand U1993 (N_1993,In_720,In_183);
and U1994 (N_1994,In_241,In_107);
nand U1995 (N_1995,In_382,In_643);
nand U1996 (N_1996,In_158,In_101);
and U1997 (N_1997,In_172,In_942);
nand U1998 (N_1998,In_171,In_968);
nor U1999 (N_1999,In_951,In_250);
nand U2000 (N_2000,In_210,In_179);
nand U2001 (N_2001,In_911,In_460);
or U2002 (N_2002,In_838,In_730);
and U2003 (N_2003,In_210,In_719);
and U2004 (N_2004,In_137,In_79);
nor U2005 (N_2005,In_461,In_712);
nand U2006 (N_2006,In_976,In_224);
and U2007 (N_2007,In_738,In_863);
nand U2008 (N_2008,In_992,In_681);
xnor U2009 (N_2009,In_494,In_375);
or U2010 (N_2010,In_637,In_678);
and U2011 (N_2011,In_451,In_924);
nand U2012 (N_2012,In_423,In_615);
and U2013 (N_2013,In_174,In_760);
and U2014 (N_2014,In_609,In_253);
or U2015 (N_2015,In_363,In_170);
or U2016 (N_2016,In_797,In_158);
and U2017 (N_2017,In_402,In_71);
and U2018 (N_2018,In_635,In_823);
or U2019 (N_2019,In_694,In_30);
nand U2020 (N_2020,In_631,In_100);
and U2021 (N_2021,In_468,In_525);
or U2022 (N_2022,In_254,In_459);
or U2023 (N_2023,In_230,In_785);
and U2024 (N_2024,In_374,In_9);
nor U2025 (N_2025,In_141,In_873);
nand U2026 (N_2026,In_277,In_451);
or U2027 (N_2027,In_658,In_134);
nor U2028 (N_2028,In_860,In_431);
and U2029 (N_2029,In_226,In_36);
or U2030 (N_2030,In_809,In_297);
or U2031 (N_2031,In_791,In_574);
or U2032 (N_2032,In_314,In_69);
or U2033 (N_2033,In_644,In_120);
xnor U2034 (N_2034,In_345,In_998);
nor U2035 (N_2035,In_993,In_220);
nor U2036 (N_2036,In_437,In_363);
nand U2037 (N_2037,In_414,In_430);
nand U2038 (N_2038,In_916,In_821);
or U2039 (N_2039,In_837,In_863);
nand U2040 (N_2040,In_495,In_529);
nand U2041 (N_2041,In_890,In_272);
nor U2042 (N_2042,In_649,In_832);
and U2043 (N_2043,In_567,In_728);
nand U2044 (N_2044,In_777,In_573);
nor U2045 (N_2045,In_825,In_65);
and U2046 (N_2046,In_472,In_291);
nor U2047 (N_2047,In_852,In_308);
or U2048 (N_2048,In_624,In_375);
or U2049 (N_2049,In_658,In_217);
nor U2050 (N_2050,In_89,In_204);
and U2051 (N_2051,In_951,In_404);
and U2052 (N_2052,In_852,In_890);
nor U2053 (N_2053,In_618,In_277);
nor U2054 (N_2054,In_41,In_870);
and U2055 (N_2055,In_843,In_566);
nor U2056 (N_2056,In_432,In_442);
and U2057 (N_2057,In_230,In_287);
and U2058 (N_2058,In_427,In_430);
nand U2059 (N_2059,In_744,In_684);
nor U2060 (N_2060,In_202,In_19);
and U2061 (N_2061,In_790,In_272);
nor U2062 (N_2062,In_739,In_170);
nor U2063 (N_2063,In_714,In_987);
or U2064 (N_2064,In_301,In_149);
and U2065 (N_2065,In_264,In_568);
nor U2066 (N_2066,In_202,In_816);
nand U2067 (N_2067,In_320,In_587);
nor U2068 (N_2068,In_958,In_729);
xnor U2069 (N_2069,In_655,In_489);
and U2070 (N_2070,In_105,In_163);
and U2071 (N_2071,In_402,In_77);
or U2072 (N_2072,In_456,In_628);
or U2073 (N_2073,In_745,In_665);
or U2074 (N_2074,In_267,In_143);
xnor U2075 (N_2075,In_507,In_148);
or U2076 (N_2076,In_283,In_883);
and U2077 (N_2077,In_45,In_116);
or U2078 (N_2078,In_604,In_261);
nor U2079 (N_2079,In_158,In_112);
or U2080 (N_2080,In_757,In_16);
nor U2081 (N_2081,In_249,In_750);
nand U2082 (N_2082,In_438,In_213);
or U2083 (N_2083,In_610,In_806);
nor U2084 (N_2084,In_348,In_675);
and U2085 (N_2085,In_931,In_619);
and U2086 (N_2086,In_498,In_274);
and U2087 (N_2087,In_438,In_342);
and U2088 (N_2088,In_845,In_828);
nor U2089 (N_2089,In_27,In_384);
and U2090 (N_2090,In_283,In_880);
and U2091 (N_2091,In_320,In_287);
nand U2092 (N_2092,In_192,In_953);
nor U2093 (N_2093,In_337,In_210);
or U2094 (N_2094,In_164,In_359);
nand U2095 (N_2095,In_928,In_131);
and U2096 (N_2096,In_971,In_658);
or U2097 (N_2097,In_60,In_162);
or U2098 (N_2098,In_385,In_788);
nand U2099 (N_2099,In_562,In_72);
nor U2100 (N_2100,In_611,In_247);
and U2101 (N_2101,In_398,In_825);
nor U2102 (N_2102,In_89,In_551);
nand U2103 (N_2103,In_2,In_824);
and U2104 (N_2104,In_31,In_887);
nor U2105 (N_2105,In_968,In_425);
nor U2106 (N_2106,In_815,In_343);
and U2107 (N_2107,In_341,In_440);
nor U2108 (N_2108,In_792,In_333);
or U2109 (N_2109,In_150,In_490);
or U2110 (N_2110,In_759,In_546);
nor U2111 (N_2111,In_396,In_173);
nand U2112 (N_2112,In_879,In_594);
and U2113 (N_2113,In_520,In_607);
nand U2114 (N_2114,In_721,In_475);
nand U2115 (N_2115,In_839,In_119);
and U2116 (N_2116,In_274,In_822);
or U2117 (N_2117,In_813,In_267);
xor U2118 (N_2118,In_405,In_449);
and U2119 (N_2119,In_395,In_811);
or U2120 (N_2120,In_243,In_389);
xor U2121 (N_2121,In_506,In_310);
nand U2122 (N_2122,In_669,In_277);
and U2123 (N_2123,In_843,In_883);
nand U2124 (N_2124,In_737,In_168);
or U2125 (N_2125,In_457,In_840);
or U2126 (N_2126,In_253,In_595);
nand U2127 (N_2127,In_156,In_917);
or U2128 (N_2128,In_847,In_700);
nand U2129 (N_2129,In_506,In_252);
xor U2130 (N_2130,In_275,In_205);
nand U2131 (N_2131,In_912,In_723);
and U2132 (N_2132,In_541,In_429);
or U2133 (N_2133,In_354,In_613);
or U2134 (N_2134,In_903,In_930);
and U2135 (N_2135,In_872,In_530);
nor U2136 (N_2136,In_302,In_361);
xnor U2137 (N_2137,In_365,In_346);
or U2138 (N_2138,In_48,In_769);
nand U2139 (N_2139,In_986,In_909);
or U2140 (N_2140,In_430,In_857);
nor U2141 (N_2141,In_966,In_501);
or U2142 (N_2142,In_359,In_67);
or U2143 (N_2143,In_830,In_631);
and U2144 (N_2144,In_831,In_209);
nor U2145 (N_2145,In_949,In_620);
and U2146 (N_2146,In_60,In_271);
nand U2147 (N_2147,In_824,In_167);
nand U2148 (N_2148,In_777,In_897);
and U2149 (N_2149,In_386,In_357);
nand U2150 (N_2150,In_96,In_952);
nor U2151 (N_2151,In_854,In_335);
or U2152 (N_2152,In_398,In_265);
or U2153 (N_2153,In_428,In_803);
nand U2154 (N_2154,In_786,In_547);
nor U2155 (N_2155,In_898,In_841);
nand U2156 (N_2156,In_856,In_974);
xor U2157 (N_2157,In_318,In_325);
nor U2158 (N_2158,In_333,In_209);
or U2159 (N_2159,In_225,In_14);
nand U2160 (N_2160,In_719,In_983);
and U2161 (N_2161,In_768,In_252);
nand U2162 (N_2162,In_395,In_314);
nor U2163 (N_2163,In_733,In_959);
nand U2164 (N_2164,In_211,In_945);
and U2165 (N_2165,In_798,In_743);
nand U2166 (N_2166,In_148,In_455);
and U2167 (N_2167,In_947,In_29);
nor U2168 (N_2168,In_999,In_904);
xor U2169 (N_2169,In_110,In_657);
or U2170 (N_2170,In_167,In_927);
nand U2171 (N_2171,In_906,In_130);
nand U2172 (N_2172,In_118,In_320);
nor U2173 (N_2173,In_688,In_107);
and U2174 (N_2174,In_857,In_876);
nand U2175 (N_2175,In_460,In_592);
and U2176 (N_2176,In_530,In_799);
or U2177 (N_2177,In_307,In_848);
and U2178 (N_2178,In_421,In_454);
or U2179 (N_2179,In_73,In_294);
and U2180 (N_2180,In_722,In_713);
or U2181 (N_2181,In_477,In_148);
or U2182 (N_2182,In_874,In_217);
nand U2183 (N_2183,In_835,In_701);
or U2184 (N_2184,In_26,In_669);
nand U2185 (N_2185,In_997,In_478);
nor U2186 (N_2186,In_146,In_271);
xor U2187 (N_2187,In_483,In_219);
nand U2188 (N_2188,In_736,In_376);
nand U2189 (N_2189,In_987,In_630);
or U2190 (N_2190,In_543,In_80);
or U2191 (N_2191,In_763,In_281);
nand U2192 (N_2192,In_791,In_247);
and U2193 (N_2193,In_914,In_703);
nor U2194 (N_2194,In_747,In_871);
and U2195 (N_2195,In_803,In_609);
or U2196 (N_2196,In_292,In_302);
nand U2197 (N_2197,In_965,In_369);
nand U2198 (N_2198,In_975,In_181);
xnor U2199 (N_2199,In_19,In_572);
and U2200 (N_2200,In_689,In_317);
and U2201 (N_2201,In_518,In_904);
and U2202 (N_2202,In_236,In_828);
and U2203 (N_2203,In_59,In_419);
or U2204 (N_2204,In_73,In_775);
or U2205 (N_2205,In_5,In_483);
and U2206 (N_2206,In_982,In_850);
xor U2207 (N_2207,In_730,In_6);
or U2208 (N_2208,In_277,In_825);
nand U2209 (N_2209,In_119,In_234);
nand U2210 (N_2210,In_332,In_404);
and U2211 (N_2211,In_24,In_508);
or U2212 (N_2212,In_388,In_150);
nor U2213 (N_2213,In_256,In_547);
nand U2214 (N_2214,In_577,In_501);
nor U2215 (N_2215,In_390,In_874);
and U2216 (N_2216,In_808,In_560);
nand U2217 (N_2217,In_555,In_310);
and U2218 (N_2218,In_523,In_982);
nor U2219 (N_2219,In_171,In_72);
or U2220 (N_2220,In_582,In_969);
nand U2221 (N_2221,In_14,In_53);
or U2222 (N_2222,In_392,In_104);
and U2223 (N_2223,In_953,In_76);
nor U2224 (N_2224,In_596,In_541);
and U2225 (N_2225,In_554,In_482);
and U2226 (N_2226,In_81,In_652);
or U2227 (N_2227,In_913,In_894);
and U2228 (N_2228,In_875,In_324);
nor U2229 (N_2229,In_839,In_815);
nand U2230 (N_2230,In_434,In_772);
nand U2231 (N_2231,In_620,In_779);
or U2232 (N_2232,In_346,In_654);
xnor U2233 (N_2233,In_155,In_933);
and U2234 (N_2234,In_250,In_737);
or U2235 (N_2235,In_690,In_115);
nor U2236 (N_2236,In_412,In_862);
and U2237 (N_2237,In_598,In_675);
nor U2238 (N_2238,In_689,In_385);
xor U2239 (N_2239,In_308,In_574);
and U2240 (N_2240,In_405,In_821);
and U2241 (N_2241,In_278,In_962);
and U2242 (N_2242,In_390,In_357);
or U2243 (N_2243,In_316,In_634);
or U2244 (N_2244,In_622,In_491);
nand U2245 (N_2245,In_694,In_761);
nand U2246 (N_2246,In_224,In_270);
or U2247 (N_2247,In_50,In_169);
xnor U2248 (N_2248,In_553,In_994);
or U2249 (N_2249,In_474,In_496);
and U2250 (N_2250,In_46,In_846);
or U2251 (N_2251,In_410,In_955);
or U2252 (N_2252,In_616,In_205);
nand U2253 (N_2253,In_350,In_937);
and U2254 (N_2254,In_144,In_652);
nand U2255 (N_2255,In_239,In_223);
nor U2256 (N_2256,In_145,In_55);
nor U2257 (N_2257,In_106,In_969);
nor U2258 (N_2258,In_743,In_464);
and U2259 (N_2259,In_875,In_373);
or U2260 (N_2260,In_800,In_591);
or U2261 (N_2261,In_426,In_111);
and U2262 (N_2262,In_372,In_882);
or U2263 (N_2263,In_114,In_987);
nor U2264 (N_2264,In_520,In_0);
or U2265 (N_2265,In_112,In_613);
and U2266 (N_2266,In_247,In_504);
or U2267 (N_2267,In_723,In_428);
or U2268 (N_2268,In_533,In_373);
nand U2269 (N_2269,In_131,In_298);
or U2270 (N_2270,In_795,In_337);
and U2271 (N_2271,In_247,In_838);
and U2272 (N_2272,In_215,In_562);
nor U2273 (N_2273,In_440,In_763);
nor U2274 (N_2274,In_14,In_198);
or U2275 (N_2275,In_569,In_6);
nor U2276 (N_2276,In_549,In_321);
or U2277 (N_2277,In_849,In_165);
and U2278 (N_2278,In_484,In_991);
and U2279 (N_2279,In_716,In_924);
nand U2280 (N_2280,In_211,In_340);
nor U2281 (N_2281,In_203,In_66);
nand U2282 (N_2282,In_523,In_541);
and U2283 (N_2283,In_152,In_149);
nor U2284 (N_2284,In_844,In_82);
or U2285 (N_2285,In_147,In_808);
nand U2286 (N_2286,In_475,In_535);
nor U2287 (N_2287,In_702,In_921);
or U2288 (N_2288,In_152,In_681);
and U2289 (N_2289,In_591,In_529);
xnor U2290 (N_2290,In_568,In_936);
nand U2291 (N_2291,In_699,In_445);
nor U2292 (N_2292,In_238,In_886);
and U2293 (N_2293,In_913,In_839);
nand U2294 (N_2294,In_252,In_186);
and U2295 (N_2295,In_526,In_367);
or U2296 (N_2296,In_897,In_634);
nand U2297 (N_2297,In_90,In_851);
nand U2298 (N_2298,In_279,In_106);
nand U2299 (N_2299,In_268,In_808);
nand U2300 (N_2300,In_517,In_506);
and U2301 (N_2301,In_896,In_816);
or U2302 (N_2302,In_999,In_801);
nand U2303 (N_2303,In_412,In_577);
nand U2304 (N_2304,In_817,In_437);
nand U2305 (N_2305,In_608,In_951);
nand U2306 (N_2306,In_286,In_31);
or U2307 (N_2307,In_378,In_258);
and U2308 (N_2308,In_807,In_196);
nor U2309 (N_2309,In_372,In_821);
and U2310 (N_2310,In_279,In_517);
and U2311 (N_2311,In_396,In_221);
or U2312 (N_2312,In_249,In_778);
nor U2313 (N_2313,In_811,In_835);
nand U2314 (N_2314,In_800,In_502);
or U2315 (N_2315,In_435,In_62);
and U2316 (N_2316,In_424,In_548);
nand U2317 (N_2317,In_267,In_850);
and U2318 (N_2318,In_256,In_983);
nand U2319 (N_2319,In_514,In_371);
and U2320 (N_2320,In_217,In_293);
nand U2321 (N_2321,In_814,In_294);
nand U2322 (N_2322,In_302,In_994);
and U2323 (N_2323,In_998,In_670);
nand U2324 (N_2324,In_456,In_994);
nor U2325 (N_2325,In_459,In_493);
or U2326 (N_2326,In_780,In_476);
nor U2327 (N_2327,In_936,In_144);
nand U2328 (N_2328,In_588,In_176);
or U2329 (N_2329,In_476,In_870);
or U2330 (N_2330,In_227,In_987);
nand U2331 (N_2331,In_255,In_603);
or U2332 (N_2332,In_556,In_620);
nor U2333 (N_2333,In_99,In_62);
nand U2334 (N_2334,In_484,In_34);
nand U2335 (N_2335,In_133,In_243);
nor U2336 (N_2336,In_483,In_865);
nor U2337 (N_2337,In_796,In_213);
and U2338 (N_2338,In_220,In_233);
or U2339 (N_2339,In_246,In_906);
or U2340 (N_2340,In_845,In_418);
nor U2341 (N_2341,In_143,In_289);
or U2342 (N_2342,In_602,In_332);
and U2343 (N_2343,In_588,In_865);
xnor U2344 (N_2344,In_705,In_667);
nor U2345 (N_2345,In_997,In_575);
nand U2346 (N_2346,In_588,In_855);
nand U2347 (N_2347,In_70,In_740);
nor U2348 (N_2348,In_114,In_720);
nor U2349 (N_2349,In_37,In_84);
and U2350 (N_2350,In_204,In_560);
and U2351 (N_2351,In_738,In_922);
and U2352 (N_2352,In_983,In_473);
or U2353 (N_2353,In_58,In_120);
and U2354 (N_2354,In_865,In_781);
or U2355 (N_2355,In_162,In_964);
nor U2356 (N_2356,In_469,In_6);
nand U2357 (N_2357,In_331,In_730);
or U2358 (N_2358,In_600,In_35);
and U2359 (N_2359,In_21,In_485);
nor U2360 (N_2360,In_165,In_123);
nor U2361 (N_2361,In_288,In_990);
nand U2362 (N_2362,In_32,In_374);
or U2363 (N_2363,In_235,In_640);
nand U2364 (N_2364,In_937,In_450);
nand U2365 (N_2365,In_43,In_610);
nor U2366 (N_2366,In_699,In_231);
and U2367 (N_2367,In_943,In_102);
nand U2368 (N_2368,In_431,In_122);
nor U2369 (N_2369,In_771,In_72);
nor U2370 (N_2370,In_733,In_484);
and U2371 (N_2371,In_558,In_962);
nand U2372 (N_2372,In_74,In_194);
or U2373 (N_2373,In_499,In_315);
or U2374 (N_2374,In_781,In_206);
or U2375 (N_2375,In_730,In_769);
nand U2376 (N_2376,In_174,In_670);
nor U2377 (N_2377,In_731,In_560);
nand U2378 (N_2378,In_972,In_604);
nand U2379 (N_2379,In_120,In_487);
or U2380 (N_2380,In_983,In_405);
xor U2381 (N_2381,In_368,In_878);
and U2382 (N_2382,In_496,In_820);
or U2383 (N_2383,In_55,In_928);
nand U2384 (N_2384,In_961,In_599);
nand U2385 (N_2385,In_208,In_385);
nand U2386 (N_2386,In_389,In_150);
or U2387 (N_2387,In_665,In_855);
xor U2388 (N_2388,In_222,In_200);
nor U2389 (N_2389,In_236,In_363);
nor U2390 (N_2390,In_912,In_702);
nor U2391 (N_2391,In_5,In_517);
nand U2392 (N_2392,In_993,In_248);
or U2393 (N_2393,In_294,In_4);
nor U2394 (N_2394,In_225,In_623);
nand U2395 (N_2395,In_129,In_892);
xnor U2396 (N_2396,In_306,In_604);
nand U2397 (N_2397,In_913,In_704);
or U2398 (N_2398,In_405,In_486);
or U2399 (N_2399,In_459,In_89);
xor U2400 (N_2400,In_888,In_482);
nor U2401 (N_2401,In_810,In_200);
xnor U2402 (N_2402,In_873,In_407);
or U2403 (N_2403,In_275,In_585);
nand U2404 (N_2404,In_48,In_612);
or U2405 (N_2405,In_221,In_849);
or U2406 (N_2406,In_329,In_720);
and U2407 (N_2407,In_523,In_865);
nor U2408 (N_2408,In_778,In_704);
and U2409 (N_2409,In_552,In_221);
xor U2410 (N_2410,In_332,In_19);
nor U2411 (N_2411,In_137,In_232);
nor U2412 (N_2412,In_280,In_597);
nand U2413 (N_2413,In_197,In_570);
xor U2414 (N_2414,In_382,In_942);
and U2415 (N_2415,In_20,In_921);
nor U2416 (N_2416,In_270,In_215);
xor U2417 (N_2417,In_73,In_454);
or U2418 (N_2418,In_463,In_856);
or U2419 (N_2419,In_371,In_281);
nand U2420 (N_2420,In_233,In_75);
and U2421 (N_2421,In_947,In_196);
nor U2422 (N_2422,In_121,In_741);
nand U2423 (N_2423,In_910,In_656);
nand U2424 (N_2424,In_736,In_155);
nor U2425 (N_2425,In_446,In_664);
nand U2426 (N_2426,In_173,In_474);
or U2427 (N_2427,In_595,In_30);
or U2428 (N_2428,In_949,In_84);
nor U2429 (N_2429,In_680,In_859);
nor U2430 (N_2430,In_899,In_801);
or U2431 (N_2431,In_113,In_18);
or U2432 (N_2432,In_415,In_802);
xnor U2433 (N_2433,In_219,In_402);
nand U2434 (N_2434,In_280,In_120);
nor U2435 (N_2435,In_746,In_72);
nor U2436 (N_2436,In_277,In_77);
nand U2437 (N_2437,In_108,In_288);
and U2438 (N_2438,In_103,In_379);
nand U2439 (N_2439,In_497,In_280);
nand U2440 (N_2440,In_832,In_537);
nor U2441 (N_2441,In_359,In_719);
nor U2442 (N_2442,In_399,In_122);
nor U2443 (N_2443,In_869,In_507);
and U2444 (N_2444,In_524,In_645);
nand U2445 (N_2445,In_78,In_793);
nand U2446 (N_2446,In_93,In_119);
nor U2447 (N_2447,In_73,In_111);
and U2448 (N_2448,In_797,In_904);
nor U2449 (N_2449,In_745,In_124);
xnor U2450 (N_2450,In_137,In_860);
nand U2451 (N_2451,In_503,In_2);
and U2452 (N_2452,In_407,In_343);
or U2453 (N_2453,In_360,In_904);
nor U2454 (N_2454,In_943,In_714);
nand U2455 (N_2455,In_568,In_412);
nand U2456 (N_2456,In_283,In_875);
or U2457 (N_2457,In_245,In_555);
nand U2458 (N_2458,In_207,In_246);
nor U2459 (N_2459,In_431,In_391);
nand U2460 (N_2460,In_23,In_908);
and U2461 (N_2461,In_245,In_452);
nand U2462 (N_2462,In_662,In_617);
nor U2463 (N_2463,In_632,In_454);
nand U2464 (N_2464,In_229,In_244);
nor U2465 (N_2465,In_497,In_606);
or U2466 (N_2466,In_8,In_723);
and U2467 (N_2467,In_342,In_562);
and U2468 (N_2468,In_85,In_964);
nand U2469 (N_2469,In_707,In_667);
and U2470 (N_2470,In_264,In_592);
or U2471 (N_2471,In_938,In_995);
nand U2472 (N_2472,In_936,In_883);
and U2473 (N_2473,In_330,In_304);
nor U2474 (N_2474,In_468,In_868);
or U2475 (N_2475,In_418,In_137);
xor U2476 (N_2476,In_500,In_258);
nand U2477 (N_2477,In_655,In_983);
nand U2478 (N_2478,In_369,In_559);
nor U2479 (N_2479,In_9,In_591);
or U2480 (N_2480,In_697,In_343);
nor U2481 (N_2481,In_730,In_976);
or U2482 (N_2482,In_952,In_547);
nor U2483 (N_2483,In_293,In_463);
nand U2484 (N_2484,In_692,In_306);
nor U2485 (N_2485,In_301,In_204);
nor U2486 (N_2486,In_206,In_62);
nand U2487 (N_2487,In_854,In_5);
or U2488 (N_2488,In_216,In_438);
or U2489 (N_2489,In_873,In_264);
or U2490 (N_2490,In_653,In_980);
or U2491 (N_2491,In_922,In_364);
and U2492 (N_2492,In_579,In_313);
or U2493 (N_2493,In_471,In_661);
nor U2494 (N_2494,In_558,In_787);
or U2495 (N_2495,In_202,In_688);
nand U2496 (N_2496,In_613,In_844);
nor U2497 (N_2497,In_838,In_304);
or U2498 (N_2498,In_59,In_322);
nand U2499 (N_2499,In_889,In_98);
or U2500 (N_2500,In_75,In_522);
and U2501 (N_2501,In_590,In_883);
or U2502 (N_2502,In_786,In_985);
and U2503 (N_2503,In_236,In_946);
nor U2504 (N_2504,In_260,In_630);
nor U2505 (N_2505,In_236,In_708);
and U2506 (N_2506,In_90,In_250);
and U2507 (N_2507,In_190,In_221);
and U2508 (N_2508,In_747,In_29);
nor U2509 (N_2509,In_920,In_270);
nand U2510 (N_2510,In_463,In_19);
or U2511 (N_2511,In_722,In_155);
nor U2512 (N_2512,In_745,In_399);
nor U2513 (N_2513,In_500,In_276);
nor U2514 (N_2514,In_360,In_274);
nor U2515 (N_2515,In_878,In_107);
or U2516 (N_2516,In_986,In_945);
and U2517 (N_2517,In_958,In_480);
nand U2518 (N_2518,In_666,In_52);
or U2519 (N_2519,In_994,In_889);
nor U2520 (N_2520,In_866,In_439);
nand U2521 (N_2521,In_813,In_556);
or U2522 (N_2522,In_117,In_321);
nor U2523 (N_2523,In_453,In_751);
nand U2524 (N_2524,In_785,In_695);
xor U2525 (N_2525,In_937,In_284);
or U2526 (N_2526,In_550,In_461);
nand U2527 (N_2527,In_579,In_329);
nand U2528 (N_2528,In_335,In_748);
or U2529 (N_2529,In_586,In_344);
or U2530 (N_2530,In_210,In_65);
and U2531 (N_2531,In_910,In_577);
nor U2532 (N_2532,In_585,In_100);
nand U2533 (N_2533,In_439,In_312);
and U2534 (N_2534,In_508,In_124);
nor U2535 (N_2535,In_461,In_291);
or U2536 (N_2536,In_7,In_293);
nand U2537 (N_2537,In_915,In_700);
nor U2538 (N_2538,In_852,In_734);
xor U2539 (N_2539,In_423,In_88);
xor U2540 (N_2540,In_838,In_142);
nand U2541 (N_2541,In_943,In_606);
nand U2542 (N_2542,In_106,In_733);
nand U2543 (N_2543,In_702,In_197);
and U2544 (N_2544,In_260,In_262);
and U2545 (N_2545,In_501,In_334);
or U2546 (N_2546,In_441,In_414);
or U2547 (N_2547,In_968,In_680);
and U2548 (N_2548,In_151,In_915);
and U2549 (N_2549,In_616,In_54);
nand U2550 (N_2550,In_170,In_840);
nor U2551 (N_2551,In_284,In_246);
nor U2552 (N_2552,In_792,In_900);
and U2553 (N_2553,In_605,In_180);
and U2554 (N_2554,In_859,In_33);
nor U2555 (N_2555,In_263,In_978);
and U2556 (N_2556,In_859,In_823);
and U2557 (N_2557,In_774,In_259);
or U2558 (N_2558,In_183,In_701);
and U2559 (N_2559,In_595,In_303);
and U2560 (N_2560,In_926,In_558);
or U2561 (N_2561,In_793,In_405);
nand U2562 (N_2562,In_45,In_236);
or U2563 (N_2563,In_374,In_399);
and U2564 (N_2564,In_836,In_205);
and U2565 (N_2565,In_421,In_709);
nor U2566 (N_2566,In_875,In_235);
or U2567 (N_2567,In_455,In_99);
or U2568 (N_2568,In_867,In_777);
or U2569 (N_2569,In_210,In_409);
nor U2570 (N_2570,In_483,In_35);
and U2571 (N_2571,In_648,In_15);
and U2572 (N_2572,In_991,In_360);
and U2573 (N_2573,In_718,In_98);
xnor U2574 (N_2574,In_934,In_531);
and U2575 (N_2575,In_313,In_36);
or U2576 (N_2576,In_463,In_397);
or U2577 (N_2577,In_492,In_969);
nand U2578 (N_2578,In_845,In_232);
or U2579 (N_2579,In_825,In_248);
nor U2580 (N_2580,In_42,In_898);
nand U2581 (N_2581,In_741,In_458);
nor U2582 (N_2582,In_479,In_905);
nor U2583 (N_2583,In_456,In_49);
or U2584 (N_2584,In_429,In_858);
nand U2585 (N_2585,In_999,In_739);
or U2586 (N_2586,In_698,In_661);
nor U2587 (N_2587,In_854,In_150);
nand U2588 (N_2588,In_335,In_557);
nand U2589 (N_2589,In_391,In_700);
nand U2590 (N_2590,In_662,In_166);
or U2591 (N_2591,In_121,In_176);
nor U2592 (N_2592,In_282,In_758);
nor U2593 (N_2593,In_191,In_255);
or U2594 (N_2594,In_592,In_959);
and U2595 (N_2595,In_867,In_395);
nand U2596 (N_2596,In_243,In_279);
and U2597 (N_2597,In_79,In_494);
and U2598 (N_2598,In_450,In_621);
and U2599 (N_2599,In_451,In_640);
or U2600 (N_2600,In_399,In_203);
nand U2601 (N_2601,In_384,In_404);
nor U2602 (N_2602,In_53,In_26);
nand U2603 (N_2603,In_526,In_277);
and U2604 (N_2604,In_417,In_226);
nor U2605 (N_2605,In_448,In_532);
and U2606 (N_2606,In_560,In_200);
nand U2607 (N_2607,In_736,In_846);
and U2608 (N_2608,In_321,In_124);
nand U2609 (N_2609,In_83,In_544);
nand U2610 (N_2610,In_389,In_432);
nor U2611 (N_2611,In_968,In_925);
and U2612 (N_2612,In_738,In_945);
and U2613 (N_2613,In_805,In_296);
or U2614 (N_2614,In_177,In_274);
nor U2615 (N_2615,In_733,In_884);
and U2616 (N_2616,In_662,In_947);
or U2617 (N_2617,In_944,In_812);
nor U2618 (N_2618,In_894,In_630);
or U2619 (N_2619,In_309,In_255);
and U2620 (N_2620,In_695,In_837);
nor U2621 (N_2621,In_492,In_632);
nand U2622 (N_2622,In_964,In_289);
nand U2623 (N_2623,In_364,In_138);
nand U2624 (N_2624,In_835,In_866);
nand U2625 (N_2625,In_979,In_482);
nand U2626 (N_2626,In_119,In_607);
and U2627 (N_2627,In_994,In_617);
and U2628 (N_2628,In_373,In_519);
and U2629 (N_2629,In_280,In_350);
nor U2630 (N_2630,In_815,In_840);
nor U2631 (N_2631,In_389,In_973);
xnor U2632 (N_2632,In_356,In_618);
or U2633 (N_2633,In_612,In_676);
nand U2634 (N_2634,In_176,In_739);
nor U2635 (N_2635,In_799,In_674);
nand U2636 (N_2636,In_352,In_410);
or U2637 (N_2637,In_581,In_467);
or U2638 (N_2638,In_377,In_257);
and U2639 (N_2639,In_451,In_110);
nor U2640 (N_2640,In_42,In_505);
and U2641 (N_2641,In_351,In_702);
xnor U2642 (N_2642,In_561,In_213);
or U2643 (N_2643,In_457,In_495);
and U2644 (N_2644,In_805,In_532);
nor U2645 (N_2645,In_745,In_31);
nand U2646 (N_2646,In_231,In_853);
or U2647 (N_2647,In_364,In_921);
or U2648 (N_2648,In_850,In_46);
or U2649 (N_2649,In_334,In_397);
and U2650 (N_2650,In_383,In_631);
or U2651 (N_2651,In_670,In_822);
nor U2652 (N_2652,In_356,In_84);
and U2653 (N_2653,In_169,In_426);
nor U2654 (N_2654,In_736,In_955);
or U2655 (N_2655,In_446,In_509);
nand U2656 (N_2656,In_683,In_667);
xnor U2657 (N_2657,In_847,In_325);
nand U2658 (N_2658,In_552,In_634);
nor U2659 (N_2659,In_277,In_830);
nor U2660 (N_2660,In_86,In_247);
nor U2661 (N_2661,In_826,In_809);
and U2662 (N_2662,In_928,In_307);
or U2663 (N_2663,In_261,In_108);
nor U2664 (N_2664,In_961,In_897);
and U2665 (N_2665,In_136,In_682);
nand U2666 (N_2666,In_309,In_517);
and U2667 (N_2667,In_994,In_804);
or U2668 (N_2668,In_722,In_772);
and U2669 (N_2669,In_161,In_309);
or U2670 (N_2670,In_16,In_847);
and U2671 (N_2671,In_550,In_102);
and U2672 (N_2672,In_316,In_262);
xor U2673 (N_2673,In_979,In_863);
nor U2674 (N_2674,In_653,In_732);
or U2675 (N_2675,In_59,In_153);
and U2676 (N_2676,In_665,In_267);
nor U2677 (N_2677,In_192,In_187);
and U2678 (N_2678,In_708,In_883);
nand U2679 (N_2679,In_363,In_795);
nand U2680 (N_2680,In_126,In_573);
nor U2681 (N_2681,In_193,In_262);
nor U2682 (N_2682,In_300,In_724);
nor U2683 (N_2683,In_580,In_203);
or U2684 (N_2684,In_762,In_360);
or U2685 (N_2685,In_51,In_774);
and U2686 (N_2686,In_872,In_801);
and U2687 (N_2687,In_977,In_161);
nor U2688 (N_2688,In_740,In_800);
and U2689 (N_2689,In_257,In_661);
and U2690 (N_2690,In_856,In_570);
nand U2691 (N_2691,In_105,In_119);
or U2692 (N_2692,In_198,In_881);
or U2693 (N_2693,In_715,In_686);
and U2694 (N_2694,In_281,In_388);
or U2695 (N_2695,In_655,In_961);
or U2696 (N_2696,In_396,In_526);
and U2697 (N_2697,In_329,In_243);
and U2698 (N_2698,In_329,In_316);
nor U2699 (N_2699,In_48,In_594);
nor U2700 (N_2700,In_27,In_647);
and U2701 (N_2701,In_360,In_86);
nor U2702 (N_2702,In_198,In_573);
and U2703 (N_2703,In_966,In_715);
or U2704 (N_2704,In_572,In_559);
or U2705 (N_2705,In_714,In_214);
nor U2706 (N_2706,In_74,In_502);
nor U2707 (N_2707,In_166,In_325);
nor U2708 (N_2708,In_270,In_389);
nor U2709 (N_2709,In_545,In_177);
xor U2710 (N_2710,In_737,In_431);
nand U2711 (N_2711,In_91,In_333);
and U2712 (N_2712,In_716,In_425);
nor U2713 (N_2713,In_891,In_503);
nor U2714 (N_2714,In_603,In_580);
nor U2715 (N_2715,In_341,In_664);
nor U2716 (N_2716,In_314,In_912);
nor U2717 (N_2717,In_198,In_884);
and U2718 (N_2718,In_837,In_482);
nand U2719 (N_2719,In_198,In_48);
or U2720 (N_2720,In_242,In_502);
xnor U2721 (N_2721,In_888,In_804);
nor U2722 (N_2722,In_791,In_104);
nand U2723 (N_2723,In_238,In_737);
or U2724 (N_2724,In_377,In_778);
nand U2725 (N_2725,In_546,In_470);
nand U2726 (N_2726,In_834,In_545);
nand U2727 (N_2727,In_400,In_41);
nor U2728 (N_2728,In_669,In_586);
and U2729 (N_2729,In_142,In_987);
or U2730 (N_2730,In_256,In_303);
and U2731 (N_2731,In_869,In_420);
nand U2732 (N_2732,In_579,In_52);
nand U2733 (N_2733,In_722,In_780);
or U2734 (N_2734,In_592,In_427);
or U2735 (N_2735,In_350,In_587);
or U2736 (N_2736,In_155,In_779);
nor U2737 (N_2737,In_524,In_86);
and U2738 (N_2738,In_325,In_791);
nand U2739 (N_2739,In_159,In_35);
or U2740 (N_2740,In_552,In_202);
nor U2741 (N_2741,In_614,In_79);
xor U2742 (N_2742,In_968,In_281);
or U2743 (N_2743,In_34,In_750);
nor U2744 (N_2744,In_680,In_230);
nor U2745 (N_2745,In_101,In_392);
nor U2746 (N_2746,In_561,In_705);
nand U2747 (N_2747,In_959,In_725);
nand U2748 (N_2748,In_689,In_352);
or U2749 (N_2749,In_301,In_106);
or U2750 (N_2750,In_433,In_640);
nand U2751 (N_2751,In_576,In_549);
nor U2752 (N_2752,In_476,In_696);
and U2753 (N_2753,In_404,In_514);
and U2754 (N_2754,In_382,In_894);
or U2755 (N_2755,In_276,In_744);
nor U2756 (N_2756,In_400,In_330);
or U2757 (N_2757,In_861,In_473);
or U2758 (N_2758,In_76,In_581);
and U2759 (N_2759,In_241,In_155);
and U2760 (N_2760,In_141,In_480);
and U2761 (N_2761,In_467,In_169);
or U2762 (N_2762,In_824,In_105);
nor U2763 (N_2763,In_238,In_239);
nor U2764 (N_2764,In_807,In_152);
and U2765 (N_2765,In_159,In_431);
xor U2766 (N_2766,In_295,In_501);
nand U2767 (N_2767,In_12,In_732);
nor U2768 (N_2768,In_515,In_73);
nand U2769 (N_2769,In_577,In_98);
or U2770 (N_2770,In_684,In_153);
nand U2771 (N_2771,In_870,In_320);
nand U2772 (N_2772,In_699,In_391);
nor U2773 (N_2773,In_148,In_631);
nor U2774 (N_2774,In_573,In_807);
and U2775 (N_2775,In_241,In_424);
nor U2776 (N_2776,In_344,In_693);
or U2777 (N_2777,In_648,In_496);
or U2778 (N_2778,In_356,In_295);
or U2779 (N_2779,In_25,In_465);
or U2780 (N_2780,In_5,In_132);
nor U2781 (N_2781,In_28,In_696);
or U2782 (N_2782,In_966,In_720);
nor U2783 (N_2783,In_786,In_963);
or U2784 (N_2784,In_634,In_639);
nand U2785 (N_2785,In_47,In_117);
nor U2786 (N_2786,In_281,In_997);
nor U2787 (N_2787,In_745,In_626);
nor U2788 (N_2788,In_961,In_230);
nand U2789 (N_2789,In_525,In_818);
nand U2790 (N_2790,In_463,In_24);
or U2791 (N_2791,In_414,In_292);
nor U2792 (N_2792,In_916,In_501);
nand U2793 (N_2793,In_28,In_765);
and U2794 (N_2794,In_23,In_873);
nand U2795 (N_2795,In_979,In_702);
nand U2796 (N_2796,In_723,In_847);
nor U2797 (N_2797,In_812,In_915);
or U2798 (N_2798,In_809,In_300);
nor U2799 (N_2799,In_928,In_7);
nand U2800 (N_2800,In_80,In_266);
or U2801 (N_2801,In_875,In_574);
or U2802 (N_2802,In_261,In_528);
and U2803 (N_2803,In_305,In_849);
nor U2804 (N_2804,In_108,In_837);
or U2805 (N_2805,In_491,In_785);
nor U2806 (N_2806,In_18,In_497);
and U2807 (N_2807,In_819,In_434);
or U2808 (N_2808,In_101,In_716);
and U2809 (N_2809,In_723,In_825);
and U2810 (N_2810,In_832,In_871);
nand U2811 (N_2811,In_542,In_451);
and U2812 (N_2812,In_807,In_423);
xnor U2813 (N_2813,In_237,In_620);
nand U2814 (N_2814,In_561,In_274);
or U2815 (N_2815,In_504,In_174);
and U2816 (N_2816,In_834,In_112);
nand U2817 (N_2817,In_609,In_0);
nand U2818 (N_2818,In_853,In_883);
and U2819 (N_2819,In_382,In_713);
or U2820 (N_2820,In_411,In_329);
and U2821 (N_2821,In_104,In_668);
or U2822 (N_2822,In_233,In_316);
nand U2823 (N_2823,In_300,In_265);
or U2824 (N_2824,In_455,In_322);
or U2825 (N_2825,In_296,In_197);
xnor U2826 (N_2826,In_463,In_474);
nor U2827 (N_2827,In_361,In_479);
or U2828 (N_2828,In_893,In_129);
and U2829 (N_2829,In_58,In_569);
or U2830 (N_2830,In_745,In_602);
nor U2831 (N_2831,In_405,In_228);
or U2832 (N_2832,In_764,In_340);
and U2833 (N_2833,In_597,In_918);
nand U2834 (N_2834,In_386,In_552);
nand U2835 (N_2835,In_509,In_365);
or U2836 (N_2836,In_469,In_641);
nand U2837 (N_2837,In_321,In_698);
nand U2838 (N_2838,In_627,In_724);
and U2839 (N_2839,In_23,In_461);
nor U2840 (N_2840,In_212,In_734);
or U2841 (N_2841,In_562,In_162);
nand U2842 (N_2842,In_122,In_133);
and U2843 (N_2843,In_66,In_1);
nand U2844 (N_2844,In_926,In_426);
nor U2845 (N_2845,In_562,In_925);
xor U2846 (N_2846,In_837,In_453);
nand U2847 (N_2847,In_320,In_394);
and U2848 (N_2848,In_300,In_502);
or U2849 (N_2849,In_945,In_130);
nand U2850 (N_2850,In_203,In_513);
and U2851 (N_2851,In_881,In_936);
or U2852 (N_2852,In_24,In_501);
nand U2853 (N_2853,In_171,In_950);
or U2854 (N_2854,In_926,In_551);
nand U2855 (N_2855,In_408,In_812);
nor U2856 (N_2856,In_977,In_248);
nor U2857 (N_2857,In_634,In_422);
or U2858 (N_2858,In_504,In_475);
nor U2859 (N_2859,In_304,In_619);
and U2860 (N_2860,In_659,In_322);
and U2861 (N_2861,In_108,In_235);
nand U2862 (N_2862,In_274,In_419);
and U2863 (N_2863,In_783,In_752);
or U2864 (N_2864,In_90,In_178);
or U2865 (N_2865,In_785,In_883);
nor U2866 (N_2866,In_298,In_63);
nor U2867 (N_2867,In_38,In_990);
nor U2868 (N_2868,In_959,In_968);
nor U2869 (N_2869,In_190,In_384);
nor U2870 (N_2870,In_980,In_906);
nor U2871 (N_2871,In_626,In_835);
xor U2872 (N_2872,In_429,In_741);
xnor U2873 (N_2873,In_836,In_593);
and U2874 (N_2874,In_687,In_891);
or U2875 (N_2875,In_773,In_330);
nor U2876 (N_2876,In_681,In_90);
xor U2877 (N_2877,In_164,In_223);
and U2878 (N_2878,In_414,In_37);
nor U2879 (N_2879,In_859,In_190);
nor U2880 (N_2880,In_920,In_922);
nor U2881 (N_2881,In_317,In_455);
or U2882 (N_2882,In_785,In_999);
nand U2883 (N_2883,In_30,In_377);
and U2884 (N_2884,In_237,In_529);
or U2885 (N_2885,In_410,In_298);
nand U2886 (N_2886,In_426,In_258);
nor U2887 (N_2887,In_869,In_782);
or U2888 (N_2888,In_446,In_298);
and U2889 (N_2889,In_600,In_310);
nor U2890 (N_2890,In_289,In_172);
nor U2891 (N_2891,In_344,In_283);
nor U2892 (N_2892,In_994,In_964);
and U2893 (N_2893,In_663,In_196);
or U2894 (N_2894,In_187,In_979);
nand U2895 (N_2895,In_257,In_31);
or U2896 (N_2896,In_993,In_7);
nand U2897 (N_2897,In_557,In_700);
or U2898 (N_2898,In_475,In_82);
and U2899 (N_2899,In_43,In_699);
nand U2900 (N_2900,In_325,In_817);
nand U2901 (N_2901,In_80,In_486);
xnor U2902 (N_2902,In_157,In_443);
and U2903 (N_2903,In_600,In_226);
and U2904 (N_2904,In_883,In_744);
nand U2905 (N_2905,In_353,In_285);
nand U2906 (N_2906,In_166,In_721);
nor U2907 (N_2907,In_835,In_870);
and U2908 (N_2908,In_71,In_976);
and U2909 (N_2909,In_723,In_287);
and U2910 (N_2910,In_652,In_714);
nor U2911 (N_2911,In_3,In_652);
nor U2912 (N_2912,In_686,In_39);
and U2913 (N_2913,In_986,In_510);
nor U2914 (N_2914,In_269,In_251);
nor U2915 (N_2915,In_85,In_867);
nand U2916 (N_2916,In_776,In_929);
or U2917 (N_2917,In_820,In_40);
or U2918 (N_2918,In_140,In_941);
xor U2919 (N_2919,In_212,In_90);
nand U2920 (N_2920,In_565,In_896);
and U2921 (N_2921,In_969,In_107);
or U2922 (N_2922,In_747,In_828);
or U2923 (N_2923,In_426,In_785);
nor U2924 (N_2924,In_585,In_327);
or U2925 (N_2925,In_52,In_826);
nand U2926 (N_2926,In_231,In_40);
nand U2927 (N_2927,In_350,In_105);
nor U2928 (N_2928,In_486,In_389);
nor U2929 (N_2929,In_587,In_856);
or U2930 (N_2930,In_123,In_99);
nand U2931 (N_2931,In_322,In_927);
nand U2932 (N_2932,In_315,In_474);
nor U2933 (N_2933,In_615,In_95);
or U2934 (N_2934,In_571,In_80);
nand U2935 (N_2935,In_714,In_344);
nor U2936 (N_2936,In_335,In_759);
nand U2937 (N_2937,In_407,In_830);
and U2938 (N_2938,In_459,In_619);
and U2939 (N_2939,In_54,In_809);
xor U2940 (N_2940,In_317,In_724);
and U2941 (N_2941,In_752,In_724);
and U2942 (N_2942,In_849,In_21);
and U2943 (N_2943,In_52,In_895);
or U2944 (N_2944,In_300,In_154);
nand U2945 (N_2945,In_745,In_857);
and U2946 (N_2946,In_484,In_521);
and U2947 (N_2947,In_852,In_738);
nand U2948 (N_2948,In_93,In_637);
and U2949 (N_2949,In_124,In_597);
nor U2950 (N_2950,In_903,In_169);
nand U2951 (N_2951,In_95,In_466);
nor U2952 (N_2952,In_155,In_487);
and U2953 (N_2953,In_986,In_567);
xor U2954 (N_2954,In_915,In_103);
and U2955 (N_2955,In_304,In_754);
or U2956 (N_2956,In_512,In_440);
nor U2957 (N_2957,In_838,In_323);
or U2958 (N_2958,In_630,In_362);
nor U2959 (N_2959,In_263,In_82);
and U2960 (N_2960,In_600,In_107);
nor U2961 (N_2961,In_532,In_625);
nor U2962 (N_2962,In_318,In_394);
nor U2963 (N_2963,In_298,In_442);
and U2964 (N_2964,In_443,In_531);
nor U2965 (N_2965,In_872,In_133);
nand U2966 (N_2966,In_60,In_749);
nor U2967 (N_2967,In_886,In_803);
or U2968 (N_2968,In_19,In_99);
nand U2969 (N_2969,In_310,In_675);
nor U2970 (N_2970,In_804,In_237);
and U2971 (N_2971,In_286,In_973);
and U2972 (N_2972,In_894,In_946);
nor U2973 (N_2973,In_536,In_946);
nand U2974 (N_2974,In_864,In_205);
nand U2975 (N_2975,In_194,In_314);
and U2976 (N_2976,In_736,In_816);
and U2977 (N_2977,In_369,In_554);
and U2978 (N_2978,In_103,In_173);
nor U2979 (N_2979,In_471,In_958);
nor U2980 (N_2980,In_741,In_956);
and U2981 (N_2981,In_650,In_764);
and U2982 (N_2982,In_75,In_861);
and U2983 (N_2983,In_671,In_328);
and U2984 (N_2984,In_346,In_373);
or U2985 (N_2985,In_337,In_881);
or U2986 (N_2986,In_100,In_64);
nor U2987 (N_2987,In_689,In_821);
nor U2988 (N_2988,In_884,In_362);
and U2989 (N_2989,In_5,In_242);
and U2990 (N_2990,In_432,In_953);
nand U2991 (N_2991,In_761,In_393);
or U2992 (N_2992,In_230,In_930);
and U2993 (N_2993,In_645,In_857);
nor U2994 (N_2994,In_425,In_813);
nand U2995 (N_2995,In_108,In_712);
and U2996 (N_2996,In_796,In_28);
or U2997 (N_2997,In_818,In_207);
nand U2998 (N_2998,In_508,In_506);
nor U2999 (N_2999,In_663,In_351);
or U3000 (N_3000,In_312,In_547);
or U3001 (N_3001,In_374,In_937);
nand U3002 (N_3002,In_664,In_317);
nor U3003 (N_3003,In_469,In_831);
xor U3004 (N_3004,In_345,In_975);
nor U3005 (N_3005,In_787,In_55);
and U3006 (N_3006,In_566,In_556);
or U3007 (N_3007,In_995,In_810);
xnor U3008 (N_3008,In_501,In_463);
nand U3009 (N_3009,In_402,In_873);
or U3010 (N_3010,In_833,In_666);
nor U3011 (N_3011,In_290,In_60);
and U3012 (N_3012,In_47,In_474);
nor U3013 (N_3013,In_403,In_303);
and U3014 (N_3014,In_119,In_100);
nand U3015 (N_3015,In_576,In_734);
or U3016 (N_3016,In_999,In_230);
and U3017 (N_3017,In_283,In_937);
xnor U3018 (N_3018,In_152,In_530);
nor U3019 (N_3019,In_635,In_850);
and U3020 (N_3020,In_171,In_846);
and U3021 (N_3021,In_920,In_35);
xor U3022 (N_3022,In_15,In_23);
nor U3023 (N_3023,In_844,In_53);
nand U3024 (N_3024,In_432,In_189);
and U3025 (N_3025,In_234,In_409);
or U3026 (N_3026,In_242,In_762);
nor U3027 (N_3027,In_608,In_298);
or U3028 (N_3028,In_116,In_4);
xor U3029 (N_3029,In_106,In_841);
or U3030 (N_3030,In_198,In_567);
and U3031 (N_3031,In_780,In_391);
nor U3032 (N_3032,In_698,In_545);
nor U3033 (N_3033,In_734,In_501);
or U3034 (N_3034,In_585,In_533);
nand U3035 (N_3035,In_116,In_919);
or U3036 (N_3036,In_46,In_657);
and U3037 (N_3037,In_763,In_147);
or U3038 (N_3038,In_988,In_456);
or U3039 (N_3039,In_531,In_904);
or U3040 (N_3040,In_86,In_884);
xnor U3041 (N_3041,In_700,In_686);
nor U3042 (N_3042,In_988,In_838);
nor U3043 (N_3043,In_31,In_682);
nor U3044 (N_3044,In_665,In_565);
or U3045 (N_3045,In_783,In_439);
or U3046 (N_3046,In_229,In_103);
or U3047 (N_3047,In_815,In_430);
and U3048 (N_3048,In_414,In_239);
or U3049 (N_3049,In_194,In_54);
or U3050 (N_3050,In_342,In_186);
nor U3051 (N_3051,In_223,In_77);
or U3052 (N_3052,In_822,In_934);
and U3053 (N_3053,In_439,In_72);
and U3054 (N_3054,In_42,In_253);
and U3055 (N_3055,In_511,In_336);
xnor U3056 (N_3056,In_354,In_133);
nand U3057 (N_3057,In_380,In_699);
or U3058 (N_3058,In_451,In_505);
and U3059 (N_3059,In_198,In_840);
nand U3060 (N_3060,In_258,In_845);
nand U3061 (N_3061,In_302,In_163);
nand U3062 (N_3062,In_645,In_633);
and U3063 (N_3063,In_99,In_396);
nor U3064 (N_3064,In_212,In_286);
or U3065 (N_3065,In_770,In_865);
and U3066 (N_3066,In_960,In_310);
nand U3067 (N_3067,In_483,In_195);
and U3068 (N_3068,In_806,In_66);
nor U3069 (N_3069,In_659,In_210);
and U3070 (N_3070,In_252,In_446);
nor U3071 (N_3071,In_268,In_836);
and U3072 (N_3072,In_222,In_96);
nand U3073 (N_3073,In_564,In_193);
nor U3074 (N_3074,In_265,In_927);
nand U3075 (N_3075,In_83,In_529);
or U3076 (N_3076,In_684,In_106);
nand U3077 (N_3077,In_864,In_348);
or U3078 (N_3078,In_544,In_418);
or U3079 (N_3079,In_547,In_847);
nor U3080 (N_3080,In_900,In_930);
nor U3081 (N_3081,In_59,In_940);
nand U3082 (N_3082,In_342,In_77);
or U3083 (N_3083,In_765,In_123);
nand U3084 (N_3084,In_978,In_782);
nor U3085 (N_3085,In_210,In_862);
or U3086 (N_3086,In_515,In_841);
nor U3087 (N_3087,In_408,In_764);
or U3088 (N_3088,In_566,In_69);
and U3089 (N_3089,In_160,In_279);
nor U3090 (N_3090,In_97,In_921);
or U3091 (N_3091,In_311,In_86);
nand U3092 (N_3092,In_196,In_78);
or U3093 (N_3093,In_652,In_193);
or U3094 (N_3094,In_140,In_744);
or U3095 (N_3095,In_323,In_552);
or U3096 (N_3096,In_300,In_174);
nand U3097 (N_3097,In_721,In_906);
nor U3098 (N_3098,In_681,In_272);
or U3099 (N_3099,In_293,In_833);
nand U3100 (N_3100,In_723,In_696);
nand U3101 (N_3101,In_845,In_352);
and U3102 (N_3102,In_846,In_137);
and U3103 (N_3103,In_359,In_918);
nand U3104 (N_3104,In_627,In_684);
and U3105 (N_3105,In_721,In_266);
and U3106 (N_3106,In_277,In_858);
nor U3107 (N_3107,In_140,In_714);
or U3108 (N_3108,In_275,In_230);
or U3109 (N_3109,In_339,In_195);
xnor U3110 (N_3110,In_412,In_383);
or U3111 (N_3111,In_12,In_29);
nand U3112 (N_3112,In_272,In_244);
and U3113 (N_3113,In_584,In_201);
nor U3114 (N_3114,In_730,In_743);
nor U3115 (N_3115,In_944,In_467);
and U3116 (N_3116,In_554,In_986);
nor U3117 (N_3117,In_671,In_503);
xnor U3118 (N_3118,In_584,In_392);
nand U3119 (N_3119,In_237,In_614);
or U3120 (N_3120,In_182,In_684);
nand U3121 (N_3121,In_601,In_791);
and U3122 (N_3122,In_669,In_463);
nand U3123 (N_3123,In_969,In_947);
nand U3124 (N_3124,In_204,In_455);
or U3125 (N_3125,In_841,In_374);
and U3126 (N_3126,In_335,In_43);
nor U3127 (N_3127,In_685,In_514);
nor U3128 (N_3128,In_955,In_930);
and U3129 (N_3129,In_619,In_598);
nand U3130 (N_3130,In_170,In_186);
and U3131 (N_3131,In_289,In_628);
nand U3132 (N_3132,In_436,In_307);
or U3133 (N_3133,In_446,In_109);
xor U3134 (N_3134,In_670,In_56);
and U3135 (N_3135,In_995,In_611);
nor U3136 (N_3136,In_308,In_487);
or U3137 (N_3137,In_654,In_150);
or U3138 (N_3138,In_526,In_210);
nor U3139 (N_3139,In_465,In_75);
and U3140 (N_3140,In_32,In_741);
and U3141 (N_3141,In_858,In_820);
nor U3142 (N_3142,In_965,In_858);
or U3143 (N_3143,In_313,In_133);
and U3144 (N_3144,In_543,In_689);
and U3145 (N_3145,In_585,In_37);
nand U3146 (N_3146,In_802,In_470);
and U3147 (N_3147,In_885,In_60);
and U3148 (N_3148,In_872,In_46);
and U3149 (N_3149,In_575,In_894);
nand U3150 (N_3150,In_1,In_576);
nand U3151 (N_3151,In_315,In_65);
or U3152 (N_3152,In_788,In_275);
or U3153 (N_3153,In_384,In_341);
nand U3154 (N_3154,In_117,In_996);
and U3155 (N_3155,In_718,In_404);
nor U3156 (N_3156,In_924,In_995);
nand U3157 (N_3157,In_958,In_474);
and U3158 (N_3158,In_731,In_714);
nor U3159 (N_3159,In_268,In_955);
nand U3160 (N_3160,In_47,In_57);
or U3161 (N_3161,In_22,In_742);
or U3162 (N_3162,In_416,In_148);
nor U3163 (N_3163,In_97,In_932);
and U3164 (N_3164,In_618,In_350);
nor U3165 (N_3165,In_913,In_844);
nand U3166 (N_3166,In_213,In_867);
or U3167 (N_3167,In_679,In_788);
or U3168 (N_3168,In_359,In_709);
nand U3169 (N_3169,In_464,In_622);
nand U3170 (N_3170,In_932,In_818);
and U3171 (N_3171,In_842,In_578);
nor U3172 (N_3172,In_587,In_302);
or U3173 (N_3173,In_795,In_434);
or U3174 (N_3174,In_987,In_498);
or U3175 (N_3175,In_718,In_634);
nand U3176 (N_3176,In_487,In_686);
xor U3177 (N_3177,In_376,In_456);
and U3178 (N_3178,In_767,In_441);
or U3179 (N_3179,In_939,In_326);
nor U3180 (N_3180,In_69,In_969);
xnor U3181 (N_3181,In_46,In_518);
nor U3182 (N_3182,In_140,In_151);
and U3183 (N_3183,In_64,In_934);
nand U3184 (N_3184,In_453,In_506);
nand U3185 (N_3185,In_854,In_922);
or U3186 (N_3186,In_895,In_771);
and U3187 (N_3187,In_252,In_800);
and U3188 (N_3188,In_779,In_246);
nand U3189 (N_3189,In_442,In_230);
or U3190 (N_3190,In_347,In_747);
nand U3191 (N_3191,In_453,In_735);
nor U3192 (N_3192,In_43,In_199);
nand U3193 (N_3193,In_422,In_943);
and U3194 (N_3194,In_659,In_235);
nor U3195 (N_3195,In_680,In_323);
nand U3196 (N_3196,In_412,In_688);
nand U3197 (N_3197,In_963,In_524);
nand U3198 (N_3198,In_64,In_858);
or U3199 (N_3199,In_571,In_39);
and U3200 (N_3200,In_467,In_167);
and U3201 (N_3201,In_405,In_100);
and U3202 (N_3202,In_180,In_5);
nor U3203 (N_3203,In_110,In_427);
or U3204 (N_3204,In_480,In_979);
or U3205 (N_3205,In_402,In_567);
nor U3206 (N_3206,In_1,In_735);
and U3207 (N_3207,In_977,In_222);
or U3208 (N_3208,In_696,In_724);
or U3209 (N_3209,In_427,In_862);
nor U3210 (N_3210,In_885,In_505);
and U3211 (N_3211,In_48,In_834);
nand U3212 (N_3212,In_108,In_973);
or U3213 (N_3213,In_544,In_384);
or U3214 (N_3214,In_969,In_754);
and U3215 (N_3215,In_965,In_785);
and U3216 (N_3216,In_755,In_611);
nand U3217 (N_3217,In_269,In_673);
nor U3218 (N_3218,In_158,In_102);
and U3219 (N_3219,In_695,In_956);
nand U3220 (N_3220,In_506,In_744);
and U3221 (N_3221,In_299,In_968);
nand U3222 (N_3222,In_510,In_617);
nor U3223 (N_3223,In_552,In_357);
or U3224 (N_3224,In_737,In_444);
and U3225 (N_3225,In_891,In_530);
and U3226 (N_3226,In_858,In_648);
or U3227 (N_3227,In_266,In_497);
and U3228 (N_3228,In_141,In_761);
nor U3229 (N_3229,In_21,In_840);
xnor U3230 (N_3230,In_101,In_662);
or U3231 (N_3231,In_808,In_780);
nand U3232 (N_3232,In_309,In_764);
and U3233 (N_3233,In_606,In_94);
and U3234 (N_3234,In_554,In_546);
and U3235 (N_3235,In_379,In_335);
nor U3236 (N_3236,In_401,In_921);
nor U3237 (N_3237,In_808,In_971);
nand U3238 (N_3238,In_740,In_838);
or U3239 (N_3239,In_896,In_852);
or U3240 (N_3240,In_602,In_802);
nor U3241 (N_3241,In_752,In_456);
nor U3242 (N_3242,In_788,In_948);
nand U3243 (N_3243,In_566,In_233);
or U3244 (N_3244,In_794,In_520);
or U3245 (N_3245,In_333,In_423);
or U3246 (N_3246,In_93,In_512);
nand U3247 (N_3247,In_783,In_998);
and U3248 (N_3248,In_69,In_176);
and U3249 (N_3249,In_777,In_131);
and U3250 (N_3250,In_467,In_766);
or U3251 (N_3251,In_90,In_935);
nor U3252 (N_3252,In_513,In_904);
nand U3253 (N_3253,In_880,In_696);
nand U3254 (N_3254,In_262,In_233);
nand U3255 (N_3255,In_926,In_98);
xnor U3256 (N_3256,In_725,In_328);
and U3257 (N_3257,In_134,In_892);
nand U3258 (N_3258,In_613,In_753);
nor U3259 (N_3259,In_877,In_600);
nand U3260 (N_3260,In_429,In_122);
nand U3261 (N_3261,In_730,In_467);
or U3262 (N_3262,In_235,In_489);
and U3263 (N_3263,In_475,In_940);
nand U3264 (N_3264,In_413,In_53);
or U3265 (N_3265,In_395,In_499);
nor U3266 (N_3266,In_269,In_522);
or U3267 (N_3267,In_50,In_298);
or U3268 (N_3268,In_632,In_51);
and U3269 (N_3269,In_471,In_659);
nor U3270 (N_3270,In_759,In_637);
and U3271 (N_3271,In_987,In_681);
or U3272 (N_3272,In_411,In_900);
and U3273 (N_3273,In_369,In_127);
nand U3274 (N_3274,In_364,In_125);
nor U3275 (N_3275,In_865,In_67);
nand U3276 (N_3276,In_935,In_607);
nor U3277 (N_3277,In_565,In_325);
or U3278 (N_3278,In_137,In_43);
nand U3279 (N_3279,In_73,In_341);
nor U3280 (N_3280,In_279,In_61);
and U3281 (N_3281,In_873,In_470);
nand U3282 (N_3282,In_192,In_75);
nand U3283 (N_3283,In_960,In_560);
or U3284 (N_3284,In_206,In_170);
and U3285 (N_3285,In_415,In_523);
or U3286 (N_3286,In_622,In_700);
and U3287 (N_3287,In_817,In_262);
and U3288 (N_3288,In_206,In_193);
or U3289 (N_3289,In_540,In_388);
nor U3290 (N_3290,In_147,In_462);
and U3291 (N_3291,In_698,In_164);
and U3292 (N_3292,In_623,In_738);
or U3293 (N_3293,In_625,In_849);
or U3294 (N_3294,In_982,In_285);
nand U3295 (N_3295,In_798,In_952);
nand U3296 (N_3296,In_439,In_908);
and U3297 (N_3297,In_340,In_520);
or U3298 (N_3298,In_1,In_365);
and U3299 (N_3299,In_801,In_530);
and U3300 (N_3300,In_895,In_638);
and U3301 (N_3301,In_384,In_652);
or U3302 (N_3302,In_531,In_401);
nand U3303 (N_3303,In_230,In_538);
or U3304 (N_3304,In_656,In_441);
or U3305 (N_3305,In_996,In_17);
nor U3306 (N_3306,In_878,In_304);
nand U3307 (N_3307,In_382,In_272);
nor U3308 (N_3308,In_741,In_84);
and U3309 (N_3309,In_804,In_459);
nand U3310 (N_3310,In_63,In_490);
nand U3311 (N_3311,In_487,In_133);
nor U3312 (N_3312,In_455,In_18);
nand U3313 (N_3313,In_352,In_930);
nand U3314 (N_3314,In_635,In_511);
nor U3315 (N_3315,In_92,In_831);
or U3316 (N_3316,In_606,In_286);
nand U3317 (N_3317,In_180,In_110);
nand U3318 (N_3318,In_948,In_185);
or U3319 (N_3319,In_568,In_953);
nand U3320 (N_3320,In_95,In_705);
xor U3321 (N_3321,In_893,In_163);
or U3322 (N_3322,In_242,In_877);
and U3323 (N_3323,In_665,In_832);
nand U3324 (N_3324,In_288,In_190);
xnor U3325 (N_3325,In_443,In_920);
nand U3326 (N_3326,In_386,In_218);
nor U3327 (N_3327,In_632,In_826);
or U3328 (N_3328,In_730,In_734);
nor U3329 (N_3329,In_134,In_783);
nor U3330 (N_3330,In_335,In_388);
or U3331 (N_3331,In_454,In_333);
or U3332 (N_3332,In_793,In_223);
and U3333 (N_3333,In_579,In_725);
or U3334 (N_3334,In_337,In_389);
and U3335 (N_3335,In_920,In_787);
nand U3336 (N_3336,In_287,In_16);
nor U3337 (N_3337,In_377,In_399);
and U3338 (N_3338,In_965,In_137);
and U3339 (N_3339,In_825,In_965);
or U3340 (N_3340,In_473,In_806);
nor U3341 (N_3341,In_800,In_495);
nand U3342 (N_3342,In_295,In_44);
and U3343 (N_3343,In_307,In_948);
nand U3344 (N_3344,In_410,In_591);
nor U3345 (N_3345,In_654,In_633);
nand U3346 (N_3346,In_707,In_220);
nand U3347 (N_3347,In_47,In_164);
nor U3348 (N_3348,In_149,In_51);
and U3349 (N_3349,In_307,In_310);
nand U3350 (N_3350,In_799,In_249);
or U3351 (N_3351,In_271,In_53);
xor U3352 (N_3352,In_859,In_494);
nand U3353 (N_3353,In_694,In_229);
xor U3354 (N_3354,In_324,In_670);
or U3355 (N_3355,In_843,In_710);
or U3356 (N_3356,In_970,In_767);
nand U3357 (N_3357,In_265,In_192);
or U3358 (N_3358,In_570,In_753);
nor U3359 (N_3359,In_626,In_642);
nor U3360 (N_3360,In_933,In_858);
nand U3361 (N_3361,In_846,In_686);
nor U3362 (N_3362,In_817,In_592);
or U3363 (N_3363,In_151,In_738);
and U3364 (N_3364,In_895,In_710);
or U3365 (N_3365,In_94,In_709);
and U3366 (N_3366,In_121,In_647);
nor U3367 (N_3367,In_70,In_276);
or U3368 (N_3368,In_713,In_898);
nor U3369 (N_3369,In_48,In_798);
nor U3370 (N_3370,In_754,In_182);
nand U3371 (N_3371,In_229,In_365);
and U3372 (N_3372,In_807,In_257);
nor U3373 (N_3373,In_81,In_567);
nand U3374 (N_3374,In_158,In_994);
nor U3375 (N_3375,In_47,In_672);
or U3376 (N_3376,In_464,In_889);
or U3377 (N_3377,In_809,In_815);
nor U3378 (N_3378,In_97,In_713);
or U3379 (N_3379,In_724,In_198);
nor U3380 (N_3380,In_60,In_924);
nand U3381 (N_3381,In_207,In_255);
nand U3382 (N_3382,In_826,In_853);
or U3383 (N_3383,In_784,In_633);
or U3384 (N_3384,In_273,In_916);
nand U3385 (N_3385,In_970,In_97);
or U3386 (N_3386,In_768,In_407);
nor U3387 (N_3387,In_332,In_14);
nand U3388 (N_3388,In_975,In_626);
or U3389 (N_3389,In_623,In_360);
nand U3390 (N_3390,In_277,In_397);
nand U3391 (N_3391,In_409,In_644);
nor U3392 (N_3392,In_13,In_841);
and U3393 (N_3393,In_237,In_907);
nand U3394 (N_3394,In_867,In_386);
nor U3395 (N_3395,In_877,In_450);
nand U3396 (N_3396,In_343,In_973);
and U3397 (N_3397,In_3,In_685);
nand U3398 (N_3398,In_694,In_110);
and U3399 (N_3399,In_75,In_446);
or U3400 (N_3400,In_2,In_891);
nor U3401 (N_3401,In_195,In_385);
nor U3402 (N_3402,In_939,In_466);
and U3403 (N_3403,In_158,In_349);
nor U3404 (N_3404,In_409,In_296);
nand U3405 (N_3405,In_130,In_56);
or U3406 (N_3406,In_266,In_978);
nand U3407 (N_3407,In_744,In_623);
nor U3408 (N_3408,In_681,In_145);
nor U3409 (N_3409,In_293,In_158);
and U3410 (N_3410,In_570,In_442);
or U3411 (N_3411,In_284,In_421);
nor U3412 (N_3412,In_64,In_486);
nand U3413 (N_3413,In_338,In_568);
and U3414 (N_3414,In_860,In_802);
and U3415 (N_3415,In_119,In_826);
nand U3416 (N_3416,In_548,In_698);
or U3417 (N_3417,In_264,In_379);
nand U3418 (N_3418,In_902,In_556);
nand U3419 (N_3419,In_324,In_70);
and U3420 (N_3420,In_389,In_101);
nor U3421 (N_3421,In_797,In_921);
and U3422 (N_3422,In_836,In_715);
nand U3423 (N_3423,In_962,In_130);
nor U3424 (N_3424,In_851,In_785);
nand U3425 (N_3425,In_523,In_542);
and U3426 (N_3426,In_191,In_33);
and U3427 (N_3427,In_347,In_866);
nor U3428 (N_3428,In_282,In_104);
and U3429 (N_3429,In_838,In_587);
or U3430 (N_3430,In_247,In_527);
or U3431 (N_3431,In_689,In_973);
nor U3432 (N_3432,In_986,In_991);
or U3433 (N_3433,In_826,In_223);
and U3434 (N_3434,In_104,In_948);
or U3435 (N_3435,In_203,In_393);
and U3436 (N_3436,In_538,In_732);
or U3437 (N_3437,In_785,In_963);
and U3438 (N_3438,In_689,In_411);
or U3439 (N_3439,In_226,In_908);
nor U3440 (N_3440,In_911,In_319);
nor U3441 (N_3441,In_763,In_404);
and U3442 (N_3442,In_420,In_413);
xnor U3443 (N_3443,In_907,In_257);
xnor U3444 (N_3444,In_669,In_889);
nand U3445 (N_3445,In_947,In_980);
and U3446 (N_3446,In_736,In_627);
nor U3447 (N_3447,In_424,In_32);
and U3448 (N_3448,In_364,In_4);
nor U3449 (N_3449,In_897,In_947);
xor U3450 (N_3450,In_153,In_515);
or U3451 (N_3451,In_860,In_620);
nand U3452 (N_3452,In_788,In_926);
nor U3453 (N_3453,In_795,In_870);
or U3454 (N_3454,In_104,In_158);
nor U3455 (N_3455,In_325,In_581);
and U3456 (N_3456,In_997,In_469);
and U3457 (N_3457,In_323,In_165);
and U3458 (N_3458,In_392,In_782);
nand U3459 (N_3459,In_316,In_244);
and U3460 (N_3460,In_500,In_69);
or U3461 (N_3461,In_209,In_342);
nor U3462 (N_3462,In_184,In_75);
or U3463 (N_3463,In_476,In_624);
and U3464 (N_3464,In_817,In_784);
nor U3465 (N_3465,In_52,In_945);
or U3466 (N_3466,In_641,In_958);
or U3467 (N_3467,In_750,In_914);
or U3468 (N_3468,In_445,In_61);
xnor U3469 (N_3469,In_616,In_694);
xnor U3470 (N_3470,In_612,In_675);
nand U3471 (N_3471,In_6,In_662);
or U3472 (N_3472,In_223,In_690);
and U3473 (N_3473,In_74,In_300);
nor U3474 (N_3474,In_335,In_232);
or U3475 (N_3475,In_85,In_134);
nor U3476 (N_3476,In_293,In_322);
nor U3477 (N_3477,In_815,In_918);
and U3478 (N_3478,In_227,In_492);
and U3479 (N_3479,In_362,In_926);
nor U3480 (N_3480,In_51,In_510);
or U3481 (N_3481,In_695,In_571);
nand U3482 (N_3482,In_595,In_829);
nor U3483 (N_3483,In_652,In_378);
and U3484 (N_3484,In_737,In_642);
or U3485 (N_3485,In_510,In_680);
and U3486 (N_3486,In_831,In_569);
and U3487 (N_3487,In_383,In_471);
nor U3488 (N_3488,In_80,In_928);
nand U3489 (N_3489,In_201,In_891);
nor U3490 (N_3490,In_268,In_205);
and U3491 (N_3491,In_141,In_227);
nand U3492 (N_3492,In_796,In_766);
or U3493 (N_3493,In_547,In_735);
and U3494 (N_3494,In_734,In_309);
or U3495 (N_3495,In_648,In_464);
and U3496 (N_3496,In_822,In_20);
nand U3497 (N_3497,In_821,In_450);
nor U3498 (N_3498,In_853,In_931);
nand U3499 (N_3499,In_459,In_927);
nand U3500 (N_3500,In_595,In_892);
or U3501 (N_3501,In_61,In_480);
nand U3502 (N_3502,In_462,In_437);
nor U3503 (N_3503,In_603,In_397);
or U3504 (N_3504,In_750,In_867);
and U3505 (N_3505,In_886,In_976);
xor U3506 (N_3506,In_553,In_498);
nand U3507 (N_3507,In_539,In_792);
or U3508 (N_3508,In_560,In_669);
and U3509 (N_3509,In_740,In_109);
and U3510 (N_3510,In_878,In_151);
nand U3511 (N_3511,In_690,In_338);
nand U3512 (N_3512,In_377,In_39);
nand U3513 (N_3513,In_495,In_265);
or U3514 (N_3514,In_940,In_77);
and U3515 (N_3515,In_789,In_912);
or U3516 (N_3516,In_650,In_642);
nand U3517 (N_3517,In_231,In_579);
xor U3518 (N_3518,In_435,In_475);
and U3519 (N_3519,In_298,In_480);
nor U3520 (N_3520,In_157,In_504);
nand U3521 (N_3521,In_237,In_246);
and U3522 (N_3522,In_114,In_783);
and U3523 (N_3523,In_207,In_142);
nor U3524 (N_3524,In_622,In_207);
nand U3525 (N_3525,In_385,In_350);
and U3526 (N_3526,In_5,In_814);
nor U3527 (N_3527,In_528,In_137);
nor U3528 (N_3528,In_327,In_454);
nand U3529 (N_3529,In_868,In_988);
nand U3530 (N_3530,In_39,In_56);
and U3531 (N_3531,In_937,In_727);
nand U3532 (N_3532,In_528,In_379);
nor U3533 (N_3533,In_633,In_82);
and U3534 (N_3534,In_389,In_798);
or U3535 (N_3535,In_188,In_163);
and U3536 (N_3536,In_666,In_302);
and U3537 (N_3537,In_753,In_369);
and U3538 (N_3538,In_23,In_632);
or U3539 (N_3539,In_887,In_147);
nor U3540 (N_3540,In_915,In_68);
or U3541 (N_3541,In_727,In_248);
and U3542 (N_3542,In_349,In_88);
xnor U3543 (N_3543,In_427,In_403);
or U3544 (N_3544,In_529,In_144);
and U3545 (N_3545,In_966,In_382);
xnor U3546 (N_3546,In_329,In_65);
nor U3547 (N_3547,In_326,In_413);
nor U3548 (N_3548,In_952,In_372);
xor U3549 (N_3549,In_800,In_773);
nor U3550 (N_3550,In_80,In_339);
or U3551 (N_3551,In_729,In_753);
nand U3552 (N_3552,In_72,In_125);
nor U3553 (N_3553,In_664,In_256);
or U3554 (N_3554,In_907,In_121);
nor U3555 (N_3555,In_831,In_137);
nand U3556 (N_3556,In_188,In_271);
and U3557 (N_3557,In_423,In_859);
nor U3558 (N_3558,In_671,In_601);
nand U3559 (N_3559,In_642,In_162);
nand U3560 (N_3560,In_620,In_688);
nor U3561 (N_3561,In_788,In_762);
nor U3562 (N_3562,In_799,In_850);
nor U3563 (N_3563,In_932,In_43);
nor U3564 (N_3564,In_124,In_711);
and U3565 (N_3565,In_408,In_469);
and U3566 (N_3566,In_759,In_202);
and U3567 (N_3567,In_536,In_767);
and U3568 (N_3568,In_333,In_555);
nand U3569 (N_3569,In_32,In_848);
or U3570 (N_3570,In_294,In_164);
and U3571 (N_3571,In_126,In_701);
or U3572 (N_3572,In_645,In_931);
nor U3573 (N_3573,In_50,In_527);
or U3574 (N_3574,In_567,In_625);
and U3575 (N_3575,In_717,In_832);
or U3576 (N_3576,In_991,In_712);
and U3577 (N_3577,In_607,In_990);
xnor U3578 (N_3578,In_532,In_426);
nand U3579 (N_3579,In_826,In_568);
nor U3580 (N_3580,In_880,In_257);
or U3581 (N_3581,In_949,In_827);
nor U3582 (N_3582,In_510,In_100);
nand U3583 (N_3583,In_184,In_866);
nor U3584 (N_3584,In_487,In_632);
nand U3585 (N_3585,In_63,In_97);
and U3586 (N_3586,In_591,In_766);
nand U3587 (N_3587,In_590,In_102);
xnor U3588 (N_3588,In_943,In_241);
and U3589 (N_3589,In_57,In_835);
and U3590 (N_3590,In_280,In_668);
nor U3591 (N_3591,In_870,In_846);
nor U3592 (N_3592,In_713,In_378);
nor U3593 (N_3593,In_754,In_229);
and U3594 (N_3594,In_769,In_929);
and U3595 (N_3595,In_106,In_600);
nor U3596 (N_3596,In_38,In_871);
or U3597 (N_3597,In_162,In_797);
or U3598 (N_3598,In_147,In_871);
nor U3599 (N_3599,In_85,In_181);
nor U3600 (N_3600,In_58,In_515);
nor U3601 (N_3601,In_691,In_867);
nand U3602 (N_3602,In_364,In_746);
or U3603 (N_3603,In_796,In_54);
nor U3604 (N_3604,In_387,In_99);
and U3605 (N_3605,In_393,In_723);
and U3606 (N_3606,In_596,In_304);
and U3607 (N_3607,In_504,In_965);
and U3608 (N_3608,In_279,In_474);
xnor U3609 (N_3609,In_803,In_171);
and U3610 (N_3610,In_5,In_476);
and U3611 (N_3611,In_8,In_16);
and U3612 (N_3612,In_846,In_720);
and U3613 (N_3613,In_544,In_774);
or U3614 (N_3614,In_891,In_763);
nor U3615 (N_3615,In_642,In_513);
nor U3616 (N_3616,In_225,In_153);
or U3617 (N_3617,In_590,In_412);
and U3618 (N_3618,In_303,In_618);
nand U3619 (N_3619,In_540,In_549);
and U3620 (N_3620,In_254,In_171);
and U3621 (N_3621,In_652,In_7);
and U3622 (N_3622,In_499,In_912);
nand U3623 (N_3623,In_886,In_937);
nand U3624 (N_3624,In_792,In_847);
nor U3625 (N_3625,In_112,In_826);
or U3626 (N_3626,In_393,In_279);
nand U3627 (N_3627,In_66,In_903);
and U3628 (N_3628,In_487,In_433);
nor U3629 (N_3629,In_679,In_561);
nand U3630 (N_3630,In_116,In_780);
and U3631 (N_3631,In_208,In_536);
nor U3632 (N_3632,In_918,In_648);
and U3633 (N_3633,In_191,In_771);
nand U3634 (N_3634,In_422,In_300);
and U3635 (N_3635,In_102,In_215);
nor U3636 (N_3636,In_893,In_331);
nand U3637 (N_3637,In_281,In_506);
nor U3638 (N_3638,In_524,In_387);
and U3639 (N_3639,In_135,In_821);
or U3640 (N_3640,In_156,In_368);
or U3641 (N_3641,In_321,In_615);
or U3642 (N_3642,In_165,In_292);
nand U3643 (N_3643,In_935,In_655);
nand U3644 (N_3644,In_303,In_907);
nand U3645 (N_3645,In_297,In_431);
and U3646 (N_3646,In_717,In_718);
nor U3647 (N_3647,In_634,In_472);
or U3648 (N_3648,In_771,In_626);
or U3649 (N_3649,In_434,In_114);
or U3650 (N_3650,In_951,In_534);
nor U3651 (N_3651,In_594,In_888);
nand U3652 (N_3652,In_446,In_563);
or U3653 (N_3653,In_860,In_746);
or U3654 (N_3654,In_373,In_94);
or U3655 (N_3655,In_390,In_771);
and U3656 (N_3656,In_21,In_305);
nor U3657 (N_3657,In_385,In_270);
nand U3658 (N_3658,In_633,In_252);
nor U3659 (N_3659,In_945,In_66);
or U3660 (N_3660,In_943,In_814);
nor U3661 (N_3661,In_569,In_690);
nand U3662 (N_3662,In_17,In_850);
or U3663 (N_3663,In_128,In_687);
nor U3664 (N_3664,In_12,In_703);
and U3665 (N_3665,In_641,In_758);
nand U3666 (N_3666,In_187,In_628);
nand U3667 (N_3667,In_964,In_121);
nor U3668 (N_3668,In_6,In_888);
nand U3669 (N_3669,In_162,In_134);
nor U3670 (N_3670,In_669,In_167);
and U3671 (N_3671,In_679,In_785);
or U3672 (N_3672,In_755,In_313);
or U3673 (N_3673,In_171,In_713);
nor U3674 (N_3674,In_882,In_869);
xor U3675 (N_3675,In_531,In_286);
nor U3676 (N_3676,In_132,In_18);
nor U3677 (N_3677,In_957,In_132);
and U3678 (N_3678,In_114,In_671);
nor U3679 (N_3679,In_77,In_351);
and U3680 (N_3680,In_140,In_972);
xnor U3681 (N_3681,In_652,In_782);
xnor U3682 (N_3682,In_511,In_125);
nand U3683 (N_3683,In_919,In_82);
or U3684 (N_3684,In_960,In_140);
and U3685 (N_3685,In_278,In_899);
nor U3686 (N_3686,In_349,In_696);
and U3687 (N_3687,In_800,In_798);
nand U3688 (N_3688,In_675,In_539);
nand U3689 (N_3689,In_254,In_386);
and U3690 (N_3690,In_482,In_460);
or U3691 (N_3691,In_737,In_718);
nand U3692 (N_3692,In_495,In_659);
nor U3693 (N_3693,In_674,In_899);
xnor U3694 (N_3694,In_243,In_75);
nor U3695 (N_3695,In_434,In_90);
nor U3696 (N_3696,In_462,In_530);
and U3697 (N_3697,In_660,In_473);
nand U3698 (N_3698,In_721,In_703);
nand U3699 (N_3699,In_25,In_498);
nor U3700 (N_3700,In_512,In_511);
nand U3701 (N_3701,In_168,In_713);
xnor U3702 (N_3702,In_856,In_454);
nand U3703 (N_3703,In_126,In_834);
nor U3704 (N_3704,In_466,In_179);
and U3705 (N_3705,In_603,In_326);
xor U3706 (N_3706,In_520,In_666);
nand U3707 (N_3707,In_66,In_577);
and U3708 (N_3708,In_389,In_452);
and U3709 (N_3709,In_800,In_280);
nand U3710 (N_3710,In_794,In_117);
nand U3711 (N_3711,In_161,In_319);
xnor U3712 (N_3712,In_24,In_346);
nand U3713 (N_3713,In_266,In_810);
nand U3714 (N_3714,In_232,In_927);
or U3715 (N_3715,In_857,In_752);
and U3716 (N_3716,In_504,In_286);
nor U3717 (N_3717,In_144,In_589);
nand U3718 (N_3718,In_1,In_33);
nand U3719 (N_3719,In_7,In_66);
nand U3720 (N_3720,In_729,In_972);
or U3721 (N_3721,In_312,In_863);
nor U3722 (N_3722,In_707,In_756);
and U3723 (N_3723,In_420,In_490);
or U3724 (N_3724,In_223,In_626);
nand U3725 (N_3725,In_158,In_775);
and U3726 (N_3726,In_952,In_419);
nand U3727 (N_3727,In_270,In_411);
nor U3728 (N_3728,In_687,In_60);
or U3729 (N_3729,In_189,In_480);
nor U3730 (N_3730,In_545,In_127);
xnor U3731 (N_3731,In_375,In_777);
nand U3732 (N_3732,In_733,In_587);
or U3733 (N_3733,In_108,In_64);
nor U3734 (N_3734,In_392,In_661);
nand U3735 (N_3735,In_26,In_450);
nand U3736 (N_3736,In_583,In_888);
nand U3737 (N_3737,In_201,In_758);
or U3738 (N_3738,In_371,In_125);
nand U3739 (N_3739,In_809,In_18);
nor U3740 (N_3740,In_902,In_594);
nor U3741 (N_3741,In_92,In_536);
and U3742 (N_3742,In_252,In_723);
nor U3743 (N_3743,In_210,In_519);
and U3744 (N_3744,In_809,In_904);
nor U3745 (N_3745,In_839,In_417);
and U3746 (N_3746,In_724,In_394);
or U3747 (N_3747,In_659,In_282);
nand U3748 (N_3748,In_232,In_548);
nor U3749 (N_3749,In_804,In_951);
nand U3750 (N_3750,In_167,In_898);
nor U3751 (N_3751,In_570,In_940);
and U3752 (N_3752,In_40,In_218);
xnor U3753 (N_3753,In_291,In_549);
nand U3754 (N_3754,In_417,In_543);
or U3755 (N_3755,In_76,In_429);
or U3756 (N_3756,In_55,In_432);
or U3757 (N_3757,In_303,In_807);
nor U3758 (N_3758,In_440,In_282);
nand U3759 (N_3759,In_861,In_438);
nor U3760 (N_3760,In_452,In_238);
or U3761 (N_3761,In_682,In_584);
and U3762 (N_3762,In_876,In_231);
nand U3763 (N_3763,In_580,In_785);
or U3764 (N_3764,In_85,In_534);
or U3765 (N_3765,In_700,In_308);
nand U3766 (N_3766,In_352,In_870);
nand U3767 (N_3767,In_265,In_672);
nand U3768 (N_3768,In_496,In_869);
nor U3769 (N_3769,In_166,In_336);
xnor U3770 (N_3770,In_437,In_778);
and U3771 (N_3771,In_272,In_84);
or U3772 (N_3772,In_276,In_44);
or U3773 (N_3773,In_812,In_808);
nor U3774 (N_3774,In_99,In_624);
or U3775 (N_3775,In_358,In_508);
nand U3776 (N_3776,In_269,In_18);
and U3777 (N_3777,In_297,In_986);
nor U3778 (N_3778,In_995,In_847);
nor U3779 (N_3779,In_415,In_689);
and U3780 (N_3780,In_341,In_315);
nand U3781 (N_3781,In_697,In_708);
or U3782 (N_3782,In_853,In_408);
nand U3783 (N_3783,In_1,In_823);
nor U3784 (N_3784,In_260,In_880);
or U3785 (N_3785,In_240,In_876);
and U3786 (N_3786,In_225,In_37);
and U3787 (N_3787,In_277,In_651);
nor U3788 (N_3788,In_139,In_175);
and U3789 (N_3789,In_906,In_878);
nand U3790 (N_3790,In_491,In_697);
or U3791 (N_3791,In_747,In_101);
and U3792 (N_3792,In_649,In_941);
or U3793 (N_3793,In_81,In_843);
and U3794 (N_3794,In_582,In_784);
and U3795 (N_3795,In_518,In_371);
nand U3796 (N_3796,In_564,In_380);
or U3797 (N_3797,In_603,In_493);
nand U3798 (N_3798,In_749,In_576);
or U3799 (N_3799,In_255,In_944);
or U3800 (N_3800,In_691,In_973);
or U3801 (N_3801,In_715,In_278);
nand U3802 (N_3802,In_847,In_550);
nand U3803 (N_3803,In_12,In_874);
nor U3804 (N_3804,In_918,In_519);
nand U3805 (N_3805,In_854,In_70);
nand U3806 (N_3806,In_333,In_185);
and U3807 (N_3807,In_739,In_518);
nor U3808 (N_3808,In_150,In_811);
or U3809 (N_3809,In_760,In_602);
or U3810 (N_3810,In_841,In_95);
and U3811 (N_3811,In_664,In_940);
nor U3812 (N_3812,In_997,In_334);
and U3813 (N_3813,In_953,In_87);
nor U3814 (N_3814,In_824,In_419);
nor U3815 (N_3815,In_276,In_335);
nand U3816 (N_3816,In_812,In_611);
and U3817 (N_3817,In_877,In_431);
nor U3818 (N_3818,In_266,In_764);
nand U3819 (N_3819,In_787,In_452);
and U3820 (N_3820,In_411,In_783);
nand U3821 (N_3821,In_96,In_522);
or U3822 (N_3822,In_310,In_663);
and U3823 (N_3823,In_351,In_866);
or U3824 (N_3824,In_701,In_148);
and U3825 (N_3825,In_550,In_477);
nand U3826 (N_3826,In_326,In_395);
or U3827 (N_3827,In_410,In_330);
and U3828 (N_3828,In_748,In_550);
and U3829 (N_3829,In_724,In_709);
or U3830 (N_3830,In_172,In_68);
nor U3831 (N_3831,In_406,In_580);
nand U3832 (N_3832,In_292,In_55);
or U3833 (N_3833,In_333,In_940);
nand U3834 (N_3834,In_918,In_224);
nor U3835 (N_3835,In_412,In_480);
and U3836 (N_3836,In_963,In_627);
and U3837 (N_3837,In_702,In_193);
and U3838 (N_3838,In_638,In_582);
nand U3839 (N_3839,In_928,In_361);
nand U3840 (N_3840,In_108,In_596);
or U3841 (N_3841,In_457,In_429);
nor U3842 (N_3842,In_379,In_20);
nor U3843 (N_3843,In_92,In_617);
and U3844 (N_3844,In_886,In_651);
nand U3845 (N_3845,In_402,In_462);
or U3846 (N_3846,In_586,In_697);
and U3847 (N_3847,In_83,In_619);
and U3848 (N_3848,In_663,In_747);
nand U3849 (N_3849,In_645,In_233);
and U3850 (N_3850,In_478,In_644);
nand U3851 (N_3851,In_758,In_998);
nand U3852 (N_3852,In_929,In_34);
and U3853 (N_3853,In_870,In_843);
or U3854 (N_3854,In_611,In_81);
or U3855 (N_3855,In_984,In_638);
nand U3856 (N_3856,In_483,In_42);
or U3857 (N_3857,In_783,In_649);
nor U3858 (N_3858,In_906,In_581);
or U3859 (N_3859,In_944,In_204);
nand U3860 (N_3860,In_923,In_6);
and U3861 (N_3861,In_412,In_586);
or U3862 (N_3862,In_456,In_960);
or U3863 (N_3863,In_224,In_993);
and U3864 (N_3864,In_808,In_160);
nand U3865 (N_3865,In_923,In_571);
or U3866 (N_3866,In_536,In_976);
and U3867 (N_3867,In_509,In_415);
xnor U3868 (N_3868,In_776,In_157);
nor U3869 (N_3869,In_110,In_273);
nand U3870 (N_3870,In_491,In_354);
or U3871 (N_3871,In_894,In_67);
nand U3872 (N_3872,In_684,In_488);
nor U3873 (N_3873,In_993,In_785);
nor U3874 (N_3874,In_382,In_563);
nand U3875 (N_3875,In_838,In_463);
and U3876 (N_3876,In_336,In_224);
nand U3877 (N_3877,In_346,In_296);
and U3878 (N_3878,In_440,In_641);
nand U3879 (N_3879,In_482,In_52);
nor U3880 (N_3880,In_360,In_698);
nor U3881 (N_3881,In_728,In_41);
nor U3882 (N_3882,In_572,In_505);
nor U3883 (N_3883,In_54,In_767);
and U3884 (N_3884,In_94,In_744);
or U3885 (N_3885,In_642,In_25);
nor U3886 (N_3886,In_587,In_785);
or U3887 (N_3887,In_573,In_9);
nand U3888 (N_3888,In_102,In_98);
nor U3889 (N_3889,In_550,In_36);
nor U3890 (N_3890,In_208,In_408);
nor U3891 (N_3891,In_35,In_213);
nor U3892 (N_3892,In_608,In_734);
nor U3893 (N_3893,In_542,In_190);
or U3894 (N_3894,In_805,In_867);
nand U3895 (N_3895,In_371,In_809);
nor U3896 (N_3896,In_383,In_994);
nor U3897 (N_3897,In_746,In_205);
or U3898 (N_3898,In_589,In_842);
or U3899 (N_3899,In_259,In_819);
nand U3900 (N_3900,In_357,In_528);
nor U3901 (N_3901,In_102,In_947);
or U3902 (N_3902,In_186,In_455);
nor U3903 (N_3903,In_462,In_150);
nand U3904 (N_3904,In_87,In_287);
xor U3905 (N_3905,In_184,In_902);
nand U3906 (N_3906,In_442,In_522);
and U3907 (N_3907,In_508,In_512);
or U3908 (N_3908,In_304,In_164);
nor U3909 (N_3909,In_500,In_52);
or U3910 (N_3910,In_105,In_56);
and U3911 (N_3911,In_756,In_470);
nand U3912 (N_3912,In_894,In_695);
or U3913 (N_3913,In_260,In_710);
nand U3914 (N_3914,In_705,In_949);
nand U3915 (N_3915,In_440,In_378);
nand U3916 (N_3916,In_992,In_117);
nand U3917 (N_3917,In_153,In_137);
and U3918 (N_3918,In_808,In_217);
or U3919 (N_3919,In_858,In_985);
nand U3920 (N_3920,In_432,In_678);
and U3921 (N_3921,In_136,In_938);
xnor U3922 (N_3922,In_130,In_331);
and U3923 (N_3923,In_67,In_862);
nand U3924 (N_3924,In_855,In_818);
nor U3925 (N_3925,In_937,In_865);
or U3926 (N_3926,In_719,In_436);
nor U3927 (N_3927,In_365,In_276);
and U3928 (N_3928,In_715,In_231);
nand U3929 (N_3929,In_658,In_483);
nand U3930 (N_3930,In_990,In_921);
or U3931 (N_3931,In_952,In_928);
nand U3932 (N_3932,In_661,In_982);
nor U3933 (N_3933,In_169,In_702);
nand U3934 (N_3934,In_65,In_190);
and U3935 (N_3935,In_456,In_886);
nand U3936 (N_3936,In_984,In_944);
xor U3937 (N_3937,In_198,In_62);
or U3938 (N_3938,In_969,In_887);
nand U3939 (N_3939,In_389,In_759);
or U3940 (N_3940,In_178,In_729);
nor U3941 (N_3941,In_921,In_388);
or U3942 (N_3942,In_706,In_980);
nand U3943 (N_3943,In_573,In_815);
or U3944 (N_3944,In_305,In_602);
and U3945 (N_3945,In_744,In_718);
nand U3946 (N_3946,In_634,In_937);
nand U3947 (N_3947,In_772,In_770);
and U3948 (N_3948,In_349,In_98);
and U3949 (N_3949,In_858,In_290);
nand U3950 (N_3950,In_281,In_0);
or U3951 (N_3951,In_106,In_527);
or U3952 (N_3952,In_856,In_353);
nor U3953 (N_3953,In_537,In_500);
and U3954 (N_3954,In_756,In_657);
nor U3955 (N_3955,In_483,In_623);
nand U3956 (N_3956,In_270,In_61);
nand U3957 (N_3957,In_285,In_312);
nor U3958 (N_3958,In_520,In_684);
or U3959 (N_3959,In_439,In_574);
and U3960 (N_3960,In_53,In_482);
xor U3961 (N_3961,In_697,In_20);
nand U3962 (N_3962,In_962,In_943);
and U3963 (N_3963,In_513,In_129);
and U3964 (N_3964,In_926,In_898);
and U3965 (N_3965,In_219,In_836);
and U3966 (N_3966,In_960,In_267);
or U3967 (N_3967,In_929,In_576);
nor U3968 (N_3968,In_813,In_535);
nand U3969 (N_3969,In_514,In_469);
nor U3970 (N_3970,In_210,In_104);
nor U3971 (N_3971,In_980,In_792);
and U3972 (N_3972,In_838,In_907);
nand U3973 (N_3973,In_11,In_936);
or U3974 (N_3974,In_724,In_13);
nand U3975 (N_3975,In_697,In_546);
or U3976 (N_3976,In_612,In_229);
nor U3977 (N_3977,In_172,In_647);
nand U3978 (N_3978,In_2,In_558);
or U3979 (N_3979,In_913,In_383);
and U3980 (N_3980,In_300,In_833);
nand U3981 (N_3981,In_492,In_255);
or U3982 (N_3982,In_880,In_380);
nor U3983 (N_3983,In_168,In_194);
nor U3984 (N_3984,In_877,In_369);
or U3985 (N_3985,In_256,In_984);
and U3986 (N_3986,In_546,In_107);
or U3987 (N_3987,In_640,In_269);
nor U3988 (N_3988,In_632,In_240);
nor U3989 (N_3989,In_360,In_507);
nand U3990 (N_3990,In_233,In_257);
and U3991 (N_3991,In_550,In_537);
nor U3992 (N_3992,In_405,In_834);
nand U3993 (N_3993,In_932,In_349);
or U3994 (N_3994,In_608,In_113);
nor U3995 (N_3995,In_199,In_723);
nor U3996 (N_3996,In_930,In_856);
nor U3997 (N_3997,In_466,In_632);
or U3998 (N_3998,In_166,In_680);
and U3999 (N_3999,In_669,In_600);
or U4000 (N_4000,In_775,In_290);
nor U4001 (N_4001,In_643,In_95);
and U4002 (N_4002,In_683,In_892);
and U4003 (N_4003,In_876,In_29);
nor U4004 (N_4004,In_262,In_421);
or U4005 (N_4005,In_546,In_229);
and U4006 (N_4006,In_750,In_682);
or U4007 (N_4007,In_804,In_46);
and U4008 (N_4008,In_56,In_137);
or U4009 (N_4009,In_126,In_664);
and U4010 (N_4010,In_112,In_896);
nand U4011 (N_4011,In_148,In_349);
nor U4012 (N_4012,In_383,In_246);
nand U4013 (N_4013,In_925,In_348);
or U4014 (N_4014,In_520,In_262);
and U4015 (N_4015,In_294,In_566);
or U4016 (N_4016,In_333,In_665);
or U4017 (N_4017,In_584,In_165);
nor U4018 (N_4018,In_479,In_164);
and U4019 (N_4019,In_27,In_771);
and U4020 (N_4020,In_266,In_601);
and U4021 (N_4021,In_594,In_416);
and U4022 (N_4022,In_886,In_955);
nor U4023 (N_4023,In_212,In_275);
or U4024 (N_4024,In_18,In_543);
nor U4025 (N_4025,In_978,In_108);
or U4026 (N_4026,In_314,In_223);
nand U4027 (N_4027,In_190,In_785);
and U4028 (N_4028,In_225,In_563);
and U4029 (N_4029,In_388,In_448);
nor U4030 (N_4030,In_639,In_662);
nor U4031 (N_4031,In_535,In_172);
and U4032 (N_4032,In_990,In_0);
and U4033 (N_4033,In_980,In_822);
or U4034 (N_4034,In_399,In_874);
and U4035 (N_4035,In_856,In_12);
nor U4036 (N_4036,In_57,In_547);
nand U4037 (N_4037,In_749,In_349);
and U4038 (N_4038,In_740,In_405);
nand U4039 (N_4039,In_463,In_176);
and U4040 (N_4040,In_742,In_111);
and U4041 (N_4041,In_254,In_323);
or U4042 (N_4042,In_587,In_820);
or U4043 (N_4043,In_865,In_698);
and U4044 (N_4044,In_926,In_594);
and U4045 (N_4045,In_869,In_148);
nor U4046 (N_4046,In_883,In_645);
and U4047 (N_4047,In_323,In_540);
or U4048 (N_4048,In_572,In_650);
nand U4049 (N_4049,In_736,In_174);
or U4050 (N_4050,In_884,In_488);
or U4051 (N_4051,In_398,In_698);
or U4052 (N_4052,In_968,In_898);
nor U4053 (N_4053,In_315,In_355);
nor U4054 (N_4054,In_249,In_549);
xor U4055 (N_4055,In_905,In_653);
nor U4056 (N_4056,In_664,In_927);
or U4057 (N_4057,In_729,In_262);
nor U4058 (N_4058,In_964,In_387);
nand U4059 (N_4059,In_786,In_559);
nand U4060 (N_4060,In_395,In_19);
or U4061 (N_4061,In_221,In_36);
nor U4062 (N_4062,In_754,In_587);
and U4063 (N_4063,In_291,In_435);
nand U4064 (N_4064,In_938,In_673);
or U4065 (N_4065,In_326,In_479);
or U4066 (N_4066,In_302,In_43);
or U4067 (N_4067,In_482,In_987);
nand U4068 (N_4068,In_576,In_797);
or U4069 (N_4069,In_356,In_861);
nand U4070 (N_4070,In_798,In_510);
nand U4071 (N_4071,In_276,In_217);
nand U4072 (N_4072,In_218,In_228);
xnor U4073 (N_4073,In_306,In_629);
xnor U4074 (N_4074,In_23,In_882);
xor U4075 (N_4075,In_590,In_725);
nor U4076 (N_4076,In_368,In_532);
nor U4077 (N_4077,In_964,In_771);
or U4078 (N_4078,In_242,In_604);
or U4079 (N_4079,In_19,In_312);
nor U4080 (N_4080,In_228,In_946);
nand U4081 (N_4081,In_997,In_381);
and U4082 (N_4082,In_903,In_97);
and U4083 (N_4083,In_65,In_47);
or U4084 (N_4084,In_109,In_387);
or U4085 (N_4085,In_9,In_282);
nand U4086 (N_4086,In_817,In_696);
nor U4087 (N_4087,In_624,In_13);
or U4088 (N_4088,In_520,In_992);
and U4089 (N_4089,In_637,In_275);
nand U4090 (N_4090,In_297,In_609);
or U4091 (N_4091,In_839,In_618);
xor U4092 (N_4092,In_462,In_358);
or U4093 (N_4093,In_855,In_571);
or U4094 (N_4094,In_195,In_384);
or U4095 (N_4095,In_546,In_824);
and U4096 (N_4096,In_758,In_714);
and U4097 (N_4097,In_828,In_87);
or U4098 (N_4098,In_336,In_916);
and U4099 (N_4099,In_580,In_999);
or U4100 (N_4100,In_273,In_8);
and U4101 (N_4101,In_583,In_454);
nand U4102 (N_4102,In_70,In_671);
nor U4103 (N_4103,In_805,In_484);
and U4104 (N_4104,In_946,In_805);
nand U4105 (N_4105,In_680,In_581);
and U4106 (N_4106,In_258,In_921);
or U4107 (N_4107,In_307,In_327);
nor U4108 (N_4108,In_296,In_179);
or U4109 (N_4109,In_601,In_171);
nand U4110 (N_4110,In_235,In_355);
and U4111 (N_4111,In_475,In_938);
and U4112 (N_4112,In_840,In_600);
nand U4113 (N_4113,In_168,In_878);
nand U4114 (N_4114,In_487,In_344);
xnor U4115 (N_4115,In_11,In_925);
nor U4116 (N_4116,In_402,In_696);
nand U4117 (N_4117,In_722,In_221);
or U4118 (N_4118,In_464,In_545);
and U4119 (N_4119,In_120,In_84);
or U4120 (N_4120,In_500,In_769);
nor U4121 (N_4121,In_602,In_922);
nor U4122 (N_4122,In_302,In_494);
or U4123 (N_4123,In_43,In_723);
nor U4124 (N_4124,In_562,In_251);
or U4125 (N_4125,In_106,In_720);
nor U4126 (N_4126,In_966,In_671);
nand U4127 (N_4127,In_5,In_576);
nor U4128 (N_4128,In_25,In_325);
nand U4129 (N_4129,In_875,In_391);
nor U4130 (N_4130,In_163,In_620);
nand U4131 (N_4131,In_753,In_512);
or U4132 (N_4132,In_326,In_545);
nand U4133 (N_4133,In_997,In_66);
or U4134 (N_4134,In_242,In_197);
nor U4135 (N_4135,In_301,In_386);
and U4136 (N_4136,In_569,In_224);
nand U4137 (N_4137,In_216,In_825);
nand U4138 (N_4138,In_187,In_180);
and U4139 (N_4139,In_652,In_816);
nand U4140 (N_4140,In_460,In_818);
nand U4141 (N_4141,In_684,In_289);
nor U4142 (N_4142,In_28,In_360);
nor U4143 (N_4143,In_227,In_640);
and U4144 (N_4144,In_406,In_233);
nand U4145 (N_4145,In_609,In_580);
or U4146 (N_4146,In_777,In_99);
nand U4147 (N_4147,In_486,In_487);
or U4148 (N_4148,In_888,In_219);
nor U4149 (N_4149,In_748,In_357);
or U4150 (N_4150,In_22,In_24);
or U4151 (N_4151,In_832,In_855);
nand U4152 (N_4152,In_321,In_950);
xnor U4153 (N_4153,In_473,In_945);
and U4154 (N_4154,In_206,In_867);
or U4155 (N_4155,In_201,In_756);
and U4156 (N_4156,In_543,In_888);
and U4157 (N_4157,In_635,In_846);
and U4158 (N_4158,In_578,In_899);
nand U4159 (N_4159,In_623,In_219);
and U4160 (N_4160,In_602,In_952);
and U4161 (N_4161,In_470,In_451);
xnor U4162 (N_4162,In_741,In_848);
and U4163 (N_4163,In_656,In_701);
and U4164 (N_4164,In_37,In_447);
nor U4165 (N_4165,In_504,In_957);
or U4166 (N_4166,In_15,In_355);
and U4167 (N_4167,In_845,In_212);
nand U4168 (N_4168,In_269,In_832);
or U4169 (N_4169,In_170,In_582);
and U4170 (N_4170,In_95,In_541);
and U4171 (N_4171,In_254,In_967);
and U4172 (N_4172,In_165,In_176);
or U4173 (N_4173,In_134,In_344);
nor U4174 (N_4174,In_365,In_684);
and U4175 (N_4175,In_18,In_222);
nor U4176 (N_4176,In_40,In_742);
or U4177 (N_4177,In_89,In_670);
nor U4178 (N_4178,In_252,In_110);
and U4179 (N_4179,In_904,In_394);
nand U4180 (N_4180,In_512,In_897);
nor U4181 (N_4181,In_853,In_786);
nand U4182 (N_4182,In_644,In_745);
and U4183 (N_4183,In_386,In_270);
or U4184 (N_4184,In_668,In_968);
nor U4185 (N_4185,In_491,In_25);
and U4186 (N_4186,In_161,In_15);
or U4187 (N_4187,In_169,In_579);
or U4188 (N_4188,In_495,In_292);
nor U4189 (N_4189,In_43,In_419);
xor U4190 (N_4190,In_620,In_799);
nor U4191 (N_4191,In_303,In_600);
nand U4192 (N_4192,In_825,In_873);
and U4193 (N_4193,In_56,In_807);
or U4194 (N_4194,In_201,In_246);
and U4195 (N_4195,In_882,In_985);
xor U4196 (N_4196,In_803,In_618);
and U4197 (N_4197,In_137,In_9);
nor U4198 (N_4198,In_906,In_836);
or U4199 (N_4199,In_738,In_440);
and U4200 (N_4200,In_353,In_103);
nand U4201 (N_4201,In_594,In_768);
or U4202 (N_4202,In_162,In_811);
or U4203 (N_4203,In_179,In_908);
or U4204 (N_4204,In_404,In_599);
nand U4205 (N_4205,In_461,In_418);
or U4206 (N_4206,In_41,In_829);
nor U4207 (N_4207,In_143,In_563);
nand U4208 (N_4208,In_426,In_182);
nor U4209 (N_4209,In_852,In_55);
or U4210 (N_4210,In_333,In_406);
and U4211 (N_4211,In_807,In_616);
nor U4212 (N_4212,In_366,In_326);
or U4213 (N_4213,In_754,In_902);
nor U4214 (N_4214,In_221,In_423);
or U4215 (N_4215,In_771,In_124);
nor U4216 (N_4216,In_22,In_611);
nand U4217 (N_4217,In_731,In_268);
nor U4218 (N_4218,In_810,In_808);
and U4219 (N_4219,In_911,In_554);
nor U4220 (N_4220,In_835,In_504);
nor U4221 (N_4221,In_616,In_178);
nor U4222 (N_4222,In_105,In_369);
nand U4223 (N_4223,In_17,In_114);
or U4224 (N_4224,In_22,In_166);
or U4225 (N_4225,In_306,In_32);
nor U4226 (N_4226,In_507,In_65);
and U4227 (N_4227,In_529,In_31);
nand U4228 (N_4228,In_577,In_772);
nor U4229 (N_4229,In_382,In_312);
and U4230 (N_4230,In_193,In_350);
or U4231 (N_4231,In_686,In_688);
nand U4232 (N_4232,In_124,In_617);
or U4233 (N_4233,In_75,In_722);
and U4234 (N_4234,In_618,In_882);
nand U4235 (N_4235,In_802,In_572);
nand U4236 (N_4236,In_193,In_743);
or U4237 (N_4237,In_713,In_770);
nand U4238 (N_4238,In_106,In_667);
nor U4239 (N_4239,In_852,In_994);
or U4240 (N_4240,In_862,In_16);
or U4241 (N_4241,In_658,In_180);
or U4242 (N_4242,In_798,In_632);
or U4243 (N_4243,In_954,In_318);
nand U4244 (N_4244,In_322,In_783);
or U4245 (N_4245,In_89,In_298);
and U4246 (N_4246,In_125,In_689);
nand U4247 (N_4247,In_283,In_548);
and U4248 (N_4248,In_761,In_753);
nand U4249 (N_4249,In_96,In_736);
nand U4250 (N_4250,In_70,In_931);
and U4251 (N_4251,In_728,In_76);
nor U4252 (N_4252,In_812,In_678);
nor U4253 (N_4253,In_493,In_983);
and U4254 (N_4254,In_163,In_100);
nand U4255 (N_4255,In_677,In_870);
xnor U4256 (N_4256,In_874,In_85);
or U4257 (N_4257,In_665,In_217);
and U4258 (N_4258,In_908,In_67);
or U4259 (N_4259,In_635,In_915);
nor U4260 (N_4260,In_722,In_167);
or U4261 (N_4261,In_257,In_692);
nor U4262 (N_4262,In_501,In_23);
or U4263 (N_4263,In_945,In_821);
nand U4264 (N_4264,In_101,In_586);
nor U4265 (N_4265,In_509,In_469);
and U4266 (N_4266,In_181,In_651);
nor U4267 (N_4267,In_804,In_755);
nand U4268 (N_4268,In_136,In_560);
or U4269 (N_4269,In_505,In_493);
nor U4270 (N_4270,In_396,In_80);
and U4271 (N_4271,In_251,In_754);
and U4272 (N_4272,In_893,In_697);
nor U4273 (N_4273,In_411,In_72);
and U4274 (N_4274,In_743,In_663);
nand U4275 (N_4275,In_967,In_359);
and U4276 (N_4276,In_522,In_224);
and U4277 (N_4277,In_894,In_161);
and U4278 (N_4278,In_517,In_757);
and U4279 (N_4279,In_411,In_782);
and U4280 (N_4280,In_946,In_297);
nand U4281 (N_4281,In_853,In_995);
nand U4282 (N_4282,In_957,In_825);
or U4283 (N_4283,In_580,In_308);
and U4284 (N_4284,In_350,In_524);
nor U4285 (N_4285,In_301,In_486);
nand U4286 (N_4286,In_184,In_550);
and U4287 (N_4287,In_586,In_334);
nor U4288 (N_4288,In_696,In_826);
nand U4289 (N_4289,In_622,In_991);
or U4290 (N_4290,In_969,In_251);
nor U4291 (N_4291,In_306,In_407);
or U4292 (N_4292,In_817,In_289);
or U4293 (N_4293,In_378,In_422);
and U4294 (N_4294,In_184,In_741);
or U4295 (N_4295,In_699,In_982);
nand U4296 (N_4296,In_233,In_788);
and U4297 (N_4297,In_675,In_43);
nand U4298 (N_4298,In_628,In_188);
nand U4299 (N_4299,In_126,In_815);
and U4300 (N_4300,In_558,In_643);
nand U4301 (N_4301,In_609,In_847);
nor U4302 (N_4302,In_307,In_809);
and U4303 (N_4303,In_714,In_326);
nand U4304 (N_4304,In_890,In_927);
nor U4305 (N_4305,In_963,In_985);
and U4306 (N_4306,In_20,In_276);
nor U4307 (N_4307,In_140,In_38);
nand U4308 (N_4308,In_362,In_569);
nor U4309 (N_4309,In_475,In_613);
nand U4310 (N_4310,In_982,In_848);
nand U4311 (N_4311,In_49,In_673);
nor U4312 (N_4312,In_852,In_894);
or U4313 (N_4313,In_187,In_918);
nor U4314 (N_4314,In_461,In_93);
and U4315 (N_4315,In_120,In_439);
nor U4316 (N_4316,In_188,In_841);
nor U4317 (N_4317,In_765,In_80);
nand U4318 (N_4318,In_892,In_317);
or U4319 (N_4319,In_734,In_357);
nor U4320 (N_4320,In_50,In_625);
or U4321 (N_4321,In_372,In_385);
and U4322 (N_4322,In_282,In_339);
and U4323 (N_4323,In_90,In_533);
nand U4324 (N_4324,In_573,In_949);
nand U4325 (N_4325,In_123,In_152);
nor U4326 (N_4326,In_546,In_440);
nor U4327 (N_4327,In_51,In_60);
or U4328 (N_4328,In_708,In_365);
nor U4329 (N_4329,In_638,In_770);
and U4330 (N_4330,In_65,In_163);
xor U4331 (N_4331,In_402,In_438);
nor U4332 (N_4332,In_676,In_967);
or U4333 (N_4333,In_466,In_692);
and U4334 (N_4334,In_601,In_793);
nor U4335 (N_4335,In_616,In_634);
nand U4336 (N_4336,In_969,In_987);
and U4337 (N_4337,In_80,In_418);
nor U4338 (N_4338,In_174,In_81);
nand U4339 (N_4339,In_976,In_199);
nor U4340 (N_4340,In_835,In_780);
nor U4341 (N_4341,In_835,In_136);
nor U4342 (N_4342,In_545,In_537);
or U4343 (N_4343,In_316,In_379);
nand U4344 (N_4344,In_230,In_903);
and U4345 (N_4345,In_414,In_611);
nor U4346 (N_4346,In_124,In_164);
nor U4347 (N_4347,In_875,In_191);
nor U4348 (N_4348,In_581,In_386);
nor U4349 (N_4349,In_926,In_263);
and U4350 (N_4350,In_381,In_266);
or U4351 (N_4351,In_884,In_536);
nor U4352 (N_4352,In_490,In_458);
and U4353 (N_4353,In_510,In_254);
nand U4354 (N_4354,In_714,In_760);
or U4355 (N_4355,In_873,In_458);
or U4356 (N_4356,In_821,In_362);
nor U4357 (N_4357,In_786,In_319);
nor U4358 (N_4358,In_109,In_363);
or U4359 (N_4359,In_76,In_923);
or U4360 (N_4360,In_816,In_876);
nand U4361 (N_4361,In_636,In_12);
or U4362 (N_4362,In_813,In_98);
and U4363 (N_4363,In_743,In_728);
nor U4364 (N_4364,In_760,In_808);
or U4365 (N_4365,In_383,In_101);
xnor U4366 (N_4366,In_452,In_417);
xnor U4367 (N_4367,In_615,In_736);
and U4368 (N_4368,In_134,In_503);
nor U4369 (N_4369,In_566,In_768);
nor U4370 (N_4370,In_552,In_640);
nor U4371 (N_4371,In_746,In_262);
nor U4372 (N_4372,In_771,In_312);
and U4373 (N_4373,In_697,In_510);
nand U4374 (N_4374,In_282,In_288);
or U4375 (N_4375,In_120,In_808);
or U4376 (N_4376,In_918,In_564);
xor U4377 (N_4377,In_0,In_127);
nor U4378 (N_4378,In_533,In_348);
and U4379 (N_4379,In_308,In_396);
and U4380 (N_4380,In_7,In_359);
nand U4381 (N_4381,In_131,In_746);
or U4382 (N_4382,In_832,In_393);
or U4383 (N_4383,In_638,In_37);
nor U4384 (N_4384,In_691,In_37);
nand U4385 (N_4385,In_244,In_967);
or U4386 (N_4386,In_839,In_324);
or U4387 (N_4387,In_667,In_372);
nand U4388 (N_4388,In_156,In_165);
nand U4389 (N_4389,In_79,In_783);
or U4390 (N_4390,In_659,In_925);
nand U4391 (N_4391,In_50,In_392);
nor U4392 (N_4392,In_650,In_629);
and U4393 (N_4393,In_203,In_24);
and U4394 (N_4394,In_256,In_315);
nor U4395 (N_4395,In_175,In_90);
nor U4396 (N_4396,In_886,In_717);
nand U4397 (N_4397,In_440,In_160);
and U4398 (N_4398,In_673,In_146);
and U4399 (N_4399,In_802,In_586);
or U4400 (N_4400,In_71,In_94);
or U4401 (N_4401,In_277,In_836);
nor U4402 (N_4402,In_238,In_19);
nor U4403 (N_4403,In_300,In_774);
or U4404 (N_4404,In_319,In_774);
nor U4405 (N_4405,In_712,In_822);
and U4406 (N_4406,In_429,In_208);
nor U4407 (N_4407,In_390,In_591);
nor U4408 (N_4408,In_523,In_45);
and U4409 (N_4409,In_617,In_73);
nor U4410 (N_4410,In_834,In_837);
nand U4411 (N_4411,In_896,In_575);
and U4412 (N_4412,In_206,In_982);
nand U4413 (N_4413,In_649,In_458);
and U4414 (N_4414,In_502,In_909);
or U4415 (N_4415,In_654,In_411);
nand U4416 (N_4416,In_150,In_637);
nor U4417 (N_4417,In_44,In_872);
or U4418 (N_4418,In_135,In_74);
nor U4419 (N_4419,In_492,In_949);
nor U4420 (N_4420,In_4,In_387);
nor U4421 (N_4421,In_127,In_418);
or U4422 (N_4422,In_327,In_309);
and U4423 (N_4423,In_95,In_756);
or U4424 (N_4424,In_139,In_509);
or U4425 (N_4425,In_764,In_480);
or U4426 (N_4426,In_989,In_386);
nand U4427 (N_4427,In_120,In_85);
or U4428 (N_4428,In_345,In_184);
and U4429 (N_4429,In_696,In_963);
nor U4430 (N_4430,In_175,In_468);
or U4431 (N_4431,In_84,In_939);
nor U4432 (N_4432,In_753,In_784);
or U4433 (N_4433,In_186,In_15);
or U4434 (N_4434,In_214,In_24);
or U4435 (N_4435,In_356,In_545);
nor U4436 (N_4436,In_79,In_949);
nor U4437 (N_4437,In_335,In_984);
nor U4438 (N_4438,In_665,In_223);
and U4439 (N_4439,In_972,In_26);
and U4440 (N_4440,In_15,In_948);
nor U4441 (N_4441,In_688,In_307);
nand U4442 (N_4442,In_728,In_605);
nand U4443 (N_4443,In_900,In_860);
nand U4444 (N_4444,In_310,In_662);
or U4445 (N_4445,In_559,In_527);
nor U4446 (N_4446,In_239,In_877);
and U4447 (N_4447,In_373,In_713);
nand U4448 (N_4448,In_223,In_641);
nor U4449 (N_4449,In_938,In_426);
or U4450 (N_4450,In_546,In_138);
nor U4451 (N_4451,In_780,In_868);
or U4452 (N_4452,In_980,In_745);
nand U4453 (N_4453,In_929,In_488);
and U4454 (N_4454,In_561,In_856);
and U4455 (N_4455,In_905,In_875);
nand U4456 (N_4456,In_498,In_299);
nor U4457 (N_4457,In_72,In_682);
nor U4458 (N_4458,In_20,In_321);
or U4459 (N_4459,In_645,In_242);
or U4460 (N_4460,In_454,In_187);
or U4461 (N_4461,In_777,In_109);
and U4462 (N_4462,In_136,In_703);
nor U4463 (N_4463,In_341,In_502);
and U4464 (N_4464,In_732,In_401);
or U4465 (N_4465,In_518,In_615);
nand U4466 (N_4466,In_270,In_584);
nand U4467 (N_4467,In_691,In_726);
or U4468 (N_4468,In_736,In_270);
or U4469 (N_4469,In_531,In_402);
nand U4470 (N_4470,In_999,In_676);
and U4471 (N_4471,In_248,In_150);
nand U4472 (N_4472,In_440,In_991);
and U4473 (N_4473,In_273,In_640);
or U4474 (N_4474,In_928,In_135);
or U4475 (N_4475,In_102,In_237);
and U4476 (N_4476,In_438,In_697);
nand U4477 (N_4477,In_51,In_127);
and U4478 (N_4478,In_28,In_371);
or U4479 (N_4479,In_567,In_294);
nand U4480 (N_4480,In_283,In_832);
and U4481 (N_4481,In_269,In_717);
nand U4482 (N_4482,In_753,In_158);
nand U4483 (N_4483,In_227,In_364);
nor U4484 (N_4484,In_503,In_77);
nand U4485 (N_4485,In_883,In_748);
and U4486 (N_4486,In_184,In_101);
nand U4487 (N_4487,In_289,In_413);
and U4488 (N_4488,In_870,In_99);
or U4489 (N_4489,In_5,In_697);
nor U4490 (N_4490,In_953,In_431);
nor U4491 (N_4491,In_802,In_694);
and U4492 (N_4492,In_869,In_714);
xor U4493 (N_4493,In_303,In_318);
or U4494 (N_4494,In_3,In_41);
nor U4495 (N_4495,In_433,In_64);
nand U4496 (N_4496,In_777,In_341);
and U4497 (N_4497,In_974,In_863);
and U4498 (N_4498,In_291,In_133);
nor U4499 (N_4499,In_363,In_309);
nand U4500 (N_4500,In_743,In_855);
and U4501 (N_4501,In_549,In_359);
xor U4502 (N_4502,In_281,In_544);
nand U4503 (N_4503,In_888,In_862);
nor U4504 (N_4504,In_924,In_477);
nand U4505 (N_4505,In_160,In_9);
and U4506 (N_4506,In_391,In_85);
nor U4507 (N_4507,In_887,In_144);
nor U4508 (N_4508,In_711,In_269);
or U4509 (N_4509,In_56,In_534);
nand U4510 (N_4510,In_384,In_838);
or U4511 (N_4511,In_675,In_412);
nor U4512 (N_4512,In_468,In_278);
or U4513 (N_4513,In_674,In_215);
or U4514 (N_4514,In_398,In_178);
and U4515 (N_4515,In_50,In_353);
or U4516 (N_4516,In_271,In_81);
or U4517 (N_4517,In_518,In_528);
and U4518 (N_4518,In_385,In_547);
nor U4519 (N_4519,In_652,In_408);
and U4520 (N_4520,In_239,In_872);
and U4521 (N_4521,In_91,In_507);
nor U4522 (N_4522,In_949,In_313);
and U4523 (N_4523,In_11,In_515);
or U4524 (N_4524,In_325,In_725);
or U4525 (N_4525,In_397,In_515);
or U4526 (N_4526,In_65,In_710);
or U4527 (N_4527,In_290,In_714);
or U4528 (N_4528,In_247,In_129);
nand U4529 (N_4529,In_979,In_139);
nand U4530 (N_4530,In_376,In_522);
or U4531 (N_4531,In_944,In_764);
nor U4532 (N_4532,In_270,In_838);
nor U4533 (N_4533,In_593,In_617);
or U4534 (N_4534,In_936,In_922);
nand U4535 (N_4535,In_340,In_705);
nor U4536 (N_4536,In_956,In_470);
or U4537 (N_4537,In_922,In_758);
nor U4538 (N_4538,In_475,In_602);
nor U4539 (N_4539,In_60,In_485);
nor U4540 (N_4540,In_951,In_843);
nor U4541 (N_4541,In_397,In_113);
or U4542 (N_4542,In_169,In_26);
or U4543 (N_4543,In_865,In_715);
nor U4544 (N_4544,In_857,In_691);
nor U4545 (N_4545,In_448,In_60);
or U4546 (N_4546,In_526,In_743);
nand U4547 (N_4547,In_473,In_423);
and U4548 (N_4548,In_43,In_557);
or U4549 (N_4549,In_906,In_153);
or U4550 (N_4550,In_70,In_65);
nor U4551 (N_4551,In_294,In_646);
nor U4552 (N_4552,In_98,In_146);
nand U4553 (N_4553,In_590,In_61);
and U4554 (N_4554,In_396,In_822);
or U4555 (N_4555,In_357,In_994);
nand U4556 (N_4556,In_848,In_892);
nor U4557 (N_4557,In_640,In_338);
nand U4558 (N_4558,In_809,In_955);
nand U4559 (N_4559,In_653,In_814);
xor U4560 (N_4560,In_916,In_299);
nor U4561 (N_4561,In_936,In_537);
or U4562 (N_4562,In_955,In_248);
nor U4563 (N_4563,In_140,In_567);
or U4564 (N_4564,In_566,In_841);
and U4565 (N_4565,In_931,In_800);
nand U4566 (N_4566,In_933,In_711);
or U4567 (N_4567,In_380,In_265);
and U4568 (N_4568,In_306,In_528);
nand U4569 (N_4569,In_145,In_253);
nand U4570 (N_4570,In_595,In_894);
nand U4571 (N_4571,In_36,In_714);
and U4572 (N_4572,In_345,In_435);
nand U4573 (N_4573,In_403,In_897);
and U4574 (N_4574,In_619,In_806);
and U4575 (N_4575,In_972,In_855);
or U4576 (N_4576,In_663,In_478);
nor U4577 (N_4577,In_903,In_558);
and U4578 (N_4578,In_921,In_282);
nand U4579 (N_4579,In_118,In_14);
nor U4580 (N_4580,In_281,In_878);
or U4581 (N_4581,In_818,In_232);
or U4582 (N_4582,In_372,In_147);
nor U4583 (N_4583,In_119,In_9);
and U4584 (N_4584,In_157,In_628);
nor U4585 (N_4585,In_736,In_563);
nand U4586 (N_4586,In_642,In_926);
nor U4587 (N_4587,In_397,In_231);
nand U4588 (N_4588,In_533,In_422);
and U4589 (N_4589,In_152,In_385);
and U4590 (N_4590,In_265,In_661);
nand U4591 (N_4591,In_878,In_130);
and U4592 (N_4592,In_507,In_89);
or U4593 (N_4593,In_283,In_696);
and U4594 (N_4594,In_978,In_162);
or U4595 (N_4595,In_257,In_312);
or U4596 (N_4596,In_520,In_406);
xnor U4597 (N_4597,In_464,In_335);
and U4598 (N_4598,In_354,In_992);
nand U4599 (N_4599,In_4,In_775);
nor U4600 (N_4600,In_670,In_82);
nand U4601 (N_4601,In_2,In_933);
nor U4602 (N_4602,In_333,In_541);
and U4603 (N_4603,In_556,In_796);
nor U4604 (N_4604,In_432,In_751);
nand U4605 (N_4605,In_619,In_328);
or U4606 (N_4606,In_870,In_790);
nand U4607 (N_4607,In_843,In_975);
or U4608 (N_4608,In_661,In_639);
nand U4609 (N_4609,In_472,In_269);
and U4610 (N_4610,In_102,In_970);
nand U4611 (N_4611,In_50,In_861);
or U4612 (N_4612,In_988,In_537);
nor U4613 (N_4613,In_353,In_749);
nor U4614 (N_4614,In_413,In_732);
nor U4615 (N_4615,In_368,In_467);
nor U4616 (N_4616,In_966,In_200);
nand U4617 (N_4617,In_928,In_769);
nand U4618 (N_4618,In_602,In_119);
and U4619 (N_4619,In_993,In_191);
nor U4620 (N_4620,In_189,In_534);
nand U4621 (N_4621,In_240,In_599);
nand U4622 (N_4622,In_830,In_0);
nand U4623 (N_4623,In_469,In_746);
nand U4624 (N_4624,In_856,In_812);
or U4625 (N_4625,In_869,In_812);
or U4626 (N_4626,In_201,In_465);
or U4627 (N_4627,In_663,In_692);
or U4628 (N_4628,In_559,In_565);
or U4629 (N_4629,In_300,In_579);
and U4630 (N_4630,In_693,In_760);
nor U4631 (N_4631,In_338,In_947);
or U4632 (N_4632,In_532,In_561);
or U4633 (N_4633,In_21,In_624);
nor U4634 (N_4634,In_524,In_860);
xnor U4635 (N_4635,In_152,In_671);
and U4636 (N_4636,In_869,In_843);
or U4637 (N_4637,In_266,In_551);
nand U4638 (N_4638,In_443,In_555);
and U4639 (N_4639,In_460,In_501);
and U4640 (N_4640,In_278,In_435);
nor U4641 (N_4641,In_298,In_10);
and U4642 (N_4642,In_292,In_277);
or U4643 (N_4643,In_944,In_825);
xor U4644 (N_4644,In_96,In_201);
nor U4645 (N_4645,In_724,In_101);
and U4646 (N_4646,In_787,In_639);
nand U4647 (N_4647,In_60,In_610);
or U4648 (N_4648,In_593,In_691);
and U4649 (N_4649,In_808,In_897);
or U4650 (N_4650,In_449,In_914);
nand U4651 (N_4651,In_467,In_857);
nand U4652 (N_4652,In_897,In_527);
nor U4653 (N_4653,In_622,In_438);
or U4654 (N_4654,In_522,In_51);
and U4655 (N_4655,In_322,In_768);
nor U4656 (N_4656,In_826,In_717);
or U4657 (N_4657,In_40,In_108);
nor U4658 (N_4658,In_607,In_503);
and U4659 (N_4659,In_468,In_810);
or U4660 (N_4660,In_253,In_454);
nand U4661 (N_4661,In_886,In_825);
nor U4662 (N_4662,In_928,In_800);
nand U4663 (N_4663,In_875,In_2);
nand U4664 (N_4664,In_760,In_923);
nand U4665 (N_4665,In_25,In_92);
nand U4666 (N_4666,In_588,In_372);
nor U4667 (N_4667,In_378,In_19);
and U4668 (N_4668,In_38,In_265);
and U4669 (N_4669,In_145,In_327);
nor U4670 (N_4670,In_57,In_343);
nor U4671 (N_4671,In_824,In_326);
nand U4672 (N_4672,In_676,In_450);
and U4673 (N_4673,In_285,In_538);
nor U4674 (N_4674,In_214,In_230);
or U4675 (N_4675,In_210,In_701);
or U4676 (N_4676,In_998,In_641);
and U4677 (N_4677,In_351,In_846);
nor U4678 (N_4678,In_910,In_387);
or U4679 (N_4679,In_264,In_267);
nor U4680 (N_4680,In_593,In_707);
nand U4681 (N_4681,In_29,In_171);
or U4682 (N_4682,In_252,In_628);
and U4683 (N_4683,In_84,In_952);
and U4684 (N_4684,In_956,In_981);
xor U4685 (N_4685,In_271,In_362);
and U4686 (N_4686,In_620,In_583);
nand U4687 (N_4687,In_480,In_970);
or U4688 (N_4688,In_38,In_370);
and U4689 (N_4689,In_124,In_402);
nor U4690 (N_4690,In_173,In_152);
or U4691 (N_4691,In_175,In_856);
nor U4692 (N_4692,In_252,In_761);
or U4693 (N_4693,In_453,In_752);
or U4694 (N_4694,In_869,In_34);
nor U4695 (N_4695,In_984,In_849);
or U4696 (N_4696,In_716,In_899);
or U4697 (N_4697,In_329,In_248);
nor U4698 (N_4698,In_989,In_743);
or U4699 (N_4699,In_119,In_233);
nand U4700 (N_4700,In_700,In_657);
nor U4701 (N_4701,In_945,In_138);
and U4702 (N_4702,In_330,In_620);
nand U4703 (N_4703,In_861,In_498);
nor U4704 (N_4704,In_408,In_969);
nand U4705 (N_4705,In_811,In_971);
and U4706 (N_4706,In_543,In_676);
xnor U4707 (N_4707,In_939,In_75);
and U4708 (N_4708,In_34,In_775);
nand U4709 (N_4709,In_840,In_336);
or U4710 (N_4710,In_54,In_423);
or U4711 (N_4711,In_929,In_182);
or U4712 (N_4712,In_924,In_847);
or U4713 (N_4713,In_536,In_331);
nor U4714 (N_4714,In_691,In_925);
nor U4715 (N_4715,In_865,In_179);
nand U4716 (N_4716,In_436,In_457);
and U4717 (N_4717,In_922,In_431);
or U4718 (N_4718,In_574,In_993);
or U4719 (N_4719,In_941,In_677);
and U4720 (N_4720,In_524,In_294);
nand U4721 (N_4721,In_607,In_969);
nor U4722 (N_4722,In_92,In_638);
nor U4723 (N_4723,In_374,In_630);
nand U4724 (N_4724,In_623,In_845);
and U4725 (N_4725,In_677,In_639);
and U4726 (N_4726,In_189,In_173);
or U4727 (N_4727,In_555,In_562);
nand U4728 (N_4728,In_673,In_874);
or U4729 (N_4729,In_767,In_45);
nand U4730 (N_4730,In_513,In_153);
nor U4731 (N_4731,In_388,In_688);
and U4732 (N_4732,In_816,In_215);
nand U4733 (N_4733,In_37,In_92);
and U4734 (N_4734,In_497,In_258);
or U4735 (N_4735,In_11,In_907);
or U4736 (N_4736,In_362,In_18);
nor U4737 (N_4737,In_542,In_729);
nor U4738 (N_4738,In_454,In_346);
or U4739 (N_4739,In_162,In_257);
nand U4740 (N_4740,In_200,In_545);
and U4741 (N_4741,In_581,In_381);
nand U4742 (N_4742,In_430,In_894);
or U4743 (N_4743,In_128,In_764);
nand U4744 (N_4744,In_752,In_391);
and U4745 (N_4745,In_106,In_513);
and U4746 (N_4746,In_318,In_888);
nor U4747 (N_4747,In_612,In_444);
and U4748 (N_4748,In_481,In_292);
nor U4749 (N_4749,In_393,In_73);
nand U4750 (N_4750,In_994,In_36);
xor U4751 (N_4751,In_922,In_976);
or U4752 (N_4752,In_733,In_226);
nand U4753 (N_4753,In_757,In_463);
and U4754 (N_4754,In_106,In_884);
and U4755 (N_4755,In_127,In_892);
and U4756 (N_4756,In_774,In_288);
nor U4757 (N_4757,In_939,In_6);
or U4758 (N_4758,In_248,In_261);
nor U4759 (N_4759,In_296,In_953);
and U4760 (N_4760,In_249,In_879);
and U4761 (N_4761,In_72,In_473);
and U4762 (N_4762,In_913,In_904);
or U4763 (N_4763,In_328,In_916);
or U4764 (N_4764,In_729,In_460);
and U4765 (N_4765,In_516,In_225);
nor U4766 (N_4766,In_965,In_106);
and U4767 (N_4767,In_934,In_265);
nand U4768 (N_4768,In_999,In_981);
nand U4769 (N_4769,In_220,In_805);
and U4770 (N_4770,In_117,In_531);
and U4771 (N_4771,In_283,In_664);
or U4772 (N_4772,In_54,In_924);
or U4773 (N_4773,In_570,In_551);
and U4774 (N_4774,In_892,In_780);
or U4775 (N_4775,In_342,In_151);
xnor U4776 (N_4776,In_162,In_881);
nand U4777 (N_4777,In_831,In_745);
and U4778 (N_4778,In_691,In_148);
or U4779 (N_4779,In_297,In_811);
xor U4780 (N_4780,In_49,In_373);
nor U4781 (N_4781,In_688,In_317);
nor U4782 (N_4782,In_149,In_925);
nor U4783 (N_4783,In_799,In_557);
nor U4784 (N_4784,In_54,In_135);
nand U4785 (N_4785,In_157,In_544);
nor U4786 (N_4786,In_153,In_721);
and U4787 (N_4787,In_926,In_948);
nand U4788 (N_4788,In_724,In_633);
and U4789 (N_4789,In_605,In_440);
xor U4790 (N_4790,In_216,In_848);
or U4791 (N_4791,In_355,In_26);
and U4792 (N_4792,In_255,In_410);
nand U4793 (N_4793,In_301,In_127);
or U4794 (N_4794,In_749,In_477);
or U4795 (N_4795,In_510,In_319);
and U4796 (N_4796,In_61,In_796);
nor U4797 (N_4797,In_91,In_571);
nand U4798 (N_4798,In_801,In_25);
nand U4799 (N_4799,In_63,In_941);
or U4800 (N_4800,In_898,In_296);
and U4801 (N_4801,In_961,In_732);
nand U4802 (N_4802,In_558,In_895);
nand U4803 (N_4803,In_721,In_352);
or U4804 (N_4804,In_609,In_787);
nand U4805 (N_4805,In_45,In_535);
or U4806 (N_4806,In_321,In_162);
and U4807 (N_4807,In_457,In_682);
nor U4808 (N_4808,In_958,In_994);
and U4809 (N_4809,In_334,In_398);
or U4810 (N_4810,In_232,In_572);
nand U4811 (N_4811,In_557,In_836);
and U4812 (N_4812,In_579,In_211);
and U4813 (N_4813,In_557,In_559);
nand U4814 (N_4814,In_998,In_899);
or U4815 (N_4815,In_472,In_205);
nor U4816 (N_4816,In_161,In_893);
nand U4817 (N_4817,In_591,In_44);
and U4818 (N_4818,In_720,In_194);
and U4819 (N_4819,In_793,In_825);
or U4820 (N_4820,In_463,In_355);
and U4821 (N_4821,In_15,In_165);
and U4822 (N_4822,In_359,In_840);
or U4823 (N_4823,In_358,In_665);
nand U4824 (N_4824,In_742,In_228);
nor U4825 (N_4825,In_174,In_474);
nor U4826 (N_4826,In_508,In_110);
nor U4827 (N_4827,In_972,In_64);
nand U4828 (N_4828,In_943,In_672);
nand U4829 (N_4829,In_558,In_641);
and U4830 (N_4830,In_777,In_648);
nand U4831 (N_4831,In_758,In_597);
or U4832 (N_4832,In_323,In_39);
or U4833 (N_4833,In_299,In_853);
nand U4834 (N_4834,In_570,In_731);
nor U4835 (N_4835,In_885,In_703);
nand U4836 (N_4836,In_689,In_797);
nor U4837 (N_4837,In_185,In_321);
and U4838 (N_4838,In_942,In_534);
nor U4839 (N_4839,In_117,In_955);
nor U4840 (N_4840,In_691,In_723);
nand U4841 (N_4841,In_664,In_266);
and U4842 (N_4842,In_950,In_298);
and U4843 (N_4843,In_675,In_929);
nand U4844 (N_4844,In_137,In_196);
or U4845 (N_4845,In_595,In_153);
and U4846 (N_4846,In_279,In_273);
and U4847 (N_4847,In_846,In_41);
nand U4848 (N_4848,In_298,In_62);
nor U4849 (N_4849,In_301,In_45);
nor U4850 (N_4850,In_272,In_212);
or U4851 (N_4851,In_318,In_875);
and U4852 (N_4852,In_17,In_870);
nor U4853 (N_4853,In_232,In_672);
or U4854 (N_4854,In_194,In_538);
and U4855 (N_4855,In_949,In_117);
and U4856 (N_4856,In_777,In_982);
nand U4857 (N_4857,In_444,In_88);
nor U4858 (N_4858,In_102,In_903);
nand U4859 (N_4859,In_269,In_870);
and U4860 (N_4860,In_642,In_240);
and U4861 (N_4861,In_553,In_318);
nand U4862 (N_4862,In_167,In_663);
nand U4863 (N_4863,In_975,In_907);
and U4864 (N_4864,In_258,In_462);
nor U4865 (N_4865,In_102,In_96);
nor U4866 (N_4866,In_144,In_769);
nand U4867 (N_4867,In_138,In_161);
nor U4868 (N_4868,In_834,In_747);
nor U4869 (N_4869,In_323,In_315);
and U4870 (N_4870,In_399,In_523);
nand U4871 (N_4871,In_173,In_259);
nand U4872 (N_4872,In_950,In_944);
nand U4873 (N_4873,In_556,In_531);
and U4874 (N_4874,In_594,In_620);
xnor U4875 (N_4875,In_121,In_583);
nor U4876 (N_4876,In_639,In_243);
and U4877 (N_4877,In_19,In_873);
nor U4878 (N_4878,In_64,In_590);
or U4879 (N_4879,In_564,In_799);
or U4880 (N_4880,In_312,In_414);
nand U4881 (N_4881,In_89,In_490);
nand U4882 (N_4882,In_755,In_277);
nand U4883 (N_4883,In_176,In_33);
or U4884 (N_4884,In_340,In_466);
nor U4885 (N_4885,In_901,In_782);
or U4886 (N_4886,In_160,In_564);
nand U4887 (N_4887,In_251,In_131);
nand U4888 (N_4888,In_236,In_313);
nor U4889 (N_4889,In_290,In_182);
nand U4890 (N_4890,In_408,In_67);
xnor U4891 (N_4891,In_779,In_274);
nand U4892 (N_4892,In_342,In_296);
nor U4893 (N_4893,In_334,In_313);
or U4894 (N_4894,In_5,In_174);
nand U4895 (N_4895,In_864,In_314);
and U4896 (N_4896,In_572,In_982);
or U4897 (N_4897,In_555,In_634);
and U4898 (N_4898,In_513,In_683);
xor U4899 (N_4899,In_495,In_468);
or U4900 (N_4900,In_707,In_249);
and U4901 (N_4901,In_824,In_265);
and U4902 (N_4902,In_787,In_47);
and U4903 (N_4903,In_911,In_75);
nor U4904 (N_4904,In_884,In_309);
and U4905 (N_4905,In_83,In_553);
nand U4906 (N_4906,In_605,In_115);
or U4907 (N_4907,In_192,In_743);
and U4908 (N_4908,In_642,In_266);
or U4909 (N_4909,In_675,In_893);
nand U4910 (N_4910,In_833,In_440);
and U4911 (N_4911,In_135,In_322);
and U4912 (N_4912,In_657,In_744);
nor U4913 (N_4913,In_575,In_515);
and U4914 (N_4914,In_782,In_379);
nor U4915 (N_4915,In_779,In_798);
nor U4916 (N_4916,In_788,In_200);
or U4917 (N_4917,In_224,In_602);
xor U4918 (N_4918,In_44,In_879);
nand U4919 (N_4919,In_466,In_829);
xnor U4920 (N_4920,In_747,In_529);
nand U4921 (N_4921,In_140,In_663);
and U4922 (N_4922,In_423,In_220);
or U4923 (N_4923,In_855,In_276);
nand U4924 (N_4924,In_319,In_479);
or U4925 (N_4925,In_336,In_323);
or U4926 (N_4926,In_819,In_22);
or U4927 (N_4927,In_32,In_56);
nand U4928 (N_4928,In_452,In_198);
nand U4929 (N_4929,In_368,In_911);
nor U4930 (N_4930,In_475,In_399);
and U4931 (N_4931,In_457,In_683);
nand U4932 (N_4932,In_278,In_807);
and U4933 (N_4933,In_867,In_620);
nand U4934 (N_4934,In_376,In_388);
nand U4935 (N_4935,In_490,In_814);
or U4936 (N_4936,In_629,In_905);
nand U4937 (N_4937,In_944,In_327);
nand U4938 (N_4938,In_613,In_968);
nand U4939 (N_4939,In_341,In_871);
nor U4940 (N_4940,In_671,In_402);
nor U4941 (N_4941,In_818,In_638);
xnor U4942 (N_4942,In_346,In_348);
or U4943 (N_4943,In_48,In_352);
and U4944 (N_4944,In_923,In_249);
nor U4945 (N_4945,In_367,In_413);
nand U4946 (N_4946,In_900,In_809);
or U4947 (N_4947,In_770,In_317);
or U4948 (N_4948,In_386,In_473);
nor U4949 (N_4949,In_374,In_719);
nor U4950 (N_4950,In_841,In_217);
or U4951 (N_4951,In_365,In_956);
or U4952 (N_4952,In_101,In_581);
and U4953 (N_4953,In_551,In_392);
nand U4954 (N_4954,In_191,In_449);
nor U4955 (N_4955,In_858,In_503);
and U4956 (N_4956,In_467,In_838);
nand U4957 (N_4957,In_647,In_295);
and U4958 (N_4958,In_21,In_245);
and U4959 (N_4959,In_940,In_481);
and U4960 (N_4960,In_375,In_428);
and U4961 (N_4961,In_93,In_415);
nand U4962 (N_4962,In_909,In_692);
or U4963 (N_4963,In_333,In_938);
nor U4964 (N_4964,In_742,In_322);
and U4965 (N_4965,In_630,In_31);
xor U4966 (N_4966,In_246,In_903);
nand U4967 (N_4967,In_115,In_6);
and U4968 (N_4968,In_915,In_601);
or U4969 (N_4969,In_658,In_688);
and U4970 (N_4970,In_296,In_984);
and U4971 (N_4971,In_321,In_410);
or U4972 (N_4972,In_271,In_232);
or U4973 (N_4973,In_744,In_269);
and U4974 (N_4974,In_658,In_446);
and U4975 (N_4975,In_784,In_361);
nand U4976 (N_4976,In_322,In_521);
nand U4977 (N_4977,In_323,In_665);
nand U4978 (N_4978,In_513,In_892);
nor U4979 (N_4979,In_755,In_7);
nand U4980 (N_4980,In_830,In_321);
and U4981 (N_4981,In_456,In_223);
or U4982 (N_4982,In_417,In_896);
nor U4983 (N_4983,In_539,In_13);
and U4984 (N_4984,In_75,In_925);
nor U4985 (N_4985,In_45,In_778);
nor U4986 (N_4986,In_698,In_924);
nor U4987 (N_4987,In_880,In_707);
nand U4988 (N_4988,In_16,In_544);
nand U4989 (N_4989,In_513,In_38);
and U4990 (N_4990,In_713,In_676);
and U4991 (N_4991,In_632,In_651);
nand U4992 (N_4992,In_737,In_23);
nand U4993 (N_4993,In_593,In_722);
and U4994 (N_4994,In_543,In_250);
nand U4995 (N_4995,In_533,In_240);
nor U4996 (N_4996,In_34,In_200);
nor U4997 (N_4997,In_1,In_332);
or U4998 (N_4998,In_664,In_747);
and U4999 (N_4999,In_863,In_29);
and U5000 (N_5000,N_1640,N_146);
or U5001 (N_5001,N_128,N_3760);
nand U5002 (N_5002,N_4116,N_2878);
and U5003 (N_5003,N_1219,N_220);
nor U5004 (N_5004,N_2554,N_350);
nand U5005 (N_5005,N_3110,N_4563);
nor U5006 (N_5006,N_145,N_2806);
nor U5007 (N_5007,N_1955,N_4872);
nor U5008 (N_5008,N_939,N_3539);
nand U5009 (N_5009,N_2803,N_3000);
nand U5010 (N_5010,N_4162,N_2312);
or U5011 (N_5011,N_1337,N_742);
and U5012 (N_5012,N_4448,N_2189);
or U5013 (N_5013,N_1517,N_243);
nand U5014 (N_5014,N_2260,N_2275);
and U5015 (N_5015,N_249,N_2195);
nand U5016 (N_5016,N_2429,N_1184);
nor U5017 (N_5017,N_2220,N_6);
or U5018 (N_5018,N_3908,N_2564);
nand U5019 (N_5019,N_4056,N_1697);
nor U5020 (N_5020,N_1606,N_4789);
nor U5021 (N_5021,N_925,N_232);
nand U5022 (N_5022,N_30,N_247);
or U5023 (N_5023,N_4510,N_3642);
nand U5024 (N_5024,N_3520,N_204);
and U5025 (N_5025,N_744,N_4029);
and U5026 (N_5026,N_639,N_3410);
or U5027 (N_5027,N_4986,N_1208);
and U5028 (N_5028,N_942,N_369);
and U5029 (N_5029,N_1406,N_3698);
nor U5030 (N_5030,N_382,N_1186);
nor U5031 (N_5031,N_1178,N_746);
and U5032 (N_5032,N_964,N_4776);
and U5033 (N_5033,N_4750,N_66);
nand U5034 (N_5034,N_3304,N_2744);
nand U5035 (N_5035,N_1297,N_1722);
nor U5036 (N_5036,N_3419,N_4012);
nor U5037 (N_5037,N_4122,N_3483);
nand U5038 (N_5038,N_279,N_2487);
nand U5039 (N_5039,N_426,N_3674);
and U5040 (N_5040,N_1616,N_4764);
and U5041 (N_5041,N_3636,N_3673);
and U5042 (N_5042,N_2194,N_2249);
nor U5043 (N_5043,N_703,N_4920);
and U5044 (N_5044,N_75,N_3852);
nor U5045 (N_5045,N_330,N_4907);
nand U5046 (N_5046,N_2417,N_2048);
nor U5047 (N_5047,N_380,N_4106);
and U5048 (N_5048,N_1596,N_251);
nand U5049 (N_5049,N_3542,N_829);
nand U5050 (N_5050,N_3396,N_3328);
nor U5051 (N_5051,N_1986,N_4609);
or U5052 (N_5052,N_2279,N_4948);
nor U5053 (N_5053,N_2158,N_549);
or U5054 (N_5054,N_4504,N_4385);
or U5055 (N_5055,N_4364,N_3060);
nand U5056 (N_5056,N_3399,N_3693);
xor U5057 (N_5057,N_4273,N_1657);
nand U5058 (N_5058,N_4757,N_4157);
xor U5059 (N_5059,N_4229,N_4585);
or U5060 (N_5060,N_2606,N_3950);
nand U5061 (N_5061,N_739,N_158);
and U5062 (N_5062,N_1272,N_4128);
nor U5063 (N_5063,N_587,N_3042);
or U5064 (N_5064,N_3055,N_2225);
nand U5065 (N_5065,N_4284,N_1529);
and U5066 (N_5066,N_3604,N_1766);
nor U5067 (N_5067,N_3815,N_3059);
nor U5068 (N_5068,N_1637,N_3930);
nor U5069 (N_5069,N_2272,N_2805);
and U5070 (N_5070,N_1591,N_954);
and U5071 (N_5071,N_4174,N_635);
nand U5072 (N_5072,N_2313,N_3474);
xor U5073 (N_5073,N_2122,N_1884);
and U5074 (N_5074,N_608,N_3416);
nand U5075 (N_5075,N_1518,N_4028);
or U5076 (N_5076,N_2435,N_3468);
and U5077 (N_5077,N_525,N_2850);
nand U5078 (N_5078,N_3865,N_2141);
nand U5079 (N_5079,N_556,N_1911);
nand U5080 (N_5080,N_818,N_120);
nor U5081 (N_5081,N_4415,N_837);
nor U5082 (N_5082,N_2540,N_4554);
and U5083 (N_5083,N_1910,N_4857);
or U5084 (N_5084,N_3592,N_1850);
or U5085 (N_5085,N_4537,N_2794);
and U5086 (N_5086,N_4485,N_4319);
and U5087 (N_5087,N_1935,N_1918);
or U5088 (N_5088,N_3885,N_1438);
or U5089 (N_5089,N_4096,N_286);
and U5090 (N_5090,N_3829,N_9);
or U5091 (N_5091,N_1959,N_3555);
and U5092 (N_5092,N_364,N_3402);
and U5093 (N_5093,N_374,N_712);
or U5094 (N_5094,N_3333,N_4092);
and U5095 (N_5095,N_3924,N_4261);
and U5096 (N_5096,N_4299,N_3712);
nand U5097 (N_5097,N_303,N_2368);
xnor U5098 (N_5098,N_2457,N_2625);
xor U5099 (N_5099,N_3945,N_2452);
and U5100 (N_5100,N_116,N_4788);
nor U5101 (N_5101,N_328,N_3692);
nor U5102 (N_5102,N_3314,N_1426);
nand U5103 (N_5103,N_2288,N_891);
nor U5104 (N_5104,N_2533,N_1803);
and U5105 (N_5105,N_1891,N_4940);
and U5106 (N_5106,N_402,N_3046);
nor U5107 (N_5107,N_1909,N_3844);
nand U5108 (N_5108,N_2952,N_1974);
nor U5109 (N_5109,N_2585,N_1994);
and U5110 (N_5110,N_1038,N_4636);
or U5111 (N_5111,N_4339,N_615);
xnor U5112 (N_5112,N_1427,N_2985);
nand U5113 (N_5113,N_1306,N_397);
or U5114 (N_5114,N_2381,N_4369);
nor U5115 (N_5115,N_1201,N_1948);
nand U5116 (N_5116,N_2923,N_4312);
nor U5117 (N_5117,N_2291,N_2180);
or U5118 (N_5118,N_2082,N_2187);
nor U5119 (N_5119,N_470,N_3500);
or U5120 (N_5120,N_606,N_1232);
or U5121 (N_5121,N_4652,N_3647);
nand U5122 (N_5122,N_4432,N_1991);
xnor U5123 (N_5123,N_3373,N_957);
or U5124 (N_5124,N_3864,N_1393);
nand U5125 (N_5125,N_3795,N_2692);
nand U5126 (N_5126,N_1726,N_782);
or U5127 (N_5127,N_4900,N_3188);
or U5128 (N_5128,N_689,N_4275);
or U5129 (N_5129,N_2682,N_179);
nand U5130 (N_5130,N_288,N_1512);
and U5131 (N_5131,N_2034,N_600);
and U5132 (N_5132,N_2166,N_3280);
or U5133 (N_5133,N_2052,N_2406);
and U5134 (N_5134,N_2138,N_616);
and U5135 (N_5135,N_3353,N_1359);
or U5136 (N_5136,N_643,N_1077);
or U5137 (N_5137,N_1624,N_3043);
nor U5138 (N_5138,N_3854,N_1716);
and U5139 (N_5139,N_432,N_3181);
and U5140 (N_5140,N_3031,N_1103);
nor U5141 (N_5141,N_3982,N_3165);
nand U5142 (N_5142,N_992,N_1441);
and U5143 (N_5143,N_3810,N_2454);
nand U5144 (N_5144,N_4131,N_3626);
and U5145 (N_5145,N_301,N_4978);
nor U5146 (N_5146,N_1837,N_2014);
nor U5147 (N_5147,N_3127,N_1746);
nand U5148 (N_5148,N_751,N_3331);
and U5149 (N_5149,N_4457,N_3337);
or U5150 (N_5150,N_353,N_4884);
and U5151 (N_5151,N_4191,N_170);
and U5152 (N_5152,N_1695,N_1318);
and U5153 (N_5153,N_593,N_3501);
nand U5154 (N_5154,N_2185,N_3888);
nand U5155 (N_5155,N_1128,N_2746);
and U5156 (N_5156,N_3870,N_300);
or U5157 (N_5157,N_3853,N_543);
nand U5158 (N_5158,N_846,N_2132);
nand U5159 (N_5159,N_3839,N_2773);
nor U5160 (N_5160,N_2366,N_2290);
nor U5161 (N_5161,N_3797,N_295);
and U5162 (N_5162,N_3837,N_2222);
or U5163 (N_5163,N_2143,N_2458);
and U5164 (N_5164,N_1666,N_2514);
and U5165 (N_5165,N_2476,N_2750);
or U5166 (N_5166,N_1217,N_655);
nand U5167 (N_5167,N_3007,N_1295);
or U5168 (N_5168,N_544,N_3411);
or U5169 (N_5169,N_1634,N_1665);
nand U5170 (N_5170,N_1333,N_4196);
or U5171 (N_5171,N_2899,N_3557);
nor U5172 (N_5172,N_1777,N_4936);
and U5173 (N_5173,N_2025,N_4340);
nand U5174 (N_5174,N_4260,N_2674);
and U5175 (N_5175,N_4151,N_2134);
and U5176 (N_5176,N_119,N_1492);
nand U5177 (N_5177,N_4947,N_2914);
or U5178 (N_5178,N_3472,N_3158);
nor U5179 (N_5179,N_2128,N_2982);
nor U5180 (N_5180,N_2922,N_918);
nand U5181 (N_5181,N_2839,N_3768);
or U5182 (N_5182,N_1002,N_1689);
nand U5183 (N_5183,N_1881,N_1549);
and U5184 (N_5184,N_3351,N_377);
nand U5185 (N_5185,N_4852,N_305);
nand U5186 (N_5186,N_1249,N_4555);
nor U5187 (N_5187,N_1494,N_4835);
or U5188 (N_5188,N_4953,N_1271);
or U5189 (N_5189,N_3040,N_24);
and U5190 (N_5190,N_2653,N_2268);
and U5191 (N_5191,N_1447,N_3841);
nor U5192 (N_5192,N_4368,N_3320);
nand U5193 (N_5193,N_699,N_1207);
and U5194 (N_5194,N_3596,N_2453);
or U5195 (N_5195,N_2154,N_3943);
nand U5196 (N_5196,N_4050,N_510);
nor U5197 (N_5197,N_3808,N_3036);
nand U5198 (N_5198,N_843,N_1875);
and U5199 (N_5199,N_2266,N_3203);
or U5200 (N_5200,N_1888,N_3905);
and U5201 (N_5201,N_2207,N_2135);
nand U5202 (N_5202,N_785,N_2933);
nor U5203 (N_5203,N_1516,N_4800);
or U5204 (N_5204,N_4291,N_1463);
nand U5205 (N_5205,N_317,N_2193);
or U5206 (N_5206,N_80,N_1280);
nor U5207 (N_5207,N_1797,N_2304);
nor U5208 (N_5208,N_4023,N_4316);
or U5209 (N_5209,N_1173,N_696);
and U5210 (N_5210,N_3807,N_2124);
nor U5211 (N_5211,N_4908,N_4198);
nand U5212 (N_5212,N_2282,N_4370);
nor U5213 (N_5213,N_1349,N_4933);
nor U5214 (N_5214,N_3791,N_1138);
nand U5215 (N_5215,N_1469,N_3132);
and U5216 (N_5216,N_2670,N_3567);
or U5217 (N_5217,N_483,N_3817);
or U5218 (N_5218,N_418,N_3428);
or U5219 (N_5219,N_1434,N_3512);
nor U5220 (N_5220,N_4854,N_1324);
nor U5221 (N_5221,N_2103,N_1413);
nand U5222 (N_5222,N_4684,N_4981);
or U5223 (N_5223,N_4803,N_870);
nor U5224 (N_5224,N_3759,N_4889);
nand U5225 (N_5225,N_2832,N_589);
or U5226 (N_5226,N_4696,N_210);
and U5227 (N_5227,N_571,N_3436);
nor U5228 (N_5228,N_2238,N_1776);
nand U5229 (N_5229,N_3183,N_4634);
and U5230 (N_5230,N_2747,N_515);
nand U5231 (N_5231,N_3715,N_786);
nor U5232 (N_5232,N_4726,N_4667);
nand U5233 (N_5233,N_3341,N_2666);
nor U5234 (N_5234,N_1912,N_3359);
nand U5235 (N_5235,N_2668,N_2203);
nor U5236 (N_5236,N_906,N_1056);
or U5237 (N_5237,N_4267,N_2816);
and U5238 (N_5238,N_2937,N_3546);
and U5239 (N_5239,N_1904,N_2579);
nor U5240 (N_5240,N_755,N_4047);
nor U5241 (N_5241,N_564,N_3024);
and U5242 (N_5242,N_4782,N_2562);
nand U5243 (N_5243,N_4780,N_2812);
or U5244 (N_5244,N_729,N_4208);
nor U5245 (N_5245,N_3556,N_3494);
nand U5246 (N_5246,N_4451,N_4120);
and U5247 (N_5247,N_3241,N_3202);
nand U5248 (N_5248,N_2019,N_2449);
nor U5249 (N_5249,N_2801,N_2432);
nand U5250 (N_5250,N_4575,N_434);
and U5251 (N_5251,N_4534,N_3931);
and U5252 (N_5252,N_4613,N_730);
or U5253 (N_5253,N_1083,N_3565);
or U5254 (N_5254,N_2792,N_695);
xor U5255 (N_5255,N_1609,N_1763);
or U5256 (N_5256,N_578,N_4837);
nor U5257 (N_5257,N_2548,N_1036);
and U5258 (N_5258,N_373,N_3834);
or U5259 (N_5259,N_706,N_3107);
nor U5260 (N_5260,N_827,N_2491);
or U5261 (N_5261,N_2863,N_1374);
and U5262 (N_5262,N_3892,N_4519);
or U5263 (N_5263,N_325,N_1230);
nand U5264 (N_5264,N_1668,N_3827);
nor U5265 (N_5265,N_1022,N_3309);
nor U5266 (N_5266,N_2398,N_4293);
or U5267 (N_5267,N_4491,N_1442);
or U5268 (N_5268,N_2797,N_4163);
nor U5269 (N_5269,N_4878,N_2036);
and U5270 (N_5270,N_1385,N_2896);
nor U5271 (N_5271,N_2441,N_1554);
and U5272 (N_5272,N_734,N_4708);
or U5273 (N_5273,N_952,N_3204);
nor U5274 (N_5274,N_1204,N_4905);
and U5275 (N_5275,N_2782,N_3691);
or U5276 (N_5276,N_2500,N_999);
and U5277 (N_5277,N_421,N_3793);
and U5278 (N_5278,N_1711,N_2661);
or U5279 (N_5279,N_1574,N_2261);
nand U5280 (N_5280,N_1021,N_1650);
or U5281 (N_5281,N_140,N_1251);
nor U5282 (N_5282,N_4910,N_4026);
or U5283 (N_5283,N_1432,N_4094);
and U5284 (N_5284,N_661,N_3889);
nor U5285 (N_5285,N_4558,N_2992);
nor U5286 (N_5286,N_1669,N_1395);
nor U5287 (N_5287,N_3992,N_1167);
or U5288 (N_5288,N_3683,N_2496);
nor U5289 (N_5289,N_1636,N_3034);
nand U5290 (N_5290,N_853,N_4975);
or U5291 (N_5291,N_2173,N_29);
and U5292 (N_5292,N_2931,N_2991);
and U5293 (N_5293,N_3401,N_104);
or U5294 (N_5294,N_4333,N_368);
nor U5295 (N_5295,N_2885,N_1563);
nor U5296 (N_5296,N_3968,N_3051);
and U5297 (N_5297,N_4816,N_64);
nand U5298 (N_5298,N_4481,N_2148);
nor U5299 (N_5299,N_799,N_4980);
nor U5300 (N_5300,N_1261,N_816);
and U5301 (N_5301,N_774,N_3851);
nand U5302 (N_5302,N_3763,N_4388);
and U5303 (N_5303,N_4183,N_2145);
or U5304 (N_5304,N_4487,N_1916);
xnor U5305 (N_5305,N_3192,N_1123);
and U5306 (N_5306,N_2883,N_2248);
and U5307 (N_5307,N_264,N_2322);
nand U5308 (N_5308,N_1628,N_4476);
or U5309 (N_5309,N_4209,N_52);
or U5310 (N_5310,N_1028,N_4843);
nor U5311 (N_5311,N_2470,N_2296);
or U5312 (N_5312,N_3171,N_4753);
and U5313 (N_5313,N_3114,N_1445);
nand U5314 (N_5314,N_4620,N_4730);
nor U5315 (N_5315,N_3371,N_248);
nor U5316 (N_5316,N_1949,N_4303);
nor U5317 (N_5317,N_2156,N_3550);
or U5318 (N_5318,N_1625,N_1470);
nand U5319 (N_5319,N_2791,N_768);
or U5320 (N_5320,N_2094,N_2607);
nor U5321 (N_5321,N_4115,N_636);
nor U5322 (N_5322,N_1926,N_1811);
and U5323 (N_5323,N_3228,N_1513);
nand U5324 (N_5324,N_2386,N_3830);
or U5325 (N_5325,N_4436,N_291);
and U5326 (N_5326,N_562,N_2735);
nor U5327 (N_5327,N_848,N_3513);
nor U5328 (N_5328,N_1162,N_4002);
xor U5329 (N_5329,N_4959,N_2512);
or U5330 (N_5330,N_3163,N_1567);
nor U5331 (N_5331,N_1176,N_561);
and U5332 (N_5332,N_2888,N_2117);
or U5333 (N_5333,N_10,N_2849);
and U5334 (N_5334,N_1125,N_4187);
nand U5335 (N_5335,N_3508,N_1188);
nand U5336 (N_5336,N_2732,N_1964);
or U5337 (N_5337,N_1132,N_3243);
and U5338 (N_5338,N_1807,N_3291);
xnor U5339 (N_5339,N_4499,N_3142);
nor U5340 (N_5340,N_4665,N_3744);
nor U5341 (N_5341,N_4527,N_117);
nor U5342 (N_5342,N_919,N_3986);
and U5343 (N_5343,N_1962,N_4969);
nor U5344 (N_5344,N_2826,N_3824);
nand U5345 (N_5345,N_2324,N_235);
nand U5346 (N_5346,N_4346,N_166);
nand U5347 (N_5347,N_3754,N_2544);
nor U5348 (N_5348,N_3521,N_2058);
or U5349 (N_5349,N_1541,N_4016);
or U5350 (N_5350,N_3719,N_1623);
nor U5351 (N_5351,N_4606,N_4917);
or U5352 (N_5352,N_4896,N_4706);
nor U5353 (N_5353,N_4222,N_3794);
nand U5354 (N_5354,N_218,N_1061);
nor U5355 (N_5355,N_2936,N_1285);
nor U5356 (N_5356,N_2032,N_3082);
nand U5357 (N_5357,N_4605,N_1829);
and U5358 (N_5358,N_1199,N_1845);
or U5359 (N_5359,N_1124,N_4348);
nor U5360 (N_5360,N_2935,N_4158);
nor U5361 (N_5361,N_3682,N_4895);
nand U5362 (N_5362,N_1989,N_2785);
xor U5363 (N_5363,N_3433,N_4366);
or U5364 (N_5364,N_1013,N_4722);
or U5365 (N_5365,N_3456,N_152);
and U5366 (N_5366,N_93,N_1334);
and U5367 (N_5367,N_792,N_2259);
or U5368 (N_5368,N_4089,N_1448);
nor U5369 (N_5369,N_4983,N_717);
nand U5370 (N_5370,N_1145,N_728);
or U5371 (N_5371,N_590,N_3222);
or U5372 (N_5372,N_73,N_4614);
nor U5373 (N_5373,N_663,N_3654);
or U5374 (N_5374,N_956,N_2305);
nand U5375 (N_5375,N_1709,N_4205);
or U5376 (N_5376,N_3767,N_1611);
or U5377 (N_5377,N_3926,N_3927);
and U5378 (N_5378,N_2077,N_1154);
and U5379 (N_5379,N_1381,N_49);
xnor U5380 (N_5380,N_3452,N_314);
nor U5381 (N_5381,N_3562,N_1235);
or U5382 (N_5382,N_2742,N_2486);
and U5383 (N_5383,N_3305,N_2258);
and U5384 (N_5384,N_0,N_2426);
nand U5385 (N_5385,N_390,N_877);
nor U5386 (N_5386,N_1630,N_4919);
or U5387 (N_5387,N_1992,N_3193);
nand U5388 (N_5388,N_1229,N_2781);
nand U5389 (N_5389,N_1403,N_4008);
or U5390 (N_5390,N_1377,N_784);
nor U5391 (N_5391,N_403,N_3529);
or U5392 (N_5392,N_4773,N_3545);
or U5393 (N_5393,N_2106,N_4700);
and U5394 (N_5394,N_3783,N_1894);
or U5395 (N_5395,N_4309,N_1198);
or U5396 (N_5396,N_3593,N_277);
nor U5397 (N_5397,N_4140,N_359);
or U5398 (N_5398,N_4195,N_1929);
nand U5399 (N_5399,N_2861,N_2722);
nand U5400 (N_5400,N_2752,N_2054);
and U5401 (N_5401,N_2617,N_4044);
nor U5402 (N_5402,N_1211,N_4215);
and U5403 (N_5403,N_1238,N_1704);
or U5404 (N_5404,N_1967,N_3573);
nand U5405 (N_5405,N_1906,N_261);
and U5406 (N_5406,N_1840,N_4898);
and U5407 (N_5407,N_3750,N_4608);
or U5408 (N_5408,N_4,N_962);
or U5409 (N_5409,N_1220,N_1528);
and U5410 (N_5410,N_3713,N_3965);
and U5411 (N_5411,N_982,N_3083);
and U5412 (N_5412,N_1237,N_2619);
or U5413 (N_5413,N_4150,N_160);
and U5414 (N_5414,N_4815,N_4517);
nand U5415 (N_5415,N_1582,N_153);
nand U5416 (N_5416,N_4313,N_4714);
nand U5417 (N_5417,N_4244,N_1682);
or U5418 (N_5418,N_1804,N_3875);
and U5419 (N_5419,N_3015,N_2380);
and U5420 (N_5420,N_775,N_1375);
nor U5421 (N_5421,N_1350,N_3677);
nor U5422 (N_5422,N_685,N_3112);
nor U5423 (N_5423,N_3105,N_3216);
nor U5424 (N_5424,N_4077,N_921);
nand U5425 (N_5425,N_1555,N_1);
nor U5426 (N_5426,N_1118,N_3258);
and U5427 (N_5427,N_2421,N_4173);
and U5428 (N_5428,N_21,N_4683);
and U5429 (N_5429,N_2358,N_896);
nand U5430 (N_5430,N_2690,N_726);
nor U5431 (N_5431,N_271,N_137);
or U5432 (N_5432,N_239,N_3669);
nor U5433 (N_5433,N_4220,N_4972);
nor U5434 (N_5434,N_1101,N_3847);
and U5435 (N_5435,N_2916,N_3524);
nor U5436 (N_5436,N_2565,N_1093);
or U5437 (N_5437,N_3278,N_3354);
and U5438 (N_5438,N_3030,N_1605);
or U5439 (N_5439,N_1717,N_4795);
and U5440 (N_5440,N_3421,N_1143);
nor U5441 (N_5441,N_2188,N_3798);
nor U5442 (N_5442,N_1033,N_1519);
or U5443 (N_5443,N_3357,N_3497);
nor U5444 (N_5444,N_28,N_842);
nor U5445 (N_5445,N_594,N_3028);
and U5446 (N_5446,N_3492,N_1245);
nand U5447 (N_5447,N_1340,N_3260);
and U5448 (N_5448,N_1079,N_4814);
xnor U5449 (N_5449,N_2957,N_1065);
nor U5450 (N_5450,N_1137,N_3406);
or U5451 (N_5451,N_3242,N_2969);
nor U5452 (N_5452,N_1740,N_1558);
and U5453 (N_5453,N_1155,N_161);
and U5454 (N_5454,N_1082,N_4631);
and U5455 (N_5455,N_1643,N_614);
nand U5456 (N_5456,N_4456,N_4724);
or U5457 (N_5457,N_3516,N_4860);
nand U5458 (N_5458,N_3934,N_121);
and U5459 (N_5459,N_3932,N_1767);
or U5460 (N_5460,N_1015,N_715);
or U5461 (N_5461,N_721,N_3417);
nor U5462 (N_5462,N_3611,N_3686);
nand U5463 (N_5463,N_1299,N_1116);
and U5464 (N_5464,N_3504,N_1510);
or U5465 (N_5465,N_159,N_1312);
and U5466 (N_5466,N_3728,N_3054);
nor U5467 (N_5467,N_931,N_2308);
or U5468 (N_5468,N_2780,N_3473);
nand U5469 (N_5469,N_1747,N_2778);
and U5470 (N_5470,N_312,N_2497);
nand U5471 (N_5471,N_3448,N_3369);
nand U5472 (N_5472,N_4253,N_2851);
nand U5473 (N_5473,N_2505,N_4167);
xor U5474 (N_5474,N_2168,N_1760);
and U5475 (N_5475,N_3469,N_4719);
or U5476 (N_5476,N_2981,N_406);
and U5477 (N_5477,N_122,N_499);
and U5478 (N_5478,N_3887,N_4955);
nor U5479 (N_5479,N_444,N_1836);
nand U5480 (N_5480,N_2416,N_495);
nor U5481 (N_5481,N_3200,N_4286);
or U5482 (N_5482,N_4587,N_1346);
nor U5483 (N_5483,N_1044,N_4512);
or U5484 (N_5484,N_3381,N_2162);
nor U5485 (N_5485,N_4574,N_2798);
and U5486 (N_5486,N_3130,N_2960);
nand U5487 (N_5487,N_1936,N_758);
and U5488 (N_5488,N_3496,N_221);
and U5489 (N_5489,N_1957,N_1857);
and U5490 (N_5490,N_3577,N_2893);
nor U5491 (N_5491,N_2196,N_1687);
nor U5492 (N_5492,N_334,N_4088);
nor U5493 (N_5493,N_1322,N_1503);
nand U5494 (N_5494,N_793,N_1886);
or U5495 (N_5495,N_4859,N_4105);
nor U5496 (N_5496,N_1421,N_4741);
and U5497 (N_5497,N_50,N_3058);
xor U5498 (N_5498,N_1815,N_3063);
or U5499 (N_5499,N_255,N_3144);
nor U5500 (N_5500,N_4746,N_551);
or U5501 (N_5501,N_167,N_724);
nand U5502 (N_5502,N_1810,N_1331);
and U5503 (N_5503,N_1043,N_4772);
nor U5504 (N_5504,N_1006,N_2285);
nor U5505 (N_5505,N_4202,N_1095);
nand U5506 (N_5506,N_1855,N_3338);
nand U5507 (N_5507,N_1693,N_1556);
and U5508 (N_5508,N_1452,N_1943);
xor U5509 (N_5509,N_1169,N_1831);
nand U5510 (N_5510,N_878,N_2270);
or U5511 (N_5511,N_823,N_7);
nor U5512 (N_5512,N_4152,N_1997);
nor U5513 (N_5513,N_1025,N_1371);
nand U5514 (N_5514,N_1805,N_4014);
or U5515 (N_5515,N_4822,N_3967);
nand U5516 (N_5516,N_3498,N_1203);
xor U5517 (N_5517,N_3566,N_2995);
and U5518 (N_5518,N_253,N_4149);
xnor U5519 (N_5519,N_3928,N_855);
nor U5520 (N_5520,N_1878,N_1287);
or U5521 (N_5521,N_2295,N_3092);
xnor U5522 (N_5522,N_3326,N_3684);
or U5523 (N_5523,N_773,N_1243);
and U5524 (N_5524,N_2367,N_4289);
or U5525 (N_5525,N_2253,N_1047);
and U5526 (N_5526,N_642,N_798);
and U5527 (N_5527,N_3788,N_1304);
and U5528 (N_5528,N_297,N_2382);
or U5529 (N_5529,N_1790,N_4989);
or U5530 (N_5530,N_2498,N_1086);
or U5531 (N_5531,N_3601,N_3707);
and U5532 (N_5532,N_4767,N_4324);
nand U5533 (N_5533,N_1182,N_3286);
or U5534 (N_5534,N_4074,N_2028);
nor U5535 (N_5535,N_361,N_2144);
nand U5536 (N_5536,N_2623,N_693);
and U5537 (N_5537,N_2315,N_960);
or U5538 (N_5538,N_1507,N_1417);
nand U5539 (N_5539,N_4707,N_3118);
and U5540 (N_5540,N_3245,N_33);
nor U5541 (N_5541,N_4839,N_2405);
and U5542 (N_5542,N_836,N_196);
and U5543 (N_5543,N_1876,N_2838);
nand U5544 (N_5544,N_4123,N_4136);
nand U5545 (N_5545,N_1999,N_948);
and U5546 (N_5546,N_584,N_3145);
and U5547 (N_5547,N_4783,N_4305);
and U5548 (N_5548,N_3348,N_518);
nor U5549 (N_5549,N_1728,N_2963);
nand U5550 (N_5550,N_4892,N_4793);
and U5551 (N_5551,N_2242,N_4893);
and U5552 (N_5552,N_519,N_1401);
nor U5553 (N_5553,N_4721,N_3288);
nor U5554 (N_5554,N_4490,N_3336);
and U5555 (N_5555,N_4740,N_565);
or U5556 (N_5556,N_3025,N_1565);
or U5557 (N_5557,N_607,N_478);
and U5558 (N_5558,N_3656,N_1681);
nand U5559 (N_5559,N_2273,N_1193);
or U5560 (N_5560,N_3460,N_3041);
nand U5561 (N_5561,N_1172,N_2684);
nor U5562 (N_5562,N_4559,N_3388);
xnor U5563 (N_5563,N_4625,N_1465);
nor U5564 (N_5564,N_1054,N_1260);
nor U5565 (N_5565,N_1920,N_2719);
and U5566 (N_5566,N_4035,N_1802);
nor U5567 (N_5567,N_4671,N_1122);
nand U5568 (N_5568,N_2113,N_2518);
and U5569 (N_5569,N_4207,N_2827);
nor U5570 (N_5570,N_3901,N_3776);
and U5571 (N_5571,N_44,N_835);
nor U5572 (N_5572,N_4292,N_3717);
or U5573 (N_5573,N_4240,N_3450);
or U5574 (N_5574,N_3721,N_2484);
or U5575 (N_5575,N_2858,N_828);
and U5576 (N_5576,N_388,N_3973);
and U5577 (N_5577,N_3451,N_4154);
or U5578 (N_5578,N_4902,N_3762);
nor U5579 (N_5579,N_2450,N_3599);
or U5580 (N_5580,N_3720,N_2064);
nand U5581 (N_5581,N_487,N_4343);
nand U5582 (N_5582,N_1097,N_2121);
and U5583 (N_5583,N_1638,N_103);
nor U5584 (N_5584,N_2672,N_2639);
nor U5585 (N_5585,N_2964,N_2620);
and U5586 (N_5586,N_201,N_1576);
nand U5587 (N_5587,N_36,N_3509);
nor U5588 (N_5588,N_3660,N_2934);
or U5589 (N_5589,N_1607,N_4318);
nor U5590 (N_5590,N_4025,N_4111);
nor U5591 (N_5591,N_4580,N_4622);
and U5592 (N_5592,N_4471,N_4429);
or U5593 (N_5593,N_2955,N_2609);
and U5594 (N_5594,N_1862,N_3948);
or U5595 (N_5595,N_4544,N_2241);
nand U5596 (N_5596,N_4751,N_1091);
and U5597 (N_5597,N_946,N_3458);
or U5598 (N_5598,N_157,N_479);
or U5599 (N_5599,N_3553,N_4478);
and U5600 (N_5600,N_238,N_1161);
nor U5601 (N_5601,N_2940,N_461);
and U5602 (N_5602,N_3072,N_1965);
nor U5603 (N_5603,N_2181,N_3963);
and U5604 (N_5604,N_4934,N_2882);
or U5605 (N_5605,N_2503,N_77);
nor U5606 (N_5606,N_2634,N_4396);
or U5607 (N_5607,N_2996,N_338);
nor U5608 (N_5608,N_3462,N_3659);
and U5609 (N_5609,N_4530,N_183);
or U5610 (N_5610,N_3734,N_2769);
or U5611 (N_5611,N_1969,N_343);
or U5612 (N_5612,N_4932,N_3666);
nor U5613 (N_5613,N_2599,N_1451);
nor U5614 (N_5614,N_4359,N_191);
and U5615 (N_5615,N_1425,N_538);
or U5616 (N_5616,N_1646,N_2578);
nand U5617 (N_5617,N_2559,N_1476);
or U5618 (N_5618,N_492,N_512);
nand U5619 (N_5619,N_735,N_4830);
nor U5620 (N_5620,N_4626,N_3733);
nor U5621 (N_5621,N_4093,N_1156);
nor U5622 (N_5622,N_407,N_4915);
and U5623 (N_5623,N_1303,N_4469);
xnor U5624 (N_5624,N_2651,N_2618);
nor U5625 (N_5625,N_1511,N_4124);
or U5626 (N_5626,N_209,N_839);
or U5627 (N_5627,N_355,N_4015);
nand U5628 (N_5628,N_4669,N_454);
nand U5629 (N_5629,N_3879,N_3989);
or U5630 (N_5630,N_2243,N_2294);
or U5631 (N_5631,N_4916,N_2705);
and U5632 (N_5632,N_3343,N_3340);
or U5633 (N_5633,N_443,N_1360);
nor U5634 (N_5634,N_2569,N_4629);
nand U5635 (N_5635,N_1615,N_3330);
nand U5636 (N_5636,N_951,N_3137);
nor U5637 (N_5637,N_4062,N_4141);
and U5638 (N_5638,N_342,N_2212);
nor U5639 (N_5639,N_1357,N_4495);
nor U5640 (N_5640,N_4545,N_4754);
nand U5641 (N_5641,N_3597,N_1200);
or U5642 (N_5642,N_2303,N_3871);
nand U5643 (N_5643,N_3860,N_2638);
and U5644 (N_5644,N_4646,N_1983);
and U5645 (N_5645,N_2921,N_1244);
xnor U5646 (N_5646,N_873,N_2023);
nor U5647 (N_5647,N_4688,N_2474);
nor U5648 (N_5648,N_1799,N_4247);
and U5649 (N_5649,N_4786,N_2235);
nor U5650 (N_5650,N_2737,N_4617);
and U5651 (N_5651,N_1764,N_453);
nand U5652 (N_5652,N_1119,N_2502);
nor U5653 (N_5653,N_3971,N_759);
or U5654 (N_5654,N_1163,N_2986);
nor U5655 (N_5655,N_1754,N_427);
nor U5656 (N_5656,N_4738,N_4112);
nor U5657 (N_5657,N_1945,N_3709);
nand U5658 (N_5658,N_4410,N_3894);
or U5659 (N_5659,N_195,N_3268);
nor U5660 (N_5660,N_4586,N_1135);
or U5661 (N_5661,N_2528,N_612);
and U5662 (N_5662,N_4524,N_2464);
nor U5663 (N_5663,N_3855,N_2396);
nor U5664 (N_5664,N_3502,N_2971);
nand U5665 (N_5665,N_1464,N_3748);
nor U5666 (N_5666,N_4287,N_2384);
nand U5667 (N_5667,N_2257,N_2099);
or U5668 (N_5668,N_129,N_3261);
and U5669 (N_5669,N_4984,N_4645);
and U5670 (N_5670,N_2111,N_4996);
nor U5671 (N_5671,N_1004,N_4618);
nor U5672 (N_5672,N_973,N_1917);
and U5673 (N_5673,N_2706,N_2631);
nor U5674 (N_5674,N_1487,N_2233);
or U5675 (N_5675,N_3212,N_3979);
nor U5676 (N_5676,N_1688,N_3857);
and U5677 (N_5677,N_3676,N_4223);
nor U5678 (N_5678,N_1859,N_90);
nor U5679 (N_5679,N_4901,N_852);
or U5680 (N_5680,N_1699,N_3446);
and U5681 (N_5681,N_967,N_4566);
nor U5682 (N_5682,N_3561,N_3065);
or U5683 (N_5683,N_2643,N_130);
nor U5684 (N_5684,N_2646,N_3897);
or U5685 (N_5685,N_1861,N_4295);
or U5686 (N_5686,N_1900,N_4551);
nand U5687 (N_5687,N_1809,N_2881);
nor U5688 (N_5688,N_601,N_4774);
or U5689 (N_5689,N_3704,N_3047);
nand U5690 (N_5690,N_4570,N_4051);
nand U5691 (N_5691,N_895,N_16);
or U5692 (N_5692,N_3878,N_1808);
nand U5693 (N_5693,N_391,N_3075);
nor U5694 (N_5694,N_1592,N_4245);
or U5695 (N_5695,N_3303,N_2447);
or U5696 (N_5696,N_226,N_1813);
or U5697 (N_5697,N_3662,N_2563);
nand U5698 (N_5698,N_599,N_2817);
or U5699 (N_5699,N_3426,N_2566);
or U5700 (N_5700,N_679,N_4562);
and U5701 (N_5701,N_207,N_4169);
and U5702 (N_5702,N_452,N_1256);
xor U5703 (N_5703,N_4756,N_3681);
nand U5704 (N_5704,N_1680,N_2570);
or U5705 (N_5705,N_4164,N_1825);
nand U5706 (N_5706,N_3429,N_3978);
and U5707 (N_5707,N_2349,N_3646);
and U5708 (N_5708,N_13,N_2151);
nand U5709 (N_5709,N_4423,N_4897);
and U5710 (N_5710,N_3861,N_2833);
nand U5711 (N_5711,N_3032,N_4031);
nand U5712 (N_5712,N_2657,N_526);
and U5713 (N_5713,N_4572,N_1062);
nand U5714 (N_5714,N_4698,N_2069);
or U5715 (N_5715,N_945,N_4383);
and U5716 (N_5716,N_3162,N_731);
nand U5717 (N_5717,N_1950,N_4326);
or U5718 (N_5718,N_420,N_3455);
nor U5719 (N_5719,N_854,N_1436);
xnor U5720 (N_5720,N_4496,N_4994);
nand U5721 (N_5721,N_3444,N_4848);
and U5722 (N_5722,N_4075,N_974);
nand U5723 (N_5723,N_3481,N_3439);
nor U5724 (N_5724,N_2445,N_888);
and U5725 (N_5725,N_67,N_988);
nor U5726 (N_5726,N_2820,N_4594);
nor U5727 (N_5727,N_4118,N_3802);
nor U5728 (N_5728,N_2845,N_3335);
and U5729 (N_5729,N_178,N_629);
or U5730 (N_5730,N_3061,N_51);
or U5731 (N_5731,N_874,N_4732);
or U5732 (N_5732,N_4479,N_3705);
nor U5733 (N_5733,N_3170,N_926);
nor U5734 (N_5734,N_4143,N_3651);
nor U5735 (N_5735,N_2192,N_63);
and U5736 (N_5736,N_4590,N_4763);
or U5737 (N_5737,N_177,N_1573);
nor U5738 (N_5738,N_638,N_348);
and U5739 (N_5739,N_4599,N_3006);
nor U5740 (N_5740,N_3738,N_4148);
or U5741 (N_5741,N_501,N_841);
or U5742 (N_5742,N_4068,N_4061);
nand U5743 (N_5743,N_560,N_2354);
nor U5744 (N_5744,N_4040,N_3459);
and U5745 (N_5745,N_4294,N_3069);
and U5746 (N_5746,N_3194,N_282);
and U5747 (N_5747,N_4812,N_2856);
or U5748 (N_5748,N_2091,N_3441);
nor U5749 (N_5749,N_644,N_4017);
and U5750 (N_5750,N_3537,N_2244);
and U5751 (N_5751,N_2541,N_4670);
nor U5752 (N_5752,N_778,N_2240);
or U5753 (N_5753,N_4034,N_3972);
nand U5754 (N_5754,N_1262,N_3607);
xnor U5755 (N_5755,N_212,N_4828);
and U5756 (N_5756,N_2030,N_634);
and U5757 (N_5757,N_278,N_4553);
or U5758 (N_5758,N_4883,N_4099);
nand U5759 (N_5759,N_4921,N_2515);
and U5760 (N_5760,N_2768,N_4644);
or U5761 (N_5761,N_1654,N_3687);
and U5762 (N_5762,N_3695,N_345);
and U5763 (N_5763,N_3758,N_1586);
nor U5764 (N_5764,N_805,N_4729);
or U5765 (N_5765,N_4227,N_3745);
or U5766 (N_5766,N_3856,N_2049);
or U5767 (N_5767,N_3347,N_1338);
nor U5768 (N_5768,N_3833,N_3322);
or U5769 (N_5769,N_1085,N_2112);
or U5770 (N_5770,N_4418,N_3638);
or U5771 (N_5771,N_1387,N_4693);
nor U5772 (N_5772,N_4421,N_4825);
nor U5773 (N_5773,N_2688,N_3874);
nor U5774 (N_5774,N_163,N_96);
and U5775 (N_5775,N_3655,N_2412);
nand U5776 (N_5776,N_3832,N_415);
or U5777 (N_5777,N_4990,N_4045);
or U5778 (N_5778,N_1410,N_318);
nand U5779 (N_5779,N_3189,N_3003);
nand U5780 (N_5780,N_2539,N_2234);
or U5781 (N_5781,N_1035,N_4443);
or U5782 (N_5782,N_1493,N_3177);
and U5783 (N_5783,N_4069,N_2376);
nand U5784 (N_5784,N_240,N_3828);
and U5785 (N_5785,N_2088,N_412);
and U5786 (N_5786,N_1788,N_4713);
nand U5787 (N_5787,N_1415,N_1474);
nand U5788 (N_5788,N_4360,N_1736);
and U5789 (N_5789,N_4095,N_1618);
xnor U5790 (N_5790,N_745,N_3530);
nor U5791 (N_5791,N_3398,N_1212);
and U5792 (N_5792,N_4962,N_3774);
and U5793 (N_5793,N_3120,N_20);
nor U5794 (N_5794,N_339,N_3997);
nor U5795 (N_5795,N_4781,N_2865);
nand U5796 (N_5796,N_1252,N_4356);
nor U5797 (N_5797,N_809,N_2205);
or U5798 (N_5798,N_770,N_417);
nor U5799 (N_5799,N_3723,N_912);
nor U5800 (N_5800,N_1267,N_1501);
or U5801 (N_5801,N_4649,N_4219);
nand U5802 (N_5802,N_1622,N_2824);
nor U5803 (N_5803,N_1914,N_3121);
or U5804 (N_5804,N_1944,N_4257);
and U5805 (N_5805,N_42,N_1651);
and U5806 (N_5806,N_1265,N_574);
and U5807 (N_5807,N_1771,N_1405);
xnor U5808 (N_5808,N_1941,N_687);
and U5809 (N_5809,N_2841,N_4965);
nor U5810 (N_5810,N_4805,N_2492);
or U5811 (N_5811,N_1189,N_2869);
nor U5812 (N_5812,N_4283,N_1844);
and U5813 (N_5813,N_802,N_112);
nor U5814 (N_5814,N_4864,N_2075);
and U5815 (N_5815,N_1956,N_3476);
nor U5816 (N_5816,N_1461,N_2387);
nand U5817 (N_5817,N_1205,N_168);
or U5818 (N_5818,N_3190,N_4941);
or U5819 (N_5819,N_4458,N_4172);
or U5820 (N_5820,N_329,N_2825);
or U5821 (N_5821,N_711,N_1223);
nor U5822 (N_5822,N_3275,N_424);
or U5823 (N_5823,N_4498,N_371);
or U5824 (N_5824,N_4778,N_26);
nand U5825 (N_5825,N_3346,N_2905);
nand U5826 (N_5826,N_1003,N_1437);
and U5827 (N_5827,N_2602,N_1462);
and U5828 (N_5828,N_2748,N_111);
or U5829 (N_5829,N_3749,N_3299);
or U5830 (N_5830,N_2409,N_3868);
or U5831 (N_5831,N_3420,N_575);
or U5832 (N_5832,N_4600,N_581);
nor U5833 (N_5833,N_620,N_3284);
and U5834 (N_5834,N_4998,N_4577);
or U5835 (N_5835,N_3215,N_1848);
and U5836 (N_5836,N_2531,N_1010);
or U5837 (N_5837,N_4914,N_2912);
or U5838 (N_5838,N_1885,N_514);
and U5839 (N_5839,N_1671,N_3307);
and U5840 (N_5840,N_1537,N_2636);
or U5841 (N_5841,N_4001,N_1031);
nand U5842 (N_5842,N_2604,N_1535);
nor U5843 (N_5843,N_413,N_933);
nand U5844 (N_5844,N_4301,N_1782);
nand U5845 (N_5845,N_3285,N_419);
nand U5846 (N_5846,N_708,N_2456);
nor U5847 (N_5847,N_4052,N_684);
and U5848 (N_5848,N_3106,N_4796);
nor U5849 (N_5849,N_2808,N_1344);
and U5850 (N_5850,N_3453,N_1632);
nor U5851 (N_5851,N_1433,N_736);
nor U5852 (N_5852,N_3334,N_1181);
or U5853 (N_5853,N_686,N_4386);
nor U5854 (N_5854,N_767,N_4616);
nand U5855 (N_5855,N_2802,N_851);
and U5856 (N_5856,N_4281,N_2632);
nand U5857 (N_5857,N_1847,N_4657);
nand U5858 (N_5858,N_3534,N_3631);
and U5859 (N_5859,N_134,N_1034);
xor U5860 (N_5860,N_882,N_475);
nand U5861 (N_5861,N_4720,N_617);
or U5862 (N_5862,N_4565,N_1473);
nand U5863 (N_5863,N_1739,N_394);
nor U5864 (N_5864,N_85,N_4258);
and U5865 (N_5865,N_4004,N_2420);
nor U5866 (N_5866,N_2199,N_4484);
and U5867 (N_5867,N_3391,N_4107);
or U5868 (N_5868,N_306,N_825);
nand U5869 (N_5869,N_1793,N_3540);
or U5870 (N_5870,N_4020,N_2932);
and U5871 (N_5871,N_3167,N_1833);
nand U5872 (N_5872,N_516,N_2810);
nor U5873 (N_5873,N_4447,N_1399);
nand U5874 (N_5874,N_4951,N_1250);
or U5875 (N_5875,N_1278,N_4547);
and U5876 (N_5876,N_3168,N_3914);
and U5877 (N_5877,N_1014,N_4166);
nand U5878 (N_5878,N_1849,N_2415);
or U5879 (N_5879,N_2866,N_3404);
and U5880 (N_5880,N_344,N_4426);
and U5881 (N_5881,N_2391,N_2090);
nand U5882 (N_5882,N_2504,N_3154);
nand U5883 (N_5883,N_3777,N_4523);
or U5884 (N_5884,N_2925,N_4702);
and U5885 (N_5885,N_972,N_349);
and U5886 (N_5886,N_1869,N_1477);
nor U5887 (N_5887,N_3780,N_3050);
nand U5888 (N_5888,N_2211,N_2645);
and U5889 (N_5889,N_31,N_1026);
nor U5890 (N_5890,N_779,N_2321);
xnor U5891 (N_5891,N_3029,N_2274);
and U5892 (N_5892,N_4540,N_2362);
and U5893 (N_5893,N_3226,N_2341);
nor U5894 (N_5894,N_4881,N_2283);
nor U5895 (N_5895,N_1332,N_1055);
nand U5896 (N_5896,N_3872,N_1481);
nand U5897 (N_5897,N_2125,N_1577);
and U5898 (N_5898,N_559,N_4063);
and U5899 (N_5899,N_1675,N_3765);
nor U5900 (N_5900,N_2494,N_2718);
or U5901 (N_5901,N_3045,N_553);
nand U5902 (N_5902,N_1099,N_602);
and U5903 (N_5903,N_4627,N_845);
nand U5904 (N_5904,N_274,N_1500);
or U5905 (N_5905,N_1164,N_626);
nand U5906 (N_5906,N_1553,N_472);
and U5907 (N_5907,N_3838,N_169);
nor U5908 (N_5908,N_1694,N_2961);
nand U5909 (N_5909,N_401,N_4849);
and U5910 (N_5910,N_4372,N_3093);
nand U5911 (N_5911,N_3023,N_4465);
nand U5912 (N_5912,N_4909,N_2667);
nor U5913 (N_5913,N_3998,N_2217);
or U5914 (N_5914,N_1744,N_1613);
or U5915 (N_5915,N_2901,N_4091);
or U5916 (N_5916,N_4794,N_3663);
and U5917 (N_5917,N_4979,N_3119);
and U5918 (N_5918,N_3801,N_2068);
nand U5919 (N_5919,N_1735,N_180);
nor U5920 (N_5920,N_2730,N_2898);
nor U5921 (N_5921,N_2938,N_2576);
or U5922 (N_5922,N_4146,N_3942);
or U5923 (N_5923,N_3994,N_4134);
and U5924 (N_5924,N_1731,N_3806);
nand U5925 (N_5925,N_3690,N_807);
or U5926 (N_5926,N_4704,N_3937);
or U5927 (N_5927,N_2483,N_2332);
xnor U5928 (N_5928,N_3511,N_4344);
and U5929 (N_5929,N_4231,N_3150);
or U5930 (N_5930,N_3716,N_336);
nand U5931 (N_5931,N_995,N_2948);
or U5932 (N_5932,N_1227,N_2093);
nor U5933 (N_5933,N_1366,N_2834);
nand U5934 (N_5934,N_4121,N_3688);
nor U5935 (N_5935,N_4176,N_1288);
or U5936 (N_5936,N_772,N_4435);
nand U5937 (N_5937,N_1515,N_771);
nand U5938 (N_5938,N_1981,N_4761);
nor U5939 (N_5939,N_302,N_3174);
and U5940 (N_5940,N_3408,N_4230);
nor U5941 (N_5941,N_1491,N_2300);
or U5942 (N_5942,N_3447,N_2286);
and U5943 (N_5943,N_704,N_4755);
or U5944 (N_5944,N_2926,N_241);
nor U5945 (N_5945,N_4779,N_1206);
nand U5946 (N_5946,N_4968,N_1631);
nand U5947 (N_5947,N_3980,N_262);
xor U5948 (N_5948,N_692,N_1583);
and U5949 (N_5949,N_1599,N_4856);
or U5950 (N_5950,N_1789,N_3378);
nor U5951 (N_5951,N_4699,N_4906);
or U5952 (N_5952,N_1961,N_2377);
nor U5953 (N_5953,N_4453,N_2943);
nor U5954 (N_5954,N_3172,N_4952);
nand U5955 (N_5955,N_3915,N_867);
or U5956 (N_5956,N_4826,N_4681);
and U5957 (N_5957,N_1547,N_2105);
or U5958 (N_5958,N_1765,N_1953);
nor U5959 (N_5959,N_1185,N_1274);
nor U5960 (N_5960,N_2226,N_1755);
nand U5961 (N_5961,N_3849,N_2717);
nand U5962 (N_5962,N_2408,N_491);
and U5963 (N_5963,N_1472,N_1670);
and U5964 (N_5964,N_4337,N_2092);
xor U5965 (N_5965,N_3615,N_1676);
or U5966 (N_5966,N_154,N_2959);
or U5967 (N_5967,N_1702,N_1738);
nor U5968 (N_5968,N_856,N_670);
nor U5969 (N_5969,N_3954,N_1192);
or U5970 (N_5970,N_2340,N_879);
nor U5971 (N_5971,N_8,N_1987);
nor U5972 (N_5972,N_4422,N_3570);
nor U5973 (N_5973,N_1977,N_2201);
nor U5974 (N_5974,N_801,N_688);
or U5975 (N_5975,N_1335,N_3831);
and U5976 (N_5976,N_1690,N_3185);
nand U5977 (N_5977,N_4821,N_3311);
nor U5978 (N_5978,N_4887,N_780);
and U5979 (N_5979,N_2840,N_3867);
and U5980 (N_5980,N_4705,N_2095);
and U5981 (N_5981,N_976,N_4725);
nand U5982 (N_5982,N_3766,N_1701);
nor U5983 (N_5983,N_1009,N_3591);
or U5984 (N_5984,N_1614,N_2459);
nand U5985 (N_5985,N_1783,N_2998);
nand U5986 (N_5986,N_1696,N_2997);
and U5987 (N_5987,N_2284,N_4018);
or U5988 (N_5988,N_2689,N_3641);
and U5989 (N_5989,N_217,N_3694);
nor U5990 (N_5990,N_2271,N_3859);
and U5991 (N_5991,N_4407,N_1550);
nand U5992 (N_5992,N_2814,N_1496);
and U5993 (N_5993,N_3151,N_2764);
or U5994 (N_5994,N_465,N_4467);
nand U5995 (N_5995,N_1450,N_2879);
and U5996 (N_5996,N_1588,N_4065);
or U5997 (N_5997,N_1115,N_4880);
nor U5998 (N_5998,N_2507,N_2110);
nand U5999 (N_5999,N_654,N_254);
and U6000 (N_6000,N_4885,N_449);
nand U6001 (N_6001,N_1170,N_1525);
or U6002 (N_6002,N_1960,N_3836);
xor U6003 (N_6003,N_497,N_1449);
or U6004 (N_6004,N_3974,N_1913);
nand U6005 (N_6005,N_716,N_2100);
nand U6006 (N_6006,N_901,N_2076);
xnor U6007 (N_6007,N_4375,N_2329);
nor U6008 (N_6008,N_3770,N_1264);
or U6009 (N_6009,N_2685,N_392);
nand U6010 (N_6010,N_628,N_585);
nor U6011 (N_6011,N_188,N_4027);
nor U6012 (N_6012,N_2221,N_4811);
nand U6013 (N_6013,N_1858,N_4988);
nor U6014 (N_6014,N_4381,N_4320);
xor U6015 (N_6015,N_4439,N_3356);
nor U6016 (N_6016,N_3589,N_3571);
or U6017 (N_6017,N_586,N_2909);
nor U6018 (N_6018,N_579,N_3387);
and U6019 (N_6019,N_3575,N_2410);
nand U6020 (N_6020,N_2289,N_583);
nor U6021 (N_6021,N_3207,N_3424);
and U6022 (N_6022,N_1698,N_3117);
xnor U6023 (N_6023,N_3377,N_4082);
nor U6024 (N_6024,N_1732,N_4926);
and U6025 (N_6025,N_3407,N_3700);
and U6026 (N_6026,N_804,N_2026);
nand U6027 (N_6027,N_457,N_1866);
and U6028 (N_6028,N_3389,N_1543);
and U6029 (N_6029,N_2359,N_3298);
and U6030 (N_6030,N_4607,N_4011);
nand U6031 (N_6031,N_4522,N_2215);
xnor U6032 (N_6032,N_2804,N_4958);
or U6033 (N_6033,N_3564,N_3862);
or U6034 (N_6034,N_4349,N_959);
and U6035 (N_6035,N_2709,N_1282);
nand U6036 (N_6036,N_2325,N_1190);
nand U6037 (N_6037,N_1408,N_304);
nand U6038 (N_6038,N_1509,N_1924);
nand U6039 (N_6039,N_1719,N_192);
or U6040 (N_6040,N_2118,N_3052);
nor U6041 (N_6041,N_1484,N_503);
or U6042 (N_6042,N_2392,N_3896);
nor U6043 (N_6043,N_1053,N_4579);
nor U6044 (N_6044,N_4674,N_283);
or U6045 (N_6045,N_3523,N_4658);
xor U6046 (N_6046,N_473,N_2978);
nor U6047 (N_6047,N_1648,N_3332);
nand U6048 (N_6048,N_4689,N_1098);
nand U6049 (N_6049,N_1196,N_1871);
and U6050 (N_6050,N_4506,N_2086);
and U6051 (N_6051,N_2107,N_1023);
nor U6052 (N_6052,N_1597,N_2999);
or U6053 (N_6053,N_3360,N_2796);
or U6054 (N_6054,N_4225,N_1129);
nor U6055 (N_6055,N_929,N_4985);
or U6056 (N_6056,N_2591,N_3657);
nand U6057 (N_6057,N_15,N_1460);
nand U6058 (N_6058,N_257,N_633);
or U6059 (N_6059,N_214,N_3365);
nand U6060 (N_6060,N_796,N_435);
nor U6061 (N_6061,N_4103,N_1791);
nand U6062 (N_6062,N_3153,N_1662);
nand U6063 (N_6063,N_3361,N_3415);
and U6064 (N_6064,N_3876,N_4310);
nand U6065 (N_6065,N_1931,N_100);
and U6066 (N_6066,N_3178,N_2894);
and U6067 (N_6067,N_1423,N_324);
nand U6068 (N_6068,N_740,N_2968);
and U6069 (N_6069,N_4875,N_494);
or U6070 (N_6070,N_224,N_2553);
or U6071 (N_6071,N_365,N_885);
or U6072 (N_6072,N_95,N_230);
nand U6073 (N_6073,N_124,N_3471);
or U6074 (N_6074,N_1927,N_4703);
or U6075 (N_6075,N_3096,N_1293);
and U6076 (N_6076,N_2438,N_831);
nor U6077 (N_6077,N_2822,N_713);
or U6078 (N_6078,N_914,N_3449);
nor U6079 (N_6079,N_3940,N_2431);
nand U6080 (N_6080,N_2126,N_4991);
nor U6081 (N_6081,N_4321,N_1570);
or U6082 (N_6082,N_2918,N_2588);
nor U6083 (N_6083,N_1471,N_624);
and U6084 (N_6084,N_2418,N_3397);
nor U6085 (N_6085,N_4824,N_3627);
nand U6086 (N_6086,N_385,N_4374);
nor U6087 (N_6087,N_2779,N_1358);
or U6088 (N_6088,N_3133,N_4650);
and U6089 (N_6089,N_863,N_989);
nand U6090 (N_6090,N_4598,N_4694);
and U6091 (N_6091,N_3062,N_4641);
nand U6092 (N_6092,N_909,N_3622);
and U6093 (N_6093,N_2754,N_4876);
nand U6094 (N_6094,N_2874,N_2652);
nor U6095 (N_6095,N_500,N_3109);
nor U6096 (N_6096,N_1674,N_4307);
nand U6097 (N_6097,N_3197,N_3623);
or U6098 (N_6098,N_366,N_216);
or U6099 (N_6099,N_4070,N_474);
nor U6100 (N_6100,N_1352,N_3009);
nor U6101 (N_6101,N_2783,N_3983);
or U6102 (N_6102,N_3301,N_2842);
nor U6103 (N_6103,N_3230,N_847);
nand U6104 (N_6104,N_3310,N_4272);
or U6105 (N_6105,N_803,N_284);
nand U6106 (N_6106,N_1273,N_2001);
or U6107 (N_6107,N_1892,N_567);
nor U6108 (N_6108,N_943,N_3625);
and U6109 (N_6109,N_3272,N_1679);
nor U6110 (N_6110,N_3624,N_1575);
or U6111 (N_6111,N_868,N_3067);
or U6112 (N_6112,N_1752,N_821);
and U6113 (N_6113,N_2269,N_1311);
xor U6114 (N_6114,N_1180,N_4503);
nand U6115 (N_6115,N_1897,N_4956);
and U6116 (N_6116,N_3653,N_3737);
or U6117 (N_6117,N_4064,N_352);
nor U6118 (N_6118,N_3076,N_4678);
nor U6119 (N_6119,N_1531,N_2989);
nand U6120 (N_6120,N_1641,N_1721);
nand U6121 (N_6121,N_2015,N_2206);
nor U6122 (N_6122,N_4797,N_530);
nand U6123 (N_6123,N_3438,N_1846);
nor U6124 (N_6124,N_534,N_1873);
and U6125 (N_6125,N_4591,N_1268);
nand U6126 (N_6126,N_3149,N_1968);
nor U6127 (N_6127,N_1925,N_916);
nand U6128 (N_6128,N_3822,N_1712);
nor U6129 (N_6129,N_1409,N_2018);
nor U6130 (N_6130,N_2584,N_285);
and U6131 (N_6131,N_3445,N_4964);
and U6132 (N_6132,N_3510,N_1963);
nand U6133 (N_6133,N_423,N_3708);
or U6134 (N_6134,N_2200,N_4325);
nor U6135 (N_6135,N_2809,N_788);
and U6136 (N_6136,N_68,N_3470);
or U6137 (N_6137,N_1656,N_1459);
nand U6138 (N_6138,N_2929,N_4855);
nand U6139 (N_6139,N_3552,N_1275);
nor U6140 (N_6140,N_3590,N_462);
nor U6141 (N_6141,N_114,N_354);
and U6142 (N_6142,N_4104,N_4648);
nor U6143 (N_6143,N_357,N_1952);
or U6144 (N_6144,N_2621,N_595);
nand U6145 (N_6145,N_4354,N_3100);
nor U6146 (N_6146,N_3221,N_3089);
nand U6147 (N_6147,N_3139,N_3730);
nor U6148 (N_6148,N_3182,N_1672);
and U6149 (N_6149,N_4596,N_1814);
nor U6150 (N_6150,N_4492,N_662);
nor U6151 (N_6151,N_2928,N_3099);
or U6152 (N_6152,N_2229,N_1479);
nor U6153 (N_6153,N_1147,N_155);
nand U6154 (N_6154,N_892,N_4387);
or U6155 (N_6155,N_966,N_1183);
and U6156 (N_6156,N_2297,N_2669);
nand U6157 (N_6157,N_1258,N_4710);
nor U6158 (N_6158,N_3551,N_4005);
or U6159 (N_6159,N_4659,N_471);
nor U6160 (N_6160,N_3409,N_3920);
and U6161 (N_6161,N_871,N_4739);
xor U6162 (N_6162,N_4171,N_2364);
nor U6163 (N_6163,N_2734,N_4331);
and U6164 (N_6164,N_4280,N_4768);
and U6165 (N_6165,N_4716,N_87);
nand U6166 (N_6166,N_2171,N_363);
nand U6167 (N_6167,N_808,N_39);
nor U6168 (N_6168,N_2000,N_1872);
xor U6169 (N_6169,N_2608,N_3921);
and U6170 (N_6170,N_3985,N_3080);
nand U6171 (N_6171,N_2399,N_1540);
xor U6172 (N_6172,N_2228,N_3081);
or U6173 (N_6173,N_202,N_294);
or U6174 (N_6174,N_791,N_4677);
or U6175 (N_6175,N_4184,N_1659);
and U6176 (N_6176,N_2157,N_3898);
nand U6177 (N_6177,N_1075,N_1045);
nand U6178 (N_6178,N_2650,N_1104);
and U6179 (N_6179,N_1762,N_1792);
nor U6180 (N_6180,N_308,N_1703);
and U6181 (N_6181,N_4300,N_934);
xnor U6182 (N_6182,N_4043,N_1440);
nand U6183 (N_6183,N_1685,N_1536);
nand U6184 (N_6184,N_1153,N_2063);
or U6185 (N_6185,N_605,N_1298);
nor U6186 (N_6186,N_27,N_181);
and U6187 (N_6187,N_375,N_3742);
nor U6188 (N_6188,N_2695,N_1990);
nor U6189 (N_6189,N_1067,N_4842);
nor U6190 (N_6190,N_4218,N_875);
and U6191 (N_6191,N_1530,N_4125);
nand U6192 (N_6192,N_983,N_3091);
or U6193 (N_6193,N_3916,N_930);
nor U6194 (N_6194,N_3206,N_1579);
or U6195 (N_6195,N_4635,N_3376);
or U6196 (N_6196,N_613,N_94);
or U6197 (N_6197,N_1354,N_25);
or U6198 (N_6198,N_4861,N_2555);
and U6199 (N_6199,N_2823,N_4395);
nor U6200 (N_6200,N_2727,N_4382);
nor U6201 (N_6201,N_2043,N_4660);
nor U6202 (N_6202,N_3259,N_1112);
nor U6203 (N_6203,N_1635,N_2059);
or U6204 (N_6204,N_2568,N_2793);
nor U6205 (N_6205,N_2330,N_3102);
nor U6206 (N_6206,N_321,N_3804);
nor U6207 (N_6207,N_190,N_135);
or U6208 (N_6208,N_2756,N_2691);
or U6209 (N_6209,N_3877,N_680);
nor U6210 (N_6210,N_4259,N_1105);
nor U6211 (N_6211,N_3488,N_3300);
or U6212 (N_6212,N_223,N_548);
or U6213 (N_6213,N_738,N_2536);
or U6214 (N_6214,N_4737,N_34);
nand U6215 (N_6215,N_3608,N_4145);
nand U6216 (N_6216,N_2580,N_4929);
and U6217 (N_6217,N_3706,N_4508);
and U6218 (N_6218,N_3544,N_815);
nand U6219 (N_6219,N_3805,N_4911);
and U6220 (N_6220,N_850,N_3423);
or U6221 (N_6221,N_3541,N_1490);
nand U6222 (N_6222,N_3293,N_464);
and U6223 (N_6223,N_4858,N_198);
nand U6224 (N_6224,N_3532,N_3403);
nor U6225 (N_6225,N_881,N_2159);
nand U6226 (N_6226,N_2170,N_4185);
and U6227 (N_6227,N_4928,N_697);
nand U6228 (N_6228,N_4053,N_2423);
and U6229 (N_6229,N_393,N_4976);
or U6230 (N_6230,N_3169,N_126);
nor U6231 (N_6231,N_832,N_1057);
and U6232 (N_6232,N_2637,N_1629);
or U6233 (N_6233,N_3254,N_979);
or U6234 (N_6234,N_4437,N_4306);
nor U6235 (N_6235,N_2314,N_482);
and U6236 (N_6236,N_2665,N_3962);
or U6237 (N_6237,N_1210,N_4308);
xnor U6238 (N_6238,N_4126,N_4021);
nor U6239 (N_6239,N_3731,N_4785);
and U6240 (N_6240,N_4505,N_2786);
or U6241 (N_6241,N_4541,N_656);
and U6242 (N_6242,N_4865,N_1984);
or U6243 (N_6243,N_1114,N_671);
nand U6244 (N_6244,N_2611,N_660);
and U6245 (N_6245,N_4322,N_4097);
and U6246 (N_6246,N_1221,N_4358);
and U6247 (N_6247,N_861,N_2630);
nand U6248 (N_6248,N_484,N_4827);
and U6249 (N_6249,N_1042,N_71);
or U6250 (N_6250,N_1110,N_2237);
or U6251 (N_6251,N_4078,N_3947);
or U6252 (N_6252,N_4130,N_1818);
nor U6253 (N_6253,N_3761,N_2758);
nor U6254 (N_6254,N_3922,N_3525);
nor U6255 (N_6255,N_1683,N_2361);
or U6256 (N_6256,N_1345,N_2080);
nor U6257 (N_6257,N_3329,N_1361);
or U6258 (N_6258,N_4963,N_3782);
nor U6259 (N_6259,N_2208,N_3547);
or U6260 (N_6260,N_3890,N_3152);
nor U6261 (N_6261,N_1226,N_4838);
or U6262 (N_6262,N_4938,N_2678);
and U6263 (N_6263,N_1029,N_4809);
or U6264 (N_6264,N_859,N_351);
or U6265 (N_6265,N_2101,N_205);
nor U6266 (N_6266,N_862,N_2369);
and U6267 (N_6267,N_4252,N_131);
and U6268 (N_6268,N_2987,N_2493);
nand U6269 (N_6269,N_540,N_4686);
and U6270 (N_6270,N_977,N_920);
nand U6271 (N_6271,N_1730,N_2109);
nand U6272 (N_6272,N_2443,N_1247);
nand U6273 (N_6273,N_4691,N_2262);
nor U6274 (N_6274,N_242,N_4073);
or U6275 (N_6275,N_1100,N_4663);
and U6276 (N_6276,N_1794,N_1404);
or U6277 (N_6277,N_3528,N_4235);
nor U6278 (N_6278,N_941,N_3548);
xnor U6279 (N_6279,N_928,N_4201);
nand U6280 (N_6280,N_3583,N_4137);
or U6281 (N_6281,N_2009,N_2182);
and U6282 (N_6282,N_3160,N_3966);
nor U6283 (N_6283,N_2788,N_4355);
nand U6284 (N_6284,N_1784,N_4412);
xnor U6285 (N_6285,N_1942,N_4651);
nor U6286 (N_6286,N_4888,N_4236);
and U6287 (N_6287,N_917,N_521);
or U6288 (N_6288,N_3952,N_3637);
nor U6289 (N_6289,N_2469,N_1930);
xor U6290 (N_6290,N_3186,N_1775);
and U6291 (N_6291,N_4182,N_781);
nor U6292 (N_6292,N_1564,N_4533);
xor U6293 (N_6293,N_3313,N_272);
xnor U6294 (N_6294,N_2967,N_940);
nor U6295 (N_6295,N_702,N_3726);
nor U6296 (N_6296,N_876,N_3585);
or U6297 (N_6297,N_968,N_2975);
or U6298 (N_6298,N_4743,N_1523);
nand U6299 (N_6299,N_1084,N_1976);
nor U6300 (N_6300,N_2337,N_144);
nand U6301 (N_6301,N_1094,N_3485);
and U6302 (N_6302,N_2726,N_3578);
xnor U6303 (N_6303,N_4328,N_4642);
or U6304 (N_6304,N_2085,N_3848);
and U6305 (N_6305,N_3386,N_2523);
nand U6306 (N_6306,N_2479,N_1242);
nor U6307 (N_6307,N_834,N_72);
or U6308 (N_6308,N_481,N_1595);
and U6309 (N_6309,N_299,N_4411);
nor U6310 (N_6310,N_1527,N_3910);
nand U6311 (N_6311,N_3988,N_1870);
and U6312 (N_6312,N_1852,N_3312);
nand U6313 (N_6313,N_748,N_1508);
and U6314 (N_6314,N_2252,N_3390);
nor U6315 (N_6315,N_2844,N_1159);
nor U6316 (N_6316,N_1522,N_3265);
nor U6317 (N_6317,N_4079,N_2603);
and U6318 (N_6318,N_83,N_3505);
and U6319 (N_6319,N_3385,N_2821);
and U6320 (N_6320,N_3506,N_3598);
nor U6321 (N_6321,N_3664,N_1816);
and U6322 (N_6322,N_2165,N_1663);
or U6323 (N_6323,N_3392,N_1988);
nor U6324 (N_6324,N_1166,N_139);
nor U6325 (N_6325,N_3796,N_4543);
or U6326 (N_6326,N_136,N_171);
nor U6327 (N_6327,N_1458,N_1414);
nand U6328 (N_6328,N_3635,N_59);
nand U6329 (N_6329,N_3427,N_1828);
nand U6330 (N_6330,N_1005,N_123);
nand U6331 (N_6331,N_320,N_2331);
nor U6332 (N_6332,N_4251,N_763);
and U6333 (N_6333,N_573,N_2318);
or U6334 (N_6334,N_1347,N_3696);
nor U6335 (N_6335,N_3008,N_322);
and U6336 (N_6336,N_710,N_4039);
and U6337 (N_6337,N_2891,N_3710);
nor U6338 (N_6338,N_1489,N_1215);
and U6339 (N_6339,N_550,N_3173);
nor U6340 (N_6340,N_4595,N_4444);
and U6341 (N_6341,N_4623,N_4332);
and U6342 (N_6342,N_2906,N_2006);
and U6343 (N_6343,N_4175,N_3559);
nor U6344 (N_6344,N_2622,N_1059);
nand U6345 (N_6345,N_4376,N_47);
xor U6346 (N_6346,N_3702,N_3618);
nand U6347 (N_6347,N_3374,N_3569);
and U6348 (N_6348,N_4791,N_4592);
and U6349 (N_6349,N_1165,N_1362);
nand U6350 (N_6350,N_496,N_2942);
or U6351 (N_6351,N_1928,N_4549);
or U6352 (N_6352,N_1339,N_4406);
xnor U6353 (N_6353,N_3884,N_3352);
or U6354 (N_6354,N_4133,N_82);
nor U6355 (N_6355,N_927,N_3955);
or U6356 (N_6356,N_92,N_502);
nand U6357 (N_6357,N_2137,N_233);
xnor U6358 (N_6358,N_4482,N_185);
and U6359 (N_6359,N_582,N_577);
and U6360 (N_6360,N_1052,N_445);
and U6361 (N_6361,N_2372,N_4760);
nand U6362 (N_6362,N_3440,N_1369);
and U6363 (N_6363,N_2892,N_2355);
and U6364 (N_6364,N_4787,N_1750);
nor U6365 (N_6365,N_46,N_4155);
or U6366 (N_6366,N_4330,N_335);
nand U6367 (N_6367,N_2654,N_2389);
and U6368 (N_6368,N_4742,N_2683);
and U6369 (N_6369,N_4602,N_346);
or U6370 (N_6370,N_508,N_2799);
or U6371 (N_6371,N_1314,N_3350);
nand U6372 (N_6372,N_591,N_3255);
or U6373 (N_6373,N_4957,N_442);
and U6374 (N_6374,N_4072,N_824);
or U6375 (N_6375,N_1294,N_3630);
and U6376 (N_6376,N_4290,N_1037);
nand U6377 (N_6377,N_597,N_298);
or U6378 (N_6378,N_4578,N_682);
nand U6379 (N_6379,N_2807,N_2467);
and U6380 (N_6380,N_1723,N_1545);
and U6381 (N_6381,N_3290,N_2946);
nor U6382 (N_6382,N_1661,N_2710);
or U6383 (N_6383,N_2872,N_2247);
and U6384 (N_6384,N_2590,N_376);
and U6385 (N_6385,N_1621,N_994);
nand U6386 (N_6386,N_2847,N_56);
or U6387 (N_6387,N_691,N_4334);
nand U6388 (N_6388,N_467,N_1946);
and U6389 (N_6389,N_2749,N_1978);
and U6390 (N_6390,N_1590,N_4548);
and U6391 (N_6391,N_1903,N_3279);
nand U6392 (N_6392,N_206,N_4144);
and U6393 (N_6393,N_3935,N_3022);
nor U6394 (N_6394,N_3113,N_2944);
or U6395 (N_6395,N_4454,N_4769);
xor U6396 (N_6396,N_1300,N_1019);
and U6397 (N_6397,N_3582,N_3201);
and U6398 (N_6398,N_3264,N_3527);
nor U6399 (N_6399,N_3225,N_2468);
nor U6400 (N_6400,N_2990,N_1276);
nor U6401 (N_6401,N_498,N_4102);
nand U6402 (N_6402,N_698,N_4353);
nor U6403 (N_6403,N_1152,N_3323);
nand U6404 (N_6404,N_2119,N_2972);
nor U6405 (N_6405,N_3253,N_3999);
or U6406 (N_6406,N_102,N_3148);
nor U6407 (N_6407,N_3616,N_596);
nand U6408 (N_6408,N_3939,N_150);
xnor U6409 (N_6409,N_3739,N_138);
nand U6410 (N_6410,N_826,N_3175);
or U6411 (N_6411,N_3680,N_3064);
and U6412 (N_6412,N_1729,N_690);
nor U6413 (N_6413,N_4317,N_2977);
nand U6414 (N_6414,N_2067,N_2614);
or U6415 (N_6415,N_2513,N_358);
and U6416 (N_6416,N_1620,N_3882);
and U6417 (N_6417,N_1604,N_757);
and U6418 (N_6418,N_2480,N_2078);
and U6419 (N_6419,N_4535,N_3621);
nand U6420 (N_6420,N_4810,N_3482);
nor U6421 (N_6421,N_2155,N_4871);
or U6422 (N_6422,N_1076,N_4971);
or U6423 (N_6423,N_3227,N_678);
nand U6424 (N_6424,N_4315,N_3558);
nor U6425 (N_6425,N_4058,N_4873);
nor U6426 (N_6426,N_1446,N_857);
nor U6427 (N_6427,N_4177,N_2292);
or U6428 (N_6428,N_3267,N_4265);
and U6429 (N_6429,N_3752,N_2379);
and U6430 (N_6430,N_237,N_3775);
nand U6431 (N_6431,N_753,N_2662);
nor U6432 (N_6432,N_997,N_4139);
nor U6433 (N_6433,N_3714,N_2951);
or U6434 (N_6434,N_2184,N_4262);
and U6435 (N_6435,N_4269,N_4192);
and U6436 (N_6436,N_4336,N_1938);
nand U6437 (N_6437,N_1418,N_315);
nor U6438 (N_6438,N_4129,N_2759);
and U6439 (N_6439,N_4846,N_337);
or U6440 (N_6440,N_3273,N_1046);
nand U6441 (N_6441,N_1985,N_3327);
nand U6442 (N_6442,N_958,N_4401);
or U6443 (N_6443,N_1151,N_4108);
nor U6444 (N_6444,N_2708,N_1106);
and U6445 (N_6445,N_35,N_2738);
nor U6446 (N_6446,N_2815,N_3779);
nand U6447 (N_6447,N_3678,N_469);
nor U6448 (N_6448,N_880,N_4655);
nand U6449 (N_6449,N_869,N_1633);
or U6450 (N_6450,N_4250,N_425);
or U6451 (N_6451,N_1581,N_2129);
and U6452 (N_6452,N_1745,N_2280);
nand U6453 (N_6453,N_422,N_133);
nand U6454 (N_6454,N_3053,N_2755);
or U6455 (N_6455,N_110,N_18);
nor U6456 (N_6456,N_2066,N_3953);
nand U6457 (N_6457,N_367,N_4851);
or U6458 (N_6458,N_3287,N_2537);
xor U6459 (N_6459,N_105,N_3658);
or U6460 (N_6460,N_3431,N_924);
nand U6461 (N_6461,N_3097,N_4960);
or U6462 (N_6462,N_60,N_203);
nor U6463 (N_6463,N_4610,N_2903);
nor U6464 (N_6464,N_1841,N_787);
nand U6465 (N_6465,N_3116,N_4413);
or U6466 (N_6466,N_2697,N_2939);
or U6467 (N_6467,N_4357,N_3362);
or U6468 (N_6468,N_2532,N_4033);
and U6469 (N_6469,N_3493,N_4509);
nand U6470 (N_6470,N_2729,N_2074);
and U6471 (N_6471,N_3125,N_379);
nand U6472 (N_6472,N_1088,N_2546);
nand U6473 (N_6473,N_4213,N_4402);
nor U6474 (N_6474,N_2534,N_1291);
and U6475 (N_6475,N_2460,N_2716);
and U6476 (N_6476,N_884,N_535);
or U6477 (N_6477,N_1030,N_3418);
nand U6478 (N_6478,N_3933,N_4612);
or U6479 (N_6479,N_3302,N_2236);
nand U6480 (N_6480,N_53,N_1327);
nand U6481 (N_6481,N_2011,N_4682);
nor U6482 (N_6482,N_1329,N_3141);
nor U6483 (N_6483,N_162,N_2227);
and U6484 (N_6484,N_4718,N_1617);
or U6485 (N_6485,N_4532,N_3480);
and U6486 (N_6486,N_3026,N_2966);
or U6487 (N_6487,N_4630,N_2714);
nor U6488 (N_6488,N_2346,N_431);
and U6489 (N_6489,N_542,N_1538);
nand U6490 (N_6490,N_362,N_4101);
nand U6491 (N_6491,N_410,N_79);
or U6492 (N_6492,N_4127,N_3843);
or U6493 (N_6493,N_399,N_4925);
and U6494 (N_6494,N_727,N_4937);
and U6495 (N_6495,N_3146,N_2680);
nor U6496 (N_6496,N_252,N_1400);
or U6497 (N_6497,N_268,N_1315);
nand U6498 (N_6498,N_143,N_4954);
and U6499 (N_6499,N_1480,N_1319);
nor U6500 (N_6500,N_1301,N_4747);
nand U6501 (N_6501,N_1179,N_3981);
or U6502 (N_6502,N_3515,N_1544);
nand U6503 (N_6503,N_3179,N_1898);
and U6504 (N_6504,N_3246,N_789);
nand U6505 (N_6505,N_2720,N_1753);
and U6506 (N_6506,N_81,N_4397);
or U6507 (N_6507,N_1498,N_4879);
or U6508 (N_6508,N_3846,N_156);
nor U6509 (N_6509,N_260,N_2520);
and U6510 (N_6510,N_776,N_3900);
nor U6511 (N_6511,N_2656,N_4621);
nand U6512 (N_6512,N_2595,N_756);
or U6513 (N_6513,N_4687,N_2097);
xor U6514 (N_6514,N_872,N_2526);
and U6515 (N_6515,N_383,N_4866);
or U6516 (N_6516,N_3283,N_4997);
nand U6517 (N_6517,N_1542,N_2941);
and U6518 (N_6518,N_3056,N_2567);
or U6519 (N_6519,N_2612,N_4672);
nand U6520 (N_6520,N_2740,N_2694);
nand U6521 (N_6521,N_1160,N_3799);
and U6522 (N_6522,N_2813,N_4564);
or U6523 (N_6523,N_2543,N_174);
or U6524 (N_6524,N_4806,N_2745);
nor U6525 (N_6525,N_3467,N_737);
or U6526 (N_6526,N_2765,N_1254);
nand U6527 (N_6527,N_4844,N_4573);
and U6528 (N_6528,N_4400,N_2172);
nor U6529 (N_6529,N_2433,N_4899);
nor U6530 (N_6530,N_4160,N_1016);
or U6531 (N_6531,N_1639,N_228);
nor U6532 (N_6532,N_3002,N_1257);
nor U6533 (N_6533,N_2463,N_2725);
nor U6534 (N_6534,N_2499,N_1214);
nor U6535 (N_6535,N_4792,N_2900);
nor U6536 (N_6536,N_2147,N_747);
or U6537 (N_6537,N_2787,N_1466);
nand U6538 (N_6538,N_4513,N_448);
nor U6539 (N_6539,N_1429,N_4363);
nor U6540 (N_6540,N_141,N_1919);
nor U6541 (N_6541,N_1024,N_1342);
nand U6542 (N_6542,N_3925,N_2223);
nor U6543 (N_6543,N_4973,N_3969);
nor U6544 (N_6544,N_2175,N_506);
nand U6545 (N_6545,N_1355,N_1411);
and U6546 (N_6546,N_2610,N_1379);
nor U6547 (N_6547,N_3956,N_1286);
and U6548 (N_6548,N_234,N_438);
and U6549 (N_6549,N_2087,N_1027);
or U6550 (N_6550,N_97,N_4377);
or U6551 (N_6551,N_108,N_4263);
or U6552 (N_6552,N_4834,N_398);
and U6553 (N_6553,N_4589,N_3987);
xnor U6554 (N_6554,N_3257,N_3344);
and U6555 (N_6555,N_991,N_3964);
or U6556 (N_6556,N_1569,N_3800);
nor U6557 (N_6557,N_2884,N_557);
nand U6558 (N_6558,N_1720,N_4135);
and U6559 (N_6559,N_4414,N_4922);
and U6560 (N_6560,N_1853,N_4084);
nor U6561 (N_6561,N_3811,N_3199);
nor U6562 (N_6562,N_4238,N_2336);
or U6563 (N_6563,N_4243,N_3465);
nor U6564 (N_6564,N_3134,N_3640);
nand U6565 (N_6565,N_2214,N_4709);
and U6566 (N_6566,N_1996,N_1078);
or U6567 (N_6567,N_222,N_1883);
or U6568 (N_6568,N_4576,N_1081);
nand U6569 (N_6569,N_3084,N_2177);
nor U6570 (N_6570,N_4935,N_2908);
nand U6571 (N_6571,N_70,N_88);
or U6572 (N_6572,N_2587,N_3549);
and U6573 (N_6573,N_2895,N_4156);
nor U6574 (N_6574,N_4483,N_2875);
nor U6575 (N_6575,N_3384,N_2605);
nand U6576 (N_6576,N_637,N_1113);
and U6577 (N_6577,N_1905,N_2310);
or U6578 (N_6578,N_4836,N_2501);
or U6579 (N_6579,N_3886,N_4080);
or U6580 (N_6580,N_4520,N_2659);
or U6581 (N_6581,N_3699,N_2149);
nor U6582 (N_6582,N_1225,N_4464);
or U6583 (N_6583,N_1041,N_4817);
or U6584 (N_6584,N_4869,N_2741);
nor U6585 (N_6585,N_4653,N_2204);
and U6586 (N_6586,N_1060,N_4511);
nor U6587 (N_6587,N_2557,N_4526);
nand U6588 (N_6588,N_3239,N_1714);
or U6589 (N_6589,N_4248,N_3414);
or U6590 (N_6590,N_2404,N_777);
or U6591 (N_6591,N_2589,N_2120);
nand U6592 (N_6592,N_1382,N_3679);
and U6593 (N_6593,N_4477,N_3895);
nor U6594 (N_6594,N_2751,N_1431);
and U6595 (N_6595,N_4038,N_1759);
nor U6596 (N_6596,N_2161,N_2299);
and U6597 (N_6597,N_900,N_3218);
nor U6598 (N_6598,N_2038,N_3);
nor U6599 (N_6599,N_969,N_1142);
and U6600 (N_6600,N_2081,N_766);
or U6601 (N_6601,N_14,N_795);
xor U6602 (N_6602,N_898,N_3176);
or U6603 (N_6603,N_208,N_386);
xor U6604 (N_6604,N_446,N_4204);
nor U6605 (N_6605,N_4604,N_1568);
or U6606 (N_6606,N_4384,N_2057);
nand U6607 (N_6607,N_844,N_1578);
or U6608 (N_6608,N_1495,N_3316);
nand U6609 (N_6609,N_1879,N_3250);
and U6610 (N_6610,N_2213,N_1277);
or U6611 (N_6611,N_2027,N_2864);
and U6612 (N_6612,N_631,N_327);
and U6613 (N_6613,N_4085,N_2256);
and U6614 (N_6614,N_2529,N_3959);
and U6615 (N_6615,N_4799,N_2434);
or U6616 (N_6616,N_2767,N_4748);
xor U6617 (N_6617,N_517,N_3413);
nor U6618 (N_6618,N_1121,N_3984);
nand U6619 (N_6619,N_4271,N_2041);
nor U6620 (N_6620,N_3213,N_3198);
xnor U6621 (N_6621,N_3425,N_341);
nor U6622 (N_6622,N_3609,N_3095);
nand U6623 (N_6623,N_38,N_2104);
or U6624 (N_6624,N_1832,N_3131);
and U6625 (N_6625,N_4067,N_2572);
and U6626 (N_6626,N_2436,N_3070);
nand U6627 (N_6627,N_151,N_1074);
nand U6628 (N_6628,N_2857,N_1177);
or U6629 (N_6629,N_3917,N_2521);
nand U6630 (N_6630,N_4723,N_1970);
nor U6631 (N_6631,N_2040,N_754);
or U6632 (N_6632,N_2712,N_3484);
nor U6633 (N_6633,N_4624,N_2472);
and U6634 (N_6634,N_4891,N_3214);
nand U6635 (N_6635,N_1966,N_1865);
nand U6636 (N_6636,N_360,N_1691);
nand U6637 (N_6637,N_2965,N_3503);
nand U6638 (N_6638,N_2679,N_902);
nor U6639 (N_6639,N_225,N_2703);
and U6640 (N_6640,N_2772,N_2167);
or U6641 (N_6641,N_3147,N_3960);
or U6642 (N_6642,N_4823,N_2397);
nor U6643 (N_6643,N_3164,N_4327);
and U6644 (N_6644,N_1539,N_1317);
nand U6645 (N_6645,N_681,N_3792);
nand U6646 (N_6646,N_1187,N_437);
or U6647 (N_6647,N_3400,N_537);
or U6648 (N_6648,N_3209,N_1922);
nand U6649 (N_6649,N_4695,N_610);
and U6650 (N_6650,N_3850,N_4488);
nor U6651 (N_6651,N_4870,N_2542);
or U6652 (N_6652,N_1090,N_3010);
or U6653 (N_6653,N_4232,N_172);
nor U6654 (N_6654,N_720,N_3195);
nand U6655 (N_6655,N_1580,N_650);
nand U6656 (N_6656,N_907,N_4654);
and U6657 (N_6657,N_2402,N_3620);
nor U6658 (N_6658,N_1365,N_3049);
nor U6659 (N_6659,N_2757,N_2700);
xor U6660 (N_6660,N_2784,N_2693);
or U6661 (N_6661,N_1087,N_118);
and U6662 (N_6662,N_23,N_4731);
or U6663 (N_6663,N_4462,N_4673);
nand U6664 (N_6664,N_694,N_1708);
or U6665 (N_6665,N_1222,N_819);
nand U6666 (N_6666,N_3367,N_2910);
nand U6667 (N_6667,N_1039,N_2350);
nand U6668 (N_6668,N_2525,N_3478);
or U6669 (N_6669,N_2342,N_965);
nand U6670 (N_6670,N_408,N_2473);
and U6671 (N_6671,N_4022,N_4568);
nand U6672 (N_6672,N_4656,N_1348);
nand U6673 (N_6673,N_2455,N_2927);
and U6674 (N_6674,N_2365,N_922);
or U6675 (N_6675,N_4486,N_576);
or U6676 (N_6676,N_2422,N_3685);
nor U6677 (N_6677,N_270,N_2715);
nand U6678 (N_6678,N_2012,N_652);
and U6679 (N_6679,N_2777,N_2994);
and U6680 (N_6680,N_1546,N_2020);
nor U6681 (N_6681,N_3880,N_1392);
nand U6682 (N_6682,N_246,N_2829);
and U6683 (N_6683,N_3380,N_2219);
nor U6684 (N_6684,N_4180,N_3595);
nor U6685 (N_6685,N_4110,N_4912);
and U6686 (N_6686,N_2907,N_2836);
nor U6687 (N_6687,N_3820,N_3129);
or U6688 (N_6688,N_4342,N_546);
nor U6689 (N_6689,N_98,N_405);
and U6690 (N_6690,N_4668,N_2574);
and U6691 (N_6691,N_1741,N_714);
and U6692 (N_6692,N_4489,N_3863);
and U6693 (N_6693,N_2024,N_659);
nor U6694 (N_6694,N_2478,N_3014);
or U6695 (N_6695,N_2311,N_3755);
or U6696 (N_6696,N_1330,N_2465);
or U6697 (N_6697,N_4468,N_4329);
and U6698 (N_6698,N_783,N_3161);
and U6699 (N_6699,N_3345,N_3038);
or U6700 (N_6700,N_2527,N_106);
and U6701 (N_6701,N_2698,N_568);
and U6702 (N_6702,N_2551,N_1649);
and U6703 (N_6703,N_2267,N_3722);
nand U6704 (N_6704,N_4264,N_4441);
nand U6705 (N_6705,N_4216,N_1453);
nand U6706 (N_6706,N_4493,N_2601);
and U6707 (N_6707,N_3324,N_883);
xnor U6708 (N_6708,N_2658,N_667);
nand U6709 (N_6709,N_182,N_4802);
nand U6710 (N_6710,N_1786,N_433);
and U6711 (N_6711,N_2245,N_2413);
or U6712 (N_6712,N_4944,N_4361);
or U6713 (N_6713,N_4399,N_949);
or U6714 (N_6714,N_4894,N_1627);
or U6715 (N_6715,N_55,N_4098);
or U6716 (N_6716,N_2915,N_48);
nand U6717 (N_6717,N_592,N_310);
xor U6718 (N_6718,N_2887,N_2016);
and U6719 (N_6719,N_1806,N_3422);
or U6720 (N_6720,N_1228,N_797);
nor U6721 (N_6721,N_2021,N_490);
or U6722 (N_6722,N_2511,N_4882);
and U6723 (N_6723,N_3395,N_4109);
and U6724 (N_6724,N_3477,N_127);
nand U6725 (N_6725,N_897,N_4203);
and U6726 (N_6726,N_1309,N_1422);
and U6727 (N_6727,N_2613,N_3990);
nand U6728 (N_6728,N_2139,N_1000);
and U6729 (N_6729,N_752,N_598);
or U6730 (N_6730,N_1108,N_640);
and U6731 (N_6731,N_2178,N_1908);
or U6732 (N_6732,N_1313,N_4393);
and U6733 (N_6733,N_814,N_4419);
and U6734 (N_6734,N_2390,N_1289);
nor U6735 (N_6735,N_3270,N_3554);
or U6736 (N_6736,N_3600,N_4777);
nand U6737 (N_6737,N_4801,N_1889);
or U6738 (N_6738,N_4571,N_4784);
or U6739 (N_6739,N_447,N_1603);
and U6740 (N_6740,N_1316,N_2481);
or U6741 (N_6741,N_1001,N_2889);
nand U6742 (N_6742,N_1283,N_1610);
nand U6743 (N_6743,N_2179,N_3747);
and U6744 (N_6744,N_4147,N_307);
or U6745 (N_6745,N_2920,N_2114);
and U6746 (N_6746,N_3612,N_3057);
nor U6747 (N_6747,N_3294,N_4425);
and U6748 (N_6748,N_1497,N_1428);
or U6749 (N_6749,N_2005,N_1982);
and U6750 (N_6750,N_1980,N_4531);
and U6751 (N_6751,N_555,N_4054);
nand U6752 (N_6752,N_3893,N_2743);
or U6753 (N_6753,N_4759,N_3236);
nand U6754 (N_6754,N_2641,N_3020);
nand U6755 (N_6755,N_2044,N_1954);
nand U6756 (N_6756,N_58,N_1902);
nor U6757 (N_6757,N_936,N_2859);
and U6758 (N_6758,N_4685,N_2902);
nand U6759 (N_6759,N_3342,N_889);
nor U6760 (N_6760,N_1233,N_3143);
nand U6761 (N_6761,N_3238,N_2644);
or U6762 (N_6762,N_3325,N_5);
or U6763 (N_6763,N_2962,N_1737);
and U6764 (N_6764,N_2440,N_3358);
nor U6765 (N_6765,N_3668,N_3823);
or U6766 (N_6766,N_69,N_1246);
nand U6767 (N_6767,N_2728,N_331);
nor U6768 (N_6768,N_2419,N_4666);
nand U6769 (N_6769,N_4440,N_625);
and U6770 (N_6770,N_4538,N_266);
nor U6771 (N_6771,N_3560,N_4268);
or U6772 (N_6772,N_1457,N_142);
or U6773 (N_6773,N_2002,N_649);
nand U6774 (N_6774,N_566,N_289);
nor U6775 (N_6775,N_2560,N_2042);
nor U6776 (N_6776,N_4567,N_3074);
nor U6777 (N_6777,N_953,N_1867);
or U6778 (N_6778,N_4389,N_4680);
nand U6779 (N_6779,N_980,N_1770);
nand U6780 (N_6780,N_3019,N_2224);
nor U6781 (N_6781,N_623,N_4179);
and U6782 (N_6782,N_3873,N_4378);
and U6783 (N_6783,N_4831,N_2007);
or U6784 (N_6784,N_4480,N_2446);
nor U6785 (N_6785,N_1150,N_292);
xnor U6786 (N_6786,N_109,N_1868);
nor U6787 (N_6787,N_3732,N_1364);
and U6788 (N_6788,N_2660,N_1407);
nor U6789 (N_6789,N_1601,N_1111);
and U6790 (N_6790,N_2471,N_3816);
nor U6791 (N_6791,N_4664,N_4638);
xnor U6792 (N_6792,N_2647,N_2370);
nor U6793 (N_6793,N_2970,N_3645);
nand U6794 (N_6794,N_3256,N_4059);
nor U6795 (N_6795,N_4212,N_429);
or U6796 (N_6796,N_428,N_4679);
nor U6797 (N_6797,N_4071,N_4153);
nand U6798 (N_6798,N_1664,N_2713);
nand U6799 (N_6799,N_2818,N_2790);
nor U6800 (N_6800,N_2627,N_2079);
or U6801 (N_6801,N_3079,N_3308);
nor U6802 (N_6802,N_4542,N_915);
or U6803 (N_6803,N_3487,N_4276);
or U6804 (N_6804,N_3282,N_528);
or U6805 (N_6805,N_3605,N_4949);
and U6806 (N_6806,N_4030,N_1915);
or U6807 (N_6807,N_507,N_3435);
nor U6808 (N_6808,N_3475,N_3735);
xor U6809 (N_6809,N_101,N_3729);
xor U6810 (N_6810,N_4048,N_3085);
nand U6811 (N_6811,N_3689,N_3223);
or U6812 (N_6812,N_485,N_2333);
and U6813 (N_6813,N_3233,N_2439);
nor U6814 (N_6814,N_3184,N_323);
nand U6815 (N_6815,N_998,N_2547);
and U6816 (N_6816,N_3461,N_1715);
or U6817 (N_6817,N_4373,N_1032);
nor U6818 (N_6818,N_2191,N_4200);
or U6819 (N_6819,N_2550,N_3724);
nor U6820 (N_6820,N_3675,N_3661);
and U6821 (N_6821,N_810,N_4628);
or U6822 (N_6822,N_1652,N_3996);
nand U6823 (N_6823,N_558,N_4228);
nand U6824 (N_6824,N_3649,N_2681);
nand U6825 (N_6825,N_2711,N_1224);
and U6826 (N_6826,N_1320,N_1713);
and U6827 (N_6827,N_1877,N_2648);
nand U6828 (N_6828,N_812,N_3909);
or U6829 (N_6829,N_3587,N_1880);
nand U6830 (N_6830,N_1248,N_2293);
and U6831 (N_6831,N_2374,N_1947);
nor U6832 (N_6832,N_3644,N_62);
nand U6833 (N_6833,N_2142,N_2582);
or U6834 (N_6834,N_1080,N_3757);
or U6835 (N_6835,N_1270,N_2811);
nor U6836 (N_6836,N_1644,N_4142);
nand U6837 (N_6837,N_3196,N_389);
nor U6838 (N_6838,N_3087,N_3219);
nor U6839 (N_6839,N_4552,N_1383);
or U6840 (N_6840,N_2209,N_4516);
nand U6841 (N_6841,N_3035,N_57);
nor U6842 (N_6842,N_3103,N_1069);
nand U6843 (N_6843,N_3906,N_1758);
and U6844 (N_6844,N_2490,N_4924);
or U6845 (N_6845,N_648,N_4392);
and U6846 (N_6846,N_1995,N_3366);
or U6847 (N_6847,N_2010,N_2046);
nor U6848 (N_6848,N_4474,N_2461);
and U6849 (N_6849,N_3602,N_4507);
nand U6850 (N_6850,N_4087,N_3249);
nor U6851 (N_6851,N_4611,N_1502);
and U6852 (N_6852,N_2378,N_2558);
or U6853 (N_6853,N_2890,N_3138);
and U6854 (N_6854,N_3784,N_2753);
nand U6855 (N_6855,N_4819,N_1842);
or U6856 (N_6856,N_627,N_2400);
nand U6857 (N_6857,N_2190,N_2846);
and U6858 (N_6858,N_4178,N_4114);
nor U6859 (N_6859,N_333,N_4569);
nand U6860 (N_6860,N_2629,N_4847);
xnor U6861 (N_6861,N_2877,N_2345);
and U6862 (N_6862,N_2265,N_1089);
and U6863 (N_6863,N_701,N_668);
nor U6864 (N_6864,N_3224,N_3155);
nand U6865 (N_6865,N_2800,N_3703);
or U6866 (N_6866,N_1801,N_3526);
and U6867 (N_6867,N_3088,N_3490);
or U6868 (N_6868,N_4942,N_199);
nor U6869 (N_6869,N_2198,N_1174);
or U6870 (N_6870,N_316,N_41);
or U6871 (N_6871,N_3442,N_2);
nor U6872 (N_6872,N_3753,N_4242);
and U6873 (N_6873,N_1499,N_2375);
or U6874 (N_6874,N_3628,N_45);
or U6875 (N_6875,N_1571,N_4282);
and U6876 (N_6876,N_1561,N_4675);
nand U6877 (N_6877,N_4460,N_2037);
nand U6878 (N_6878,N_1430,N_1824);
nand U6879 (N_6879,N_3671,N_2724);
nor U6880 (N_6880,N_4853,N_4138);
and U6881 (N_6881,N_4311,N_148);
nor U6882 (N_6882,N_529,N_1821);
nor U6883 (N_6883,N_3697,N_458);
or U6884 (N_6884,N_1456,N_762);
nand U6885 (N_6885,N_1467,N_2642);
and U6886 (N_6886,N_3903,N_3787);
or U6887 (N_6887,N_2466,N_3317);
or U6888 (N_6888,N_4832,N_1827);
or U6889 (N_6889,N_2351,N_4514);
nand U6890 (N_6890,N_480,N_707);
or U6891 (N_6891,N_3489,N_4371);
nand U6892 (N_6892,N_1951,N_2089);
nor U6893 (N_6893,N_3536,N_3711);
or U6894 (N_6894,N_4939,N_1899);
or U6895 (N_6895,N_4643,N_466);
or U6896 (N_6896,N_1975,N_4950);
nand U6897 (N_6897,N_1718,N_1667);
and U6898 (N_6898,N_1854,N_1234);
and U6899 (N_6899,N_630,N_1589);
xnor U6900 (N_6900,N_4314,N_40);
or U6901 (N_6901,N_3018,N_2596);
nor U6902 (N_6902,N_1923,N_2347);
nand U6903 (N_6903,N_2335,N_4992);
nand U6904 (N_6904,N_2835,N_4877);
and U6905 (N_6905,N_4165,N_3126);
nand U6906 (N_6906,N_2230,N_1168);
and U6907 (N_6907,N_430,N_732);
nand U6908 (N_6908,N_937,N_1171);
and U6909 (N_6909,N_2428,N_3736);
nand U6910 (N_6910,N_3576,N_91);
or U6911 (N_6911,N_2677,N_3454);
or U6912 (N_6912,N_1102,N_3995);
nor U6913 (N_6913,N_1475,N_1455);
nand U6914 (N_6914,N_3180,N_2218);
xor U6915 (N_6915,N_1070,N_865);
xnor U6916 (N_6916,N_4193,N_1336);
nor U6917 (N_6917,N_2974,N_3771);
nand U6918 (N_6918,N_4715,N_3809);
nor U6919 (N_6919,N_1018,N_2592);
nand U6920 (N_6920,N_2031,N_4159);
nor U6921 (N_6921,N_750,N_231);
or U6922 (N_6922,N_1363,N_1134);
nor U6923 (N_6923,N_2352,N_2911);
and U6924 (N_6924,N_4521,N_3613);
nor U6925 (N_6925,N_4217,N_887);
nand U6926 (N_6926,N_905,N_840);
nor U6927 (N_6927,N_1971,N_2904);
and U6928 (N_6928,N_3021,N_1388);
and U6929 (N_6929,N_2871,N_2239);
and U6930 (N_6930,N_2357,N_860);
nor U6931 (N_6931,N_1993,N_4961);
nand U6932 (N_6932,N_2721,N_2263);
nand U6933 (N_6933,N_1934,N_3315);
or U6934 (N_6934,N_886,N_3538);
nor U6935 (N_6935,N_3044,N_2640);
and U6936 (N_6936,N_646,N_3991);
and U6937 (N_6937,N_2298,N_4042);
nand U6938 (N_6938,N_2356,N_2169);
nor U6939 (N_6939,N_1040,N_4536);
or U6940 (N_6940,N_4868,N_4745);
and U6941 (N_6941,N_2437,N_1748);
nor U6942 (N_6942,N_2039,N_1133);
nand U6943 (N_6943,N_441,N_4550);
or U6944 (N_6944,N_4752,N_1864);
xnor U6945 (N_6945,N_4736,N_4818);
nor U6946 (N_6946,N_132,N_2702);
nor U6947 (N_6947,N_3883,N_4804);
and U6948 (N_6948,N_4214,N_1368);
nand U6949 (N_6949,N_3746,N_3191);
or U6950 (N_6950,N_676,N_1725);
nor U6951 (N_6951,N_1860,N_263);
nor U6952 (N_6952,N_4640,N_3372);
and U6953 (N_6953,N_54,N_2264);
or U6954 (N_6954,N_1895,N_3869);
and U6955 (N_6955,N_2136,N_1307);
or U6956 (N_6956,N_3306,N_2070);
or U6957 (N_6957,N_4239,N_1533);
and U6958 (N_6958,N_4662,N_1241);
xor U6959 (N_6959,N_760,N_1653);
nor U6960 (N_6960,N_2084,N_17);
or U6961 (N_6961,N_910,N_4237);
nor U6962 (N_6962,N_1284,N_1302);
nand U6963 (N_6963,N_4090,N_1882);
nor U6964 (N_6964,N_1148,N_2897);
nand U6965 (N_6965,N_522,N_3434);
or U6966 (N_6966,N_1787,N_3370);
or U6967 (N_6967,N_1548,N_396);
nor U6968 (N_6968,N_2739,N_1593);
nor U6969 (N_6969,N_4701,N_3918);
nand U6970 (N_6970,N_2383,N_563);
and U6971 (N_6971,N_2687,N_4274);
or U6972 (N_6972,N_2508,N_511);
or U6973 (N_6973,N_4132,N_2108);
nand U6974 (N_6974,N_1823,N_194);
and U6975 (N_6975,N_2953,N_864);
and U6976 (N_6976,N_4863,N_1524);
nand U6977 (N_6977,N_2127,N_2343);
or U6978 (N_6978,N_3667,N_3665);
or U6979 (N_6979,N_267,N_1937);
nand U6980 (N_6980,N_3232,N_3457);
nor U6981 (N_6981,N_1608,N_653);
and U6982 (N_6982,N_4181,N_4431);
nor U6983 (N_6983,N_3187,N_3005);
or U6984 (N_6984,N_3951,N_1958);
nand U6985 (N_6985,N_622,N_2594);
nand U6986 (N_6986,N_1587,N_1488);
or U6987 (N_6987,N_4734,N_4661);
and U6988 (N_6988,N_2017,N_4867);
or U6989 (N_6989,N_996,N_4982);
nand U6990 (N_6990,N_245,N_1454);
nor U6991 (N_6991,N_2676,N_1678);
nor U6992 (N_6992,N_2956,N_3517);
and U6993 (N_6993,N_4009,N_666);
and U6994 (N_6994,N_3491,N_3858);
nor U6995 (N_6995,N_3614,N_2102);
and U6996 (N_6996,N_3355,N_276);
and U6997 (N_6997,N_2733,N_2373);
or U6998 (N_6998,N_3321,N_4987);
nor U6999 (N_6999,N_269,N_2530);
nor U7000 (N_7000,N_1398,N_1817);
nand U7001 (N_7001,N_4302,N_2984);
nor U7002 (N_7002,N_4829,N_3094);
nand U7003 (N_7003,N_733,N_4430);
or U7004 (N_7004,N_1236,N_2976);
and U7005 (N_7005,N_4603,N_3580);
nand U7006 (N_7006,N_4037,N_2153);
nor U7007 (N_7007,N_4255,N_1785);
nor U7008 (N_7008,N_4367,N_811);
or U7009 (N_7009,N_1372,N_4076);
or U7010 (N_7010,N_741,N_2309);
nor U7011 (N_7011,N_664,N_1660);
nand U7012 (N_7012,N_2360,N_1269);
nand U7013 (N_7013,N_532,N_2980);
and U7014 (N_7014,N_2696,N_197);
or U7015 (N_7015,N_4197,N_4727);
nor U7016 (N_7016,N_3803,N_2442);
nand U7017 (N_7017,N_3881,N_1376);
nor U7018 (N_7018,N_1520,N_1356);
nor U7019 (N_7019,N_1779,N_913);
nor U7020 (N_7020,N_765,N_213);
nor U7021 (N_7021,N_2615,N_4013);
or U7022 (N_7022,N_1890,N_4445);
xnor U7023 (N_7023,N_4515,N_3781);
xor U7024 (N_7024,N_1851,N_1402);
nand U7025 (N_7025,N_4408,N_3944);
nor U7026 (N_7026,N_817,N_813);
or U7027 (N_7027,N_4995,N_381);
and U7028 (N_7028,N_3012,N_4862);
or U7029 (N_7029,N_3101,N_259);
and U7030 (N_7030,N_2462,N_2029);
and U7031 (N_7031,N_4676,N_4501);
and U7032 (N_7032,N_340,N_2913);
and U7033 (N_7033,N_2843,N_3240);
nand U7034 (N_7034,N_1483,N_2451);
nand U7035 (N_7035,N_378,N_908);
nor U7036 (N_7036,N_4199,N_4833);
nand U7037 (N_7037,N_3725,N_4711);
nor U7038 (N_7038,N_1412,N_2958);
and U7039 (N_7039,N_2232,N_3718);
nand U7040 (N_7040,N_22,N_3789);
or U7041 (N_7041,N_1296,N_4475);
and U7042 (N_7042,N_115,N_3518);
nand U7043 (N_7043,N_935,N_1856);
or U7044 (N_7044,N_2055,N_2326);
or U7045 (N_7045,N_1157,N_2763);
and U7046 (N_7046,N_4931,N_961);
nand U7047 (N_7047,N_570,N_4904);
and U7048 (N_7048,N_4466,N_440);
nor U7049 (N_7049,N_2174,N_2633);
nor U7050 (N_7050,N_3632,N_1139);
and U7051 (N_7051,N_3247,N_990);
nand U7052 (N_7052,N_790,N_2571);
or U7053 (N_7053,N_651,N_2287);
nand U7054 (N_7054,N_4190,N_4210);
nor U7055 (N_7055,N_4206,N_3297);
nor U7056 (N_7056,N_4390,N_76);
nand U7057 (N_7057,N_4352,N_3899);
nand U7058 (N_7058,N_1907,N_1109);
nand U7059 (N_7059,N_3211,N_1647);
nor U7060 (N_7060,N_2056,N_281);
nand U7061 (N_7061,N_2096,N_4930);
nand U7062 (N_7062,N_4086,N_545);
and U7063 (N_7063,N_2053,N_2317);
and U7064 (N_7064,N_227,N_2062);
or U7065 (N_7065,N_2098,N_456);
xnor U7066 (N_7066,N_3840,N_1896);
or U7067 (N_7067,N_2363,N_4285);
and U7068 (N_7068,N_1305,N_3701);
or U7069 (N_7069,N_603,N_4556);
and U7070 (N_7070,N_4270,N_523);
nand U7071 (N_7071,N_572,N_3229);
and U7072 (N_7072,N_3349,N_1706);
xnor U7073 (N_7073,N_1136,N_1710);
or U7074 (N_7074,N_1011,N_4463);
nand U7075 (N_7075,N_4024,N_3670);
and U7076 (N_7076,N_1822,N_1063);
or U7077 (N_7077,N_3825,N_1839);
or U7078 (N_7078,N_287,N_3535);
or U7079 (N_7079,N_1068,N_2246);
or U7080 (N_7080,N_84,N_74);
nand U7081 (N_7081,N_2699,N_673);
nand U7082 (N_7082,N_3507,N_1146);
xor U7083 (N_7083,N_219,N_725);
and U7084 (N_7084,N_3606,N_3013);
or U7085 (N_7085,N_3588,N_4518);
or U7086 (N_7086,N_4398,N_4379);
or U7087 (N_7087,N_3375,N_2831);
nand U7088 (N_7088,N_3756,N_2131);
xnor U7089 (N_7089,N_1768,N_4601);
nand U7090 (N_7090,N_1051,N_4697);
nor U7091 (N_7091,N_2047,N_677);
and U7092 (N_7092,N_2761,N_1940);
or U7093 (N_7093,N_4119,N_486);
nand U7094 (N_7094,N_2071,N_533);
or U7095 (N_7095,N_2254,N_2488);
nand U7096 (N_7096,N_193,N_3786);
and U7097 (N_7097,N_3672,N_2334);
nor U7098 (N_7098,N_2577,N_1292);
or U7099 (N_7099,N_4036,N_3004);
nand U7100 (N_7100,N_4615,N_3826);
and U7101 (N_7101,N_718,N_1328);
and U7102 (N_7102,N_1202,N_3866);
nor U7103 (N_7103,N_4211,N_2395);
and U7104 (N_7104,N_4323,N_3208);
nor U7105 (N_7105,N_1144,N_4424);
and U7106 (N_7106,N_2338,N_3586);
nand U7107 (N_7107,N_4999,N_4266);
nand U7108 (N_7108,N_4420,N_1486);
and U7109 (N_7109,N_4560,N_4194);
or U7110 (N_7110,N_1826,N_400);
xnor U7111 (N_7111,N_2388,N_806);
nor U7112 (N_7112,N_468,N_2035);
or U7113 (N_7113,N_3572,N_2947);
and U7114 (N_7114,N_1534,N_672);
and U7115 (N_7115,N_1064,N_319);
nand U7116 (N_7116,N_3495,N_1939);
nand U7117 (N_7117,N_3639,N_3929);
and U7118 (N_7118,N_1658,N_2628);
or U7119 (N_7119,N_1532,N_2150);
and U7120 (N_7120,N_1468,N_4766);
and U7121 (N_7121,N_3078,N_3650);
or U7122 (N_7122,N_2255,N_4690);
nor U7123 (N_7123,N_3437,N_665);
and U7124 (N_7124,N_4840,N_3364);
nor U7125 (N_7125,N_4966,N_459);
xnor U7126 (N_7126,N_4918,N_200);
nand U7127 (N_7127,N_3251,N_2277);
or U7128 (N_7128,N_761,N_436);
or U7129 (N_7129,N_2862,N_416);
nor U7130 (N_7130,N_4758,N_2231);
nor U7131 (N_7131,N_1820,N_3479);
nor U7132 (N_7132,N_4427,N_2586);
and U7133 (N_7133,N_722,N_1394);
and U7134 (N_7134,N_1933,N_3842);
or U7135 (N_7135,N_1008,N_539);
or U7136 (N_7136,N_1602,N_1073);
nand U7137 (N_7137,N_830,N_2186);
nand U7138 (N_7138,N_2123,N_3970);
xor U7139 (N_7139,N_3252,N_489);
or U7140 (N_7140,N_4945,N_3156);
or U7141 (N_7141,N_3263,N_1439);
nor U7142 (N_7142,N_4765,N_3958);
or U7143 (N_7143,N_1072,N_311);
nand U7144 (N_7144,N_4790,N_347);
or U7145 (N_7145,N_3648,N_4298);
or U7146 (N_7146,N_175,N_2411);
nand U7147 (N_7147,N_2323,N_2973);
nor U7148 (N_7148,N_187,N_2424);
and U7149 (N_7149,N_2008,N_1308);
nor U7150 (N_7150,N_2414,N_769);
nor U7151 (N_7151,N_3814,N_3318);
or U7152 (N_7152,N_1733,N_618);
and U7153 (N_7153,N_256,N_1370);
nand U7154 (N_7154,N_4234,N_2624);
or U7155 (N_7155,N_723,N_513);
and U7156 (N_7156,N_1830,N_2830);
or U7157 (N_7157,N_3039,N_4639);
nand U7158 (N_7158,N_985,N_2597);
nor U7159 (N_7159,N_1584,N_4304);
nor U7160 (N_7160,N_4632,N_3563);
nand U7161 (N_7161,N_794,N_2160);
and U7162 (N_7162,N_4452,N_3957);
nand U7163 (N_7163,N_838,N_3073);
and U7164 (N_7164,N_609,N_2945);
nand U7165 (N_7165,N_963,N_2549);
and U7166 (N_7166,N_89,N_2140);
nor U7167 (N_7167,N_3522,N_1140);
and U7168 (N_7168,N_2183,N_4497);
and U7169 (N_7169,N_1835,N_2873);
and U7170 (N_7170,N_32,N_1259);
nor U7171 (N_7171,N_3764,N_3432);
or U7172 (N_7172,N_4170,N_554);
nand U7173 (N_7173,N_3743,N_541);
nand U7174 (N_7174,N_3961,N_1893);
nand U7175 (N_7175,N_3382,N_4461);
nand U7176 (N_7176,N_2983,N_4347);
nor U7177 (N_7177,N_4874,N_2448);
nor U7178 (N_7178,N_4351,N_4974);
and U7179 (N_7179,N_2004,N_2524);
nor U7180 (N_7180,N_955,N_3790);
nor U7181 (N_7181,N_981,N_2065);
and U7182 (N_7182,N_3271,N_1096);
nand U7183 (N_7183,N_2482,N_2516);
nand U7184 (N_7184,N_1263,N_1367);
and U7185 (N_7185,N_2302,N_309);
nor U7186 (N_7186,N_2306,N_1727);
or U7187 (N_7187,N_2760,N_1973);
nand U7188 (N_7188,N_1780,N_1416);
or U7189 (N_7189,N_2707,N_3581);
nor U7190 (N_7190,N_536,N_1612);
or U7191 (N_7191,N_384,N_2022);
and U7192 (N_7192,N_4100,N_1560);
or U7193 (N_7193,N_3584,N_250);
nand U7194 (N_7194,N_3751,N_1386);
nor U7195 (N_7195,N_4735,N_4226);
or U7196 (N_7196,N_923,N_4224);
or U7197 (N_7197,N_4113,N_2789);
nor U7198 (N_7198,N_476,N_296);
and U7199 (N_7199,N_451,N_3157);
xor U7200 (N_7200,N_455,N_833);
or U7201 (N_7201,N_3136,N_1552);
or U7202 (N_7202,N_43,N_326);
nor U7203 (N_7203,N_904,N_2855);
nand U7204 (N_7204,N_3610,N_1504);
nand U7205 (N_7205,N_2033,N_1812);
nor U7206 (N_7206,N_1700,N_1756);
and U7207 (N_7207,N_1557,N_1600);
nand U7208 (N_7208,N_1435,N_2870);
or U7209 (N_7209,N_2686,N_4528);
nor U7210 (N_7210,N_3244,N_1209);
nor U7211 (N_7211,N_2176,N_4588);
or U7212 (N_7212,N_3281,N_849);
and U7213 (N_7213,N_99,N_2477);
nor U7214 (N_7214,N_1048,N_4256);
nor U7215 (N_7215,N_4189,N_4161);
nor U7216 (N_7216,N_2545,N_1863);
nor U7217 (N_7217,N_1216,N_719);
nand U7218 (N_7218,N_4117,N_477);
nor U7219 (N_7219,N_505,N_3111);
and U7220 (N_7220,N_3835,N_4288);
nor U7221 (N_7221,N_1921,N_4055);
nor U7222 (N_7222,N_1585,N_4391);
nand U7223 (N_7223,N_588,N_4409);
nor U7224 (N_7224,N_4771,N_3235);
and U7225 (N_7225,N_3902,N_3993);
and U7226 (N_7226,N_2766,N_683);
nor U7227 (N_7227,N_2950,N_1798);
or U7228 (N_7228,N_411,N_2573);
or U7229 (N_7229,N_4913,N_4380);
nand U7230 (N_7230,N_4529,N_993);
and U7231 (N_7231,N_1598,N_1772);
nor U7232 (N_7232,N_3077,N_1378);
or U7233 (N_7233,N_3430,N_669);
or U7234 (N_7234,N_2538,N_2251);
nand U7235 (N_7235,N_1397,N_107);
nor U7236 (N_7236,N_2819,N_4584);
or U7237 (N_7237,N_3122,N_4438);
nand U7238 (N_7238,N_1050,N_3913);
nand U7239 (N_7239,N_2301,N_2307);
nand U7240 (N_7240,N_709,N_370);
nand U7241 (N_7241,N_2848,N_11);
nor U7242 (N_7242,N_2919,N_176);
nand U7243 (N_7243,N_978,N_147);
and U7244 (N_7244,N_1485,N_1551);
nor U7245 (N_7245,N_3217,N_1838);
and U7246 (N_7246,N_2770,N_2485);
and U7247 (N_7247,N_1396,N_3912);
and U7248 (N_7248,N_3821,N_2130);
nor U7249 (N_7249,N_4886,N_1281);
or U7250 (N_7250,N_4923,N_4647);
nor U7251 (N_7251,N_2509,N_3037);
nand U7252 (N_7252,N_2731,N_3634);
or U7253 (N_7253,N_2152,N_2671);
nor U7254 (N_7254,N_4927,N_2876);
and U7255 (N_7255,N_2673,N_1506);
and U7256 (N_7256,N_2771,N_2701);
nand U7257 (N_7257,N_1175,N_3393);
or U7258 (N_7258,N_1197,N_2216);
nand U7259 (N_7259,N_2371,N_4470);
and U7260 (N_7260,N_1353,N_3629);
nand U7261 (N_7261,N_3740,N_4007);
nor U7262 (N_7262,N_3946,N_184);
nand U7263 (N_7263,N_1049,N_3123);
nand U7264 (N_7264,N_1834,N_986);
nor U7265 (N_7265,N_647,N_1932);
or U7266 (N_7266,N_1424,N_3159);
or U7267 (N_7267,N_65,N_3923);
and U7268 (N_7268,N_3135,N_2626);
nor U7269 (N_7269,N_4692,N_822);
nor U7270 (N_7270,N_86,N_1751);
or U7271 (N_7271,N_4459,N_657);
nand U7272 (N_7272,N_3363,N_1795);
nor U7273 (N_7273,N_4057,N_2050);
nor U7274 (N_7274,N_4993,N_12);
and U7275 (N_7275,N_4807,N_2593);
or U7276 (N_7276,N_404,N_2083);
nand U7277 (N_7277,N_4744,N_749);
or U7278 (N_7278,N_3533,N_2795);
or U7279 (N_7279,N_2348,N_439);
xor U7280 (N_7280,N_3594,N_3778);
nor U7281 (N_7281,N_2060,N_3514);
or U7282 (N_7282,N_211,N_1266);
nand U7283 (N_7283,N_236,N_61);
or U7284 (N_7284,N_4405,N_4417);
nor U7285 (N_7285,N_4186,N_2664);
or U7286 (N_7286,N_971,N_2949);
nor U7287 (N_7287,N_504,N_2556);
nor U7288 (N_7288,N_705,N_3248);
nor U7289 (N_7289,N_2979,N_2704);
and U7290 (N_7290,N_1444,N_1757);
or U7291 (N_7291,N_1677,N_493);
nand U7292 (N_7292,N_313,N_3574);
and U7293 (N_7293,N_950,N_2489);
nor U7294 (N_7294,N_764,N_488);
or U7295 (N_7295,N_4850,N_4502);
nor U7296 (N_7296,N_3619,N_2860);
nor U7297 (N_7297,N_450,N_4728);
or U7298 (N_7298,N_1800,N_641);
or U7299 (N_7299,N_2316,N_1012);
or U7300 (N_7300,N_4943,N_2510);
nand U7301 (N_7301,N_4041,N_2519);
and U7302 (N_7302,N_1773,N_463);
nand U7303 (N_7303,N_1673,N_4946);
and U7304 (N_7304,N_899,N_2116);
nor U7305 (N_7305,N_4450,N_4539);
or U7306 (N_7306,N_3499,N_2886);
and U7307 (N_7307,N_3269,N_3234);
and U7308 (N_7308,N_1724,N_3812);
nand U7309 (N_7309,N_258,N_4060);
nand U7310 (N_7310,N_1420,N_1734);
nor U7311 (N_7311,N_1195,N_2583);
xor U7312 (N_7312,N_4717,N_4903);
and U7313 (N_7313,N_3262,N_4583);
and U7314 (N_7314,N_1692,N_4350);
and U7315 (N_7315,N_3274,N_4597);
or U7316 (N_7316,N_1686,N_4221);
or U7317 (N_7317,N_1781,N_3086);
or U7318 (N_7318,N_2146,N_4712);
or U7319 (N_7319,N_186,N_1351);
or U7320 (N_7320,N_3405,N_3785);
nor U7321 (N_7321,N_1443,N_4345);
nor U7322 (N_7322,N_3292,N_149);
nor U7323 (N_7323,N_2115,N_4083);
and U7324 (N_7324,N_1239,N_4046);
nor U7325 (N_7325,N_4188,N_2774);
and U7326 (N_7326,N_3124,N_2762);
and U7327 (N_7327,N_4977,N_4032);
or U7328 (N_7328,N_4561,N_1769);
or U7329 (N_7329,N_2868,N_3464);
nand U7330 (N_7330,N_2675,N_1092);
or U7331 (N_7331,N_743,N_189);
or U7332 (N_7332,N_414,N_1684);
or U7333 (N_7333,N_3727,N_2401);
nand U7334 (N_7334,N_932,N_3617);
and U7335 (N_7335,N_4049,N_2319);
or U7336 (N_7336,N_4338,N_3098);
nor U7337 (N_7337,N_2930,N_2276);
nor U7338 (N_7338,N_4249,N_4000);
and U7339 (N_7339,N_2133,N_3090);
nand U7340 (N_7340,N_1290,N_1514);
xnor U7341 (N_7341,N_1253,N_1384);
and U7342 (N_7342,N_4775,N_2776);
nor U7343 (N_7343,N_2561,N_1373);
nor U7344 (N_7344,N_2736,N_903);
or U7345 (N_7345,N_4557,N_4278);
and U7346 (N_7346,N_372,N_4633);
or U7347 (N_7347,N_2281,N_37);
and U7348 (N_7348,N_3220,N_2988);
and U7349 (N_7349,N_3975,N_1130);
nand U7350 (N_7350,N_4546,N_4593);
or U7351 (N_7351,N_3643,N_619);
or U7352 (N_7352,N_2328,N_2425);
nand U7353 (N_7353,N_552,N_3941);
or U7354 (N_7354,N_2210,N_2339);
nand U7355 (N_7355,N_3016,N_4967);
nor U7356 (N_7356,N_2061,N_820);
nand U7357 (N_7357,N_2506,N_1323);
nor U7358 (N_7358,N_1482,N_3772);
nor U7359 (N_7359,N_2327,N_2045);
and U7360 (N_7360,N_524,N_1007);
or U7361 (N_7361,N_947,N_675);
or U7362 (N_7362,N_1979,N_4335);
or U7363 (N_7363,N_1017,N_893);
or U7364 (N_7364,N_2880,N_2320);
nor U7365 (N_7365,N_3845,N_3001);
nor U7366 (N_7366,N_2475,N_4394);
nor U7367 (N_7367,N_3904,N_3319);
nand U7368 (N_7368,N_2013,N_1478);
nor U7369 (N_7369,N_2600,N_275);
or U7370 (N_7370,N_4637,N_531);
nand U7371 (N_7371,N_3531,N_3276);
or U7372 (N_7372,N_4473,N_1141);
and U7373 (N_7373,N_165,N_113);
and U7374 (N_7374,N_4619,N_3048);
nor U7375 (N_7375,N_2854,N_1126);
nand U7376 (N_7376,N_2775,N_1107);
and U7377 (N_7377,N_984,N_3011);
or U7378 (N_7378,N_332,N_520);
nand U7379 (N_7379,N_1341,N_1194);
or U7380 (N_7380,N_4081,N_1240);
nor U7381 (N_7381,N_1131,N_3017);
nor U7382 (N_7382,N_4442,N_1389);
or U7383 (N_7383,N_2197,N_800);
or U7384 (N_7384,N_4500,N_3295);
and U7385 (N_7385,N_1127,N_293);
or U7386 (N_7386,N_1626,N_4813);
and U7387 (N_7387,N_1774,N_894);
nand U7388 (N_7388,N_632,N_2385);
nor U7389 (N_7389,N_1819,N_4428);
and U7390 (N_7390,N_4798,N_2003);
or U7391 (N_7391,N_700,N_2073);
and U7392 (N_7392,N_1594,N_1058);
and U7393 (N_7393,N_645,N_1380);
nor U7394 (N_7394,N_2867,N_3463);
and U7395 (N_7395,N_409,N_173);
or U7396 (N_7396,N_4403,N_265);
nor U7397 (N_7397,N_4890,N_2522);
nor U7398 (N_7398,N_2163,N_2407);
nand U7399 (N_7399,N_2663,N_1391);
or U7400 (N_7400,N_4970,N_1998);
and U7401 (N_7401,N_580,N_1743);
nand U7402 (N_7402,N_3603,N_1343);
or U7403 (N_7403,N_3068,N_3104);
nand U7404 (N_7404,N_3443,N_2393);
and U7405 (N_7405,N_3891,N_4749);
nand U7406 (N_7406,N_1655,N_4003);
and U7407 (N_7407,N_4472,N_3579);
or U7408 (N_7408,N_2852,N_215);
xor U7409 (N_7409,N_3071,N_1562);
nand U7410 (N_7410,N_164,N_1742);
and U7411 (N_7411,N_1642,N_3938);
nor U7412 (N_7412,N_290,N_3033);
nor U7413 (N_7413,N_2924,N_2535);
nor U7414 (N_7414,N_4845,N_1566);
and U7415 (N_7415,N_3210,N_125);
nand U7416 (N_7416,N_3027,N_3394);
and U7417 (N_7417,N_1218,N_4820);
nand U7418 (N_7418,N_1749,N_4494);
and U7419 (N_7419,N_356,N_1843);
and U7420 (N_7420,N_4066,N_460);
and U7421 (N_7421,N_3813,N_2051);
and U7422 (N_7422,N_1326,N_604);
and U7423 (N_7423,N_1796,N_1149);
nor U7424 (N_7424,N_2837,N_1526);
or U7425 (N_7425,N_3108,N_395);
or U7426 (N_7426,N_3115,N_3296);
nor U7427 (N_7427,N_3907,N_4362);
and U7428 (N_7428,N_4241,N_611);
and U7429 (N_7429,N_2444,N_4279);
nand U7430 (N_7430,N_3339,N_1559);
nand U7431 (N_7431,N_1213,N_2495);
or U7432 (N_7432,N_4433,N_2353);
nand U7433 (N_7433,N_1325,N_1619);
and U7434 (N_7434,N_4449,N_4446);
and U7435 (N_7435,N_2403,N_2828);
and U7436 (N_7436,N_2655,N_3128);
nand U7437 (N_7437,N_4581,N_2430);
nand U7438 (N_7438,N_944,N_4762);
nand U7439 (N_7439,N_1778,N_4525);
nand U7440 (N_7440,N_3412,N_1321);
or U7441 (N_7441,N_938,N_4246);
nand U7442 (N_7442,N_1310,N_2517);
and U7443 (N_7443,N_4297,N_2616);
nor U7444 (N_7444,N_3976,N_1120);
and U7445 (N_7445,N_3277,N_970);
nor U7446 (N_7446,N_987,N_569);
or U7447 (N_7447,N_2993,N_4233);
or U7448 (N_7448,N_621,N_4733);
or U7449 (N_7449,N_3633,N_2278);
and U7450 (N_7450,N_3741,N_4404);
and U7451 (N_7451,N_3936,N_3266);
nand U7452 (N_7452,N_3383,N_547);
nor U7453 (N_7453,N_2250,N_890);
or U7454 (N_7454,N_1707,N_3231);
and U7455 (N_7455,N_4010,N_2164);
and U7456 (N_7456,N_1231,N_3066);
and U7457 (N_7457,N_280,N_3519);
nand U7458 (N_7458,N_4434,N_273);
and U7459 (N_7459,N_4841,N_3949);
nor U7460 (N_7460,N_3769,N_3379);
nand U7461 (N_7461,N_3289,N_4168);
nor U7462 (N_7462,N_3140,N_1191);
or U7463 (N_7463,N_1158,N_1901);
and U7464 (N_7464,N_3977,N_2575);
xnor U7465 (N_7465,N_1117,N_4808);
nor U7466 (N_7466,N_2344,N_2552);
and U7467 (N_7467,N_3166,N_3568);
nand U7468 (N_7468,N_4455,N_2723);
nand U7469 (N_7469,N_3205,N_3819);
or U7470 (N_7470,N_658,N_4770);
nor U7471 (N_7471,N_2954,N_2635);
nand U7472 (N_7472,N_2394,N_1066);
nor U7473 (N_7473,N_78,N_4254);
or U7474 (N_7474,N_2917,N_1972);
and U7475 (N_7475,N_3919,N_1645);
nand U7476 (N_7476,N_4006,N_527);
and U7477 (N_7477,N_19,N_1572);
xor U7478 (N_7478,N_1505,N_674);
and U7479 (N_7479,N_2072,N_3911);
nand U7480 (N_7480,N_244,N_4296);
nand U7481 (N_7481,N_4365,N_2649);
or U7482 (N_7482,N_2427,N_4582);
and U7483 (N_7483,N_1521,N_3237);
nand U7484 (N_7484,N_2853,N_3368);
nor U7485 (N_7485,N_1887,N_2598);
and U7486 (N_7486,N_2202,N_3486);
nand U7487 (N_7487,N_3773,N_3466);
nor U7488 (N_7488,N_387,N_1390);
nand U7489 (N_7489,N_1020,N_4277);
nand U7490 (N_7490,N_2581,N_229);
nor U7491 (N_7491,N_975,N_3818);
and U7492 (N_7492,N_1761,N_1419);
nor U7493 (N_7493,N_1705,N_866);
xor U7494 (N_7494,N_3652,N_1071);
or U7495 (N_7495,N_1279,N_4341);
and U7496 (N_7496,N_1874,N_4416);
nor U7497 (N_7497,N_509,N_3543);
nand U7498 (N_7498,N_858,N_911);
nor U7499 (N_7499,N_4019,N_1255);
nand U7500 (N_7500,N_2298,N_2547);
and U7501 (N_7501,N_4576,N_1614);
and U7502 (N_7502,N_573,N_1016);
nor U7503 (N_7503,N_2374,N_966);
nand U7504 (N_7504,N_4973,N_1032);
and U7505 (N_7505,N_1997,N_3480);
nand U7506 (N_7506,N_1213,N_4261);
or U7507 (N_7507,N_1763,N_2774);
or U7508 (N_7508,N_2638,N_4402);
nor U7509 (N_7509,N_1392,N_929);
nand U7510 (N_7510,N_2091,N_1274);
or U7511 (N_7511,N_1618,N_1420);
nand U7512 (N_7512,N_3273,N_4884);
nor U7513 (N_7513,N_1426,N_978);
and U7514 (N_7514,N_1160,N_1144);
nor U7515 (N_7515,N_209,N_1822);
nor U7516 (N_7516,N_2572,N_2843);
nand U7517 (N_7517,N_880,N_969);
nand U7518 (N_7518,N_4841,N_4967);
nand U7519 (N_7519,N_1436,N_3041);
nor U7520 (N_7520,N_2272,N_31);
nand U7521 (N_7521,N_2138,N_2811);
nor U7522 (N_7522,N_3676,N_1823);
and U7523 (N_7523,N_695,N_2541);
nor U7524 (N_7524,N_472,N_1707);
and U7525 (N_7525,N_3244,N_3461);
nor U7526 (N_7526,N_52,N_2205);
and U7527 (N_7527,N_4699,N_607);
and U7528 (N_7528,N_488,N_1807);
nand U7529 (N_7529,N_1060,N_3337);
nor U7530 (N_7530,N_645,N_3409);
or U7531 (N_7531,N_1889,N_1087);
nor U7532 (N_7532,N_4516,N_1370);
and U7533 (N_7533,N_206,N_4394);
and U7534 (N_7534,N_207,N_3759);
nand U7535 (N_7535,N_4392,N_3439);
nand U7536 (N_7536,N_1625,N_2263);
nand U7537 (N_7537,N_2615,N_3289);
and U7538 (N_7538,N_803,N_1882);
xnor U7539 (N_7539,N_3190,N_230);
or U7540 (N_7540,N_262,N_354);
or U7541 (N_7541,N_3095,N_979);
and U7542 (N_7542,N_3164,N_3252);
nand U7543 (N_7543,N_821,N_1892);
nand U7544 (N_7544,N_3569,N_171);
xor U7545 (N_7545,N_2222,N_601);
and U7546 (N_7546,N_940,N_223);
nor U7547 (N_7547,N_811,N_4329);
or U7548 (N_7548,N_946,N_2139);
and U7549 (N_7549,N_2664,N_208);
or U7550 (N_7550,N_1589,N_3124);
nand U7551 (N_7551,N_277,N_2280);
nand U7552 (N_7552,N_4360,N_895);
and U7553 (N_7553,N_947,N_894);
nor U7554 (N_7554,N_4499,N_4157);
nand U7555 (N_7555,N_519,N_1909);
or U7556 (N_7556,N_4576,N_3550);
or U7557 (N_7557,N_2514,N_1151);
nor U7558 (N_7558,N_3356,N_1261);
nor U7559 (N_7559,N_4324,N_2949);
nor U7560 (N_7560,N_4518,N_1302);
and U7561 (N_7561,N_891,N_1989);
nor U7562 (N_7562,N_4357,N_10);
nor U7563 (N_7563,N_720,N_2475);
nand U7564 (N_7564,N_4345,N_4442);
and U7565 (N_7565,N_2280,N_1879);
or U7566 (N_7566,N_2364,N_3951);
and U7567 (N_7567,N_2228,N_3643);
and U7568 (N_7568,N_4353,N_1637);
nor U7569 (N_7569,N_4687,N_3362);
nor U7570 (N_7570,N_1459,N_2291);
nand U7571 (N_7571,N_2153,N_3623);
nand U7572 (N_7572,N_2305,N_1020);
nand U7573 (N_7573,N_4888,N_3424);
or U7574 (N_7574,N_4155,N_3188);
xnor U7575 (N_7575,N_4309,N_3900);
or U7576 (N_7576,N_2236,N_2998);
nor U7577 (N_7577,N_3953,N_1865);
nand U7578 (N_7578,N_2013,N_538);
and U7579 (N_7579,N_3058,N_3705);
nand U7580 (N_7580,N_4663,N_54);
and U7581 (N_7581,N_394,N_3522);
nor U7582 (N_7582,N_619,N_518);
nor U7583 (N_7583,N_122,N_2178);
and U7584 (N_7584,N_3975,N_3750);
and U7585 (N_7585,N_3444,N_4030);
nand U7586 (N_7586,N_28,N_4375);
or U7587 (N_7587,N_1397,N_4746);
nand U7588 (N_7588,N_2825,N_506);
or U7589 (N_7589,N_236,N_1290);
and U7590 (N_7590,N_3033,N_4769);
nand U7591 (N_7591,N_3485,N_1245);
or U7592 (N_7592,N_498,N_1331);
and U7593 (N_7593,N_1302,N_3818);
nor U7594 (N_7594,N_1998,N_4632);
and U7595 (N_7595,N_2057,N_2823);
or U7596 (N_7596,N_476,N_3453);
nand U7597 (N_7597,N_1726,N_1308);
and U7598 (N_7598,N_2459,N_2787);
nor U7599 (N_7599,N_474,N_4426);
and U7600 (N_7600,N_1524,N_2569);
and U7601 (N_7601,N_1193,N_275);
and U7602 (N_7602,N_2895,N_1692);
or U7603 (N_7603,N_2057,N_4022);
and U7604 (N_7604,N_1925,N_727);
nor U7605 (N_7605,N_3725,N_73);
nor U7606 (N_7606,N_501,N_1183);
nand U7607 (N_7607,N_1200,N_4070);
nand U7608 (N_7608,N_2708,N_4070);
nand U7609 (N_7609,N_645,N_4729);
and U7610 (N_7610,N_2536,N_2538);
or U7611 (N_7611,N_1549,N_300);
nor U7612 (N_7612,N_4385,N_367);
nand U7613 (N_7613,N_4413,N_926);
nor U7614 (N_7614,N_4653,N_1613);
or U7615 (N_7615,N_1478,N_1551);
nor U7616 (N_7616,N_2009,N_3302);
nor U7617 (N_7617,N_1161,N_1466);
nor U7618 (N_7618,N_3175,N_3168);
nand U7619 (N_7619,N_341,N_947);
or U7620 (N_7620,N_2143,N_3467);
or U7621 (N_7621,N_195,N_3634);
and U7622 (N_7622,N_4455,N_237);
or U7623 (N_7623,N_4626,N_182);
or U7624 (N_7624,N_3187,N_718);
or U7625 (N_7625,N_3625,N_2010);
nor U7626 (N_7626,N_1295,N_2612);
or U7627 (N_7627,N_2358,N_3259);
and U7628 (N_7628,N_2076,N_2438);
and U7629 (N_7629,N_285,N_1348);
or U7630 (N_7630,N_4821,N_1147);
nor U7631 (N_7631,N_1421,N_3837);
xor U7632 (N_7632,N_3036,N_68);
or U7633 (N_7633,N_1781,N_4734);
xnor U7634 (N_7634,N_2331,N_184);
or U7635 (N_7635,N_255,N_3757);
nand U7636 (N_7636,N_620,N_3431);
and U7637 (N_7637,N_2182,N_2753);
nand U7638 (N_7638,N_1557,N_2901);
or U7639 (N_7639,N_2777,N_1495);
nand U7640 (N_7640,N_4033,N_4557);
or U7641 (N_7641,N_3439,N_330);
nor U7642 (N_7642,N_1695,N_3778);
or U7643 (N_7643,N_1666,N_1935);
nand U7644 (N_7644,N_1930,N_4521);
and U7645 (N_7645,N_3351,N_4691);
and U7646 (N_7646,N_4225,N_3610);
nand U7647 (N_7647,N_4327,N_2812);
nand U7648 (N_7648,N_4867,N_2893);
or U7649 (N_7649,N_1540,N_1230);
and U7650 (N_7650,N_1164,N_4839);
and U7651 (N_7651,N_1244,N_1819);
nand U7652 (N_7652,N_3513,N_3172);
and U7653 (N_7653,N_4207,N_208);
and U7654 (N_7654,N_9,N_4763);
nand U7655 (N_7655,N_2895,N_1117);
and U7656 (N_7656,N_3263,N_1605);
nand U7657 (N_7657,N_1963,N_1585);
or U7658 (N_7658,N_4080,N_4431);
or U7659 (N_7659,N_1535,N_370);
and U7660 (N_7660,N_4553,N_440);
and U7661 (N_7661,N_4606,N_2515);
or U7662 (N_7662,N_3044,N_2719);
nand U7663 (N_7663,N_4891,N_2350);
and U7664 (N_7664,N_4494,N_1678);
nor U7665 (N_7665,N_4709,N_1223);
or U7666 (N_7666,N_1474,N_4811);
or U7667 (N_7667,N_2086,N_3303);
and U7668 (N_7668,N_2227,N_1970);
nand U7669 (N_7669,N_944,N_3536);
nor U7670 (N_7670,N_3875,N_4171);
nand U7671 (N_7671,N_460,N_4279);
nand U7672 (N_7672,N_4005,N_3372);
nor U7673 (N_7673,N_2213,N_747);
and U7674 (N_7674,N_4228,N_1653);
and U7675 (N_7675,N_2637,N_3101);
nor U7676 (N_7676,N_2703,N_407);
or U7677 (N_7677,N_2234,N_4491);
or U7678 (N_7678,N_2692,N_3696);
nand U7679 (N_7679,N_3255,N_966);
nor U7680 (N_7680,N_2063,N_608);
and U7681 (N_7681,N_2689,N_2048);
or U7682 (N_7682,N_104,N_143);
or U7683 (N_7683,N_3193,N_4133);
nand U7684 (N_7684,N_3013,N_4686);
nand U7685 (N_7685,N_2665,N_3065);
or U7686 (N_7686,N_4884,N_4141);
or U7687 (N_7687,N_873,N_2093);
nand U7688 (N_7688,N_2979,N_2820);
or U7689 (N_7689,N_4333,N_2962);
or U7690 (N_7690,N_4045,N_520);
nand U7691 (N_7691,N_4190,N_507);
and U7692 (N_7692,N_2876,N_1029);
or U7693 (N_7693,N_702,N_2538);
and U7694 (N_7694,N_3973,N_594);
or U7695 (N_7695,N_3281,N_2199);
nand U7696 (N_7696,N_946,N_2607);
xor U7697 (N_7697,N_3185,N_1069);
nor U7698 (N_7698,N_300,N_4731);
nand U7699 (N_7699,N_691,N_982);
and U7700 (N_7700,N_4208,N_1961);
nor U7701 (N_7701,N_1265,N_298);
and U7702 (N_7702,N_4224,N_1546);
and U7703 (N_7703,N_488,N_1019);
nand U7704 (N_7704,N_562,N_4460);
nor U7705 (N_7705,N_1771,N_3732);
nor U7706 (N_7706,N_2249,N_807);
nand U7707 (N_7707,N_31,N_2621);
or U7708 (N_7708,N_4751,N_1663);
nor U7709 (N_7709,N_1596,N_2832);
nor U7710 (N_7710,N_603,N_2520);
or U7711 (N_7711,N_2231,N_766);
and U7712 (N_7712,N_2346,N_1648);
nor U7713 (N_7713,N_1356,N_4469);
or U7714 (N_7714,N_4274,N_2007);
and U7715 (N_7715,N_3364,N_4986);
nand U7716 (N_7716,N_4416,N_3866);
and U7717 (N_7717,N_1745,N_2107);
nand U7718 (N_7718,N_1950,N_999);
nor U7719 (N_7719,N_2347,N_3099);
xnor U7720 (N_7720,N_4945,N_2705);
nand U7721 (N_7721,N_2843,N_372);
or U7722 (N_7722,N_2197,N_4021);
or U7723 (N_7723,N_211,N_374);
or U7724 (N_7724,N_2436,N_1195);
xnor U7725 (N_7725,N_3245,N_2310);
nand U7726 (N_7726,N_280,N_3539);
and U7727 (N_7727,N_3460,N_4731);
nor U7728 (N_7728,N_3926,N_4425);
or U7729 (N_7729,N_2342,N_4142);
xnor U7730 (N_7730,N_3958,N_2622);
or U7731 (N_7731,N_4639,N_1646);
and U7732 (N_7732,N_2060,N_1971);
nor U7733 (N_7733,N_443,N_2614);
nand U7734 (N_7734,N_2192,N_4908);
or U7735 (N_7735,N_4503,N_615);
or U7736 (N_7736,N_404,N_4477);
nand U7737 (N_7737,N_895,N_3404);
nor U7738 (N_7738,N_959,N_3136);
nand U7739 (N_7739,N_639,N_2416);
or U7740 (N_7740,N_2747,N_1134);
and U7741 (N_7741,N_2851,N_2581);
nand U7742 (N_7742,N_4552,N_2472);
or U7743 (N_7743,N_2633,N_2532);
or U7744 (N_7744,N_3742,N_1724);
or U7745 (N_7745,N_3332,N_924);
or U7746 (N_7746,N_4094,N_4835);
or U7747 (N_7747,N_2208,N_2470);
or U7748 (N_7748,N_4354,N_1854);
or U7749 (N_7749,N_347,N_3673);
or U7750 (N_7750,N_4299,N_4978);
and U7751 (N_7751,N_3609,N_4061);
and U7752 (N_7752,N_4576,N_3800);
and U7753 (N_7753,N_139,N_3467);
nand U7754 (N_7754,N_2133,N_126);
nor U7755 (N_7755,N_58,N_3223);
and U7756 (N_7756,N_4044,N_4577);
and U7757 (N_7757,N_1339,N_1276);
nand U7758 (N_7758,N_3723,N_3804);
and U7759 (N_7759,N_4390,N_87);
nand U7760 (N_7760,N_4169,N_3879);
or U7761 (N_7761,N_3352,N_209);
and U7762 (N_7762,N_4666,N_2369);
nand U7763 (N_7763,N_661,N_345);
or U7764 (N_7764,N_2611,N_4241);
and U7765 (N_7765,N_3434,N_3419);
and U7766 (N_7766,N_3876,N_3344);
nand U7767 (N_7767,N_2168,N_1658);
or U7768 (N_7768,N_1035,N_4057);
nand U7769 (N_7769,N_1471,N_706);
or U7770 (N_7770,N_1221,N_2985);
xor U7771 (N_7771,N_3064,N_4811);
or U7772 (N_7772,N_905,N_4105);
nor U7773 (N_7773,N_4274,N_2531);
and U7774 (N_7774,N_1410,N_2782);
or U7775 (N_7775,N_4758,N_4528);
nand U7776 (N_7776,N_1471,N_2610);
or U7777 (N_7777,N_1224,N_188);
or U7778 (N_7778,N_3415,N_2815);
nor U7779 (N_7779,N_666,N_979);
nand U7780 (N_7780,N_2177,N_2108);
or U7781 (N_7781,N_1365,N_485);
nor U7782 (N_7782,N_3782,N_2345);
nand U7783 (N_7783,N_838,N_4181);
or U7784 (N_7784,N_2380,N_2144);
nand U7785 (N_7785,N_1243,N_2161);
and U7786 (N_7786,N_2012,N_2245);
and U7787 (N_7787,N_1771,N_3028);
nand U7788 (N_7788,N_4952,N_2652);
nand U7789 (N_7789,N_2371,N_4293);
and U7790 (N_7790,N_4420,N_187);
and U7791 (N_7791,N_3932,N_2632);
nand U7792 (N_7792,N_2583,N_4765);
nand U7793 (N_7793,N_1325,N_3560);
nand U7794 (N_7794,N_2154,N_1361);
nor U7795 (N_7795,N_4426,N_2636);
or U7796 (N_7796,N_4639,N_328);
and U7797 (N_7797,N_128,N_2683);
xnor U7798 (N_7798,N_2726,N_3401);
nand U7799 (N_7799,N_3531,N_4849);
or U7800 (N_7800,N_4664,N_3122);
and U7801 (N_7801,N_2580,N_1121);
nor U7802 (N_7802,N_53,N_721);
and U7803 (N_7803,N_2510,N_1651);
or U7804 (N_7804,N_2110,N_2902);
or U7805 (N_7805,N_3146,N_2180);
nor U7806 (N_7806,N_4199,N_4185);
and U7807 (N_7807,N_1325,N_320);
nand U7808 (N_7808,N_2288,N_2143);
xnor U7809 (N_7809,N_1456,N_3938);
nor U7810 (N_7810,N_4026,N_4604);
and U7811 (N_7811,N_702,N_2487);
or U7812 (N_7812,N_1262,N_1276);
and U7813 (N_7813,N_511,N_1543);
and U7814 (N_7814,N_4644,N_4610);
nand U7815 (N_7815,N_1900,N_4649);
nand U7816 (N_7816,N_183,N_644);
nor U7817 (N_7817,N_3657,N_289);
nor U7818 (N_7818,N_2468,N_4212);
or U7819 (N_7819,N_1036,N_2203);
nand U7820 (N_7820,N_1397,N_2623);
or U7821 (N_7821,N_2910,N_2348);
and U7822 (N_7822,N_1244,N_3064);
or U7823 (N_7823,N_1977,N_4249);
nand U7824 (N_7824,N_4788,N_2311);
or U7825 (N_7825,N_974,N_3314);
or U7826 (N_7826,N_2408,N_2701);
or U7827 (N_7827,N_2723,N_2536);
nand U7828 (N_7828,N_2525,N_4717);
and U7829 (N_7829,N_1752,N_2267);
nor U7830 (N_7830,N_4893,N_4515);
or U7831 (N_7831,N_4052,N_1313);
nand U7832 (N_7832,N_1872,N_1052);
nor U7833 (N_7833,N_132,N_4995);
or U7834 (N_7834,N_3214,N_172);
nand U7835 (N_7835,N_2886,N_61);
nand U7836 (N_7836,N_974,N_3827);
nand U7837 (N_7837,N_1857,N_856);
or U7838 (N_7838,N_4525,N_1068);
nor U7839 (N_7839,N_2627,N_4522);
and U7840 (N_7840,N_4577,N_480);
nor U7841 (N_7841,N_3865,N_1103);
nor U7842 (N_7842,N_938,N_3078);
or U7843 (N_7843,N_4879,N_3641);
or U7844 (N_7844,N_3472,N_973);
or U7845 (N_7845,N_2386,N_1820);
nand U7846 (N_7846,N_1716,N_3360);
or U7847 (N_7847,N_477,N_1562);
and U7848 (N_7848,N_2175,N_1974);
nor U7849 (N_7849,N_4340,N_3842);
nor U7850 (N_7850,N_203,N_3190);
nor U7851 (N_7851,N_721,N_1283);
and U7852 (N_7852,N_3538,N_2559);
nand U7853 (N_7853,N_743,N_2426);
or U7854 (N_7854,N_385,N_718);
nand U7855 (N_7855,N_4885,N_4076);
and U7856 (N_7856,N_2016,N_605);
xor U7857 (N_7857,N_4555,N_4066);
nand U7858 (N_7858,N_940,N_2782);
nand U7859 (N_7859,N_2317,N_3349);
nor U7860 (N_7860,N_2298,N_2283);
xor U7861 (N_7861,N_1483,N_841);
or U7862 (N_7862,N_865,N_115);
or U7863 (N_7863,N_3485,N_3490);
xnor U7864 (N_7864,N_2145,N_2767);
and U7865 (N_7865,N_3636,N_2219);
nand U7866 (N_7866,N_3569,N_1237);
nand U7867 (N_7867,N_4186,N_3975);
nand U7868 (N_7868,N_880,N_709);
or U7869 (N_7869,N_560,N_3441);
nand U7870 (N_7870,N_3297,N_1930);
nor U7871 (N_7871,N_2548,N_3498);
nor U7872 (N_7872,N_3024,N_2698);
or U7873 (N_7873,N_2810,N_4268);
nor U7874 (N_7874,N_569,N_2773);
nand U7875 (N_7875,N_1750,N_3013);
nor U7876 (N_7876,N_1053,N_3600);
and U7877 (N_7877,N_4177,N_366);
nand U7878 (N_7878,N_1101,N_3355);
or U7879 (N_7879,N_3281,N_3199);
or U7880 (N_7880,N_3727,N_1385);
or U7881 (N_7881,N_421,N_3257);
nand U7882 (N_7882,N_3177,N_3900);
or U7883 (N_7883,N_2119,N_4174);
or U7884 (N_7884,N_1859,N_1326);
or U7885 (N_7885,N_4937,N_854);
and U7886 (N_7886,N_1234,N_1219);
and U7887 (N_7887,N_850,N_3809);
nor U7888 (N_7888,N_1557,N_4766);
or U7889 (N_7889,N_4839,N_1075);
nand U7890 (N_7890,N_4182,N_2765);
nand U7891 (N_7891,N_1169,N_4676);
nand U7892 (N_7892,N_2084,N_3246);
nor U7893 (N_7893,N_3010,N_4321);
xor U7894 (N_7894,N_504,N_372);
nor U7895 (N_7895,N_3940,N_521);
and U7896 (N_7896,N_1287,N_1396);
nand U7897 (N_7897,N_1768,N_363);
or U7898 (N_7898,N_2644,N_4191);
and U7899 (N_7899,N_3773,N_2538);
nor U7900 (N_7900,N_2390,N_3245);
nand U7901 (N_7901,N_3891,N_1743);
nand U7902 (N_7902,N_3562,N_1467);
nand U7903 (N_7903,N_1901,N_939);
and U7904 (N_7904,N_4610,N_258);
nand U7905 (N_7905,N_1202,N_2328);
nand U7906 (N_7906,N_1139,N_3437);
and U7907 (N_7907,N_2398,N_3688);
or U7908 (N_7908,N_1350,N_514);
and U7909 (N_7909,N_3566,N_4350);
nor U7910 (N_7910,N_4591,N_1812);
or U7911 (N_7911,N_2372,N_4667);
and U7912 (N_7912,N_4183,N_3174);
nand U7913 (N_7913,N_1405,N_2315);
nand U7914 (N_7914,N_1139,N_2332);
nor U7915 (N_7915,N_4985,N_3795);
nor U7916 (N_7916,N_3144,N_621);
and U7917 (N_7917,N_4908,N_2653);
nand U7918 (N_7918,N_4960,N_1353);
or U7919 (N_7919,N_3591,N_2856);
or U7920 (N_7920,N_3429,N_3134);
nor U7921 (N_7921,N_3839,N_115);
or U7922 (N_7922,N_1262,N_361);
nand U7923 (N_7923,N_3284,N_218);
or U7924 (N_7924,N_1099,N_3213);
xor U7925 (N_7925,N_1205,N_2910);
nor U7926 (N_7926,N_2068,N_1725);
and U7927 (N_7927,N_383,N_173);
and U7928 (N_7928,N_4572,N_4093);
nor U7929 (N_7929,N_2925,N_3304);
or U7930 (N_7930,N_3890,N_2093);
or U7931 (N_7931,N_2831,N_3855);
and U7932 (N_7932,N_465,N_984);
nand U7933 (N_7933,N_106,N_2105);
nor U7934 (N_7934,N_1149,N_3623);
nand U7935 (N_7935,N_1530,N_4658);
nand U7936 (N_7936,N_4751,N_3027);
nand U7937 (N_7937,N_4691,N_2956);
nor U7938 (N_7938,N_173,N_862);
nand U7939 (N_7939,N_3561,N_165);
or U7940 (N_7940,N_861,N_4243);
nand U7941 (N_7941,N_674,N_2115);
nand U7942 (N_7942,N_535,N_1612);
or U7943 (N_7943,N_70,N_1707);
nor U7944 (N_7944,N_3121,N_4251);
and U7945 (N_7945,N_4447,N_3876);
nand U7946 (N_7946,N_3707,N_3465);
xor U7947 (N_7947,N_2473,N_3947);
or U7948 (N_7948,N_928,N_2569);
nand U7949 (N_7949,N_2525,N_181);
and U7950 (N_7950,N_3844,N_559);
or U7951 (N_7951,N_1055,N_2464);
or U7952 (N_7952,N_4250,N_1054);
and U7953 (N_7953,N_3011,N_2211);
nand U7954 (N_7954,N_2901,N_4119);
or U7955 (N_7955,N_4522,N_3289);
nor U7956 (N_7956,N_3999,N_138);
nor U7957 (N_7957,N_232,N_385);
or U7958 (N_7958,N_4426,N_2571);
and U7959 (N_7959,N_296,N_2805);
nor U7960 (N_7960,N_1999,N_4972);
or U7961 (N_7961,N_4564,N_4517);
or U7962 (N_7962,N_47,N_933);
nor U7963 (N_7963,N_345,N_3686);
nor U7964 (N_7964,N_2288,N_1123);
nor U7965 (N_7965,N_2711,N_2803);
nor U7966 (N_7966,N_1032,N_3510);
or U7967 (N_7967,N_4901,N_1331);
nand U7968 (N_7968,N_1021,N_1297);
or U7969 (N_7969,N_2068,N_3657);
nor U7970 (N_7970,N_274,N_3398);
nor U7971 (N_7971,N_972,N_3394);
nand U7972 (N_7972,N_4694,N_3086);
nor U7973 (N_7973,N_176,N_1953);
nor U7974 (N_7974,N_933,N_4787);
and U7975 (N_7975,N_2592,N_1739);
nor U7976 (N_7976,N_1646,N_3524);
nand U7977 (N_7977,N_558,N_3022);
and U7978 (N_7978,N_798,N_3624);
or U7979 (N_7979,N_1338,N_464);
and U7980 (N_7980,N_2354,N_2268);
nand U7981 (N_7981,N_3591,N_3157);
nand U7982 (N_7982,N_2068,N_4142);
nand U7983 (N_7983,N_2528,N_4911);
and U7984 (N_7984,N_3744,N_218);
and U7985 (N_7985,N_3433,N_2767);
or U7986 (N_7986,N_3335,N_1452);
xor U7987 (N_7987,N_2012,N_2602);
nor U7988 (N_7988,N_3244,N_1645);
and U7989 (N_7989,N_2290,N_221);
nor U7990 (N_7990,N_4168,N_321);
nand U7991 (N_7991,N_4379,N_4924);
nand U7992 (N_7992,N_1409,N_462);
nand U7993 (N_7993,N_472,N_3346);
nor U7994 (N_7994,N_182,N_4431);
or U7995 (N_7995,N_2365,N_4068);
nand U7996 (N_7996,N_3895,N_2539);
nor U7997 (N_7997,N_2116,N_1042);
nand U7998 (N_7998,N_4223,N_2516);
and U7999 (N_7999,N_3561,N_3542);
or U8000 (N_8000,N_795,N_3301);
nand U8001 (N_8001,N_4922,N_4230);
and U8002 (N_8002,N_1420,N_4473);
and U8003 (N_8003,N_2555,N_391);
nand U8004 (N_8004,N_2008,N_4730);
nand U8005 (N_8005,N_3958,N_3073);
and U8006 (N_8006,N_4582,N_371);
and U8007 (N_8007,N_440,N_4873);
nor U8008 (N_8008,N_1867,N_1424);
or U8009 (N_8009,N_4985,N_3267);
and U8010 (N_8010,N_3888,N_3007);
and U8011 (N_8011,N_4374,N_1466);
nand U8012 (N_8012,N_3803,N_2859);
nor U8013 (N_8013,N_1452,N_4067);
and U8014 (N_8014,N_1864,N_2723);
or U8015 (N_8015,N_351,N_1713);
and U8016 (N_8016,N_3024,N_1271);
nor U8017 (N_8017,N_1387,N_1888);
and U8018 (N_8018,N_19,N_3571);
and U8019 (N_8019,N_513,N_2400);
nand U8020 (N_8020,N_1437,N_891);
nor U8021 (N_8021,N_3160,N_1147);
and U8022 (N_8022,N_3899,N_1928);
nand U8023 (N_8023,N_1157,N_498);
xnor U8024 (N_8024,N_3044,N_955);
nor U8025 (N_8025,N_843,N_2674);
nand U8026 (N_8026,N_4289,N_1982);
nand U8027 (N_8027,N_2596,N_660);
or U8028 (N_8028,N_3,N_4375);
nand U8029 (N_8029,N_984,N_2574);
nand U8030 (N_8030,N_1732,N_2599);
nand U8031 (N_8031,N_1979,N_4939);
nor U8032 (N_8032,N_3300,N_4164);
and U8033 (N_8033,N_4656,N_3074);
or U8034 (N_8034,N_3481,N_3294);
and U8035 (N_8035,N_3727,N_1553);
nand U8036 (N_8036,N_436,N_617);
nor U8037 (N_8037,N_4903,N_4411);
and U8038 (N_8038,N_1630,N_2475);
or U8039 (N_8039,N_4348,N_2335);
and U8040 (N_8040,N_1608,N_4340);
nor U8041 (N_8041,N_1856,N_3892);
nand U8042 (N_8042,N_1145,N_1758);
or U8043 (N_8043,N_1848,N_2450);
nor U8044 (N_8044,N_2127,N_4064);
nand U8045 (N_8045,N_3479,N_2103);
nor U8046 (N_8046,N_2166,N_4002);
nand U8047 (N_8047,N_2947,N_1738);
or U8048 (N_8048,N_2169,N_2322);
nand U8049 (N_8049,N_359,N_2817);
nor U8050 (N_8050,N_2663,N_3235);
nand U8051 (N_8051,N_1735,N_3554);
nand U8052 (N_8052,N_4915,N_4639);
nand U8053 (N_8053,N_1817,N_1271);
or U8054 (N_8054,N_487,N_467);
or U8055 (N_8055,N_217,N_1071);
xnor U8056 (N_8056,N_1594,N_1389);
or U8057 (N_8057,N_3924,N_1307);
nand U8058 (N_8058,N_735,N_868);
nand U8059 (N_8059,N_1451,N_4044);
or U8060 (N_8060,N_3434,N_1388);
and U8061 (N_8061,N_3016,N_1502);
nor U8062 (N_8062,N_1368,N_4762);
nand U8063 (N_8063,N_3878,N_4180);
or U8064 (N_8064,N_4650,N_4857);
or U8065 (N_8065,N_2367,N_2114);
or U8066 (N_8066,N_3273,N_3667);
and U8067 (N_8067,N_2098,N_1567);
or U8068 (N_8068,N_1935,N_2141);
nor U8069 (N_8069,N_1637,N_2727);
and U8070 (N_8070,N_1216,N_664);
nor U8071 (N_8071,N_1010,N_543);
and U8072 (N_8072,N_521,N_3418);
nand U8073 (N_8073,N_4110,N_2912);
xnor U8074 (N_8074,N_72,N_342);
nor U8075 (N_8075,N_1285,N_2115);
nand U8076 (N_8076,N_538,N_229);
and U8077 (N_8077,N_2068,N_4901);
and U8078 (N_8078,N_948,N_1429);
nor U8079 (N_8079,N_4322,N_3772);
nor U8080 (N_8080,N_4869,N_4282);
or U8081 (N_8081,N_2713,N_4748);
nand U8082 (N_8082,N_3638,N_4974);
or U8083 (N_8083,N_77,N_4940);
or U8084 (N_8084,N_3395,N_336);
and U8085 (N_8085,N_4125,N_3230);
or U8086 (N_8086,N_198,N_346);
nand U8087 (N_8087,N_1422,N_4229);
or U8088 (N_8088,N_1525,N_4832);
nand U8089 (N_8089,N_3732,N_3023);
nor U8090 (N_8090,N_4239,N_2843);
or U8091 (N_8091,N_1761,N_907);
and U8092 (N_8092,N_3303,N_1495);
or U8093 (N_8093,N_1368,N_4152);
or U8094 (N_8094,N_978,N_2054);
or U8095 (N_8095,N_526,N_403);
nand U8096 (N_8096,N_2045,N_1065);
xnor U8097 (N_8097,N_857,N_2509);
nand U8098 (N_8098,N_2417,N_1044);
and U8099 (N_8099,N_1074,N_59);
nand U8100 (N_8100,N_120,N_2634);
nor U8101 (N_8101,N_3207,N_1959);
nand U8102 (N_8102,N_628,N_2081);
nand U8103 (N_8103,N_1399,N_3281);
nand U8104 (N_8104,N_4702,N_3672);
or U8105 (N_8105,N_69,N_926);
and U8106 (N_8106,N_3055,N_3376);
nor U8107 (N_8107,N_2384,N_3645);
nand U8108 (N_8108,N_3584,N_4589);
or U8109 (N_8109,N_900,N_2263);
nand U8110 (N_8110,N_3390,N_4428);
nor U8111 (N_8111,N_2390,N_1708);
xor U8112 (N_8112,N_377,N_639);
or U8113 (N_8113,N_62,N_3540);
and U8114 (N_8114,N_154,N_2143);
or U8115 (N_8115,N_4334,N_2461);
or U8116 (N_8116,N_4565,N_757);
or U8117 (N_8117,N_241,N_3143);
nand U8118 (N_8118,N_1421,N_2436);
and U8119 (N_8119,N_3112,N_1041);
and U8120 (N_8120,N_254,N_1989);
or U8121 (N_8121,N_1017,N_4688);
nor U8122 (N_8122,N_3886,N_4524);
nand U8123 (N_8123,N_928,N_864);
nand U8124 (N_8124,N_1847,N_2268);
or U8125 (N_8125,N_4708,N_554);
nor U8126 (N_8126,N_227,N_844);
and U8127 (N_8127,N_1102,N_1945);
or U8128 (N_8128,N_1097,N_2882);
or U8129 (N_8129,N_2484,N_4741);
or U8130 (N_8130,N_4614,N_336);
nor U8131 (N_8131,N_4751,N_4421);
nand U8132 (N_8132,N_2885,N_1564);
or U8133 (N_8133,N_3172,N_2514);
nand U8134 (N_8134,N_2025,N_1748);
nand U8135 (N_8135,N_2588,N_3273);
and U8136 (N_8136,N_4033,N_1035);
nor U8137 (N_8137,N_1459,N_4089);
nand U8138 (N_8138,N_1282,N_1613);
and U8139 (N_8139,N_2038,N_1367);
nor U8140 (N_8140,N_2009,N_1448);
nand U8141 (N_8141,N_3472,N_1860);
nand U8142 (N_8142,N_4673,N_3864);
nor U8143 (N_8143,N_2238,N_1137);
and U8144 (N_8144,N_3567,N_4393);
and U8145 (N_8145,N_3777,N_1913);
and U8146 (N_8146,N_4985,N_2486);
nand U8147 (N_8147,N_2254,N_2825);
nor U8148 (N_8148,N_2749,N_577);
or U8149 (N_8149,N_2374,N_2667);
and U8150 (N_8150,N_4014,N_4161);
nand U8151 (N_8151,N_1252,N_1013);
or U8152 (N_8152,N_1546,N_1202);
or U8153 (N_8153,N_3843,N_853);
and U8154 (N_8154,N_3477,N_2231);
and U8155 (N_8155,N_4390,N_3797);
nor U8156 (N_8156,N_1300,N_3536);
or U8157 (N_8157,N_59,N_3097);
or U8158 (N_8158,N_3908,N_1791);
nand U8159 (N_8159,N_4928,N_2164);
nor U8160 (N_8160,N_734,N_3506);
or U8161 (N_8161,N_691,N_1921);
and U8162 (N_8162,N_365,N_4611);
or U8163 (N_8163,N_1628,N_1452);
xnor U8164 (N_8164,N_3501,N_3989);
and U8165 (N_8165,N_1690,N_3582);
nand U8166 (N_8166,N_762,N_4366);
and U8167 (N_8167,N_116,N_801);
nand U8168 (N_8168,N_2578,N_4638);
nor U8169 (N_8169,N_4921,N_3808);
or U8170 (N_8170,N_3939,N_1924);
nand U8171 (N_8171,N_4344,N_3377);
nor U8172 (N_8172,N_2759,N_2452);
nor U8173 (N_8173,N_586,N_4767);
nand U8174 (N_8174,N_2088,N_4137);
nand U8175 (N_8175,N_2207,N_2841);
nor U8176 (N_8176,N_1768,N_3942);
nor U8177 (N_8177,N_1349,N_1359);
or U8178 (N_8178,N_1996,N_4962);
or U8179 (N_8179,N_4666,N_2360);
or U8180 (N_8180,N_802,N_1399);
or U8181 (N_8181,N_4348,N_441);
nor U8182 (N_8182,N_949,N_3636);
nand U8183 (N_8183,N_3267,N_3517);
nand U8184 (N_8184,N_790,N_146);
nor U8185 (N_8185,N_2347,N_4173);
nor U8186 (N_8186,N_3590,N_1213);
nand U8187 (N_8187,N_4696,N_135);
nand U8188 (N_8188,N_3347,N_3613);
nand U8189 (N_8189,N_2217,N_3302);
nor U8190 (N_8190,N_4871,N_1735);
and U8191 (N_8191,N_2648,N_2137);
and U8192 (N_8192,N_3272,N_1106);
nand U8193 (N_8193,N_4420,N_3796);
nand U8194 (N_8194,N_1596,N_838);
nor U8195 (N_8195,N_4430,N_3474);
and U8196 (N_8196,N_1221,N_2849);
or U8197 (N_8197,N_935,N_576);
nand U8198 (N_8198,N_1364,N_1572);
nor U8199 (N_8199,N_500,N_1049);
and U8200 (N_8200,N_1544,N_1248);
and U8201 (N_8201,N_4435,N_4671);
nor U8202 (N_8202,N_3359,N_159);
xnor U8203 (N_8203,N_3868,N_4685);
and U8204 (N_8204,N_875,N_4602);
nand U8205 (N_8205,N_648,N_3736);
or U8206 (N_8206,N_2735,N_280);
nor U8207 (N_8207,N_1236,N_1617);
nand U8208 (N_8208,N_4188,N_3399);
or U8209 (N_8209,N_2677,N_825);
and U8210 (N_8210,N_1038,N_2991);
nand U8211 (N_8211,N_2269,N_645);
nor U8212 (N_8212,N_1633,N_1860);
and U8213 (N_8213,N_4324,N_1357);
or U8214 (N_8214,N_1018,N_3587);
nand U8215 (N_8215,N_333,N_1412);
or U8216 (N_8216,N_2957,N_2517);
nand U8217 (N_8217,N_272,N_3707);
and U8218 (N_8218,N_3437,N_2733);
and U8219 (N_8219,N_4956,N_3009);
nor U8220 (N_8220,N_1651,N_2468);
nand U8221 (N_8221,N_4988,N_3906);
or U8222 (N_8222,N_4209,N_2092);
nand U8223 (N_8223,N_3042,N_3125);
nand U8224 (N_8224,N_3732,N_2667);
nor U8225 (N_8225,N_1394,N_1951);
and U8226 (N_8226,N_246,N_1237);
nand U8227 (N_8227,N_3279,N_4329);
and U8228 (N_8228,N_1664,N_3699);
or U8229 (N_8229,N_3950,N_2015);
and U8230 (N_8230,N_3572,N_3600);
and U8231 (N_8231,N_3052,N_1486);
nor U8232 (N_8232,N_3222,N_1611);
nand U8233 (N_8233,N_4330,N_1556);
nor U8234 (N_8234,N_2906,N_772);
nand U8235 (N_8235,N_3919,N_4109);
nand U8236 (N_8236,N_2063,N_2822);
and U8237 (N_8237,N_434,N_56);
or U8238 (N_8238,N_44,N_497);
nor U8239 (N_8239,N_1588,N_4817);
or U8240 (N_8240,N_372,N_2566);
and U8241 (N_8241,N_3943,N_129);
nor U8242 (N_8242,N_1164,N_1463);
and U8243 (N_8243,N_4922,N_644);
nand U8244 (N_8244,N_1095,N_3395);
nor U8245 (N_8245,N_1466,N_490);
nor U8246 (N_8246,N_2707,N_3172);
nor U8247 (N_8247,N_1389,N_623);
or U8248 (N_8248,N_2828,N_1450);
and U8249 (N_8249,N_2446,N_463);
nand U8250 (N_8250,N_2306,N_4455);
nor U8251 (N_8251,N_2082,N_3456);
or U8252 (N_8252,N_205,N_1941);
or U8253 (N_8253,N_3656,N_1120);
nor U8254 (N_8254,N_3406,N_4555);
nor U8255 (N_8255,N_1494,N_4661);
or U8256 (N_8256,N_2190,N_311);
nand U8257 (N_8257,N_3801,N_2693);
or U8258 (N_8258,N_1151,N_3614);
or U8259 (N_8259,N_1017,N_3811);
xor U8260 (N_8260,N_3580,N_3391);
and U8261 (N_8261,N_3976,N_2747);
and U8262 (N_8262,N_1784,N_1726);
xor U8263 (N_8263,N_4125,N_195);
xor U8264 (N_8264,N_782,N_381);
and U8265 (N_8265,N_4494,N_709);
nor U8266 (N_8266,N_3347,N_2735);
and U8267 (N_8267,N_4142,N_4724);
and U8268 (N_8268,N_1874,N_1094);
nor U8269 (N_8269,N_2682,N_4922);
and U8270 (N_8270,N_3752,N_2352);
and U8271 (N_8271,N_4228,N_4726);
nor U8272 (N_8272,N_2026,N_4517);
nand U8273 (N_8273,N_4050,N_279);
nor U8274 (N_8274,N_932,N_3789);
nand U8275 (N_8275,N_676,N_2807);
nor U8276 (N_8276,N_423,N_560);
nor U8277 (N_8277,N_4706,N_3805);
nand U8278 (N_8278,N_878,N_2454);
nor U8279 (N_8279,N_553,N_1611);
nand U8280 (N_8280,N_1723,N_4260);
nor U8281 (N_8281,N_3358,N_3615);
and U8282 (N_8282,N_4332,N_540);
and U8283 (N_8283,N_1001,N_932);
xor U8284 (N_8284,N_3314,N_4984);
or U8285 (N_8285,N_1987,N_2033);
and U8286 (N_8286,N_2646,N_4024);
nor U8287 (N_8287,N_1719,N_4663);
and U8288 (N_8288,N_812,N_4223);
nor U8289 (N_8289,N_1114,N_272);
or U8290 (N_8290,N_4476,N_1586);
and U8291 (N_8291,N_882,N_4686);
nor U8292 (N_8292,N_121,N_2603);
nor U8293 (N_8293,N_4504,N_2243);
and U8294 (N_8294,N_3162,N_3187);
or U8295 (N_8295,N_533,N_877);
or U8296 (N_8296,N_3911,N_3385);
nand U8297 (N_8297,N_1288,N_2127);
and U8298 (N_8298,N_3979,N_4470);
or U8299 (N_8299,N_4670,N_216);
and U8300 (N_8300,N_1228,N_3813);
nor U8301 (N_8301,N_4359,N_1866);
nand U8302 (N_8302,N_1278,N_1076);
or U8303 (N_8303,N_4892,N_3717);
nor U8304 (N_8304,N_4846,N_714);
nor U8305 (N_8305,N_812,N_1471);
nand U8306 (N_8306,N_4768,N_4294);
and U8307 (N_8307,N_4785,N_3735);
nor U8308 (N_8308,N_125,N_855);
nand U8309 (N_8309,N_3005,N_935);
nor U8310 (N_8310,N_2866,N_3415);
nor U8311 (N_8311,N_8,N_601);
nor U8312 (N_8312,N_4951,N_2253);
and U8313 (N_8313,N_2343,N_2629);
or U8314 (N_8314,N_822,N_333);
and U8315 (N_8315,N_4207,N_2166);
and U8316 (N_8316,N_248,N_2510);
and U8317 (N_8317,N_2895,N_2874);
or U8318 (N_8318,N_1977,N_1462);
and U8319 (N_8319,N_3366,N_3085);
nor U8320 (N_8320,N_263,N_3017);
nor U8321 (N_8321,N_192,N_390);
nand U8322 (N_8322,N_4180,N_3836);
nor U8323 (N_8323,N_1663,N_642);
or U8324 (N_8324,N_431,N_692);
xnor U8325 (N_8325,N_4864,N_2802);
nor U8326 (N_8326,N_2413,N_2133);
and U8327 (N_8327,N_3680,N_4448);
nand U8328 (N_8328,N_2804,N_1033);
and U8329 (N_8329,N_3639,N_1222);
nand U8330 (N_8330,N_2370,N_2944);
nand U8331 (N_8331,N_3975,N_2999);
or U8332 (N_8332,N_687,N_3346);
or U8333 (N_8333,N_3014,N_2874);
and U8334 (N_8334,N_1391,N_490);
or U8335 (N_8335,N_3854,N_2362);
nand U8336 (N_8336,N_2452,N_1394);
nor U8337 (N_8337,N_1130,N_2482);
nand U8338 (N_8338,N_3259,N_3102);
nand U8339 (N_8339,N_2536,N_4073);
nand U8340 (N_8340,N_3960,N_4784);
nand U8341 (N_8341,N_242,N_4191);
or U8342 (N_8342,N_4638,N_315);
nor U8343 (N_8343,N_1412,N_1298);
nor U8344 (N_8344,N_732,N_3162);
or U8345 (N_8345,N_1699,N_4950);
or U8346 (N_8346,N_651,N_458);
or U8347 (N_8347,N_3364,N_1386);
nor U8348 (N_8348,N_1887,N_4263);
or U8349 (N_8349,N_183,N_1805);
and U8350 (N_8350,N_3217,N_1150);
nand U8351 (N_8351,N_2174,N_592);
and U8352 (N_8352,N_4165,N_4132);
nand U8353 (N_8353,N_4109,N_3989);
or U8354 (N_8354,N_3016,N_4288);
or U8355 (N_8355,N_2087,N_1305);
nor U8356 (N_8356,N_3789,N_3934);
or U8357 (N_8357,N_3127,N_3583);
and U8358 (N_8358,N_2140,N_4288);
xor U8359 (N_8359,N_2262,N_1514);
or U8360 (N_8360,N_2021,N_32);
and U8361 (N_8361,N_3595,N_1573);
nor U8362 (N_8362,N_3223,N_101);
nor U8363 (N_8363,N_349,N_1193);
nor U8364 (N_8364,N_1953,N_3757);
nor U8365 (N_8365,N_4828,N_1339);
and U8366 (N_8366,N_2190,N_1944);
and U8367 (N_8367,N_4139,N_1583);
nor U8368 (N_8368,N_4872,N_1916);
nand U8369 (N_8369,N_3215,N_358);
nor U8370 (N_8370,N_2535,N_2295);
nor U8371 (N_8371,N_1849,N_561);
or U8372 (N_8372,N_2572,N_2218);
nand U8373 (N_8373,N_4337,N_123);
nand U8374 (N_8374,N_3993,N_3850);
and U8375 (N_8375,N_560,N_4528);
nand U8376 (N_8376,N_265,N_4372);
nand U8377 (N_8377,N_1069,N_3108);
xnor U8378 (N_8378,N_75,N_4187);
nor U8379 (N_8379,N_1465,N_2453);
or U8380 (N_8380,N_4024,N_2851);
nand U8381 (N_8381,N_3547,N_4329);
nor U8382 (N_8382,N_4845,N_4888);
nor U8383 (N_8383,N_133,N_722);
nor U8384 (N_8384,N_3286,N_4672);
nand U8385 (N_8385,N_1939,N_3599);
nor U8386 (N_8386,N_1150,N_796);
nor U8387 (N_8387,N_1951,N_1247);
nand U8388 (N_8388,N_2312,N_873);
or U8389 (N_8389,N_4961,N_2338);
and U8390 (N_8390,N_3143,N_1003);
and U8391 (N_8391,N_4430,N_1114);
and U8392 (N_8392,N_1101,N_462);
or U8393 (N_8393,N_2972,N_151);
nor U8394 (N_8394,N_3098,N_2522);
nor U8395 (N_8395,N_2417,N_3527);
and U8396 (N_8396,N_1441,N_4160);
or U8397 (N_8397,N_2084,N_1587);
or U8398 (N_8398,N_828,N_160);
or U8399 (N_8399,N_233,N_2504);
and U8400 (N_8400,N_4899,N_41);
nor U8401 (N_8401,N_4726,N_709);
xor U8402 (N_8402,N_1759,N_2004);
or U8403 (N_8403,N_3458,N_1524);
nor U8404 (N_8404,N_4641,N_3108);
or U8405 (N_8405,N_688,N_4453);
or U8406 (N_8406,N_4486,N_4495);
and U8407 (N_8407,N_1104,N_2153);
nand U8408 (N_8408,N_998,N_1003);
and U8409 (N_8409,N_1123,N_602);
nor U8410 (N_8410,N_3507,N_2198);
nor U8411 (N_8411,N_4389,N_2021);
nor U8412 (N_8412,N_4935,N_4139);
nor U8413 (N_8413,N_4420,N_721);
or U8414 (N_8414,N_4917,N_2020);
nand U8415 (N_8415,N_2096,N_1396);
nand U8416 (N_8416,N_986,N_3718);
or U8417 (N_8417,N_3861,N_3477);
and U8418 (N_8418,N_2760,N_1876);
and U8419 (N_8419,N_1448,N_4881);
xor U8420 (N_8420,N_213,N_2901);
nand U8421 (N_8421,N_1114,N_4757);
nand U8422 (N_8422,N_935,N_2823);
nand U8423 (N_8423,N_781,N_4916);
nor U8424 (N_8424,N_48,N_1650);
or U8425 (N_8425,N_1820,N_1138);
and U8426 (N_8426,N_858,N_146);
nand U8427 (N_8427,N_1658,N_3139);
nor U8428 (N_8428,N_3336,N_78);
or U8429 (N_8429,N_860,N_755);
nand U8430 (N_8430,N_2676,N_784);
nor U8431 (N_8431,N_2273,N_1203);
nand U8432 (N_8432,N_138,N_3731);
and U8433 (N_8433,N_753,N_2409);
nand U8434 (N_8434,N_3025,N_2223);
or U8435 (N_8435,N_3222,N_427);
nor U8436 (N_8436,N_968,N_2378);
nand U8437 (N_8437,N_4222,N_3851);
xor U8438 (N_8438,N_679,N_1143);
nand U8439 (N_8439,N_336,N_4988);
nand U8440 (N_8440,N_1613,N_3080);
xnor U8441 (N_8441,N_639,N_3968);
or U8442 (N_8442,N_4908,N_463);
or U8443 (N_8443,N_1712,N_4237);
nand U8444 (N_8444,N_34,N_2998);
and U8445 (N_8445,N_3624,N_526);
or U8446 (N_8446,N_1062,N_3038);
nor U8447 (N_8447,N_4276,N_2733);
nor U8448 (N_8448,N_3025,N_874);
nor U8449 (N_8449,N_2569,N_1482);
nor U8450 (N_8450,N_452,N_3596);
nor U8451 (N_8451,N_721,N_4057);
or U8452 (N_8452,N_1744,N_1449);
nand U8453 (N_8453,N_352,N_3444);
nand U8454 (N_8454,N_1974,N_1279);
or U8455 (N_8455,N_2857,N_797);
nand U8456 (N_8456,N_4718,N_167);
and U8457 (N_8457,N_3749,N_4528);
or U8458 (N_8458,N_210,N_872);
nor U8459 (N_8459,N_1624,N_2860);
nor U8460 (N_8460,N_724,N_4426);
xor U8461 (N_8461,N_4858,N_785);
nand U8462 (N_8462,N_4543,N_4765);
nor U8463 (N_8463,N_2765,N_4883);
or U8464 (N_8464,N_1909,N_4725);
nor U8465 (N_8465,N_1423,N_4731);
nand U8466 (N_8466,N_86,N_1490);
and U8467 (N_8467,N_4758,N_1272);
nor U8468 (N_8468,N_2421,N_2819);
or U8469 (N_8469,N_2112,N_4710);
or U8470 (N_8470,N_2733,N_2056);
nor U8471 (N_8471,N_4077,N_1526);
nand U8472 (N_8472,N_1339,N_403);
or U8473 (N_8473,N_4355,N_4287);
and U8474 (N_8474,N_3780,N_2830);
nand U8475 (N_8475,N_493,N_3078);
or U8476 (N_8476,N_3975,N_4509);
xnor U8477 (N_8477,N_3933,N_2439);
nor U8478 (N_8478,N_2286,N_1832);
and U8479 (N_8479,N_1033,N_2096);
xnor U8480 (N_8480,N_3039,N_4389);
and U8481 (N_8481,N_3751,N_4225);
or U8482 (N_8482,N_945,N_3207);
or U8483 (N_8483,N_4741,N_1954);
and U8484 (N_8484,N_399,N_2051);
nand U8485 (N_8485,N_2143,N_2414);
nor U8486 (N_8486,N_2623,N_603);
and U8487 (N_8487,N_4285,N_1885);
xnor U8488 (N_8488,N_3852,N_2838);
nor U8489 (N_8489,N_1767,N_63);
and U8490 (N_8490,N_4331,N_1879);
nand U8491 (N_8491,N_1872,N_1205);
nor U8492 (N_8492,N_673,N_1741);
xor U8493 (N_8493,N_4598,N_4951);
nand U8494 (N_8494,N_1922,N_2958);
and U8495 (N_8495,N_759,N_3970);
nand U8496 (N_8496,N_3003,N_2346);
and U8497 (N_8497,N_4470,N_4964);
or U8498 (N_8498,N_4893,N_2479);
nand U8499 (N_8499,N_28,N_1479);
nor U8500 (N_8500,N_795,N_4530);
nand U8501 (N_8501,N_282,N_4745);
xor U8502 (N_8502,N_1338,N_683);
nand U8503 (N_8503,N_3902,N_2004);
nor U8504 (N_8504,N_4354,N_1089);
nor U8505 (N_8505,N_3576,N_4651);
and U8506 (N_8506,N_4324,N_4826);
and U8507 (N_8507,N_3142,N_541);
or U8508 (N_8508,N_1401,N_3857);
or U8509 (N_8509,N_3414,N_4139);
and U8510 (N_8510,N_3985,N_1941);
or U8511 (N_8511,N_1078,N_3700);
nand U8512 (N_8512,N_3522,N_3227);
nor U8513 (N_8513,N_2559,N_4656);
nand U8514 (N_8514,N_2660,N_1386);
nand U8515 (N_8515,N_3253,N_2095);
and U8516 (N_8516,N_2770,N_37);
xor U8517 (N_8517,N_2551,N_4794);
nor U8518 (N_8518,N_1774,N_2325);
nor U8519 (N_8519,N_1994,N_4733);
nor U8520 (N_8520,N_972,N_4309);
xor U8521 (N_8521,N_1725,N_1659);
nor U8522 (N_8522,N_3772,N_80);
nor U8523 (N_8523,N_4779,N_4813);
nand U8524 (N_8524,N_2252,N_4799);
nand U8525 (N_8525,N_2854,N_4124);
nand U8526 (N_8526,N_1146,N_997);
or U8527 (N_8527,N_3944,N_404);
nand U8528 (N_8528,N_3097,N_3426);
nand U8529 (N_8529,N_234,N_2826);
nor U8530 (N_8530,N_2648,N_1757);
or U8531 (N_8531,N_2341,N_1335);
nand U8532 (N_8532,N_86,N_270);
and U8533 (N_8533,N_2762,N_1470);
nand U8534 (N_8534,N_1939,N_243);
or U8535 (N_8535,N_2403,N_4911);
and U8536 (N_8536,N_2748,N_2899);
or U8537 (N_8537,N_4980,N_4846);
nand U8538 (N_8538,N_3723,N_4386);
and U8539 (N_8539,N_3074,N_3385);
and U8540 (N_8540,N_2066,N_3137);
or U8541 (N_8541,N_2597,N_2497);
and U8542 (N_8542,N_2591,N_1867);
and U8543 (N_8543,N_2224,N_4436);
or U8544 (N_8544,N_4925,N_1027);
nand U8545 (N_8545,N_2525,N_778);
nand U8546 (N_8546,N_2632,N_1848);
nand U8547 (N_8547,N_2863,N_497);
nand U8548 (N_8548,N_589,N_4640);
or U8549 (N_8549,N_40,N_2594);
nand U8550 (N_8550,N_469,N_2949);
or U8551 (N_8551,N_2226,N_2411);
or U8552 (N_8552,N_2955,N_601);
or U8553 (N_8553,N_1474,N_1116);
and U8554 (N_8554,N_1706,N_1399);
nor U8555 (N_8555,N_3747,N_338);
nand U8556 (N_8556,N_3462,N_4353);
nand U8557 (N_8557,N_1666,N_4228);
and U8558 (N_8558,N_621,N_2884);
nor U8559 (N_8559,N_2644,N_3297);
and U8560 (N_8560,N_287,N_3946);
nor U8561 (N_8561,N_1095,N_3787);
nor U8562 (N_8562,N_3363,N_3834);
and U8563 (N_8563,N_4527,N_3526);
nand U8564 (N_8564,N_4498,N_767);
nor U8565 (N_8565,N_50,N_1150);
and U8566 (N_8566,N_2073,N_2837);
nor U8567 (N_8567,N_4933,N_1754);
and U8568 (N_8568,N_3772,N_2103);
and U8569 (N_8569,N_3287,N_3232);
or U8570 (N_8570,N_1160,N_3821);
nor U8571 (N_8571,N_529,N_3595);
nor U8572 (N_8572,N_3292,N_3144);
and U8573 (N_8573,N_4087,N_3357);
and U8574 (N_8574,N_1680,N_4666);
or U8575 (N_8575,N_4573,N_448);
nor U8576 (N_8576,N_4686,N_3246);
or U8577 (N_8577,N_3666,N_1989);
nor U8578 (N_8578,N_929,N_3304);
or U8579 (N_8579,N_3691,N_3752);
nand U8580 (N_8580,N_499,N_2060);
or U8581 (N_8581,N_1203,N_4011);
or U8582 (N_8582,N_588,N_3073);
and U8583 (N_8583,N_4913,N_1119);
nand U8584 (N_8584,N_1101,N_2433);
or U8585 (N_8585,N_497,N_995);
or U8586 (N_8586,N_899,N_2739);
nand U8587 (N_8587,N_1314,N_3899);
and U8588 (N_8588,N_1736,N_1992);
or U8589 (N_8589,N_4120,N_4757);
and U8590 (N_8590,N_1199,N_1185);
and U8591 (N_8591,N_1339,N_2744);
and U8592 (N_8592,N_1620,N_4322);
or U8593 (N_8593,N_3013,N_1161);
and U8594 (N_8594,N_2511,N_40);
and U8595 (N_8595,N_4756,N_4626);
xnor U8596 (N_8596,N_3140,N_616);
nand U8597 (N_8597,N_207,N_2894);
and U8598 (N_8598,N_3916,N_1281);
nand U8599 (N_8599,N_3931,N_3356);
and U8600 (N_8600,N_4943,N_2168);
or U8601 (N_8601,N_4565,N_4105);
or U8602 (N_8602,N_4119,N_3369);
and U8603 (N_8603,N_340,N_3892);
or U8604 (N_8604,N_4675,N_1884);
xor U8605 (N_8605,N_3351,N_3149);
nand U8606 (N_8606,N_2842,N_3220);
xor U8607 (N_8607,N_1892,N_940);
nor U8608 (N_8608,N_792,N_1639);
or U8609 (N_8609,N_751,N_3185);
nor U8610 (N_8610,N_2547,N_2593);
nand U8611 (N_8611,N_1769,N_4571);
xor U8612 (N_8612,N_4763,N_463);
nor U8613 (N_8613,N_836,N_3778);
nor U8614 (N_8614,N_2823,N_817);
or U8615 (N_8615,N_2571,N_3103);
and U8616 (N_8616,N_972,N_1133);
nand U8617 (N_8617,N_1828,N_447);
and U8618 (N_8618,N_1280,N_1789);
xor U8619 (N_8619,N_1003,N_40);
and U8620 (N_8620,N_3433,N_2445);
nor U8621 (N_8621,N_690,N_744);
nand U8622 (N_8622,N_4501,N_4072);
nor U8623 (N_8623,N_4546,N_701);
nand U8624 (N_8624,N_2106,N_3181);
nand U8625 (N_8625,N_4194,N_996);
nor U8626 (N_8626,N_4845,N_4836);
and U8627 (N_8627,N_2409,N_1863);
nand U8628 (N_8628,N_1414,N_4774);
and U8629 (N_8629,N_4033,N_3770);
or U8630 (N_8630,N_3736,N_1925);
or U8631 (N_8631,N_2497,N_4051);
xnor U8632 (N_8632,N_1278,N_4277);
nor U8633 (N_8633,N_3581,N_4111);
and U8634 (N_8634,N_1764,N_285);
nor U8635 (N_8635,N_4875,N_1352);
and U8636 (N_8636,N_4985,N_4329);
or U8637 (N_8637,N_2772,N_1047);
and U8638 (N_8638,N_3116,N_2121);
nand U8639 (N_8639,N_1055,N_1942);
xnor U8640 (N_8640,N_3572,N_1600);
nor U8641 (N_8641,N_285,N_4678);
xor U8642 (N_8642,N_2681,N_3375);
and U8643 (N_8643,N_857,N_4672);
or U8644 (N_8644,N_3157,N_3421);
and U8645 (N_8645,N_1384,N_1729);
nor U8646 (N_8646,N_2101,N_2580);
and U8647 (N_8647,N_3307,N_3730);
nand U8648 (N_8648,N_2555,N_4575);
or U8649 (N_8649,N_3493,N_1245);
and U8650 (N_8650,N_4462,N_4796);
nand U8651 (N_8651,N_279,N_3188);
nand U8652 (N_8652,N_740,N_1336);
or U8653 (N_8653,N_1333,N_1384);
nand U8654 (N_8654,N_4040,N_2826);
or U8655 (N_8655,N_3675,N_3257);
or U8656 (N_8656,N_84,N_2494);
and U8657 (N_8657,N_1854,N_1166);
or U8658 (N_8658,N_1349,N_1019);
nor U8659 (N_8659,N_513,N_664);
nand U8660 (N_8660,N_3400,N_2384);
nor U8661 (N_8661,N_319,N_2023);
or U8662 (N_8662,N_1634,N_1661);
and U8663 (N_8663,N_504,N_2452);
nand U8664 (N_8664,N_180,N_2764);
and U8665 (N_8665,N_1445,N_3432);
and U8666 (N_8666,N_4905,N_282);
and U8667 (N_8667,N_757,N_1586);
or U8668 (N_8668,N_1539,N_2894);
nand U8669 (N_8669,N_3241,N_2924);
nor U8670 (N_8670,N_494,N_2630);
or U8671 (N_8671,N_4802,N_1751);
or U8672 (N_8672,N_3796,N_1563);
nor U8673 (N_8673,N_2805,N_268);
nor U8674 (N_8674,N_278,N_1180);
xnor U8675 (N_8675,N_1186,N_1293);
or U8676 (N_8676,N_418,N_2737);
or U8677 (N_8677,N_3762,N_1424);
or U8678 (N_8678,N_1913,N_57);
or U8679 (N_8679,N_682,N_425);
or U8680 (N_8680,N_4505,N_1134);
or U8681 (N_8681,N_4069,N_1072);
nor U8682 (N_8682,N_47,N_1295);
nor U8683 (N_8683,N_177,N_3022);
or U8684 (N_8684,N_3850,N_2581);
nand U8685 (N_8685,N_3422,N_2962);
nor U8686 (N_8686,N_2027,N_2130);
nand U8687 (N_8687,N_593,N_4749);
nor U8688 (N_8688,N_2415,N_4893);
nor U8689 (N_8689,N_4224,N_1439);
nor U8690 (N_8690,N_2062,N_1055);
nand U8691 (N_8691,N_2664,N_3958);
nand U8692 (N_8692,N_4533,N_3056);
or U8693 (N_8693,N_4427,N_74);
nor U8694 (N_8694,N_3992,N_2538);
nor U8695 (N_8695,N_3656,N_4497);
and U8696 (N_8696,N_3981,N_4582);
or U8697 (N_8697,N_1,N_2130);
and U8698 (N_8698,N_3972,N_1290);
and U8699 (N_8699,N_3664,N_730);
or U8700 (N_8700,N_3489,N_4341);
and U8701 (N_8701,N_1930,N_3681);
nand U8702 (N_8702,N_4001,N_1375);
or U8703 (N_8703,N_2493,N_4631);
and U8704 (N_8704,N_282,N_4651);
and U8705 (N_8705,N_1172,N_3547);
nor U8706 (N_8706,N_1183,N_2141);
or U8707 (N_8707,N_1685,N_701);
and U8708 (N_8708,N_2206,N_362);
and U8709 (N_8709,N_1238,N_2347);
nand U8710 (N_8710,N_4058,N_2300);
nor U8711 (N_8711,N_4665,N_2391);
nand U8712 (N_8712,N_3723,N_4726);
or U8713 (N_8713,N_2070,N_213);
or U8714 (N_8714,N_3713,N_4938);
nand U8715 (N_8715,N_2912,N_1263);
and U8716 (N_8716,N_2876,N_718);
and U8717 (N_8717,N_3078,N_917);
and U8718 (N_8718,N_1554,N_992);
or U8719 (N_8719,N_617,N_653);
nand U8720 (N_8720,N_377,N_1730);
nand U8721 (N_8721,N_92,N_1103);
xor U8722 (N_8722,N_987,N_1988);
or U8723 (N_8723,N_3321,N_2617);
and U8724 (N_8724,N_4699,N_3684);
nor U8725 (N_8725,N_2015,N_4149);
nand U8726 (N_8726,N_4732,N_3102);
nand U8727 (N_8727,N_1662,N_2964);
nand U8728 (N_8728,N_1091,N_1934);
nor U8729 (N_8729,N_467,N_4378);
or U8730 (N_8730,N_898,N_1935);
nor U8731 (N_8731,N_4426,N_380);
and U8732 (N_8732,N_1177,N_3535);
nand U8733 (N_8733,N_220,N_838);
and U8734 (N_8734,N_4972,N_4331);
nand U8735 (N_8735,N_4896,N_2564);
nor U8736 (N_8736,N_1264,N_475);
nand U8737 (N_8737,N_914,N_2817);
and U8738 (N_8738,N_4487,N_4063);
and U8739 (N_8739,N_241,N_1142);
nor U8740 (N_8740,N_345,N_4032);
nor U8741 (N_8741,N_895,N_1134);
or U8742 (N_8742,N_3069,N_3298);
and U8743 (N_8743,N_1791,N_4356);
or U8744 (N_8744,N_3023,N_4948);
nand U8745 (N_8745,N_4565,N_2064);
nor U8746 (N_8746,N_918,N_3322);
or U8747 (N_8747,N_1497,N_699);
xor U8748 (N_8748,N_1966,N_530);
and U8749 (N_8749,N_3101,N_125);
nand U8750 (N_8750,N_505,N_1138);
nor U8751 (N_8751,N_4855,N_4288);
nand U8752 (N_8752,N_823,N_3325);
nand U8753 (N_8753,N_338,N_144);
or U8754 (N_8754,N_2843,N_2416);
nand U8755 (N_8755,N_1595,N_1808);
and U8756 (N_8756,N_2571,N_4708);
nand U8757 (N_8757,N_1445,N_792);
nor U8758 (N_8758,N_3096,N_1641);
or U8759 (N_8759,N_1,N_507);
nor U8760 (N_8760,N_2496,N_3730);
nor U8761 (N_8761,N_3190,N_963);
or U8762 (N_8762,N_3598,N_2846);
nand U8763 (N_8763,N_4669,N_3706);
nand U8764 (N_8764,N_4890,N_362);
xnor U8765 (N_8765,N_3808,N_4826);
nand U8766 (N_8766,N_973,N_2486);
nor U8767 (N_8767,N_654,N_2826);
nand U8768 (N_8768,N_3369,N_4137);
nor U8769 (N_8769,N_4700,N_3305);
nand U8770 (N_8770,N_3575,N_3695);
and U8771 (N_8771,N_4062,N_3676);
or U8772 (N_8772,N_4346,N_4596);
and U8773 (N_8773,N_753,N_299);
or U8774 (N_8774,N_4693,N_3158);
and U8775 (N_8775,N_3385,N_3455);
nand U8776 (N_8776,N_4397,N_2356);
and U8777 (N_8777,N_1717,N_4756);
and U8778 (N_8778,N_2460,N_2330);
xor U8779 (N_8779,N_1034,N_1765);
and U8780 (N_8780,N_3253,N_66);
or U8781 (N_8781,N_4008,N_4571);
and U8782 (N_8782,N_4565,N_3005);
and U8783 (N_8783,N_4744,N_841);
xor U8784 (N_8784,N_3456,N_2879);
or U8785 (N_8785,N_4691,N_4004);
nor U8786 (N_8786,N_2967,N_3231);
nor U8787 (N_8787,N_3882,N_1058);
or U8788 (N_8788,N_2220,N_1386);
nand U8789 (N_8789,N_4449,N_2059);
or U8790 (N_8790,N_4907,N_753);
nor U8791 (N_8791,N_819,N_3387);
and U8792 (N_8792,N_739,N_3513);
and U8793 (N_8793,N_2897,N_3659);
nand U8794 (N_8794,N_1740,N_4697);
nand U8795 (N_8795,N_1055,N_4025);
and U8796 (N_8796,N_4041,N_3188);
nor U8797 (N_8797,N_4508,N_819);
or U8798 (N_8798,N_737,N_1190);
and U8799 (N_8799,N_4291,N_4351);
and U8800 (N_8800,N_3962,N_4586);
and U8801 (N_8801,N_2637,N_2339);
nand U8802 (N_8802,N_3521,N_1093);
nand U8803 (N_8803,N_2371,N_797);
or U8804 (N_8804,N_664,N_3588);
nor U8805 (N_8805,N_2427,N_4419);
nand U8806 (N_8806,N_2290,N_3128);
nand U8807 (N_8807,N_1542,N_346);
and U8808 (N_8808,N_4235,N_3014);
and U8809 (N_8809,N_732,N_3295);
nor U8810 (N_8810,N_3372,N_2395);
or U8811 (N_8811,N_1309,N_1067);
or U8812 (N_8812,N_4716,N_1476);
nand U8813 (N_8813,N_1425,N_1568);
xor U8814 (N_8814,N_4095,N_832);
and U8815 (N_8815,N_2835,N_3925);
nor U8816 (N_8816,N_1629,N_4947);
or U8817 (N_8817,N_1185,N_4445);
or U8818 (N_8818,N_2832,N_2614);
nand U8819 (N_8819,N_994,N_312);
and U8820 (N_8820,N_4184,N_2513);
and U8821 (N_8821,N_878,N_2903);
nor U8822 (N_8822,N_695,N_4649);
or U8823 (N_8823,N_99,N_856);
or U8824 (N_8824,N_2815,N_3692);
nor U8825 (N_8825,N_1857,N_399);
nor U8826 (N_8826,N_1058,N_215);
and U8827 (N_8827,N_4188,N_1471);
nor U8828 (N_8828,N_3775,N_321);
nor U8829 (N_8829,N_1593,N_1312);
and U8830 (N_8830,N_147,N_4274);
nand U8831 (N_8831,N_3229,N_741);
nor U8832 (N_8832,N_668,N_1150);
or U8833 (N_8833,N_3649,N_4438);
nor U8834 (N_8834,N_3405,N_1584);
or U8835 (N_8835,N_1255,N_3431);
and U8836 (N_8836,N_2167,N_3643);
or U8837 (N_8837,N_4891,N_337);
nor U8838 (N_8838,N_157,N_2711);
nand U8839 (N_8839,N_2904,N_61);
and U8840 (N_8840,N_2108,N_338);
nand U8841 (N_8841,N_1249,N_2253);
nand U8842 (N_8842,N_1490,N_3402);
nor U8843 (N_8843,N_1154,N_1721);
or U8844 (N_8844,N_4245,N_4024);
or U8845 (N_8845,N_3834,N_3204);
nor U8846 (N_8846,N_4352,N_7);
nand U8847 (N_8847,N_3341,N_3320);
and U8848 (N_8848,N_359,N_2971);
nor U8849 (N_8849,N_1760,N_1223);
nand U8850 (N_8850,N_1053,N_2565);
nand U8851 (N_8851,N_1376,N_3741);
or U8852 (N_8852,N_1032,N_1618);
nand U8853 (N_8853,N_4933,N_3982);
nand U8854 (N_8854,N_3416,N_1747);
or U8855 (N_8855,N_2664,N_2929);
nand U8856 (N_8856,N_2944,N_4146);
and U8857 (N_8857,N_516,N_3553);
nand U8858 (N_8858,N_3647,N_1021);
or U8859 (N_8859,N_4645,N_23);
nor U8860 (N_8860,N_4566,N_3776);
nand U8861 (N_8861,N_2493,N_1519);
or U8862 (N_8862,N_3442,N_4899);
nor U8863 (N_8863,N_392,N_1184);
or U8864 (N_8864,N_965,N_3291);
nand U8865 (N_8865,N_4287,N_4557);
nor U8866 (N_8866,N_1978,N_143);
nor U8867 (N_8867,N_132,N_1240);
nand U8868 (N_8868,N_4825,N_917);
or U8869 (N_8869,N_3691,N_1321);
and U8870 (N_8870,N_2215,N_2493);
and U8871 (N_8871,N_3055,N_2911);
nor U8872 (N_8872,N_934,N_2746);
and U8873 (N_8873,N_666,N_241);
nor U8874 (N_8874,N_4655,N_4076);
nor U8875 (N_8875,N_337,N_1466);
nor U8876 (N_8876,N_4511,N_4210);
or U8877 (N_8877,N_2558,N_2022);
or U8878 (N_8878,N_4143,N_3265);
nor U8879 (N_8879,N_4220,N_1754);
and U8880 (N_8880,N_2708,N_3630);
nor U8881 (N_8881,N_4854,N_2215);
and U8882 (N_8882,N_726,N_936);
and U8883 (N_8883,N_639,N_3059);
and U8884 (N_8884,N_852,N_1110);
nor U8885 (N_8885,N_1254,N_1906);
or U8886 (N_8886,N_548,N_3128);
nand U8887 (N_8887,N_2409,N_145);
nand U8888 (N_8888,N_1788,N_208);
and U8889 (N_8889,N_4393,N_2403);
nand U8890 (N_8890,N_716,N_479);
and U8891 (N_8891,N_145,N_584);
nor U8892 (N_8892,N_863,N_4883);
nor U8893 (N_8893,N_4316,N_3355);
and U8894 (N_8894,N_4428,N_2384);
nor U8895 (N_8895,N_3460,N_3413);
and U8896 (N_8896,N_4691,N_972);
or U8897 (N_8897,N_4662,N_1757);
or U8898 (N_8898,N_4854,N_1743);
nand U8899 (N_8899,N_4376,N_4226);
nor U8900 (N_8900,N_899,N_3628);
nand U8901 (N_8901,N_3908,N_1243);
and U8902 (N_8902,N_2191,N_2534);
or U8903 (N_8903,N_743,N_1942);
nand U8904 (N_8904,N_199,N_654);
and U8905 (N_8905,N_4913,N_986);
or U8906 (N_8906,N_1542,N_350);
nand U8907 (N_8907,N_1896,N_978);
and U8908 (N_8908,N_4239,N_451);
nand U8909 (N_8909,N_3290,N_1988);
nand U8910 (N_8910,N_2872,N_3179);
nor U8911 (N_8911,N_4454,N_2433);
nor U8912 (N_8912,N_2673,N_391);
and U8913 (N_8913,N_92,N_4015);
or U8914 (N_8914,N_3983,N_4331);
nand U8915 (N_8915,N_3316,N_1713);
or U8916 (N_8916,N_4774,N_2904);
nor U8917 (N_8917,N_4934,N_467);
or U8918 (N_8918,N_4342,N_1777);
nor U8919 (N_8919,N_4305,N_2754);
xor U8920 (N_8920,N_159,N_2254);
nor U8921 (N_8921,N_4903,N_4952);
or U8922 (N_8922,N_1555,N_4742);
nor U8923 (N_8923,N_1878,N_3724);
nand U8924 (N_8924,N_3170,N_788);
or U8925 (N_8925,N_2493,N_3291);
nor U8926 (N_8926,N_3283,N_4386);
or U8927 (N_8927,N_3087,N_97);
nor U8928 (N_8928,N_3511,N_2882);
or U8929 (N_8929,N_133,N_3740);
xor U8930 (N_8930,N_1123,N_1764);
and U8931 (N_8931,N_3062,N_3444);
nor U8932 (N_8932,N_4323,N_4298);
xnor U8933 (N_8933,N_2588,N_464);
or U8934 (N_8934,N_4792,N_2078);
or U8935 (N_8935,N_3881,N_107);
or U8936 (N_8936,N_2188,N_4666);
nand U8937 (N_8937,N_1460,N_4980);
nand U8938 (N_8938,N_3627,N_602);
or U8939 (N_8939,N_3516,N_3519);
nor U8940 (N_8940,N_2701,N_3780);
or U8941 (N_8941,N_1540,N_4555);
nor U8942 (N_8942,N_2107,N_4944);
nand U8943 (N_8943,N_1213,N_3681);
nand U8944 (N_8944,N_4690,N_596);
and U8945 (N_8945,N_4995,N_2812);
nor U8946 (N_8946,N_2720,N_3278);
or U8947 (N_8947,N_3691,N_4933);
and U8948 (N_8948,N_1557,N_3397);
nand U8949 (N_8949,N_3129,N_4558);
and U8950 (N_8950,N_3917,N_1188);
xor U8951 (N_8951,N_3041,N_936);
and U8952 (N_8952,N_1710,N_676);
and U8953 (N_8953,N_1571,N_3149);
nor U8954 (N_8954,N_1055,N_2158);
nand U8955 (N_8955,N_3224,N_1279);
and U8956 (N_8956,N_37,N_3643);
or U8957 (N_8957,N_4260,N_893);
or U8958 (N_8958,N_2162,N_4964);
or U8959 (N_8959,N_4690,N_3338);
nand U8960 (N_8960,N_1416,N_3129);
nand U8961 (N_8961,N_480,N_4945);
nor U8962 (N_8962,N_4285,N_3178);
nor U8963 (N_8963,N_2194,N_2016);
and U8964 (N_8964,N_976,N_2728);
nor U8965 (N_8965,N_1004,N_2615);
nand U8966 (N_8966,N_4644,N_769);
nand U8967 (N_8967,N_3749,N_2436);
or U8968 (N_8968,N_4159,N_3930);
or U8969 (N_8969,N_817,N_3385);
or U8970 (N_8970,N_3231,N_4463);
and U8971 (N_8971,N_1180,N_2196);
and U8972 (N_8972,N_1453,N_890);
xor U8973 (N_8973,N_3435,N_4867);
or U8974 (N_8974,N_3085,N_2653);
or U8975 (N_8975,N_1303,N_1763);
nor U8976 (N_8976,N_4060,N_2055);
nand U8977 (N_8977,N_1804,N_540);
nor U8978 (N_8978,N_3039,N_4941);
nand U8979 (N_8979,N_3458,N_2409);
nand U8980 (N_8980,N_3332,N_3540);
nor U8981 (N_8981,N_4814,N_3958);
nor U8982 (N_8982,N_1789,N_551);
nor U8983 (N_8983,N_3760,N_311);
and U8984 (N_8984,N_2673,N_565);
nor U8985 (N_8985,N_434,N_1858);
and U8986 (N_8986,N_4526,N_3667);
nor U8987 (N_8987,N_1453,N_1480);
nor U8988 (N_8988,N_739,N_3866);
nor U8989 (N_8989,N_1651,N_2985);
and U8990 (N_8990,N_460,N_1646);
nor U8991 (N_8991,N_1130,N_4313);
nor U8992 (N_8992,N_3820,N_4337);
and U8993 (N_8993,N_2292,N_734);
nand U8994 (N_8994,N_1070,N_4663);
nor U8995 (N_8995,N_4605,N_2586);
nor U8996 (N_8996,N_326,N_45);
or U8997 (N_8997,N_4613,N_48);
or U8998 (N_8998,N_4321,N_2595);
nand U8999 (N_8999,N_3517,N_4964);
nand U9000 (N_9000,N_3787,N_120);
or U9001 (N_9001,N_152,N_1251);
and U9002 (N_9002,N_4376,N_3692);
xor U9003 (N_9003,N_4654,N_2742);
and U9004 (N_9004,N_1446,N_3195);
nor U9005 (N_9005,N_2464,N_406);
xnor U9006 (N_9006,N_4524,N_2537);
and U9007 (N_9007,N_4333,N_816);
nor U9008 (N_9008,N_3583,N_4331);
nor U9009 (N_9009,N_2528,N_1299);
or U9010 (N_9010,N_3512,N_1984);
nand U9011 (N_9011,N_4976,N_1283);
xnor U9012 (N_9012,N_3378,N_2871);
and U9013 (N_9013,N_126,N_2412);
or U9014 (N_9014,N_2389,N_1214);
and U9015 (N_9015,N_3784,N_4560);
or U9016 (N_9016,N_3549,N_3419);
or U9017 (N_9017,N_2175,N_684);
nand U9018 (N_9018,N_2762,N_794);
nor U9019 (N_9019,N_2932,N_1574);
and U9020 (N_9020,N_3970,N_2662);
or U9021 (N_9021,N_4254,N_3215);
nand U9022 (N_9022,N_1012,N_4604);
or U9023 (N_9023,N_787,N_650);
and U9024 (N_9024,N_1236,N_4272);
nor U9025 (N_9025,N_3466,N_1889);
or U9026 (N_9026,N_1435,N_1874);
nor U9027 (N_9027,N_1828,N_3613);
or U9028 (N_9028,N_2309,N_2833);
or U9029 (N_9029,N_2089,N_2406);
or U9030 (N_9030,N_4545,N_763);
and U9031 (N_9031,N_1561,N_2517);
nor U9032 (N_9032,N_4098,N_4437);
and U9033 (N_9033,N_2716,N_2183);
and U9034 (N_9034,N_1946,N_3574);
or U9035 (N_9035,N_37,N_2554);
nor U9036 (N_9036,N_247,N_1516);
or U9037 (N_9037,N_2847,N_831);
nor U9038 (N_9038,N_1567,N_4902);
or U9039 (N_9039,N_925,N_3593);
or U9040 (N_9040,N_3317,N_405);
nand U9041 (N_9041,N_3799,N_4403);
or U9042 (N_9042,N_1289,N_88);
and U9043 (N_9043,N_980,N_3971);
nand U9044 (N_9044,N_4459,N_4948);
or U9045 (N_9045,N_3925,N_2006);
nand U9046 (N_9046,N_4151,N_1042);
and U9047 (N_9047,N_4759,N_4981);
nor U9048 (N_9048,N_2633,N_1907);
nand U9049 (N_9049,N_1605,N_2366);
nand U9050 (N_9050,N_1318,N_4201);
and U9051 (N_9051,N_4592,N_1646);
nand U9052 (N_9052,N_4318,N_4660);
or U9053 (N_9053,N_4431,N_3657);
xnor U9054 (N_9054,N_1455,N_2962);
nand U9055 (N_9055,N_1829,N_1676);
xnor U9056 (N_9056,N_3419,N_3450);
nor U9057 (N_9057,N_2302,N_6);
nand U9058 (N_9058,N_3120,N_1349);
nor U9059 (N_9059,N_4270,N_2010);
or U9060 (N_9060,N_3387,N_3171);
nand U9061 (N_9061,N_4085,N_1622);
and U9062 (N_9062,N_414,N_394);
nor U9063 (N_9063,N_4208,N_2481);
nor U9064 (N_9064,N_3643,N_3899);
nand U9065 (N_9065,N_2673,N_4973);
or U9066 (N_9066,N_1488,N_1463);
nor U9067 (N_9067,N_293,N_1095);
nor U9068 (N_9068,N_236,N_1550);
nor U9069 (N_9069,N_4760,N_4670);
and U9070 (N_9070,N_2046,N_3175);
nor U9071 (N_9071,N_934,N_930);
nor U9072 (N_9072,N_276,N_4566);
and U9073 (N_9073,N_1432,N_4101);
nor U9074 (N_9074,N_111,N_773);
or U9075 (N_9075,N_2613,N_124);
nand U9076 (N_9076,N_3757,N_4935);
nor U9077 (N_9077,N_3227,N_917);
nand U9078 (N_9078,N_4359,N_2005);
nand U9079 (N_9079,N_4062,N_2844);
and U9080 (N_9080,N_2876,N_2863);
nor U9081 (N_9081,N_1752,N_1253);
or U9082 (N_9082,N_2450,N_643);
or U9083 (N_9083,N_4624,N_3134);
nor U9084 (N_9084,N_4226,N_699);
nor U9085 (N_9085,N_911,N_3097);
or U9086 (N_9086,N_1238,N_1980);
and U9087 (N_9087,N_269,N_4263);
and U9088 (N_9088,N_354,N_2938);
xnor U9089 (N_9089,N_1309,N_4349);
or U9090 (N_9090,N_722,N_3791);
or U9091 (N_9091,N_4381,N_1115);
nor U9092 (N_9092,N_3851,N_4392);
or U9093 (N_9093,N_4357,N_3949);
and U9094 (N_9094,N_1832,N_3356);
and U9095 (N_9095,N_3114,N_3866);
nand U9096 (N_9096,N_1101,N_3000);
nor U9097 (N_9097,N_1126,N_4251);
nand U9098 (N_9098,N_1341,N_332);
nor U9099 (N_9099,N_4293,N_67);
and U9100 (N_9100,N_4367,N_1556);
or U9101 (N_9101,N_509,N_1384);
or U9102 (N_9102,N_4104,N_2233);
nand U9103 (N_9103,N_4755,N_4805);
or U9104 (N_9104,N_3992,N_3933);
or U9105 (N_9105,N_276,N_196);
or U9106 (N_9106,N_4425,N_922);
and U9107 (N_9107,N_1878,N_1508);
nor U9108 (N_9108,N_4116,N_4214);
nor U9109 (N_9109,N_4251,N_1334);
and U9110 (N_9110,N_339,N_4512);
nand U9111 (N_9111,N_141,N_3511);
and U9112 (N_9112,N_3003,N_3996);
or U9113 (N_9113,N_2169,N_2962);
nor U9114 (N_9114,N_3987,N_4949);
or U9115 (N_9115,N_2681,N_4616);
nor U9116 (N_9116,N_2956,N_1997);
nor U9117 (N_9117,N_3869,N_3440);
or U9118 (N_9118,N_3530,N_901);
xor U9119 (N_9119,N_4348,N_730);
nand U9120 (N_9120,N_4903,N_2683);
or U9121 (N_9121,N_3880,N_3028);
or U9122 (N_9122,N_1390,N_232);
nor U9123 (N_9123,N_2710,N_4542);
or U9124 (N_9124,N_3364,N_193);
and U9125 (N_9125,N_4961,N_2447);
nor U9126 (N_9126,N_1330,N_4011);
nor U9127 (N_9127,N_3263,N_1820);
nor U9128 (N_9128,N_226,N_552);
xor U9129 (N_9129,N_1954,N_4093);
nand U9130 (N_9130,N_3335,N_293);
or U9131 (N_9131,N_582,N_4851);
nor U9132 (N_9132,N_4250,N_456);
and U9133 (N_9133,N_1913,N_1070);
and U9134 (N_9134,N_1993,N_412);
nor U9135 (N_9135,N_3165,N_4376);
or U9136 (N_9136,N_2898,N_2384);
nor U9137 (N_9137,N_2992,N_1138);
nor U9138 (N_9138,N_988,N_4784);
and U9139 (N_9139,N_190,N_3191);
nor U9140 (N_9140,N_1001,N_2558);
and U9141 (N_9141,N_2975,N_270);
or U9142 (N_9142,N_3592,N_181);
nand U9143 (N_9143,N_1279,N_4663);
xnor U9144 (N_9144,N_473,N_4896);
or U9145 (N_9145,N_1517,N_1793);
nand U9146 (N_9146,N_1063,N_4397);
xor U9147 (N_9147,N_4233,N_4355);
nor U9148 (N_9148,N_2267,N_2809);
nand U9149 (N_9149,N_4340,N_4610);
nor U9150 (N_9150,N_843,N_4190);
or U9151 (N_9151,N_1424,N_1111);
and U9152 (N_9152,N_2427,N_2583);
and U9153 (N_9153,N_1867,N_3739);
or U9154 (N_9154,N_1027,N_1739);
nand U9155 (N_9155,N_3594,N_640);
and U9156 (N_9156,N_2634,N_1932);
nand U9157 (N_9157,N_1526,N_407);
or U9158 (N_9158,N_8,N_1290);
nand U9159 (N_9159,N_2101,N_4279);
or U9160 (N_9160,N_4745,N_1491);
nand U9161 (N_9161,N_2142,N_149);
nand U9162 (N_9162,N_4157,N_1482);
or U9163 (N_9163,N_4659,N_4760);
or U9164 (N_9164,N_2762,N_4869);
nor U9165 (N_9165,N_1074,N_4503);
or U9166 (N_9166,N_871,N_4382);
and U9167 (N_9167,N_3045,N_2105);
or U9168 (N_9168,N_1114,N_1797);
or U9169 (N_9169,N_2901,N_1066);
and U9170 (N_9170,N_1373,N_2346);
nand U9171 (N_9171,N_2626,N_2018);
and U9172 (N_9172,N_2851,N_924);
or U9173 (N_9173,N_2600,N_1062);
nor U9174 (N_9174,N_2776,N_474);
nor U9175 (N_9175,N_2350,N_3875);
nand U9176 (N_9176,N_3862,N_695);
and U9177 (N_9177,N_3972,N_2222);
or U9178 (N_9178,N_396,N_536);
nor U9179 (N_9179,N_4814,N_1983);
nand U9180 (N_9180,N_2534,N_3295);
and U9181 (N_9181,N_3036,N_2861);
nand U9182 (N_9182,N_880,N_1785);
and U9183 (N_9183,N_1687,N_4671);
nor U9184 (N_9184,N_4591,N_4365);
nor U9185 (N_9185,N_865,N_1600);
or U9186 (N_9186,N_291,N_100);
or U9187 (N_9187,N_2923,N_4640);
or U9188 (N_9188,N_1743,N_3952);
or U9189 (N_9189,N_3928,N_3390);
nor U9190 (N_9190,N_1193,N_3375);
or U9191 (N_9191,N_3782,N_1234);
or U9192 (N_9192,N_2003,N_4742);
or U9193 (N_9193,N_3101,N_1000);
and U9194 (N_9194,N_4463,N_4229);
nor U9195 (N_9195,N_876,N_4644);
nor U9196 (N_9196,N_4055,N_2998);
and U9197 (N_9197,N_4042,N_4021);
or U9198 (N_9198,N_51,N_1561);
nor U9199 (N_9199,N_206,N_2950);
nand U9200 (N_9200,N_937,N_4635);
or U9201 (N_9201,N_2711,N_4760);
nor U9202 (N_9202,N_2681,N_4520);
xor U9203 (N_9203,N_3584,N_2407);
or U9204 (N_9204,N_4563,N_433);
or U9205 (N_9205,N_3575,N_1924);
nor U9206 (N_9206,N_1623,N_2088);
or U9207 (N_9207,N_3776,N_266);
and U9208 (N_9208,N_1903,N_2415);
nand U9209 (N_9209,N_2324,N_2465);
nand U9210 (N_9210,N_1455,N_1548);
or U9211 (N_9211,N_206,N_3625);
xnor U9212 (N_9212,N_1851,N_4911);
and U9213 (N_9213,N_2883,N_4274);
or U9214 (N_9214,N_655,N_2963);
or U9215 (N_9215,N_4248,N_2347);
and U9216 (N_9216,N_3586,N_3504);
nor U9217 (N_9217,N_639,N_75);
nand U9218 (N_9218,N_1475,N_2792);
and U9219 (N_9219,N_814,N_3618);
nor U9220 (N_9220,N_3674,N_4369);
nor U9221 (N_9221,N_4240,N_809);
or U9222 (N_9222,N_2236,N_859);
nand U9223 (N_9223,N_4638,N_1580);
and U9224 (N_9224,N_413,N_2272);
or U9225 (N_9225,N_768,N_2614);
nand U9226 (N_9226,N_2039,N_2743);
and U9227 (N_9227,N_3559,N_2130);
and U9228 (N_9228,N_2470,N_3407);
and U9229 (N_9229,N_4853,N_942);
or U9230 (N_9230,N_1525,N_1327);
nor U9231 (N_9231,N_2502,N_4313);
nand U9232 (N_9232,N_2327,N_1127);
nor U9233 (N_9233,N_4150,N_1975);
and U9234 (N_9234,N_2847,N_1179);
or U9235 (N_9235,N_1302,N_837);
nor U9236 (N_9236,N_2179,N_23);
or U9237 (N_9237,N_1858,N_1712);
and U9238 (N_9238,N_2045,N_939);
nor U9239 (N_9239,N_4092,N_2104);
nor U9240 (N_9240,N_678,N_368);
and U9241 (N_9241,N_11,N_4263);
or U9242 (N_9242,N_2536,N_2456);
nand U9243 (N_9243,N_2519,N_3227);
and U9244 (N_9244,N_1140,N_180);
nand U9245 (N_9245,N_761,N_3599);
nand U9246 (N_9246,N_1481,N_308);
or U9247 (N_9247,N_594,N_2989);
and U9248 (N_9248,N_1286,N_77);
or U9249 (N_9249,N_4724,N_2277);
nand U9250 (N_9250,N_4281,N_4703);
nor U9251 (N_9251,N_154,N_2721);
and U9252 (N_9252,N_1710,N_2119);
or U9253 (N_9253,N_2739,N_3200);
and U9254 (N_9254,N_1370,N_446);
and U9255 (N_9255,N_4810,N_1985);
nand U9256 (N_9256,N_4224,N_2079);
nor U9257 (N_9257,N_4445,N_408);
nor U9258 (N_9258,N_1552,N_3102);
xor U9259 (N_9259,N_4651,N_4578);
or U9260 (N_9260,N_361,N_4245);
and U9261 (N_9261,N_3794,N_3207);
nor U9262 (N_9262,N_2466,N_829);
nor U9263 (N_9263,N_456,N_4452);
nand U9264 (N_9264,N_81,N_4433);
nor U9265 (N_9265,N_4524,N_4547);
nor U9266 (N_9266,N_2592,N_603);
or U9267 (N_9267,N_3184,N_2180);
and U9268 (N_9268,N_950,N_1364);
and U9269 (N_9269,N_3536,N_301);
nor U9270 (N_9270,N_2342,N_1857);
nand U9271 (N_9271,N_674,N_4212);
and U9272 (N_9272,N_1384,N_1474);
nor U9273 (N_9273,N_2196,N_4302);
nand U9274 (N_9274,N_778,N_1256);
or U9275 (N_9275,N_4285,N_920);
nor U9276 (N_9276,N_913,N_3911);
and U9277 (N_9277,N_1201,N_4739);
nor U9278 (N_9278,N_3825,N_1174);
nand U9279 (N_9279,N_3169,N_512);
and U9280 (N_9280,N_4451,N_1422);
nand U9281 (N_9281,N_2591,N_27);
or U9282 (N_9282,N_2007,N_431);
nand U9283 (N_9283,N_4893,N_4098);
or U9284 (N_9284,N_1440,N_1733);
and U9285 (N_9285,N_2722,N_4793);
nor U9286 (N_9286,N_1670,N_2830);
or U9287 (N_9287,N_1653,N_2601);
and U9288 (N_9288,N_2609,N_2246);
nor U9289 (N_9289,N_3894,N_3120);
nor U9290 (N_9290,N_3879,N_4376);
and U9291 (N_9291,N_1162,N_77);
nand U9292 (N_9292,N_2575,N_4835);
nand U9293 (N_9293,N_1251,N_984);
nand U9294 (N_9294,N_2081,N_4544);
nand U9295 (N_9295,N_2356,N_4527);
and U9296 (N_9296,N_2051,N_4638);
nor U9297 (N_9297,N_1404,N_1294);
or U9298 (N_9298,N_2167,N_1804);
or U9299 (N_9299,N_3470,N_1847);
and U9300 (N_9300,N_240,N_1112);
nand U9301 (N_9301,N_4589,N_766);
or U9302 (N_9302,N_3452,N_2933);
nand U9303 (N_9303,N_4102,N_1849);
nand U9304 (N_9304,N_4730,N_4903);
nand U9305 (N_9305,N_4698,N_2044);
or U9306 (N_9306,N_1424,N_3652);
nand U9307 (N_9307,N_1491,N_3860);
and U9308 (N_9308,N_2840,N_987);
nand U9309 (N_9309,N_4937,N_1322);
nor U9310 (N_9310,N_3857,N_3757);
nor U9311 (N_9311,N_2003,N_1972);
nand U9312 (N_9312,N_1375,N_2620);
nor U9313 (N_9313,N_2333,N_1455);
nand U9314 (N_9314,N_663,N_1416);
and U9315 (N_9315,N_1857,N_2117);
and U9316 (N_9316,N_4586,N_2661);
nand U9317 (N_9317,N_782,N_1294);
or U9318 (N_9318,N_220,N_803);
nor U9319 (N_9319,N_3328,N_3954);
nand U9320 (N_9320,N_3748,N_3263);
nor U9321 (N_9321,N_4831,N_2203);
nor U9322 (N_9322,N_4228,N_1608);
or U9323 (N_9323,N_617,N_4743);
nor U9324 (N_9324,N_3614,N_4599);
nand U9325 (N_9325,N_758,N_66);
nand U9326 (N_9326,N_1623,N_2165);
nor U9327 (N_9327,N_2476,N_1300);
or U9328 (N_9328,N_4614,N_3682);
xor U9329 (N_9329,N_2383,N_4748);
or U9330 (N_9330,N_2533,N_1896);
nand U9331 (N_9331,N_1426,N_3699);
and U9332 (N_9332,N_4692,N_27);
xor U9333 (N_9333,N_3006,N_2518);
and U9334 (N_9334,N_865,N_2095);
nand U9335 (N_9335,N_645,N_3574);
or U9336 (N_9336,N_840,N_2801);
or U9337 (N_9337,N_1608,N_3752);
and U9338 (N_9338,N_2299,N_1480);
or U9339 (N_9339,N_3462,N_1030);
nand U9340 (N_9340,N_1169,N_2217);
nand U9341 (N_9341,N_522,N_851);
or U9342 (N_9342,N_530,N_4313);
xor U9343 (N_9343,N_2311,N_980);
and U9344 (N_9344,N_3632,N_2783);
or U9345 (N_9345,N_2158,N_2327);
nor U9346 (N_9346,N_987,N_4289);
nor U9347 (N_9347,N_4478,N_1352);
and U9348 (N_9348,N_4983,N_4962);
or U9349 (N_9349,N_2299,N_3971);
nor U9350 (N_9350,N_4991,N_1687);
and U9351 (N_9351,N_4285,N_547);
nand U9352 (N_9352,N_31,N_3862);
or U9353 (N_9353,N_1305,N_4351);
nor U9354 (N_9354,N_850,N_2145);
nor U9355 (N_9355,N_2759,N_2982);
or U9356 (N_9356,N_2065,N_1374);
and U9357 (N_9357,N_602,N_4721);
or U9358 (N_9358,N_2717,N_2116);
nor U9359 (N_9359,N_4395,N_1053);
and U9360 (N_9360,N_377,N_2113);
nor U9361 (N_9361,N_1530,N_3381);
and U9362 (N_9362,N_4418,N_2478);
xor U9363 (N_9363,N_4297,N_2760);
or U9364 (N_9364,N_950,N_1509);
and U9365 (N_9365,N_1649,N_4634);
nand U9366 (N_9366,N_4013,N_2105);
and U9367 (N_9367,N_4401,N_2383);
and U9368 (N_9368,N_1550,N_4635);
and U9369 (N_9369,N_2043,N_3893);
or U9370 (N_9370,N_4640,N_3808);
nand U9371 (N_9371,N_205,N_2005);
nor U9372 (N_9372,N_949,N_4217);
and U9373 (N_9373,N_4956,N_1726);
and U9374 (N_9374,N_2276,N_2123);
nor U9375 (N_9375,N_3305,N_2184);
and U9376 (N_9376,N_3910,N_1788);
nor U9377 (N_9377,N_4744,N_833);
or U9378 (N_9378,N_3968,N_485);
nand U9379 (N_9379,N_3891,N_2877);
or U9380 (N_9380,N_4413,N_3270);
or U9381 (N_9381,N_3803,N_1228);
and U9382 (N_9382,N_776,N_3034);
and U9383 (N_9383,N_4514,N_4063);
nor U9384 (N_9384,N_3372,N_4572);
or U9385 (N_9385,N_4418,N_1291);
xor U9386 (N_9386,N_4689,N_2223);
and U9387 (N_9387,N_3680,N_736);
and U9388 (N_9388,N_0,N_2241);
xnor U9389 (N_9389,N_4720,N_3891);
nor U9390 (N_9390,N_3235,N_1673);
xor U9391 (N_9391,N_2386,N_1249);
nor U9392 (N_9392,N_370,N_843);
nor U9393 (N_9393,N_3544,N_4644);
xnor U9394 (N_9394,N_832,N_2808);
and U9395 (N_9395,N_828,N_130);
or U9396 (N_9396,N_185,N_4753);
and U9397 (N_9397,N_840,N_2254);
or U9398 (N_9398,N_3074,N_2303);
nand U9399 (N_9399,N_1563,N_4267);
xnor U9400 (N_9400,N_3746,N_3043);
xor U9401 (N_9401,N_1581,N_2873);
and U9402 (N_9402,N_4812,N_3776);
nor U9403 (N_9403,N_2719,N_4911);
and U9404 (N_9404,N_4087,N_42);
nand U9405 (N_9405,N_1853,N_4229);
or U9406 (N_9406,N_4732,N_4469);
and U9407 (N_9407,N_2202,N_1615);
and U9408 (N_9408,N_4720,N_3552);
and U9409 (N_9409,N_1279,N_249);
nand U9410 (N_9410,N_2192,N_2573);
nand U9411 (N_9411,N_3201,N_4596);
nand U9412 (N_9412,N_4565,N_423);
and U9413 (N_9413,N_462,N_2764);
or U9414 (N_9414,N_1430,N_1607);
or U9415 (N_9415,N_563,N_38);
or U9416 (N_9416,N_1028,N_1833);
and U9417 (N_9417,N_2898,N_688);
nor U9418 (N_9418,N_3300,N_3496);
nand U9419 (N_9419,N_641,N_1299);
or U9420 (N_9420,N_3412,N_2855);
or U9421 (N_9421,N_1982,N_4287);
nor U9422 (N_9422,N_979,N_1019);
nand U9423 (N_9423,N_3080,N_3349);
or U9424 (N_9424,N_4661,N_4909);
nor U9425 (N_9425,N_4621,N_2472);
and U9426 (N_9426,N_210,N_4019);
nand U9427 (N_9427,N_1072,N_3672);
and U9428 (N_9428,N_849,N_3839);
or U9429 (N_9429,N_3169,N_1045);
nor U9430 (N_9430,N_2394,N_3341);
nand U9431 (N_9431,N_4048,N_4002);
nor U9432 (N_9432,N_3219,N_2778);
and U9433 (N_9433,N_2520,N_153);
nand U9434 (N_9434,N_2170,N_4742);
or U9435 (N_9435,N_2742,N_1125);
and U9436 (N_9436,N_118,N_4794);
or U9437 (N_9437,N_689,N_1405);
nand U9438 (N_9438,N_3978,N_4622);
and U9439 (N_9439,N_721,N_4607);
nor U9440 (N_9440,N_1501,N_4382);
or U9441 (N_9441,N_1860,N_697);
nand U9442 (N_9442,N_1234,N_4975);
or U9443 (N_9443,N_3625,N_780);
or U9444 (N_9444,N_3276,N_2302);
or U9445 (N_9445,N_2885,N_4575);
and U9446 (N_9446,N_1498,N_394);
or U9447 (N_9447,N_4188,N_1);
or U9448 (N_9448,N_509,N_333);
and U9449 (N_9449,N_3246,N_3121);
and U9450 (N_9450,N_760,N_946);
or U9451 (N_9451,N_3227,N_2249);
or U9452 (N_9452,N_4612,N_68);
nor U9453 (N_9453,N_3036,N_367);
nand U9454 (N_9454,N_473,N_4779);
or U9455 (N_9455,N_3636,N_2104);
nand U9456 (N_9456,N_1031,N_1276);
and U9457 (N_9457,N_4293,N_2336);
nand U9458 (N_9458,N_870,N_1317);
and U9459 (N_9459,N_2280,N_769);
nand U9460 (N_9460,N_1519,N_4647);
nor U9461 (N_9461,N_82,N_516);
nor U9462 (N_9462,N_3558,N_925);
nand U9463 (N_9463,N_3389,N_1097);
or U9464 (N_9464,N_4143,N_1610);
nor U9465 (N_9465,N_4557,N_4121);
or U9466 (N_9466,N_1474,N_4045);
nand U9467 (N_9467,N_779,N_210);
and U9468 (N_9468,N_4206,N_3895);
or U9469 (N_9469,N_177,N_1817);
and U9470 (N_9470,N_1550,N_4080);
nor U9471 (N_9471,N_2817,N_2382);
or U9472 (N_9472,N_1914,N_4239);
nand U9473 (N_9473,N_3991,N_2885);
or U9474 (N_9474,N_790,N_1807);
and U9475 (N_9475,N_2512,N_4280);
nor U9476 (N_9476,N_1892,N_3821);
or U9477 (N_9477,N_1099,N_3640);
nor U9478 (N_9478,N_4461,N_4508);
xnor U9479 (N_9479,N_1568,N_4951);
and U9480 (N_9480,N_1666,N_990);
and U9481 (N_9481,N_4092,N_4973);
and U9482 (N_9482,N_4337,N_776);
or U9483 (N_9483,N_423,N_2890);
nor U9484 (N_9484,N_1485,N_4134);
xor U9485 (N_9485,N_2108,N_2291);
nand U9486 (N_9486,N_3338,N_1242);
and U9487 (N_9487,N_2100,N_3134);
nor U9488 (N_9488,N_3387,N_2637);
and U9489 (N_9489,N_3859,N_4269);
and U9490 (N_9490,N_4225,N_3609);
and U9491 (N_9491,N_3969,N_774);
and U9492 (N_9492,N_3454,N_1996);
xnor U9493 (N_9493,N_2577,N_3860);
nor U9494 (N_9494,N_1777,N_2482);
nand U9495 (N_9495,N_4547,N_1640);
or U9496 (N_9496,N_3084,N_855);
or U9497 (N_9497,N_2807,N_2768);
or U9498 (N_9498,N_3516,N_717);
and U9499 (N_9499,N_2524,N_4319);
or U9500 (N_9500,N_3837,N_4965);
and U9501 (N_9501,N_2913,N_1796);
xnor U9502 (N_9502,N_613,N_1791);
and U9503 (N_9503,N_4300,N_1034);
nand U9504 (N_9504,N_366,N_3425);
nor U9505 (N_9505,N_641,N_196);
nand U9506 (N_9506,N_686,N_2994);
or U9507 (N_9507,N_2336,N_4576);
nand U9508 (N_9508,N_1218,N_4302);
nand U9509 (N_9509,N_937,N_4731);
nand U9510 (N_9510,N_1529,N_4031);
nand U9511 (N_9511,N_961,N_2707);
nor U9512 (N_9512,N_982,N_113);
or U9513 (N_9513,N_1553,N_2208);
and U9514 (N_9514,N_2136,N_1728);
nand U9515 (N_9515,N_1240,N_3142);
and U9516 (N_9516,N_1619,N_3435);
nor U9517 (N_9517,N_2493,N_3952);
or U9518 (N_9518,N_2581,N_4775);
nor U9519 (N_9519,N_3323,N_803);
nand U9520 (N_9520,N_4217,N_106);
and U9521 (N_9521,N_1186,N_3471);
nand U9522 (N_9522,N_4245,N_1512);
and U9523 (N_9523,N_3597,N_2974);
nor U9524 (N_9524,N_4534,N_7);
nand U9525 (N_9525,N_2035,N_3112);
nand U9526 (N_9526,N_1297,N_753);
or U9527 (N_9527,N_3308,N_1120);
or U9528 (N_9528,N_1712,N_1096);
nor U9529 (N_9529,N_4993,N_4870);
nor U9530 (N_9530,N_4662,N_3045);
nor U9531 (N_9531,N_4736,N_2974);
or U9532 (N_9532,N_2915,N_3779);
nor U9533 (N_9533,N_2380,N_3359);
nand U9534 (N_9534,N_1938,N_1329);
nand U9535 (N_9535,N_1209,N_4433);
or U9536 (N_9536,N_1776,N_1059);
or U9537 (N_9537,N_1228,N_3570);
nand U9538 (N_9538,N_4164,N_3977);
and U9539 (N_9539,N_1170,N_134);
and U9540 (N_9540,N_334,N_4415);
nand U9541 (N_9541,N_1668,N_2623);
nand U9542 (N_9542,N_4740,N_1631);
and U9543 (N_9543,N_696,N_4836);
nand U9544 (N_9544,N_2691,N_1613);
nand U9545 (N_9545,N_3089,N_1160);
nand U9546 (N_9546,N_3744,N_49);
and U9547 (N_9547,N_329,N_733);
nor U9548 (N_9548,N_4682,N_3084);
or U9549 (N_9549,N_4799,N_4685);
or U9550 (N_9550,N_943,N_3468);
nand U9551 (N_9551,N_4826,N_4266);
or U9552 (N_9552,N_3308,N_2431);
nor U9553 (N_9553,N_4169,N_2263);
and U9554 (N_9554,N_775,N_4120);
and U9555 (N_9555,N_3152,N_2543);
nor U9556 (N_9556,N_1196,N_1027);
or U9557 (N_9557,N_1071,N_3258);
and U9558 (N_9558,N_2263,N_296);
nor U9559 (N_9559,N_1325,N_1777);
nand U9560 (N_9560,N_3237,N_4795);
nand U9561 (N_9561,N_1579,N_3150);
nor U9562 (N_9562,N_3242,N_4770);
nor U9563 (N_9563,N_2457,N_4677);
nand U9564 (N_9564,N_1744,N_626);
or U9565 (N_9565,N_2525,N_4523);
nand U9566 (N_9566,N_3683,N_4919);
and U9567 (N_9567,N_984,N_3329);
nor U9568 (N_9568,N_866,N_1229);
nand U9569 (N_9569,N_2848,N_4672);
nor U9570 (N_9570,N_2720,N_3751);
and U9571 (N_9571,N_934,N_2732);
and U9572 (N_9572,N_2127,N_3037);
nand U9573 (N_9573,N_1426,N_3562);
nand U9574 (N_9574,N_1693,N_2100);
nor U9575 (N_9575,N_3962,N_3495);
nand U9576 (N_9576,N_3988,N_2406);
or U9577 (N_9577,N_556,N_1296);
or U9578 (N_9578,N_4171,N_3565);
nor U9579 (N_9579,N_3278,N_1093);
nand U9580 (N_9580,N_410,N_4270);
nor U9581 (N_9581,N_3674,N_3417);
and U9582 (N_9582,N_274,N_2503);
nand U9583 (N_9583,N_2576,N_4525);
nand U9584 (N_9584,N_1802,N_1537);
nand U9585 (N_9585,N_1408,N_1220);
and U9586 (N_9586,N_4669,N_4700);
and U9587 (N_9587,N_1266,N_1611);
or U9588 (N_9588,N_1085,N_4665);
and U9589 (N_9589,N_2903,N_875);
xnor U9590 (N_9590,N_2216,N_1788);
xnor U9591 (N_9591,N_1511,N_1281);
or U9592 (N_9592,N_2453,N_2859);
and U9593 (N_9593,N_4447,N_2332);
nor U9594 (N_9594,N_2623,N_4555);
or U9595 (N_9595,N_2889,N_2151);
or U9596 (N_9596,N_1247,N_662);
or U9597 (N_9597,N_431,N_2522);
or U9598 (N_9598,N_3159,N_2667);
nor U9599 (N_9599,N_3992,N_1428);
xor U9600 (N_9600,N_3493,N_4959);
nor U9601 (N_9601,N_4491,N_3207);
or U9602 (N_9602,N_1952,N_3804);
nor U9603 (N_9603,N_4390,N_2059);
nand U9604 (N_9604,N_556,N_2270);
nand U9605 (N_9605,N_2528,N_2389);
and U9606 (N_9606,N_3865,N_1084);
or U9607 (N_9607,N_2931,N_560);
nand U9608 (N_9608,N_4614,N_1500);
nand U9609 (N_9609,N_2158,N_2136);
or U9610 (N_9610,N_3990,N_546);
nand U9611 (N_9611,N_2014,N_3245);
or U9612 (N_9612,N_1729,N_2283);
nand U9613 (N_9613,N_1867,N_4860);
and U9614 (N_9614,N_4683,N_1833);
and U9615 (N_9615,N_2781,N_213);
nor U9616 (N_9616,N_3542,N_1211);
or U9617 (N_9617,N_2365,N_1108);
and U9618 (N_9618,N_448,N_1667);
nor U9619 (N_9619,N_3267,N_1084);
or U9620 (N_9620,N_4910,N_2523);
or U9621 (N_9621,N_2819,N_2085);
nand U9622 (N_9622,N_933,N_2754);
nor U9623 (N_9623,N_2778,N_4224);
and U9624 (N_9624,N_2380,N_1667);
or U9625 (N_9625,N_1850,N_3880);
nand U9626 (N_9626,N_1386,N_4799);
nor U9627 (N_9627,N_3818,N_871);
or U9628 (N_9628,N_3154,N_1609);
xnor U9629 (N_9629,N_3118,N_1566);
and U9630 (N_9630,N_4364,N_1827);
or U9631 (N_9631,N_4051,N_4998);
nor U9632 (N_9632,N_4350,N_999);
and U9633 (N_9633,N_757,N_2312);
nor U9634 (N_9634,N_2941,N_3329);
or U9635 (N_9635,N_4467,N_4428);
and U9636 (N_9636,N_2240,N_4985);
nand U9637 (N_9637,N_1255,N_3425);
or U9638 (N_9638,N_3534,N_2070);
or U9639 (N_9639,N_1286,N_2235);
or U9640 (N_9640,N_339,N_1556);
or U9641 (N_9641,N_4208,N_4062);
nor U9642 (N_9642,N_4237,N_1922);
or U9643 (N_9643,N_4595,N_2132);
or U9644 (N_9644,N_1945,N_69);
nand U9645 (N_9645,N_4617,N_869);
or U9646 (N_9646,N_4923,N_3962);
nand U9647 (N_9647,N_1330,N_987);
nor U9648 (N_9648,N_2604,N_2741);
and U9649 (N_9649,N_628,N_2117);
or U9650 (N_9650,N_2715,N_4830);
or U9651 (N_9651,N_784,N_1346);
nor U9652 (N_9652,N_234,N_2536);
nand U9653 (N_9653,N_663,N_3287);
or U9654 (N_9654,N_2180,N_1836);
nand U9655 (N_9655,N_4215,N_2137);
and U9656 (N_9656,N_2241,N_4012);
or U9657 (N_9657,N_4982,N_2005);
and U9658 (N_9658,N_445,N_3099);
nor U9659 (N_9659,N_1691,N_3150);
or U9660 (N_9660,N_2523,N_451);
and U9661 (N_9661,N_1527,N_3216);
xor U9662 (N_9662,N_2653,N_3227);
and U9663 (N_9663,N_628,N_2552);
and U9664 (N_9664,N_1693,N_1887);
nand U9665 (N_9665,N_1949,N_2557);
nor U9666 (N_9666,N_3204,N_2661);
and U9667 (N_9667,N_4209,N_2416);
nand U9668 (N_9668,N_2237,N_644);
nand U9669 (N_9669,N_3782,N_1024);
nor U9670 (N_9670,N_3308,N_995);
xor U9671 (N_9671,N_1079,N_3770);
and U9672 (N_9672,N_1254,N_2146);
nor U9673 (N_9673,N_771,N_57);
and U9674 (N_9674,N_677,N_988);
and U9675 (N_9675,N_1185,N_4910);
nand U9676 (N_9676,N_1487,N_393);
nor U9677 (N_9677,N_430,N_1732);
nor U9678 (N_9678,N_2358,N_4857);
or U9679 (N_9679,N_3058,N_3983);
nor U9680 (N_9680,N_3978,N_3488);
nand U9681 (N_9681,N_1866,N_3599);
or U9682 (N_9682,N_1737,N_16);
nor U9683 (N_9683,N_4787,N_4581);
nand U9684 (N_9684,N_1002,N_1547);
or U9685 (N_9685,N_3875,N_1732);
nand U9686 (N_9686,N_1001,N_1723);
and U9687 (N_9687,N_906,N_869);
or U9688 (N_9688,N_891,N_3212);
nand U9689 (N_9689,N_3966,N_477);
nand U9690 (N_9690,N_880,N_2895);
nor U9691 (N_9691,N_2229,N_3719);
or U9692 (N_9692,N_4761,N_4559);
or U9693 (N_9693,N_4899,N_1470);
nor U9694 (N_9694,N_1118,N_4390);
or U9695 (N_9695,N_3181,N_1449);
nor U9696 (N_9696,N_199,N_2801);
nand U9697 (N_9697,N_3597,N_4158);
or U9698 (N_9698,N_4464,N_1463);
or U9699 (N_9699,N_671,N_3661);
or U9700 (N_9700,N_916,N_708);
nand U9701 (N_9701,N_258,N_4216);
or U9702 (N_9702,N_1578,N_2030);
nand U9703 (N_9703,N_2629,N_1465);
nand U9704 (N_9704,N_688,N_221);
nand U9705 (N_9705,N_1270,N_937);
nor U9706 (N_9706,N_1307,N_4335);
or U9707 (N_9707,N_2209,N_3441);
nand U9708 (N_9708,N_3489,N_2751);
nand U9709 (N_9709,N_2443,N_2988);
and U9710 (N_9710,N_1109,N_3519);
nor U9711 (N_9711,N_3572,N_4443);
nor U9712 (N_9712,N_3676,N_1438);
or U9713 (N_9713,N_1288,N_2593);
nand U9714 (N_9714,N_1280,N_4377);
or U9715 (N_9715,N_376,N_222);
and U9716 (N_9716,N_1944,N_407);
or U9717 (N_9717,N_4819,N_280);
and U9718 (N_9718,N_588,N_4606);
nand U9719 (N_9719,N_926,N_1807);
or U9720 (N_9720,N_1828,N_4);
nand U9721 (N_9721,N_129,N_2797);
nor U9722 (N_9722,N_1850,N_1956);
nor U9723 (N_9723,N_3402,N_3106);
and U9724 (N_9724,N_2921,N_3571);
nor U9725 (N_9725,N_2424,N_1861);
nor U9726 (N_9726,N_2170,N_2067);
or U9727 (N_9727,N_3509,N_4666);
nor U9728 (N_9728,N_2908,N_993);
nor U9729 (N_9729,N_4530,N_3270);
and U9730 (N_9730,N_4146,N_4107);
and U9731 (N_9731,N_689,N_1687);
nand U9732 (N_9732,N_2430,N_4341);
or U9733 (N_9733,N_2084,N_2160);
and U9734 (N_9734,N_964,N_2172);
or U9735 (N_9735,N_606,N_3348);
nand U9736 (N_9736,N_1060,N_671);
and U9737 (N_9737,N_4269,N_3848);
or U9738 (N_9738,N_3319,N_2860);
nor U9739 (N_9739,N_1308,N_802);
nand U9740 (N_9740,N_145,N_1297);
nor U9741 (N_9741,N_3470,N_2136);
nand U9742 (N_9742,N_722,N_4410);
and U9743 (N_9743,N_3636,N_3876);
nor U9744 (N_9744,N_1536,N_4254);
and U9745 (N_9745,N_1147,N_2863);
or U9746 (N_9746,N_4224,N_182);
nor U9747 (N_9747,N_222,N_1491);
nor U9748 (N_9748,N_3839,N_1559);
and U9749 (N_9749,N_3156,N_4721);
or U9750 (N_9750,N_2537,N_1281);
nand U9751 (N_9751,N_669,N_1223);
or U9752 (N_9752,N_2372,N_1754);
or U9753 (N_9753,N_600,N_3320);
or U9754 (N_9754,N_4372,N_1739);
and U9755 (N_9755,N_4420,N_4297);
nor U9756 (N_9756,N_1269,N_3829);
nand U9757 (N_9757,N_2708,N_445);
nor U9758 (N_9758,N_1651,N_486);
and U9759 (N_9759,N_3598,N_233);
or U9760 (N_9760,N_1556,N_2390);
and U9761 (N_9761,N_310,N_125);
and U9762 (N_9762,N_1732,N_3128);
nor U9763 (N_9763,N_1869,N_2280);
xor U9764 (N_9764,N_1478,N_4026);
or U9765 (N_9765,N_3228,N_2731);
or U9766 (N_9766,N_1866,N_3939);
and U9767 (N_9767,N_1313,N_4015);
xnor U9768 (N_9768,N_3596,N_1356);
or U9769 (N_9769,N_394,N_1981);
and U9770 (N_9770,N_303,N_4307);
or U9771 (N_9771,N_791,N_1092);
nand U9772 (N_9772,N_2208,N_1405);
nand U9773 (N_9773,N_2221,N_4862);
or U9774 (N_9774,N_2060,N_2378);
or U9775 (N_9775,N_298,N_1779);
xnor U9776 (N_9776,N_1608,N_1217);
nand U9777 (N_9777,N_1857,N_970);
nor U9778 (N_9778,N_1673,N_2988);
and U9779 (N_9779,N_1782,N_995);
and U9780 (N_9780,N_2267,N_182);
or U9781 (N_9781,N_470,N_4842);
and U9782 (N_9782,N_1236,N_3602);
and U9783 (N_9783,N_3308,N_4571);
xnor U9784 (N_9784,N_2502,N_2517);
nor U9785 (N_9785,N_1098,N_4431);
and U9786 (N_9786,N_3748,N_2316);
nor U9787 (N_9787,N_4209,N_516);
and U9788 (N_9788,N_4768,N_654);
and U9789 (N_9789,N_4675,N_2896);
nand U9790 (N_9790,N_4563,N_4145);
or U9791 (N_9791,N_3454,N_3902);
or U9792 (N_9792,N_2916,N_1850);
nor U9793 (N_9793,N_1686,N_4047);
or U9794 (N_9794,N_2932,N_2966);
and U9795 (N_9795,N_943,N_3607);
nor U9796 (N_9796,N_2136,N_714);
nand U9797 (N_9797,N_875,N_3543);
nand U9798 (N_9798,N_585,N_1948);
nand U9799 (N_9799,N_3837,N_3876);
or U9800 (N_9800,N_3482,N_1536);
or U9801 (N_9801,N_1191,N_2766);
nand U9802 (N_9802,N_2897,N_3874);
or U9803 (N_9803,N_1051,N_1424);
or U9804 (N_9804,N_4122,N_4738);
and U9805 (N_9805,N_3729,N_1311);
nor U9806 (N_9806,N_4736,N_2897);
or U9807 (N_9807,N_1269,N_1555);
nand U9808 (N_9808,N_2681,N_1966);
nand U9809 (N_9809,N_1284,N_1647);
nor U9810 (N_9810,N_494,N_3290);
nand U9811 (N_9811,N_4040,N_4324);
nand U9812 (N_9812,N_1082,N_430);
nand U9813 (N_9813,N_4760,N_1256);
nand U9814 (N_9814,N_1493,N_4759);
or U9815 (N_9815,N_4915,N_4051);
and U9816 (N_9816,N_1244,N_4264);
nand U9817 (N_9817,N_604,N_2155);
or U9818 (N_9818,N_3615,N_2078);
nand U9819 (N_9819,N_2860,N_1390);
or U9820 (N_9820,N_4827,N_675);
and U9821 (N_9821,N_2675,N_1077);
and U9822 (N_9822,N_2373,N_2628);
or U9823 (N_9823,N_738,N_4705);
or U9824 (N_9824,N_4203,N_1287);
nor U9825 (N_9825,N_3150,N_2698);
nor U9826 (N_9826,N_391,N_4240);
nor U9827 (N_9827,N_811,N_80);
and U9828 (N_9828,N_4042,N_2797);
nor U9829 (N_9829,N_1460,N_130);
nand U9830 (N_9830,N_1754,N_11);
and U9831 (N_9831,N_51,N_4724);
nand U9832 (N_9832,N_2854,N_4246);
nand U9833 (N_9833,N_592,N_1059);
nand U9834 (N_9834,N_4603,N_618);
nand U9835 (N_9835,N_4429,N_2538);
nor U9836 (N_9836,N_4655,N_4467);
and U9837 (N_9837,N_898,N_3740);
and U9838 (N_9838,N_233,N_374);
xnor U9839 (N_9839,N_942,N_2854);
nand U9840 (N_9840,N_2166,N_82);
or U9841 (N_9841,N_1436,N_2434);
and U9842 (N_9842,N_1765,N_216);
nand U9843 (N_9843,N_3109,N_4107);
or U9844 (N_9844,N_2870,N_1184);
and U9845 (N_9845,N_198,N_2345);
nand U9846 (N_9846,N_4959,N_4503);
nor U9847 (N_9847,N_1868,N_98);
or U9848 (N_9848,N_1028,N_1431);
and U9849 (N_9849,N_3303,N_3574);
nand U9850 (N_9850,N_4177,N_710);
or U9851 (N_9851,N_2279,N_1847);
or U9852 (N_9852,N_92,N_3643);
or U9853 (N_9853,N_4919,N_3656);
xnor U9854 (N_9854,N_2505,N_3666);
or U9855 (N_9855,N_1239,N_2555);
and U9856 (N_9856,N_2518,N_33);
or U9857 (N_9857,N_202,N_2863);
nor U9858 (N_9858,N_650,N_1829);
or U9859 (N_9859,N_1220,N_328);
nand U9860 (N_9860,N_750,N_917);
nor U9861 (N_9861,N_1187,N_4672);
nor U9862 (N_9862,N_837,N_902);
nand U9863 (N_9863,N_796,N_2080);
and U9864 (N_9864,N_312,N_1924);
or U9865 (N_9865,N_2382,N_4501);
and U9866 (N_9866,N_1338,N_2412);
nand U9867 (N_9867,N_2081,N_757);
and U9868 (N_9868,N_4243,N_853);
and U9869 (N_9869,N_1638,N_1452);
or U9870 (N_9870,N_993,N_649);
or U9871 (N_9871,N_99,N_2938);
nor U9872 (N_9872,N_2823,N_2291);
nor U9873 (N_9873,N_3505,N_3997);
nor U9874 (N_9874,N_1978,N_3772);
or U9875 (N_9875,N_3588,N_4614);
nand U9876 (N_9876,N_2069,N_1953);
or U9877 (N_9877,N_303,N_1409);
or U9878 (N_9878,N_1446,N_382);
or U9879 (N_9879,N_4922,N_1903);
and U9880 (N_9880,N_3603,N_483);
nand U9881 (N_9881,N_1208,N_4289);
nor U9882 (N_9882,N_2085,N_628);
nor U9883 (N_9883,N_823,N_711);
and U9884 (N_9884,N_872,N_795);
or U9885 (N_9885,N_2917,N_1715);
nand U9886 (N_9886,N_669,N_3333);
nor U9887 (N_9887,N_2740,N_109);
nand U9888 (N_9888,N_4257,N_361);
nand U9889 (N_9889,N_3861,N_4806);
or U9890 (N_9890,N_1201,N_2631);
nor U9891 (N_9891,N_3988,N_2984);
or U9892 (N_9892,N_4505,N_1275);
nor U9893 (N_9893,N_3963,N_953);
and U9894 (N_9894,N_4417,N_1103);
and U9895 (N_9895,N_3442,N_3915);
xor U9896 (N_9896,N_1100,N_4790);
and U9897 (N_9897,N_3079,N_2073);
nor U9898 (N_9898,N_2764,N_4792);
nor U9899 (N_9899,N_735,N_1880);
or U9900 (N_9900,N_2055,N_4707);
nor U9901 (N_9901,N_2380,N_2963);
nor U9902 (N_9902,N_1986,N_3132);
and U9903 (N_9903,N_871,N_3887);
nor U9904 (N_9904,N_3214,N_3809);
nor U9905 (N_9905,N_632,N_3498);
nor U9906 (N_9906,N_2276,N_1395);
nand U9907 (N_9907,N_973,N_3093);
or U9908 (N_9908,N_998,N_3886);
nor U9909 (N_9909,N_4574,N_1890);
nand U9910 (N_9910,N_1623,N_1330);
nor U9911 (N_9911,N_2923,N_4205);
or U9912 (N_9912,N_4341,N_2566);
nand U9913 (N_9913,N_512,N_613);
nor U9914 (N_9914,N_1405,N_4911);
nor U9915 (N_9915,N_433,N_2058);
nand U9916 (N_9916,N_4176,N_3754);
and U9917 (N_9917,N_4357,N_4306);
nor U9918 (N_9918,N_2861,N_704);
or U9919 (N_9919,N_999,N_4786);
nand U9920 (N_9920,N_214,N_1091);
nor U9921 (N_9921,N_4173,N_3081);
xor U9922 (N_9922,N_4891,N_3687);
nand U9923 (N_9923,N_1737,N_131);
nand U9924 (N_9924,N_2523,N_1127);
and U9925 (N_9925,N_3230,N_2659);
nand U9926 (N_9926,N_2062,N_3508);
and U9927 (N_9927,N_2122,N_4636);
and U9928 (N_9928,N_585,N_4109);
or U9929 (N_9929,N_1309,N_4020);
nand U9930 (N_9930,N_2501,N_1508);
and U9931 (N_9931,N_331,N_323);
nand U9932 (N_9932,N_3556,N_3696);
and U9933 (N_9933,N_3046,N_4360);
or U9934 (N_9934,N_1512,N_92);
nand U9935 (N_9935,N_749,N_2382);
nand U9936 (N_9936,N_3461,N_1200);
and U9937 (N_9937,N_3100,N_4329);
or U9938 (N_9938,N_263,N_3405);
and U9939 (N_9939,N_4645,N_2408);
nor U9940 (N_9940,N_3298,N_2848);
or U9941 (N_9941,N_2767,N_2937);
nor U9942 (N_9942,N_2282,N_4614);
and U9943 (N_9943,N_4863,N_4486);
or U9944 (N_9944,N_1912,N_4041);
nand U9945 (N_9945,N_4812,N_2743);
nor U9946 (N_9946,N_4177,N_126);
or U9947 (N_9947,N_2795,N_3760);
nor U9948 (N_9948,N_3968,N_3976);
nor U9949 (N_9949,N_4834,N_35);
nor U9950 (N_9950,N_1,N_3288);
and U9951 (N_9951,N_2879,N_4209);
nand U9952 (N_9952,N_2208,N_3784);
and U9953 (N_9953,N_622,N_2555);
nor U9954 (N_9954,N_2384,N_3016);
and U9955 (N_9955,N_1464,N_1914);
nand U9956 (N_9956,N_4298,N_1470);
nand U9957 (N_9957,N_4316,N_880);
nand U9958 (N_9958,N_1848,N_2558);
and U9959 (N_9959,N_96,N_239);
nand U9960 (N_9960,N_1066,N_1626);
or U9961 (N_9961,N_1201,N_2561);
nand U9962 (N_9962,N_2114,N_1404);
or U9963 (N_9963,N_955,N_2760);
and U9964 (N_9964,N_1664,N_984);
and U9965 (N_9965,N_4300,N_4265);
or U9966 (N_9966,N_738,N_42);
nor U9967 (N_9967,N_3689,N_1280);
nor U9968 (N_9968,N_103,N_222);
and U9969 (N_9969,N_750,N_2873);
xnor U9970 (N_9970,N_3916,N_3150);
and U9971 (N_9971,N_4736,N_4967);
and U9972 (N_9972,N_358,N_3656);
nand U9973 (N_9973,N_825,N_3051);
or U9974 (N_9974,N_958,N_4896);
nand U9975 (N_9975,N_1668,N_4823);
xor U9976 (N_9976,N_3633,N_2260);
nor U9977 (N_9977,N_1949,N_4208);
nor U9978 (N_9978,N_2217,N_27);
nand U9979 (N_9979,N_122,N_542);
and U9980 (N_9980,N_742,N_2121);
nor U9981 (N_9981,N_2852,N_4404);
nor U9982 (N_9982,N_2759,N_3379);
nor U9983 (N_9983,N_2529,N_2141);
nor U9984 (N_9984,N_2005,N_1621);
nor U9985 (N_9985,N_4140,N_4646);
and U9986 (N_9986,N_1568,N_1612);
nor U9987 (N_9987,N_3608,N_2038);
nor U9988 (N_9988,N_1016,N_358);
or U9989 (N_9989,N_1404,N_4257);
or U9990 (N_9990,N_210,N_1755);
and U9991 (N_9991,N_1271,N_1432);
xor U9992 (N_9992,N_3604,N_2860);
nand U9993 (N_9993,N_4757,N_1513);
or U9994 (N_9994,N_471,N_48);
and U9995 (N_9995,N_3964,N_84);
xor U9996 (N_9996,N_3899,N_1106);
and U9997 (N_9997,N_110,N_853);
and U9998 (N_9998,N_4425,N_4213);
and U9999 (N_9999,N_962,N_518);
or UO_0 (O_0,N_8979,N_6369);
and UO_1 (O_1,N_5949,N_9217);
nand UO_2 (O_2,N_5396,N_8101);
and UO_3 (O_3,N_6889,N_6033);
nor UO_4 (O_4,N_5716,N_6988);
and UO_5 (O_5,N_7960,N_9543);
and UO_6 (O_6,N_8581,N_7421);
and UO_7 (O_7,N_7236,N_7874);
nand UO_8 (O_8,N_9233,N_7533);
and UO_9 (O_9,N_5237,N_7402);
and UO_10 (O_10,N_8721,N_7870);
nand UO_11 (O_11,N_5824,N_6362);
and UO_12 (O_12,N_9979,N_9446);
nor UO_13 (O_13,N_7086,N_8245);
or UO_14 (O_14,N_7843,N_8593);
or UO_15 (O_15,N_6302,N_9262);
and UO_16 (O_16,N_6591,N_8433);
or UO_17 (O_17,N_7876,N_7329);
xnor UO_18 (O_18,N_7169,N_8076);
nor UO_19 (O_19,N_5791,N_6703);
and UO_20 (O_20,N_9824,N_8132);
nand UO_21 (O_21,N_8665,N_6566);
and UO_22 (O_22,N_7748,N_5991);
and UO_23 (O_23,N_5082,N_9925);
and UO_24 (O_24,N_8153,N_6247);
and UO_25 (O_25,N_9365,N_7644);
or UO_26 (O_26,N_6307,N_6572);
nand UO_27 (O_27,N_8779,N_6261);
nor UO_28 (O_28,N_9959,N_9159);
and UO_29 (O_29,N_7635,N_8464);
nand UO_30 (O_30,N_5461,N_6286);
nor UO_31 (O_31,N_5935,N_5581);
and UO_32 (O_32,N_5756,N_6767);
nor UO_33 (O_33,N_9278,N_6169);
nand UO_34 (O_34,N_9862,N_8940);
or UO_35 (O_35,N_6366,N_8919);
or UO_36 (O_36,N_7217,N_7336);
nand UO_37 (O_37,N_8297,N_9506);
and UO_38 (O_38,N_8074,N_5537);
or UO_39 (O_39,N_8009,N_8769);
or UO_40 (O_40,N_9668,N_9267);
nor UO_41 (O_41,N_7722,N_6221);
or UO_42 (O_42,N_8950,N_8482);
nand UO_43 (O_43,N_5902,N_7553);
nor UO_44 (O_44,N_9142,N_5897);
and UO_45 (O_45,N_5688,N_7377);
nor UO_46 (O_46,N_9508,N_6244);
nor UO_47 (O_47,N_9708,N_7199);
and UO_48 (O_48,N_7090,N_9151);
or UO_49 (O_49,N_9968,N_9647);
or UO_50 (O_50,N_9721,N_9438);
and UO_51 (O_51,N_7363,N_9333);
or UO_52 (O_52,N_8576,N_5334);
nand UO_53 (O_53,N_9081,N_9232);
and UO_54 (O_54,N_5706,N_6390);
or UO_55 (O_55,N_6877,N_7252);
or UO_56 (O_56,N_8641,N_7456);
nor UO_57 (O_57,N_8532,N_6742);
or UO_58 (O_58,N_8264,N_5435);
or UO_59 (O_59,N_8923,N_9753);
and UO_60 (O_60,N_9436,N_8107);
nand UO_61 (O_61,N_7404,N_7504);
or UO_62 (O_62,N_6167,N_6431);
or UO_63 (O_63,N_9252,N_9409);
xnor UO_64 (O_64,N_5227,N_8275);
nand UO_65 (O_65,N_5523,N_6330);
nand UO_66 (O_66,N_5649,N_8881);
nor UO_67 (O_67,N_8835,N_6250);
or UO_68 (O_68,N_9288,N_8172);
or UO_69 (O_69,N_6429,N_8765);
or UO_70 (O_70,N_8840,N_8333);
nand UO_71 (O_71,N_9105,N_8853);
nor UO_72 (O_72,N_9330,N_8423);
nand UO_73 (O_73,N_8303,N_8270);
nand UO_74 (O_74,N_6803,N_9226);
and UO_75 (O_75,N_6711,N_9241);
nor UO_76 (O_76,N_9903,N_5573);
and UO_77 (O_77,N_9879,N_6031);
nor UO_78 (O_78,N_8763,N_5731);
and UO_79 (O_79,N_5768,N_6718);
or UO_80 (O_80,N_8471,N_5369);
nor UO_81 (O_81,N_8796,N_7364);
and UO_82 (O_82,N_5661,N_6935);
or UO_83 (O_83,N_6149,N_7952);
and UO_84 (O_84,N_7743,N_7825);
nand UO_85 (O_85,N_8003,N_9440);
or UO_86 (O_86,N_6937,N_5878);
or UO_87 (O_87,N_5595,N_9191);
and UO_88 (O_88,N_6394,N_6065);
nor UO_89 (O_89,N_9421,N_9514);
or UO_90 (O_90,N_9189,N_7940);
and UO_91 (O_91,N_9738,N_9633);
nor UO_92 (O_92,N_8858,N_6683);
and UO_93 (O_93,N_8319,N_7557);
and UO_94 (O_94,N_9482,N_5597);
nand UO_95 (O_95,N_9162,N_8693);
and UO_96 (O_96,N_6507,N_8238);
nand UO_97 (O_97,N_5327,N_7758);
xnor UO_98 (O_98,N_9383,N_5676);
or UO_99 (O_99,N_5041,N_7712);
and UO_100 (O_100,N_5772,N_8239);
or UO_101 (O_101,N_5097,N_6246);
or UO_102 (O_102,N_6376,N_9125);
nor UO_103 (O_103,N_5978,N_5958);
and UO_104 (O_104,N_6562,N_9304);
or UO_105 (O_105,N_9507,N_6652);
and UO_106 (O_106,N_7450,N_7684);
and UO_107 (O_107,N_8951,N_5501);
or UO_108 (O_108,N_8300,N_6967);
nand UO_109 (O_109,N_9868,N_7446);
nand UO_110 (O_110,N_7076,N_7358);
and UO_111 (O_111,N_5497,N_5149);
and UO_112 (O_112,N_6229,N_9059);
or UO_113 (O_113,N_8887,N_8267);
and UO_114 (O_114,N_9133,N_6921);
nand UO_115 (O_115,N_7801,N_6207);
and UO_116 (O_116,N_5359,N_5083);
and UO_117 (O_117,N_7146,N_8903);
or UO_118 (O_118,N_6492,N_5663);
nand UO_119 (O_119,N_9951,N_9223);
nand UO_120 (O_120,N_8006,N_7859);
nor UO_121 (O_121,N_9788,N_8383);
xor UO_122 (O_122,N_7028,N_8805);
and UO_123 (O_123,N_5107,N_9521);
or UO_124 (O_124,N_6144,N_6318);
nor UO_125 (O_125,N_7137,N_5785);
nand UO_126 (O_126,N_6336,N_7772);
nor UO_127 (O_127,N_6327,N_8220);
or UO_128 (O_128,N_6470,N_5431);
and UO_129 (O_129,N_6345,N_9510);
nand UO_130 (O_130,N_5516,N_7079);
nor UO_131 (O_131,N_5728,N_5314);
nor UO_132 (O_132,N_7344,N_5637);
nand UO_133 (O_133,N_8515,N_6792);
nand UO_134 (O_134,N_8188,N_6373);
nor UO_135 (O_135,N_5952,N_9840);
and UO_136 (O_136,N_7820,N_8386);
nor UO_137 (O_137,N_9749,N_7560);
and UO_138 (O_138,N_9856,N_7800);
nand UO_139 (O_139,N_7389,N_7571);
and UO_140 (O_140,N_7341,N_7257);
nand UO_141 (O_141,N_5384,N_7755);
nand UO_142 (O_142,N_5410,N_9895);
nor UO_143 (O_143,N_7395,N_8806);
or UO_144 (O_144,N_8612,N_5889);
nand UO_145 (O_145,N_9695,N_9805);
and UO_146 (O_146,N_9572,N_7632);
xnor UO_147 (O_147,N_9042,N_5591);
nor UO_148 (O_148,N_5784,N_7045);
nor UO_149 (O_149,N_5631,N_6610);
and UO_150 (O_150,N_8705,N_8256);
nand UO_151 (O_151,N_9131,N_8589);
nor UO_152 (O_152,N_6177,N_7454);
nand UO_153 (O_153,N_8831,N_9764);
and UO_154 (O_154,N_7426,N_8616);
and UO_155 (O_155,N_6981,N_6191);
nor UO_156 (O_156,N_5158,N_8553);
xor UO_157 (O_157,N_6280,N_7115);
and UO_158 (O_158,N_5802,N_7905);
or UO_159 (O_159,N_5129,N_9311);
or UO_160 (O_160,N_9201,N_9718);
nand UO_161 (O_161,N_5152,N_7459);
xor UO_162 (O_162,N_9424,N_9816);
nand UO_163 (O_163,N_8167,N_8711);
nor UO_164 (O_164,N_6148,N_7597);
or UO_165 (O_165,N_5013,N_9161);
or UO_166 (O_166,N_6700,N_5858);
or UO_167 (O_167,N_7056,N_7925);
and UO_168 (O_168,N_8541,N_6795);
nor UO_169 (O_169,N_9571,N_5279);
or UO_170 (O_170,N_5941,N_5580);
or UO_171 (O_171,N_8056,N_8102);
nor UO_172 (O_172,N_9858,N_6186);
and UO_173 (O_173,N_6434,N_8041);
or UO_174 (O_174,N_7084,N_5912);
nand UO_175 (O_175,N_8223,N_5895);
or UO_176 (O_176,N_5634,N_7443);
nor UO_177 (O_177,N_6857,N_5504);
nor UO_178 (O_178,N_7166,N_6267);
or UO_179 (O_179,N_5686,N_6577);
nand UO_180 (O_180,N_5016,N_9564);
or UO_181 (O_181,N_8160,N_8224);
or UO_182 (O_182,N_9696,N_7305);
and UO_183 (O_183,N_9080,N_6759);
nand UO_184 (O_184,N_8993,N_9725);
nand UO_185 (O_185,N_9489,N_7039);
or UO_186 (O_186,N_8703,N_5172);
and UO_187 (O_187,N_5287,N_5293);
or UO_188 (O_188,N_5707,N_7243);
nand UO_189 (O_189,N_6090,N_5916);
nor UO_190 (O_190,N_8361,N_9643);
nor UO_191 (O_191,N_9882,N_9944);
nand UO_192 (O_192,N_8656,N_5040);
nand UO_193 (O_193,N_5989,N_5827);
nand UO_194 (O_194,N_5307,N_5252);
nand UO_195 (O_195,N_6242,N_6290);
nor UO_196 (O_196,N_6059,N_9209);
or UO_197 (O_197,N_9876,N_8856);
and UO_198 (O_198,N_8859,N_7883);
or UO_199 (O_199,N_5726,N_9836);
or UO_200 (O_200,N_7120,N_8370);
nand UO_201 (O_201,N_5179,N_8213);
nand UO_202 (O_202,N_7599,N_9070);
nand UO_203 (O_203,N_8533,N_6188);
nor UO_204 (O_204,N_8020,N_9040);
and UO_205 (O_205,N_6984,N_9634);
and UO_206 (O_206,N_8425,N_8653);
nand UO_207 (O_207,N_5363,N_6934);
nand UO_208 (O_208,N_9974,N_8566);
nor UO_209 (O_209,N_8897,N_5202);
and UO_210 (O_210,N_7240,N_5515);
nor UO_211 (O_211,N_8501,N_9605);
and UO_212 (O_212,N_5799,N_8271);
or UO_213 (O_213,N_6841,N_6162);
and UO_214 (O_214,N_6054,N_5062);
and UO_215 (O_215,N_5459,N_6717);
nor UO_216 (O_216,N_9274,N_5224);
or UO_217 (O_217,N_8755,N_5348);
nor UO_218 (O_218,N_7624,N_5727);
or UO_219 (O_219,N_6449,N_7078);
and UO_220 (O_220,N_5841,N_8373);
and UO_221 (O_221,N_8985,N_5930);
nor UO_222 (O_222,N_8643,N_7046);
nor UO_223 (O_223,N_8196,N_8842);
nand UO_224 (O_224,N_5965,N_6605);
nand UO_225 (O_225,N_5993,N_6198);
or UO_226 (O_226,N_7150,N_5052);
nand UO_227 (O_227,N_7666,N_7921);
and UO_228 (O_228,N_7927,N_8837);
and UO_229 (O_229,N_6740,N_8565);
nand UO_230 (O_230,N_9752,N_8594);
and UO_231 (O_231,N_6808,N_8659);
nor UO_232 (O_232,N_5692,N_9684);
nor UO_233 (O_233,N_8371,N_9362);
and UO_234 (O_234,N_9639,N_8442);
nor UO_235 (O_235,N_7152,N_9065);
nand UO_236 (O_236,N_5651,N_7912);
and UO_237 (O_237,N_9017,N_8269);
nand UO_238 (O_238,N_7982,N_5994);
and UO_239 (O_239,N_8149,N_8427);
nand UO_240 (O_240,N_8084,N_6420);
and UO_241 (O_241,N_7623,N_9327);
and UO_242 (O_242,N_9577,N_6046);
nand UO_243 (O_243,N_5406,N_7068);
nor UO_244 (O_244,N_9670,N_8709);
xor UO_245 (O_245,N_5366,N_8935);
and UO_246 (O_246,N_6611,N_8323);
xnor UO_247 (O_247,N_5980,N_9272);
and UO_248 (O_248,N_8799,N_9989);
or UO_249 (O_249,N_5429,N_7251);
nand UO_250 (O_250,N_9594,N_5923);
and UO_251 (O_251,N_6209,N_9030);
nor UO_252 (O_252,N_9686,N_8480);
nor UO_253 (O_253,N_9320,N_6077);
nor UO_254 (O_254,N_7384,N_5301);
nand UO_255 (O_255,N_8699,N_9891);
nand UO_256 (O_256,N_5191,N_5722);
and UO_257 (O_257,N_6108,N_5351);
nor UO_258 (O_258,N_7824,N_9911);
nand UO_259 (O_259,N_6707,N_6498);
or UO_260 (O_260,N_9978,N_6404);
nand UO_261 (O_261,N_7027,N_8100);
and UO_262 (O_262,N_7142,N_6453);
and UO_263 (O_263,N_9427,N_5423);
or UO_264 (O_264,N_5975,N_7953);
and UO_265 (O_265,N_8850,N_8405);
nor UO_266 (O_266,N_9908,N_9047);
xnor UO_267 (O_267,N_9529,N_8684);
nand UO_268 (O_268,N_5848,N_6796);
or UO_269 (O_269,N_9385,N_8393);
or UO_270 (O_270,N_9098,N_6002);
nand UO_271 (O_271,N_6102,N_9039);
and UO_272 (O_272,N_7822,N_5639);
and UO_273 (O_273,N_7873,N_6617);
nand UO_274 (O_274,N_8816,N_5166);
nand UO_275 (O_275,N_8868,N_6416);
nor UO_276 (O_276,N_8675,N_8946);
and UO_277 (O_277,N_7269,N_6216);
and UO_278 (O_278,N_5161,N_5102);
or UO_279 (O_279,N_8322,N_6650);
nor UO_280 (O_280,N_5373,N_5701);
or UO_281 (O_281,N_6654,N_9784);
and UO_282 (O_282,N_8986,N_6526);
nand UO_283 (O_283,N_8955,N_9261);
and UO_284 (O_284,N_7819,N_9905);
nand UO_285 (O_285,N_7962,N_8775);
nand UO_286 (O_286,N_7531,N_9181);
or UO_287 (O_287,N_5517,N_6061);
and UO_288 (O_288,N_5818,N_6490);
nor UO_289 (O_289,N_9803,N_6159);
nor UO_290 (O_290,N_7810,N_7091);
xnor UO_291 (O_291,N_7815,N_7841);
nand UO_292 (O_292,N_7528,N_6398);
or UO_293 (O_293,N_7225,N_8141);
nor UO_294 (O_294,N_9986,N_9192);
or UO_295 (O_295,N_5682,N_7609);
nor UO_296 (O_296,N_6530,N_6713);
or UO_297 (O_297,N_6051,N_6866);
nor UO_298 (O_298,N_9126,N_6294);
xor UO_299 (O_299,N_7737,N_8970);
nor UO_300 (O_300,N_5766,N_5583);
and UO_301 (O_301,N_7136,N_9539);
and UO_302 (O_302,N_8683,N_5472);
and UO_303 (O_303,N_5266,N_7832);
nor UO_304 (O_304,N_8580,N_7787);
and UO_305 (O_305,N_8920,N_5554);
and UO_306 (O_306,N_8522,N_7193);
and UO_307 (O_307,N_7019,N_7203);
or UO_308 (O_308,N_7963,N_8750);
nor UO_309 (O_309,N_6953,N_5807);
nor UO_310 (O_310,N_6377,N_8272);
and UO_311 (O_311,N_8745,N_7176);
or UO_312 (O_312,N_9516,N_9992);
nand UO_313 (O_313,N_9407,N_9560);
nor UO_314 (O_314,N_5112,N_8928);
nand UO_315 (O_315,N_8385,N_5896);
nor UO_316 (O_316,N_7968,N_7435);
nor UO_317 (O_317,N_6608,N_7971);
and UO_318 (O_318,N_6231,N_8800);
nor UO_319 (O_319,N_5934,N_6137);
and UO_320 (O_320,N_6777,N_5590);
nand UO_321 (O_321,N_5913,N_7995);
nor UO_322 (O_322,N_9100,N_8600);
or UO_323 (O_323,N_9437,N_5925);
or UO_324 (O_324,N_6880,N_9088);
and UO_325 (O_325,N_6779,N_7965);
or UO_326 (O_326,N_5561,N_7309);
nor UO_327 (O_327,N_8441,N_5608);
xnor UO_328 (O_328,N_9687,N_5270);
and UO_329 (O_329,N_5338,N_8191);
and UO_330 (O_330,N_5263,N_9214);
nand UO_331 (O_331,N_7584,N_5641);
and UO_332 (O_332,N_9839,N_5255);
or UO_333 (O_333,N_9674,N_9745);
or UO_334 (O_334,N_5236,N_7161);
and UO_335 (O_335,N_8134,N_7029);
nor UO_336 (O_336,N_8921,N_6641);
nand UO_337 (O_337,N_9473,N_8866);
nor UO_338 (O_338,N_9225,N_5687);
and UO_339 (O_339,N_7768,N_5817);
nand UO_340 (O_340,N_5335,N_7319);
or UO_341 (O_341,N_7696,N_5921);
and UO_342 (O_342,N_6933,N_7837);
or UO_343 (O_343,N_9342,N_5806);
or UO_344 (O_344,N_5260,N_6821);
or UO_345 (O_345,N_8915,N_8730);
and UO_346 (O_346,N_9820,N_8652);
nand UO_347 (O_347,N_7659,N_9294);
or UO_348 (O_348,N_9747,N_8157);
nand UO_349 (O_349,N_7299,N_9254);
or UO_350 (O_350,N_5028,N_8378);
xor UO_351 (O_351,N_9505,N_8590);
nor UO_352 (O_352,N_8926,N_8013);
and UO_353 (O_353,N_9022,N_6949);
or UO_354 (O_354,N_5049,N_9380);
and UO_355 (O_355,N_7101,N_7865);
or UO_356 (O_356,N_5108,N_7186);
and UO_357 (O_357,N_9555,N_7174);
nand UO_358 (O_358,N_8391,N_9283);
nand UO_359 (O_359,N_6311,N_5006);
nand UO_360 (O_360,N_9980,N_9432);
or UO_361 (O_361,N_9512,N_6830);
nor UO_362 (O_362,N_7324,N_6657);
and UO_363 (O_363,N_9425,N_6747);
nor UO_364 (O_364,N_5466,N_6262);
and UO_365 (O_365,N_8889,N_7525);
or UO_366 (O_366,N_6252,N_6359);
nor UO_367 (O_367,N_6271,N_9822);
nor UO_368 (O_368,N_8793,N_9907);
nor UO_369 (O_369,N_6248,N_9650);
nand UO_370 (O_370,N_7283,N_5098);
nand UO_371 (O_371,N_6043,N_5759);
nand UO_372 (O_372,N_8045,N_9912);
nor UO_373 (O_373,N_6133,N_5340);
or UO_374 (O_374,N_6797,N_8636);
nor UO_375 (O_375,N_6491,N_8714);
nor UO_376 (O_376,N_6638,N_6210);
or UO_377 (O_377,N_9459,N_5380);
or UO_378 (O_378,N_6472,N_8552);
and UO_379 (O_379,N_7219,N_6279);
nand UO_380 (O_380,N_5222,N_7407);
nor UO_381 (O_381,N_9336,N_6460);
xor UO_382 (O_382,N_9878,N_6999);
and UO_383 (O_383,N_9266,N_8389);
xor UO_384 (O_384,N_7907,N_5578);
nor UO_385 (O_385,N_8343,N_5213);
nor UO_386 (O_386,N_6706,N_8731);
nor UO_387 (O_387,N_7228,N_8424);
and UO_388 (O_388,N_8626,N_9293);
nand UO_389 (O_389,N_9163,N_6556);
nor UO_390 (O_390,N_9682,N_6092);
and UO_391 (O_391,N_8771,N_6097);
nor UO_392 (O_392,N_6426,N_7569);
nor UO_393 (O_393,N_9183,N_5710);
nand UO_394 (O_394,N_9689,N_7185);
nand UO_395 (O_395,N_9503,N_7158);
nand UO_396 (O_396,N_8688,N_8225);
nor UO_397 (O_397,N_6213,N_5058);
and UO_398 (O_398,N_6128,N_5027);
and UO_399 (O_399,N_8492,N_5265);
and UO_400 (O_400,N_6423,N_9522);
and UO_401 (O_401,N_5942,N_5449);
nand UO_402 (O_402,N_8432,N_7479);
or UO_403 (O_403,N_5919,N_7556);
and UO_404 (O_404,N_7314,N_9534);
nor UO_405 (O_405,N_9073,N_5821);
and UO_406 (O_406,N_9137,N_5683);
nand UO_407 (O_407,N_9298,N_7213);
or UO_408 (O_408,N_6926,N_9949);
and UO_409 (O_409,N_9200,N_8161);
nand UO_410 (O_410,N_9468,N_9476);
or UO_411 (O_411,N_6755,N_7049);
or UO_412 (O_412,N_9210,N_7445);
nor UO_413 (O_413,N_7725,N_5903);
nand UO_414 (O_414,N_8106,N_6537);
and UO_415 (O_415,N_6201,N_7035);
or UO_416 (O_416,N_5375,N_9664);
and UO_417 (O_417,N_9110,N_8820);
and UO_418 (O_418,N_8379,N_6528);
or UO_419 (O_419,N_6337,N_8824);
nor UO_420 (O_420,N_9276,N_8209);
or UO_421 (O_421,N_6884,N_9203);
and UO_422 (O_422,N_6299,N_7495);
and UO_423 (O_423,N_6892,N_5709);
nor UO_424 (O_424,N_9082,N_8570);
or UO_425 (O_425,N_8934,N_6275);
nand UO_426 (O_426,N_8283,N_5568);
or UO_427 (O_427,N_6313,N_5001);
nand UO_428 (O_428,N_5485,N_9826);
nand UO_429 (O_429,N_5283,N_8890);
or UO_430 (O_430,N_5051,N_7750);
nand UO_431 (O_431,N_5664,N_6558);
or UO_432 (O_432,N_5267,N_6833);
xor UO_433 (O_433,N_6098,N_7596);
nor UO_434 (O_434,N_6687,N_5215);
nor UO_435 (O_435,N_6485,N_5690);
nor UO_436 (O_436,N_9370,N_9319);
nand UO_437 (O_437,N_6397,N_6352);
or UO_438 (O_438,N_9626,N_5014);
nor UO_439 (O_439,N_6936,N_6588);
and UO_440 (O_440,N_6073,N_8024);
nor UO_441 (O_441,N_6752,N_7325);
and UO_442 (O_442,N_6818,N_7429);
nand UO_443 (O_443,N_5086,N_5600);
or UO_444 (O_444,N_9896,N_5046);
nor UO_445 (O_445,N_5090,N_5387);
and UO_446 (O_446,N_8304,N_5189);
nor UO_447 (O_447,N_5737,N_7694);
nand UO_448 (O_448,N_8154,N_5182);
nand UO_449 (O_449,N_5869,N_9874);
and UO_450 (O_450,N_8320,N_5636);
nand UO_451 (O_451,N_5966,N_5160);
nor UO_452 (O_452,N_6415,N_9917);
nand UO_453 (O_453,N_5996,N_9631);
and UO_454 (O_454,N_6199,N_8963);
and UO_455 (O_455,N_9453,N_8764);
or UO_456 (O_456,N_9953,N_5196);
nor UO_457 (O_457,N_9230,N_7579);
and UO_458 (O_458,N_9118,N_6673);
or UO_459 (O_459,N_5496,N_5899);
and UO_460 (O_460,N_7785,N_7582);
nor UO_461 (O_461,N_8156,N_7945);
nor UO_462 (O_462,N_7272,N_9601);
or UO_463 (O_463,N_6789,N_6563);
and UO_464 (O_464,N_7262,N_9545);
or UO_465 (O_465,N_7537,N_5801);
and UO_466 (O_466,N_7040,N_9454);
nand UO_467 (O_467,N_8218,N_9335);
and UO_468 (O_468,N_6200,N_9569);
and UO_469 (O_469,N_8344,N_6075);
nor UO_470 (O_470,N_9024,N_6726);
or UO_471 (O_471,N_7671,N_7653);
or UO_472 (O_472,N_8097,N_5383);
nor UO_473 (O_473,N_7390,N_6625);
nor UO_474 (O_474,N_7226,N_8757);
and UO_475 (O_475,N_7719,N_8354);
or UO_476 (O_476,N_9711,N_9158);
and UO_477 (O_477,N_6804,N_7096);
xor UO_478 (O_478,N_5330,N_9646);
nand UO_479 (O_479,N_9263,N_6419);
or UO_480 (O_480,N_8548,N_9838);
nor UO_481 (O_481,N_9871,N_9072);
nand UO_482 (O_482,N_5368,N_5938);
or UO_483 (O_483,N_8147,N_6517);
nor UO_484 (O_484,N_8095,N_8011);
nor UO_485 (O_485,N_5456,N_7451);
nor UO_486 (O_486,N_6754,N_7440);
or UO_487 (O_487,N_8529,N_7187);
xor UO_488 (O_488,N_9443,N_5810);
and UO_489 (O_489,N_7351,N_8706);
nor UO_490 (O_490,N_9921,N_7189);
or UO_491 (O_491,N_7220,N_7254);
and UO_492 (O_492,N_9617,N_6545);
xor UO_493 (O_493,N_5615,N_8374);
nor UO_494 (O_494,N_7458,N_8110);
nor UO_495 (O_495,N_6353,N_9374);
and UO_496 (O_496,N_9754,N_8166);
or UO_497 (O_497,N_8178,N_8353);
or UO_498 (O_498,N_7474,N_6206);
or UO_499 (O_499,N_7833,N_8395);
nor UO_500 (O_500,N_7598,N_8788);
and UO_501 (O_501,N_8292,N_7904);
and UO_502 (O_502,N_9958,N_8143);
nand UO_503 (O_503,N_5719,N_9596);
nand UO_504 (O_504,N_5592,N_7542);
and UO_505 (O_505,N_9352,N_6195);
nand UO_506 (O_506,N_6270,N_6447);
nand UO_507 (O_507,N_6698,N_8766);
nand UO_508 (O_508,N_8217,N_5240);
or UO_509 (O_509,N_6793,N_6595);
nor UO_510 (O_510,N_5199,N_9005);
nand UO_511 (O_511,N_5490,N_6996);
nand UO_512 (O_512,N_6913,N_9852);
nor UO_513 (O_513,N_7036,N_9593);
or UO_514 (O_514,N_9041,N_7909);
nor UO_515 (O_515,N_9216,N_5851);
or UO_516 (O_516,N_6235,N_6619);
nor UO_517 (O_517,N_7881,N_8598);
nand UO_518 (O_518,N_6770,N_5769);
or UO_519 (O_519,N_7061,N_8728);
and UO_520 (O_520,N_6987,N_7861);
and UO_521 (O_521,N_8782,N_5574);
and UO_522 (O_522,N_7930,N_6568);
and UO_523 (O_523,N_8211,N_9970);
nor UO_524 (O_524,N_9472,N_8628);
and UO_525 (O_525,N_5681,N_6350);
and UO_526 (O_526,N_7742,N_6281);
nor UO_527 (O_527,N_6406,N_6859);
and UO_528 (O_528,N_8250,N_8847);
or UO_529 (O_529,N_5657,N_9984);
and UO_530 (O_530,N_5447,N_8342);
nand UO_531 (O_531,N_9597,N_5282);
nor UO_532 (O_532,N_8384,N_7562);
nand UO_533 (O_533,N_6664,N_5742);
or UO_534 (O_534,N_8136,N_6041);
nand UO_535 (O_535,N_6672,N_9045);
nand UO_536 (O_536,N_9056,N_8929);
nor UO_537 (O_537,N_9627,N_6237);
nor UO_538 (O_538,N_9186,N_6539);
and UO_539 (O_539,N_8968,N_8192);
nor UO_540 (O_540,N_8436,N_8954);
nor UO_541 (O_541,N_6761,N_7172);
or UO_542 (O_542,N_7268,N_6741);
nand UO_543 (O_543,N_9077,N_8927);
nor UO_544 (O_544,N_5655,N_7882);
nand UO_545 (O_545,N_5866,N_7288);
nor UO_546 (O_546,N_9782,N_6646);
xor UO_547 (O_547,N_6565,N_9463);
nor UO_548 (O_548,N_8826,N_5473);
or UO_549 (O_549,N_7880,N_7475);
nand UO_550 (O_550,N_8666,N_7846);
or UO_551 (O_551,N_7898,N_9060);
nand UO_552 (O_552,N_8719,N_9574);
nand UO_553 (O_553,N_9735,N_7924);
nand UO_554 (O_554,N_8004,N_9685);
or UO_555 (O_555,N_7724,N_6737);
nor UO_556 (O_556,N_7729,N_7333);
nor UO_557 (O_557,N_9699,N_6962);
nand UO_558 (O_558,N_9566,N_7042);
nor UO_559 (O_559,N_6659,N_7778);
nand UO_560 (O_560,N_9511,N_9598);
or UO_561 (O_561,N_6685,N_5572);
or UO_562 (O_562,N_6335,N_8702);
and UO_563 (O_563,N_7196,N_8822);
nand UO_564 (O_564,N_7655,N_9099);
nor UO_565 (O_565,N_7627,N_6994);
or UO_566 (O_566,N_8242,N_6955);
nor UO_567 (O_567,N_5816,N_9389);
nand UO_568 (O_568,N_9635,N_9930);
and UO_569 (O_569,N_8049,N_8689);
nand UO_570 (O_570,N_7552,N_8390);
nor UO_571 (O_571,N_7987,N_6442);
and UO_572 (O_572,N_6760,N_5395);
nor UO_573 (O_573,N_5783,N_7503);
and UO_574 (O_574,N_9354,N_7799);
and UO_575 (O_575,N_7093,N_8294);
or UO_576 (O_576,N_6395,N_9413);
or UO_577 (O_577,N_7295,N_9676);
and UO_578 (O_578,N_9393,N_5735);
xor UO_579 (O_579,N_6630,N_8263);
nand UO_580 (O_580,N_9498,N_5929);
nor UO_581 (O_581,N_9844,N_8618);
nor UO_582 (O_582,N_9085,N_9014);
or UO_583 (O_583,N_7053,N_8276);
and UO_584 (O_584,N_5969,N_5017);
nor UO_585 (O_585,N_8933,N_9168);
nor UO_586 (O_586,N_6917,N_7327);
or UO_587 (O_587,N_9355,N_8495);
nor UO_588 (O_588,N_6719,N_9860);
or UO_589 (O_589,N_5920,N_9548);
nor UO_590 (O_590,N_5880,N_9999);
or UO_591 (O_591,N_6405,N_5788);
nor UO_592 (O_592,N_6438,N_9902);
and UO_593 (O_593,N_7985,N_9090);
nand UO_594 (O_594,N_7530,N_7679);
xnor UO_595 (O_595,N_5141,N_9845);
or UO_596 (O_596,N_9751,N_7978);
and UO_597 (O_597,N_7369,N_6348);
nand UO_598 (O_598,N_5217,N_9124);
nor UO_599 (O_599,N_6251,N_6511);
and UO_600 (O_600,N_6298,N_8028);
or UO_601 (O_601,N_6466,N_6096);
or UO_602 (O_602,N_9557,N_7949);
xnor UO_603 (O_603,N_5436,N_8620);
nor UO_604 (O_604,N_7178,N_8609);
and UO_605 (O_605,N_9649,N_5111);
xnor UO_606 (O_606,N_5365,N_9706);
nor UO_607 (O_607,N_8232,N_5274);
nor UO_608 (O_608,N_9579,N_9870);
nor UO_609 (O_609,N_8647,N_5875);
and UO_610 (O_610,N_8284,N_6482);
nand UO_611 (O_611,N_6071,N_6746);
and UO_612 (O_612,N_6037,N_7480);
nand UO_613 (O_613,N_6204,N_5493);
or UO_614 (O_614,N_7687,N_8642);
xnor UO_615 (O_615,N_9755,N_6871);
nand UO_616 (O_616,N_5462,N_9416);
nand UO_617 (O_617,N_6003,N_5891);
nor UO_618 (O_618,N_6541,N_7069);
nor UO_619 (O_619,N_5594,N_7567);
or UO_620 (O_620,N_8981,N_7678);
and UO_621 (O_621,N_6822,N_5342);
nor UO_622 (O_622,N_8679,N_7681);
and UO_623 (O_623,N_7011,N_5022);
nand UO_624 (O_624,N_5355,N_8854);
nor UO_625 (O_625,N_9196,N_8090);
and UO_626 (O_626,N_6399,N_8623);
nand UO_627 (O_627,N_5535,N_9589);
nand UO_628 (O_628,N_9390,N_6142);
and UO_629 (O_629,N_8054,N_6553);
or UO_630 (O_630,N_8372,N_8470);
or UO_631 (O_631,N_6751,N_7055);
and UO_632 (O_632,N_6998,N_7807);
or UO_633 (O_633,N_8302,N_9337);
and UO_634 (O_634,N_9957,N_5494);
and UO_635 (O_635,N_9198,N_9928);
nor UO_636 (O_636,N_9734,N_8561);
nand UO_637 (O_637,N_7796,N_8059);
or UO_638 (O_638,N_5394,N_8739);
or UO_639 (O_639,N_8111,N_5489);
nand UO_640 (O_640,N_6047,N_5671);
nand UO_641 (O_641,N_8259,N_7103);
and UO_642 (O_642,N_7326,N_6131);
and UO_643 (O_643,N_9205,N_8958);
nor UO_644 (O_644,N_7568,N_7918);
nor UO_645 (O_645,N_6219,N_6674);
nand UO_646 (O_646,N_6058,N_7948);
nand UO_647 (O_647,N_9306,N_9258);
or UO_648 (O_648,N_6074,N_7195);
nor UO_649 (O_649,N_8340,N_7897);
nor UO_650 (O_650,N_7469,N_5855);
or UO_651 (O_651,N_7818,N_5453);
nor UO_652 (O_652,N_5415,N_8130);
nor UO_653 (O_653,N_6001,N_5886);
xnor UO_654 (O_654,N_8525,N_6836);
nor UO_655 (O_655,N_6493,N_6205);
and UO_656 (O_656,N_5020,N_9843);
nor UO_657 (O_657,N_7455,N_9495);
nand UO_658 (O_658,N_7134,N_8603);
and UO_659 (O_659,N_5749,N_7500);
and UO_660 (O_660,N_8261,N_6124);
nand UO_661 (O_661,N_5566,N_9817);
nand UO_662 (O_662,N_6042,N_7767);
nand UO_663 (O_663,N_8037,N_5770);
and UO_664 (O_664,N_5029,N_8588);
nor UO_665 (O_665,N_5377,N_9069);
nand UO_666 (O_666,N_9260,N_6916);
or UO_667 (O_667,N_8936,N_7463);
nand UO_668 (O_668,N_8852,N_8124);
and UO_669 (O_669,N_6379,N_6139);
nand UO_670 (O_670,N_8645,N_8734);
and UO_671 (O_671,N_6243,N_7770);
nand UO_672 (O_672,N_5757,N_9128);
and UO_673 (O_673,N_6766,N_6529);
nor UO_674 (O_674,N_6441,N_5445);
and UO_675 (O_675,N_9947,N_8352);
nor UO_676 (O_676,N_5065,N_5246);
nand UO_677 (O_677,N_5571,N_7845);
or UO_678 (O_678,N_9229,N_9693);
and UO_679 (O_679,N_8406,N_7082);
and UO_680 (O_680,N_6109,N_9910);
and UO_681 (O_681,N_7895,N_7348);
nand UO_682 (O_682,N_9667,N_8549);
xor UO_683 (O_683,N_7140,N_5977);
nor UO_684 (O_684,N_5642,N_9883);
or UO_685 (O_685,N_6695,N_6677);
and UO_686 (O_686,N_5219,N_5048);
nand UO_687 (O_687,N_7110,N_7603);
nor UO_688 (O_688,N_6848,N_7063);
xnor UO_689 (O_689,N_7581,N_6222);
nand UO_690 (O_690,N_7776,N_7608);
nand UO_691 (O_691,N_9368,N_7752);
and UO_692 (O_692,N_6354,N_5559);
nor UO_693 (O_693,N_9280,N_5853);
and UO_694 (O_694,N_8376,N_9867);
or UO_695 (O_695,N_7282,N_6820);
and UO_696 (O_696,N_6970,N_6501);
or UO_697 (O_697,N_5840,N_5209);
and UO_698 (O_698,N_8965,N_7587);
nand UO_699 (O_699,N_6499,N_9392);
nand UO_700 (O_700,N_6784,N_8058);
nand UO_701 (O_701,N_8219,N_6634);
nor UO_702 (O_702,N_9558,N_9541);
nand UO_703 (O_703,N_9873,N_9950);
xnor UO_704 (O_704,N_5238,N_9250);
or UO_705 (O_705,N_9236,N_5843);
nor UO_706 (O_706,N_6138,N_6383);
nor UO_707 (O_707,N_9265,N_7200);
xnor UO_708 (O_708,N_7313,N_8321);
and UO_709 (O_709,N_8328,N_7153);
nand UO_710 (O_710,N_6518,N_5185);
nor UO_711 (O_711,N_6032,N_9079);
nand UO_712 (O_712,N_5987,N_8168);
nand UO_713 (O_713,N_9717,N_5542);
nand UO_714 (O_714,N_9769,N_9051);
or UO_715 (O_715,N_5990,N_9760);
nand UO_716 (O_716,N_9094,N_8531);
and UO_717 (O_717,N_5842,N_7018);
xor UO_718 (O_718,N_8885,N_9991);
nand UO_719 (O_719,N_9012,N_8843);
nand UO_720 (O_720,N_7099,N_6557);
xnor UO_721 (O_721,N_6328,N_8040);
nor UO_722 (O_722,N_9264,N_9743);
nand UO_723 (O_723,N_8025,N_7676);
nand UO_724 (O_724,N_6932,N_6739);
or UO_725 (O_725,N_8438,N_9884);
and UO_726 (O_726,N_6851,N_5964);
and UO_727 (O_727,N_6874,N_9640);
and UO_728 (O_728,N_9898,N_6488);
nand UO_729 (O_729,N_6048,N_5518);
nand UO_730 (O_730,N_9026,N_9532);
nor UO_731 (O_731,N_6029,N_9790);
or UO_732 (O_732,N_7002,N_8687);
or UO_733 (O_733,N_8610,N_5943);
nand UO_734 (O_734,N_8158,N_6110);
nand UO_735 (O_735,N_9386,N_6669);
or UO_736 (O_736,N_8611,N_5230);
or UO_737 (O_737,N_8216,N_9006);
and UO_738 (O_738,N_8065,N_6412);
and UO_739 (O_739,N_5003,N_9307);
and UO_740 (O_740,N_7991,N_9602);
nor UO_741 (O_741,N_7374,N_8131);
or UO_742 (O_742,N_6644,N_5820);
or UO_743 (O_743,N_6855,N_5063);
nand UO_744 (O_744,N_9952,N_5695);
or UO_745 (O_745,N_8942,N_7774);
nand UO_746 (O_746,N_7419,N_7160);
and UO_747 (O_747,N_7779,N_6268);
nand UO_748 (O_748,N_5125,N_9945);
nor UO_749 (O_749,N_7113,N_5474);
nand UO_750 (O_750,N_8296,N_7518);
or UO_751 (O_751,N_7009,N_8285);
or UO_752 (O_752,N_9691,N_5280);
nor UO_753 (O_753,N_5705,N_5164);
nor UO_754 (O_754,N_7216,N_6505);
and UO_755 (O_755,N_7735,N_7320);
nand UO_756 (O_756,N_7311,N_6860);
nand UO_757 (O_757,N_5643,N_7230);
nor UO_758 (O_758,N_5352,N_7397);
nand UO_759 (O_759,N_7836,N_6208);
nand UO_760 (O_760,N_6941,N_9247);
nand UO_761 (O_761,N_5220,N_7616);
xnor UO_762 (O_762,N_5519,N_8697);
nor UO_763 (O_763,N_5606,N_6951);
nor UO_764 (O_764,N_9955,N_5834);
nor UO_765 (O_765,N_8366,N_7929);
and UO_766 (O_766,N_8901,N_7376);
or UO_767 (O_767,N_9075,N_5849);
nor UO_768 (O_768,N_9702,N_8474);
and UO_769 (O_769,N_5915,N_9943);
and UO_770 (O_770,N_6481,N_5741);
nand UO_771 (O_771,N_5463,N_5060);
and UO_772 (O_772,N_8447,N_5997);
or UO_773 (O_773,N_7919,N_8877);
nor UO_774 (O_774,N_9672,N_5844);
nor UO_775 (O_775,N_9965,N_5370);
nor UO_776 (O_776,N_8639,N_6643);
xor UO_777 (O_777,N_9218,N_7278);
nand UO_778 (O_778,N_6831,N_9360);
nand UO_779 (O_779,N_6487,N_5959);
nand UO_780 (O_780,N_8150,N_9400);
nor UO_781 (O_781,N_6944,N_5667);
nor UO_782 (O_782,N_9614,N_8674);
nor UO_783 (O_783,N_9810,N_7647);
nor UO_784 (O_784,N_6842,N_8808);
nor UO_785 (O_785,N_5337,N_9101);
nand UO_786 (O_786,N_9134,N_5239);
nand UO_787 (O_787,N_8126,N_8747);
or UO_788 (O_788,N_7698,N_8513);
or UO_789 (O_789,N_6062,N_6560);
nand UO_790 (O_790,N_5744,N_8089);
and UO_791 (O_791,N_9814,N_8922);
nand UO_792 (O_792,N_8607,N_8537);
nor UO_793 (O_793,N_6714,N_5025);
or UO_794 (O_794,N_5290,N_5150);
and UO_795 (O_795,N_6989,N_7723);
nor UO_796 (O_796,N_9391,N_9146);
and UO_797 (O_797,N_7127,N_9913);
nand UO_798 (O_798,N_9182,N_9055);
nor UO_799 (O_799,N_5151,N_8672);
nor UO_800 (O_800,N_6118,N_6226);
and UO_801 (O_801,N_8668,N_9690);
and UO_802 (O_802,N_9477,N_9519);
and UO_803 (O_803,N_9972,N_8367);
nand UO_804 (O_804,N_5398,N_7322);
nand UO_805 (O_805,N_8918,N_8108);
or UO_806 (O_806,N_9969,N_6115);
and UO_807 (O_807,N_9864,N_8704);
nand UO_808 (O_808,N_7959,N_9929);
and UO_809 (O_809,N_8099,N_7592);
and UO_810 (O_810,N_8857,N_6947);
and UO_811 (O_811,N_5319,N_6346);
nor UO_812 (O_812,N_5184,N_6901);
or UO_813 (O_813,N_5901,N_8983);
and UO_814 (O_814,N_8737,N_8274);
and UO_815 (O_815,N_6166,N_8175);
nor UO_816 (O_816,N_9301,N_8578);
and UO_817 (O_817,N_9071,N_6868);
nor UO_818 (O_818,N_8287,N_8236);
xnor UO_819 (O_819,N_5488,N_9709);
or UO_820 (O_820,N_6645,N_5945);
nor UO_821 (O_821,N_8499,N_7260);
nor UO_822 (O_822,N_7667,N_7703);
nand UO_823 (O_823,N_9089,N_7301);
and UO_824 (O_824,N_8712,N_8094);
and UO_825 (O_825,N_8430,N_9113);
nand UO_826 (O_826,N_7749,N_8122);
nor UO_827 (O_827,N_5838,N_9914);
or UO_828 (O_828,N_8802,N_6072);
nand UO_829 (O_829,N_7433,N_8836);
nand UO_830 (O_830,N_6662,N_9116);
nor UO_831 (O_831,N_8664,N_8151);
nor UO_832 (O_832,N_8871,N_5067);
nor UO_833 (O_833,N_5514,N_9785);
or UO_834 (O_834,N_8187,N_9257);
or UO_835 (O_835,N_5777,N_8008);
and UO_836 (O_836,N_5193,N_5781);
and UO_837 (O_837,N_9474,N_7964);
nor UO_838 (O_838,N_9781,N_7492);
and UO_839 (O_839,N_8032,N_7478);
nand UO_840 (O_840,N_5558,N_7208);
nand UO_841 (O_841,N_9778,N_7920);
nand UO_842 (O_842,N_9623,N_7037);
or UO_843 (O_843,N_8199,N_9490);
and UO_844 (O_844,N_9993,N_9147);
nand UO_845 (O_845,N_7422,N_7420);
or UO_846 (O_846,N_5326,N_8087);
nand UO_847 (O_847,N_6068,N_7984);
nor UO_848 (O_848,N_7276,N_8356);
nand UO_849 (O_849,N_8001,N_9414);
and UO_850 (O_850,N_8307,N_6215);
or UO_851 (O_851,N_8000,N_7379);
and UO_852 (O_852,N_7591,N_5629);
or UO_853 (O_853,N_5988,N_8301);
or UO_854 (O_854,N_5539,N_7375);
and UO_855 (O_855,N_7908,N_5170);
nand UO_856 (O_856,N_7092,N_7323);
nand UO_857 (O_857,N_8544,N_7400);
nand UO_858 (O_858,N_6990,N_6295);
nand UO_859 (O_859,N_8723,N_5582);
or UO_860 (O_860,N_6601,N_6574);
or UO_861 (O_861,N_7168,N_7163);
nor UO_862 (O_862,N_9420,N_8493);
and UO_863 (O_863,N_6593,N_5534);
and UO_864 (O_864,N_6757,N_8349);
xor UO_865 (O_865,N_6063,N_7131);
and UO_866 (O_866,N_9197,N_7438);
nor UO_867 (O_867,N_8527,N_6858);
xnor UO_868 (O_868,N_9976,N_7860);
nand UO_869 (O_869,N_5587,N_8892);
nor UO_870 (O_870,N_7246,N_5208);
nor UO_871 (O_871,N_9758,N_6602);
nand UO_872 (O_872,N_5506,N_7403);
or UO_873 (O_873,N_9846,N_8562);
nor UO_874 (O_874,N_9481,N_5399);
nand UO_875 (O_875,N_7903,N_8494);
nor UO_876 (O_876,N_7222,N_6692);
or UO_877 (O_877,N_6056,N_6292);
nor UO_878 (O_878,N_9553,N_5124);
or UO_879 (O_879,N_9430,N_9479);
nand UO_880 (O_880,N_9204,N_6338);
nor UO_881 (O_881,N_5907,N_6607);
or UO_882 (O_882,N_9659,N_7651);
and UO_883 (O_883,N_5531,N_8152);
or UO_884 (O_884,N_7893,N_5653);
nor UO_885 (O_885,N_7378,N_7354);
nand UO_886 (O_886,N_9245,N_9015);
and UO_887 (O_887,N_7662,N_5668);
nand UO_888 (O_888,N_6417,N_6018);
or UO_889 (O_889,N_9422,N_9314);
and UO_890 (O_890,N_9184,N_7621);
nand UO_891 (O_891,N_9603,N_8518);
or UO_892 (O_892,N_8953,N_8825);
nand UO_893 (O_893,N_5119,N_7380);
or UO_894 (O_894,N_8995,N_9550);
and UO_895 (O_895,N_6035,N_7637);
nand UO_896 (O_896,N_6122,N_9592);
nor UO_897 (O_897,N_9114,N_5998);
nand UO_898 (O_898,N_5389,N_6512);
and UO_899 (O_899,N_5679,N_7177);
or UO_900 (O_900,N_7813,N_9967);
nor UO_901 (O_901,N_8924,N_6017);
nand UO_902 (O_902,N_7315,N_7794);
or UO_903 (O_903,N_7448,N_6184);
and UO_904 (O_904,N_7241,N_7126);
nand UO_905 (O_905,N_9043,N_7346);
or UO_906 (O_906,N_8144,N_7915);
nor UO_907 (O_907,N_5708,N_6854);
and UO_908 (O_908,N_7031,N_6614);
nor UO_909 (O_909,N_8861,N_7209);
nor UO_910 (O_910,N_9405,N_7708);
nor UO_911 (O_911,N_8446,N_5797);
nand UO_912 (O_912,N_7872,N_6708);
nand UO_913 (O_913,N_5361,N_7547);
nand UO_914 (O_914,N_6401,N_9450);
nor UO_915 (O_915,N_9536,N_5305);
or UO_916 (O_916,N_7756,N_7231);
nand UO_917 (O_917,N_8557,N_9087);
and UO_918 (O_918,N_6392,N_5096);
and UO_919 (O_919,N_6915,N_7757);
and UO_920 (O_920,N_9620,N_7851);
and UO_921 (O_921,N_6895,N_8907);
nand UO_922 (O_922,N_7015,N_8893);
nor UO_923 (O_923,N_6790,N_9323);
and UO_924 (O_924,N_5624,N_8186);
or UO_925 (O_925,N_6743,N_9715);
nand UO_926 (O_926,N_7786,N_9990);
and UO_927 (O_927,N_9977,N_6800);
nand UO_928 (O_928,N_9068,N_9458);
or UO_929 (O_929,N_9295,N_7133);
or UO_930 (O_930,N_9255,N_6155);
nand UO_931 (O_931,N_9487,N_6315);
nand UO_932 (O_932,N_8726,N_8363);
nand UO_933 (O_933,N_8883,N_5502);
nand UO_934 (O_934,N_9399,N_8046);
nand UO_935 (O_935,N_5693,N_5257);
nor UO_936 (O_936,N_8967,N_5424);
and UO_937 (O_937,N_9732,N_9524);
nand UO_938 (O_938,N_6886,N_8488);
and UO_939 (O_939,N_5284,N_5670);
nand UO_940 (O_940,N_7535,N_9185);
nand UO_941 (O_941,N_9435,N_6829);
nor UO_942 (O_942,N_6088,N_5074);
or UO_943 (O_943,N_5421,N_6832);
nor UO_944 (O_944,N_5736,N_9356);
and UO_945 (O_945,N_7297,N_7957);
nor UO_946 (O_946,N_5458,N_5200);
and UO_947 (O_947,N_6196,N_5117);
and UO_948 (O_948,N_7808,N_7878);
or UO_949 (O_949,N_9886,N_5499);
and UO_950 (O_950,N_8911,N_6320);
or UO_951 (O_951,N_6686,N_8663);
and UO_952 (O_952,N_7289,N_7817);
and UO_953 (O_953,N_7000,N_9542);
nor UO_954 (O_954,N_5190,N_8680);
nor UO_955 (O_955,N_9783,N_5527);
nor UO_956 (O_956,N_5143,N_6727);
or UO_957 (O_957,N_9271,N_7398);
nor UO_958 (O_958,N_7764,N_9066);
nand UO_959 (O_959,N_6296,N_6635);
or UO_960 (O_960,N_7052,N_9954);
and UO_961 (O_961,N_5450,N_6902);
nand UO_962 (O_962,N_9417,N_5773);
and UO_963 (O_963,N_7901,N_8587);
nand UO_964 (O_964,N_9363,N_9936);
and UO_965 (O_965,N_6534,N_5900);
nor UO_966 (O_966,N_5142,N_7956);
nand UO_967 (O_967,N_7308,N_5155);
or UO_968 (O_968,N_5354,N_9448);
nor UO_969 (O_969,N_9308,N_6523);
and UO_970 (O_970,N_7253,N_7702);
nand UO_971 (O_971,N_9019,N_7148);
and UO_972 (O_972,N_5469,N_7157);
nor UO_973 (O_973,N_9765,N_9552);
nor UO_974 (O_974,N_5951,N_7490);
and UO_975 (O_975,N_5638,N_8210);
or UO_976 (O_976,N_5680,N_7021);
or UO_977 (O_977,N_9402,N_6496);
nand UO_978 (O_978,N_9451,N_7534);
nor UO_979 (O_979,N_6632,N_9888);
nand UO_980 (O_980,N_5898,N_8539);
nand UO_981 (O_981,N_6161,N_8179);
or UO_982 (O_982,N_8748,N_8966);
xnor UO_983 (O_983,N_6146,N_6658);
nand UO_984 (O_984,N_9934,N_7156);
nand UO_985 (O_985,N_6773,N_5656);
nand UO_986 (O_986,N_6347,N_6225);
nor UO_987 (O_987,N_8569,N_7159);
or UO_988 (O_988,N_6573,N_8039);
or UO_989 (O_989,N_8073,N_9981);
or UO_990 (O_990,N_5787,N_8556);
nor UO_991 (O_991,N_8579,N_6130);
nor UO_992 (O_992,N_7436,N_5931);
nand UO_993 (O_993,N_8795,N_9835);
nand UO_994 (O_994,N_7491,N_9243);
nor UO_995 (O_995,N_6084,N_9819);
and UO_996 (O_996,N_7207,N_9375);
nor UO_997 (O_997,N_6569,N_6324);
nor UO_998 (O_998,N_5121,N_9004);
or UO_999 (O_999,N_8540,N_8060);
nand UO_1000 (O_1000,N_7141,N_9036);
nand UO_1001 (O_1001,N_6590,N_8984);
nand UO_1002 (O_1002,N_5053,N_7020);
nand UO_1003 (O_1003,N_7215,N_9554);
nand UO_1004 (O_1004,N_5599,N_6765);
and UO_1005 (O_1005,N_8227,N_5830);
nand UO_1006 (O_1006,N_7633,N_6069);
nand UO_1007 (O_1007,N_8183,N_8952);
nand UO_1008 (O_1008,N_7700,N_6126);
or UO_1009 (O_1009,N_8878,N_7452);
or UO_1010 (O_1010,N_5520,N_8075);
or UO_1011 (O_1011,N_9831,N_9731);
nand UO_1012 (O_1012,N_5000,N_6106);
and UO_1013 (O_1013,N_9767,N_8448);
nor UO_1014 (O_1014,N_8508,N_9551);
nand UO_1015 (O_1015,N_5026,N_7541);
xor UO_1016 (O_1016,N_6699,N_5541);
and UO_1017 (O_1017,N_8767,N_7913);
nand UO_1018 (O_1018,N_5721,N_9418);
or UO_1019 (O_1019,N_8485,N_7888);
or UO_1020 (O_1020,N_5294,N_5388);
nor UO_1021 (O_1021,N_9750,N_5893);
nor UO_1022 (O_1022,N_6647,N_6087);
nor UO_1023 (O_1023,N_5440,N_6370);
nand UO_1024 (O_1024,N_7902,N_8939);
nor UO_1025 (O_1025,N_8418,N_6356);
nand UO_1026 (O_1026,N_8635,N_6258);
and UO_1027 (O_1027,N_7075,N_7466);
or UO_1028 (O_1028,N_7821,N_8725);
nor UO_1029 (O_1029,N_9494,N_5614);
nand UO_1030 (O_1030,N_8638,N_9329);
and UO_1031 (O_1031,N_5264,N_5645);
nor UO_1032 (O_1032,N_6158,N_7938);
nand UO_1033 (O_1033,N_9048,N_9431);
or UO_1034 (O_1034,N_8949,N_9946);
nor UO_1035 (O_1035,N_5229,N_8568);
nor UO_1036 (O_1036,N_7249,N_5479);
and UO_1037 (O_1037,N_5870,N_7165);
xnor UO_1038 (O_1038,N_8512,N_8477);
nor UO_1039 (O_1039,N_5244,N_6326);
nor UO_1040 (O_1040,N_7064,N_5647);
nand UO_1041 (O_1041,N_7430,N_5024);
nand UO_1042 (O_1042,N_5564,N_6826);
and UO_1043 (O_1043,N_5691,N_8558);
and UO_1044 (O_1044,N_9493,N_8956);
nor UO_1045 (O_1045,N_6305,N_6716);
nand UO_1046 (O_1046,N_6202,N_9108);
nor UO_1047 (O_1047,N_7060,N_9530);
nor UO_1048 (O_1048,N_9927,N_8971);
and UO_1049 (O_1049,N_9310,N_5498);
or UO_1050 (O_1050,N_9439,N_8048);
or UO_1051 (O_1051,N_9996,N_5666);
xnor UO_1052 (O_1052,N_6303,N_6532);
and UO_1053 (O_1053,N_5295,N_8451);
nor UO_1054 (O_1054,N_8335,N_5702);
nand UO_1055 (O_1055,N_5181,N_6536);
nor UO_1056 (O_1056,N_6277,N_7612);
or UO_1057 (O_1057,N_9484,N_9662);
nor UO_1058 (O_1058,N_5094,N_5882);
xnor UO_1059 (O_1059,N_8817,N_6547);
or UO_1060 (O_1060,N_6157,N_8500);
or UO_1061 (O_1061,N_6991,N_8404);
or UO_1062 (O_1062,N_8633,N_6756);
or UO_1063 (O_1063,N_8925,N_7224);
nand UO_1064 (O_1064,N_9242,N_8103);
and UO_1065 (O_1065,N_7292,N_7746);
and UO_1066 (O_1066,N_9195,N_8358);
nor UO_1067 (O_1067,N_9568,N_6825);
nand UO_1068 (O_1068,N_7366,N_6807);
nand UO_1069 (O_1069,N_7626,N_7586);
and UO_1070 (O_1070,N_9491,N_7606);
and UO_1071 (O_1071,N_7847,N_5101);
and UO_1072 (O_1072,N_8387,N_9478);
or UO_1073 (O_1073,N_9680,N_7431);
and UO_1074 (O_1074,N_7235,N_8575);
or UO_1075 (O_1075,N_7527,N_9549);
nor UO_1076 (O_1076,N_7601,N_6019);
nor UO_1077 (O_1077,N_9619,N_7871);
nand UO_1078 (O_1078,N_5932,N_9607);
nand UO_1079 (O_1079,N_6471,N_5390);
or UO_1080 (O_1080,N_8450,N_5536);
nor UO_1081 (O_1081,N_6812,N_5173);
xnor UO_1082 (O_1082,N_6132,N_9889);
or UO_1083 (O_1083,N_8458,N_5308);
nor UO_1084 (O_1084,N_5963,N_6885);
or UO_1085 (O_1085,N_8169,N_5508);
and UO_1086 (O_1086,N_8722,N_5640);
or UO_1087 (O_1087,N_5760,N_8876);
or UO_1088 (O_1088,N_9762,N_5613);
and UO_1089 (O_1089,N_6211,N_8394);
nor UO_1090 (O_1090,N_7640,N_8809);
and UO_1091 (O_1091,N_5126,N_6958);
nor UO_1092 (O_1092,N_6091,N_8761);
or UO_1093 (O_1093,N_5625,N_9848);
nor UO_1094 (O_1094,N_9611,N_9713);
nor UO_1095 (O_1095,N_8978,N_6127);
or UO_1096 (O_1096,N_7033,N_5852);
nor UO_1097 (O_1097,N_9677,N_9624);
nor UO_1098 (O_1098,N_9666,N_6374);
and UO_1099 (O_1099,N_6549,N_6220);
and UO_1100 (O_1100,N_9692,N_8535);
and UO_1101 (O_1101,N_6738,N_9841);
nand UO_1102 (O_1102,N_6256,N_8787);
and UO_1103 (O_1103,N_6141,N_7615);
nor UO_1104 (O_1104,N_8240,N_5703);
or UO_1105 (O_1105,N_9813,N_8165);
and UO_1106 (O_1106,N_8511,N_9461);
nor UO_1107 (O_1107,N_8669,N_8397);
nor UO_1108 (O_1108,N_9341,N_9429);
nor UO_1109 (O_1109,N_7958,N_7360);
or UO_1110 (O_1110,N_8174,N_9339);
and UO_1111 (O_1111,N_6769,N_8346);
nand UO_1112 (O_1112,N_5364,N_9096);
nand UO_1113 (O_1113,N_7281,N_8204);
and UO_1114 (O_1114,N_9050,N_6814);
nor UO_1115 (O_1115,N_7394,N_6170);
or UO_1116 (O_1116,N_8415,N_5767);
or UO_1117 (O_1117,N_7937,N_5792);
nand UO_1118 (O_1118,N_7386,N_9595);
and UO_1119 (O_1119,N_6064,N_5804);
nand UO_1120 (O_1120,N_9447,N_9705);
and UO_1121 (O_1121,N_9170,N_8496);
nand UO_1122 (O_1122,N_7514,N_7751);
or UO_1123 (O_1123,N_8902,N_7566);
nand UO_1124 (O_1124,N_8908,N_9138);
xor UO_1125 (O_1125,N_5177,N_7143);
and UO_1126 (O_1126,N_6355,N_7094);
nor UO_1127 (O_1127,N_7976,N_9923);
or UO_1128 (O_1128,N_9289,N_6923);
or UO_1129 (O_1129,N_9786,N_7731);
nand UO_1130 (O_1130,N_5467,N_7368);
and UO_1131 (O_1131,N_5313,N_6596);
or UO_1132 (O_1132,N_6334,N_7149);
and UO_1133 (O_1133,N_6385,N_7524);
or UO_1134 (O_1134,N_5092,N_5524);
nand UO_1135 (O_1135,N_6655,N_9997);
nor UO_1136 (O_1136,N_9324,N_6897);
nor UO_1137 (O_1137,N_5464,N_5234);
nand UO_1138 (O_1138,N_5733,N_9139);
or UO_1139 (O_1139,N_5755,N_8773);
nor UO_1140 (O_1140,N_6123,N_9793);
and UO_1141 (O_1141,N_5135,N_8584);
or UO_1142 (O_1142,N_8194,N_7338);
nor UO_1143 (O_1143,N_6870,N_7634);
nor UO_1144 (O_1144,N_6010,N_9240);
or UO_1145 (O_1145,N_6107,N_9795);
nand UO_1146 (O_1146,N_6621,N_9933);
nand UO_1147 (O_1147,N_7710,N_9869);
and UO_1148 (O_1148,N_8338,N_8234);
or UO_1149 (O_1149,N_6129,N_7372);
and UO_1150 (O_1150,N_9415,N_6758);
nand UO_1151 (O_1151,N_9533,N_7544);
or UO_1152 (O_1152,N_6734,N_8720);
and UO_1153 (O_1153,N_8869,N_8115);
and UO_1154 (O_1154,N_8435,N_9857);
and UO_1155 (O_1155,N_8254,N_7980);
or UO_1156 (O_1156,N_6331,N_9590);
or UO_1157 (O_1157,N_6276,N_6351);
nor UO_1158 (O_1158,N_7408,N_5206);
nor UO_1159 (O_1159,N_8862,N_5937);
and UO_1160 (O_1160,N_6791,N_8472);
nand UO_1161 (O_1161,N_7337,N_7499);
nor UO_1162 (O_1162,N_6389,N_5007);
nand UO_1163 (O_1163,N_9035,N_7050);
or UO_1164 (O_1164,N_8064,N_5598);
nor UO_1165 (O_1165,N_6444,N_9573);
and UO_1166 (O_1166,N_9406,N_6616);
or UO_1167 (O_1167,N_8667,N_5033);
nand UO_1168 (O_1168,N_9612,N_5859);
and UO_1169 (O_1169,N_8022,N_8181);
nor UO_1170 (O_1170,N_9575,N_5857);
nand UO_1171 (O_1171,N_7287,N_5725);
nor UO_1172 (O_1172,N_6817,N_6846);
nor UO_1173 (O_1173,N_9671,N_7951);
nand UO_1174 (O_1174,N_7997,N_9821);
or UO_1175 (O_1175,N_5790,N_6181);
nor UO_1176 (O_1176,N_5616,N_7432);
or UO_1177 (O_1177,N_8388,N_8524);
or UO_1178 (O_1178,N_6052,N_8455);
nor UO_1179 (O_1179,N_9305,N_5763);
nor UO_1180 (O_1180,N_7387,N_8377);
or UO_1181 (O_1181,N_5601,N_5761);
nor UO_1182 (O_1182,N_5652,N_8573);
and UO_1183 (O_1183,N_5904,N_8708);
nor UO_1184 (O_1184,N_6375,N_9829);
and UO_1185 (O_1185,N_6038,N_9588);
or UO_1186 (O_1186,N_6959,N_8804);
nand UO_1187 (O_1187,N_5087,N_5819);
nand UO_1188 (O_1188,N_6461,N_8621);
and UO_1189 (O_1189,N_8369,N_5095);
nand UO_1190 (O_1190,N_7788,N_9499);
nor UO_1191 (O_1191,N_5259,N_5194);
nor UO_1192 (O_1192,N_6725,N_8707);
or UO_1193 (O_1193,N_9220,N_6554);
and UO_1194 (O_1194,N_9733,N_6116);
nand UO_1195 (O_1195,N_8476,N_6516);
and UO_1196 (O_1196,N_9369,N_7577);
or UO_1197 (O_1197,N_8744,N_6105);
nor UO_1198 (O_1198,N_8945,N_8604);
nor UO_1199 (O_1199,N_8785,N_7564);
or UO_1200 (O_1200,N_5176,N_6007);
nand UO_1201 (O_1201,N_8507,N_9523);
nor UO_1202 (O_1202,N_8466,N_7382);
and UO_1203 (O_1203,N_7353,N_9483);
nor UO_1204 (O_1204,N_9851,N_6005);
and UO_1205 (O_1205,N_6613,N_8128);
and UO_1206 (O_1206,N_9467,N_7906);
and UO_1207 (O_1207,N_5303,N_6049);
or UO_1208 (O_1208,N_5336,N_6384);
nand UO_1209 (O_1209,N_6968,N_8880);
and UO_1210 (O_1210,N_5021,N_9651);
or UO_1211 (O_1211,N_8235,N_6024);
or UO_1212 (O_1212,N_6721,N_8070);
nand UO_1213 (O_1213,N_8135,N_8146);
and UO_1214 (O_1214,N_5269,N_5409);
and UO_1215 (O_1215,N_5633,N_5922);
nand UO_1216 (O_1216,N_6435,N_6361);
or UO_1217 (O_1217,N_6559,N_7367);
nand UO_1218 (O_1218,N_5778,N_9576);
nor UO_1219 (O_1219,N_5019,N_7388);
and UO_1220 (O_1220,N_9906,N_9853);
nor UO_1221 (O_1221,N_7877,N_7886);
nor UO_1222 (O_1222,N_8798,N_8913);
or UO_1223 (O_1223,N_5433,N_9259);
nor UO_1224 (O_1224,N_9287,N_7392);
nor UO_1225 (O_1225,N_5066,N_7760);
and UO_1226 (O_1226,N_5427,N_7947);
nand UO_1227 (O_1227,N_9518,N_9582);
nor UO_1228 (O_1228,N_6014,N_5350);
nand UO_1229 (O_1229,N_9351,N_5298);
or UO_1230 (O_1230,N_5588,N_5057);
and UO_1231 (O_1231,N_7184,N_9663);
xor UO_1232 (O_1232,N_7179,N_8546);
nand UO_1233 (O_1233,N_8080,N_7793);
nand UO_1234 (O_1234,N_9636,N_6381);
nor UO_1235 (O_1235,N_8682,N_5232);
nor UO_1236 (O_1236,N_8602,N_7081);
and UO_1237 (O_1237,N_9412,N_5732);
nand UO_1238 (O_1238,N_6508,N_5381);
or UO_1239 (O_1239,N_8519,N_5353);
or UO_1240 (O_1240,N_6147,N_7932);
nand UO_1241 (O_1241,N_7371,N_9500);
nand UO_1242 (O_1242,N_5400,N_5521);
or UO_1243 (O_1243,N_8976,N_7483);
and UO_1244 (O_1244,N_8014,N_5443);
or UO_1245 (O_1245,N_7280,N_6942);
nor UO_1246 (O_1246,N_5414,N_6656);
nor UO_1247 (O_1247,N_8988,N_9995);
and UO_1248 (O_1248,N_6463,N_8786);
or UO_1249 (O_1249,N_5402,N_8119);
and UO_1250 (O_1250,N_5251,N_8162);
nor UO_1251 (O_1251,N_5927,N_5628);
nor UO_1252 (O_1252,N_8462,N_6151);
and UO_1253 (O_1253,N_6329,N_5268);
or UO_1254 (O_1254,N_7147,N_5675);
and UO_1255 (O_1255,N_9932,N_6358);
or UO_1256 (O_1256,N_7682,N_6945);
or UO_1257 (O_1257,N_6724,N_9394);
nand UO_1258 (O_1258,N_5751,N_9567);
or UO_1259 (O_1259,N_6477,N_7370);
and UO_1260 (O_1260,N_8774,N_8752);
nor UO_1261 (O_1261,N_8489,N_7931);
nor UO_1262 (O_1262,N_6066,N_7803);
nor UO_1263 (O_1263,N_8964,N_9083);
or UO_1264 (O_1264,N_8082,N_9002);
and UO_1265 (O_1265,N_8459,N_7227);
nand UO_1266 (O_1266,N_6319,N_6548);
and UO_1267 (O_1267,N_6585,N_5970);
nor UO_1268 (O_1268,N_5002,N_9053);
nand UO_1269 (O_1269,N_7789,N_5862);
nand UO_1270 (O_1270,N_7639,N_6189);
nand UO_1271 (O_1271,N_5323,N_9759);
nor UO_1272 (O_1272,N_8781,N_7205);
or UO_1273 (O_1273,N_6120,N_6907);
or UO_1274 (O_1274,N_5231,N_7783);
and UO_1275 (O_1275,N_8504,N_8262);
nand UO_1276 (O_1276,N_5509,N_7355);
nor UO_1277 (O_1277,N_9740,N_9504);
nor UO_1278 (O_1278,N_5256,N_5064);
or UO_1279 (O_1279,N_9093,N_7600);
and UO_1280 (O_1280,N_5144,N_5358);
nor UO_1281 (O_1281,N_8221,N_6993);
nor UO_1282 (O_1282,N_7164,N_9078);
nand UO_1283 (O_1283,N_8849,N_5699);
nand UO_1284 (O_1284,N_8855,N_5872);
or UO_1285 (O_1285,N_7739,N_5617);
and UO_1286 (O_1286,N_8758,N_7933);
and UO_1287 (O_1287,N_5646,N_7797);
nor UO_1288 (O_1288,N_6134,N_7928);
and UO_1289 (O_1289,N_6121,N_9313);
or UO_1290 (O_1290,N_6227,N_9629);
and UO_1291 (O_1291,N_6104,N_8931);
nand UO_1292 (O_1292,N_6171,N_7532);
or UO_1293 (O_1293,N_9982,N_7273);
nand UO_1294 (O_1294,N_9547,N_7521);
or UO_1295 (O_1295,N_6633,N_9897);
nor UO_1296 (O_1296,N_6604,N_6111);
or UO_1297 (O_1297,N_8605,N_8246);
nor UO_1298 (O_1298,N_9007,N_6609);
and UO_1299 (O_1299,N_6422,N_7411);
and UO_1300 (O_1300,N_5320,N_9849);
and UO_1301 (O_1301,N_9540,N_7828);
nand UO_1302 (O_1302,N_5630,N_8206);
and UO_1303 (O_1303,N_9309,N_7414);
nand UO_1304 (O_1304,N_7294,N_9855);
nor UO_1305 (O_1305,N_8832,N_9284);
or UO_1306 (O_1306,N_8671,N_8033);
and UO_1307 (O_1307,N_6462,N_7210);
xnor UO_1308 (O_1308,N_7012,N_8293);
or UO_1309 (O_1309,N_6458,N_6637);
nor UO_1310 (O_1310,N_6622,N_7334);
nand UO_1311 (O_1311,N_9123,N_8421);
nand UO_1312 (O_1312,N_7862,N_6238);
xor UO_1313 (O_1313,N_8121,N_9460);
nor UO_1314 (O_1314,N_6236,N_9084);
or UO_1315 (O_1315,N_8930,N_8754);
and UO_1316 (O_1316,N_9515,N_8125);
and UO_1317 (O_1317,N_7399,N_9669);
nor UO_1318 (O_1318,N_9894,N_8357);
or UO_1319 (O_1319,N_8117,N_9772);
nand UO_1320 (O_1320,N_7638,N_6691);
nand UO_1321 (O_1321,N_7284,N_7508);
or UO_1322 (O_1322,N_8426,N_8685);
nand UO_1323 (O_1323,N_5304,N_7858);
or UO_1324 (O_1324,N_6363,N_6232);
nand UO_1325 (O_1325,N_5724,N_6852);
and UO_1326 (O_1326,N_8844,N_5420);
and UO_1327 (O_1327,N_6094,N_7270);
nand UO_1328 (O_1328,N_6709,N_5526);
and UO_1329 (O_1329,N_9025,N_6615);
or UO_1330 (O_1330,N_6805,N_7391);
and UO_1331 (O_1331,N_6733,N_8443);
nand UO_1332 (O_1332,N_9956,N_8874);
nor UO_1333 (O_1333,N_7175,N_7946);
nand UO_1334 (O_1334,N_7194,N_5444);
nor UO_1335 (O_1335,N_6815,N_6679);
nor UO_1336 (O_1336,N_9456,N_9719);
nand UO_1337 (O_1337,N_6624,N_8644);
and UO_1338 (O_1338,N_6978,N_7006);
nand UO_1339 (O_1339,N_6407,N_9591);
nor UO_1340 (O_1340,N_5586,N_7975);
nand UO_1341 (O_1341,N_8846,N_7088);
and UO_1342 (O_1342,N_8982,N_7087);
and UO_1343 (O_1343,N_8205,N_5253);
nand UO_1344 (O_1344,N_9269,N_9325);
or UO_1345 (O_1345,N_8497,N_7385);
nor UO_1346 (O_1346,N_6575,N_5070);
or UO_1347 (O_1347,N_9653,N_6543);
nor UO_1348 (O_1348,N_8969,N_6954);
nor UO_1349 (O_1349,N_9966,N_8870);
xnor UO_1350 (O_1350,N_5482,N_9791);
and UO_1351 (O_1351,N_7424,N_6274);
nor UO_1352 (O_1352,N_8351,N_7003);
nor UO_1353 (O_1353,N_5296,N_6454);
nand UO_1354 (O_1354,N_6310,N_9939);
nor UO_1355 (O_1355,N_6627,N_6086);
or UO_1356 (O_1356,N_5322,N_8990);
or UO_1357 (O_1357,N_6388,N_8444);
and UO_1358 (O_1358,N_8093,N_8738);
nor UO_1359 (O_1359,N_9251,N_6982);
or UO_1360 (O_1360,N_5192,N_5281);
xor UO_1361 (O_1361,N_8646,N_5947);
nor UO_1362 (O_1362,N_6112,N_7685);
nand UO_1363 (O_1363,N_7672,N_9948);
nor UO_1364 (O_1364,N_7001,N_8347);
nand UO_1365 (O_1365,N_6787,N_7520);
or UO_1366 (O_1366,N_7151,N_8614);
nand UO_1367 (O_1367,N_6618,N_9097);
and UO_1368 (O_1368,N_8185,N_5867);
or UO_1369 (O_1369,N_7842,N_9618);
nand UO_1370 (O_1370,N_8947,N_5560);
nand UO_1371 (O_1371,N_8914,N_7505);
or UO_1372 (O_1372,N_5106,N_5981);
nor UO_1373 (O_1373,N_8879,N_8606);
or UO_1374 (O_1374,N_5043,N_7468);
nand UO_1375 (O_1375,N_6600,N_6293);
and UO_1376 (O_1376,N_7010,N_6774);
or UO_1377 (O_1377,N_7038,N_6173);
nand UO_1378 (O_1378,N_5452,N_7244);
or UO_1379 (O_1379,N_7198,N_8330);
nand UO_1380 (O_1380,N_5250,N_5285);
nor UO_1381 (O_1381,N_7668,N_5487);
nand UO_1382 (O_1382,N_7780,N_5345);
or UO_1383 (O_1383,N_8251,N_8096);
or UO_1384 (O_1384,N_5602,N_5563);
and UO_1385 (O_1385,N_8909,N_7298);
nand UO_1386 (O_1386,N_5957,N_8465);
nor UO_1387 (O_1387,N_6838,N_7067);
and UO_1388 (O_1388,N_9153,N_5876);
nand UO_1389 (O_1389,N_6136,N_8027);
and UO_1390 (O_1390,N_8088,N_8563);
nor UO_1391 (O_1391,N_7487,N_9716);
or UO_1392 (O_1392,N_5579,N_7663);
and UO_1393 (O_1393,N_8715,N_5347);
nand UO_1394 (O_1394,N_6020,N_8171);
and UO_1395 (O_1395,N_9610,N_7999);
nand UO_1396 (O_1396,N_6976,N_8896);
nand UO_1397 (O_1397,N_9172,N_7080);
nor UO_1398 (O_1398,N_5116,N_7416);
nor UO_1399 (O_1399,N_5914,N_7361);
nand UO_1400 (O_1400,N_9290,N_6612);
or UO_1401 (O_1401,N_5113,N_6586);
or UO_1402 (O_1402,N_5047,N_5622);
or UO_1403 (O_1403,N_5954,N_7119);
nand UO_1404 (O_1404,N_9160,N_8208);
and UO_1405 (O_1405,N_9975,N_9544);
nand UO_1406 (O_1406,N_8673,N_5739);
nand UO_1407 (O_1407,N_7025,N_5407);
nor UO_1408 (O_1408,N_6969,N_5926);
and UO_1409 (O_1409,N_6266,N_9800);
and UO_1410 (O_1410,N_6257,N_6550);
nor UO_1411 (O_1411,N_7083,N_7022);
nand UO_1412 (O_1412,N_7669,N_6806);
nand UO_1413 (O_1413,N_6382,N_6016);
nand UO_1414 (O_1414,N_9779,N_8142);
or UO_1415 (O_1415,N_8314,N_5317);
and UO_1416 (O_1416,N_8716,N_5476);
nand UO_1417 (O_1417,N_6930,N_5310);
and UO_1418 (O_1418,N_8190,N_8700);
and UO_1419 (O_1419,N_7190,N_7855);
and UO_1420 (O_1420,N_9207,N_7102);
nor UO_1421 (O_1421,N_8081,N_7412);
nand UO_1422 (O_1422,N_7116,N_7264);
xnor UO_1423 (O_1423,N_7464,N_8298);
nand UO_1424 (O_1424,N_5805,N_8991);
nand UO_1425 (O_1425,N_6689,N_9655);
and UO_1426 (O_1426,N_8975,N_8051);
nor UO_1427 (O_1427,N_6952,N_9398);
and UO_1428 (O_1428,N_6223,N_8770);
or UO_1429 (O_1429,N_5877,N_6060);
nand UO_1430 (O_1430,N_8906,N_6768);
or UO_1431 (O_1431,N_7004,N_6479);
nand UO_1432 (O_1432,N_6410,N_7885);
nor UO_1433 (O_1433,N_5546,N_8821);
nand UO_1434 (O_1434,N_7673,N_8034);
nand UO_1435 (O_1435,N_8164,N_5288);
or UO_1436 (O_1436,N_5329,N_5962);
and UO_1437 (O_1437,N_5753,N_8055);
nor UO_1438 (O_1438,N_5131,N_5316);
and UO_1439 (O_1439,N_8661,N_6440);
nand UO_1440 (O_1440,N_9013,N_9885);
nor UO_1441 (O_1441,N_7771,N_5812);
or UO_1442 (O_1442,N_7889,N_9292);
nor UO_1443 (O_1443,N_9221,N_9960);
xor UO_1444 (O_1444,N_7107,N_6697);
nand UO_1445 (O_1445,N_5248,N_8180);
nor UO_1446 (O_1446,N_7900,N_7917);
nand UO_1447 (O_1447,N_9694,N_9441);
nor UO_1448 (O_1448,N_9919,N_7104);
nand UO_1449 (O_1449,N_7977,N_7652);
nor UO_1450 (O_1450,N_9606,N_9642);
and UO_1451 (O_1451,N_5948,N_8554);
nand UO_1452 (O_1452,N_5277,N_5140);
and UO_1453 (O_1453,N_5127,N_9585);
nor UO_1454 (O_1454,N_5110,N_8506);
nand UO_1455 (O_1455,N_5454,N_5118);
and UO_1456 (O_1456,N_6728,N_6816);
and UO_1457 (O_1457,N_5609,N_7515);
and UO_1458 (O_1458,N_7381,N_5318);
nor UO_1459 (O_1459,N_9061,N_7356);
nor UO_1460 (O_1460,N_5887,N_8741);
and UO_1461 (O_1461,N_9167,N_7580);
nor UO_1462 (O_1462,N_6628,N_7869);
or UO_1463 (O_1463,N_5892,N_9373);
nand UO_1464 (O_1464,N_9942,N_8686);
and UO_1465 (O_1465,N_9376,N_9935);
or UO_1466 (O_1466,N_9031,N_7265);
nor UO_1467 (O_1467,N_8184,N_7271);
nor UO_1468 (O_1468,N_9707,N_6224);
nand UO_1469 (O_1469,N_8457,N_8545);
or UO_1470 (O_1470,N_8895,N_6135);
xnor UO_1471 (O_1471,N_5145,N_5385);
or UO_1472 (O_1472,N_7720,N_8534);
and UO_1473 (O_1473,N_7303,N_5660);
or UO_1474 (O_1474,N_6000,N_5297);
nand UO_1475 (O_1475,N_8018,N_5529);
or UO_1476 (O_1476,N_8505,N_7790);
nand UO_1477 (O_1477,N_8768,N_8201);
nor UO_1478 (O_1478,N_6079,N_8735);
or UO_1479 (O_1479,N_9092,N_8962);
nand UO_1480 (O_1480,N_5813,N_6015);
or UO_1481 (O_1481,N_9722,N_5315);
nand UO_1482 (O_1482,N_5153,N_5576);
nor UO_1483 (O_1483,N_5346,N_6918);
or UO_1484 (O_1484,N_5405,N_7509);
xor UO_1485 (O_1485,N_5552,N_5911);
or UO_1486 (O_1486,N_6651,N_5023);
nor UO_1487 (O_1487,N_9353,N_6780);
nand UO_1488 (O_1488,N_8736,N_6891);
and UO_1489 (O_1489,N_8996,N_9102);
and UO_1490 (O_1490,N_7373,N_5861);
and UO_1491 (O_1491,N_8202,N_9615);
nor UO_1492 (O_1492,N_6456,N_7809);
or UO_1493 (O_1493,N_8713,N_6486);
xnor UO_1494 (O_1494,N_7513,N_7706);
or UO_1495 (O_1495,N_9739,N_9176);
nand UO_1496 (O_1496,N_9496,N_7849);
or UO_1497 (O_1497,N_9973,N_5956);
and UO_1498 (O_1498,N_7654,N_6045);
and UO_1499 (O_1499,N_6450,N_5495);
endmodule