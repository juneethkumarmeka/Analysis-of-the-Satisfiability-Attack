module basic_1500_15000_2000_75_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_366,In_190);
or U1 (N_1,In_663,In_1371);
nand U2 (N_2,In_170,In_443);
nor U3 (N_3,In_886,In_744);
or U4 (N_4,In_371,In_924);
nand U5 (N_5,In_1463,In_119);
xor U6 (N_6,In_1257,In_1474);
or U7 (N_7,In_1281,In_932);
nor U8 (N_8,In_125,In_234);
nand U9 (N_9,In_894,In_1422);
and U10 (N_10,In_318,In_1129);
and U11 (N_11,In_281,In_931);
and U12 (N_12,In_474,In_923);
nor U13 (N_13,In_565,In_973);
nor U14 (N_14,In_479,In_835);
nand U15 (N_15,In_809,In_1189);
or U16 (N_16,In_159,In_1019);
nand U17 (N_17,In_647,In_437);
or U18 (N_18,In_1133,In_562);
xor U19 (N_19,In_899,In_669);
xor U20 (N_20,In_867,In_107);
nand U21 (N_21,In_1253,In_950);
nor U22 (N_22,In_72,In_1159);
or U23 (N_23,In_1218,In_1476);
or U24 (N_24,In_675,In_510);
nor U25 (N_25,In_703,In_676);
xor U26 (N_26,In_1302,In_941);
or U27 (N_27,In_1293,In_713);
or U28 (N_28,In_247,In_65);
nor U29 (N_29,In_458,In_633);
nand U30 (N_30,In_477,In_674);
nor U31 (N_31,In_512,In_909);
nor U32 (N_32,In_87,In_200);
nor U33 (N_33,In_1263,In_433);
and U34 (N_34,In_354,In_1195);
nor U35 (N_35,In_786,In_1052);
xnor U36 (N_36,In_819,In_729);
nand U37 (N_37,In_784,In_333);
xnor U38 (N_38,In_517,In_895);
or U39 (N_39,In_834,In_148);
and U40 (N_40,In_901,In_1336);
nand U41 (N_41,In_1036,In_1341);
nor U42 (N_42,In_974,In_1110);
nor U43 (N_43,In_1228,In_1241);
nand U44 (N_44,In_276,In_731);
or U45 (N_45,In_967,In_79);
nand U46 (N_46,In_1149,In_1437);
and U47 (N_47,In_765,In_601);
and U48 (N_48,In_1456,In_163);
or U49 (N_49,In_722,In_736);
or U50 (N_50,In_586,In_797);
nand U51 (N_51,In_617,In_456);
and U52 (N_52,In_441,In_825);
or U53 (N_53,In_1069,In_488);
nand U54 (N_54,In_235,In_1374);
nand U55 (N_55,In_139,In_432);
or U56 (N_56,In_501,In_1358);
nand U57 (N_57,In_944,In_1327);
nand U58 (N_58,In_1247,In_10);
nor U59 (N_59,In_261,In_680);
or U60 (N_60,In_589,In_648);
xnor U61 (N_61,In_363,In_1215);
nor U62 (N_62,In_677,In_1322);
and U63 (N_63,In_316,In_1481);
nand U64 (N_64,In_1396,In_298);
nand U65 (N_65,In_120,In_31);
nand U66 (N_66,In_26,In_440);
nor U67 (N_67,In_382,In_7);
and U68 (N_68,In_618,In_632);
nand U69 (N_69,In_1389,In_1136);
or U70 (N_70,In_449,In_915);
and U71 (N_71,In_1059,In_1352);
nor U72 (N_72,In_523,In_112);
nand U73 (N_73,In_704,In_1060);
nand U74 (N_74,In_1089,In_447);
nand U75 (N_75,In_138,In_1032);
or U76 (N_76,In_612,In_860);
nor U77 (N_77,In_1350,In_564);
and U78 (N_78,In_1066,In_368);
nor U79 (N_79,In_885,In_1109);
or U80 (N_80,In_845,In_104);
or U81 (N_81,In_375,In_1193);
and U82 (N_82,In_1353,In_1154);
nand U83 (N_83,In_34,In_192);
nor U84 (N_84,In_219,In_233);
nor U85 (N_85,In_1412,In_408);
nand U86 (N_86,In_659,In_228);
nand U87 (N_87,In_1268,In_478);
xor U88 (N_88,In_1120,In_728);
or U89 (N_89,In_715,In_1273);
nand U90 (N_90,In_146,In_579);
nor U91 (N_91,In_239,In_407);
and U92 (N_92,In_779,In_196);
nand U93 (N_93,In_852,In_166);
and U94 (N_94,In_550,In_455);
nand U95 (N_95,In_288,In_790);
and U96 (N_96,In_900,In_1030);
and U97 (N_97,In_1178,In_1102);
and U98 (N_98,In_1416,In_19);
and U99 (N_99,In_1187,In_1419);
or U100 (N_100,In_623,In_39);
and U101 (N_101,In_370,In_1013);
nand U102 (N_102,In_1483,In_379);
nor U103 (N_103,In_716,In_1104);
and U104 (N_104,In_723,In_544);
and U105 (N_105,In_324,In_329);
nor U106 (N_106,In_1184,In_727);
nor U107 (N_107,In_806,In_1289);
or U108 (N_108,In_547,In_1306);
and U109 (N_109,In_184,In_266);
or U110 (N_110,In_1359,In_301);
nor U111 (N_111,In_693,In_429);
and U112 (N_112,In_740,In_1124);
and U113 (N_113,In_921,In_1497);
nand U114 (N_114,In_1064,In_1079);
and U115 (N_115,In_210,In_29);
and U116 (N_116,In_188,In_545);
nor U117 (N_117,In_587,In_975);
and U118 (N_118,In_661,In_1487);
or U119 (N_119,In_1294,In_1356);
and U120 (N_120,In_250,In_347);
or U121 (N_121,In_1369,In_448);
xor U122 (N_122,In_1223,In_1261);
xor U123 (N_123,In_1084,In_1333);
nand U124 (N_124,In_452,In_927);
nand U125 (N_125,In_1311,In_1291);
nand U126 (N_126,In_492,In_853);
and U127 (N_127,In_113,In_62);
nand U128 (N_128,In_1464,In_516);
nor U129 (N_129,In_115,In_257);
or U130 (N_130,In_995,In_70);
or U131 (N_131,In_751,In_757);
nand U132 (N_132,In_572,In_52);
and U133 (N_133,In_286,In_1330);
and U134 (N_134,In_1192,In_1450);
and U135 (N_135,In_529,In_454);
and U136 (N_136,In_936,In_665);
or U137 (N_137,In_773,In_1017);
or U138 (N_138,In_891,In_588);
and U139 (N_139,In_285,In_1251);
and U140 (N_140,In_1403,In_1424);
xnor U141 (N_141,In_1298,In_1145);
nand U142 (N_142,In_307,In_692);
nand U143 (N_143,In_220,In_842);
and U144 (N_144,In_493,In_871);
nor U145 (N_145,In_582,In_342);
xor U146 (N_146,In_1329,In_1367);
or U147 (N_147,In_502,In_896);
or U148 (N_148,In_350,In_1351);
nor U149 (N_149,In_642,In_424);
nand U150 (N_150,In_850,In_1346);
nor U151 (N_151,In_1132,In_1307);
nand U152 (N_152,In_935,In_914);
nand U153 (N_153,In_338,In_848);
nand U154 (N_154,In_1174,In_1284);
nor U155 (N_155,In_947,In_241);
nor U156 (N_156,In_1026,In_992);
nor U157 (N_157,In_212,In_1146);
and U158 (N_158,In_1209,In_951);
or U159 (N_159,In_621,In_1397);
nor U160 (N_160,In_1452,In_348);
and U161 (N_161,In_627,In_280);
nor U162 (N_162,In_8,In_778);
and U163 (N_163,In_925,In_262);
or U164 (N_164,In_1206,In_1020);
nor U165 (N_165,In_697,In_360);
and U166 (N_166,In_748,In_426);
and U167 (N_167,In_635,In_327);
nor U168 (N_168,In_801,In_1155);
and U169 (N_169,In_737,In_785);
nand U170 (N_170,In_741,In_533);
and U171 (N_171,In_1141,In_1015);
or U172 (N_172,In_1049,In_222);
nand U173 (N_173,In_1318,In_268);
nor U174 (N_174,In_671,In_710);
nor U175 (N_175,In_733,In_607);
and U176 (N_176,In_643,In_884);
and U177 (N_177,In_1343,In_933);
nand U178 (N_178,In_263,In_1055);
nand U179 (N_179,In_962,In_171);
nor U180 (N_180,In_1144,In_386);
nor U181 (N_181,In_98,In_609);
nand U182 (N_182,In_1401,In_450);
nand U183 (N_183,In_1494,In_172);
nand U184 (N_184,In_1267,In_614);
nor U185 (N_185,In_144,In_417);
and U186 (N_186,In_994,In_574);
nand U187 (N_187,In_684,In_1349);
and U188 (N_188,In_1075,In_345);
nand U189 (N_189,In_1377,In_1116);
and U190 (N_190,In_521,In_175);
nand U191 (N_191,In_875,In_705);
or U192 (N_192,In_1085,In_151);
nor U193 (N_193,In_513,In_961);
and U194 (N_194,In_945,In_1037);
xor U195 (N_195,In_794,In_1387);
and U196 (N_196,In_1199,In_176);
nor U197 (N_197,In_1469,In_993);
or U198 (N_198,In_1114,In_396);
xor U199 (N_199,In_1150,In_832);
nand U200 (N_200,In_583,In_165);
xnor U201 (N_201,In_224,In_349);
nand U202 (N_202,In_137,In_1347);
and U203 (N_203,In_1345,In_63);
and U204 (N_204,In_490,In_1001);
or U205 (N_205,In_917,In_260);
nand U206 (N_206,In_53,In_73);
nand U207 (N_207,In_334,N_59);
nor U208 (N_208,N_117,In_1400);
nor U209 (N_209,N_133,In_484);
or U210 (N_210,In_831,In_485);
nand U211 (N_211,In_546,In_71);
or U212 (N_212,In_289,In_1477);
nor U213 (N_213,In_804,In_240);
nor U214 (N_214,In_1460,In_272);
or U215 (N_215,N_11,In_1137);
nor U216 (N_216,In_497,In_1453);
nor U217 (N_217,N_189,In_77);
or U218 (N_218,In_1384,N_28);
nor U219 (N_219,In_907,In_712);
or U220 (N_220,In_463,In_1443);
nor U221 (N_221,In_655,In_1073);
nor U222 (N_222,In_827,In_134);
nor U223 (N_223,In_37,In_543);
nand U224 (N_224,In_1444,In_1210);
or U225 (N_225,In_796,In_101);
nand U226 (N_226,In_873,In_561);
nor U227 (N_227,In_1185,In_1092);
and U228 (N_228,In_387,In_956);
or U229 (N_229,In_1088,In_21);
nand U230 (N_230,In_1007,In_1131);
and U231 (N_231,In_640,In_602);
xor U232 (N_232,N_125,In_649);
or U233 (N_233,In_1264,In_1279);
nor U234 (N_234,In_194,In_326);
and U235 (N_235,In_179,In_570);
nor U236 (N_236,N_174,In_960);
nand U237 (N_237,N_169,In_472);
nand U238 (N_238,In_168,In_195);
nand U239 (N_239,In_341,N_22);
nor U240 (N_240,In_149,In_1182);
and U241 (N_241,N_53,N_74);
nor U242 (N_242,In_594,In_381);
or U243 (N_243,In_721,In_390);
nand U244 (N_244,In_1004,In_1214);
and U245 (N_245,In_913,In_469);
and U246 (N_246,N_27,In_1287);
xnor U247 (N_247,In_82,In_1062);
and U248 (N_248,N_149,N_67);
nand U249 (N_249,In_1372,In_1246);
or U250 (N_250,In_279,N_194);
nor U251 (N_251,In_1386,In_598);
xor U252 (N_252,In_1418,In_187);
and U253 (N_253,N_36,In_1034);
nor U254 (N_254,In_1233,N_134);
nor U255 (N_255,In_916,In_1083);
nor U256 (N_256,In_66,In_500);
nand U257 (N_257,In_1362,In_208);
nor U258 (N_258,In_799,In_527);
xnor U259 (N_259,In_776,In_76);
and U260 (N_260,In_116,In_628);
nor U261 (N_261,In_434,N_138);
nor U262 (N_262,In_59,In_937);
xnor U263 (N_263,N_47,In_1411);
or U264 (N_264,In_296,N_55);
nand U265 (N_265,In_352,In_613);
or U266 (N_266,In_664,In_616);
nor U267 (N_267,In_47,N_165);
nor U268 (N_268,In_23,In_1440);
nand U269 (N_269,In_103,In_768);
nor U270 (N_270,In_435,In_560);
and U271 (N_271,In_274,In_1225);
xor U272 (N_272,N_162,In_245);
nor U273 (N_273,In_511,N_105);
nand U274 (N_274,In_254,In_393);
nand U275 (N_275,In_963,In_634);
and U276 (N_276,In_812,In_1172);
nand U277 (N_277,In_238,In_889);
or U278 (N_278,In_1243,In_946);
nand U279 (N_279,In_385,In_494);
or U280 (N_280,In_998,N_135);
or U281 (N_281,In_1312,In_491);
xor U282 (N_282,In_177,In_650);
or U283 (N_283,In_725,In_1006);
xnor U284 (N_284,In_780,N_51);
or U285 (N_285,In_402,In_344);
nor U286 (N_286,In_556,In_1258);
or U287 (N_287,In_506,In_590);
nand U288 (N_288,In_864,N_72);
nand U289 (N_289,In_255,N_15);
nand U290 (N_290,In_844,In_207);
or U291 (N_291,In_652,In_1191);
and U292 (N_292,In_611,In_299);
and U293 (N_293,In_708,In_226);
nor U294 (N_294,In_1454,In_753);
nand U295 (N_295,In_1489,In_557);
and U296 (N_296,In_531,In_1157);
nor U297 (N_297,In_1045,In_278);
and U298 (N_298,In_707,N_0);
nand U299 (N_299,In_1467,In_1388);
and U300 (N_300,In_833,N_127);
and U301 (N_301,In_1262,In_840);
xor U302 (N_302,In_1099,In_1236);
or U303 (N_303,In_1479,N_92);
or U304 (N_304,In_930,In_256);
or U305 (N_305,In_199,In_678);
or U306 (N_306,In_297,In_320);
nor U307 (N_307,In_660,In_567);
and U308 (N_308,In_686,In_185);
or U309 (N_309,N_183,In_987);
and U310 (N_310,In_391,In_215);
nand U311 (N_311,In_969,In_696);
nand U312 (N_312,In_604,In_1410);
nand U313 (N_313,In_1103,In_308);
or U314 (N_314,N_140,In_1320);
nor U315 (N_315,In_752,In_656);
nand U316 (N_316,In_481,N_101);
nor U317 (N_317,In_857,In_911);
xor U318 (N_318,In_668,In_92);
nor U319 (N_319,N_75,In_174);
or U320 (N_320,In_1301,In_624);
and U321 (N_321,In_1082,In_411);
and U322 (N_322,In_1138,In_15);
nor U323 (N_323,In_27,In_672);
nor U324 (N_324,In_117,In_405);
and U325 (N_325,In_340,In_1275);
xor U326 (N_326,In_595,In_1065);
xor U327 (N_327,In_20,N_193);
nand U328 (N_328,In_1090,In_1237);
nand U329 (N_329,In_223,In_1196);
nor U330 (N_330,In_421,In_1376);
nand U331 (N_331,In_549,In_745);
or U332 (N_332,In_783,N_52);
xnor U333 (N_333,In_1119,In_1162);
nand U334 (N_334,N_102,In_558);
xor U335 (N_335,In_1285,In_84);
or U336 (N_336,In_1429,In_1143);
or U337 (N_337,N_197,In_483);
nand U338 (N_338,In_1283,In_398);
and U339 (N_339,N_77,In_577);
nand U340 (N_340,In_1470,In_28);
or U341 (N_341,In_1295,In_133);
nand U342 (N_342,In_1466,N_2);
nand U343 (N_343,In_1039,In_1057);
xnor U344 (N_344,In_136,In_46);
and U345 (N_345,In_305,In_221);
nor U346 (N_346,In_1364,In_807);
and U347 (N_347,In_395,In_859);
and U348 (N_348,In_217,In_1380);
nor U349 (N_349,In_36,In_18);
and U350 (N_350,In_232,In_1449);
nor U351 (N_351,In_302,In_1153);
or U352 (N_352,In_5,In_1435);
nor U353 (N_353,In_294,N_49);
nand U354 (N_354,In_979,In_1002);
nor U355 (N_355,N_89,N_91);
nor U356 (N_356,In_108,In_213);
or U357 (N_357,In_1363,In_803);
nand U358 (N_358,In_1357,In_1127);
nand U359 (N_359,In_265,In_620);
or U360 (N_360,N_50,In_69);
and U361 (N_361,In_400,In_1304);
or U362 (N_362,N_199,In_126);
and U363 (N_363,In_571,In_1296);
or U364 (N_364,In_1220,In_482);
or U365 (N_365,In_1239,In_45);
or U366 (N_366,N_42,In_563);
and U367 (N_367,In_35,N_64);
or U368 (N_368,N_124,In_1230);
or U369 (N_369,In_95,In_958);
nor U370 (N_370,In_473,In_61);
or U371 (N_371,In_282,N_48);
nor U372 (N_372,In_1278,N_98);
xnor U373 (N_373,In_795,In_1331);
or U374 (N_374,In_682,In_1023);
nor U375 (N_375,In_1061,N_122);
or U376 (N_376,In_141,In_1365);
or U377 (N_377,In_1378,In_1234);
and U378 (N_378,In_81,N_34);
and U379 (N_379,In_952,In_756);
nor U380 (N_380,In_626,In_1095);
xnor U381 (N_381,In_1360,In_374);
nor U382 (N_382,N_30,In_1171);
nor U383 (N_383,In_145,In_462);
nand U384 (N_384,N_70,In_685);
nor U385 (N_385,In_193,In_1126);
and U386 (N_386,In_1167,In_681);
and U387 (N_387,In_1370,In_619);
nor U388 (N_388,In_1417,In_1334);
nand U389 (N_389,N_198,N_9);
or U390 (N_390,In_657,In_903);
nand U391 (N_391,In_415,In_759);
nand U392 (N_392,In_989,In_769);
xor U393 (N_393,In_243,N_188);
nor U394 (N_394,In_540,N_35);
nand U395 (N_395,N_14,N_7);
nor U396 (N_396,N_29,N_45);
or U397 (N_397,In_33,In_158);
xnor U398 (N_398,In_526,In_1130);
xnor U399 (N_399,In_4,N_137);
and U400 (N_400,N_159,In_1314);
nor U401 (N_401,N_399,In_377);
nor U402 (N_402,In_427,In_180);
xnor U403 (N_403,In_743,In_425);
xor U404 (N_404,In_629,In_991);
nand U405 (N_405,In_597,In_418);
or U406 (N_406,N_314,In_823);
xnor U407 (N_407,In_1063,N_362);
and U408 (N_408,In_225,In_1499);
nor U409 (N_409,N_300,In_1248);
xor U410 (N_410,In_881,N_249);
nand U411 (N_411,In_1299,N_171);
or U412 (N_412,N_252,In_110);
and U413 (N_413,In_460,N_132);
nor U414 (N_414,In_496,In_181);
nor U415 (N_415,In_314,In_416);
nand U416 (N_416,In_855,In_1393);
xnor U417 (N_417,N_379,In_1379);
nand U418 (N_418,In_1112,In_800);
or U419 (N_419,In_155,In_74);
nand U420 (N_420,In_1269,In_514);
nand U421 (N_421,In_1458,In_537);
nand U422 (N_422,In_1074,In_406);
nand U423 (N_423,In_1337,In_1425);
and U424 (N_424,In_948,In_972);
or U425 (N_425,In_1255,N_378);
or U426 (N_426,N_222,In_706);
nor U427 (N_427,In_1271,N_93);
or U428 (N_428,N_347,In_161);
and U429 (N_429,In_1414,In_264);
xnor U430 (N_430,In_878,In_695);
and U431 (N_431,N_373,In_267);
and U432 (N_432,N_106,N_353);
nor U433 (N_433,In_1406,In_548);
and U434 (N_434,In_43,N_395);
and U435 (N_435,N_380,In_788);
or U436 (N_436,N_358,In_1219);
xnor U437 (N_437,In_1402,In_464);
xor U438 (N_438,In_167,In_1047);
or U439 (N_439,N_278,N_218);
nor U440 (N_440,N_361,In_40);
nor U441 (N_441,N_153,N_230);
nor U442 (N_442,In_1491,In_205);
and U443 (N_443,In_880,In_1028);
and U444 (N_444,In_820,N_295);
xnor U445 (N_445,In_68,N_343);
and U446 (N_446,In_1398,In_843);
nor U447 (N_447,In_592,In_690);
nand U448 (N_448,In_1290,In_717);
and U449 (N_449,In_1113,N_186);
or U450 (N_450,In_1040,In_249);
nand U451 (N_451,In_926,N_282);
and U452 (N_452,In_755,In_1);
nor U453 (N_453,N_385,In_1160);
or U454 (N_454,In_346,In_1348);
nor U455 (N_455,N_33,N_116);
xor U456 (N_456,In_593,In_96);
or U457 (N_457,In_310,In_413);
xnor U458 (N_458,In_498,In_1022);
nor U459 (N_459,In_837,In_1170);
or U460 (N_460,In_331,N_184);
nand U461 (N_461,N_291,N_224);
nor U462 (N_462,In_442,In_1031);
and U463 (N_463,N_391,In_1197);
nand U464 (N_464,In_1316,In_1381);
nor U465 (N_465,In_1216,In_9);
xor U466 (N_466,In_897,In_439);
and U467 (N_467,In_836,N_119);
and U468 (N_468,In_153,In_761);
xnor U469 (N_469,N_150,In_1313);
nand U470 (N_470,N_76,N_350);
and U471 (N_471,In_879,N_173);
nand U472 (N_472,N_368,N_397);
or U473 (N_473,In_216,In_738);
nand U474 (N_474,In_688,In_1208);
and U475 (N_475,In_358,N_60);
or U476 (N_476,N_235,In_1176);
nand U477 (N_477,N_147,In_1300);
nand U478 (N_478,In_525,N_144);
nor U479 (N_479,N_264,N_136);
nand U480 (N_480,N_242,In_929);
or U481 (N_481,In_714,In_1122);
or U482 (N_482,In_575,In_55);
nand U483 (N_483,In_323,N_236);
or U484 (N_484,In_1142,In_476);
and U485 (N_485,N_247,In_569);
and U486 (N_486,In_332,In_1207);
or U487 (N_487,N_352,N_152);
nor U488 (N_488,N_366,In_97);
xnor U489 (N_489,In_730,N_387);
and U490 (N_490,In_465,In_541);
and U491 (N_491,N_294,In_130);
or U492 (N_492,N_317,In_898);
and U493 (N_493,In_57,In_1277);
nor U494 (N_494,In_639,In_698);
and U495 (N_495,In_814,In_1498);
nand U496 (N_496,In_143,In_910);
and U497 (N_497,N_219,In_636);
or U498 (N_498,In_581,In_351);
and U499 (N_499,In_760,N_348);
or U500 (N_500,N_258,In_466);
xor U501 (N_501,In_1106,In_1152);
xnor U502 (N_502,In_404,In_1226);
nor U503 (N_503,In_388,N_297);
nor U504 (N_504,N_69,In_24);
nor U505 (N_505,N_143,In_1096);
nand U506 (N_506,In_830,In_309);
nand U507 (N_507,In_14,In_41);
and U508 (N_508,In_976,In_1280);
nor U509 (N_509,In_965,In_293);
or U510 (N_510,N_337,In_520);
and U511 (N_511,In_644,In_882);
nand U512 (N_512,In_78,N_316);
nor U513 (N_513,In_129,In_1173);
nand U514 (N_514,In_1077,In_410);
nor U515 (N_515,In_983,In_1319);
nor U516 (N_516,In_1430,In_1025);
and U517 (N_517,N_240,In_1121);
nor U518 (N_518,N_179,N_231);
and U519 (N_519,In_461,In_12);
xor U520 (N_520,In_777,In_446);
nand U521 (N_521,In_851,In_128);
nand U522 (N_522,N_142,N_312);
and U523 (N_523,In_1010,In_58);
or U524 (N_524,N_205,In_793);
nand U525 (N_525,In_539,In_670);
and U526 (N_526,In_487,In_522);
and U527 (N_527,In_808,N_326);
and U528 (N_528,N_296,N_96);
nand U529 (N_529,In_1442,In_912);
xor U530 (N_530,In_821,N_283);
nor U531 (N_531,N_24,In_306);
or U532 (N_532,N_123,In_423);
or U533 (N_533,In_438,In_489);
and U534 (N_534,N_71,N_232);
nor U535 (N_535,N_213,N_129);
nand U536 (N_536,N_202,In_874);
nand U537 (N_537,N_248,In_1164);
and U538 (N_538,In_709,N_141);
nor U539 (N_539,In_152,In_1148);
or U540 (N_540,In_1405,In_378);
and U541 (N_541,In_362,In_1231);
nor U542 (N_542,N_372,N_86);
and U543 (N_543,N_177,In_480);
nand U544 (N_544,N_8,In_519);
nor U545 (N_545,In_876,In_980);
or U546 (N_546,In_1086,In_1324);
or U547 (N_547,N_255,In_771);
nor U548 (N_548,In_99,In_1471);
and U549 (N_549,N_374,In_142);
nand U550 (N_550,In_813,N_304);
or U551 (N_551,In_1448,N_307);
or U552 (N_552,In_1433,N_246);
xor U553 (N_553,In_905,In_1305);
nand U554 (N_554,N_241,In_230);
xor U555 (N_555,N_207,N_371);
nand U556 (N_556,In_353,N_327);
and U557 (N_557,N_356,N_229);
and U558 (N_558,N_275,In_44);
nand U559 (N_559,In_573,In_719);
nor U560 (N_560,In_1035,N_280);
or U561 (N_561,In_1097,In_638);
nand U562 (N_562,In_258,In_524);
xnor U563 (N_563,In_237,In_1181);
nand U564 (N_564,In_1492,N_388);
and U565 (N_565,In_1229,N_345);
nor U566 (N_566,In_1203,In_412);
nor U567 (N_567,In_336,In_1420);
or U568 (N_568,In_870,In_666);
nor U569 (N_569,N_244,N_341);
or U570 (N_570,In_1366,In_1413);
nand U571 (N_571,In_868,N_256);
nor U572 (N_572,In_1332,In_856);
and U573 (N_573,In_1067,In_1081);
xor U574 (N_574,N_313,N_225);
nand U575 (N_575,N_292,In_3);
or U576 (N_576,N_80,In_1436);
xor U577 (N_577,In_1188,In_1391);
nor U578 (N_578,In_826,N_267);
nand U579 (N_579,In_1321,In_1242);
and U580 (N_580,In_475,N_145);
nand U581 (N_581,In_1441,In_106);
and U582 (N_582,In_1240,In_1468);
nand U583 (N_583,N_262,N_40);
nand U584 (N_584,N_299,N_243);
or U585 (N_585,In_162,In_1408);
or U586 (N_586,N_208,N_156);
and U587 (N_587,In_253,In_1180);
xor U588 (N_588,In_532,In_922);
or U589 (N_589,N_112,In_1115);
nand U590 (N_590,In_1472,In_954);
or U591 (N_591,N_344,In_1179);
and U592 (N_592,N_331,In_1339);
and U593 (N_593,In_691,In_1016);
or U594 (N_594,In_858,In_1204);
nor U595 (N_595,In_603,In_322);
or U596 (N_596,In_1043,N_118);
nand U597 (N_597,In_1438,In_1222);
xnor U598 (N_598,In_887,N_18);
xnor U599 (N_599,In_343,In_1070);
nor U600 (N_600,In_1147,In_367);
nand U601 (N_601,N_212,N_32);
xnor U602 (N_602,N_130,N_166);
nand U603 (N_603,In_542,N_178);
or U604 (N_604,N_411,In_735);
and U605 (N_605,In_982,In_271);
and U606 (N_606,N_417,In_747);
or U607 (N_607,N_220,In_1375);
xnor U608 (N_608,N_285,In_1014);
and U609 (N_609,N_100,In_2);
xor U610 (N_610,N_492,In_86);
nor U611 (N_611,In_1111,N_447);
nor U612 (N_612,N_302,In_1166);
and U613 (N_613,N_384,N_108);
xor U614 (N_614,N_265,In_315);
or U615 (N_615,In_1100,N_554);
nand U616 (N_616,N_154,In_1286);
and U617 (N_617,N_479,N_386);
or U618 (N_618,In_509,In_1183);
or U619 (N_619,In_732,In_270);
nor U620 (N_620,N_115,N_454);
and U621 (N_621,In_1093,In_403);
nand U622 (N_622,In_746,N_558);
and U623 (N_623,N_393,N_227);
nand U624 (N_624,N_531,N_505);
nand U625 (N_625,N_415,In_1427);
nor U626 (N_626,In_508,N_563);
nand U627 (N_627,In_50,N_585);
nor U628 (N_628,N_214,In_1309);
nor U629 (N_629,In_1457,In_1217);
or U630 (N_630,In_920,In_1266);
nand U631 (N_631,In_67,In_399);
nand U632 (N_632,N_587,In_1276);
xor U633 (N_633,In_109,N_588);
nor U634 (N_634,In_100,In_147);
nor U635 (N_635,In_1428,In_54);
nand U636 (N_636,N_37,N_467);
or U637 (N_637,In_311,N_310);
nand U638 (N_638,N_576,In_164);
nor U639 (N_639,N_572,In_1000);
nor U640 (N_640,N_309,In_553);
and U641 (N_641,N_84,In_118);
xnor U642 (N_642,In_419,In_1009);
nor U643 (N_643,N_477,N_209);
xor U644 (N_644,In_445,In_596);
xnor U645 (N_645,N_210,In_1482);
or U646 (N_646,N_419,In_1335);
nor U647 (N_647,In_1445,N_553);
nand U648 (N_648,In_1087,N_223);
nand U649 (N_649,N_38,In_1399);
or U650 (N_650,In_940,N_161);
and U651 (N_651,In_699,In_290);
or U652 (N_652,In_397,In_124);
and U653 (N_653,In_1169,In_1395);
and U654 (N_654,In_1165,N_99);
or U655 (N_655,In_990,In_1018);
nor U656 (N_656,N_437,N_190);
or U657 (N_657,In_1190,In_22);
nand U658 (N_658,In_824,N_578);
nor U659 (N_659,N_109,In_453);
or U660 (N_660,In_883,In_470);
and U661 (N_661,In_1323,N_557);
or U662 (N_662,In_892,N_293);
or U663 (N_663,N_590,N_435);
and U664 (N_664,N_425,In_1259);
nor U665 (N_665,N_398,N_511);
nor U666 (N_666,In_227,N_521);
and U667 (N_667,In_662,N_465);
and U668 (N_668,N_216,In_495);
or U669 (N_669,In_409,N_128);
and U670 (N_670,N_104,N_286);
nor U671 (N_671,In_838,In_1446);
and U672 (N_672,N_476,N_570);
nand U673 (N_673,N_168,N_176);
nor U674 (N_674,In_13,In_157);
and U675 (N_675,N_259,In_1317);
or U676 (N_676,N_20,N_540);
or U677 (N_677,N_460,N_598);
nor U678 (N_678,In_888,N_439);
nand U679 (N_679,In_300,In_383);
nand U680 (N_680,N_273,N_541);
nand U681 (N_681,N_167,In_615);
and U682 (N_682,In_32,In_938);
and U683 (N_683,N_305,N_381);
or U684 (N_684,N_396,N_192);
nand U685 (N_685,In_658,In_414);
nor U686 (N_686,N_83,In_1213);
or U687 (N_687,In_105,In_1053);
and U688 (N_688,N_306,In_1272);
and U689 (N_689,In_16,In_275);
or U690 (N_690,N_349,In_865);
nor U691 (N_691,In_1244,In_325);
and U692 (N_692,N_320,In_312);
and U693 (N_693,In_111,N_333);
nand U694 (N_694,In_599,N_446);
or U695 (N_695,N_418,N_329);
or U696 (N_696,In_64,In_90);
or U697 (N_697,N_448,N_403);
and U698 (N_698,N_595,N_560);
nand U699 (N_699,N_360,N_409);
nor U700 (N_700,N_462,N_405);
or U701 (N_701,In_1252,In_284);
nand U702 (N_702,N_475,N_114);
nor U703 (N_703,In_248,In_361);
nand U704 (N_704,In_203,N_66);
nor U705 (N_705,In_292,N_526);
and U706 (N_706,N_269,In_1068);
xnor U707 (N_707,In_372,N_440);
nor U708 (N_708,In_1308,In_631);
or U709 (N_709,N_311,In_1260);
or U710 (N_710,In_1158,In_1373);
nand U711 (N_711,N_336,N_443);
or U712 (N_712,N_82,In_645);
or U713 (N_713,In_1139,In_1194);
and U714 (N_714,N_324,In_1238);
and U715 (N_715,In_750,In_467);
or U716 (N_716,In_1005,N_516);
and U717 (N_717,In_273,N_537);
nand U718 (N_718,In_1496,N_318);
or U719 (N_719,N_288,In_1056);
or U720 (N_720,N_148,N_568);
xnor U721 (N_721,In_173,In_1368);
nor U722 (N_722,In_1415,In_772);
and U723 (N_723,N_376,N_470);
nor U724 (N_724,In_943,N_23);
or U725 (N_725,In_1198,In_904);
nand U726 (N_726,N_284,In_637);
or U727 (N_727,In_373,N_487);
and U728 (N_728,N_26,N_195);
nor U729 (N_729,In_622,N_481);
xnor U730 (N_730,N_517,In_121);
nand U731 (N_731,In_919,In_1042);
nand U732 (N_732,N_200,In_357);
and U733 (N_733,N_529,In_38);
or U734 (N_734,N_346,In_93);
nand U735 (N_735,In_60,N_315);
nor U736 (N_736,In_849,In_444);
or U737 (N_737,In_767,In_1392);
or U738 (N_738,N_95,N_85);
nor U739 (N_739,N_453,In_140);
xor U740 (N_740,N_416,N_518);
xnor U741 (N_741,N_498,In_646);
or U742 (N_742,N_555,In_1488);
nor U743 (N_743,N_533,In_123);
or U744 (N_744,In_1485,N_25);
and U745 (N_745,In_11,N_163);
or U746 (N_746,In_828,N_4);
or U747 (N_747,In_1024,N_463);
nand U748 (N_748,N_527,In_214);
xnor U749 (N_749,N_103,N_61);
and U750 (N_750,In_1094,N_484);
nor U751 (N_751,In_503,N_420);
nor U752 (N_752,In_1407,In_1012);
nand U753 (N_753,In_328,In_811);
nand U754 (N_754,N_522,In_1227);
and U755 (N_755,In_726,In_1338);
and U756 (N_756,In_754,In_667);
or U757 (N_757,In_287,In_186);
nor U758 (N_758,In_206,N_363);
or U759 (N_759,In_242,In_1249);
nor U760 (N_760,In_829,N_340);
nor U761 (N_761,In_981,N_211);
and U762 (N_762,In_1212,In_641);
or U763 (N_763,In_359,In_770);
nor U764 (N_764,In_1340,In_782);
nor U765 (N_765,In_966,In_955);
and U766 (N_766,In_1303,In_88);
or U767 (N_767,In_1270,In_798);
nor U768 (N_768,In_80,N_274);
nand U769 (N_769,In_997,N_31);
xor U770 (N_770,N_504,N_277);
or U771 (N_771,N_196,In_75);
and U772 (N_772,In_499,N_523);
xor U773 (N_773,N_441,In_1409);
nor U774 (N_774,In_555,In_700);
xnor U775 (N_775,N_412,N_458);
nor U776 (N_776,N_430,N_543);
and U777 (N_777,In_1151,In_1354);
nand U778 (N_778,In_939,N_263);
nand U779 (N_779,N_328,In_1265);
nor U780 (N_780,In_160,In_365);
or U781 (N_781,In_854,N_469);
nor U782 (N_782,In_85,N_421);
nand U783 (N_783,In_1098,In_1385);
and U784 (N_784,N_63,N_355);
nand U785 (N_785,In_89,N_164);
and U786 (N_786,N_586,N_383);
nand U787 (N_787,In_1245,N_459);
nand U788 (N_788,In_580,N_429);
nor U789 (N_789,N_488,In_384);
or U790 (N_790,In_1484,N_468);
nand U791 (N_791,N_581,In_1254);
nor U792 (N_792,N_206,In_459);
nor U793 (N_793,N_251,N_234);
nor U794 (N_794,In_1342,In_1041);
and U795 (N_795,In_673,In_568);
nor U796 (N_796,In_1051,In_1490);
nor U797 (N_797,In_246,In_608);
or U798 (N_798,In_718,In_724);
nor U799 (N_799,N_266,N_509);
nor U800 (N_800,In_1462,In_317);
nor U801 (N_801,N_564,In_1486);
nand U802 (N_802,N_611,In_775);
or U803 (N_803,In_304,In_749);
nor U804 (N_804,N_643,N_375);
nor U805 (N_805,N_754,In_277);
nand U806 (N_806,In_1058,N_616);
or U807 (N_807,N_745,N_428);
xor U808 (N_808,In_295,N_39);
nor U809 (N_809,N_749,In_178);
nand U810 (N_810,N_290,In_1326);
nor U811 (N_811,N_609,N_499);
xor U812 (N_812,N_624,In_1423);
nor U813 (N_813,N_94,In_83);
nor U814 (N_814,N_591,N_741);
nand U815 (N_815,In_376,N_753);
or U816 (N_816,In_1076,In_1315);
and U817 (N_817,N_694,In_1175);
nand U818 (N_818,N_682,N_545);
nor U819 (N_819,N_260,N_473);
and U820 (N_820,In_25,In_505);
or U821 (N_821,In_585,N_617);
or U822 (N_822,In_986,In_49);
nand U823 (N_823,In_1232,In_1382);
or U824 (N_824,N_464,N_548);
nor U825 (N_825,N_646,In_131);
and U826 (N_826,N_270,In_1201);
nand U827 (N_827,N_621,N_257);
nor U828 (N_828,In_701,In_1021);
xnor U829 (N_829,N_704,N_569);
nand U830 (N_830,In_1071,N_452);
and U831 (N_831,In_451,In_428);
or U832 (N_832,N_746,N_737);
or U833 (N_833,N_444,N_325);
and U834 (N_834,N_698,N_81);
nand U835 (N_835,In_739,N_744);
nand U836 (N_836,In_1459,N_427);
or U837 (N_837,In_1495,N_279);
nor U838 (N_838,N_684,N_674);
nand U839 (N_839,N_319,In_436);
and U840 (N_840,N_774,N_732);
or U841 (N_841,N_619,N_413);
nand U842 (N_842,In_1383,N_608);
nor U843 (N_843,N_677,N_514);
and U844 (N_844,N_606,N_351);
and U845 (N_845,N_17,N_759);
xor U846 (N_846,N_673,N_323);
nor U847 (N_847,N_618,In_1493);
and U848 (N_848,N_664,In_816);
nor U849 (N_849,In_303,N_65);
nand U850 (N_850,In_530,N_457);
xnor U851 (N_851,In_1355,N_491);
nand U852 (N_852,N_490,In_1426);
xor U853 (N_853,N_612,N_638);
or U854 (N_854,N_728,N_705);
nand U855 (N_855,N_726,N_559);
or U856 (N_856,N_637,N_767);
nor U857 (N_857,N_394,In_576);
and U858 (N_858,N_215,N_710);
and U859 (N_859,In_209,In_1038);
xnor U860 (N_860,N_644,In_252);
xnor U861 (N_861,N_524,N_721);
nand U862 (N_862,N_734,N_632);
xor U863 (N_863,In_791,In_1118);
nand U864 (N_864,N_406,In_339);
and U865 (N_865,N_512,N_658);
and U866 (N_866,N_238,In_389);
nor U867 (N_867,N_339,N_500);
xor U868 (N_868,N_436,N_596);
nor U869 (N_869,N_422,In_1390);
nand U870 (N_870,In_1256,In_999);
nor U871 (N_871,N_107,In_610);
and U872 (N_872,N_589,N_782);
nand U873 (N_873,N_730,N_679);
or U874 (N_874,N_332,N_696);
nand U875 (N_875,N_656,In_846);
nand U876 (N_876,N_780,In_1361);
nor U877 (N_877,N_731,N_335);
nand U878 (N_878,N_445,N_46);
nand U879 (N_879,N_433,N_87);
nand U880 (N_880,N_503,N_594);
or U881 (N_881,In_1288,In_251);
or U882 (N_882,N_68,In_394);
and U883 (N_883,N_659,N_401);
nor U884 (N_884,N_359,In_762);
or U885 (N_885,In_1478,N_478);
or U886 (N_886,N_78,N_640);
xor U887 (N_887,In_319,N_57);
and U888 (N_888,In_957,In_1200);
nor U889 (N_889,N_424,N_623);
nor U890 (N_890,N_582,In_1054);
or U891 (N_891,N_146,In_122);
nand U892 (N_892,N_709,In_802);
or U893 (N_893,In_313,N_699);
nand U894 (N_894,N_90,N_797);
and U895 (N_895,N_508,N_700);
nand U896 (N_896,In_1224,In_877);
nand U897 (N_897,N_180,N_170);
or U898 (N_898,N_472,In_114);
nor U899 (N_899,In_988,N_56);
and U900 (N_900,In_507,N_276);
nor U901 (N_901,N_707,In_1177);
or U902 (N_902,In_1044,N_725);
xnor U903 (N_903,N_228,In_486);
and U904 (N_904,In_51,In_1205);
nor U905 (N_905,In_863,N_486);
and U906 (N_906,N_766,N_613);
or U907 (N_907,In_908,In_17);
xor U908 (N_908,In_1186,N_793);
nor U909 (N_909,N_466,N_442);
or U910 (N_910,N_271,In_1101);
nand U911 (N_911,In_847,N_407);
nor U912 (N_912,N_691,N_650);
or U913 (N_913,N_706,In_758);
xor U914 (N_914,N_301,In_970);
and U915 (N_915,In_763,In_890);
or U916 (N_916,N_685,N_423);
nand U917 (N_917,In_1250,In_1328);
and U918 (N_918,N_321,N_338);
nor U919 (N_919,N_182,N_233);
or U920 (N_920,N_97,N_226);
or U921 (N_921,In_1046,N_729);
and U922 (N_922,In_559,N_583);
or U923 (N_923,In_1421,N_739);
nand U924 (N_924,N_719,N_438);
or U925 (N_925,In_605,N_298);
nand U926 (N_926,N_636,In_1008);
nor U927 (N_927,In_1048,In_1344);
nor U928 (N_928,N_538,N_546);
or U929 (N_929,N_599,N_456);
nand U930 (N_930,N_711,N_703);
nand U931 (N_931,In_1211,In_431);
or U932 (N_932,In_789,N_642);
xor U933 (N_933,N_547,In_606);
nor U934 (N_934,N_649,In_1107);
nor U935 (N_935,N_772,N_788);
xnor U936 (N_936,In_720,N_482);
or U937 (N_937,N_392,In_337);
and U938 (N_938,In_1091,N_54);
or U939 (N_939,In_422,In_1140);
nor U940 (N_940,In_764,In_653);
and U941 (N_941,N_308,N_354);
or U942 (N_942,N_217,N_552);
nand U943 (N_943,N_785,In_1394);
or U944 (N_944,N_687,In_1135);
or U945 (N_945,In_1168,In_654);
nand U946 (N_946,In_985,N_743);
and U947 (N_947,In_689,N_760);
or U948 (N_948,N_480,In_906);
and U949 (N_949,N_510,N_798);
and U950 (N_950,In_380,N_634);
or U951 (N_951,In_996,N_614);
xor U952 (N_952,In_964,In_1123);
nand U953 (N_953,N_735,N_501);
or U954 (N_954,N_534,In_694);
nand U955 (N_955,In_330,N_628);
and U956 (N_956,In_1163,In_551);
xor U957 (N_957,In_202,N_334);
and U958 (N_958,N_775,In_528);
or U959 (N_959,N_752,N_414);
nor U960 (N_960,N_626,N_689);
nor U961 (N_961,N_544,N_672);
nor U962 (N_962,N_203,N_779);
or U963 (N_963,N_404,In_711);
and U964 (N_964,N_474,In_91);
and U965 (N_965,In_918,In_1455);
or U966 (N_966,In_56,In_1432);
and U967 (N_967,In_150,N_790);
and U968 (N_968,N_693,In_869);
nand U969 (N_969,N_432,In_335);
nor U970 (N_970,In_420,N_641);
xor U971 (N_971,N_761,In_515);
xnor U972 (N_972,N_377,N_556);
nand U973 (N_973,In_211,N_660);
nand U974 (N_974,N_16,In_401);
or U975 (N_975,In_841,N_254);
and U976 (N_976,In_742,In_1475);
or U977 (N_977,N_712,In_1310);
nor U978 (N_978,N_5,In_1292);
and U979 (N_979,N_520,In_584);
nor U980 (N_980,N_157,N_126);
and U981 (N_981,N_740,N_191);
and U982 (N_982,N_663,In_6);
or U983 (N_983,N_722,N_528);
nor U984 (N_984,N_670,N_539);
nor U985 (N_985,In_355,In_244);
nor U986 (N_986,In_1325,In_902);
nor U987 (N_987,In_1134,N_365);
nand U988 (N_988,N_580,In_1480);
nor U989 (N_989,In_683,In_552);
nand U990 (N_990,In_127,N_724);
nand U991 (N_991,N_43,N_683);
and U992 (N_992,N_653,In_862);
nand U993 (N_993,N_357,N_577);
or U994 (N_994,In_554,In_154);
nor U995 (N_995,N_513,N_151);
or U996 (N_996,N_622,N_605);
nand U997 (N_997,In_1128,N_221);
xnor U998 (N_998,In_1282,N_625);
and U999 (N_999,N_647,In_1297);
or U1000 (N_1000,N_885,N_155);
nand U1001 (N_1001,N_822,In_534);
and U1002 (N_1002,N_542,N_869);
nand U1003 (N_1003,In_928,In_356);
or U1004 (N_1004,N_967,N_73);
xor U1005 (N_1005,N_751,N_874);
nor U1006 (N_1006,In_504,In_591);
nand U1007 (N_1007,N_801,N_808);
nor U1008 (N_1008,In_1050,In_817);
or U1009 (N_1009,N_855,N_938);
or U1010 (N_1010,In_1202,In_978);
nand U1011 (N_1011,N_714,N_342);
nand U1012 (N_1012,N_662,N_844);
nor U1013 (N_1013,N_973,N_550);
nor U1014 (N_1014,N_812,N_930);
and U1015 (N_1015,N_676,N_768);
xnor U1016 (N_1016,N_668,In_132);
nand U1017 (N_1017,N_41,N_811);
nand U1018 (N_1018,N_821,N_971);
and U1019 (N_1019,N_830,N_449);
xnor U1020 (N_1020,N_678,N_573);
nand U1021 (N_1021,In_182,In_231);
nor U1022 (N_1022,In_169,N_44);
nand U1023 (N_1023,N_849,N_532);
and U1024 (N_1024,In_984,N_681);
and U1025 (N_1025,In_1003,N_450);
and U1026 (N_1026,In_578,N_692);
nor U1027 (N_1027,N_976,In_197);
and U1028 (N_1028,N_245,N_680);
nand U1029 (N_1029,N_940,N_771);
and U1030 (N_1030,N_922,N_551);
nand U1031 (N_1031,N_695,N_965);
and U1032 (N_1032,N_856,In_1434);
nor U1033 (N_1033,In_839,In_94);
or U1034 (N_1034,N_952,N_382);
and U1035 (N_1035,N_455,N_817);
nor U1036 (N_1036,N_877,N_838);
nor U1037 (N_1037,N_268,N_633);
nand U1038 (N_1038,In_1105,N_895);
and U1039 (N_1039,N_651,N_842);
or U1040 (N_1040,N_597,N_181);
nand U1041 (N_1041,In_1033,N_717);
xor U1042 (N_1042,N_854,In_1461);
nand U1043 (N_1043,N_963,In_959);
or U1044 (N_1044,In_600,N_783);
nor U1045 (N_1045,N_648,In_535);
or U1046 (N_1046,In_392,N_639);
or U1047 (N_1047,N_859,N_370);
nor U1048 (N_1048,N_507,N_756);
nand U1049 (N_1049,N_851,In_1029);
nand U1050 (N_1050,N_897,In_651);
nor U1051 (N_1051,N_287,N_887);
and U1052 (N_1052,N_955,In_183);
nand U1053 (N_1053,N_201,N_836);
nor U1054 (N_1054,N_718,In_822);
and U1055 (N_1055,N_862,In_30);
and U1056 (N_1056,In_866,N_289);
and U1057 (N_1057,In_1117,N_992);
or U1058 (N_1058,N_571,N_924);
nor U1059 (N_1059,N_742,N_402);
and U1060 (N_1060,N_786,In_1011);
nand U1061 (N_1061,N_878,In_430);
nand U1062 (N_1062,N_937,In_1072);
nor U1063 (N_1063,N_565,In_291);
and U1064 (N_1064,N_912,N_765);
nand U1065 (N_1065,N_6,N_939);
or U1066 (N_1066,In_1125,N_600);
and U1067 (N_1067,N_871,N_904);
or U1068 (N_1068,N_431,N_876);
and U1069 (N_1069,N_655,In_518);
nor U1070 (N_1070,N_863,N_928);
nor U1071 (N_1071,N_956,N_873);
nor U1072 (N_1072,N_400,In_815);
and U1073 (N_1073,N_485,N_715);
or U1074 (N_1074,N_716,N_21);
xor U1075 (N_1075,N_120,N_629);
or U1076 (N_1076,In_1161,N_850);
and U1077 (N_1077,N_567,N_755);
and U1078 (N_1078,In_566,N_894);
and U1079 (N_1079,N_889,In_625);
nand U1080 (N_1080,N_870,N_110);
and U1081 (N_1081,N_839,N_915);
nand U1082 (N_1082,N_575,N_872);
nand U1083 (N_1083,In_1439,In_949);
nand U1084 (N_1084,N_875,N_175);
nand U1085 (N_1085,N_172,N_635);
nand U1086 (N_1086,N_997,N_579);
and U1087 (N_1087,N_10,N_910);
nor U1088 (N_1088,N_493,N_802);
nor U1089 (N_1089,N_891,N_330);
nand U1090 (N_1090,In_229,N_281);
or U1091 (N_1091,N_367,In_48);
or U1092 (N_1092,In_189,In_204);
nor U1093 (N_1093,N_261,N_620);
or U1094 (N_1094,N_820,N_561);
nand U1095 (N_1095,N_495,N_426);
nor U1096 (N_1096,N_630,N_847);
or U1097 (N_1097,N_602,N_671);
or U1098 (N_1098,N_893,In_1078);
nand U1099 (N_1099,In_805,N_815);
or U1100 (N_1100,N_389,N_549);
nor U1101 (N_1101,N_451,N_914);
and U1102 (N_1102,N_949,N_747);
or U1103 (N_1103,N_654,N_951);
or U1104 (N_1104,N_974,In_1431);
nor U1105 (N_1105,N_62,In_953);
nand U1106 (N_1106,N_733,In_766);
and U1107 (N_1107,N_322,N_701);
or U1108 (N_1108,N_805,N_111);
nor U1109 (N_1109,N_113,N_994);
or U1110 (N_1110,N_926,N_607);
xor U1111 (N_1111,N_784,N_879);
or U1112 (N_1112,In_198,N_979);
and U1113 (N_1113,N_702,N_947);
and U1114 (N_1114,N_860,N_795);
nand U1115 (N_1115,N_978,In_1465);
and U1116 (N_1116,N_601,N_935);
and U1117 (N_1117,N_763,N_943);
nand U1118 (N_1118,N_932,In_321);
xor U1119 (N_1119,N_483,In_968);
and U1120 (N_1120,N_945,N_713);
nand U1121 (N_1121,N_789,N_840);
nand U1122 (N_1122,N_390,N_250);
and U1123 (N_1123,N_886,N_806);
xor U1124 (N_1124,N_661,N_903);
nor U1125 (N_1125,N_834,N_237);
xor U1126 (N_1126,N_669,In_1274);
and U1127 (N_1127,N_434,N_566);
xnor U1128 (N_1128,N_920,N_816);
nand U1129 (N_1129,In_942,N_899);
or U1130 (N_1130,N_948,N_461);
xor U1131 (N_1131,N_962,N_884);
and U1132 (N_1132,N_835,In_269);
or U1133 (N_1133,N_921,N_160);
nor U1134 (N_1134,N_204,N_905);
or U1135 (N_1135,In_283,N_954);
or U1136 (N_1136,N_890,N_907);
xor U1137 (N_1137,In_42,N_666);
and U1138 (N_1138,N_986,N_708);
nand U1139 (N_1139,In_536,N_927);
nor U1140 (N_1140,N_158,In_457);
or U1141 (N_1141,N_645,N_867);
nor U1142 (N_1142,N_883,N_946);
nor U1143 (N_1143,N_911,N_750);
and U1144 (N_1144,N_970,N_828);
nor U1145 (N_1145,In_538,N_530);
nor U1146 (N_1146,N_762,In_218);
nor U1147 (N_1147,N_690,N_3);
nor U1148 (N_1148,N_832,N_813);
nand U1149 (N_1149,N_996,In_0);
nand U1150 (N_1150,N_975,N_757);
nor U1151 (N_1151,N_989,N_984);
nor U1152 (N_1152,N_665,N_868);
xnor U1153 (N_1153,N_991,N_824);
nor U1154 (N_1154,N_791,In_1080);
nand U1155 (N_1155,N_1,N_736);
nor U1156 (N_1156,N_615,N_852);
and U1157 (N_1157,N_776,N_506);
nand U1158 (N_1158,In_1108,N_593);
nor U1159 (N_1159,N_688,N_998);
or U1160 (N_1160,N_525,In_1235);
xor U1161 (N_1161,In_818,In_734);
and U1162 (N_1162,N_494,N_770);
and U1163 (N_1163,N_898,N_906);
or U1164 (N_1164,N_866,N_121);
or U1165 (N_1165,N_892,In_364);
or U1166 (N_1166,N_803,In_201);
and U1167 (N_1167,N_592,N_471);
nor U1168 (N_1168,N_995,N_908);
nand U1169 (N_1169,N_913,N_727);
nand U1170 (N_1170,N_535,N_853);
nand U1171 (N_1171,N_968,In_1027);
or U1172 (N_1172,N_769,In_1156);
or U1173 (N_1173,N_778,N_804);
and U1174 (N_1174,N_758,N_631);
nor U1175 (N_1175,N_833,N_604);
and U1176 (N_1176,N_675,N_253);
and U1177 (N_1177,N_794,N_972);
or U1178 (N_1178,N_865,In_934);
nor U1179 (N_1179,N_826,N_969);
and U1180 (N_1180,N_896,N_861);
nand U1181 (N_1181,In_872,N_985);
nand U1182 (N_1182,N_723,N_819);
nand U1183 (N_1183,N_944,N_857);
nor U1184 (N_1184,In_702,In_977);
nand U1185 (N_1185,N_79,N_831);
or U1186 (N_1186,N_187,N_515);
nor U1187 (N_1187,N_697,N_796);
and U1188 (N_1188,N_686,N_942);
xor U1189 (N_1189,N_814,N_364);
nor U1190 (N_1190,N_610,In_1447);
and U1191 (N_1191,N_843,N_958);
and U1192 (N_1192,N_272,In_156);
xnor U1193 (N_1193,In_893,N_909);
nand U1194 (N_1194,N_916,N_827);
or U1195 (N_1195,N_933,N_810);
and U1196 (N_1196,In_861,N_792);
nor U1197 (N_1197,In_781,In_1451);
nand U1198 (N_1198,N_901,N_408);
or U1199 (N_1199,N_845,N_931);
or U1200 (N_1200,N_1137,N_410);
and U1201 (N_1201,N_1131,N_1014);
and U1202 (N_1202,N_1028,N_1093);
nand U1203 (N_1203,N_1063,N_950);
or U1204 (N_1204,N_917,N_929);
and U1205 (N_1205,N_1142,In_369);
or U1206 (N_1206,N_1118,N_1192);
nor U1207 (N_1207,N_959,N_1174);
nand U1208 (N_1208,N_781,N_1038);
nor U1209 (N_1209,N_1166,N_1160);
nand U1210 (N_1210,N_1196,N_497);
or U1211 (N_1211,N_1022,N_1066);
nand U1212 (N_1212,N_19,N_1170);
xor U1213 (N_1213,N_1065,N_1102);
xnor U1214 (N_1214,N_848,N_1047);
nor U1215 (N_1215,N_1026,N_1191);
nand U1216 (N_1216,N_1112,N_1108);
or U1217 (N_1217,N_1129,N_1147);
or U1218 (N_1218,N_574,N_1056);
and U1219 (N_1219,N_1075,N_1091);
or U1220 (N_1220,N_1182,N_1043);
or U1221 (N_1221,N_1099,N_841);
nand U1222 (N_1222,N_1069,N_502);
nand U1223 (N_1223,N_1036,N_1155);
and U1224 (N_1224,N_1079,N_239);
and U1225 (N_1225,N_1039,N_1133);
or U1226 (N_1226,N_1123,In_191);
nor U1227 (N_1227,In_630,In_102);
or U1228 (N_1228,N_1175,N_1134);
nor U1229 (N_1229,N_1144,N_1105);
or U1230 (N_1230,N_1163,In_259);
and U1231 (N_1231,In_468,N_1013);
and U1232 (N_1232,N_1148,N_1157);
or U1233 (N_1233,N_1130,N_1121);
or U1234 (N_1234,N_1045,N_799);
and U1235 (N_1235,N_1169,N_1081);
nand U1236 (N_1236,N_1084,N_1010);
nor U1237 (N_1237,N_1187,In_787);
and U1238 (N_1238,N_1100,N_900);
nand U1239 (N_1239,N_1083,N_1058);
and U1240 (N_1240,N_1179,N_1150);
nor U1241 (N_1241,In_1221,N_1041);
nor U1242 (N_1242,N_1011,N_1019);
and U1243 (N_1243,N_627,N_800);
nor U1244 (N_1244,N_13,N_966);
and U1245 (N_1245,N_823,N_864);
nor U1246 (N_1246,N_809,N_1034);
nor U1247 (N_1247,N_1141,N_1124);
and U1248 (N_1248,N_919,N_1113);
nor U1249 (N_1249,N_934,N_1178);
nor U1250 (N_1250,N_58,N_1127);
nand U1251 (N_1251,N_1165,N_1051);
and U1252 (N_1252,N_1031,N_990);
nand U1253 (N_1253,N_1024,N_1195);
xnor U1254 (N_1254,N_787,In_774);
nand U1255 (N_1255,N_1005,N_1061);
and U1256 (N_1256,N_1185,N_1159);
or U1257 (N_1257,N_1085,N_1009);
xor U1258 (N_1258,In_236,N_846);
nand U1259 (N_1259,N_1197,N_1015);
or U1260 (N_1260,N_825,N_584);
and U1261 (N_1261,N_1186,N_1003);
or U1262 (N_1262,N_1000,N_1128);
or U1263 (N_1263,N_88,N_185);
nor U1264 (N_1264,N_1153,N_1149);
nor U1265 (N_1265,N_738,N_1111);
nor U1266 (N_1266,N_1004,N_1177);
and U1267 (N_1267,N_1189,N_1119);
and U1268 (N_1268,N_139,N_1062);
nand U1269 (N_1269,N_941,In_135);
nand U1270 (N_1270,N_993,In_792);
and U1271 (N_1271,N_1046,N_562);
nor U1272 (N_1272,N_818,N_12);
xnor U1273 (N_1273,N_1073,N_1089);
nand U1274 (N_1274,In_471,N_1035);
or U1275 (N_1275,N_1135,N_1146);
nor U1276 (N_1276,N_1162,N_667);
and U1277 (N_1277,N_1098,N_1161);
nor U1278 (N_1278,N_1193,N_1082);
or U1279 (N_1279,N_1152,N_1122);
nand U1280 (N_1280,N_1188,N_1030);
xor U1281 (N_1281,N_1095,N_1064);
or U1282 (N_1282,N_1020,N_1067);
and U1283 (N_1283,N_1060,N_1044);
xor U1284 (N_1284,N_964,N_1183);
nand U1285 (N_1285,N_1094,N_1007);
xnor U1286 (N_1286,N_657,N_1103);
nand U1287 (N_1287,N_1145,N_369);
and U1288 (N_1288,N_1198,N_720);
and U1289 (N_1289,N_1037,N_1057);
and U1290 (N_1290,N_496,N_829);
nor U1291 (N_1291,N_1068,N_981);
and U1292 (N_1292,N_999,N_1027);
nand U1293 (N_1293,N_1109,N_881);
or U1294 (N_1294,N_1143,N_489);
and U1295 (N_1295,N_1114,N_777);
nor U1296 (N_1296,N_1072,N_988);
and U1297 (N_1297,N_603,N_1126);
or U1298 (N_1298,N_1052,N_1139);
and U1299 (N_1299,N_1097,N_957);
xor U1300 (N_1300,N_1017,N_977);
and U1301 (N_1301,N_858,In_679);
nor U1302 (N_1302,N_1042,N_1086);
or U1303 (N_1303,N_987,N_1107);
nor U1304 (N_1304,N_1025,N_1117);
nand U1305 (N_1305,N_1054,N_1055);
nand U1306 (N_1306,N_1087,N_980);
xor U1307 (N_1307,N_1012,N_1059);
or U1308 (N_1308,N_1154,N_1074);
nor U1309 (N_1309,N_882,In_687);
nor U1310 (N_1310,N_837,N_1176);
xor U1311 (N_1311,N_748,N_1190);
nand U1312 (N_1312,N_536,N_936);
xor U1313 (N_1313,N_1110,N_1125);
and U1314 (N_1314,N_1008,N_1001);
nand U1315 (N_1315,N_1115,N_1048);
nor U1316 (N_1316,N_1173,N_888);
and U1317 (N_1317,N_1172,N_1002);
nor U1318 (N_1318,N_1078,N_1049);
nand U1319 (N_1319,N_923,N_902);
nand U1320 (N_1320,N_961,N_807);
nor U1321 (N_1321,N_1021,N_1040);
nor U1322 (N_1322,N_1180,N_1033);
nand U1323 (N_1323,N_982,N_519);
and U1324 (N_1324,N_1168,N_918);
or U1325 (N_1325,N_1096,In_1404);
xor U1326 (N_1326,N_1092,N_1006);
and U1327 (N_1327,N_1023,N_1120);
or U1328 (N_1328,N_925,N_1151);
nor U1329 (N_1329,N_953,N_1140);
nand U1330 (N_1330,N_1032,N_1076);
nor U1331 (N_1331,N_1029,N_1101);
or U1332 (N_1332,N_1071,N_1070);
nor U1333 (N_1333,N_652,In_971);
xor U1334 (N_1334,N_1053,N_1016);
or U1335 (N_1335,N_1156,N_1167);
or U1336 (N_1336,In_810,N_1199);
nand U1337 (N_1337,N_1080,N_1088);
nand U1338 (N_1338,N_1158,N_1138);
nand U1339 (N_1339,N_1050,N_1171);
nand U1340 (N_1340,N_1018,N_1181);
or U1341 (N_1341,In_1473,N_1164);
nand U1342 (N_1342,N_764,N_1077);
and U1343 (N_1343,N_1104,N_1106);
nand U1344 (N_1344,N_1136,N_131);
xor U1345 (N_1345,N_1116,N_960);
and U1346 (N_1346,N_1090,N_1132);
nand U1347 (N_1347,N_1184,N_983);
nor U1348 (N_1348,N_1194,N_773);
nand U1349 (N_1349,N_303,N_880);
or U1350 (N_1350,N_1041,N_1104);
or U1351 (N_1351,N_1123,N_980);
nand U1352 (N_1352,N_1090,N_966);
nor U1353 (N_1353,N_1024,N_1149);
xor U1354 (N_1354,N_1016,N_748);
or U1355 (N_1355,N_1125,N_1051);
and U1356 (N_1356,N_1087,In_191);
or U1357 (N_1357,N_489,N_1018);
nor U1358 (N_1358,N_1040,N_1000);
nand U1359 (N_1359,N_1000,In_369);
nand U1360 (N_1360,N_562,N_1076);
and U1361 (N_1361,N_1142,N_1100);
nand U1362 (N_1362,N_1171,In_1473);
or U1363 (N_1363,N_1076,N_1148);
nor U1364 (N_1364,N_1038,N_1109);
nand U1365 (N_1365,N_1199,N_1120);
and U1366 (N_1366,N_1155,N_980);
nand U1367 (N_1367,N_980,N_1171);
nand U1368 (N_1368,N_139,N_1185);
and U1369 (N_1369,N_1009,N_1035);
and U1370 (N_1370,N_1079,N_1015);
and U1371 (N_1371,N_1134,N_496);
or U1372 (N_1372,N_139,N_1171);
and U1373 (N_1373,N_1135,N_800);
nand U1374 (N_1374,N_1036,N_858);
nand U1375 (N_1375,N_1064,N_627);
xnor U1376 (N_1376,In_468,In_810);
nand U1377 (N_1377,N_1160,N_1176);
nor U1378 (N_1378,N_1108,N_1098);
nor U1379 (N_1379,N_19,N_1139);
nor U1380 (N_1380,N_1174,N_864);
nor U1381 (N_1381,N_1188,N_1166);
or U1382 (N_1382,N_1106,N_1115);
nor U1383 (N_1383,N_1142,N_959);
nor U1384 (N_1384,N_1102,N_1034);
or U1385 (N_1385,N_1086,N_1187);
or U1386 (N_1386,N_1007,N_1148);
or U1387 (N_1387,N_1175,N_1079);
nand U1388 (N_1388,N_1063,N_1089);
or U1389 (N_1389,N_1089,N_1018);
nor U1390 (N_1390,N_1091,N_1120);
xor U1391 (N_1391,N_139,N_1175);
nor U1392 (N_1392,N_562,N_131);
nand U1393 (N_1393,N_1112,N_1188);
nand U1394 (N_1394,N_1079,N_1033);
nor U1395 (N_1395,N_1080,N_1123);
nor U1396 (N_1396,N_12,In_1221);
nor U1397 (N_1397,N_574,N_1175);
and U1398 (N_1398,N_1002,N_953);
and U1399 (N_1399,N_807,N_950);
xnor U1400 (N_1400,N_1397,N_1323);
or U1401 (N_1401,N_1254,N_1393);
or U1402 (N_1402,N_1211,N_1280);
or U1403 (N_1403,N_1225,N_1246);
and U1404 (N_1404,N_1299,N_1292);
nor U1405 (N_1405,N_1353,N_1286);
and U1406 (N_1406,N_1378,N_1228);
and U1407 (N_1407,N_1210,N_1373);
nor U1408 (N_1408,N_1328,N_1383);
nor U1409 (N_1409,N_1252,N_1304);
nand U1410 (N_1410,N_1321,N_1239);
nand U1411 (N_1411,N_1255,N_1291);
or U1412 (N_1412,N_1282,N_1352);
nor U1413 (N_1413,N_1266,N_1376);
nand U1414 (N_1414,N_1315,N_1271);
nor U1415 (N_1415,N_1256,N_1333);
xor U1416 (N_1416,N_1369,N_1263);
or U1417 (N_1417,N_1267,N_1327);
nor U1418 (N_1418,N_1275,N_1285);
nand U1419 (N_1419,N_1388,N_1350);
xnor U1420 (N_1420,N_1231,N_1355);
nor U1421 (N_1421,N_1365,N_1374);
and U1422 (N_1422,N_1340,N_1386);
and U1423 (N_1423,N_1213,N_1250);
nand U1424 (N_1424,N_1346,N_1313);
nand U1425 (N_1425,N_1284,N_1335);
xnor U1426 (N_1426,N_1202,N_1314);
nor U1427 (N_1427,N_1216,N_1243);
and U1428 (N_1428,N_1351,N_1311);
nor U1429 (N_1429,N_1370,N_1223);
and U1430 (N_1430,N_1205,N_1208);
nor U1431 (N_1431,N_1343,N_1371);
and U1432 (N_1432,N_1363,N_1203);
xor U1433 (N_1433,N_1245,N_1262);
and U1434 (N_1434,N_1310,N_1317);
or U1435 (N_1435,N_1390,N_1392);
and U1436 (N_1436,N_1247,N_1366);
nor U1437 (N_1437,N_1272,N_1395);
nand U1438 (N_1438,N_1394,N_1385);
nor U1439 (N_1439,N_1226,N_1207);
or U1440 (N_1440,N_1229,N_1359);
nor U1441 (N_1441,N_1294,N_1230);
nor U1442 (N_1442,N_1269,N_1259);
nor U1443 (N_1443,N_1288,N_1354);
or U1444 (N_1444,N_1204,N_1206);
nand U1445 (N_1445,N_1377,N_1325);
or U1446 (N_1446,N_1362,N_1358);
or U1447 (N_1447,N_1347,N_1212);
and U1448 (N_1448,N_1227,N_1372);
nand U1449 (N_1449,N_1233,N_1289);
or U1450 (N_1450,N_1274,N_1217);
nor U1451 (N_1451,N_1232,N_1221);
nand U1452 (N_1452,N_1242,N_1306);
nand U1453 (N_1453,N_1326,N_1375);
and U1454 (N_1454,N_1257,N_1222);
or U1455 (N_1455,N_1300,N_1384);
or U1456 (N_1456,N_1268,N_1215);
nand U1457 (N_1457,N_1324,N_1399);
or U1458 (N_1458,N_1200,N_1312);
and U1459 (N_1459,N_1293,N_1302);
nand U1460 (N_1460,N_1336,N_1330);
or U1461 (N_1461,N_1281,N_1261);
nor U1462 (N_1462,N_1339,N_1342);
nor U1463 (N_1463,N_1290,N_1277);
xnor U1464 (N_1464,N_1236,N_1244);
nor U1465 (N_1465,N_1367,N_1381);
nor U1466 (N_1466,N_1318,N_1276);
nor U1467 (N_1467,N_1331,N_1298);
and U1468 (N_1468,N_1389,N_1320);
nand U1469 (N_1469,N_1332,N_1224);
nand U1470 (N_1470,N_1237,N_1341);
and U1471 (N_1471,N_1308,N_1270);
or U1472 (N_1472,N_1219,N_1248);
or U1473 (N_1473,N_1348,N_1238);
and U1474 (N_1474,N_1218,N_1214);
or U1475 (N_1475,N_1361,N_1265);
and U1476 (N_1476,N_1279,N_1209);
nand U1477 (N_1477,N_1316,N_1258);
or U1478 (N_1478,N_1241,N_1338);
and U1479 (N_1479,N_1387,N_1360);
or U1480 (N_1480,N_1349,N_1380);
nand U1481 (N_1481,N_1297,N_1337);
nand U1482 (N_1482,N_1357,N_1260);
and U1483 (N_1483,N_1287,N_1382);
nand U1484 (N_1484,N_1398,N_1307);
or U1485 (N_1485,N_1379,N_1296);
nand U1486 (N_1486,N_1283,N_1391);
and U1487 (N_1487,N_1396,N_1364);
and U1488 (N_1488,N_1249,N_1273);
xnor U1489 (N_1489,N_1235,N_1301);
and U1490 (N_1490,N_1251,N_1303);
xor U1491 (N_1491,N_1278,N_1345);
nor U1492 (N_1492,N_1334,N_1344);
and U1493 (N_1493,N_1309,N_1295);
nand U1494 (N_1494,N_1322,N_1253);
and U1495 (N_1495,N_1368,N_1305);
and U1496 (N_1496,N_1201,N_1220);
or U1497 (N_1497,N_1240,N_1319);
nor U1498 (N_1498,N_1234,N_1356);
nor U1499 (N_1499,N_1264,N_1329);
and U1500 (N_1500,N_1252,N_1396);
or U1501 (N_1501,N_1290,N_1216);
nor U1502 (N_1502,N_1290,N_1303);
nor U1503 (N_1503,N_1231,N_1311);
nand U1504 (N_1504,N_1292,N_1304);
or U1505 (N_1505,N_1305,N_1317);
and U1506 (N_1506,N_1209,N_1284);
nand U1507 (N_1507,N_1211,N_1305);
xnor U1508 (N_1508,N_1247,N_1203);
and U1509 (N_1509,N_1393,N_1332);
or U1510 (N_1510,N_1238,N_1316);
nand U1511 (N_1511,N_1234,N_1360);
nor U1512 (N_1512,N_1395,N_1238);
nor U1513 (N_1513,N_1211,N_1272);
nor U1514 (N_1514,N_1204,N_1262);
xnor U1515 (N_1515,N_1349,N_1301);
nor U1516 (N_1516,N_1318,N_1344);
nor U1517 (N_1517,N_1397,N_1305);
nand U1518 (N_1518,N_1282,N_1226);
nor U1519 (N_1519,N_1231,N_1392);
nand U1520 (N_1520,N_1259,N_1397);
nand U1521 (N_1521,N_1375,N_1234);
or U1522 (N_1522,N_1250,N_1378);
and U1523 (N_1523,N_1305,N_1385);
or U1524 (N_1524,N_1346,N_1275);
nor U1525 (N_1525,N_1216,N_1378);
xnor U1526 (N_1526,N_1376,N_1283);
or U1527 (N_1527,N_1265,N_1268);
nand U1528 (N_1528,N_1374,N_1390);
nor U1529 (N_1529,N_1328,N_1320);
nand U1530 (N_1530,N_1372,N_1280);
nand U1531 (N_1531,N_1203,N_1254);
xnor U1532 (N_1532,N_1350,N_1329);
nand U1533 (N_1533,N_1326,N_1236);
and U1534 (N_1534,N_1377,N_1364);
nand U1535 (N_1535,N_1284,N_1277);
nor U1536 (N_1536,N_1347,N_1246);
and U1537 (N_1537,N_1262,N_1218);
nor U1538 (N_1538,N_1272,N_1319);
and U1539 (N_1539,N_1354,N_1389);
nand U1540 (N_1540,N_1371,N_1203);
and U1541 (N_1541,N_1363,N_1319);
and U1542 (N_1542,N_1291,N_1268);
or U1543 (N_1543,N_1370,N_1212);
or U1544 (N_1544,N_1363,N_1242);
and U1545 (N_1545,N_1207,N_1359);
and U1546 (N_1546,N_1224,N_1212);
and U1547 (N_1547,N_1236,N_1338);
nand U1548 (N_1548,N_1379,N_1365);
nor U1549 (N_1549,N_1347,N_1344);
or U1550 (N_1550,N_1281,N_1392);
nor U1551 (N_1551,N_1209,N_1392);
and U1552 (N_1552,N_1271,N_1288);
and U1553 (N_1553,N_1342,N_1382);
nand U1554 (N_1554,N_1240,N_1247);
or U1555 (N_1555,N_1325,N_1239);
nand U1556 (N_1556,N_1281,N_1356);
nand U1557 (N_1557,N_1305,N_1379);
or U1558 (N_1558,N_1382,N_1236);
nor U1559 (N_1559,N_1388,N_1331);
or U1560 (N_1560,N_1253,N_1341);
nand U1561 (N_1561,N_1346,N_1231);
or U1562 (N_1562,N_1319,N_1388);
nand U1563 (N_1563,N_1296,N_1298);
nor U1564 (N_1564,N_1363,N_1280);
and U1565 (N_1565,N_1293,N_1310);
or U1566 (N_1566,N_1348,N_1245);
and U1567 (N_1567,N_1283,N_1237);
and U1568 (N_1568,N_1326,N_1309);
nor U1569 (N_1569,N_1342,N_1368);
nand U1570 (N_1570,N_1235,N_1304);
and U1571 (N_1571,N_1256,N_1208);
or U1572 (N_1572,N_1249,N_1365);
and U1573 (N_1573,N_1272,N_1214);
nand U1574 (N_1574,N_1249,N_1339);
nand U1575 (N_1575,N_1221,N_1333);
xnor U1576 (N_1576,N_1324,N_1210);
or U1577 (N_1577,N_1333,N_1376);
nand U1578 (N_1578,N_1319,N_1236);
nand U1579 (N_1579,N_1389,N_1252);
or U1580 (N_1580,N_1347,N_1376);
xnor U1581 (N_1581,N_1333,N_1239);
nand U1582 (N_1582,N_1269,N_1300);
nand U1583 (N_1583,N_1340,N_1269);
or U1584 (N_1584,N_1301,N_1230);
or U1585 (N_1585,N_1227,N_1247);
nand U1586 (N_1586,N_1287,N_1311);
and U1587 (N_1587,N_1349,N_1342);
xnor U1588 (N_1588,N_1397,N_1380);
or U1589 (N_1589,N_1345,N_1261);
or U1590 (N_1590,N_1335,N_1310);
nor U1591 (N_1591,N_1270,N_1255);
or U1592 (N_1592,N_1361,N_1312);
and U1593 (N_1593,N_1288,N_1314);
nand U1594 (N_1594,N_1283,N_1224);
nand U1595 (N_1595,N_1362,N_1329);
and U1596 (N_1596,N_1390,N_1235);
nor U1597 (N_1597,N_1327,N_1315);
nor U1598 (N_1598,N_1223,N_1255);
nand U1599 (N_1599,N_1298,N_1203);
nor U1600 (N_1600,N_1467,N_1476);
and U1601 (N_1601,N_1464,N_1479);
nand U1602 (N_1602,N_1552,N_1412);
and U1603 (N_1603,N_1572,N_1598);
and U1604 (N_1604,N_1516,N_1430);
nor U1605 (N_1605,N_1514,N_1558);
nand U1606 (N_1606,N_1589,N_1526);
nor U1607 (N_1607,N_1454,N_1532);
nor U1608 (N_1608,N_1455,N_1594);
nor U1609 (N_1609,N_1521,N_1474);
nor U1610 (N_1610,N_1425,N_1563);
nor U1611 (N_1611,N_1446,N_1411);
xor U1612 (N_1612,N_1562,N_1555);
or U1613 (N_1613,N_1596,N_1488);
and U1614 (N_1614,N_1568,N_1544);
or U1615 (N_1615,N_1546,N_1583);
xnor U1616 (N_1616,N_1553,N_1566);
xor U1617 (N_1617,N_1484,N_1409);
and U1618 (N_1618,N_1591,N_1577);
xor U1619 (N_1619,N_1402,N_1441);
nor U1620 (N_1620,N_1404,N_1584);
nor U1621 (N_1621,N_1472,N_1469);
nor U1622 (N_1622,N_1590,N_1510);
or U1623 (N_1623,N_1452,N_1501);
and U1624 (N_1624,N_1458,N_1406);
nor U1625 (N_1625,N_1439,N_1509);
or U1626 (N_1626,N_1459,N_1473);
or U1627 (N_1627,N_1530,N_1560);
nor U1628 (N_1628,N_1426,N_1448);
nand U1629 (N_1629,N_1528,N_1585);
xnor U1630 (N_1630,N_1453,N_1445);
nor U1631 (N_1631,N_1486,N_1400);
nand U1632 (N_1632,N_1414,N_1434);
nand U1633 (N_1633,N_1432,N_1468);
nor U1634 (N_1634,N_1511,N_1408);
nand U1635 (N_1635,N_1498,N_1569);
and U1636 (N_1636,N_1461,N_1531);
nor U1637 (N_1637,N_1597,N_1418);
or U1638 (N_1638,N_1524,N_1493);
and U1639 (N_1639,N_1465,N_1559);
nand U1640 (N_1640,N_1547,N_1576);
and U1641 (N_1641,N_1462,N_1429);
nand U1642 (N_1642,N_1415,N_1470);
and U1643 (N_1643,N_1595,N_1548);
nand U1644 (N_1644,N_1580,N_1499);
or U1645 (N_1645,N_1512,N_1539);
nand U1646 (N_1646,N_1503,N_1575);
xnor U1647 (N_1647,N_1423,N_1450);
nor U1648 (N_1648,N_1478,N_1490);
and U1649 (N_1649,N_1574,N_1534);
nand U1650 (N_1650,N_1401,N_1554);
nand U1651 (N_1651,N_1550,N_1403);
nand U1652 (N_1652,N_1485,N_1567);
nor U1653 (N_1653,N_1570,N_1556);
and U1654 (N_1654,N_1471,N_1542);
or U1655 (N_1655,N_1435,N_1447);
nor U1656 (N_1656,N_1578,N_1494);
nor U1657 (N_1657,N_1571,N_1424);
nand U1658 (N_1658,N_1482,N_1508);
and U1659 (N_1659,N_1599,N_1500);
and U1660 (N_1660,N_1419,N_1422);
nor U1661 (N_1661,N_1517,N_1565);
nor U1662 (N_1662,N_1525,N_1410);
xnor U1663 (N_1663,N_1449,N_1438);
or U1664 (N_1664,N_1475,N_1495);
or U1665 (N_1665,N_1579,N_1480);
or U1666 (N_1666,N_1523,N_1431);
and U1667 (N_1667,N_1551,N_1491);
nor U1668 (N_1668,N_1513,N_1545);
nand U1669 (N_1669,N_1443,N_1515);
and U1670 (N_1670,N_1483,N_1538);
nand U1671 (N_1671,N_1540,N_1405);
nand U1672 (N_1672,N_1536,N_1502);
nor U1673 (N_1673,N_1433,N_1421);
nor U1674 (N_1674,N_1504,N_1587);
nor U1675 (N_1675,N_1573,N_1477);
and U1676 (N_1676,N_1507,N_1420);
or U1677 (N_1677,N_1588,N_1535);
nor U1678 (N_1678,N_1487,N_1537);
xnor U1679 (N_1679,N_1442,N_1413);
and U1680 (N_1680,N_1543,N_1586);
or U1681 (N_1681,N_1451,N_1437);
and U1682 (N_1682,N_1527,N_1557);
nand U1683 (N_1683,N_1456,N_1549);
and U1684 (N_1684,N_1463,N_1520);
nor U1685 (N_1685,N_1506,N_1460);
or U1686 (N_1686,N_1593,N_1417);
nor U1687 (N_1687,N_1496,N_1466);
nor U1688 (N_1688,N_1561,N_1407);
nand U1689 (N_1689,N_1436,N_1444);
or U1690 (N_1690,N_1533,N_1492);
xor U1691 (N_1691,N_1427,N_1428);
and U1692 (N_1692,N_1564,N_1489);
nor U1693 (N_1693,N_1522,N_1519);
nor U1694 (N_1694,N_1497,N_1529);
and U1695 (N_1695,N_1592,N_1457);
nand U1696 (N_1696,N_1481,N_1581);
nor U1697 (N_1697,N_1582,N_1541);
nor U1698 (N_1698,N_1440,N_1505);
and U1699 (N_1699,N_1416,N_1518);
and U1700 (N_1700,N_1519,N_1579);
nand U1701 (N_1701,N_1565,N_1493);
and U1702 (N_1702,N_1429,N_1515);
or U1703 (N_1703,N_1442,N_1474);
xnor U1704 (N_1704,N_1522,N_1545);
nand U1705 (N_1705,N_1499,N_1469);
xor U1706 (N_1706,N_1531,N_1554);
or U1707 (N_1707,N_1511,N_1471);
or U1708 (N_1708,N_1583,N_1526);
nor U1709 (N_1709,N_1527,N_1424);
nand U1710 (N_1710,N_1468,N_1579);
xor U1711 (N_1711,N_1540,N_1409);
nor U1712 (N_1712,N_1445,N_1573);
and U1713 (N_1713,N_1435,N_1567);
xor U1714 (N_1714,N_1503,N_1506);
nand U1715 (N_1715,N_1504,N_1469);
nor U1716 (N_1716,N_1562,N_1567);
or U1717 (N_1717,N_1545,N_1597);
or U1718 (N_1718,N_1497,N_1475);
nor U1719 (N_1719,N_1500,N_1455);
or U1720 (N_1720,N_1454,N_1418);
or U1721 (N_1721,N_1553,N_1458);
nand U1722 (N_1722,N_1494,N_1553);
nor U1723 (N_1723,N_1560,N_1413);
nor U1724 (N_1724,N_1572,N_1514);
nand U1725 (N_1725,N_1490,N_1565);
and U1726 (N_1726,N_1446,N_1561);
nor U1727 (N_1727,N_1485,N_1573);
xnor U1728 (N_1728,N_1439,N_1472);
and U1729 (N_1729,N_1597,N_1533);
nand U1730 (N_1730,N_1468,N_1590);
nand U1731 (N_1731,N_1526,N_1580);
nor U1732 (N_1732,N_1533,N_1544);
nor U1733 (N_1733,N_1537,N_1426);
nor U1734 (N_1734,N_1499,N_1528);
nor U1735 (N_1735,N_1592,N_1506);
xnor U1736 (N_1736,N_1595,N_1464);
nand U1737 (N_1737,N_1401,N_1446);
and U1738 (N_1738,N_1433,N_1477);
and U1739 (N_1739,N_1527,N_1410);
and U1740 (N_1740,N_1440,N_1510);
or U1741 (N_1741,N_1477,N_1565);
or U1742 (N_1742,N_1416,N_1590);
xor U1743 (N_1743,N_1539,N_1563);
nand U1744 (N_1744,N_1559,N_1431);
nor U1745 (N_1745,N_1596,N_1425);
xnor U1746 (N_1746,N_1596,N_1464);
or U1747 (N_1747,N_1457,N_1553);
and U1748 (N_1748,N_1401,N_1549);
nand U1749 (N_1749,N_1413,N_1553);
and U1750 (N_1750,N_1410,N_1496);
nand U1751 (N_1751,N_1507,N_1527);
nor U1752 (N_1752,N_1413,N_1434);
nand U1753 (N_1753,N_1569,N_1587);
and U1754 (N_1754,N_1594,N_1565);
nand U1755 (N_1755,N_1427,N_1519);
and U1756 (N_1756,N_1532,N_1405);
nor U1757 (N_1757,N_1556,N_1457);
nor U1758 (N_1758,N_1579,N_1438);
nor U1759 (N_1759,N_1530,N_1455);
and U1760 (N_1760,N_1515,N_1478);
and U1761 (N_1761,N_1528,N_1458);
and U1762 (N_1762,N_1470,N_1524);
or U1763 (N_1763,N_1504,N_1466);
nor U1764 (N_1764,N_1410,N_1416);
xor U1765 (N_1765,N_1568,N_1412);
or U1766 (N_1766,N_1454,N_1489);
nand U1767 (N_1767,N_1524,N_1459);
nor U1768 (N_1768,N_1535,N_1483);
nand U1769 (N_1769,N_1431,N_1542);
nand U1770 (N_1770,N_1443,N_1585);
or U1771 (N_1771,N_1558,N_1492);
and U1772 (N_1772,N_1522,N_1410);
nor U1773 (N_1773,N_1441,N_1419);
or U1774 (N_1774,N_1591,N_1457);
and U1775 (N_1775,N_1424,N_1493);
nor U1776 (N_1776,N_1400,N_1542);
or U1777 (N_1777,N_1486,N_1565);
xor U1778 (N_1778,N_1489,N_1558);
or U1779 (N_1779,N_1563,N_1442);
nor U1780 (N_1780,N_1579,N_1556);
and U1781 (N_1781,N_1571,N_1518);
and U1782 (N_1782,N_1443,N_1582);
or U1783 (N_1783,N_1557,N_1516);
xnor U1784 (N_1784,N_1588,N_1560);
nand U1785 (N_1785,N_1458,N_1401);
nor U1786 (N_1786,N_1480,N_1586);
and U1787 (N_1787,N_1443,N_1490);
nor U1788 (N_1788,N_1544,N_1449);
or U1789 (N_1789,N_1546,N_1554);
and U1790 (N_1790,N_1436,N_1560);
and U1791 (N_1791,N_1504,N_1502);
or U1792 (N_1792,N_1589,N_1598);
nor U1793 (N_1793,N_1496,N_1561);
nand U1794 (N_1794,N_1594,N_1598);
and U1795 (N_1795,N_1494,N_1434);
nor U1796 (N_1796,N_1401,N_1553);
nand U1797 (N_1797,N_1424,N_1488);
xnor U1798 (N_1798,N_1589,N_1512);
nand U1799 (N_1799,N_1471,N_1545);
nor U1800 (N_1800,N_1723,N_1708);
or U1801 (N_1801,N_1693,N_1638);
xnor U1802 (N_1802,N_1667,N_1771);
nor U1803 (N_1803,N_1730,N_1753);
nand U1804 (N_1804,N_1651,N_1738);
nor U1805 (N_1805,N_1684,N_1650);
or U1806 (N_1806,N_1659,N_1647);
and U1807 (N_1807,N_1774,N_1645);
nor U1808 (N_1808,N_1787,N_1688);
or U1809 (N_1809,N_1782,N_1766);
nand U1810 (N_1810,N_1664,N_1672);
nor U1811 (N_1811,N_1656,N_1663);
nor U1812 (N_1812,N_1754,N_1660);
or U1813 (N_1813,N_1750,N_1704);
and U1814 (N_1814,N_1669,N_1763);
or U1815 (N_1815,N_1791,N_1760);
nor U1816 (N_1816,N_1628,N_1713);
or U1817 (N_1817,N_1728,N_1602);
and U1818 (N_1818,N_1739,N_1797);
nor U1819 (N_1819,N_1712,N_1700);
or U1820 (N_1820,N_1743,N_1625);
xor U1821 (N_1821,N_1691,N_1703);
or U1822 (N_1822,N_1758,N_1634);
nand U1823 (N_1823,N_1781,N_1720);
nand U1824 (N_1824,N_1749,N_1779);
or U1825 (N_1825,N_1614,N_1642);
nand U1826 (N_1826,N_1671,N_1610);
nor U1827 (N_1827,N_1711,N_1715);
nor U1828 (N_1828,N_1780,N_1694);
nor U1829 (N_1829,N_1777,N_1640);
or U1830 (N_1830,N_1626,N_1689);
nor U1831 (N_1831,N_1662,N_1658);
or U1832 (N_1832,N_1615,N_1717);
and U1833 (N_1833,N_1621,N_1727);
nand U1834 (N_1834,N_1605,N_1761);
and U1835 (N_1835,N_1646,N_1709);
or U1836 (N_1836,N_1746,N_1632);
nor U1837 (N_1837,N_1710,N_1795);
nor U1838 (N_1838,N_1606,N_1719);
nor U1839 (N_1839,N_1769,N_1794);
nand U1840 (N_1840,N_1724,N_1695);
xor U1841 (N_1841,N_1751,N_1613);
nor U1842 (N_1842,N_1764,N_1740);
and U1843 (N_1843,N_1698,N_1648);
nor U1844 (N_1844,N_1798,N_1643);
and U1845 (N_1845,N_1603,N_1745);
or U1846 (N_1846,N_1734,N_1661);
nand U1847 (N_1847,N_1776,N_1668);
or U1848 (N_1848,N_1696,N_1726);
and U1849 (N_1849,N_1762,N_1619);
nand U1850 (N_1850,N_1670,N_1759);
xor U1851 (N_1851,N_1630,N_1692);
and U1852 (N_1852,N_1639,N_1756);
and U1853 (N_1853,N_1673,N_1778);
or U1854 (N_1854,N_1600,N_1631);
and U1855 (N_1855,N_1636,N_1683);
and U1856 (N_1856,N_1623,N_1737);
or U1857 (N_1857,N_1767,N_1652);
nor U1858 (N_1858,N_1706,N_1624);
or U1859 (N_1859,N_1616,N_1792);
nor U1860 (N_1860,N_1609,N_1747);
nor U1861 (N_1861,N_1686,N_1665);
and U1862 (N_1862,N_1680,N_1783);
or U1863 (N_1863,N_1718,N_1620);
nor U1864 (N_1864,N_1770,N_1666);
or U1865 (N_1865,N_1702,N_1654);
or U1866 (N_1866,N_1629,N_1607);
or U1867 (N_1867,N_1752,N_1641);
nor U1868 (N_1868,N_1784,N_1681);
and U1869 (N_1869,N_1608,N_1655);
nand U1870 (N_1870,N_1678,N_1796);
and U1871 (N_1871,N_1675,N_1799);
and U1872 (N_1872,N_1627,N_1772);
nand U1873 (N_1873,N_1785,N_1657);
or U1874 (N_1874,N_1611,N_1676);
and U1875 (N_1875,N_1635,N_1790);
and U1876 (N_1876,N_1765,N_1775);
or U1877 (N_1877,N_1682,N_1788);
nor U1878 (N_1878,N_1729,N_1741);
nand U1879 (N_1879,N_1707,N_1721);
xor U1880 (N_1880,N_1725,N_1679);
nand U1881 (N_1881,N_1768,N_1755);
nor U1882 (N_1882,N_1612,N_1617);
and U1883 (N_1883,N_1644,N_1622);
nor U1884 (N_1884,N_1649,N_1735);
and U1885 (N_1885,N_1786,N_1697);
xor U1886 (N_1886,N_1601,N_1705);
xor U1887 (N_1887,N_1732,N_1742);
xnor U1888 (N_1888,N_1748,N_1618);
nand U1889 (N_1889,N_1793,N_1789);
nand U1890 (N_1890,N_1653,N_1685);
or U1891 (N_1891,N_1690,N_1674);
nand U1892 (N_1892,N_1699,N_1714);
nand U1893 (N_1893,N_1637,N_1731);
nand U1894 (N_1894,N_1757,N_1604);
nor U1895 (N_1895,N_1736,N_1701);
nand U1896 (N_1896,N_1733,N_1633);
and U1897 (N_1897,N_1722,N_1687);
nand U1898 (N_1898,N_1744,N_1677);
nand U1899 (N_1899,N_1716,N_1773);
nand U1900 (N_1900,N_1665,N_1715);
nor U1901 (N_1901,N_1799,N_1629);
or U1902 (N_1902,N_1600,N_1763);
or U1903 (N_1903,N_1621,N_1728);
xnor U1904 (N_1904,N_1651,N_1685);
nand U1905 (N_1905,N_1768,N_1671);
and U1906 (N_1906,N_1644,N_1663);
nand U1907 (N_1907,N_1608,N_1710);
and U1908 (N_1908,N_1673,N_1735);
nor U1909 (N_1909,N_1750,N_1610);
and U1910 (N_1910,N_1703,N_1662);
xor U1911 (N_1911,N_1768,N_1794);
xor U1912 (N_1912,N_1665,N_1643);
nand U1913 (N_1913,N_1649,N_1622);
and U1914 (N_1914,N_1645,N_1672);
nor U1915 (N_1915,N_1781,N_1749);
or U1916 (N_1916,N_1639,N_1799);
and U1917 (N_1917,N_1797,N_1682);
nor U1918 (N_1918,N_1727,N_1619);
or U1919 (N_1919,N_1691,N_1639);
nor U1920 (N_1920,N_1740,N_1773);
and U1921 (N_1921,N_1781,N_1649);
nand U1922 (N_1922,N_1712,N_1791);
nor U1923 (N_1923,N_1787,N_1730);
and U1924 (N_1924,N_1725,N_1790);
and U1925 (N_1925,N_1699,N_1753);
nand U1926 (N_1926,N_1637,N_1659);
nor U1927 (N_1927,N_1639,N_1690);
or U1928 (N_1928,N_1706,N_1691);
and U1929 (N_1929,N_1745,N_1779);
nand U1930 (N_1930,N_1675,N_1691);
nand U1931 (N_1931,N_1739,N_1658);
nand U1932 (N_1932,N_1729,N_1721);
nand U1933 (N_1933,N_1731,N_1756);
and U1934 (N_1934,N_1638,N_1642);
and U1935 (N_1935,N_1690,N_1697);
or U1936 (N_1936,N_1700,N_1793);
xor U1937 (N_1937,N_1793,N_1715);
or U1938 (N_1938,N_1655,N_1778);
xor U1939 (N_1939,N_1776,N_1766);
nor U1940 (N_1940,N_1727,N_1620);
nor U1941 (N_1941,N_1687,N_1667);
or U1942 (N_1942,N_1772,N_1660);
and U1943 (N_1943,N_1684,N_1777);
or U1944 (N_1944,N_1600,N_1774);
nor U1945 (N_1945,N_1789,N_1605);
nor U1946 (N_1946,N_1695,N_1608);
or U1947 (N_1947,N_1780,N_1739);
nor U1948 (N_1948,N_1702,N_1630);
nand U1949 (N_1949,N_1634,N_1607);
or U1950 (N_1950,N_1617,N_1732);
or U1951 (N_1951,N_1704,N_1725);
nor U1952 (N_1952,N_1700,N_1772);
xnor U1953 (N_1953,N_1650,N_1713);
and U1954 (N_1954,N_1751,N_1719);
or U1955 (N_1955,N_1773,N_1708);
nand U1956 (N_1956,N_1667,N_1712);
nand U1957 (N_1957,N_1780,N_1775);
nand U1958 (N_1958,N_1767,N_1780);
nor U1959 (N_1959,N_1720,N_1692);
nor U1960 (N_1960,N_1752,N_1748);
and U1961 (N_1961,N_1637,N_1762);
xor U1962 (N_1962,N_1664,N_1701);
nor U1963 (N_1963,N_1766,N_1779);
and U1964 (N_1964,N_1731,N_1645);
and U1965 (N_1965,N_1758,N_1644);
or U1966 (N_1966,N_1602,N_1702);
and U1967 (N_1967,N_1751,N_1614);
nand U1968 (N_1968,N_1768,N_1700);
and U1969 (N_1969,N_1623,N_1686);
nand U1970 (N_1970,N_1785,N_1737);
or U1971 (N_1971,N_1748,N_1705);
xor U1972 (N_1972,N_1616,N_1724);
or U1973 (N_1973,N_1700,N_1688);
and U1974 (N_1974,N_1725,N_1783);
and U1975 (N_1975,N_1770,N_1631);
nand U1976 (N_1976,N_1600,N_1602);
nand U1977 (N_1977,N_1607,N_1760);
or U1978 (N_1978,N_1759,N_1760);
nand U1979 (N_1979,N_1624,N_1731);
and U1980 (N_1980,N_1722,N_1620);
nand U1981 (N_1981,N_1649,N_1710);
nor U1982 (N_1982,N_1672,N_1715);
or U1983 (N_1983,N_1705,N_1676);
or U1984 (N_1984,N_1747,N_1657);
or U1985 (N_1985,N_1763,N_1741);
xor U1986 (N_1986,N_1798,N_1637);
nor U1987 (N_1987,N_1699,N_1709);
and U1988 (N_1988,N_1792,N_1697);
nand U1989 (N_1989,N_1679,N_1791);
nand U1990 (N_1990,N_1625,N_1717);
or U1991 (N_1991,N_1707,N_1735);
nor U1992 (N_1992,N_1668,N_1693);
nand U1993 (N_1993,N_1721,N_1671);
nand U1994 (N_1994,N_1738,N_1713);
nand U1995 (N_1995,N_1733,N_1741);
nand U1996 (N_1996,N_1733,N_1651);
nor U1997 (N_1997,N_1677,N_1651);
and U1998 (N_1998,N_1775,N_1707);
or U1999 (N_1999,N_1789,N_1766);
or U2000 (N_2000,N_1958,N_1811);
nor U2001 (N_2001,N_1857,N_1942);
xnor U2002 (N_2002,N_1880,N_1921);
nor U2003 (N_2003,N_1978,N_1931);
or U2004 (N_2004,N_1974,N_1887);
nor U2005 (N_2005,N_1806,N_1877);
nand U2006 (N_2006,N_1849,N_1839);
nand U2007 (N_2007,N_1935,N_1982);
nand U2008 (N_2008,N_1813,N_1818);
and U2009 (N_2009,N_1967,N_1843);
nand U2010 (N_2010,N_1841,N_1976);
nand U2011 (N_2011,N_1896,N_1916);
nor U2012 (N_2012,N_1973,N_1847);
nand U2013 (N_2013,N_1885,N_1977);
nand U2014 (N_2014,N_1985,N_1927);
nor U2015 (N_2015,N_1999,N_1997);
or U2016 (N_2016,N_1986,N_1914);
nor U2017 (N_2017,N_1901,N_1953);
and U2018 (N_2018,N_1956,N_1913);
nand U2019 (N_2019,N_1981,N_1949);
or U2020 (N_2020,N_1966,N_1906);
nor U2021 (N_2021,N_1915,N_1988);
and U2022 (N_2022,N_1894,N_1874);
or U2023 (N_2023,N_1941,N_1882);
and U2024 (N_2024,N_1859,N_1808);
nand U2025 (N_2025,N_1917,N_1904);
and U2026 (N_2026,N_1911,N_1893);
and U2027 (N_2027,N_1844,N_1993);
nor U2028 (N_2028,N_1952,N_1903);
nand U2029 (N_2029,N_1828,N_1970);
nand U2030 (N_2030,N_1838,N_1898);
and U2031 (N_2031,N_1872,N_1825);
nor U2032 (N_2032,N_1922,N_1855);
nand U2033 (N_2033,N_1902,N_1946);
and U2034 (N_2034,N_1814,N_1868);
or U2035 (N_2035,N_1819,N_1939);
or U2036 (N_2036,N_1856,N_1969);
or U2037 (N_2037,N_1905,N_1960);
and U2038 (N_2038,N_1832,N_1860);
nor U2039 (N_2039,N_1979,N_1842);
and U2040 (N_2040,N_1823,N_1907);
and U2041 (N_2041,N_1957,N_1807);
and U2042 (N_2042,N_1987,N_1983);
or U2043 (N_2043,N_1912,N_1802);
nor U2044 (N_2044,N_1940,N_1918);
nand U2045 (N_2045,N_1937,N_1889);
nor U2046 (N_2046,N_1833,N_1925);
or U2047 (N_2047,N_1870,N_1845);
nor U2048 (N_2048,N_1884,N_1920);
nor U2049 (N_2049,N_1871,N_1876);
nand U2050 (N_2050,N_1895,N_1869);
nand U2051 (N_2051,N_1950,N_1848);
nand U2052 (N_2052,N_1955,N_1980);
or U2053 (N_2053,N_1899,N_1824);
and U2054 (N_2054,N_1908,N_1968);
and U2055 (N_2055,N_1867,N_1883);
nor U2056 (N_2056,N_1989,N_1801);
or U2057 (N_2057,N_1829,N_1810);
nor U2058 (N_2058,N_1864,N_1850);
or U2059 (N_2059,N_1831,N_1826);
nand U2060 (N_2060,N_1984,N_1944);
or U2061 (N_2061,N_1892,N_1800);
nor U2062 (N_2062,N_1804,N_1900);
nor U2063 (N_2063,N_1962,N_1865);
nand U2064 (N_2064,N_1861,N_1835);
and U2065 (N_2065,N_1858,N_1992);
or U2066 (N_2066,N_1852,N_1951);
and U2067 (N_2067,N_1875,N_1878);
nand U2068 (N_2068,N_1821,N_1866);
nor U2069 (N_2069,N_1924,N_1990);
and U2070 (N_2070,N_1954,N_1890);
nor U2071 (N_2071,N_1995,N_1961);
nor U2072 (N_2072,N_1827,N_1873);
nand U2073 (N_2073,N_1936,N_1948);
nand U2074 (N_2074,N_1972,N_1945);
nand U2075 (N_2075,N_1971,N_1854);
and U2076 (N_2076,N_1963,N_1933);
nor U2077 (N_2077,N_1923,N_1932);
or U2078 (N_2078,N_1817,N_1846);
and U2079 (N_2079,N_1809,N_1879);
nor U2080 (N_2080,N_1805,N_1919);
or U2081 (N_2081,N_1851,N_1815);
or U2082 (N_2082,N_1840,N_1928);
xor U2083 (N_2083,N_1886,N_1965);
and U2084 (N_2084,N_1930,N_1991);
and U2085 (N_2085,N_1964,N_1897);
or U2086 (N_2086,N_1943,N_1959);
nand U2087 (N_2087,N_1888,N_1837);
and U2088 (N_2088,N_1994,N_1934);
nand U2089 (N_2089,N_1938,N_1820);
nor U2090 (N_2090,N_1803,N_1862);
or U2091 (N_2091,N_1812,N_1881);
or U2092 (N_2092,N_1926,N_1836);
nor U2093 (N_2093,N_1909,N_1998);
nand U2094 (N_2094,N_1996,N_1891);
nor U2095 (N_2095,N_1947,N_1834);
nor U2096 (N_2096,N_1830,N_1816);
nor U2097 (N_2097,N_1910,N_1853);
nor U2098 (N_2098,N_1822,N_1975);
nand U2099 (N_2099,N_1929,N_1863);
nand U2100 (N_2100,N_1883,N_1988);
nor U2101 (N_2101,N_1832,N_1974);
nor U2102 (N_2102,N_1804,N_1997);
nor U2103 (N_2103,N_1934,N_1944);
nand U2104 (N_2104,N_1814,N_1984);
or U2105 (N_2105,N_1915,N_1908);
or U2106 (N_2106,N_1990,N_1816);
or U2107 (N_2107,N_1995,N_1970);
or U2108 (N_2108,N_1825,N_1908);
nor U2109 (N_2109,N_1860,N_1856);
nor U2110 (N_2110,N_1858,N_1863);
nor U2111 (N_2111,N_1864,N_1806);
xnor U2112 (N_2112,N_1913,N_1925);
nor U2113 (N_2113,N_1846,N_1903);
and U2114 (N_2114,N_1962,N_1908);
and U2115 (N_2115,N_1826,N_1899);
nand U2116 (N_2116,N_1959,N_1892);
nor U2117 (N_2117,N_1934,N_1899);
nand U2118 (N_2118,N_1804,N_1884);
or U2119 (N_2119,N_1925,N_1970);
and U2120 (N_2120,N_1848,N_1932);
or U2121 (N_2121,N_1822,N_1878);
nor U2122 (N_2122,N_1956,N_1844);
xor U2123 (N_2123,N_1930,N_1885);
nor U2124 (N_2124,N_1877,N_1878);
nor U2125 (N_2125,N_1807,N_1843);
nor U2126 (N_2126,N_1862,N_1889);
nor U2127 (N_2127,N_1872,N_1954);
nor U2128 (N_2128,N_1845,N_1972);
or U2129 (N_2129,N_1819,N_1803);
nor U2130 (N_2130,N_1998,N_1913);
and U2131 (N_2131,N_1971,N_1891);
or U2132 (N_2132,N_1948,N_1849);
nor U2133 (N_2133,N_1932,N_1987);
nand U2134 (N_2134,N_1972,N_1837);
nand U2135 (N_2135,N_1957,N_1983);
and U2136 (N_2136,N_1979,N_1886);
nor U2137 (N_2137,N_1997,N_1937);
xor U2138 (N_2138,N_1871,N_1831);
or U2139 (N_2139,N_1802,N_1923);
or U2140 (N_2140,N_1857,N_1992);
or U2141 (N_2141,N_1901,N_1964);
and U2142 (N_2142,N_1847,N_1957);
xnor U2143 (N_2143,N_1994,N_1926);
nor U2144 (N_2144,N_1906,N_1821);
nand U2145 (N_2145,N_1962,N_1850);
or U2146 (N_2146,N_1827,N_1886);
xnor U2147 (N_2147,N_1896,N_1847);
xor U2148 (N_2148,N_1975,N_1908);
nand U2149 (N_2149,N_1975,N_1902);
nor U2150 (N_2150,N_1959,N_1887);
nand U2151 (N_2151,N_1850,N_1859);
and U2152 (N_2152,N_1967,N_1942);
nand U2153 (N_2153,N_1999,N_1822);
xnor U2154 (N_2154,N_1888,N_1944);
nor U2155 (N_2155,N_1984,N_1922);
and U2156 (N_2156,N_1887,N_1860);
or U2157 (N_2157,N_1825,N_1940);
nand U2158 (N_2158,N_1838,N_1943);
xnor U2159 (N_2159,N_1891,N_1960);
or U2160 (N_2160,N_1961,N_1935);
nand U2161 (N_2161,N_1843,N_1859);
or U2162 (N_2162,N_1936,N_1866);
nand U2163 (N_2163,N_1828,N_1902);
nor U2164 (N_2164,N_1812,N_1977);
or U2165 (N_2165,N_1996,N_1994);
and U2166 (N_2166,N_1810,N_1805);
nand U2167 (N_2167,N_1890,N_1923);
nand U2168 (N_2168,N_1917,N_1977);
xor U2169 (N_2169,N_1913,N_1877);
nor U2170 (N_2170,N_1803,N_1900);
or U2171 (N_2171,N_1905,N_1910);
xor U2172 (N_2172,N_1902,N_1900);
or U2173 (N_2173,N_1991,N_1967);
or U2174 (N_2174,N_1918,N_1898);
and U2175 (N_2175,N_1871,N_1858);
nand U2176 (N_2176,N_1963,N_1875);
nor U2177 (N_2177,N_1854,N_1847);
xnor U2178 (N_2178,N_1997,N_1984);
nor U2179 (N_2179,N_1811,N_1942);
nand U2180 (N_2180,N_1849,N_1990);
xor U2181 (N_2181,N_1914,N_1972);
and U2182 (N_2182,N_1983,N_1933);
nor U2183 (N_2183,N_1937,N_1959);
and U2184 (N_2184,N_1815,N_1915);
nor U2185 (N_2185,N_1958,N_1991);
or U2186 (N_2186,N_1834,N_1822);
xor U2187 (N_2187,N_1954,N_1865);
nor U2188 (N_2188,N_1989,N_1937);
nor U2189 (N_2189,N_1946,N_1839);
xor U2190 (N_2190,N_1879,N_1833);
nand U2191 (N_2191,N_1982,N_1865);
xnor U2192 (N_2192,N_1902,N_1958);
or U2193 (N_2193,N_1804,N_1920);
or U2194 (N_2194,N_1944,N_1924);
or U2195 (N_2195,N_1800,N_1901);
and U2196 (N_2196,N_1804,N_1849);
and U2197 (N_2197,N_1893,N_1925);
and U2198 (N_2198,N_1973,N_1857);
nor U2199 (N_2199,N_1821,N_1926);
or U2200 (N_2200,N_2115,N_2171);
and U2201 (N_2201,N_2148,N_2190);
nand U2202 (N_2202,N_2129,N_2189);
nand U2203 (N_2203,N_2094,N_2144);
nand U2204 (N_2204,N_2128,N_2176);
xor U2205 (N_2205,N_2028,N_2068);
and U2206 (N_2206,N_2073,N_2136);
or U2207 (N_2207,N_2184,N_2177);
nand U2208 (N_2208,N_2080,N_2143);
and U2209 (N_2209,N_2172,N_2105);
nand U2210 (N_2210,N_2012,N_2085);
nand U2211 (N_2211,N_2159,N_2065);
or U2212 (N_2212,N_2084,N_2037);
or U2213 (N_2213,N_2179,N_2081);
nand U2214 (N_2214,N_2016,N_2147);
or U2215 (N_2215,N_2022,N_2072);
or U2216 (N_2216,N_2170,N_2041);
nand U2217 (N_2217,N_2131,N_2063);
and U2218 (N_2218,N_2157,N_2007);
or U2219 (N_2219,N_2130,N_2161);
or U2220 (N_2220,N_2062,N_2024);
nand U2221 (N_2221,N_2122,N_2111);
or U2222 (N_2222,N_2025,N_2079);
nand U2223 (N_2223,N_2142,N_2059);
or U2224 (N_2224,N_2017,N_2118);
nand U2225 (N_2225,N_2107,N_2175);
nor U2226 (N_2226,N_2164,N_2069);
and U2227 (N_2227,N_2152,N_2074);
nor U2228 (N_2228,N_2027,N_2004);
nor U2229 (N_2229,N_2197,N_2087);
or U2230 (N_2230,N_2139,N_2061);
and U2231 (N_2231,N_2067,N_2088);
xor U2232 (N_2232,N_2199,N_2106);
nor U2233 (N_2233,N_2052,N_2011);
or U2234 (N_2234,N_2009,N_2021);
nor U2235 (N_2235,N_2098,N_2187);
or U2236 (N_2236,N_2082,N_2178);
and U2237 (N_2237,N_2047,N_2035);
nand U2238 (N_2238,N_2043,N_2174);
nor U2239 (N_2239,N_2093,N_2051);
or U2240 (N_2240,N_2154,N_2044);
and U2241 (N_2241,N_2185,N_2146);
nand U2242 (N_2242,N_2019,N_2023);
and U2243 (N_2243,N_2020,N_2173);
nand U2244 (N_2244,N_2018,N_2191);
or U2245 (N_2245,N_2076,N_2150);
xor U2246 (N_2246,N_2145,N_2137);
or U2247 (N_2247,N_2015,N_2101);
nand U2248 (N_2248,N_2169,N_2092);
nand U2249 (N_2249,N_2100,N_2158);
and U2250 (N_2250,N_2095,N_2055);
nand U2251 (N_2251,N_2029,N_2151);
and U2252 (N_2252,N_2010,N_2167);
nor U2253 (N_2253,N_2003,N_2031);
nor U2254 (N_2254,N_2075,N_2099);
xor U2255 (N_2255,N_2034,N_2060);
nor U2256 (N_2256,N_2089,N_2077);
nor U2257 (N_2257,N_2127,N_2198);
nor U2258 (N_2258,N_2156,N_2193);
nand U2259 (N_2259,N_2163,N_2186);
nor U2260 (N_2260,N_2183,N_2117);
nand U2261 (N_2261,N_2125,N_2086);
or U2262 (N_2262,N_2194,N_2056);
nand U2263 (N_2263,N_2195,N_2053);
nand U2264 (N_2264,N_2066,N_2039);
xor U2265 (N_2265,N_2181,N_2054);
nand U2266 (N_2266,N_2132,N_2070);
and U2267 (N_2267,N_2114,N_2124);
and U2268 (N_2268,N_2149,N_2045);
and U2269 (N_2269,N_2182,N_2071);
and U2270 (N_2270,N_2155,N_2033);
nand U2271 (N_2271,N_2196,N_2097);
xnor U2272 (N_2272,N_2000,N_2102);
xnor U2273 (N_2273,N_2112,N_2001);
nor U2274 (N_2274,N_2160,N_2096);
and U2275 (N_2275,N_2110,N_2002);
or U2276 (N_2276,N_2113,N_2040);
nor U2277 (N_2277,N_2109,N_2188);
and U2278 (N_2278,N_2141,N_2083);
nor U2279 (N_2279,N_2165,N_2030);
nor U2280 (N_2280,N_2135,N_2126);
or U2281 (N_2281,N_2108,N_2032);
xnor U2282 (N_2282,N_2013,N_2046);
and U2283 (N_2283,N_2133,N_2049);
and U2284 (N_2284,N_2057,N_2121);
nor U2285 (N_2285,N_2014,N_2103);
and U2286 (N_2286,N_2134,N_2180);
nor U2287 (N_2287,N_2050,N_2153);
nor U2288 (N_2288,N_2008,N_2091);
and U2289 (N_2289,N_2120,N_2140);
nand U2290 (N_2290,N_2006,N_2192);
nor U2291 (N_2291,N_2038,N_2090);
nor U2292 (N_2292,N_2042,N_2162);
and U2293 (N_2293,N_2168,N_2026);
or U2294 (N_2294,N_2058,N_2138);
and U2295 (N_2295,N_2078,N_2005);
nand U2296 (N_2296,N_2123,N_2166);
or U2297 (N_2297,N_2119,N_2036);
xor U2298 (N_2298,N_2104,N_2048);
or U2299 (N_2299,N_2116,N_2064);
nor U2300 (N_2300,N_2030,N_2010);
or U2301 (N_2301,N_2166,N_2036);
nand U2302 (N_2302,N_2061,N_2056);
nand U2303 (N_2303,N_2160,N_2063);
or U2304 (N_2304,N_2102,N_2113);
nand U2305 (N_2305,N_2013,N_2102);
and U2306 (N_2306,N_2110,N_2029);
xor U2307 (N_2307,N_2087,N_2074);
nor U2308 (N_2308,N_2150,N_2120);
nand U2309 (N_2309,N_2022,N_2177);
and U2310 (N_2310,N_2176,N_2019);
nand U2311 (N_2311,N_2115,N_2125);
nand U2312 (N_2312,N_2174,N_2135);
nor U2313 (N_2313,N_2148,N_2053);
nand U2314 (N_2314,N_2176,N_2038);
nor U2315 (N_2315,N_2087,N_2184);
nor U2316 (N_2316,N_2099,N_2091);
and U2317 (N_2317,N_2046,N_2083);
or U2318 (N_2318,N_2110,N_2018);
xnor U2319 (N_2319,N_2028,N_2063);
nor U2320 (N_2320,N_2011,N_2191);
nand U2321 (N_2321,N_2005,N_2023);
xnor U2322 (N_2322,N_2191,N_2172);
xor U2323 (N_2323,N_2091,N_2053);
nor U2324 (N_2324,N_2109,N_2063);
or U2325 (N_2325,N_2164,N_2151);
and U2326 (N_2326,N_2041,N_2085);
or U2327 (N_2327,N_2126,N_2141);
or U2328 (N_2328,N_2071,N_2140);
nand U2329 (N_2329,N_2184,N_2195);
nor U2330 (N_2330,N_2001,N_2133);
or U2331 (N_2331,N_2175,N_2172);
and U2332 (N_2332,N_2187,N_2143);
nand U2333 (N_2333,N_2157,N_2096);
nand U2334 (N_2334,N_2099,N_2019);
or U2335 (N_2335,N_2140,N_2176);
and U2336 (N_2336,N_2087,N_2013);
and U2337 (N_2337,N_2025,N_2067);
nand U2338 (N_2338,N_2174,N_2199);
and U2339 (N_2339,N_2170,N_2175);
nand U2340 (N_2340,N_2016,N_2021);
nand U2341 (N_2341,N_2190,N_2115);
or U2342 (N_2342,N_2075,N_2027);
and U2343 (N_2343,N_2024,N_2081);
xnor U2344 (N_2344,N_2063,N_2172);
nand U2345 (N_2345,N_2133,N_2005);
nor U2346 (N_2346,N_2054,N_2057);
and U2347 (N_2347,N_2105,N_2129);
nand U2348 (N_2348,N_2099,N_2059);
xor U2349 (N_2349,N_2067,N_2022);
and U2350 (N_2350,N_2165,N_2162);
and U2351 (N_2351,N_2037,N_2199);
and U2352 (N_2352,N_2054,N_2096);
and U2353 (N_2353,N_2125,N_2024);
nand U2354 (N_2354,N_2044,N_2127);
nand U2355 (N_2355,N_2096,N_2004);
nor U2356 (N_2356,N_2056,N_2116);
and U2357 (N_2357,N_2067,N_2008);
nor U2358 (N_2358,N_2194,N_2068);
nor U2359 (N_2359,N_2022,N_2172);
nand U2360 (N_2360,N_2174,N_2002);
nor U2361 (N_2361,N_2169,N_2163);
nand U2362 (N_2362,N_2121,N_2124);
or U2363 (N_2363,N_2013,N_2092);
nor U2364 (N_2364,N_2028,N_2001);
nor U2365 (N_2365,N_2057,N_2098);
xnor U2366 (N_2366,N_2091,N_2197);
nand U2367 (N_2367,N_2092,N_2123);
nand U2368 (N_2368,N_2069,N_2044);
xor U2369 (N_2369,N_2141,N_2179);
or U2370 (N_2370,N_2085,N_2082);
and U2371 (N_2371,N_2154,N_2185);
or U2372 (N_2372,N_2094,N_2079);
or U2373 (N_2373,N_2127,N_2023);
and U2374 (N_2374,N_2178,N_2028);
xor U2375 (N_2375,N_2049,N_2045);
or U2376 (N_2376,N_2082,N_2142);
and U2377 (N_2377,N_2122,N_2057);
or U2378 (N_2378,N_2018,N_2082);
or U2379 (N_2379,N_2083,N_2137);
nand U2380 (N_2380,N_2026,N_2126);
nor U2381 (N_2381,N_2080,N_2057);
nand U2382 (N_2382,N_2001,N_2010);
or U2383 (N_2383,N_2062,N_2115);
xnor U2384 (N_2384,N_2003,N_2155);
xor U2385 (N_2385,N_2149,N_2198);
or U2386 (N_2386,N_2197,N_2159);
or U2387 (N_2387,N_2031,N_2041);
and U2388 (N_2388,N_2124,N_2108);
nor U2389 (N_2389,N_2142,N_2174);
nor U2390 (N_2390,N_2076,N_2160);
nor U2391 (N_2391,N_2094,N_2183);
nand U2392 (N_2392,N_2177,N_2193);
and U2393 (N_2393,N_2053,N_2038);
nor U2394 (N_2394,N_2179,N_2084);
nand U2395 (N_2395,N_2129,N_2120);
and U2396 (N_2396,N_2142,N_2136);
nand U2397 (N_2397,N_2102,N_2016);
nor U2398 (N_2398,N_2176,N_2136);
or U2399 (N_2399,N_2092,N_2096);
nand U2400 (N_2400,N_2388,N_2296);
or U2401 (N_2401,N_2295,N_2214);
nor U2402 (N_2402,N_2323,N_2217);
nand U2403 (N_2403,N_2391,N_2208);
or U2404 (N_2404,N_2396,N_2286);
xnor U2405 (N_2405,N_2368,N_2205);
nand U2406 (N_2406,N_2316,N_2293);
xnor U2407 (N_2407,N_2276,N_2247);
and U2408 (N_2408,N_2256,N_2399);
and U2409 (N_2409,N_2343,N_2290);
nor U2410 (N_2410,N_2223,N_2375);
or U2411 (N_2411,N_2255,N_2338);
or U2412 (N_2412,N_2230,N_2377);
or U2413 (N_2413,N_2303,N_2280);
nor U2414 (N_2414,N_2392,N_2267);
or U2415 (N_2415,N_2398,N_2304);
or U2416 (N_2416,N_2306,N_2355);
and U2417 (N_2417,N_2271,N_2327);
and U2418 (N_2418,N_2237,N_2227);
or U2419 (N_2419,N_2228,N_2213);
nor U2420 (N_2420,N_2333,N_2281);
or U2421 (N_2421,N_2261,N_2337);
xor U2422 (N_2422,N_2229,N_2361);
xor U2423 (N_2423,N_2331,N_2283);
nor U2424 (N_2424,N_2352,N_2294);
nor U2425 (N_2425,N_2339,N_2394);
or U2426 (N_2426,N_2358,N_2359);
nand U2427 (N_2427,N_2373,N_2322);
and U2428 (N_2428,N_2384,N_2330);
and U2429 (N_2429,N_2221,N_2200);
or U2430 (N_2430,N_2393,N_2360);
xor U2431 (N_2431,N_2204,N_2285);
or U2432 (N_2432,N_2313,N_2209);
nand U2433 (N_2433,N_2297,N_2272);
and U2434 (N_2434,N_2279,N_2312);
or U2435 (N_2435,N_2282,N_2334);
xnor U2436 (N_2436,N_2242,N_2284);
nand U2437 (N_2437,N_2351,N_2371);
nand U2438 (N_2438,N_2252,N_2219);
and U2439 (N_2439,N_2349,N_2348);
and U2440 (N_2440,N_2385,N_2268);
nand U2441 (N_2441,N_2344,N_2326);
xnor U2442 (N_2442,N_2357,N_2215);
or U2443 (N_2443,N_2259,N_2300);
nor U2444 (N_2444,N_2234,N_2308);
and U2445 (N_2445,N_2389,N_2233);
and U2446 (N_2446,N_2329,N_2305);
and U2447 (N_2447,N_2321,N_2243);
and U2448 (N_2448,N_2369,N_2277);
or U2449 (N_2449,N_2235,N_2244);
or U2450 (N_2450,N_2395,N_2264);
or U2451 (N_2451,N_2382,N_2380);
and U2452 (N_2452,N_2232,N_2202);
nor U2453 (N_2453,N_2212,N_2315);
nor U2454 (N_2454,N_2250,N_2301);
nand U2455 (N_2455,N_2288,N_2206);
nand U2456 (N_2456,N_2291,N_2220);
nand U2457 (N_2457,N_2275,N_2254);
or U2458 (N_2458,N_2287,N_2336);
or U2459 (N_2459,N_2211,N_2363);
or U2460 (N_2460,N_2367,N_2278);
and U2461 (N_2461,N_2362,N_2332);
xnor U2462 (N_2462,N_2347,N_2241);
nand U2463 (N_2463,N_2201,N_2397);
or U2464 (N_2464,N_2390,N_2335);
nor U2465 (N_2465,N_2299,N_2249);
and U2466 (N_2466,N_2263,N_2222);
and U2467 (N_2467,N_2274,N_2381);
nand U2468 (N_2468,N_2314,N_2273);
or U2469 (N_2469,N_2342,N_2302);
or U2470 (N_2470,N_2386,N_2262);
or U2471 (N_2471,N_2246,N_2311);
or U2472 (N_2472,N_2245,N_2370);
nor U2473 (N_2473,N_2260,N_2318);
or U2474 (N_2474,N_2238,N_2251);
and U2475 (N_2475,N_2226,N_2346);
nand U2476 (N_2476,N_2340,N_2218);
and U2477 (N_2477,N_2270,N_2258);
xor U2478 (N_2478,N_2265,N_2269);
or U2479 (N_2479,N_2248,N_2203);
nand U2480 (N_2480,N_2225,N_2231);
nand U2481 (N_2481,N_2345,N_2257);
xor U2482 (N_2482,N_2309,N_2210);
or U2483 (N_2483,N_2207,N_2240);
or U2484 (N_2484,N_2324,N_2378);
or U2485 (N_2485,N_2292,N_2350);
nor U2486 (N_2486,N_2310,N_2239);
and U2487 (N_2487,N_2365,N_2320);
or U2488 (N_2488,N_2383,N_2376);
or U2489 (N_2489,N_2364,N_2353);
and U2490 (N_2490,N_2307,N_2356);
xor U2491 (N_2491,N_2289,N_2298);
or U2492 (N_2492,N_2372,N_2354);
or U2493 (N_2493,N_2317,N_2216);
nor U2494 (N_2494,N_2379,N_2236);
and U2495 (N_2495,N_2328,N_2341);
or U2496 (N_2496,N_2325,N_2319);
and U2497 (N_2497,N_2253,N_2387);
xor U2498 (N_2498,N_2374,N_2366);
nand U2499 (N_2499,N_2224,N_2266);
nor U2500 (N_2500,N_2367,N_2222);
or U2501 (N_2501,N_2204,N_2311);
nand U2502 (N_2502,N_2305,N_2294);
nand U2503 (N_2503,N_2338,N_2252);
nor U2504 (N_2504,N_2396,N_2331);
and U2505 (N_2505,N_2382,N_2372);
or U2506 (N_2506,N_2210,N_2248);
or U2507 (N_2507,N_2242,N_2301);
or U2508 (N_2508,N_2376,N_2308);
nand U2509 (N_2509,N_2324,N_2340);
nand U2510 (N_2510,N_2336,N_2349);
nor U2511 (N_2511,N_2286,N_2248);
and U2512 (N_2512,N_2252,N_2352);
nor U2513 (N_2513,N_2323,N_2333);
nand U2514 (N_2514,N_2249,N_2241);
nand U2515 (N_2515,N_2365,N_2364);
or U2516 (N_2516,N_2324,N_2342);
and U2517 (N_2517,N_2237,N_2345);
nand U2518 (N_2518,N_2333,N_2363);
and U2519 (N_2519,N_2305,N_2288);
and U2520 (N_2520,N_2255,N_2316);
nand U2521 (N_2521,N_2314,N_2256);
nand U2522 (N_2522,N_2252,N_2282);
nor U2523 (N_2523,N_2277,N_2395);
nor U2524 (N_2524,N_2269,N_2251);
nand U2525 (N_2525,N_2221,N_2305);
nand U2526 (N_2526,N_2351,N_2202);
or U2527 (N_2527,N_2369,N_2386);
nor U2528 (N_2528,N_2308,N_2322);
and U2529 (N_2529,N_2304,N_2331);
xor U2530 (N_2530,N_2357,N_2231);
nor U2531 (N_2531,N_2324,N_2362);
nor U2532 (N_2532,N_2389,N_2351);
and U2533 (N_2533,N_2215,N_2211);
nand U2534 (N_2534,N_2283,N_2299);
nor U2535 (N_2535,N_2244,N_2207);
nand U2536 (N_2536,N_2386,N_2266);
and U2537 (N_2537,N_2340,N_2345);
nor U2538 (N_2538,N_2226,N_2219);
nand U2539 (N_2539,N_2295,N_2274);
or U2540 (N_2540,N_2206,N_2330);
or U2541 (N_2541,N_2248,N_2307);
or U2542 (N_2542,N_2359,N_2298);
xnor U2543 (N_2543,N_2291,N_2380);
xnor U2544 (N_2544,N_2223,N_2346);
and U2545 (N_2545,N_2335,N_2250);
or U2546 (N_2546,N_2375,N_2345);
xor U2547 (N_2547,N_2390,N_2233);
and U2548 (N_2548,N_2372,N_2344);
nor U2549 (N_2549,N_2302,N_2277);
nor U2550 (N_2550,N_2371,N_2385);
nand U2551 (N_2551,N_2297,N_2316);
nand U2552 (N_2552,N_2383,N_2327);
xnor U2553 (N_2553,N_2301,N_2385);
and U2554 (N_2554,N_2356,N_2234);
or U2555 (N_2555,N_2389,N_2305);
and U2556 (N_2556,N_2298,N_2369);
nand U2557 (N_2557,N_2225,N_2362);
or U2558 (N_2558,N_2394,N_2281);
nor U2559 (N_2559,N_2389,N_2227);
or U2560 (N_2560,N_2352,N_2377);
nand U2561 (N_2561,N_2278,N_2384);
and U2562 (N_2562,N_2281,N_2384);
or U2563 (N_2563,N_2270,N_2211);
or U2564 (N_2564,N_2358,N_2242);
or U2565 (N_2565,N_2358,N_2208);
nor U2566 (N_2566,N_2379,N_2296);
nor U2567 (N_2567,N_2240,N_2203);
and U2568 (N_2568,N_2285,N_2290);
nor U2569 (N_2569,N_2243,N_2283);
xor U2570 (N_2570,N_2273,N_2305);
nor U2571 (N_2571,N_2368,N_2245);
nor U2572 (N_2572,N_2227,N_2280);
or U2573 (N_2573,N_2208,N_2377);
nor U2574 (N_2574,N_2399,N_2293);
or U2575 (N_2575,N_2239,N_2252);
or U2576 (N_2576,N_2391,N_2374);
nor U2577 (N_2577,N_2272,N_2363);
or U2578 (N_2578,N_2250,N_2297);
nand U2579 (N_2579,N_2240,N_2331);
and U2580 (N_2580,N_2367,N_2387);
or U2581 (N_2581,N_2254,N_2330);
and U2582 (N_2582,N_2211,N_2319);
and U2583 (N_2583,N_2257,N_2300);
and U2584 (N_2584,N_2336,N_2243);
xnor U2585 (N_2585,N_2381,N_2360);
or U2586 (N_2586,N_2247,N_2395);
nor U2587 (N_2587,N_2302,N_2373);
and U2588 (N_2588,N_2397,N_2393);
or U2589 (N_2589,N_2341,N_2348);
or U2590 (N_2590,N_2237,N_2201);
or U2591 (N_2591,N_2391,N_2315);
nor U2592 (N_2592,N_2387,N_2241);
nand U2593 (N_2593,N_2320,N_2301);
and U2594 (N_2594,N_2311,N_2217);
nor U2595 (N_2595,N_2296,N_2390);
or U2596 (N_2596,N_2321,N_2275);
xor U2597 (N_2597,N_2260,N_2306);
xor U2598 (N_2598,N_2364,N_2324);
nor U2599 (N_2599,N_2288,N_2281);
and U2600 (N_2600,N_2549,N_2461);
nor U2601 (N_2601,N_2544,N_2522);
xor U2602 (N_2602,N_2473,N_2494);
or U2603 (N_2603,N_2576,N_2593);
xnor U2604 (N_2604,N_2451,N_2442);
nor U2605 (N_2605,N_2424,N_2571);
and U2606 (N_2606,N_2495,N_2501);
or U2607 (N_2607,N_2467,N_2508);
nand U2608 (N_2608,N_2539,N_2560);
or U2609 (N_2609,N_2546,N_2489);
xnor U2610 (N_2610,N_2587,N_2496);
nand U2611 (N_2611,N_2579,N_2499);
nand U2612 (N_2612,N_2476,N_2582);
and U2613 (N_2613,N_2401,N_2464);
and U2614 (N_2614,N_2471,N_2525);
nand U2615 (N_2615,N_2446,N_2417);
nand U2616 (N_2616,N_2553,N_2488);
nor U2617 (N_2617,N_2574,N_2416);
and U2618 (N_2618,N_2521,N_2443);
or U2619 (N_2619,N_2447,N_2459);
nand U2620 (N_2620,N_2487,N_2518);
nand U2621 (N_2621,N_2482,N_2445);
nor U2622 (N_2622,N_2523,N_2430);
nand U2623 (N_2623,N_2586,N_2463);
or U2624 (N_2624,N_2529,N_2510);
nand U2625 (N_2625,N_2419,N_2456);
nor U2626 (N_2626,N_2462,N_2444);
or U2627 (N_2627,N_2583,N_2598);
nor U2628 (N_2628,N_2502,N_2441);
and U2629 (N_2629,N_2493,N_2405);
xor U2630 (N_2630,N_2517,N_2475);
xnor U2631 (N_2631,N_2584,N_2513);
nand U2632 (N_2632,N_2474,N_2407);
nand U2633 (N_2633,N_2599,N_2557);
nor U2634 (N_2634,N_2519,N_2434);
nand U2635 (N_2635,N_2590,N_2594);
and U2636 (N_2636,N_2437,N_2452);
and U2637 (N_2637,N_2588,N_2409);
nand U2638 (N_2638,N_2477,N_2575);
or U2639 (N_2639,N_2486,N_2428);
xor U2640 (N_2640,N_2431,N_2478);
nor U2641 (N_2641,N_2465,N_2535);
and U2642 (N_2642,N_2559,N_2433);
and U2643 (N_2643,N_2564,N_2570);
and U2644 (N_2644,N_2404,N_2460);
and U2645 (N_2645,N_2505,N_2506);
nor U2646 (N_2646,N_2497,N_2568);
or U2647 (N_2647,N_2412,N_2562);
and U2648 (N_2648,N_2527,N_2438);
xor U2649 (N_2649,N_2455,N_2402);
nand U2650 (N_2650,N_2516,N_2453);
or U2651 (N_2651,N_2484,N_2410);
or U2652 (N_2652,N_2439,N_2545);
nand U2653 (N_2653,N_2472,N_2418);
nand U2654 (N_2654,N_2569,N_2563);
nor U2655 (N_2655,N_2403,N_2432);
nand U2656 (N_2656,N_2534,N_2481);
or U2657 (N_2657,N_2556,N_2512);
nand U2658 (N_2658,N_2425,N_2573);
and U2659 (N_2659,N_2555,N_2585);
nor U2660 (N_2660,N_2581,N_2507);
xnor U2661 (N_2661,N_2530,N_2547);
nand U2662 (N_2662,N_2448,N_2427);
nand U2663 (N_2663,N_2578,N_2440);
nand U2664 (N_2664,N_2454,N_2526);
nand U2665 (N_2665,N_2408,N_2426);
xor U2666 (N_2666,N_2551,N_2531);
nand U2667 (N_2667,N_2491,N_2595);
nand U2668 (N_2668,N_2550,N_2542);
and U2669 (N_2669,N_2537,N_2483);
nand U2670 (N_2670,N_2580,N_2450);
nor U2671 (N_2671,N_2498,N_2515);
or U2672 (N_2672,N_2492,N_2420);
or U2673 (N_2673,N_2533,N_2415);
and U2674 (N_2674,N_2532,N_2567);
nand U2675 (N_2675,N_2485,N_2457);
xor U2676 (N_2676,N_2514,N_2435);
and U2677 (N_2677,N_2591,N_2466);
or U2678 (N_2678,N_2429,N_2421);
nor U2679 (N_2679,N_2423,N_2436);
nand U2680 (N_2680,N_2414,N_2528);
or U2681 (N_2681,N_2538,N_2552);
nor U2682 (N_2682,N_2589,N_2548);
nand U2683 (N_2683,N_2558,N_2449);
and U2684 (N_2684,N_2503,N_2596);
xnor U2685 (N_2685,N_2572,N_2480);
nor U2686 (N_2686,N_2561,N_2504);
and U2687 (N_2687,N_2411,N_2566);
nand U2688 (N_2688,N_2406,N_2470);
nand U2689 (N_2689,N_2422,N_2400);
or U2690 (N_2690,N_2500,N_2458);
nand U2691 (N_2691,N_2536,N_2511);
or U2692 (N_2692,N_2541,N_2469);
or U2693 (N_2693,N_2524,N_2597);
and U2694 (N_2694,N_2543,N_2479);
or U2695 (N_2695,N_2413,N_2577);
nand U2696 (N_2696,N_2468,N_2565);
nand U2697 (N_2697,N_2490,N_2520);
or U2698 (N_2698,N_2554,N_2509);
xnor U2699 (N_2699,N_2592,N_2540);
or U2700 (N_2700,N_2439,N_2407);
nor U2701 (N_2701,N_2509,N_2543);
or U2702 (N_2702,N_2566,N_2450);
or U2703 (N_2703,N_2578,N_2416);
or U2704 (N_2704,N_2596,N_2417);
nand U2705 (N_2705,N_2556,N_2475);
nand U2706 (N_2706,N_2568,N_2489);
and U2707 (N_2707,N_2468,N_2596);
nand U2708 (N_2708,N_2408,N_2570);
and U2709 (N_2709,N_2578,N_2552);
and U2710 (N_2710,N_2571,N_2553);
nand U2711 (N_2711,N_2476,N_2414);
or U2712 (N_2712,N_2588,N_2571);
xor U2713 (N_2713,N_2452,N_2459);
or U2714 (N_2714,N_2419,N_2479);
or U2715 (N_2715,N_2547,N_2538);
or U2716 (N_2716,N_2522,N_2514);
and U2717 (N_2717,N_2503,N_2529);
nor U2718 (N_2718,N_2549,N_2450);
or U2719 (N_2719,N_2573,N_2441);
nand U2720 (N_2720,N_2536,N_2417);
xnor U2721 (N_2721,N_2497,N_2534);
xor U2722 (N_2722,N_2528,N_2454);
and U2723 (N_2723,N_2574,N_2478);
nor U2724 (N_2724,N_2435,N_2480);
nor U2725 (N_2725,N_2417,N_2509);
and U2726 (N_2726,N_2450,N_2475);
nor U2727 (N_2727,N_2451,N_2566);
nand U2728 (N_2728,N_2525,N_2540);
nand U2729 (N_2729,N_2585,N_2552);
nor U2730 (N_2730,N_2599,N_2598);
and U2731 (N_2731,N_2455,N_2438);
xor U2732 (N_2732,N_2507,N_2440);
nand U2733 (N_2733,N_2591,N_2518);
nor U2734 (N_2734,N_2537,N_2497);
xnor U2735 (N_2735,N_2597,N_2476);
xor U2736 (N_2736,N_2596,N_2550);
and U2737 (N_2737,N_2481,N_2556);
or U2738 (N_2738,N_2436,N_2567);
xnor U2739 (N_2739,N_2444,N_2524);
xor U2740 (N_2740,N_2534,N_2595);
or U2741 (N_2741,N_2431,N_2575);
nand U2742 (N_2742,N_2440,N_2537);
or U2743 (N_2743,N_2418,N_2441);
or U2744 (N_2744,N_2489,N_2514);
nor U2745 (N_2745,N_2556,N_2412);
and U2746 (N_2746,N_2574,N_2571);
nand U2747 (N_2747,N_2466,N_2442);
or U2748 (N_2748,N_2592,N_2517);
and U2749 (N_2749,N_2523,N_2434);
or U2750 (N_2750,N_2529,N_2536);
and U2751 (N_2751,N_2420,N_2536);
nand U2752 (N_2752,N_2403,N_2477);
nand U2753 (N_2753,N_2479,N_2557);
nand U2754 (N_2754,N_2497,N_2456);
and U2755 (N_2755,N_2454,N_2543);
and U2756 (N_2756,N_2560,N_2563);
nand U2757 (N_2757,N_2442,N_2549);
or U2758 (N_2758,N_2585,N_2414);
and U2759 (N_2759,N_2469,N_2461);
nand U2760 (N_2760,N_2421,N_2414);
nand U2761 (N_2761,N_2570,N_2454);
nand U2762 (N_2762,N_2582,N_2448);
nor U2763 (N_2763,N_2433,N_2461);
nand U2764 (N_2764,N_2457,N_2510);
nor U2765 (N_2765,N_2599,N_2470);
or U2766 (N_2766,N_2423,N_2549);
and U2767 (N_2767,N_2504,N_2583);
and U2768 (N_2768,N_2414,N_2595);
nor U2769 (N_2769,N_2594,N_2491);
or U2770 (N_2770,N_2446,N_2406);
nor U2771 (N_2771,N_2476,N_2568);
nand U2772 (N_2772,N_2558,N_2456);
nand U2773 (N_2773,N_2481,N_2507);
and U2774 (N_2774,N_2408,N_2482);
nor U2775 (N_2775,N_2586,N_2410);
nor U2776 (N_2776,N_2479,N_2416);
nor U2777 (N_2777,N_2407,N_2507);
or U2778 (N_2778,N_2446,N_2405);
and U2779 (N_2779,N_2547,N_2469);
nor U2780 (N_2780,N_2469,N_2453);
or U2781 (N_2781,N_2589,N_2456);
nand U2782 (N_2782,N_2549,N_2493);
or U2783 (N_2783,N_2566,N_2534);
nand U2784 (N_2784,N_2428,N_2484);
or U2785 (N_2785,N_2599,N_2430);
nor U2786 (N_2786,N_2509,N_2580);
or U2787 (N_2787,N_2597,N_2548);
nand U2788 (N_2788,N_2473,N_2491);
nand U2789 (N_2789,N_2496,N_2422);
nor U2790 (N_2790,N_2568,N_2406);
nor U2791 (N_2791,N_2585,N_2500);
and U2792 (N_2792,N_2470,N_2565);
nor U2793 (N_2793,N_2426,N_2528);
xor U2794 (N_2794,N_2442,N_2441);
nor U2795 (N_2795,N_2469,N_2540);
nand U2796 (N_2796,N_2480,N_2519);
xnor U2797 (N_2797,N_2413,N_2557);
xnor U2798 (N_2798,N_2488,N_2484);
nor U2799 (N_2799,N_2429,N_2459);
or U2800 (N_2800,N_2775,N_2653);
nor U2801 (N_2801,N_2747,N_2708);
and U2802 (N_2802,N_2763,N_2724);
nor U2803 (N_2803,N_2664,N_2673);
nor U2804 (N_2804,N_2699,N_2760);
or U2805 (N_2805,N_2703,N_2646);
nand U2806 (N_2806,N_2726,N_2773);
and U2807 (N_2807,N_2737,N_2752);
nor U2808 (N_2808,N_2636,N_2743);
or U2809 (N_2809,N_2615,N_2767);
nor U2810 (N_2810,N_2797,N_2643);
nand U2811 (N_2811,N_2634,N_2793);
nor U2812 (N_2812,N_2651,N_2672);
nor U2813 (N_2813,N_2740,N_2776);
nor U2814 (N_2814,N_2621,N_2670);
and U2815 (N_2815,N_2676,N_2766);
and U2816 (N_2816,N_2730,N_2603);
nor U2817 (N_2817,N_2770,N_2729);
and U2818 (N_2818,N_2781,N_2756);
and U2819 (N_2819,N_2602,N_2750);
and U2820 (N_2820,N_2655,N_2614);
nor U2821 (N_2821,N_2665,N_2685);
nand U2822 (N_2822,N_2725,N_2748);
nor U2823 (N_2823,N_2642,N_2698);
or U2824 (N_2824,N_2680,N_2610);
nor U2825 (N_2825,N_2689,N_2608);
nand U2826 (N_2826,N_2732,N_2789);
nand U2827 (N_2827,N_2735,N_2717);
nand U2828 (N_2828,N_2690,N_2624);
and U2829 (N_2829,N_2761,N_2728);
nand U2830 (N_2830,N_2707,N_2683);
nor U2831 (N_2831,N_2782,N_2710);
nor U2832 (N_2832,N_2607,N_2609);
or U2833 (N_2833,N_2669,N_2681);
or U2834 (N_2834,N_2796,N_2674);
xor U2835 (N_2835,N_2757,N_2704);
nor U2836 (N_2836,N_2696,N_2666);
nand U2837 (N_2837,N_2633,N_2627);
and U2838 (N_2838,N_2723,N_2618);
nand U2839 (N_2839,N_2600,N_2650);
nor U2840 (N_2840,N_2783,N_2749);
nor U2841 (N_2841,N_2733,N_2679);
nor U2842 (N_2842,N_2738,N_2617);
or U2843 (N_2843,N_2641,N_2758);
and U2844 (N_2844,N_2741,N_2660);
and U2845 (N_2845,N_2755,N_2606);
or U2846 (N_2846,N_2658,N_2754);
or U2847 (N_2847,N_2739,N_2788);
nand U2848 (N_2848,N_2719,N_2709);
or U2849 (N_2849,N_2605,N_2632);
nor U2850 (N_2850,N_2791,N_2677);
xor U2851 (N_2851,N_2722,N_2716);
xor U2852 (N_2852,N_2684,N_2645);
nand U2853 (N_2853,N_2718,N_2780);
or U2854 (N_2854,N_2695,N_2612);
and U2855 (N_2855,N_2713,N_2746);
nand U2856 (N_2856,N_2771,N_2795);
nor U2857 (N_2857,N_2769,N_2668);
nand U2858 (N_2858,N_2778,N_2619);
xor U2859 (N_2859,N_2692,N_2630);
nor U2860 (N_2860,N_2711,N_2639);
and U2861 (N_2861,N_2714,N_2628);
or U2862 (N_2862,N_2626,N_2648);
nor U2863 (N_2863,N_2623,N_2790);
nor U2864 (N_2864,N_2687,N_2667);
and U2865 (N_2865,N_2745,N_2662);
xnor U2866 (N_2866,N_2720,N_2691);
nor U2867 (N_2867,N_2682,N_2694);
or U2868 (N_2868,N_2751,N_2649);
or U2869 (N_2869,N_2647,N_2787);
nor U2870 (N_2870,N_2652,N_2765);
and U2871 (N_2871,N_2635,N_2779);
or U2872 (N_2872,N_2742,N_2759);
xor U2873 (N_2873,N_2762,N_2753);
nand U2874 (N_2874,N_2727,N_2622);
nor U2875 (N_2875,N_2659,N_2798);
nor U2876 (N_2876,N_2774,N_2706);
nor U2877 (N_2877,N_2705,N_2712);
or U2878 (N_2878,N_2701,N_2693);
nor U2879 (N_2879,N_2637,N_2764);
nor U2880 (N_2880,N_2772,N_2736);
nor U2881 (N_2881,N_2785,N_2768);
xor U2882 (N_2882,N_2663,N_2616);
nand U2883 (N_2883,N_2625,N_2644);
and U2884 (N_2884,N_2799,N_2792);
nor U2885 (N_2885,N_2744,N_2784);
nand U2886 (N_2886,N_2629,N_2601);
or U2887 (N_2887,N_2734,N_2777);
or U2888 (N_2888,N_2638,N_2611);
or U2889 (N_2889,N_2671,N_2794);
and U2890 (N_2890,N_2700,N_2697);
nor U2891 (N_2891,N_2654,N_2721);
nand U2892 (N_2892,N_2786,N_2678);
and U2893 (N_2893,N_2620,N_2686);
xor U2894 (N_2894,N_2657,N_2640);
nor U2895 (N_2895,N_2604,N_2656);
and U2896 (N_2896,N_2661,N_2702);
nor U2897 (N_2897,N_2675,N_2613);
xor U2898 (N_2898,N_2688,N_2631);
and U2899 (N_2899,N_2731,N_2715);
xor U2900 (N_2900,N_2683,N_2637);
and U2901 (N_2901,N_2668,N_2609);
nor U2902 (N_2902,N_2620,N_2609);
nand U2903 (N_2903,N_2699,N_2794);
and U2904 (N_2904,N_2794,N_2775);
xor U2905 (N_2905,N_2716,N_2766);
and U2906 (N_2906,N_2685,N_2799);
nand U2907 (N_2907,N_2789,N_2666);
nand U2908 (N_2908,N_2773,N_2660);
and U2909 (N_2909,N_2600,N_2617);
and U2910 (N_2910,N_2681,N_2648);
nor U2911 (N_2911,N_2659,N_2663);
nor U2912 (N_2912,N_2766,N_2669);
nand U2913 (N_2913,N_2775,N_2777);
nor U2914 (N_2914,N_2697,N_2642);
and U2915 (N_2915,N_2799,N_2724);
and U2916 (N_2916,N_2623,N_2799);
nor U2917 (N_2917,N_2748,N_2641);
nand U2918 (N_2918,N_2722,N_2715);
and U2919 (N_2919,N_2697,N_2618);
and U2920 (N_2920,N_2603,N_2607);
or U2921 (N_2921,N_2690,N_2646);
or U2922 (N_2922,N_2696,N_2691);
nor U2923 (N_2923,N_2755,N_2699);
nor U2924 (N_2924,N_2622,N_2686);
nor U2925 (N_2925,N_2693,N_2790);
nor U2926 (N_2926,N_2662,N_2666);
and U2927 (N_2927,N_2708,N_2794);
xnor U2928 (N_2928,N_2799,N_2768);
or U2929 (N_2929,N_2780,N_2771);
nand U2930 (N_2930,N_2701,N_2799);
nor U2931 (N_2931,N_2645,N_2738);
or U2932 (N_2932,N_2712,N_2722);
and U2933 (N_2933,N_2755,N_2731);
nor U2934 (N_2934,N_2752,N_2712);
or U2935 (N_2935,N_2706,N_2703);
or U2936 (N_2936,N_2758,N_2625);
nand U2937 (N_2937,N_2728,N_2704);
nor U2938 (N_2938,N_2670,N_2693);
or U2939 (N_2939,N_2688,N_2732);
nand U2940 (N_2940,N_2634,N_2623);
or U2941 (N_2941,N_2799,N_2720);
or U2942 (N_2942,N_2645,N_2663);
nand U2943 (N_2943,N_2735,N_2701);
and U2944 (N_2944,N_2795,N_2735);
xnor U2945 (N_2945,N_2654,N_2642);
nand U2946 (N_2946,N_2752,N_2649);
nor U2947 (N_2947,N_2698,N_2771);
nor U2948 (N_2948,N_2701,N_2761);
xor U2949 (N_2949,N_2673,N_2689);
or U2950 (N_2950,N_2781,N_2614);
xor U2951 (N_2951,N_2729,N_2668);
and U2952 (N_2952,N_2720,N_2778);
nor U2953 (N_2953,N_2622,N_2710);
or U2954 (N_2954,N_2795,N_2648);
and U2955 (N_2955,N_2688,N_2621);
xnor U2956 (N_2956,N_2608,N_2659);
nand U2957 (N_2957,N_2673,N_2654);
nand U2958 (N_2958,N_2746,N_2653);
or U2959 (N_2959,N_2625,N_2662);
and U2960 (N_2960,N_2778,N_2623);
and U2961 (N_2961,N_2779,N_2655);
xor U2962 (N_2962,N_2603,N_2753);
and U2963 (N_2963,N_2722,N_2797);
xor U2964 (N_2964,N_2629,N_2787);
xnor U2965 (N_2965,N_2646,N_2727);
or U2966 (N_2966,N_2768,N_2788);
or U2967 (N_2967,N_2650,N_2792);
or U2968 (N_2968,N_2668,N_2636);
nor U2969 (N_2969,N_2795,N_2794);
nor U2970 (N_2970,N_2760,N_2713);
or U2971 (N_2971,N_2753,N_2715);
nor U2972 (N_2972,N_2629,N_2765);
or U2973 (N_2973,N_2642,N_2622);
nand U2974 (N_2974,N_2707,N_2652);
nor U2975 (N_2975,N_2744,N_2691);
nor U2976 (N_2976,N_2743,N_2756);
or U2977 (N_2977,N_2677,N_2691);
nand U2978 (N_2978,N_2781,N_2752);
xor U2979 (N_2979,N_2784,N_2759);
and U2980 (N_2980,N_2789,N_2730);
nand U2981 (N_2981,N_2685,N_2676);
nor U2982 (N_2982,N_2656,N_2706);
nand U2983 (N_2983,N_2631,N_2725);
nor U2984 (N_2984,N_2723,N_2710);
or U2985 (N_2985,N_2647,N_2618);
nor U2986 (N_2986,N_2613,N_2757);
nand U2987 (N_2987,N_2732,N_2667);
nor U2988 (N_2988,N_2792,N_2798);
nand U2989 (N_2989,N_2625,N_2667);
or U2990 (N_2990,N_2786,N_2681);
nand U2991 (N_2991,N_2763,N_2707);
and U2992 (N_2992,N_2610,N_2688);
and U2993 (N_2993,N_2716,N_2619);
nand U2994 (N_2994,N_2718,N_2767);
and U2995 (N_2995,N_2703,N_2675);
and U2996 (N_2996,N_2739,N_2795);
and U2997 (N_2997,N_2673,N_2626);
nor U2998 (N_2998,N_2706,N_2627);
or U2999 (N_2999,N_2704,N_2624);
and U3000 (N_3000,N_2926,N_2808);
xnor U3001 (N_3001,N_2901,N_2958);
and U3002 (N_3002,N_2845,N_2805);
and U3003 (N_3003,N_2983,N_2948);
nand U3004 (N_3004,N_2955,N_2832);
nor U3005 (N_3005,N_2849,N_2954);
nor U3006 (N_3006,N_2892,N_2991);
nand U3007 (N_3007,N_2807,N_2820);
xor U3008 (N_3008,N_2887,N_2800);
nand U3009 (N_3009,N_2905,N_2931);
xor U3010 (N_3010,N_2930,N_2912);
and U3011 (N_3011,N_2816,N_2866);
nor U3012 (N_3012,N_2921,N_2852);
nand U3013 (N_3013,N_2864,N_2994);
and U3014 (N_3014,N_2821,N_2969);
nor U3015 (N_3015,N_2967,N_2950);
nand U3016 (N_3016,N_2959,N_2996);
or U3017 (N_3017,N_2970,N_2987);
nand U3018 (N_3018,N_2842,N_2916);
xnor U3019 (N_3019,N_2982,N_2939);
nor U3020 (N_3020,N_2839,N_2928);
nor U3021 (N_3021,N_2848,N_2992);
and U3022 (N_3022,N_2968,N_2846);
nand U3023 (N_3023,N_2896,N_2876);
and U3024 (N_3024,N_2833,N_2999);
and U3025 (N_3025,N_2953,N_2934);
and U3026 (N_3026,N_2838,N_2927);
nor U3027 (N_3027,N_2988,N_2853);
nor U3028 (N_3028,N_2998,N_2925);
nand U3029 (N_3029,N_2837,N_2936);
nor U3030 (N_3030,N_2872,N_2875);
nor U3031 (N_3031,N_2865,N_2840);
nor U3032 (N_3032,N_2903,N_2803);
xnor U3033 (N_3033,N_2888,N_2918);
nand U3034 (N_3034,N_2861,N_2862);
and U3035 (N_3035,N_2924,N_2834);
or U3036 (N_3036,N_2985,N_2801);
or U3037 (N_3037,N_2917,N_2871);
nand U3038 (N_3038,N_2910,N_2806);
nor U3039 (N_3039,N_2886,N_2858);
and U3040 (N_3040,N_2895,N_2913);
nand U3041 (N_3041,N_2824,N_2880);
or U3042 (N_3042,N_2812,N_2810);
xor U3043 (N_3043,N_2965,N_2981);
nor U3044 (N_3044,N_2818,N_2831);
nand U3045 (N_3045,N_2919,N_2822);
nor U3046 (N_3046,N_2972,N_2836);
xor U3047 (N_3047,N_2851,N_2827);
nor U3048 (N_3048,N_2932,N_2922);
nand U3049 (N_3049,N_2937,N_2802);
and U3050 (N_3050,N_2859,N_2945);
nor U3051 (N_3051,N_2975,N_2980);
nand U3052 (N_3052,N_2949,N_2835);
or U3053 (N_3053,N_2877,N_2946);
and U3054 (N_3054,N_2863,N_2941);
nor U3055 (N_3055,N_2828,N_2860);
nor U3056 (N_3056,N_2898,N_2973);
and U3057 (N_3057,N_2993,N_2885);
nor U3058 (N_3058,N_2890,N_2811);
and U3059 (N_3059,N_2889,N_2881);
and U3060 (N_3060,N_2900,N_2868);
and U3061 (N_3061,N_2979,N_2947);
and U3062 (N_3062,N_2929,N_2915);
or U3063 (N_3063,N_2984,N_2944);
or U3064 (N_3064,N_2914,N_2844);
or U3065 (N_3065,N_2809,N_2964);
nor U3066 (N_3066,N_2943,N_2935);
nand U3067 (N_3067,N_2904,N_2908);
xor U3068 (N_3068,N_2951,N_2823);
nor U3069 (N_3069,N_2867,N_2976);
nand U3070 (N_3070,N_2879,N_2971);
and U3071 (N_3071,N_2902,N_2826);
nor U3072 (N_3072,N_2986,N_2894);
or U3073 (N_3073,N_2883,N_2974);
and U3074 (N_3074,N_2966,N_2893);
nor U3075 (N_3075,N_2813,N_2957);
and U3076 (N_3076,N_2899,N_2874);
and U3077 (N_3077,N_2920,N_2873);
nor U3078 (N_3078,N_2830,N_2847);
nor U3079 (N_3079,N_2978,N_2963);
or U3080 (N_3080,N_2884,N_2850);
nor U3081 (N_3081,N_2841,N_2878);
and U3082 (N_3082,N_2854,N_2819);
xor U3083 (N_3083,N_2961,N_2815);
nor U3084 (N_3084,N_2960,N_2829);
nor U3085 (N_3085,N_2855,N_2843);
and U3086 (N_3086,N_2857,N_2962);
xor U3087 (N_3087,N_2897,N_2956);
nand U3088 (N_3088,N_2923,N_2869);
and U3089 (N_3089,N_2909,N_2989);
and U3090 (N_3090,N_2940,N_2907);
and U3091 (N_3091,N_2804,N_2942);
and U3092 (N_3092,N_2911,N_2906);
nor U3093 (N_3093,N_2817,N_2856);
or U3094 (N_3094,N_2825,N_2870);
nand U3095 (N_3095,N_2977,N_2891);
and U3096 (N_3096,N_2938,N_2952);
nand U3097 (N_3097,N_2933,N_2995);
nor U3098 (N_3098,N_2990,N_2882);
and U3099 (N_3099,N_2997,N_2814);
nor U3100 (N_3100,N_2984,N_2962);
and U3101 (N_3101,N_2827,N_2902);
xnor U3102 (N_3102,N_2985,N_2928);
nor U3103 (N_3103,N_2879,N_2916);
nor U3104 (N_3104,N_2836,N_2843);
nor U3105 (N_3105,N_2993,N_2865);
or U3106 (N_3106,N_2932,N_2843);
nand U3107 (N_3107,N_2913,N_2899);
and U3108 (N_3108,N_2801,N_2847);
and U3109 (N_3109,N_2966,N_2837);
and U3110 (N_3110,N_2987,N_2861);
and U3111 (N_3111,N_2903,N_2827);
nand U3112 (N_3112,N_2853,N_2818);
xnor U3113 (N_3113,N_2903,N_2851);
nor U3114 (N_3114,N_2882,N_2902);
nand U3115 (N_3115,N_2857,N_2918);
nor U3116 (N_3116,N_2907,N_2910);
and U3117 (N_3117,N_2835,N_2824);
nor U3118 (N_3118,N_2824,N_2899);
or U3119 (N_3119,N_2822,N_2927);
xnor U3120 (N_3120,N_2904,N_2901);
and U3121 (N_3121,N_2973,N_2891);
or U3122 (N_3122,N_2976,N_2852);
nand U3123 (N_3123,N_2935,N_2960);
and U3124 (N_3124,N_2940,N_2877);
or U3125 (N_3125,N_2857,N_2867);
nand U3126 (N_3126,N_2910,N_2857);
or U3127 (N_3127,N_2882,N_2981);
nor U3128 (N_3128,N_2873,N_2828);
nand U3129 (N_3129,N_2905,N_2821);
or U3130 (N_3130,N_2976,N_2848);
nand U3131 (N_3131,N_2806,N_2903);
and U3132 (N_3132,N_2950,N_2951);
nand U3133 (N_3133,N_2986,N_2996);
nor U3134 (N_3134,N_2982,N_2997);
and U3135 (N_3135,N_2830,N_2870);
and U3136 (N_3136,N_2965,N_2836);
nand U3137 (N_3137,N_2867,N_2982);
or U3138 (N_3138,N_2823,N_2828);
and U3139 (N_3139,N_2856,N_2993);
or U3140 (N_3140,N_2945,N_2982);
nand U3141 (N_3141,N_2906,N_2853);
or U3142 (N_3142,N_2928,N_2933);
nor U3143 (N_3143,N_2999,N_2929);
nand U3144 (N_3144,N_2915,N_2814);
and U3145 (N_3145,N_2897,N_2872);
xnor U3146 (N_3146,N_2938,N_2908);
xnor U3147 (N_3147,N_2816,N_2954);
nor U3148 (N_3148,N_2804,N_2895);
and U3149 (N_3149,N_2986,N_2846);
nand U3150 (N_3150,N_2810,N_2840);
and U3151 (N_3151,N_2829,N_2885);
and U3152 (N_3152,N_2971,N_2949);
nand U3153 (N_3153,N_2874,N_2904);
nand U3154 (N_3154,N_2858,N_2846);
nand U3155 (N_3155,N_2816,N_2840);
nor U3156 (N_3156,N_2815,N_2872);
nor U3157 (N_3157,N_2925,N_2857);
xnor U3158 (N_3158,N_2808,N_2923);
nand U3159 (N_3159,N_2972,N_2806);
and U3160 (N_3160,N_2965,N_2966);
nor U3161 (N_3161,N_2952,N_2826);
nor U3162 (N_3162,N_2816,N_2834);
and U3163 (N_3163,N_2924,N_2854);
nand U3164 (N_3164,N_2866,N_2897);
nand U3165 (N_3165,N_2839,N_2887);
nor U3166 (N_3166,N_2908,N_2815);
nand U3167 (N_3167,N_2847,N_2928);
or U3168 (N_3168,N_2983,N_2927);
nor U3169 (N_3169,N_2853,N_2907);
xnor U3170 (N_3170,N_2901,N_2851);
nand U3171 (N_3171,N_2981,N_2855);
or U3172 (N_3172,N_2887,N_2922);
nor U3173 (N_3173,N_2895,N_2832);
and U3174 (N_3174,N_2890,N_2937);
nor U3175 (N_3175,N_2923,N_2852);
xnor U3176 (N_3176,N_2958,N_2847);
nand U3177 (N_3177,N_2934,N_2998);
xnor U3178 (N_3178,N_2848,N_2940);
xnor U3179 (N_3179,N_2827,N_2980);
or U3180 (N_3180,N_2943,N_2940);
and U3181 (N_3181,N_2860,N_2835);
nor U3182 (N_3182,N_2821,N_2894);
nand U3183 (N_3183,N_2820,N_2819);
nand U3184 (N_3184,N_2857,N_2974);
nor U3185 (N_3185,N_2803,N_2833);
nand U3186 (N_3186,N_2814,N_2863);
nor U3187 (N_3187,N_2976,N_2835);
nand U3188 (N_3188,N_2931,N_2854);
or U3189 (N_3189,N_2957,N_2845);
xnor U3190 (N_3190,N_2912,N_2800);
xor U3191 (N_3191,N_2916,N_2848);
nand U3192 (N_3192,N_2889,N_2963);
or U3193 (N_3193,N_2826,N_2815);
nor U3194 (N_3194,N_2877,N_2965);
and U3195 (N_3195,N_2846,N_2811);
nand U3196 (N_3196,N_2987,N_2868);
or U3197 (N_3197,N_2934,N_2948);
or U3198 (N_3198,N_2898,N_2803);
or U3199 (N_3199,N_2935,N_2921);
nor U3200 (N_3200,N_3111,N_3071);
nand U3201 (N_3201,N_3005,N_3123);
nand U3202 (N_3202,N_3021,N_3053);
and U3203 (N_3203,N_3184,N_3116);
xnor U3204 (N_3204,N_3019,N_3155);
or U3205 (N_3205,N_3008,N_3161);
nand U3206 (N_3206,N_3108,N_3121);
nand U3207 (N_3207,N_3105,N_3074);
and U3208 (N_3208,N_3082,N_3139);
or U3209 (N_3209,N_3001,N_3157);
nor U3210 (N_3210,N_3078,N_3158);
or U3211 (N_3211,N_3007,N_3093);
and U3212 (N_3212,N_3138,N_3022);
nor U3213 (N_3213,N_3118,N_3065);
nor U3214 (N_3214,N_3058,N_3133);
nand U3215 (N_3215,N_3024,N_3183);
and U3216 (N_3216,N_3143,N_3057);
or U3217 (N_3217,N_3044,N_3012);
or U3218 (N_3218,N_3179,N_3145);
and U3219 (N_3219,N_3195,N_3085);
and U3220 (N_3220,N_3120,N_3172);
nor U3221 (N_3221,N_3055,N_3064);
nor U3222 (N_3222,N_3102,N_3114);
and U3223 (N_3223,N_3156,N_3162);
nor U3224 (N_3224,N_3177,N_3091);
or U3225 (N_3225,N_3199,N_3198);
or U3226 (N_3226,N_3170,N_3174);
nor U3227 (N_3227,N_3049,N_3169);
nor U3228 (N_3228,N_3164,N_3081);
or U3229 (N_3229,N_3115,N_3073);
xnor U3230 (N_3230,N_3038,N_3059);
nor U3231 (N_3231,N_3186,N_3188);
or U3232 (N_3232,N_3016,N_3029);
nand U3233 (N_3233,N_3094,N_3051);
or U3234 (N_3234,N_3002,N_3176);
nand U3235 (N_3235,N_3086,N_3084);
and U3236 (N_3236,N_3066,N_3144);
xor U3237 (N_3237,N_3089,N_3150);
or U3238 (N_3238,N_3072,N_3095);
or U3239 (N_3239,N_3042,N_3100);
nand U3240 (N_3240,N_3032,N_3031);
and U3241 (N_3241,N_3087,N_3125);
nand U3242 (N_3242,N_3110,N_3165);
and U3243 (N_3243,N_3026,N_3122);
nor U3244 (N_3244,N_3182,N_3126);
and U3245 (N_3245,N_3140,N_3017);
nor U3246 (N_3246,N_3061,N_3068);
or U3247 (N_3247,N_3023,N_3043);
and U3248 (N_3248,N_3197,N_3141);
nand U3249 (N_3249,N_3039,N_3027);
and U3250 (N_3250,N_3171,N_3113);
nand U3251 (N_3251,N_3062,N_3040);
nor U3252 (N_3252,N_3135,N_3018);
and U3253 (N_3253,N_3104,N_3028);
nor U3254 (N_3254,N_3079,N_3025);
and U3255 (N_3255,N_3099,N_3088);
xor U3256 (N_3256,N_3180,N_3033);
xor U3257 (N_3257,N_3098,N_3075);
nand U3258 (N_3258,N_3127,N_3154);
and U3259 (N_3259,N_3148,N_3096);
or U3260 (N_3260,N_3142,N_3151);
and U3261 (N_3261,N_3112,N_3146);
or U3262 (N_3262,N_3175,N_3119);
or U3263 (N_3263,N_3192,N_3054);
and U3264 (N_3264,N_3067,N_3130);
and U3265 (N_3265,N_3106,N_3129);
or U3266 (N_3266,N_3006,N_3196);
and U3267 (N_3267,N_3009,N_3034);
nor U3268 (N_3268,N_3041,N_3004);
and U3269 (N_3269,N_3101,N_3134);
or U3270 (N_3270,N_3046,N_3163);
and U3271 (N_3271,N_3076,N_3069);
xnor U3272 (N_3272,N_3160,N_3070);
nand U3273 (N_3273,N_3083,N_3036);
nand U3274 (N_3274,N_3097,N_3050);
and U3275 (N_3275,N_3137,N_3077);
or U3276 (N_3276,N_3152,N_3149);
or U3277 (N_3277,N_3153,N_3159);
nand U3278 (N_3278,N_3030,N_3013);
nand U3279 (N_3279,N_3092,N_3037);
nor U3280 (N_3280,N_3173,N_3168);
nand U3281 (N_3281,N_3190,N_3187);
and U3282 (N_3282,N_3003,N_3147);
and U3283 (N_3283,N_3193,N_3056);
nand U3284 (N_3284,N_3048,N_3080);
xnor U3285 (N_3285,N_3045,N_3191);
nor U3286 (N_3286,N_3063,N_3117);
nand U3287 (N_3287,N_3136,N_3047);
and U3288 (N_3288,N_3178,N_3181);
and U3289 (N_3289,N_3020,N_3015);
or U3290 (N_3290,N_3166,N_3132);
and U3291 (N_3291,N_3124,N_3035);
nand U3292 (N_3292,N_3131,N_3194);
or U3293 (N_3293,N_3185,N_3000);
and U3294 (N_3294,N_3060,N_3010);
and U3295 (N_3295,N_3167,N_3189);
nor U3296 (N_3296,N_3011,N_3107);
nor U3297 (N_3297,N_3128,N_3103);
and U3298 (N_3298,N_3052,N_3109);
nand U3299 (N_3299,N_3090,N_3014);
nor U3300 (N_3300,N_3170,N_3008);
xor U3301 (N_3301,N_3191,N_3168);
and U3302 (N_3302,N_3160,N_3071);
nand U3303 (N_3303,N_3098,N_3184);
or U3304 (N_3304,N_3139,N_3019);
or U3305 (N_3305,N_3002,N_3137);
nand U3306 (N_3306,N_3038,N_3146);
and U3307 (N_3307,N_3006,N_3173);
nand U3308 (N_3308,N_3049,N_3109);
and U3309 (N_3309,N_3002,N_3054);
and U3310 (N_3310,N_3031,N_3124);
nand U3311 (N_3311,N_3143,N_3056);
xor U3312 (N_3312,N_3044,N_3188);
and U3313 (N_3313,N_3051,N_3088);
and U3314 (N_3314,N_3006,N_3026);
nand U3315 (N_3315,N_3116,N_3064);
nor U3316 (N_3316,N_3059,N_3144);
and U3317 (N_3317,N_3168,N_3174);
nor U3318 (N_3318,N_3011,N_3189);
nand U3319 (N_3319,N_3040,N_3167);
or U3320 (N_3320,N_3008,N_3071);
or U3321 (N_3321,N_3115,N_3186);
nand U3322 (N_3322,N_3077,N_3023);
nand U3323 (N_3323,N_3199,N_3082);
and U3324 (N_3324,N_3080,N_3167);
or U3325 (N_3325,N_3058,N_3186);
nand U3326 (N_3326,N_3153,N_3051);
and U3327 (N_3327,N_3193,N_3112);
and U3328 (N_3328,N_3060,N_3084);
nand U3329 (N_3329,N_3054,N_3115);
and U3330 (N_3330,N_3101,N_3188);
and U3331 (N_3331,N_3041,N_3012);
nand U3332 (N_3332,N_3049,N_3059);
nand U3333 (N_3333,N_3139,N_3179);
and U3334 (N_3334,N_3021,N_3056);
and U3335 (N_3335,N_3130,N_3147);
or U3336 (N_3336,N_3016,N_3074);
nor U3337 (N_3337,N_3168,N_3084);
and U3338 (N_3338,N_3147,N_3085);
nand U3339 (N_3339,N_3098,N_3180);
or U3340 (N_3340,N_3121,N_3079);
nand U3341 (N_3341,N_3032,N_3083);
and U3342 (N_3342,N_3139,N_3133);
xnor U3343 (N_3343,N_3086,N_3130);
or U3344 (N_3344,N_3179,N_3042);
and U3345 (N_3345,N_3167,N_3007);
or U3346 (N_3346,N_3086,N_3046);
nand U3347 (N_3347,N_3168,N_3158);
nor U3348 (N_3348,N_3051,N_3150);
nor U3349 (N_3349,N_3086,N_3015);
and U3350 (N_3350,N_3188,N_3182);
and U3351 (N_3351,N_3094,N_3103);
and U3352 (N_3352,N_3159,N_3024);
and U3353 (N_3353,N_3075,N_3192);
xnor U3354 (N_3354,N_3013,N_3088);
nand U3355 (N_3355,N_3125,N_3092);
and U3356 (N_3356,N_3152,N_3086);
nor U3357 (N_3357,N_3092,N_3155);
nor U3358 (N_3358,N_3073,N_3000);
and U3359 (N_3359,N_3046,N_3075);
or U3360 (N_3360,N_3063,N_3027);
and U3361 (N_3361,N_3129,N_3104);
or U3362 (N_3362,N_3117,N_3066);
and U3363 (N_3363,N_3027,N_3107);
nor U3364 (N_3364,N_3165,N_3168);
xor U3365 (N_3365,N_3018,N_3120);
or U3366 (N_3366,N_3057,N_3055);
and U3367 (N_3367,N_3094,N_3168);
or U3368 (N_3368,N_3016,N_3132);
or U3369 (N_3369,N_3086,N_3021);
and U3370 (N_3370,N_3025,N_3006);
nand U3371 (N_3371,N_3182,N_3016);
xor U3372 (N_3372,N_3195,N_3002);
nor U3373 (N_3373,N_3150,N_3185);
and U3374 (N_3374,N_3110,N_3187);
xor U3375 (N_3375,N_3181,N_3119);
nand U3376 (N_3376,N_3128,N_3038);
nor U3377 (N_3377,N_3159,N_3156);
or U3378 (N_3378,N_3014,N_3009);
nand U3379 (N_3379,N_3186,N_3135);
and U3380 (N_3380,N_3066,N_3033);
or U3381 (N_3381,N_3074,N_3134);
or U3382 (N_3382,N_3077,N_3027);
or U3383 (N_3383,N_3101,N_3172);
or U3384 (N_3384,N_3171,N_3181);
or U3385 (N_3385,N_3167,N_3005);
and U3386 (N_3386,N_3115,N_3017);
nand U3387 (N_3387,N_3163,N_3022);
xnor U3388 (N_3388,N_3080,N_3055);
nand U3389 (N_3389,N_3143,N_3085);
xnor U3390 (N_3390,N_3168,N_3079);
nand U3391 (N_3391,N_3099,N_3175);
xor U3392 (N_3392,N_3155,N_3008);
nor U3393 (N_3393,N_3086,N_3114);
and U3394 (N_3394,N_3092,N_3168);
nor U3395 (N_3395,N_3076,N_3129);
xor U3396 (N_3396,N_3129,N_3047);
nand U3397 (N_3397,N_3176,N_3061);
nand U3398 (N_3398,N_3154,N_3010);
nor U3399 (N_3399,N_3076,N_3050);
nand U3400 (N_3400,N_3204,N_3252);
xnor U3401 (N_3401,N_3337,N_3275);
nand U3402 (N_3402,N_3300,N_3269);
nor U3403 (N_3403,N_3302,N_3293);
xnor U3404 (N_3404,N_3336,N_3355);
xor U3405 (N_3405,N_3299,N_3289);
xnor U3406 (N_3406,N_3345,N_3283);
and U3407 (N_3407,N_3365,N_3236);
nand U3408 (N_3408,N_3344,N_3328);
and U3409 (N_3409,N_3231,N_3317);
and U3410 (N_3410,N_3377,N_3376);
and U3411 (N_3411,N_3330,N_3214);
and U3412 (N_3412,N_3284,N_3303);
nand U3413 (N_3413,N_3335,N_3371);
nand U3414 (N_3414,N_3260,N_3381);
nand U3415 (N_3415,N_3228,N_3280);
and U3416 (N_3416,N_3395,N_3202);
and U3417 (N_3417,N_3287,N_3205);
or U3418 (N_3418,N_3351,N_3346);
nand U3419 (N_3419,N_3398,N_3232);
nand U3420 (N_3420,N_3243,N_3257);
nand U3421 (N_3421,N_3313,N_3307);
or U3422 (N_3422,N_3209,N_3250);
nand U3423 (N_3423,N_3273,N_3315);
nor U3424 (N_3424,N_3279,N_3352);
nand U3425 (N_3425,N_3251,N_3271);
and U3426 (N_3426,N_3255,N_3217);
and U3427 (N_3427,N_3341,N_3382);
and U3428 (N_3428,N_3226,N_3241);
and U3429 (N_3429,N_3294,N_3270);
nor U3430 (N_3430,N_3379,N_3316);
nor U3431 (N_3431,N_3334,N_3372);
and U3432 (N_3432,N_3218,N_3342);
and U3433 (N_3433,N_3314,N_3399);
or U3434 (N_3434,N_3210,N_3272);
nand U3435 (N_3435,N_3348,N_3235);
nor U3436 (N_3436,N_3396,N_3246);
nand U3437 (N_3437,N_3301,N_3309);
nand U3438 (N_3438,N_3224,N_3230);
nor U3439 (N_3439,N_3333,N_3350);
xnor U3440 (N_3440,N_3207,N_3208);
and U3441 (N_3441,N_3215,N_3362);
xor U3442 (N_3442,N_3206,N_3237);
xnor U3443 (N_3443,N_3201,N_3331);
or U3444 (N_3444,N_3332,N_3353);
nor U3445 (N_3445,N_3385,N_3364);
nor U3446 (N_3446,N_3292,N_3378);
or U3447 (N_3447,N_3325,N_3295);
and U3448 (N_3448,N_3291,N_3388);
nand U3449 (N_3449,N_3222,N_3264);
nand U3450 (N_3450,N_3373,N_3323);
or U3451 (N_3451,N_3339,N_3220);
or U3452 (N_3452,N_3312,N_3389);
xnor U3453 (N_3453,N_3391,N_3225);
or U3454 (N_3454,N_3253,N_3261);
nor U3455 (N_3455,N_3256,N_3211);
nand U3456 (N_3456,N_3296,N_3240);
or U3457 (N_3457,N_3239,N_3259);
nand U3458 (N_3458,N_3213,N_3340);
and U3459 (N_3459,N_3266,N_3258);
and U3460 (N_3460,N_3282,N_3227);
and U3461 (N_3461,N_3268,N_3212);
nor U3462 (N_3462,N_3276,N_3308);
nand U3463 (N_3463,N_3216,N_3393);
or U3464 (N_3464,N_3367,N_3358);
nor U3465 (N_3465,N_3265,N_3356);
nand U3466 (N_3466,N_3326,N_3380);
nand U3467 (N_3467,N_3360,N_3278);
nor U3468 (N_3468,N_3368,N_3329);
nand U3469 (N_3469,N_3200,N_3277);
nand U3470 (N_3470,N_3392,N_3286);
or U3471 (N_3471,N_3263,N_3375);
nand U3472 (N_3472,N_3361,N_3238);
or U3473 (N_3473,N_3384,N_3249);
nor U3474 (N_3474,N_3248,N_3394);
nor U3475 (N_3475,N_3319,N_3244);
and U3476 (N_3476,N_3318,N_3359);
nor U3477 (N_3477,N_3387,N_3290);
xnor U3478 (N_3478,N_3305,N_3233);
nor U3479 (N_3479,N_3321,N_3297);
or U3480 (N_3480,N_3310,N_3322);
and U3481 (N_3481,N_3254,N_3320);
and U3482 (N_3482,N_3370,N_3203);
xor U3483 (N_3483,N_3285,N_3229);
or U3484 (N_3484,N_3369,N_3349);
nor U3485 (N_3485,N_3223,N_3374);
nand U3486 (N_3486,N_3363,N_3247);
nor U3487 (N_3487,N_3221,N_3267);
and U3488 (N_3488,N_3397,N_3347);
and U3489 (N_3489,N_3366,N_3390);
and U3490 (N_3490,N_3304,N_3354);
or U3491 (N_3491,N_3245,N_3324);
and U3492 (N_3492,N_3298,N_3234);
and U3493 (N_3493,N_3262,N_3288);
xor U3494 (N_3494,N_3383,N_3311);
or U3495 (N_3495,N_3327,N_3242);
and U3496 (N_3496,N_3281,N_3338);
nor U3497 (N_3497,N_3357,N_3343);
or U3498 (N_3498,N_3386,N_3274);
or U3499 (N_3499,N_3306,N_3219);
nand U3500 (N_3500,N_3266,N_3337);
nand U3501 (N_3501,N_3280,N_3207);
nor U3502 (N_3502,N_3362,N_3344);
nand U3503 (N_3503,N_3332,N_3247);
nand U3504 (N_3504,N_3397,N_3364);
nor U3505 (N_3505,N_3388,N_3315);
and U3506 (N_3506,N_3292,N_3274);
nor U3507 (N_3507,N_3214,N_3267);
and U3508 (N_3508,N_3353,N_3315);
nor U3509 (N_3509,N_3387,N_3382);
or U3510 (N_3510,N_3318,N_3252);
or U3511 (N_3511,N_3279,N_3203);
nand U3512 (N_3512,N_3259,N_3283);
and U3513 (N_3513,N_3259,N_3270);
nor U3514 (N_3514,N_3221,N_3237);
or U3515 (N_3515,N_3220,N_3232);
nor U3516 (N_3516,N_3295,N_3365);
nor U3517 (N_3517,N_3250,N_3346);
or U3518 (N_3518,N_3265,N_3354);
or U3519 (N_3519,N_3301,N_3359);
xor U3520 (N_3520,N_3375,N_3231);
xnor U3521 (N_3521,N_3332,N_3297);
and U3522 (N_3522,N_3363,N_3362);
and U3523 (N_3523,N_3260,N_3312);
xnor U3524 (N_3524,N_3350,N_3204);
or U3525 (N_3525,N_3316,N_3373);
or U3526 (N_3526,N_3334,N_3292);
nand U3527 (N_3527,N_3309,N_3398);
nand U3528 (N_3528,N_3397,N_3226);
nand U3529 (N_3529,N_3287,N_3391);
or U3530 (N_3530,N_3374,N_3263);
and U3531 (N_3531,N_3276,N_3346);
and U3532 (N_3532,N_3234,N_3351);
nand U3533 (N_3533,N_3239,N_3392);
nor U3534 (N_3534,N_3222,N_3279);
nand U3535 (N_3535,N_3359,N_3316);
nor U3536 (N_3536,N_3321,N_3271);
xnor U3537 (N_3537,N_3208,N_3258);
or U3538 (N_3538,N_3320,N_3337);
and U3539 (N_3539,N_3355,N_3347);
or U3540 (N_3540,N_3209,N_3394);
or U3541 (N_3541,N_3283,N_3328);
and U3542 (N_3542,N_3254,N_3317);
or U3543 (N_3543,N_3332,N_3339);
xnor U3544 (N_3544,N_3240,N_3264);
and U3545 (N_3545,N_3397,N_3204);
nor U3546 (N_3546,N_3361,N_3303);
and U3547 (N_3547,N_3360,N_3354);
or U3548 (N_3548,N_3230,N_3316);
xor U3549 (N_3549,N_3245,N_3303);
xor U3550 (N_3550,N_3231,N_3370);
nor U3551 (N_3551,N_3201,N_3205);
xor U3552 (N_3552,N_3293,N_3350);
or U3553 (N_3553,N_3339,N_3207);
nand U3554 (N_3554,N_3308,N_3340);
or U3555 (N_3555,N_3234,N_3317);
and U3556 (N_3556,N_3230,N_3233);
and U3557 (N_3557,N_3284,N_3254);
nor U3558 (N_3558,N_3222,N_3212);
nand U3559 (N_3559,N_3277,N_3385);
nand U3560 (N_3560,N_3283,N_3204);
nand U3561 (N_3561,N_3290,N_3217);
nor U3562 (N_3562,N_3301,N_3263);
and U3563 (N_3563,N_3235,N_3244);
and U3564 (N_3564,N_3280,N_3250);
or U3565 (N_3565,N_3234,N_3399);
nand U3566 (N_3566,N_3253,N_3394);
and U3567 (N_3567,N_3374,N_3319);
nand U3568 (N_3568,N_3290,N_3208);
and U3569 (N_3569,N_3323,N_3249);
nand U3570 (N_3570,N_3257,N_3392);
nor U3571 (N_3571,N_3380,N_3278);
nand U3572 (N_3572,N_3358,N_3323);
nand U3573 (N_3573,N_3263,N_3272);
xor U3574 (N_3574,N_3335,N_3313);
nor U3575 (N_3575,N_3222,N_3246);
and U3576 (N_3576,N_3264,N_3250);
and U3577 (N_3577,N_3317,N_3252);
or U3578 (N_3578,N_3283,N_3334);
or U3579 (N_3579,N_3364,N_3362);
nor U3580 (N_3580,N_3335,N_3299);
or U3581 (N_3581,N_3271,N_3394);
or U3582 (N_3582,N_3348,N_3272);
nor U3583 (N_3583,N_3367,N_3382);
nand U3584 (N_3584,N_3274,N_3381);
or U3585 (N_3585,N_3255,N_3330);
nor U3586 (N_3586,N_3217,N_3397);
or U3587 (N_3587,N_3200,N_3312);
nor U3588 (N_3588,N_3289,N_3362);
nand U3589 (N_3589,N_3259,N_3202);
nand U3590 (N_3590,N_3280,N_3265);
and U3591 (N_3591,N_3220,N_3324);
xor U3592 (N_3592,N_3299,N_3328);
or U3593 (N_3593,N_3339,N_3248);
xnor U3594 (N_3594,N_3297,N_3339);
or U3595 (N_3595,N_3319,N_3252);
nor U3596 (N_3596,N_3343,N_3224);
nand U3597 (N_3597,N_3384,N_3230);
nor U3598 (N_3598,N_3277,N_3211);
and U3599 (N_3599,N_3294,N_3221);
xnor U3600 (N_3600,N_3551,N_3594);
nand U3601 (N_3601,N_3452,N_3510);
or U3602 (N_3602,N_3514,N_3417);
xor U3603 (N_3603,N_3506,N_3497);
and U3604 (N_3604,N_3424,N_3517);
nand U3605 (N_3605,N_3498,N_3410);
nor U3606 (N_3606,N_3531,N_3472);
nor U3607 (N_3607,N_3556,N_3580);
nand U3608 (N_3608,N_3496,N_3574);
nor U3609 (N_3609,N_3470,N_3445);
or U3610 (N_3610,N_3520,N_3555);
xnor U3611 (N_3611,N_3414,N_3469);
or U3612 (N_3612,N_3489,N_3546);
or U3613 (N_3613,N_3586,N_3494);
nand U3614 (N_3614,N_3433,N_3473);
and U3615 (N_3615,N_3513,N_3420);
nand U3616 (N_3616,N_3553,N_3522);
nor U3617 (N_3617,N_3461,N_3593);
and U3618 (N_3618,N_3563,N_3579);
nor U3619 (N_3619,N_3464,N_3523);
nand U3620 (N_3620,N_3495,N_3416);
and U3621 (N_3621,N_3462,N_3566);
or U3622 (N_3622,N_3584,N_3519);
and U3623 (N_3623,N_3577,N_3587);
nor U3624 (N_3624,N_3441,N_3509);
nor U3625 (N_3625,N_3434,N_3507);
and U3626 (N_3626,N_3467,N_3515);
nand U3627 (N_3627,N_3481,N_3528);
nand U3628 (N_3628,N_3501,N_3478);
nor U3629 (N_3629,N_3570,N_3552);
and U3630 (N_3630,N_3431,N_3599);
or U3631 (N_3631,N_3540,N_3482);
xnor U3632 (N_3632,N_3560,N_3533);
nand U3633 (N_3633,N_3585,N_3572);
and U3634 (N_3634,N_3526,N_3554);
xnor U3635 (N_3635,N_3457,N_3402);
xor U3636 (N_3636,N_3548,N_3407);
nor U3637 (N_3637,N_3581,N_3530);
and U3638 (N_3638,N_3409,N_3449);
or U3639 (N_3639,N_3471,N_3539);
or U3640 (N_3640,N_3408,N_3400);
nand U3641 (N_3641,N_3588,N_3479);
nand U3642 (N_3642,N_3592,N_3569);
nor U3643 (N_3643,N_3578,N_3484);
or U3644 (N_3644,N_3442,N_3536);
nand U3645 (N_3645,N_3568,N_3550);
nor U3646 (N_3646,N_3589,N_3521);
or U3647 (N_3647,N_3440,N_3465);
nor U3648 (N_3648,N_3456,N_3450);
xor U3649 (N_3649,N_3518,N_3541);
nand U3650 (N_3650,N_3524,N_3538);
and U3651 (N_3651,N_3547,N_3545);
xnor U3652 (N_3652,N_3418,N_3525);
and U3653 (N_3653,N_3483,N_3542);
and U3654 (N_3654,N_3534,N_3564);
nor U3655 (N_3655,N_3595,N_3544);
and U3656 (N_3656,N_3425,N_3591);
nor U3657 (N_3657,N_3446,N_3590);
nand U3658 (N_3658,N_3537,N_3435);
and U3659 (N_3659,N_3490,N_3411);
nand U3660 (N_3660,N_3432,N_3403);
and U3661 (N_3661,N_3573,N_3406);
xnor U3662 (N_3662,N_3502,N_3582);
and U3663 (N_3663,N_3576,N_3447);
nor U3664 (N_3664,N_3468,N_3421);
or U3665 (N_3665,N_3437,N_3529);
nand U3666 (N_3666,N_3413,N_3558);
or U3667 (N_3667,N_3429,N_3565);
and U3668 (N_3668,N_3444,N_3448);
or U3669 (N_3669,N_3598,N_3428);
or U3670 (N_3670,N_3476,N_3549);
nor U3671 (N_3671,N_3493,N_3485);
nor U3672 (N_3672,N_3597,N_3415);
nand U3673 (N_3673,N_3527,N_3405);
or U3674 (N_3674,N_3487,N_3412);
or U3675 (N_3675,N_3500,N_3453);
xnor U3676 (N_3676,N_3532,N_3423);
and U3677 (N_3677,N_3426,N_3427);
and U3678 (N_3678,N_3443,N_3477);
and U3679 (N_3679,N_3562,N_3488);
and U3680 (N_3680,N_3454,N_3575);
or U3681 (N_3681,N_3559,N_3512);
nor U3682 (N_3682,N_3596,N_3475);
and U3683 (N_3683,N_3463,N_3571);
or U3684 (N_3684,N_3466,N_3543);
nor U3685 (N_3685,N_3583,N_3504);
nor U3686 (N_3686,N_3535,N_3511);
and U3687 (N_3687,N_3567,N_3436);
xnor U3688 (N_3688,N_3505,N_3401);
xnor U3689 (N_3689,N_3430,N_3516);
or U3690 (N_3690,N_3459,N_3491);
and U3691 (N_3691,N_3451,N_3474);
nor U3692 (N_3692,N_3458,N_3508);
xnor U3693 (N_3693,N_3422,N_3499);
nand U3694 (N_3694,N_3486,N_3561);
or U3695 (N_3695,N_3492,N_3438);
and U3696 (N_3696,N_3439,N_3419);
and U3697 (N_3697,N_3460,N_3557);
nor U3698 (N_3698,N_3480,N_3503);
xor U3699 (N_3699,N_3455,N_3404);
nor U3700 (N_3700,N_3466,N_3541);
or U3701 (N_3701,N_3471,N_3472);
and U3702 (N_3702,N_3502,N_3400);
or U3703 (N_3703,N_3534,N_3557);
nand U3704 (N_3704,N_3414,N_3505);
nand U3705 (N_3705,N_3425,N_3494);
nand U3706 (N_3706,N_3524,N_3504);
and U3707 (N_3707,N_3474,N_3486);
and U3708 (N_3708,N_3465,N_3446);
and U3709 (N_3709,N_3440,N_3563);
or U3710 (N_3710,N_3524,N_3511);
nor U3711 (N_3711,N_3446,N_3480);
nand U3712 (N_3712,N_3408,N_3528);
nand U3713 (N_3713,N_3557,N_3527);
or U3714 (N_3714,N_3430,N_3537);
nor U3715 (N_3715,N_3457,N_3507);
or U3716 (N_3716,N_3410,N_3539);
nor U3717 (N_3717,N_3596,N_3442);
nand U3718 (N_3718,N_3468,N_3496);
and U3719 (N_3719,N_3446,N_3441);
xor U3720 (N_3720,N_3515,N_3477);
and U3721 (N_3721,N_3466,N_3438);
or U3722 (N_3722,N_3516,N_3543);
and U3723 (N_3723,N_3516,N_3483);
nand U3724 (N_3724,N_3565,N_3448);
xor U3725 (N_3725,N_3486,N_3525);
or U3726 (N_3726,N_3422,N_3554);
nor U3727 (N_3727,N_3515,N_3497);
nand U3728 (N_3728,N_3556,N_3454);
and U3729 (N_3729,N_3476,N_3508);
nand U3730 (N_3730,N_3410,N_3554);
nor U3731 (N_3731,N_3585,N_3437);
nor U3732 (N_3732,N_3534,N_3489);
or U3733 (N_3733,N_3580,N_3529);
or U3734 (N_3734,N_3505,N_3591);
or U3735 (N_3735,N_3582,N_3432);
nand U3736 (N_3736,N_3466,N_3444);
nor U3737 (N_3737,N_3462,N_3510);
or U3738 (N_3738,N_3513,N_3430);
xor U3739 (N_3739,N_3431,N_3516);
and U3740 (N_3740,N_3439,N_3590);
nand U3741 (N_3741,N_3593,N_3525);
and U3742 (N_3742,N_3401,N_3457);
or U3743 (N_3743,N_3406,N_3501);
or U3744 (N_3744,N_3469,N_3455);
nor U3745 (N_3745,N_3527,N_3531);
or U3746 (N_3746,N_3464,N_3435);
nor U3747 (N_3747,N_3589,N_3430);
or U3748 (N_3748,N_3483,N_3465);
nor U3749 (N_3749,N_3424,N_3559);
xor U3750 (N_3750,N_3413,N_3563);
or U3751 (N_3751,N_3559,N_3577);
and U3752 (N_3752,N_3461,N_3541);
and U3753 (N_3753,N_3467,N_3512);
nand U3754 (N_3754,N_3502,N_3480);
and U3755 (N_3755,N_3583,N_3429);
nand U3756 (N_3756,N_3436,N_3412);
or U3757 (N_3757,N_3478,N_3563);
and U3758 (N_3758,N_3479,N_3501);
or U3759 (N_3759,N_3555,N_3597);
nand U3760 (N_3760,N_3548,N_3489);
and U3761 (N_3761,N_3547,N_3460);
nand U3762 (N_3762,N_3515,N_3431);
or U3763 (N_3763,N_3561,N_3441);
nand U3764 (N_3764,N_3505,N_3584);
and U3765 (N_3765,N_3554,N_3444);
nor U3766 (N_3766,N_3400,N_3517);
and U3767 (N_3767,N_3406,N_3414);
and U3768 (N_3768,N_3511,N_3421);
nor U3769 (N_3769,N_3419,N_3433);
nor U3770 (N_3770,N_3407,N_3490);
nor U3771 (N_3771,N_3560,N_3595);
and U3772 (N_3772,N_3400,N_3415);
nor U3773 (N_3773,N_3444,N_3531);
nand U3774 (N_3774,N_3462,N_3523);
xnor U3775 (N_3775,N_3499,N_3498);
nor U3776 (N_3776,N_3572,N_3573);
and U3777 (N_3777,N_3463,N_3585);
nor U3778 (N_3778,N_3428,N_3565);
and U3779 (N_3779,N_3405,N_3530);
xnor U3780 (N_3780,N_3489,N_3402);
nand U3781 (N_3781,N_3472,N_3458);
nor U3782 (N_3782,N_3539,N_3488);
xor U3783 (N_3783,N_3476,N_3414);
nor U3784 (N_3784,N_3524,N_3432);
xor U3785 (N_3785,N_3532,N_3576);
or U3786 (N_3786,N_3485,N_3599);
xnor U3787 (N_3787,N_3428,N_3483);
or U3788 (N_3788,N_3538,N_3565);
nor U3789 (N_3789,N_3581,N_3414);
nand U3790 (N_3790,N_3577,N_3474);
and U3791 (N_3791,N_3561,N_3472);
xnor U3792 (N_3792,N_3426,N_3490);
xnor U3793 (N_3793,N_3510,N_3405);
xor U3794 (N_3794,N_3483,N_3543);
and U3795 (N_3795,N_3598,N_3527);
xnor U3796 (N_3796,N_3464,N_3478);
nor U3797 (N_3797,N_3508,N_3527);
nand U3798 (N_3798,N_3509,N_3415);
or U3799 (N_3799,N_3495,N_3515);
or U3800 (N_3800,N_3756,N_3695);
nor U3801 (N_3801,N_3788,N_3650);
nand U3802 (N_3802,N_3630,N_3662);
nand U3803 (N_3803,N_3626,N_3785);
nor U3804 (N_3804,N_3734,N_3703);
and U3805 (N_3805,N_3745,N_3791);
nand U3806 (N_3806,N_3665,N_3746);
or U3807 (N_3807,N_3739,N_3713);
or U3808 (N_3808,N_3749,N_3609);
and U3809 (N_3809,N_3750,N_3670);
nor U3810 (N_3810,N_3751,N_3760);
nand U3811 (N_3811,N_3731,N_3774);
nor U3812 (N_3812,N_3709,N_3730);
nand U3813 (N_3813,N_3712,N_3759);
and U3814 (N_3814,N_3754,N_3762);
nor U3815 (N_3815,N_3702,N_3685);
and U3816 (N_3816,N_3629,N_3641);
nand U3817 (N_3817,N_3725,N_3614);
and U3818 (N_3818,N_3761,N_3744);
or U3819 (N_3819,N_3763,N_3663);
or U3820 (N_3820,N_3655,N_3622);
and U3821 (N_3821,N_3607,N_3621);
and U3822 (N_3822,N_3603,N_3741);
or U3823 (N_3823,N_3639,N_3775);
nand U3824 (N_3824,N_3707,N_3779);
nand U3825 (N_3825,N_3729,N_3782);
nor U3826 (N_3826,N_3638,N_3642);
nor U3827 (N_3827,N_3792,N_3628);
or U3828 (N_3828,N_3675,N_3631);
or U3829 (N_3829,N_3780,N_3740);
or U3830 (N_3830,N_3611,N_3752);
or U3831 (N_3831,N_3627,N_3795);
nor U3832 (N_3832,N_3689,N_3764);
and U3833 (N_3833,N_3719,N_3748);
and U3834 (N_3834,N_3784,N_3742);
or U3835 (N_3835,N_3700,N_3776);
and U3836 (N_3836,N_3677,N_3651);
nor U3837 (N_3837,N_3717,N_3654);
nand U3838 (N_3838,N_3796,N_3623);
nand U3839 (N_3839,N_3755,N_3687);
or U3840 (N_3840,N_3694,N_3757);
nor U3841 (N_3841,N_3600,N_3772);
and U3842 (N_3842,N_3679,N_3718);
nand U3843 (N_3843,N_3794,N_3653);
or U3844 (N_3844,N_3688,N_3736);
nand U3845 (N_3845,N_3649,N_3758);
nor U3846 (N_3846,N_3692,N_3624);
nor U3847 (N_3847,N_3714,N_3681);
xor U3848 (N_3848,N_3724,N_3766);
nor U3849 (N_3849,N_3643,N_3684);
or U3850 (N_3850,N_3723,N_3698);
or U3851 (N_3851,N_3733,N_3747);
xor U3852 (N_3852,N_3632,N_3738);
nand U3853 (N_3853,N_3678,N_3706);
nand U3854 (N_3854,N_3767,N_3682);
nor U3855 (N_3855,N_3640,N_3727);
xor U3856 (N_3856,N_3652,N_3674);
nor U3857 (N_3857,N_3625,N_3606);
and U3858 (N_3858,N_3783,N_3657);
or U3859 (N_3859,N_3798,N_3722);
and U3860 (N_3860,N_3769,N_3683);
or U3861 (N_3861,N_3720,N_3721);
nor U3862 (N_3862,N_3634,N_3633);
and U3863 (N_3863,N_3799,N_3770);
xor U3864 (N_3864,N_3680,N_3789);
or U3865 (N_3865,N_3610,N_3615);
and U3866 (N_3866,N_3786,N_3648);
nand U3867 (N_3867,N_3690,N_3601);
and U3868 (N_3868,N_3671,N_3735);
nor U3869 (N_3869,N_3656,N_3604);
nand U3870 (N_3870,N_3691,N_3699);
nor U3871 (N_3871,N_3697,N_3768);
nor U3872 (N_3872,N_3612,N_3602);
nand U3873 (N_3873,N_3696,N_3647);
nor U3874 (N_3874,N_3705,N_3704);
and U3875 (N_3875,N_3773,N_3668);
nor U3876 (N_3876,N_3732,N_3660);
xnor U3877 (N_3877,N_3726,N_3636);
nor U3878 (N_3878,N_3753,N_3728);
or U3879 (N_3879,N_3737,N_3608);
nor U3880 (N_3880,N_3646,N_3667);
xor U3881 (N_3881,N_3661,N_3618);
nand U3882 (N_3882,N_3616,N_3777);
xnor U3883 (N_3883,N_3710,N_3666);
or U3884 (N_3884,N_3613,N_3701);
or U3885 (N_3885,N_3790,N_3664);
or U3886 (N_3886,N_3645,N_3669);
or U3887 (N_3887,N_3676,N_3771);
and U3888 (N_3888,N_3644,N_3605);
nand U3889 (N_3889,N_3715,N_3778);
and U3890 (N_3890,N_3797,N_3716);
xor U3891 (N_3891,N_3781,N_3659);
or U3892 (N_3892,N_3743,N_3708);
nand U3893 (N_3893,N_3711,N_3673);
nand U3894 (N_3894,N_3686,N_3787);
or U3895 (N_3895,N_3617,N_3619);
nor U3896 (N_3896,N_3620,N_3693);
nor U3897 (N_3897,N_3672,N_3793);
nor U3898 (N_3898,N_3658,N_3635);
xnor U3899 (N_3899,N_3637,N_3765);
nor U3900 (N_3900,N_3688,N_3673);
and U3901 (N_3901,N_3694,N_3742);
or U3902 (N_3902,N_3705,N_3732);
xnor U3903 (N_3903,N_3767,N_3685);
nand U3904 (N_3904,N_3784,N_3616);
nor U3905 (N_3905,N_3746,N_3734);
xnor U3906 (N_3906,N_3666,N_3689);
nor U3907 (N_3907,N_3742,N_3647);
or U3908 (N_3908,N_3616,N_3682);
and U3909 (N_3909,N_3606,N_3697);
nand U3910 (N_3910,N_3784,N_3631);
nand U3911 (N_3911,N_3787,N_3744);
or U3912 (N_3912,N_3754,N_3716);
and U3913 (N_3913,N_3661,N_3615);
nand U3914 (N_3914,N_3655,N_3698);
nor U3915 (N_3915,N_3771,N_3715);
nand U3916 (N_3916,N_3673,N_3685);
nor U3917 (N_3917,N_3733,N_3667);
nor U3918 (N_3918,N_3779,N_3686);
xor U3919 (N_3919,N_3781,N_3729);
nand U3920 (N_3920,N_3736,N_3718);
nand U3921 (N_3921,N_3772,N_3696);
and U3922 (N_3922,N_3656,N_3679);
nor U3923 (N_3923,N_3777,N_3682);
nand U3924 (N_3924,N_3790,N_3643);
nor U3925 (N_3925,N_3626,N_3623);
and U3926 (N_3926,N_3787,N_3723);
xor U3927 (N_3927,N_3668,N_3666);
nor U3928 (N_3928,N_3606,N_3687);
and U3929 (N_3929,N_3755,N_3667);
or U3930 (N_3930,N_3694,N_3631);
nand U3931 (N_3931,N_3671,N_3726);
nor U3932 (N_3932,N_3650,N_3733);
nor U3933 (N_3933,N_3733,N_3744);
and U3934 (N_3934,N_3693,N_3642);
or U3935 (N_3935,N_3686,N_3753);
and U3936 (N_3936,N_3644,N_3789);
or U3937 (N_3937,N_3680,N_3783);
and U3938 (N_3938,N_3696,N_3717);
and U3939 (N_3939,N_3771,N_3779);
nor U3940 (N_3940,N_3620,N_3719);
or U3941 (N_3941,N_3722,N_3671);
nand U3942 (N_3942,N_3735,N_3792);
nor U3943 (N_3943,N_3771,N_3756);
nand U3944 (N_3944,N_3605,N_3772);
xor U3945 (N_3945,N_3792,N_3633);
and U3946 (N_3946,N_3770,N_3689);
or U3947 (N_3947,N_3646,N_3721);
and U3948 (N_3948,N_3676,N_3759);
or U3949 (N_3949,N_3617,N_3607);
nor U3950 (N_3950,N_3732,N_3739);
nand U3951 (N_3951,N_3740,N_3692);
and U3952 (N_3952,N_3640,N_3602);
nor U3953 (N_3953,N_3643,N_3698);
nor U3954 (N_3954,N_3720,N_3785);
xor U3955 (N_3955,N_3649,N_3651);
and U3956 (N_3956,N_3706,N_3775);
nor U3957 (N_3957,N_3729,N_3633);
nor U3958 (N_3958,N_3775,N_3668);
xor U3959 (N_3959,N_3638,N_3773);
nand U3960 (N_3960,N_3769,N_3776);
nor U3961 (N_3961,N_3653,N_3609);
nor U3962 (N_3962,N_3791,N_3611);
nor U3963 (N_3963,N_3725,N_3693);
nor U3964 (N_3964,N_3649,N_3659);
nor U3965 (N_3965,N_3616,N_3704);
or U3966 (N_3966,N_3757,N_3619);
and U3967 (N_3967,N_3668,N_3746);
and U3968 (N_3968,N_3631,N_3707);
xnor U3969 (N_3969,N_3639,N_3634);
xnor U3970 (N_3970,N_3622,N_3608);
and U3971 (N_3971,N_3610,N_3729);
nor U3972 (N_3972,N_3734,N_3621);
and U3973 (N_3973,N_3689,N_3778);
and U3974 (N_3974,N_3754,N_3764);
xor U3975 (N_3975,N_3743,N_3707);
and U3976 (N_3976,N_3795,N_3684);
nand U3977 (N_3977,N_3623,N_3797);
nor U3978 (N_3978,N_3722,N_3745);
or U3979 (N_3979,N_3666,N_3698);
or U3980 (N_3980,N_3681,N_3617);
nor U3981 (N_3981,N_3671,N_3728);
nand U3982 (N_3982,N_3778,N_3608);
nor U3983 (N_3983,N_3776,N_3601);
nand U3984 (N_3984,N_3626,N_3767);
nand U3985 (N_3985,N_3774,N_3684);
or U3986 (N_3986,N_3643,N_3759);
nor U3987 (N_3987,N_3629,N_3644);
or U3988 (N_3988,N_3649,N_3755);
or U3989 (N_3989,N_3623,N_3633);
or U3990 (N_3990,N_3621,N_3615);
and U3991 (N_3991,N_3676,N_3632);
nand U3992 (N_3992,N_3795,N_3779);
nand U3993 (N_3993,N_3601,N_3664);
nand U3994 (N_3994,N_3639,N_3706);
or U3995 (N_3995,N_3609,N_3700);
nor U3996 (N_3996,N_3735,N_3688);
or U3997 (N_3997,N_3684,N_3664);
and U3998 (N_3998,N_3648,N_3675);
nor U3999 (N_3999,N_3615,N_3731);
xnor U4000 (N_4000,N_3939,N_3825);
nand U4001 (N_4001,N_3852,N_3897);
nor U4002 (N_4002,N_3883,N_3966);
xor U4003 (N_4003,N_3962,N_3974);
nand U4004 (N_4004,N_3955,N_3860);
or U4005 (N_4005,N_3877,N_3970);
nor U4006 (N_4006,N_3922,N_3906);
or U4007 (N_4007,N_3928,N_3868);
and U4008 (N_4008,N_3921,N_3943);
nor U4009 (N_4009,N_3808,N_3947);
and U4010 (N_4010,N_3936,N_3926);
xor U4011 (N_4011,N_3836,N_3875);
nor U4012 (N_4012,N_3944,N_3803);
nor U4013 (N_4013,N_3923,N_3824);
nor U4014 (N_4014,N_3841,N_3855);
xor U4015 (N_4015,N_3806,N_3804);
or U4016 (N_4016,N_3994,N_3931);
or U4017 (N_4017,N_3916,N_3827);
and U4018 (N_4018,N_3905,N_3859);
or U4019 (N_4019,N_3961,N_3856);
or U4020 (N_4020,N_3832,N_3898);
or U4021 (N_4021,N_3862,N_3821);
or U4022 (N_4022,N_3951,N_3918);
and U4023 (N_4023,N_3884,N_3880);
nand U4024 (N_4024,N_3828,N_3982);
nand U4025 (N_4025,N_3989,N_3847);
nand U4026 (N_4026,N_3935,N_3963);
nand U4027 (N_4027,N_3829,N_3911);
or U4028 (N_4028,N_3891,N_3991);
or U4029 (N_4029,N_3849,N_3844);
or U4030 (N_4030,N_3919,N_3881);
and U4031 (N_4031,N_3810,N_3975);
or U4032 (N_4032,N_3950,N_3822);
nand U4033 (N_4033,N_3997,N_3899);
xor U4034 (N_4034,N_3959,N_3873);
xnor U4035 (N_4035,N_3814,N_3861);
nand U4036 (N_4036,N_3909,N_3858);
or U4037 (N_4037,N_3826,N_3996);
nor U4038 (N_4038,N_3917,N_3887);
nor U4039 (N_4039,N_3937,N_3864);
and U4040 (N_4040,N_3817,N_3967);
nand U4041 (N_4041,N_3910,N_3818);
nand U4042 (N_4042,N_3846,N_3851);
or U4043 (N_4043,N_3995,N_3903);
or U4044 (N_4044,N_3807,N_3964);
nand U4045 (N_4045,N_3865,N_3908);
nor U4046 (N_4046,N_3973,N_3972);
and U4047 (N_4047,N_3956,N_3907);
or U4048 (N_4048,N_3889,N_3820);
nand U4049 (N_4049,N_3998,N_3977);
nand U4050 (N_4050,N_3968,N_3914);
or U4051 (N_4051,N_3981,N_3870);
nor U4052 (N_4052,N_3850,N_3954);
and U4053 (N_4053,N_3815,N_3837);
or U4054 (N_4054,N_3900,N_3894);
or U4055 (N_4055,N_3801,N_3871);
xor U4056 (N_4056,N_3854,N_3800);
nor U4057 (N_4057,N_3857,N_3863);
xnor U4058 (N_4058,N_3893,N_3874);
and U4059 (N_4059,N_3838,N_3969);
xor U4060 (N_4060,N_3942,N_3872);
nor U4061 (N_4061,N_3915,N_3979);
nand U4062 (N_4062,N_3882,N_3888);
nand U4063 (N_4063,N_3960,N_3802);
nor U4064 (N_4064,N_3992,N_3990);
xnor U4065 (N_4065,N_3987,N_3833);
nand U4066 (N_4066,N_3843,N_3924);
nand U4067 (N_4067,N_3890,N_3819);
nand U4068 (N_4068,N_3830,N_3834);
nor U4069 (N_4069,N_3980,N_3886);
and U4070 (N_4070,N_3876,N_3848);
xnor U4071 (N_4071,N_3985,N_3938);
and U4072 (N_4072,N_3971,N_3993);
nor U4073 (N_4073,N_3945,N_3983);
xor U4074 (N_4074,N_3927,N_3999);
nand U4075 (N_4075,N_3816,N_3984);
nand U4076 (N_4076,N_3813,N_3958);
and U4077 (N_4077,N_3934,N_3831);
nor U4078 (N_4078,N_3840,N_3940);
nand U4079 (N_4079,N_3948,N_3866);
nand U4080 (N_4080,N_3913,N_3952);
nand U4081 (N_4081,N_3941,N_3845);
nand U4082 (N_4082,N_3929,N_3895);
or U4083 (N_4083,N_3853,N_3812);
and U4084 (N_4084,N_3885,N_3811);
nor U4085 (N_4085,N_3878,N_3932);
nor U4086 (N_4086,N_3879,N_3869);
and U4087 (N_4087,N_3835,N_3933);
or U4088 (N_4088,N_3930,N_3957);
or U4089 (N_4089,N_3867,N_3842);
and U4090 (N_4090,N_3976,N_3946);
or U4091 (N_4091,N_3839,N_3892);
nand U4092 (N_4092,N_3920,N_3986);
or U4093 (N_4093,N_3925,N_3949);
or U4094 (N_4094,N_3805,N_3953);
nor U4095 (N_4095,N_3904,N_3901);
or U4096 (N_4096,N_3912,N_3965);
xor U4097 (N_4097,N_3902,N_3896);
xnor U4098 (N_4098,N_3823,N_3988);
and U4099 (N_4099,N_3809,N_3978);
nand U4100 (N_4100,N_3940,N_3947);
and U4101 (N_4101,N_3884,N_3923);
nand U4102 (N_4102,N_3995,N_3877);
nand U4103 (N_4103,N_3929,N_3837);
nand U4104 (N_4104,N_3940,N_3926);
nor U4105 (N_4105,N_3945,N_3985);
and U4106 (N_4106,N_3992,N_3865);
nand U4107 (N_4107,N_3899,N_3864);
or U4108 (N_4108,N_3861,N_3956);
nor U4109 (N_4109,N_3998,N_3890);
nand U4110 (N_4110,N_3890,N_3996);
nand U4111 (N_4111,N_3856,N_3909);
or U4112 (N_4112,N_3818,N_3986);
nand U4113 (N_4113,N_3931,N_3979);
and U4114 (N_4114,N_3972,N_3800);
nor U4115 (N_4115,N_3818,N_3800);
nor U4116 (N_4116,N_3967,N_3802);
nor U4117 (N_4117,N_3875,N_3951);
and U4118 (N_4118,N_3963,N_3876);
and U4119 (N_4119,N_3899,N_3966);
and U4120 (N_4120,N_3992,N_3946);
and U4121 (N_4121,N_3914,N_3910);
xor U4122 (N_4122,N_3911,N_3856);
nand U4123 (N_4123,N_3857,N_3952);
and U4124 (N_4124,N_3809,N_3863);
xnor U4125 (N_4125,N_3935,N_3893);
or U4126 (N_4126,N_3896,N_3840);
or U4127 (N_4127,N_3822,N_3867);
xor U4128 (N_4128,N_3924,N_3811);
nand U4129 (N_4129,N_3931,N_3980);
and U4130 (N_4130,N_3936,N_3873);
or U4131 (N_4131,N_3986,N_3983);
or U4132 (N_4132,N_3970,N_3903);
or U4133 (N_4133,N_3945,N_3953);
and U4134 (N_4134,N_3946,N_3895);
or U4135 (N_4135,N_3940,N_3993);
nand U4136 (N_4136,N_3859,N_3846);
or U4137 (N_4137,N_3846,N_3943);
nand U4138 (N_4138,N_3808,N_3800);
and U4139 (N_4139,N_3815,N_3992);
xnor U4140 (N_4140,N_3880,N_3932);
and U4141 (N_4141,N_3930,N_3986);
nor U4142 (N_4142,N_3960,N_3825);
or U4143 (N_4143,N_3938,N_3856);
or U4144 (N_4144,N_3953,N_3827);
nor U4145 (N_4145,N_3954,N_3974);
and U4146 (N_4146,N_3876,N_3817);
and U4147 (N_4147,N_3885,N_3883);
or U4148 (N_4148,N_3893,N_3866);
nand U4149 (N_4149,N_3808,N_3861);
or U4150 (N_4150,N_3852,N_3842);
or U4151 (N_4151,N_3939,N_3951);
xor U4152 (N_4152,N_3945,N_3984);
or U4153 (N_4153,N_3841,N_3830);
xor U4154 (N_4154,N_3954,N_3976);
or U4155 (N_4155,N_3815,N_3871);
and U4156 (N_4156,N_3838,N_3953);
nand U4157 (N_4157,N_3938,N_3874);
and U4158 (N_4158,N_3845,N_3981);
and U4159 (N_4159,N_3958,N_3932);
and U4160 (N_4160,N_3834,N_3947);
nand U4161 (N_4161,N_3936,N_3858);
nor U4162 (N_4162,N_3976,N_3923);
or U4163 (N_4163,N_3896,N_3885);
xnor U4164 (N_4164,N_3930,N_3822);
xor U4165 (N_4165,N_3872,N_3931);
nand U4166 (N_4166,N_3996,N_3948);
nor U4167 (N_4167,N_3826,N_3879);
or U4168 (N_4168,N_3877,N_3845);
xor U4169 (N_4169,N_3826,N_3975);
xnor U4170 (N_4170,N_3897,N_3995);
and U4171 (N_4171,N_3996,N_3984);
and U4172 (N_4172,N_3842,N_3935);
or U4173 (N_4173,N_3987,N_3955);
nor U4174 (N_4174,N_3899,N_3885);
or U4175 (N_4175,N_3810,N_3900);
nor U4176 (N_4176,N_3804,N_3867);
nand U4177 (N_4177,N_3928,N_3934);
or U4178 (N_4178,N_3934,N_3915);
or U4179 (N_4179,N_3809,N_3902);
nand U4180 (N_4180,N_3965,N_3956);
nand U4181 (N_4181,N_3923,N_3867);
nor U4182 (N_4182,N_3820,N_3957);
or U4183 (N_4183,N_3927,N_3892);
or U4184 (N_4184,N_3914,N_3949);
xor U4185 (N_4185,N_3878,N_3875);
and U4186 (N_4186,N_3811,N_3809);
nand U4187 (N_4187,N_3841,N_3984);
and U4188 (N_4188,N_3943,N_3910);
or U4189 (N_4189,N_3812,N_3955);
nor U4190 (N_4190,N_3929,N_3834);
and U4191 (N_4191,N_3803,N_3830);
and U4192 (N_4192,N_3821,N_3873);
xnor U4193 (N_4193,N_3911,N_3946);
and U4194 (N_4194,N_3971,N_3863);
xnor U4195 (N_4195,N_3844,N_3856);
nor U4196 (N_4196,N_3816,N_3971);
nor U4197 (N_4197,N_3896,N_3800);
and U4198 (N_4198,N_3870,N_3931);
xnor U4199 (N_4199,N_3919,N_3802);
nand U4200 (N_4200,N_4182,N_4195);
xor U4201 (N_4201,N_4095,N_4157);
xor U4202 (N_4202,N_4057,N_4076);
nor U4203 (N_4203,N_4001,N_4176);
nor U4204 (N_4204,N_4169,N_4102);
and U4205 (N_4205,N_4135,N_4181);
and U4206 (N_4206,N_4144,N_4131);
or U4207 (N_4207,N_4086,N_4140);
nand U4208 (N_4208,N_4036,N_4160);
nor U4209 (N_4209,N_4198,N_4089);
and U4210 (N_4210,N_4109,N_4009);
nand U4211 (N_4211,N_4012,N_4165);
nor U4212 (N_4212,N_4087,N_4013);
nor U4213 (N_4213,N_4055,N_4024);
or U4214 (N_4214,N_4121,N_4171);
nor U4215 (N_4215,N_4143,N_4004);
xnor U4216 (N_4216,N_4032,N_4052);
nand U4217 (N_4217,N_4005,N_4147);
and U4218 (N_4218,N_4120,N_4007);
nand U4219 (N_4219,N_4138,N_4065);
and U4220 (N_4220,N_4041,N_4038);
nor U4221 (N_4221,N_4101,N_4134);
or U4222 (N_4222,N_4019,N_4119);
nor U4223 (N_4223,N_4022,N_4092);
and U4224 (N_4224,N_4063,N_4192);
xnor U4225 (N_4225,N_4015,N_4100);
and U4226 (N_4226,N_4110,N_4081);
nor U4227 (N_4227,N_4096,N_4163);
nand U4228 (N_4228,N_4193,N_4028);
nand U4229 (N_4229,N_4091,N_4014);
and U4230 (N_4230,N_4117,N_4021);
xor U4231 (N_4231,N_4060,N_4061);
xnor U4232 (N_4232,N_4035,N_4141);
or U4233 (N_4233,N_4187,N_4085);
and U4234 (N_4234,N_4072,N_4127);
or U4235 (N_4235,N_4034,N_4067);
and U4236 (N_4236,N_4166,N_4040);
nor U4237 (N_4237,N_4175,N_4045);
and U4238 (N_4238,N_4106,N_4158);
or U4239 (N_4239,N_4044,N_4118);
nand U4240 (N_4240,N_4130,N_4042);
xnor U4241 (N_4241,N_4185,N_4070);
nand U4242 (N_4242,N_4133,N_4008);
or U4243 (N_4243,N_4199,N_4029);
or U4244 (N_4244,N_4173,N_4184);
and U4245 (N_4245,N_4016,N_4071);
or U4246 (N_4246,N_4142,N_4030);
nor U4247 (N_4247,N_4050,N_4159);
or U4248 (N_4248,N_4105,N_4123);
and U4249 (N_4249,N_4126,N_4053);
nand U4250 (N_4250,N_4078,N_4162);
nand U4251 (N_4251,N_4116,N_4124);
nand U4252 (N_4252,N_4046,N_4064);
xor U4253 (N_4253,N_4066,N_4049);
or U4254 (N_4254,N_4114,N_4167);
and U4255 (N_4255,N_4023,N_4002);
nand U4256 (N_4256,N_4068,N_4088);
nor U4257 (N_4257,N_4098,N_4062);
xnor U4258 (N_4258,N_4168,N_4020);
nor U4259 (N_4259,N_4018,N_4103);
or U4260 (N_4260,N_4025,N_4075);
or U4261 (N_4261,N_4097,N_4190);
xnor U4262 (N_4262,N_4188,N_4073);
and U4263 (N_4263,N_4145,N_4149);
nor U4264 (N_4264,N_4189,N_4139);
or U4265 (N_4265,N_4113,N_4197);
or U4266 (N_4266,N_4054,N_4154);
or U4267 (N_4267,N_4058,N_4152);
nand U4268 (N_4268,N_4172,N_4153);
and U4269 (N_4269,N_4177,N_4079);
or U4270 (N_4270,N_4136,N_4122);
nor U4271 (N_4271,N_4137,N_4074);
nor U4272 (N_4272,N_4115,N_4011);
or U4273 (N_4273,N_4128,N_4170);
or U4274 (N_4274,N_4069,N_4183);
nor U4275 (N_4275,N_4056,N_4174);
or U4276 (N_4276,N_4082,N_4047);
and U4277 (N_4277,N_4010,N_4051);
and U4278 (N_4278,N_4039,N_4108);
and U4279 (N_4279,N_4148,N_4099);
and U4280 (N_4280,N_4083,N_4006);
or U4281 (N_4281,N_4093,N_4196);
or U4282 (N_4282,N_4129,N_4178);
and U4283 (N_4283,N_4080,N_4027);
xnor U4284 (N_4284,N_4179,N_4107);
nand U4285 (N_4285,N_4017,N_4094);
and U4286 (N_4286,N_4161,N_4003);
and U4287 (N_4287,N_4132,N_4186);
or U4288 (N_4288,N_4146,N_4090);
nand U4289 (N_4289,N_4164,N_4150);
nand U4290 (N_4290,N_4048,N_4033);
nand U4291 (N_4291,N_4037,N_4000);
nand U4292 (N_4292,N_4031,N_4077);
nor U4293 (N_4293,N_4155,N_4125);
nand U4294 (N_4294,N_4156,N_4191);
or U4295 (N_4295,N_4059,N_4104);
xor U4296 (N_4296,N_4084,N_4180);
or U4297 (N_4297,N_4112,N_4043);
and U4298 (N_4298,N_4111,N_4194);
and U4299 (N_4299,N_4151,N_4026);
nor U4300 (N_4300,N_4053,N_4030);
xnor U4301 (N_4301,N_4039,N_4080);
nor U4302 (N_4302,N_4154,N_4084);
nand U4303 (N_4303,N_4034,N_4050);
or U4304 (N_4304,N_4006,N_4140);
or U4305 (N_4305,N_4092,N_4153);
or U4306 (N_4306,N_4001,N_4008);
nand U4307 (N_4307,N_4145,N_4047);
or U4308 (N_4308,N_4114,N_4004);
or U4309 (N_4309,N_4157,N_4130);
and U4310 (N_4310,N_4043,N_4141);
nor U4311 (N_4311,N_4191,N_4149);
nor U4312 (N_4312,N_4006,N_4195);
nand U4313 (N_4313,N_4132,N_4143);
or U4314 (N_4314,N_4128,N_4143);
or U4315 (N_4315,N_4075,N_4198);
and U4316 (N_4316,N_4023,N_4057);
xnor U4317 (N_4317,N_4092,N_4023);
xnor U4318 (N_4318,N_4099,N_4009);
nand U4319 (N_4319,N_4087,N_4141);
and U4320 (N_4320,N_4049,N_4008);
nand U4321 (N_4321,N_4146,N_4087);
nand U4322 (N_4322,N_4183,N_4041);
nand U4323 (N_4323,N_4177,N_4004);
and U4324 (N_4324,N_4118,N_4176);
nor U4325 (N_4325,N_4167,N_4056);
nand U4326 (N_4326,N_4169,N_4054);
xnor U4327 (N_4327,N_4143,N_4043);
or U4328 (N_4328,N_4191,N_4028);
or U4329 (N_4329,N_4104,N_4067);
nand U4330 (N_4330,N_4040,N_4031);
xor U4331 (N_4331,N_4044,N_4092);
and U4332 (N_4332,N_4177,N_4014);
and U4333 (N_4333,N_4074,N_4007);
nand U4334 (N_4334,N_4006,N_4183);
or U4335 (N_4335,N_4173,N_4118);
xor U4336 (N_4336,N_4005,N_4160);
nor U4337 (N_4337,N_4069,N_4019);
nor U4338 (N_4338,N_4095,N_4025);
and U4339 (N_4339,N_4141,N_4060);
nor U4340 (N_4340,N_4124,N_4178);
nand U4341 (N_4341,N_4036,N_4073);
nand U4342 (N_4342,N_4096,N_4199);
nand U4343 (N_4343,N_4195,N_4147);
or U4344 (N_4344,N_4146,N_4151);
and U4345 (N_4345,N_4006,N_4096);
nand U4346 (N_4346,N_4163,N_4133);
xor U4347 (N_4347,N_4053,N_4152);
or U4348 (N_4348,N_4103,N_4162);
or U4349 (N_4349,N_4017,N_4161);
and U4350 (N_4350,N_4198,N_4070);
xor U4351 (N_4351,N_4182,N_4001);
or U4352 (N_4352,N_4108,N_4027);
nand U4353 (N_4353,N_4081,N_4189);
and U4354 (N_4354,N_4134,N_4007);
and U4355 (N_4355,N_4199,N_4054);
nand U4356 (N_4356,N_4090,N_4005);
and U4357 (N_4357,N_4060,N_4092);
and U4358 (N_4358,N_4045,N_4002);
nand U4359 (N_4359,N_4102,N_4160);
nor U4360 (N_4360,N_4159,N_4177);
or U4361 (N_4361,N_4136,N_4058);
nor U4362 (N_4362,N_4196,N_4121);
nand U4363 (N_4363,N_4090,N_4085);
and U4364 (N_4364,N_4133,N_4063);
nand U4365 (N_4365,N_4087,N_4088);
nor U4366 (N_4366,N_4047,N_4028);
nand U4367 (N_4367,N_4098,N_4055);
nor U4368 (N_4368,N_4176,N_4134);
or U4369 (N_4369,N_4179,N_4073);
xnor U4370 (N_4370,N_4124,N_4073);
nand U4371 (N_4371,N_4086,N_4012);
and U4372 (N_4372,N_4007,N_4031);
nor U4373 (N_4373,N_4161,N_4141);
nand U4374 (N_4374,N_4119,N_4048);
nand U4375 (N_4375,N_4009,N_4158);
nor U4376 (N_4376,N_4012,N_4069);
nor U4377 (N_4377,N_4059,N_4193);
nor U4378 (N_4378,N_4019,N_4011);
or U4379 (N_4379,N_4172,N_4035);
nor U4380 (N_4380,N_4047,N_4128);
and U4381 (N_4381,N_4083,N_4192);
nor U4382 (N_4382,N_4013,N_4062);
nand U4383 (N_4383,N_4054,N_4001);
nor U4384 (N_4384,N_4183,N_4025);
nand U4385 (N_4385,N_4195,N_4070);
and U4386 (N_4386,N_4119,N_4070);
or U4387 (N_4387,N_4028,N_4013);
nand U4388 (N_4388,N_4051,N_4197);
nand U4389 (N_4389,N_4131,N_4062);
nor U4390 (N_4390,N_4048,N_4181);
or U4391 (N_4391,N_4170,N_4121);
xnor U4392 (N_4392,N_4037,N_4120);
and U4393 (N_4393,N_4037,N_4163);
xor U4394 (N_4394,N_4093,N_4112);
xnor U4395 (N_4395,N_4102,N_4101);
nand U4396 (N_4396,N_4171,N_4156);
and U4397 (N_4397,N_4104,N_4113);
nand U4398 (N_4398,N_4179,N_4042);
or U4399 (N_4399,N_4047,N_4095);
xnor U4400 (N_4400,N_4262,N_4303);
nand U4401 (N_4401,N_4286,N_4231);
nor U4402 (N_4402,N_4397,N_4298);
or U4403 (N_4403,N_4355,N_4240);
or U4404 (N_4404,N_4249,N_4315);
or U4405 (N_4405,N_4297,N_4385);
nand U4406 (N_4406,N_4273,N_4274);
xnor U4407 (N_4407,N_4346,N_4311);
and U4408 (N_4408,N_4215,N_4388);
nor U4409 (N_4409,N_4328,N_4370);
or U4410 (N_4410,N_4381,N_4225);
nand U4411 (N_4411,N_4335,N_4205);
nand U4412 (N_4412,N_4354,N_4226);
and U4413 (N_4413,N_4280,N_4258);
or U4414 (N_4414,N_4253,N_4259);
nand U4415 (N_4415,N_4268,N_4221);
or U4416 (N_4416,N_4382,N_4372);
nor U4417 (N_4417,N_4317,N_4306);
and U4418 (N_4418,N_4344,N_4362);
or U4419 (N_4419,N_4348,N_4284);
and U4420 (N_4420,N_4389,N_4236);
and U4421 (N_4421,N_4237,N_4364);
and U4422 (N_4422,N_4287,N_4216);
nand U4423 (N_4423,N_4230,N_4310);
or U4424 (N_4424,N_4209,N_4363);
and U4425 (N_4425,N_4368,N_4282);
and U4426 (N_4426,N_4392,N_4265);
nand U4427 (N_4427,N_4279,N_4341);
nand U4428 (N_4428,N_4312,N_4386);
or U4429 (N_4429,N_4380,N_4203);
and U4430 (N_4430,N_4396,N_4260);
and U4431 (N_4431,N_4376,N_4309);
nor U4432 (N_4432,N_4299,N_4232);
xnor U4433 (N_4433,N_4349,N_4246);
and U4434 (N_4434,N_4339,N_4263);
and U4435 (N_4435,N_4331,N_4296);
nand U4436 (N_4436,N_4242,N_4393);
or U4437 (N_4437,N_4318,N_4308);
and U4438 (N_4438,N_4247,N_4321);
nand U4439 (N_4439,N_4320,N_4357);
and U4440 (N_4440,N_4360,N_4227);
and U4441 (N_4441,N_4300,N_4301);
and U4442 (N_4442,N_4330,N_4379);
nand U4443 (N_4443,N_4342,N_4324);
nor U4444 (N_4444,N_4222,N_4367);
nand U4445 (N_4445,N_4254,N_4238);
nand U4446 (N_4446,N_4234,N_4394);
nand U4447 (N_4447,N_4319,N_4369);
nand U4448 (N_4448,N_4356,N_4275);
xor U4449 (N_4449,N_4395,N_4200);
nand U4450 (N_4450,N_4257,N_4206);
and U4451 (N_4451,N_4314,N_4293);
and U4452 (N_4452,N_4269,N_4289);
nor U4453 (N_4453,N_4340,N_4207);
nand U4454 (N_4454,N_4325,N_4212);
or U4455 (N_4455,N_4345,N_4223);
nor U4456 (N_4456,N_4202,N_4337);
nor U4457 (N_4457,N_4305,N_4307);
nand U4458 (N_4458,N_4229,N_4267);
nand U4459 (N_4459,N_4359,N_4391);
nand U4460 (N_4460,N_4373,N_4220);
or U4461 (N_4461,N_4323,N_4343);
or U4462 (N_4462,N_4375,N_4217);
xor U4463 (N_4463,N_4304,N_4350);
or U4464 (N_4464,N_4250,N_4295);
or U4465 (N_4465,N_4248,N_4384);
nor U4466 (N_4466,N_4288,N_4292);
and U4467 (N_4467,N_4374,N_4351);
and U4468 (N_4468,N_4290,N_4252);
nand U4469 (N_4469,N_4233,N_4239);
nand U4470 (N_4470,N_4329,N_4211);
nor U4471 (N_4471,N_4264,N_4201);
and U4472 (N_4472,N_4285,N_4399);
nand U4473 (N_4473,N_4366,N_4218);
and U4474 (N_4474,N_4358,N_4316);
or U4475 (N_4475,N_4210,N_4302);
or U4476 (N_4476,N_4332,N_4353);
nor U4477 (N_4477,N_4291,N_4228);
nor U4478 (N_4478,N_4322,N_4213);
xor U4479 (N_4479,N_4241,N_4398);
nor U4480 (N_4480,N_4270,N_4333);
nand U4481 (N_4481,N_4387,N_4271);
nand U4482 (N_4482,N_4283,N_4361);
or U4483 (N_4483,N_4272,N_4336);
nand U4484 (N_4484,N_4245,N_4208);
nor U4485 (N_4485,N_4390,N_4378);
nand U4486 (N_4486,N_4214,N_4204);
nand U4487 (N_4487,N_4281,N_4327);
or U4488 (N_4488,N_4371,N_4243);
nand U4489 (N_4489,N_4365,N_4347);
and U4490 (N_4490,N_4266,N_4219);
nor U4491 (N_4491,N_4255,N_4251);
nor U4492 (N_4492,N_4352,N_4377);
nand U4493 (N_4493,N_4278,N_4261);
nor U4494 (N_4494,N_4277,N_4326);
and U4495 (N_4495,N_4276,N_4256);
nand U4496 (N_4496,N_4334,N_4294);
and U4497 (N_4497,N_4235,N_4313);
nand U4498 (N_4498,N_4224,N_4338);
and U4499 (N_4499,N_4244,N_4383);
and U4500 (N_4500,N_4299,N_4217);
or U4501 (N_4501,N_4307,N_4252);
and U4502 (N_4502,N_4394,N_4288);
or U4503 (N_4503,N_4212,N_4257);
nor U4504 (N_4504,N_4291,N_4276);
or U4505 (N_4505,N_4382,N_4275);
and U4506 (N_4506,N_4373,N_4381);
or U4507 (N_4507,N_4258,N_4244);
nor U4508 (N_4508,N_4344,N_4338);
nor U4509 (N_4509,N_4200,N_4286);
or U4510 (N_4510,N_4353,N_4399);
or U4511 (N_4511,N_4394,N_4341);
or U4512 (N_4512,N_4205,N_4394);
nand U4513 (N_4513,N_4368,N_4234);
nand U4514 (N_4514,N_4238,N_4356);
nand U4515 (N_4515,N_4233,N_4323);
nor U4516 (N_4516,N_4326,N_4399);
xnor U4517 (N_4517,N_4363,N_4269);
or U4518 (N_4518,N_4284,N_4246);
xnor U4519 (N_4519,N_4317,N_4260);
or U4520 (N_4520,N_4266,N_4263);
nor U4521 (N_4521,N_4271,N_4261);
or U4522 (N_4522,N_4207,N_4210);
nor U4523 (N_4523,N_4315,N_4261);
or U4524 (N_4524,N_4348,N_4283);
xnor U4525 (N_4525,N_4293,N_4251);
nor U4526 (N_4526,N_4393,N_4248);
and U4527 (N_4527,N_4396,N_4200);
nand U4528 (N_4528,N_4214,N_4341);
nor U4529 (N_4529,N_4339,N_4317);
or U4530 (N_4530,N_4384,N_4292);
and U4531 (N_4531,N_4249,N_4252);
xor U4532 (N_4532,N_4265,N_4313);
and U4533 (N_4533,N_4280,N_4224);
nand U4534 (N_4534,N_4335,N_4268);
or U4535 (N_4535,N_4348,N_4350);
nor U4536 (N_4536,N_4232,N_4251);
nand U4537 (N_4537,N_4348,N_4220);
nor U4538 (N_4538,N_4266,N_4356);
or U4539 (N_4539,N_4287,N_4253);
and U4540 (N_4540,N_4254,N_4244);
nand U4541 (N_4541,N_4332,N_4321);
or U4542 (N_4542,N_4278,N_4351);
or U4543 (N_4543,N_4230,N_4339);
and U4544 (N_4544,N_4234,N_4318);
or U4545 (N_4545,N_4212,N_4346);
and U4546 (N_4546,N_4353,N_4349);
and U4547 (N_4547,N_4393,N_4324);
or U4548 (N_4548,N_4388,N_4211);
nand U4549 (N_4549,N_4320,N_4229);
or U4550 (N_4550,N_4227,N_4365);
xor U4551 (N_4551,N_4369,N_4241);
or U4552 (N_4552,N_4393,N_4383);
nand U4553 (N_4553,N_4248,N_4275);
or U4554 (N_4554,N_4321,N_4239);
or U4555 (N_4555,N_4294,N_4262);
and U4556 (N_4556,N_4375,N_4215);
nand U4557 (N_4557,N_4231,N_4310);
or U4558 (N_4558,N_4277,N_4206);
or U4559 (N_4559,N_4323,N_4284);
nor U4560 (N_4560,N_4399,N_4319);
nand U4561 (N_4561,N_4385,N_4376);
or U4562 (N_4562,N_4329,N_4316);
or U4563 (N_4563,N_4344,N_4392);
nor U4564 (N_4564,N_4254,N_4241);
and U4565 (N_4565,N_4386,N_4286);
or U4566 (N_4566,N_4207,N_4347);
and U4567 (N_4567,N_4226,N_4361);
nor U4568 (N_4568,N_4376,N_4262);
or U4569 (N_4569,N_4221,N_4206);
xnor U4570 (N_4570,N_4337,N_4382);
xnor U4571 (N_4571,N_4200,N_4382);
or U4572 (N_4572,N_4304,N_4278);
and U4573 (N_4573,N_4303,N_4306);
or U4574 (N_4574,N_4335,N_4249);
or U4575 (N_4575,N_4353,N_4207);
and U4576 (N_4576,N_4275,N_4228);
nor U4577 (N_4577,N_4325,N_4231);
xor U4578 (N_4578,N_4230,N_4262);
nand U4579 (N_4579,N_4339,N_4328);
and U4580 (N_4580,N_4360,N_4333);
nand U4581 (N_4581,N_4282,N_4322);
or U4582 (N_4582,N_4382,N_4307);
or U4583 (N_4583,N_4265,N_4285);
nor U4584 (N_4584,N_4387,N_4265);
and U4585 (N_4585,N_4248,N_4276);
or U4586 (N_4586,N_4252,N_4251);
or U4587 (N_4587,N_4383,N_4360);
or U4588 (N_4588,N_4282,N_4274);
or U4589 (N_4589,N_4202,N_4379);
and U4590 (N_4590,N_4309,N_4269);
nand U4591 (N_4591,N_4226,N_4289);
and U4592 (N_4592,N_4266,N_4304);
xor U4593 (N_4593,N_4364,N_4224);
and U4594 (N_4594,N_4349,N_4398);
nand U4595 (N_4595,N_4249,N_4391);
xor U4596 (N_4596,N_4258,N_4221);
nand U4597 (N_4597,N_4268,N_4274);
nand U4598 (N_4598,N_4379,N_4358);
and U4599 (N_4599,N_4371,N_4365);
or U4600 (N_4600,N_4427,N_4595);
or U4601 (N_4601,N_4446,N_4458);
or U4602 (N_4602,N_4429,N_4565);
nor U4603 (N_4603,N_4538,N_4419);
or U4604 (N_4604,N_4477,N_4467);
nand U4605 (N_4605,N_4455,N_4574);
and U4606 (N_4606,N_4556,N_4557);
nand U4607 (N_4607,N_4480,N_4560);
nor U4608 (N_4608,N_4412,N_4451);
nor U4609 (N_4609,N_4562,N_4555);
nor U4610 (N_4610,N_4591,N_4571);
nand U4611 (N_4611,N_4553,N_4402);
nor U4612 (N_4612,N_4434,N_4468);
or U4613 (N_4613,N_4413,N_4541);
nand U4614 (N_4614,N_4437,N_4483);
nand U4615 (N_4615,N_4463,N_4513);
nand U4616 (N_4616,N_4542,N_4425);
and U4617 (N_4617,N_4456,N_4426);
and U4618 (N_4618,N_4523,N_4465);
or U4619 (N_4619,N_4473,N_4487);
or U4620 (N_4620,N_4432,N_4439);
and U4621 (N_4621,N_4423,N_4422);
and U4622 (N_4622,N_4415,N_4593);
or U4623 (N_4623,N_4549,N_4525);
nor U4624 (N_4624,N_4436,N_4433);
nand U4625 (N_4625,N_4494,N_4405);
or U4626 (N_4626,N_4492,N_4497);
nand U4627 (N_4627,N_4502,N_4520);
nand U4628 (N_4628,N_4450,N_4597);
and U4629 (N_4629,N_4469,N_4506);
xor U4630 (N_4630,N_4532,N_4537);
and U4631 (N_4631,N_4596,N_4488);
nand U4632 (N_4632,N_4585,N_4519);
nor U4633 (N_4633,N_4454,N_4536);
xnor U4634 (N_4634,N_4457,N_4576);
or U4635 (N_4635,N_4577,N_4581);
nor U4636 (N_4636,N_4440,N_4448);
nor U4637 (N_4637,N_4543,N_4496);
or U4638 (N_4638,N_4478,N_4526);
and U4639 (N_4639,N_4476,N_4414);
nor U4640 (N_4640,N_4438,N_4512);
and U4641 (N_4641,N_4464,N_4420);
and U4642 (N_4642,N_4548,N_4418);
nand U4643 (N_4643,N_4504,N_4507);
nor U4644 (N_4644,N_4442,N_4407);
nor U4645 (N_4645,N_4550,N_4509);
and U4646 (N_4646,N_4474,N_4529);
nand U4647 (N_4647,N_4599,N_4401);
xnor U4648 (N_4648,N_4499,N_4472);
nor U4649 (N_4649,N_4563,N_4530);
nor U4650 (N_4650,N_4587,N_4447);
or U4651 (N_4651,N_4598,N_4408);
nand U4652 (N_4652,N_4482,N_4424);
nor U4653 (N_4653,N_4475,N_4552);
nand U4654 (N_4654,N_4441,N_4431);
nor U4655 (N_4655,N_4453,N_4570);
nor U4656 (N_4656,N_4489,N_4582);
nor U4657 (N_4657,N_4527,N_4445);
or U4658 (N_4658,N_4522,N_4470);
nor U4659 (N_4659,N_4539,N_4449);
and U4660 (N_4660,N_4462,N_4511);
nor U4661 (N_4661,N_4533,N_4471);
or U4662 (N_4662,N_4421,N_4528);
or U4663 (N_4663,N_4443,N_4569);
or U4664 (N_4664,N_4510,N_4589);
and U4665 (N_4665,N_4564,N_4517);
nand U4666 (N_4666,N_4400,N_4410);
nand U4667 (N_4667,N_4580,N_4579);
and U4668 (N_4668,N_4521,N_4491);
xor U4669 (N_4669,N_4459,N_4505);
nor U4670 (N_4670,N_4561,N_4404);
or U4671 (N_4671,N_4518,N_4594);
and U4672 (N_4672,N_4573,N_4444);
and U4673 (N_4673,N_4551,N_4508);
nand U4674 (N_4674,N_4495,N_4583);
xor U4675 (N_4675,N_4461,N_4409);
nor U4676 (N_4676,N_4411,N_4558);
nand U4677 (N_4677,N_4584,N_4544);
nand U4678 (N_4678,N_4484,N_4590);
and U4679 (N_4679,N_4545,N_4578);
nor U4680 (N_4680,N_4524,N_4416);
or U4681 (N_4681,N_4452,N_4428);
xor U4682 (N_4682,N_4575,N_4479);
xor U4683 (N_4683,N_4430,N_4486);
nor U4684 (N_4684,N_4592,N_4481);
nor U4685 (N_4685,N_4406,N_4466);
xnor U4686 (N_4686,N_4403,N_4586);
xor U4687 (N_4687,N_4588,N_4503);
nor U4688 (N_4688,N_4572,N_4500);
xor U4689 (N_4689,N_4490,N_4559);
and U4690 (N_4690,N_4515,N_4501);
nor U4691 (N_4691,N_4485,N_4514);
nor U4692 (N_4692,N_4534,N_4417);
nor U4693 (N_4693,N_4567,N_4547);
and U4694 (N_4694,N_4516,N_4554);
nand U4695 (N_4695,N_4460,N_4493);
and U4696 (N_4696,N_4546,N_4498);
or U4697 (N_4697,N_4535,N_4568);
xnor U4698 (N_4698,N_4435,N_4540);
nand U4699 (N_4699,N_4566,N_4531);
and U4700 (N_4700,N_4575,N_4416);
nor U4701 (N_4701,N_4527,N_4405);
xnor U4702 (N_4702,N_4575,N_4520);
or U4703 (N_4703,N_4422,N_4575);
nand U4704 (N_4704,N_4402,N_4500);
xor U4705 (N_4705,N_4424,N_4552);
nor U4706 (N_4706,N_4454,N_4481);
xnor U4707 (N_4707,N_4543,N_4501);
nand U4708 (N_4708,N_4500,N_4527);
or U4709 (N_4709,N_4427,N_4574);
and U4710 (N_4710,N_4456,N_4410);
nand U4711 (N_4711,N_4401,N_4496);
nor U4712 (N_4712,N_4530,N_4588);
nand U4713 (N_4713,N_4592,N_4569);
nor U4714 (N_4714,N_4557,N_4497);
and U4715 (N_4715,N_4526,N_4415);
or U4716 (N_4716,N_4559,N_4580);
nor U4717 (N_4717,N_4419,N_4590);
nor U4718 (N_4718,N_4522,N_4594);
nand U4719 (N_4719,N_4435,N_4496);
or U4720 (N_4720,N_4526,N_4406);
and U4721 (N_4721,N_4492,N_4462);
nand U4722 (N_4722,N_4533,N_4535);
nand U4723 (N_4723,N_4540,N_4503);
and U4724 (N_4724,N_4442,N_4516);
nor U4725 (N_4725,N_4496,N_4439);
and U4726 (N_4726,N_4576,N_4529);
and U4727 (N_4727,N_4584,N_4449);
nor U4728 (N_4728,N_4566,N_4501);
nand U4729 (N_4729,N_4545,N_4488);
xor U4730 (N_4730,N_4550,N_4567);
nor U4731 (N_4731,N_4486,N_4533);
and U4732 (N_4732,N_4424,N_4562);
or U4733 (N_4733,N_4591,N_4519);
nand U4734 (N_4734,N_4492,N_4542);
nor U4735 (N_4735,N_4521,N_4578);
and U4736 (N_4736,N_4464,N_4418);
and U4737 (N_4737,N_4458,N_4420);
nand U4738 (N_4738,N_4426,N_4591);
nor U4739 (N_4739,N_4562,N_4539);
or U4740 (N_4740,N_4453,N_4492);
nand U4741 (N_4741,N_4591,N_4558);
or U4742 (N_4742,N_4487,N_4433);
nor U4743 (N_4743,N_4441,N_4590);
nor U4744 (N_4744,N_4537,N_4417);
nor U4745 (N_4745,N_4500,N_4412);
nor U4746 (N_4746,N_4524,N_4512);
nand U4747 (N_4747,N_4568,N_4444);
nand U4748 (N_4748,N_4466,N_4554);
nor U4749 (N_4749,N_4527,N_4523);
and U4750 (N_4750,N_4527,N_4494);
or U4751 (N_4751,N_4507,N_4556);
and U4752 (N_4752,N_4574,N_4505);
and U4753 (N_4753,N_4448,N_4539);
and U4754 (N_4754,N_4477,N_4516);
nor U4755 (N_4755,N_4441,N_4537);
xnor U4756 (N_4756,N_4443,N_4492);
nand U4757 (N_4757,N_4433,N_4547);
or U4758 (N_4758,N_4500,N_4496);
nand U4759 (N_4759,N_4532,N_4538);
nor U4760 (N_4760,N_4430,N_4474);
nor U4761 (N_4761,N_4444,N_4539);
nand U4762 (N_4762,N_4583,N_4530);
nor U4763 (N_4763,N_4595,N_4559);
or U4764 (N_4764,N_4510,N_4519);
nor U4765 (N_4765,N_4402,N_4449);
or U4766 (N_4766,N_4508,N_4498);
and U4767 (N_4767,N_4526,N_4545);
nand U4768 (N_4768,N_4544,N_4449);
or U4769 (N_4769,N_4598,N_4496);
nor U4770 (N_4770,N_4423,N_4457);
or U4771 (N_4771,N_4544,N_4591);
and U4772 (N_4772,N_4577,N_4596);
nor U4773 (N_4773,N_4416,N_4491);
or U4774 (N_4774,N_4428,N_4559);
nand U4775 (N_4775,N_4453,N_4483);
nand U4776 (N_4776,N_4474,N_4579);
xnor U4777 (N_4777,N_4430,N_4472);
or U4778 (N_4778,N_4491,N_4573);
and U4779 (N_4779,N_4502,N_4407);
nand U4780 (N_4780,N_4520,N_4418);
or U4781 (N_4781,N_4518,N_4472);
or U4782 (N_4782,N_4571,N_4451);
nand U4783 (N_4783,N_4408,N_4538);
and U4784 (N_4784,N_4576,N_4519);
nor U4785 (N_4785,N_4509,N_4532);
nor U4786 (N_4786,N_4563,N_4426);
nor U4787 (N_4787,N_4586,N_4592);
and U4788 (N_4788,N_4477,N_4539);
and U4789 (N_4789,N_4467,N_4555);
nand U4790 (N_4790,N_4445,N_4502);
nand U4791 (N_4791,N_4450,N_4451);
nor U4792 (N_4792,N_4406,N_4574);
nor U4793 (N_4793,N_4493,N_4477);
xor U4794 (N_4794,N_4432,N_4561);
and U4795 (N_4795,N_4422,N_4430);
xnor U4796 (N_4796,N_4411,N_4436);
nor U4797 (N_4797,N_4449,N_4421);
or U4798 (N_4798,N_4436,N_4552);
and U4799 (N_4799,N_4500,N_4567);
nor U4800 (N_4800,N_4789,N_4700);
nand U4801 (N_4801,N_4792,N_4723);
or U4802 (N_4802,N_4771,N_4683);
xor U4803 (N_4803,N_4704,N_4641);
nor U4804 (N_4804,N_4712,N_4757);
or U4805 (N_4805,N_4628,N_4664);
nand U4806 (N_4806,N_4740,N_4797);
xnor U4807 (N_4807,N_4629,N_4763);
and U4808 (N_4808,N_4733,N_4752);
nor U4809 (N_4809,N_4724,N_4761);
nor U4810 (N_4810,N_4601,N_4710);
nand U4811 (N_4811,N_4671,N_4748);
nor U4812 (N_4812,N_4637,N_4735);
and U4813 (N_4813,N_4702,N_4624);
nor U4814 (N_4814,N_4619,N_4756);
or U4815 (N_4815,N_4686,N_4753);
and U4816 (N_4816,N_4666,N_4796);
and U4817 (N_4817,N_4726,N_4688);
xor U4818 (N_4818,N_4680,N_4722);
nor U4819 (N_4819,N_4721,N_4694);
nand U4820 (N_4820,N_4685,N_4750);
and U4821 (N_4821,N_4614,N_4747);
nand U4822 (N_4822,N_4741,N_4779);
nor U4823 (N_4823,N_4785,N_4746);
and U4824 (N_4824,N_4784,N_4633);
or U4825 (N_4825,N_4720,N_4703);
or U4826 (N_4826,N_4626,N_4689);
and U4827 (N_4827,N_4657,N_4602);
nor U4828 (N_4828,N_4608,N_4681);
nand U4829 (N_4829,N_4783,N_4714);
nor U4830 (N_4830,N_4701,N_4667);
nand U4831 (N_4831,N_4679,N_4764);
nor U4832 (N_4832,N_4780,N_4794);
nand U4833 (N_4833,N_4618,N_4604);
or U4834 (N_4834,N_4622,N_4744);
nand U4835 (N_4835,N_4661,N_4799);
nor U4836 (N_4836,N_4776,N_4670);
and U4837 (N_4837,N_4616,N_4660);
or U4838 (N_4838,N_4684,N_4692);
or U4839 (N_4839,N_4737,N_4791);
and U4840 (N_4840,N_4715,N_4603);
nand U4841 (N_4841,N_4758,N_4662);
nand U4842 (N_4842,N_4705,N_4690);
or U4843 (N_4843,N_4613,N_4668);
or U4844 (N_4844,N_4609,N_4621);
nor U4845 (N_4845,N_4730,N_4765);
or U4846 (N_4846,N_4650,N_4617);
or U4847 (N_4847,N_4777,N_4658);
nor U4848 (N_4848,N_4638,N_4644);
or U4849 (N_4849,N_4652,N_4787);
nor U4850 (N_4850,N_4646,N_4636);
nor U4851 (N_4851,N_4788,N_4620);
and U4852 (N_4852,N_4699,N_4762);
nor U4853 (N_4853,N_4623,N_4745);
nand U4854 (N_4854,N_4639,N_4647);
nand U4855 (N_4855,N_4768,N_4775);
nor U4856 (N_4856,N_4611,N_4728);
xnor U4857 (N_4857,N_4798,N_4709);
or U4858 (N_4858,N_4736,N_4738);
nor U4859 (N_4859,N_4760,N_4786);
nand U4860 (N_4860,N_4653,N_4790);
and U4861 (N_4861,N_4673,N_4742);
nand U4862 (N_4862,N_4631,N_4600);
and U4863 (N_4863,N_4677,N_4635);
nor U4864 (N_4864,N_4725,N_4642);
nor U4865 (N_4865,N_4610,N_4678);
nand U4866 (N_4866,N_4687,N_4605);
nor U4867 (N_4867,N_4693,N_4732);
nand U4868 (N_4868,N_4612,N_4706);
nor U4869 (N_4869,N_4774,N_4675);
nand U4870 (N_4870,N_4755,N_4691);
nor U4871 (N_4871,N_4734,N_4770);
xor U4872 (N_4872,N_4648,N_4711);
or U4873 (N_4873,N_4698,N_4759);
nand U4874 (N_4874,N_4716,N_4754);
or U4875 (N_4875,N_4766,N_4665);
xnor U4876 (N_4876,N_4729,N_4708);
nand U4877 (N_4877,N_4749,N_4615);
and U4878 (N_4878,N_4773,N_4696);
nor U4879 (N_4879,N_4718,N_4676);
nor U4880 (N_4880,N_4713,N_4731);
or U4881 (N_4881,N_4634,N_4627);
or U4882 (N_4882,N_4649,N_4663);
nor U4883 (N_4883,N_4655,N_4682);
and U4884 (N_4884,N_4606,N_4607);
nand U4885 (N_4885,N_4659,N_4778);
nand U4886 (N_4886,N_4669,N_4625);
nor U4887 (N_4887,N_4769,N_4654);
or U4888 (N_4888,N_4697,N_4632);
nor U4889 (N_4889,N_4656,N_4782);
and U4890 (N_4890,N_4793,N_4707);
nor U4891 (N_4891,N_4695,N_4630);
nand U4892 (N_4892,N_4643,N_4719);
nor U4893 (N_4893,N_4672,N_4739);
xnor U4894 (N_4894,N_4781,N_4674);
nand U4895 (N_4895,N_4767,N_4751);
and U4896 (N_4896,N_4727,N_4743);
and U4897 (N_4897,N_4795,N_4645);
nor U4898 (N_4898,N_4651,N_4772);
and U4899 (N_4899,N_4640,N_4717);
and U4900 (N_4900,N_4640,N_4795);
nor U4901 (N_4901,N_4735,N_4786);
or U4902 (N_4902,N_4664,N_4727);
and U4903 (N_4903,N_4620,N_4680);
and U4904 (N_4904,N_4770,N_4616);
nor U4905 (N_4905,N_4743,N_4636);
or U4906 (N_4906,N_4658,N_4775);
or U4907 (N_4907,N_4788,N_4698);
or U4908 (N_4908,N_4726,N_4750);
and U4909 (N_4909,N_4775,N_4743);
nor U4910 (N_4910,N_4688,N_4698);
nor U4911 (N_4911,N_4600,N_4796);
or U4912 (N_4912,N_4661,N_4678);
and U4913 (N_4913,N_4707,N_4726);
nor U4914 (N_4914,N_4792,N_4783);
or U4915 (N_4915,N_4730,N_4752);
nor U4916 (N_4916,N_4646,N_4680);
and U4917 (N_4917,N_4756,N_4709);
nor U4918 (N_4918,N_4736,N_4705);
or U4919 (N_4919,N_4620,N_4645);
nor U4920 (N_4920,N_4726,N_4737);
nor U4921 (N_4921,N_4775,N_4791);
or U4922 (N_4922,N_4615,N_4699);
or U4923 (N_4923,N_4740,N_4720);
xor U4924 (N_4924,N_4778,N_4791);
nand U4925 (N_4925,N_4794,N_4601);
nand U4926 (N_4926,N_4665,N_4691);
nor U4927 (N_4927,N_4609,N_4769);
and U4928 (N_4928,N_4661,N_4610);
nand U4929 (N_4929,N_4743,N_4746);
nand U4930 (N_4930,N_4737,N_4710);
nand U4931 (N_4931,N_4647,N_4616);
nand U4932 (N_4932,N_4639,N_4760);
or U4933 (N_4933,N_4735,N_4756);
and U4934 (N_4934,N_4603,N_4672);
nor U4935 (N_4935,N_4684,N_4614);
nand U4936 (N_4936,N_4794,N_4730);
xor U4937 (N_4937,N_4708,N_4765);
nor U4938 (N_4938,N_4705,N_4622);
nor U4939 (N_4939,N_4763,N_4686);
and U4940 (N_4940,N_4786,N_4754);
nor U4941 (N_4941,N_4771,N_4743);
nand U4942 (N_4942,N_4710,N_4706);
or U4943 (N_4943,N_4600,N_4681);
or U4944 (N_4944,N_4648,N_4682);
xor U4945 (N_4945,N_4662,N_4776);
nor U4946 (N_4946,N_4635,N_4757);
or U4947 (N_4947,N_4697,N_4714);
and U4948 (N_4948,N_4639,N_4756);
and U4949 (N_4949,N_4701,N_4732);
or U4950 (N_4950,N_4644,N_4730);
xor U4951 (N_4951,N_4600,N_4692);
or U4952 (N_4952,N_4704,N_4697);
xnor U4953 (N_4953,N_4729,N_4657);
nor U4954 (N_4954,N_4631,N_4634);
nor U4955 (N_4955,N_4762,N_4640);
and U4956 (N_4956,N_4749,N_4716);
nand U4957 (N_4957,N_4762,N_4703);
and U4958 (N_4958,N_4615,N_4712);
nor U4959 (N_4959,N_4684,N_4657);
nor U4960 (N_4960,N_4638,N_4724);
and U4961 (N_4961,N_4669,N_4701);
nand U4962 (N_4962,N_4680,N_4609);
nor U4963 (N_4963,N_4739,N_4688);
nor U4964 (N_4964,N_4700,N_4694);
or U4965 (N_4965,N_4614,N_4707);
xnor U4966 (N_4966,N_4611,N_4667);
nor U4967 (N_4967,N_4742,N_4621);
or U4968 (N_4968,N_4782,N_4700);
nand U4969 (N_4969,N_4779,N_4688);
nor U4970 (N_4970,N_4726,N_4788);
or U4971 (N_4971,N_4631,N_4636);
nor U4972 (N_4972,N_4768,N_4714);
and U4973 (N_4973,N_4675,N_4743);
nor U4974 (N_4974,N_4619,N_4674);
nand U4975 (N_4975,N_4718,N_4692);
or U4976 (N_4976,N_4714,N_4610);
nand U4977 (N_4977,N_4761,N_4799);
and U4978 (N_4978,N_4697,N_4673);
and U4979 (N_4979,N_4644,N_4683);
or U4980 (N_4980,N_4666,N_4668);
xor U4981 (N_4981,N_4694,N_4792);
or U4982 (N_4982,N_4656,N_4760);
nor U4983 (N_4983,N_4626,N_4666);
nand U4984 (N_4984,N_4669,N_4764);
nor U4985 (N_4985,N_4798,N_4692);
or U4986 (N_4986,N_4729,N_4618);
xnor U4987 (N_4987,N_4612,N_4781);
and U4988 (N_4988,N_4762,N_4750);
or U4989 (N_4989,N_4782,N_4611);
nand U4990 (N_4990,N_4686,N_4621);
xnor U4991 (N_4991,N_4620,N_4781);
xor U4992 (N_4992,N_4751,N_4747);
and U4993 (N_4993,N_4650,N_4608);
or U4994 (N_4994,N_4758,N_4785);
or U4995 (N_4995,N_4604,N_4710);
and U4996 (N_4996,N_4688,N_4670);
nand U4997 (N_4997,N_4658,N_4600);
nand U4998 (N_4998,N_4650,N_4682);
nor U4999 (N_4999,N_4649,N_4675);
nor U5000 (N_5000,N_4850,N_4984);
nand U5001 (N_5001,N_4953,N_4907);
nor U5002 (N_5002,N_4937,N_4902);
xnor U5003 (N_5003,N_4814,N_4932);
and U5004 (N_5004,N_4912,N_4964);
nand U5005 (N_5005,N_4894,N_4927);
xnor U5006 (N_5006,N_4839,N_4972);
and U5007 (N_5007,N_4891,N_4822);
nand U5008 (N_5008,N_4834,N_4817);
and U5009 (N_5009,N_4826,N_4848);
nor U5010 (N_5010,N_4926,N_4840);
xnor U5011 (N_5011,N_4919,N_4830);
and U5012 (N_5012,N_4829,N_4863);
or U5013 (N_5013,N_4847,N_4955);
nor U5014 (N_5014,N_4924,N_4938);
nor U5015 (N_5015,N_4877,N_4900);
or U5016 (N_5016,N_4857,N_4844);
xnor U5017 (N_5017,N_4883,N_4842);
nor U5018 (N_5018,N_4841,N_4890);
or U5019 (N_5019,N_4983,N_4828);
nand U5020 (N_5020,N_4884,N_4929);
xor U5021 (N_5021,N_4947,N_4946);
or U5022 (N_5022,N_4976,N_4968);
or U5023 (N_5023,N_4978,N_4933);
xor U5024 (N_5024,N_4885,N_4922);
nor U5025 (N_5025,N_4889,N_4951);
nand U5026 (N_5026,N_4981,N_4806);
nor U5027 (N_5027,N_4990,N_4905);
nand U5028 (N_5028,N_4893,N_4858);
or U5029 (N_5029,N_4918,N_4813);
nor U5030 (N_5030,N_4914,N_4895);
and U5031 (N_5031,N_4838,N_4899);
and U5032 (N_5032,N_4939,N_4818);
or U5033 (N_5033,N_4974,N_4872);
nand U5034 (N_5034,N_4945,N_4888);
and U5035 (N_5035,N_4908,N_4961);
nand U5036 (N_5036,N_4851,N_4920);
nand U5037 (N_5037,N_4879,N_4915);
and U5038 (N_5038,N_4835,N_4913);
nand U5039 (N_5039,N_4950,N_4956);
nor U5040 (N_5040,N_4831,N_4959);
and U5041 (N_5041,N_4896,N_4866);
or U5042 (N_5042,N_4948,N_4910);
nand U5043 (N_5043,N_4874,N_4960);
or U5044 (N_5044,N_4800,N_4886);
and U5045 (N_5045,N_4986,N_4864);
xnor U5046 (N_5046,N_4867,N_4827);
and U5047 (N_5047,N_4940,N_4821);
nand U5048 (N_5048,N_4909,N_4965);
nor U5049 (N_5049,N_4837,N_4871);
or U5050 (N_5050,N_4811,N_4878);
or U5051 (N_5051,N_4943,N_4931);
or U5052 (N_5052,N_4917,N_4944);
nor U5053 (N_5053,N_4880,N_4941);
and U5054 (N_5054,N_4928,N_4936);
and U5055 (N_5055,N_4952,N_4954);
and U5056 (N_5056,N_4985,N_4816);
nand U5057 (N_5057,N_4824,N_4916);
or U5058 (N_5058,N_4865,N_4906);
nor U5059 (N_5059,N_4875,N_4805);
nand U5060 (N_5060,N_4833,N_4998);
and U5061 (N_5061,N_4809,N_4819);
nor U5062 (N_5062,N_4855,N_4854);
nand U5063 (N_5063,N_4949,N_4987);
or U5064 (N_5064,N_4992,N_4887);
nand U5065 (N_5065,N_4815,N_4958);
xor U5066 (N_5066,N_4963,N_4930);
nand U5067 (N_5067,N_4832,N_4966);
xor U5068 (N_5068,N_4923,N_4808);
nor U5069 (N_5069,N_4971,N_4970);
nor U5070 (N_5070,N_4861,N_4802);
nand U5071 (N_5071,N_4846,N_4820);
and U5072 (N_5072,N_4934,N_4935);
or U5073 (N_5073,N_4810,N_4942);
and U5074 (N_5074,N_4973,N_4999);
and U5075 (N_5075,N_4925,N_4882);
nand U5076 (N_5076,N_4993,N_4969);
and U5077 (N_5077,N_4996,N_4921);
and U5078 (N_5078,N_4904,N_4823);
and U5079 (N_5079,N_4967,N_4991);
or U5080 (N_5080,N_4997,N_4898);
nor U5081 (N_5081,N_4836,N_4980);
nor U5082 (N_5082,N_4903,N_4812);
nand U5083 (N_5083,N_4901,N_4862);
and U5084 (N_5084,N_4859,N_4911);
or U5085 (N_5085,N_4849,N_4989);
nor U5086 (N_5086,N_4856,N_4843);
nand U5087 (N_5087,N_4860,N_4852);
nand U5088 (N_5088,N_4881,N_4825);
or U5089 (N_5089,N_4869,N_4982);
and U5090 (N_5090,N_4957,N_4845);
nand U5091 (N_5091,N_4994,N_4807);
nand U5092 (N_5092,N_4892,N_4876);
nor U5093 (N_5093,N_4873,N_4975);
and U5094 (N_5094,N_4962,N_4979);
or U5095 (N_5095,N_4868,N_4853);
and U5096 (N_5096,N_4995,N_4870);
or U5097 (N_5097,N_4897,N_4803);
xor U5098 (N_5098,N_4977,N_4988);
nor U5099 (N_5099,N_4804,N_4801);
and U5100 (N_5100,N_4950,N_4902);
nand U5101 (N_5101,N_4816,N_4923);
nor U5102 (N_5102,N_4859,N_4880);
nand U5103 (N_5103,N_4987,N_4961);
nand U5104 (N_5104,N_4984,N_4874);
nand U5105 (N_5105,N_4933,N_4991);
nor U5106 (N_5106,N_4841,N_4871);
nand U5107 (N_5107,N_4894,N_4897);
or U5108 (N_5108,N_4867,N_4918);
or U5109 (N_5109,N_4804,N_4870);
and U5110 (N_5110,N_4886,N_4893);
or U5111 (N_5111,N_4887,N_4834);
nor U5112 (N_5112,N_4961,N_4878);
nand U5113 (N_5113,N_4983,N_4947);
and U5114 (N_5114,N_4842,N_4888);
or U5115 (N_5115,N_4989,N_4964);
and U5116 (N_5116,N_4942,N_4918);
nand U5117 (N_5117,N_4834,N_4881);
or U5118 (N_5118,N_4987,N_4813);
and U5119 (N_5119,N_4918,N_4845);
nand U5120 (N_5120,N_4992,N_4840);
or U5121 (N_5121,N_4934,N_4844);
nor U5122 (N_5122,N_4895,N_4916);
nor U5123 (N_5123,N_4881,N_4869);
xor U5124 (N_5124,N_4818,N_4813);
or U5125 (N_5125,N_4826,N_4868);
or U5126 (N_5126,N_4916,N_4835);
nor U5127 (N_5127,N_4958,N_4944);
nor U5128 (N_5128,N_4800,N_4944);
nor U5129 (N_5129,N_4997,N_4965);
or U5130 (N_5130,N_4924,N_4994);
xor U5131 (N_5131,N_4802,N_4990);
and U5132 (N_5132,N_4865,N_4981);
nor U5133 (N_5133,N_4941,N_4841);
or U5134 (N_5134,N_4932,N_4948);
xor U5135 (N_5135,N_4982,N_4810);
or U5136 (N_5136,N_4925,N_4861);
and U5137 (N_5137,N_4850,N_4884);
and U5138 (N_5138,N_4882,N_4893);
or U5139 (N_5139,N_4950,N_4928);
and U5140 (N_5140,N_4801,N_4834);
and U5141 (N_5141,N_4824,N_4964);
xnor U5142 (N_5142,N_4818,N_4904);
nand U5143 (N_5143,N_4829,N_4819);
nand U5144 (N_5144,N_4848,N_4816);
or U5145 (N_5145,N_4817,N_4989);
and U5146 (N_5146,N_4881,N_4909);
nand U5147 (N_5147,N_4855,N_4880);
or U5148 (N_5148,N_4978,N_4948);
or U5149 (N_5149,N_4995,N_4826);
and U5150 (N_5150,N_4992,N_4925);
and U5151 (N_5151,N_4825,N_4912);
and U5152 (N_5152,N_4990,N_4942);
or U5153 (N_5153,N_4946,N_4979);
nand U5154 (N_5154,N_4803,N_4925);
nand U5155 (N_5155,N_4917,N_4807);
nor U5156 (N_5156,N_4968,N_4884);
or U5157 (N_5157,N_4957,N_4865);
and U5158 (N_5158,N_4886,N_4844);
and U5159 (N_5159,N_4972,N_4802);
nor U5160 (N_5160,N_4999,N_4967);
or U5161 (N_5161,N_4888,N_4846);
nor U5162 (N_5162,N_4852,N_4930);
nand U5163 (N_5163,N_4906,N_4813);
or U5164 (N_5164,N_4968,N_4817);
nand U5165 (N_5165,N_4943,N_4824);
nand U5166 (N_5166,N_4858,N_4847);
nor U5167 (N_5167,N_4860,N_4882);
nor U5168 (N_5168,N_4817,N_4990);
or U5169 (N_5169,N_4934,N_4845);
or U5170 (N_5170,N_4962,N_4887);
or U5171 (N_5171,N_4982,N_4941);
and U5172 (N_5172,N_4993,N_4924);
nor U5173 (N_5173,N_4991,N_4964);
and U5174 (N_5174,N_4990,N_4957);
or U5175 (N_5175,N_4938,N_4880);
and U5176 (N_5176,N_4805,N_4977);
or U5177 (N_5177,N_4872,N_4897);
or U5178 (N_5178,N_4994,N_4923);
and U5179 (N_5179,N_4873,N_4805);
or U5180 (N_5180,N_4844,N_4918);
nand U5181 (N_5181,N_4943,N_4932);
and U5182 (N_5182,N_4859,N_4945);
xor U5183 (N_5183,N_4959,N_4906);
or U5184 (N_5184,N_4942,N_4963);
or U5185 (N_5185,N_4819,N_4832);
nand U5186 (N_5186,N_4805,N_4847);
nand U5187 (N_5187,N_4811,N_4844);
nor U5188 (N_5188,N_4892,N_4891);
or U5189 (N_5189,N_4840,N_4920);
nor U5190 (N_5190,N_4904,N_4844);
xnor U5191 (N_5191,N_4922,N_4881);
xor U5192 (N_5192,N_4994,N_4987);
nor U5193 (N_5193,N_4877,N_4995);
nor U5194 (N_5194,N_4958,N_4985);
nand U5195 (N_5195,N_4890,N_4949);
xnor U5196 (N_5196,N_4905,N_4899);
nor U5197 (N_5197,N_4904,N_4857);
nor U5198 (N_5198,N_4838,N_4925);
and U5199 (N_5199,N_4837,N_4939);
or U5200 (N_5200,N_5005,N_5048);
and U5201 (N_5201,N_5180,N_5027);
xnor U5202 (N_5202,N_5078,N_5198);
and U5203 (N_5203,N_5083,N_5117);
and U5204 (N_5204,N_5060,N_5131);
or U5205 (N_5205,N_5140,N_5050);
and U5206 (N_5206,N_5167,N_5188);
or U5207 (N_5207,N_5105,N_5199);
or U5208 (N_5208,N_5042,N_5181);
xor U5209 (N_5209,N_5161,N_5061);
nand U5210 (N_5210,N_5046,N_5107);
and U5211 (N_5211,N_5079,N_5119);
nand U5212 (N_5212,N_5082,N_5157);
and U5213 (N_5213,N_5103,N_5065);
or U5214 (N_5214,N_5186,N_5018);
nand U5215 (N_5215,N_5165,N_5011);
or U5216 (N_5216,N_5139,N_5156);
and U5217 (N_5217,N_5002,N_5182);
nor U5218 (N_5218,N_5033,N_5035);
or U5219 (N_5219,N_5192,N_5125);
xor U5220 (N_5220,N_5054,N_5108);
nor U5221 (N_5221,N_5170,N_5090);
or U5222 (N_5222,N_5190,N_5135);
and U5223 (N_5223,N_5178,N_5123);
nand U5224 (N_5224,N_5066,N_5089);
or U5225 (N_5225,N_5067,N_5038);
and U5226 (N_5226,N_5051,N_5129);
or U5227 (N_5227,N_5019,N_5100);
nand U5228 (N_5228,N_5132,N_5145);
and U5229 (N_5229,N_5091,N_5008);
nand U5230 (N_5230,N_5183,N_5115);
nand U5231 (N_5231,N_5000,N_5168);
or U5232 (N_5232,N_5014,N_5137);
nor U5233 (N_5233,N_5146,N_5080);
and U5234 (N_5234,N_5133,N_5104);
nand U5235 (N_5235,N_5013,N_5193);
and U5236 (N_5236,N_5149,N_5074);
nand U5237 (N_5237,N_5085,N_5023);
xor U5238 (N_5238,N_5053,N_5073);
xnor U5239 (N_5239,N_5185,N_5092);
xnor U5240 (N_5240,N_5062,N_5001);
and U5241 (N_5241,N_5154,N_5166);
nand U5242 (N_5242,N_5072,N_5026);
or U5243 (N_5243,N_5110,N_5003);
or U5244 (N_5244,N_5141,N_5086);
nor U5245 (N_5245,N_5017,N_5142);
nand U5246 (N_5246,N_5195,N_5127);
nor U5247 (N_5247,N_5111,N_5098);
nand U5248 (N_5248,N_5196,N_5102);
xnor U5249 (N_5249,N_5136,N_5016);
and U5250 (N_5250,N_5025,N_5116);
nor U5251 (N_5251,N_5034,N_5112);
nand U5252 (N_5252,N_5101,N_5134);
nor U5253 (N_5253,N_5020,N_5055);
nor U5254 (N_5254,N_5088,N_5172);
nor U5255 (N_5255,N_5138,N_5120);
and U5256 (N_5256,N_5121,N_5064);
and U5257 (N_5257,N_5151,N_5063);
and U5258 (N_5258,N_5099,N_5028);
nor U5259 (N_5259,N_5056,N_5175);
and U5260 (N_5260,N_5007,N_5049);
and U5261 (N_5261,N_5191,N_5009);
nor U5262 (N_5262,N_5094,N_5030);
nor U5263 (N_5263,N_5032,N_5147);
xnor U5264 (N_5264,N_5189,N_5163);
nor U5265 (N_5265,N_5171,N_5126);
nand U5266 (N_5266,N_5118,N_5084);
nand U5267 (N_5267,N_5077,N_5047);
xnor U5268 (N_5268,N_5184,N_5076);
and U5269 (N_5269,N_5070,N_5164);
or U5270 (N_5270,N_5113,N_5057);
xor U5271 (N_5271,N_5155,N_5162);
xnor U5272 (N_5272,N_5031,N_5024);
or U5273 (N_5273,N_5158,N_5177);
nor U5274 (N_5274,N_5152,N_5037);
nand U5275 (N_5275,N_5148,N_5039);
and U5276 (N_5276,N_5052,N_5097);
and U5277 (N_5277,N_5122,N_5095);
nor U5278 (N_5278,N_5015,N_5169);
or U5279 (N_5279,N_5176,N_5160);
or U5280 (N_5280,N_5109,N_5075);
nor U5281 (N_5281,N_5106,N_5006);
nor U5282 (N_5282,N_5114,N_5150);
xor U5283 (N_5283,N_5045,N_5144);
and U5284 (N_5284,N_5174,N_5124);
or U5285 (N_5285,N_5093,N_5004);
nor U5286 (N_5286,N_5040,N_5197);
nor U5287 (N_5287,N_5041,N_5012);
and U5288 (N_5288,N_5153,N_5179);
xnor U5289 (N_5289,N_5081,N_5173);
and U5290 (N_5290,N_5043,N_5029);
nor U5291 (N_5291,N_5096,N_5021);
and U5292 (N_5292,N_5059,N_5143);
xnor U5293 (N_5293,N_5010,N_5187);
nor U5294 (N_5294,N_5194,N_5068);
nor U5295 (N_5295,N_5159,N_5022);
nand U5296 (N_5296,N_5071,N_5058);
nor U5297 (N_5297,N_5044,N_5087);
or U5298 (N_5298,N_5036,N_5130);
and U5299 (N_5299,N_5069,N_5128);
or U5300 (N_5300,N_5059,N_5109);
and U5301 (N_5301,N_5028,N_5044);
nor U5302 (N_5302,N_5006,N_5156);
or U5303 (N_5303,N_5131,N_5005);
xor U5304 (N_5304,N_5065,N_5053);
and U5305 (N_5305,N_5161,N_5159);
or U5306 (N_5306,N_5075,N_5069);
or U5307 (N_5307,N_5169,N_5010);
xnor U5308 (N_5308,N_5122,N_5104);
nand U5309 (N_5309,N_5071,N_5052);
and U5310 (N_5310,N_5058,N_5033);
nand U5311 (N_5311,N_5083,N_5189);
or U5312 (N_5312,N_5097,N_5146);
or U5313 (N_5313,N_5101,N_5008);
nand U5314 (N_5314,N_5188,N_5123);
or U5315 (N_5315,N_5146,N_5085);
or U5316 (N_5316,N_5152,N_5004);
nor U5317 (N_5317,N_5033,N_5193);
nand U5318 (N_5318,N_5057,N_5044);
nand U5319 (N_5319,N_5084,N_5073);
nor U5320 (N_5320,N_5129,N_5034);
nor U5321 (N_5321,N_5132,N_5185);
xor U5322 (N_5322,N_5014,N_5001);
or U5323 (N_5323,N_5109,N_5025);
or U5324 (N_5324,N_5197,N_5185);
and U5325 (N_5325,N_5103,N_5133);
xnor U5326 (N_5326,N_5066,N_5185);
and U5327 (N_5327,N_5097,N_5001);
or U5328 (N_5328,N_5112,N_5080);
nand U5329 (N_5329,N_5082,N_5011);
or U5330 (N_5330,N_5068,N_5162);
or U5331 (N_5331,N_5086,N_5124);
and U5332 (N_5332,N_5045,N_5182);
xor U5333 (N_5333,N_5171,N_5072);
nor U5334 (N_5334,N_5065,N_5059);
and U5335 (N_5335,N_5046,N_5019);
or U5336 (N_5336,N_5036,N_5063);
nor U5337 (N_5337,N_5144,N_5132);
and U5338 (N_5338,N_5042,N_5135);
nor U5339 (N_5339,N_5104,N_5099);
nor U5340 (N_5340,N_5036,N_5067);
or U5341 (N_5341,N_5169,N_5156);
xor U5342 (N_5342,N_5063,N_5130);
and U5343 (N_5343,N_5029,N_5006);
and U5344 (N_5344,N_5018,N_5112);
or U5345 (N_5345,N_5038,N_5035);
nor U5346 (N_5346,N_5059,N_5190);
nor U5347 (N_5347,N_5177,N_5067);
or U5348 (N_5348,N_5077,N_5022);
nand U5349 (N_5349,N_5185,N_5193);
or U5350 (N_5350,N_5143,N_5139);
nor U5351 (N_5351,N_5153,N_5090);
nor U5352 (N_5352,N_5025,N_5087);
or U5353 (N_5353,N_5029,N_5008);
or U5354 (N_5354,N_5036,N_5188);
nand U5355 (N_5355,N_5025,N_5108);
nor U5356 (N_5356,N_5010,N_5180);
and U5357 (N_5357,N_5163,N_5129);
or U5358 (N_5358,N_5190,N_5048);
or U5359 (N_5359,N_5070,N_5069);
and U5360 (N_5360,N_5035,N_5175);
nor U5361 (N_5361,N_5096,N_5005);
or U5362 (N_5362,N_5087,N_5100);
nand U5363 (N_5363,N_5137,N_5093);
nor U5364 (N_5364,N_5141,N_5118);
nor U5365 (N_5365,N_5108,N_5177);
or U5366 (N_5366,N_5079,N_5025);
nand U5367 (N_5367,N_5062,N_5036);
nand U5368 (N_5368,N_5133,N_5187);
nand U5369 (N_5369,N_5132,N_5119);
nor U5370 (N_5370,N_5050,N_5149);
nand U5371 (N_5371,N_5007,N_5186);
and U5372 (N_5372,N_5007,N_5089);
or U5373 (N_5373,N_5070,N_5192);
or U5374 (N_5374,N_5157,N_5150);
or U5375 (N_5375,N_5082,N_5028);
and U5376 (N_5376,N_5198,N_5077);
xnor U5377 (N_5377,N_5190,N_5045);
or U5378 (N_5378,N_5076,N_5117);
nor U5379 (N_5379,N_5115,N_5136);
nor U5380 (N_5380,N_5161,N_5078);
nand U5381 (N_5381,N_5066,N_5178);
nand U5382 (N_5382,N_5191,N_5115);
and U5383 (N_5383,N_5098,N_5123);
and U5384 (N_5384,N_5158,N_5098);
nor U5385 (N_5385,N_5041,N_5037);
or U5386 (N_5386,N_5082,N_5044);
or U5387 (N_5387,N_5142,N_5042);
and U5388 (N_5388,N_5172,N_5049);
nor U5389 (N_5389,N_5175,N_5148);
and U5390 (N_5390,N_5093,N_5044);
xor U5391 (N_5391,N_5124,N_5109);
and U5392 (N_5392,N_5024,N_5160);
nor U5393 (N_5393,N_5085,N_5165);
or U5394 (N_5394,N_5037,N_5142);
or U5395 (N_5395,N_5179,N_5013);
nor U5396 (N_5396,N_5066,N_5014);
or U5397 (N_5397,N_5047,N_5035);
nor U5398 (N_5398,N_5179,N_5023);
xor U5399 (N_5399,N_5117,N_5120);
or U5400 (N_5400,N_5238,N_5294);
nor U5401 (N_5401,N_5299,N_5276);
nor U5402 (N_5402,N_5392,N_5279);
nand U5403 (N_5403,N_5233,N_5267);
and U5404 (N_5404,N_5337,N_5202);
nor U5405 (N_5405,N_5311,N_5380);
nor U5406 (N_5406,N_5338,N_5257);
nand U5407 (N_5407,N_5229,N_5307);
nand U5408 (N_5408,N_5240,N_5212);
or U5409 (N_5409,N_5230,N_5353);
or U5410 (N_5410,N_5272,N_5351);
and U5411 (N_5411,N_5269,N_5378);
nand U5412 (N_5412,N_5358,N_5331);
or U5413 (N_5413,N_5201,N_5357);
xnor U5414 (N_5414,N_5200,N_5205);
xnor U5415 (N_5415,N_5322,N_5333);
or U5416 (N_5416,N_5398,N_5381);
and U5417 (N_5417,N_5298,N_5330);
and U5418 (N_5418,N_5312,N_5232);
nor U5419 (N_5419,N_5255,N_5215);
and U5420 (N_5420,N_5296,N_5341);
nor U5421 (N_5421,N_5317,N_5313);
nor U5422 (N_5422,N_5391,N_5239);
or U5423 (N_5423,N_5211,N_5264);
nand U5424 (N_5424,N_5304,N_5268);
and U5425 (N_5425,N_5302,N_5350);
and U5426 (N_5426,N_5310,N_5334);
xnor U5427 (N_5427,N_5289,N_5342);
and U5428 (N_5428,N_5308,N_5250);
nor U5429 (N_5429,N_5323,N_5325);
nand U5430 (N_5430,N_5343,N_5374);
nand U5431 (N_5431,N_5260,N_5251);
nor U5432 (N_5432,N_5214,N_5383);
and U5433 (N_5433,N_5277,N_5258);
or U5434 (N_5434,N_5319,N_5320);
nor U5435 (N_5435,N_5221,N_5370);
or U5436 (N_5436,N_5244,N_5373);
and U5437 (N_5437,N_5228,N_5284);
and U5438 (N_5438,N_5339,N_5309);
nand U5439 (N_5439,N_5399,N_5223);
nor U5440 (N_5440,N_5281,N_5261);
nor U5441 (N_5441,N_5292,N_5359);
nand U5442 (N_5442,N_5216,N_5278);
nand U5443 (N_5443,N_5242,N_5219);
and U5444 (N_5444,N_5336,N_5354);
or U5445 (N_5445,N_5300,N_5389);
xor U5446 (N_5446,N_5280,N_5248);
nand U5447 (N_5447,N_5328,N_5210);
and U5448 (N_5448,N_5273,N_5345);
nand U5449 (N_5449,N_5327,N_5224);
nand U5450 (N_5450,N_5235,N_5335);
nand U5451 (N_5451,N_5388,N_5288);
or U5452 (N_5452,N_5301,N_5234);
xnor U5453 (N_5453,N_5326,N_5316);
or U5454 (N_5454,N_5290,N_5254);
and U5455 (N_5455,N_5218,N_5225);
or U5456 (N_5456,N_5237,N_5365);
nand U5457 (N_5457,N_5368,N_5249);
xnor U5458 (N_5458,N_5367,N_5241);
and U5459 (N_5459,N_5285,N_5377);
nand U5460 (N_5460,N_5376,N_5375);
nand U5461 (N_5461,N_5259,N_5347);
and U5462 (N_5462,N_5245,N_5386);
or U5463 (N_5463,N_5203,N_5348);
and U5464 (N_5464,N_5329,N_5283);
or U5465 (N_5465,N_5332,N_5209);
or U5466 (N_5466,N_5395,N_5387);
nand U5467 (N_5467,N_5303,N_5396);
nor U5468 (N_5468,N_5355,N_5371);
or U5469 (N_5469,N_5295,N_5393);
nand U5470 (N_5470,N_5364,N_5226);
nand U5471 (N_5471,N_5222,N_5340);
or U5472 (N_5472,N_5220,N_5291);
nand U5473 (N_5473,N_5306,N_5372);
xnor U5474 (N_5474,N_5363,N_5382);
or U5475 (N_5475,N_5270,N_5256);
and U5476 (N_5476,N_5263,N_5394);
nand U5477 (N_5477,N_5390,N_5246);
and U5478 (N_5478,N_5213,N_5344);
nand U5479 (N_5479,N_5282,N_5236);
or U5480 (N_5480,N_5253,N_5362);
or U5481 (N_5481,N_5321,N_5384);
nor U5482 (N_5482,N_5265,N_5231);
nor U5483 (N_5483,N_5208,N_5262);
nor U5484 (N_5484,N_5352,N_5318);
nand U5485 (N_5485,N_5274,N_5346);
nor U5486 (N_5486,N_5266,N_5349);
and U5487 (N_5487,N_5324,N_5252);
and U5488 (N_5488,N_5397,N_5287);
nor U5489 (N_5489,N_5305,N_5297);
nand U5490 (N_5490,N_5369,N_5385);
and U5491 (N_5491,N_5275,N_5207);
and U5492 (N_5492,N_5293,N_5204);
xor U5493 (N_5493,N_5217,N_5227);
nor U5494 (N_5494,N_5314,N_5243);
nand U5495 (N_5495,N_5315,N_5206);
nand U5496 (N_5496,N_5361,N_5271);
and U5497 (N_5497,N_5379,N_5360);
or U5498 (N_5498,N_5247,N_5366);
or U5499 (N_5499,N_5286,N_5356);
or U5500 (N_5500,N_5377,N_5375);
and U5501 (N_5501,N_5256,N_5218);
nand U5502 (N_5502,N_5250,N_5314);
xnor U5503 (N_5503,N_5341,N_5248);
nand U5504 (N_5504,N_5332,N_5294);
nor U5505 (N_5505,N_5326,N_5318);
nand U5506 (N_5506,N_5337,N_5367);
xor U5507 (N_5507,N_5349,N_5376);
xnor U5508 (N_5508,N_5331,N_5396);
or U5509 (N_5509,N_5202,N_5257);
and U5510 (N_5510,N_5268,N_5240);
or U5511 (N_5511,N_5239,N_5367);
or U5512 (N_5512,N_5249,N_5310);
nand U5513 (N_5513,N_5300,N_5231);
and U5514 (N_5514,N_5353,N_5225);
or U5515 (N_5515,N_5391,N_5231);
and U5516 (N_5516,N_5251,N_5344);
nor U5517 (N_5517,N_5239,N_5376);
and U5518 (N_5518,N_5239,N_5295);
and U5519 (N_5519,N_5315,N_5276);
nor U5520 (N_5520,N_5243,N_5364);
nand U5521 (N_5521,N_5361,N_5318);
or U5522 (N_5522,N_5399,N_5389);
nor U5523 (N_5523,N_5236,N_5211);
and U5524 (N_5524,N_5303,N_5234);
nand U5525 (N_5525,N_5313,N_5218);
or U5526 (N_5526,N_5337,N_5289);
xnor U5527 (N_5527,N_5213,N_5386);
and U5528 (N_5528,N_5364,N_5327);
nor U5529 (N_5529,N_5311,N_5350);
nor U5530 (N_5530,N_5277,N_5283);
nor U5531 (N_5531,N_5323,N_5291);
or U5532 (N_5532,N_5385,N_5262);
or U5533 (N_5533,N_5205,N_5247);
nor U5534 (N_5534,N_5212,N_5276);
and U5535 (N_5535,N_5275,N_5242);
or U5536 (N_5536,N_5353,N_5348);
and U5537 (N_5537,N_5272,N_5344);
nor U5538 (N_5538,N_5257,N_5235);
nand U5539 (N_5539,N_5394,N_5350);
or U5540 (N_5540,N_5393,N_5388);
nor U5541 (N_5541,N_5250,N_5249);
or U5542 (N_5542,N_5273,N_5361);
and U5543 (N_5543,N_5302,N_5295);
nor U5544 (N_5544,N_5293,N_5326);
and U5545 (N_5545,N_5226,N_5241);
nor U5546 (N_5546,N_5280,N_5345);
and U5547 (N_5547,N_5382,N_5391);
or U5548 (N_5548,N_5270,N_5207);
nand U5549 (N_5549,N_5361,N_5215);
xnor U5550 (N_5550,N_5394,N_5387);
nor U5551 (N_5551,N_5242,N_5317);
nor U5552 (N_5552,N_5344,N_5273);
and U5553 (N_5553,N_5282,N_5223);
nand U5554 (N_5554,N_5377,N_5242);
or U5555 (N_5555,N_5344,N_5226);
or U5556 (N_5556,N_5286,N_5382);
and U5557 (N_5557,N_5313,N_5338);
nor U5558 (N_5558,N_5391,N_5224);
and U5559 (N_5559,N_5255,N_5323);
nor U5560 (N_5560,N_5347,N_5320);
nand U5561 (N_5561,N_5221,N_5311);
nor U5562 (N_5562,N_5229,N_5315);
nand U5563 (N_5563,N_5311,N_5296);
or U5564 (N_5564,N_5371,N_5234);
and U5565 (N_5565,N_5359,N_5394);
or U5566 (N_5566,N_5356,N_5294);
or U5567 (N_5567,N_5251,N_5218);
and U5568 (N_5568,N_5314,N_5266);
nor U5569 (N_5569,N_5311,N_5391);
and U5570 (N_5570,N_5274,N_5304);
and U5571 (N_5571,N_5364,N_5223);
or U5572 (N_5572,N_5316,N_5211);
and U5573 (N_5573,N_5252,N_5288);
nand U5574 (N_5574,N_5258,N_5240);
nor U5575 (N_5575,N_5226,N_5376);
nor U5576 (N_5576,N_5354,N_5320);
nor U5577 (N_5577,N_5277,N_5361);
nand U5578 (N_5578,N_5221,N_5281);
and U5579 (N_5579,N_5376,N_5275);
xnor U5580 (N_5580,N_5313,N_5211);
nor U5581 (N_5581,N_5246,N_5344);
nand U5582 (N_5582,N_5345,N_5396);
or U5583 (N_5583,N_5240,N_5360);
nor U5584 (N_5584,N_5204,N_5215);
nor U5585 (N_5585,N_5376,N_5296);
nand U5586 (N_5586,N_5365,N_5394);
and U5587 (N_5587,N_5310,N_5343);
and U5588 (N_5588,N_5373,N_5339);
and U5589 (N_5589,N_5236,N_5227);
or U5590 (N_5590,N_5315,N_5288);
nand U5591 (N_5591,N_5225,N_5359);
nand U5592 (N_5592,N_5258,N_5252);
and U5593 (N_5593,N_5235,N_5282);
nor U5594 (N_5594,N_5381,N_5242);
and U5595 (N_5595,N_5325,N_5376);
nor U5596 (N_5596,N_5268,N_5237);
and U5597 (N_5597,N_5242,N_5353);
and U5598 (N_5598,N_5246,N_5209);
and U5599 (N_5599,N_5224,N_5207);
or U5600 (N_5600,N_5429,N_5466);
or U5601 (N_5601,N_5578,N_5444);
nand U5602 (N_5602,N_5596,N_5582);
and U5603 (N_5603,N_5563,N_5531);
or U5604 (N_5604,N_5455,N_5499);
nor U5605 (N_5605,N_5513,N_5526);
or U5606 (N_5606,N_5400,N_5458);
xnor U5607 (N_5607,N_5445,N_5450);
or U5608 (N_5608,N_5503,N_5476);
or U5609 (N_5609,N_5575,N_5443);
or U5610 (N_5610,N_5464,N_5518);
nor U5611 (N_5611,N_5527,N_5406);
and U5612 (N_5612,N_5501,N_5416);
and U5613 (N_5613,N_5423,N_5440);
xnor U5614 (N_5614,N_5534,N_5477);
and U5615 (N_5615,N_5419,N_5481);
nor U5616 (N_5616,N_5583,N_5593);
nand U5617 (N_5617,N_5425,N_5421);
nor U5618 (N_5618,N_5556,N_5576);
or U5619 (N_5619,N_5492,N_5505);
or U5620 (N_5620,N_5407,N_5474);
and U5621 (N_5621,N_5415,N_5432);
and U5622 (N_5622,N_5412,N_5472);
or U5623 (N_5623,N_5469,N_5523);
or U5624 (N_5624,N_5514,N_5540);
and U5625 (N_5625,N_5581,N_5572);
nor U5626 (N_5626,N_5524,N_5473);
or U5627 (N_5627,N_5414,N_5403);
or U5628 (N_5628,N_5555,N_5426);
nand U5629 (N_5629,N_5528,N_5533);
or U5630 (N_5630,N_5559,N_5589);
nor U5631 (N_5631,N_5401,N_5408);
or U5632 (N_5632,N_5545,N_5584);
xor U5633 (N_5633,N_5479,N_5577);
and U5634 (N_5634,N_5436,N_5552);
nand U5635 (N_5635,N_5405,N_5497);
nand U5636 (N_5636,N_5439,N_5550);
nand U5637 (N_5637,N_5538,N_5571);
or U5638 (N_5638,N_5585,N_5428);
and U5639 (N_5639,N_5542,N_5547);
or U5640 (N_5640,N_5516,N_5482);
xor U5641 (N_5641,N_5539,N_5548);
and U5642 (N_5642,N_5586,N_5484);
nor U5643 (N_5643,N_5509,N_5488);
xnor U5644 (N_5644,N_5475,N_5420);
and U5645 (N_5645,N_5459,N_5553);
or U5646 (N_5646,N_5448,N_5591);
or U5647 (N_5647,N_5438,N_5506);
and U5648 (N_5648,N_5561,N_5430);
nand U5649 (N_5649,N_5410,N_5532);
nand U5650 (N_5650,N_5489,N_5504);
nand U5651 (N_5651,N_5595,N_5590);
or U5652 (N_5652,N_5560,N_5562);
nor U5653 (N_5653,N_5465,N_5508);
nand U5654 (N_5654,N_5525,N_5454);
or U5655 (N_5655,N_5433,N_5483);
nand U5656 (N_5656,N_5570,N_5543);
or U5657 (N_5657,N_5512,N_5537);
nand U5658 (N_5658,N_5530,N_5541);
and U5659 (N_5659,N_5404,N_5413);
and U5660 (N_5660,N_5544,N_5486);
and U5661 (N_5661,N_5424,N_5554);
and U5662 (N_5662,N_5587,N_5434);
nor U5663 (N_5663,N_5485,N_5471);
or U5664 (N_5664,N_5568,N_5460);
nor U5665 (N_5665,N_5456,N_5449);
xor U5666 (N_5666,N_5565,N_5487);
or U5667 (N_5667,N_5529,N_5567);
and U5668 (N_5668,N_5470,N_5442);
and U5669 (N_5669,N_5409,N_5549);
nor U5670 (N_5670,N_5510,N_5422);
nand U5671 (N_5671,N_5517,N_5557);
or U5672 (N_5672,N_5495,N_5494);
or U5673 (N_5673,N_5411,N_5515);
nand U5674 (N_5674,N_5579,N_5500);
and U5675 (N_5675,N_5599,N_5463);
xnor U5676 (N_5676,N_5431,N_5519);
or U5677 (N_5677,N_5551,N_5480);
or U5678 (N_5678,N_5592,N_5435);
nor U5679 (N_5679,N_5468,N_5490);
xor U5680 (N_5680,N_5511,N_5597);
nand U5681 (N_5681,N_5453,N_5564);
nor U5682 (N_5682,N_5418,N_5447);
xor U5683 (N_5683,N_5402,N_5521);
nand U5684 (N_5684,N_5457,N_5451);
or U5685 (N_5685,N_5594,N_5441);
nor U5686 (N_5686,N_5574,N_5461);
or U5687 (N_5687,N_5498,N_5536);
and U5688 (N_5688,N_5520,N_5588);
or U5689 (N_5689,N_5546,N_5446);
and U5690 (N_5690,N_5507,N_5462);
xor U5691 (N_5691,N_5493,N_5467);
nand U5692 (N_5692,N_5437,N_5522);
nand U5693 (N_5693,N_5569,N_5566);
nand U5694 (N_5694,N_5478,N_5427);
and U5695 (N_5695,N_5452,N_5580);
nor U5696 (N_5696,N_5417,N_5558);
nand U5697 (N_5697,N_5598,N_5491);
nor U5698 (N_5698,N_5573,N_5535);
or U5699 (N_5699,N_5496,N_5502);
nand U5700 (N_5700,N_5419,N_5590);
nand U5701 (N_5701,N_5476,N_5465);
xor U5702 (N_5702,N_5416,N_5581);
and U5703 (N_5703,N_5441,N_5516);
nand U5704 (N_5704,N_5430,N_5521);
nor U5705 (N_5705,N_5595,N_5571);
or U5706 (N_5706,N_5471,N_5540);
or U5707 (N_5707,N_5401,N_5435);
nor U5708 (N_5708,N_5494,N_5547);
or U5709 (N_5709,N_5498,N_5460);
nand U5710 (N_5710,N_5510,N_5417);
nor U5711 (N_5711,N_5583,N_5532);
xor U5712 (N_5712,N_5571,N_5577);
or U5713 (N_5713,N_5576,N_5432);
and U5714 (N_5714,N_5443,N_5590);
and U5715 (N_5715,N_5530,N_5461);
and U5716 (N_5716,N_5568,N_5567);
and U5717 (N_5717,N_5490,N_5410);
and U5718 (N_5718,N_5579,N_5564);
nor U5719 (N_5719,N_5436,N_5524);
nor U5720 (N_5720,N_5575,N_5474);
and U5721 (N_5721,N_5453,N_5532);
nand U5722 (N_5722,N_5466,N_5587);
and U5723 (N_5723,N_5515,N_5546);
xnor U5724 (N_5724,N_5514,N_5562);
or U5725 (N_5725,N_5507,N_5501);
nor U5726 (N_5726,N_5510,N_5475);
nor U5727 (N_5727,N_5457,N_5481);
and U5728 (N_5728,N_5527,N_5553);
nor U5729 (N_5729,N_5531,N_5495);
xor U5730 (N_5730,N_5444,N_5551);
xnor U5731 (N_5731,N_5471,N_5400);
and U5732 (N_5732,N_5538,N_5553);
and U5733 (N_5733,N_5465,N_5477);
and U5734 (N_5734,N_5550,N_5501);
nand U5735 (N_5735,N_5441,N_5487);
xor U5736 (N_5736,N_5426,N_5445);
and U5737 (N_5737,N_5460,N_5449);
nand U5738 (N_5738,N_5454,N_5410);
nand U5739 (N_5739,N_5521,N_5451);
and U5740 (N_5740,N_5458,N_5515);
or U5741 (N_5741,N_5497,N_5515);
nand U5742 (N_5742,N_5414,N_5562);
nand U5743 (N_5743,N_5488,N_5572);
nand U5744 (N_5744,N_5458,N_5416);
nor U5745 (N_5745,N_5591,N_5524);
nand U5746 (N_5746,N_5595,N_5488);
or U5747 (N_5747,N_5521,N_5514);
nor U5748 (N_5748,N_5515,N_5483);
or U5749 (N_5749,N_5481,N_5586);
nor U5750 (N_5750,N_5572,N_5408);
nor U5751 (N_5751,N_5479,N_5549);
nand U5752 (N_5752,N_5556,N_5599);
xor U5753 (N_5753,N_5528,N_5540);
and U5754 (N_5754,N_5426,N_5525);
and U5755 (N_5755,N_5567,N_5466);
or U5756 (N_5756,N_5546,N_5584);
or U5757 (N_5757,N_5428,N_5409);
and U5758 (N_5758,N_5423,N_5584);
or U5759 (N_5759,N_5457,N_5563);
nand U5760 (N_5760,N_5458,N_5412);
nor U5761 (N_5761,N_5400,N_5499);
and U5762 (N_5762,N_5457,N_5484);
nor U5763 (N_5763,N_5553,N_5586);
or U5764 (N_5764,N_5499,N_5555);
and U5765 (N_5765,N_5531,N_5501);
or U5766 (N_5766,N_5437,N_5545);
and U5767 (N_5767,N_5575,N_5420);
and U5768 (N_5768,N_5445,N_5457);
or U5769 (N_5769,N_5597,N_5501);
nor U5770 (N_5770,N_5438,N_5535);
xnor U5771 (N_5771,N_5588,N_5502);
or U5772 (N_5772,N_5447,N_5429);
nor U5773 (N_5773,N_5534,N_5565);
nor U5774 (N_5774,N_5404,N_5480);
or U5775 (N_5775,N_5546,N_5552);
nor U5776 (N_5776,N_5466,N_5589);
xnor U5777 (N_5777,N_5461,N_5473);
nor U5778 (N_5778,N_5466,N_5556);
nand U5779 (N_5779,N_5524,N_5460);
nor U5780 (N_5780,N_5556,N_5583);
nor U5781 (N_5781,N_5479,N_5556);
nand U5782 (N_5782,N_5444,N_5480);
nor U5783 (N_5783,N_5444,N_5555);
nand U5784 (N_5784,N_5494,N_5477);
nand U5785 (N_5785,N_5464,N_5430);
nand U5786 (N_5786,N_5417,N_5496);
nor U5787 (N_5787,N_5407,N_5522);
nor U5788 (N_5788,N_5450,N_5459);
nor U5789 (N_5789,N_5419,N_5462);
or U5790 (N_5790,N_5423,N_5443);
or U5791 (N_5791,N_5406,N_5525);
nand U5792 (N_5792,N_5496,N_5432);
or U5793 (N_5793,N_5472,N_5582);
nor U5794 (N_5794,N_5509,N_5595);
and U5795 (N_5795,N_5446,N_5592);
xor U5796 (N_5796,N_5428,N_5591);
nor U5797 (N_5797,N_5545,N_5443);
xnor U5798 (N_5798,N_5581,N_5400);
nand U5799 (N_5799,N_5406,N_5407);
nand U5800 (N_5800,N_5775,N_5684);
or U5801 (N_5801,N_5773,N_5638);
and U5802 (N_5802,N_5739,N_5676);
or U5803 (N_5803,N_5659,N_5604);
and U5804 (N_5804,N_5751,N_5704);
nand U5805 (N_5805,N_5727,N_5621);
or U5806 (N_5806,N_5647,N_5677);
or U5807 (N_5807,N_5787,N_5744);
and U5808 (N_5808,N_5678,N_5754);
and U5809 (N_5809,N_5767,N_5792);
nand U5810 (N_5810,N_5639,N_5634);
nand U5811 (N_5811,N_5761,N_5709);
and U5812 (N_5812,N_5642,N_5680);
or U5813 (N_5813,N_5645,N_5672);
or U5814 (N_5814,N_5731,N_5603);
nor U5815 (N_5815,N_5774,N_5636);
xor U5816 (N_5816,N_5786,N_5609);
nor U5817 (N_5817,N_5785,N_5610);
xnor U5818 (N_5818,N_5681,N_5656);
nor U5819 (N_5819,N_5652,N_5762);
and U5820 (N_5820,N_5625,N_5798);
nor U5821 (N_5821,N_5705,N_5673);
nand U5822 (N_5822,N_5766,N_5768);
nor U5823 (N_5823,N_5674,N_5640);
xnor U5824 (N_5824,N_5740,N_5696);
and U5825 (N_5825,N_5752,N_5714);
and U5826 (N_5826,N_5675,N_5772);
nand U5827 (N_5827,N_5613,N_5755);
nand U5828 (N_5828,N_5793,N_5790);
nor U5829 (N_5829,N_5628,N_5671);
and U5830 (N_5830,N_5760,N_5701);
and U5831 (N_5831,N_5765,N_5661);
or U5832 (N_5832,N_5602,N_5637);
nor U5833 (N_5833,N_5641,N_5719);
nor U5834 (N_5834,N_5745,N_5713);
nor U5835 (N_5835,N_5716,N_5718);
or U5836 (N_5836,N_5615,N_5794);
nor U5837 (N_5837,N_5670,N_5758);
nor U5838 (N_5838,N_5729,N_5777);
nor U5839 (N_5839,N_5753,N_5695);
or U5840 (N_5840,N_5683,N_5730);
and U5841 (N_5841,N_5618,N_5622);
and U5842 (N_5842,N_5707,N_5653);
nor U5843 (N_5843,N_5699,N_5749);
or U5844 (N_5844,N_5608,N_5698);
nand U5845 (N_5845,N_5644,N_5779);
xnor U5846 (N_5846,N_5735,N_5624);
nand U5847 (N_5847,N_5650,N_5726);
and U5848 (N_5848,N_5692,N_5697);
nor U5849 (N_5849,N_5776,N_5756);
nand U5850 (N_5850,N_5666,N_5791);
nor U5851 (N_5851,N_5788,N_5799);
and U5852 (N_5852,N_5643,N_5629);
nand U5853 (N_5853,N_5658,N_5736);
or U5854 (N_5854,N_5626,N_5728);
and U5855 (N_5855,N_5606,N_5664);
or U5856 (N_5856,N_5743,N_5738);
or U5857 (N_5857,N_5685,N_5660);
or U5858 (N_5858,N_5654,N_5764);
nor U5859 (N_5859,N_5667,N_5657);
or U5860 (N_5860,N_5627,N_5665);
or U5861 (N_5861,N_5796,N_5620);
nand U5862 (N_5862,N_5607,N_5689);
nand U5863 (N_5863,N_5703,N_5781);
and U5864 (N_5864,N_5797,N_5711);
nand U5865 (N_5865,N_5605,N_5690);
or U5866 (N_5866,N_5601,N_5700);
or U5867 (N_5867,N_5721,N_5795);
nor U5868 (N_5868,N_5693,N_5770);
or U5869 (N_5869,N_5710,N_5668);
nor U5870 (N_5870,N_5663,N_5631);
and U5871 (N_5871,N_5746,N_5734);
and U5872 (N_5872,N_5778,N_5783);
and U5873 (N_5873,N_5702,N_5635);
or U5874 (N_5874,N_5619,N_5682);
or U5875 (N_5875,N_5763,N_5662);
and U5876 (N_5876,N_5687,N_5617);
nand U5877 (N_5877,N_5612,N_5722);
or U5878 (N_5878,N_5679,N_5616);
and U5879 (N_5879,N_5623,N_5769);
and U5880 (N_5880,N_5780,N_5720);
and U5881 (N_5881,N_5748,N_5789);
and U5882 (N_5882,N_5630,N_5648);
or U5883 (N_5883,N_5611,N_5750);
and U5884 (N_5884,N_5691,N_5632);
nor U5885 (N_5885,N_5694,N_5715);
and U5886 (N_5886,N_5724,N_5686);
and U5887 (N_5887,N_5651,N_5614);
nor U5888 (N_5888,N_5723,N_5633);
nand U5889 (N_5889,N_5712,N_5737);
nor U5890 (N_5890,N_5669,N_5771);
and U5891 (N_5891,N_5733,N_5706);
nand U5892 (N_5892,N_5725,N_5784);
nor U5893 (N_5893,N_5688,N_5757);
or U5894 (N_5894,N_5742,N_5741);
nor U5895 (N_5895,N_5782,N_5732);
or U5896 (N_5896,N_5759,N_5708);
and U5897 (N_5897,N_5649,N_5646);
nor U5898 (N_5898,N_5717,N_5655);
nand U5899 (N_5899,N_5600,N_5747);
and U5900 (N_5900,N_5603,N_5795);
nand U5901 (N_5901,N_5699,N_5732);
or U5902 (N_5902,N_5711,N_5751);
and U5903 (N_5903,N_5679,N_5615);
nand U5904 (N_5904,N_5611,N_5721);
nand U5905 (N_5905,N_5792,N_5690);
or U5906 (N_5906,N_5687,N_5762);
xor U5907 (N_5907,N_5612,N_5762);
nor U5908 (N_5908,N_5632,N_5612);
or U5909 (N_5909,N_5737,N_5652);
and U5910 (N_5910,N_5785,N_5728);
nor U5911 (N_5911,N_5654,N_5631);
nand U5912 (N_5912,N_5683,N_5687);
and U5913 (N_5913,N_5715,N_5636);
nor U5914 (N_5914,N_5750,N_5757);
nor U5915 (N_5915,N_5712,N_5618);
nor U5916 (N_5916,N_5716,N_5793);
nor U5917 (N_5917,N_5774,N_5627);
or U5918 (N_5918,N_5701,N_5631);
xnor U5919 (N_5919,N_5697,N_5631);
or U5920 (N_5920,N_5603,N_5677);
xnor U5921 (N_5921,N_5749,N_5785);
nor U5922 (N_5922,N_5787,N_5713);
nor U5923 (N_5923,N_5601,N_5687);
nor U5924 (N_5924,N_5604,N_5601);
and U5925 (N_5925,N_5696,N_5616);
and U5926 (N_5926,N_5663,N_5636);
or U5927 (N_5927,N_5793,N_5795);
nand U5928 (N_5928,N_5695,N_5787);
and U5929 (N_5929,N_5664,N_5789);
and U5930 (N_5930,N_5633,N_5769);
or U5931 (N_5931,N_5607,N_5732);
and U5932 (N_5932,N_5668,N_5643);
and U5933 (N_5933,N_5721,N_5620);
xnor U5934 (N_5934,N_5678,N_5600);
xor U5935 (N_5935,N_5638,N_5771);
and U5936 (N_5936,N_5660,N_5692);
or U5937 (N_5937,N_5695,N_5703);
and U5938 (N_5938,N_5644,N_5708);
nand U5939 (N_5939,N_5716,N_5614);
and U5940 (N_5940,N_5628,N_5617);
and U5941 (N_5941,N_5735,N_5609);
nand U5942 (N_5942,N_5606,N_5635);
nor U5943 (N_5943,N_5628,N_5607);
or U5944 (N_5944,N_5612,N_5754);
or U5945 (N_5945,N_5751,N_5703);
and U5946 (N_5946,N_5683,N_5640);
and U5947 (N_5947,N_5627,N_5682);
and U5948 (N_5948,N_5695,N_5772);
or U5949 (N_5949,N_5716,N_5708);
nand U5950 (N_5950,N_5752,N_5763);
xor U5951 (N_5951,N_5653,N_5686);
and U5952 (N_5952,N_5690,N_5664);
and U5953 (N_5953,N_5604,N_5768);
nor U5954 (N_5954,N_5772,N_5605);
and U5955 (N_5955,N_5629,N_5695);
or U5956 (N_5956,N_5730,N_5689);
nand U5957 (N_5957,N_5633,N_5713);
or U5958 (N_5958,N_5620,N_5605);
and U5959 (N_5959,N_5742,N_5714);
or U5960 (N_5960,N_5705,N_5609);
nand U5961 (N_5961,N_5734,N_5660);
or U5962 (N_5962,N_5778,N_5761);
or U5963 (N_5963,N_5693,N_5664);
or U5964 (N_5964,N_5776,N_5602);
xor U5965 (N_5965,N_5649,N_5765);
and U5966 (N_5966,N_5699,N_5642);
and U5967 (N_5967,N_5766,N_5718);
nand U5968 (N_5968,N_5751,N_5629);
nand U5969 (N_5969,N_5662,N_5720);
and U5970 (N_5970,N_5637,N_5723);
and U5971 (N_5971,N_5662,N_5653);
and U5972 (N_5972,N_5719,N_5709);
and U5973 (N_5973,N_5714,N_5710);
nand U5974 (N_5974,N_5692,N_5713);
nand U5975 (N_5975,N_5691,N_5715);
and U5976 (N_5976,N_5750,N_5607);
and U5977 (N_5977,N_5717,N_5662);
and U5978 (N_5978,N_5742,N_5683);
and U5979 (N_5979,N_5683,N_5724);
or U5980 (N_5980,N_5744,N_5749);
or U5981 (N_5981,N_5771,N_5657);
nor U5982 (N_5982,N_5764,N_5687);
xor U5983 (N_5983,N_5749,N_5734);
or U5984 (N_5984,N_5665,N_5656);
xnor U5985 (N_5985,N_5763,N_5780);
nor U5986 (N_5986,N_5713,N_5781);
nor U5987 (N_5987,N_5615,N_5759);
nand U5988 (N_5988,N_5644,N_5667);
or U5989 (N_5989,N_5610,N_5708);
nor U5990 (N_5990,N_5665,N_5631);
nand U5991 (N_5991,N_5635,N_5685);
or U5992 (N_5992,N_5686,N_5773);
nor U5993 (N_5993,N_5663,N_5722);
nor U5994 (N_5994,N_5631,N_5651);
nand U5995 (N_5995,N_5644,N_5714);
or U5996 (N_5996,N_5691,N_5654);
nand U5997 (N_5997,N_5658,N_5672);
nor U5998 (N_5998,N_5683,N_5738);
and U5999 (N_5999,N_5725,N_5792);
nor U6000 (N_6000,N_5964,N_5850);
nor U6001 (N_6001,N_5913,N_5827);
and U6002 (N_6002,N_5917,N_5871);
and U6003 (N_6003,N_5943,N_5938);
nor U6004 (N_6004,N_5960,N_5941);
or U6005 (N_6005,N_5956,N_5816);
and U6006 (N_6006,N_5823,N_5987);
nor U6007 (N_6007,N_5815,N_5889);
nor U6008 (N_6008,N_5966,N_5974);
and U6009 (N_6009,N_5990,N_5958);
xor U6010 (N_6010,N_5820,N_5894);
xor U6011 (N_6011,N_5809,N_5922);
nand U6012 (N_6012,N_5931,N_5852);
or U6013 (N_6013,N_5854,N_5918);
and U6014 (N_6014,N_5861,N_5910);
or U6015 (N_6015,N_5800,N_5982);
or U6016 (N_6016,N_5991,N_5915);
and U6017 (N_6017,N_5996,N_5880);
and U6018 (N_6018,N_5881,N_5836);
xor U6019 (N_6019,N_5873,N_5972);
nand U6020 (N_6020,N_5868,N_5806);
nand U6021 (N_6021,N_5872,N_5851);
xnor U6022 (N_6022,N_5975,N_5909);
and U6023 (N_6023,N_5927,N_5884);
or U6024 (N_6024,N_5945,N_5825);
nor U6025 (N_6025,N_5988,N_5932);
nor U6026 (N_6026,N_5875,N_5858);
nand U6027 (N_6027,N_5992,N_5979);
and U6028 (N_6028,N_5807,N_5955);
nor U6029 (N_6029,N_5940,N_5834);
xnor U6030 (N_6030,N_5912,N_5828);
and U6031 (N_6031,N_5859,N_5952);
nand U6032 (N_6032,N_5993,N_5887);
nor U6033 (N_6033,N_5950,N_5926);
or U6034 (N_6034,N_5997,N_5830);
nand U6035 (N_6035,N_5892,N_5846);
and U6036 (N_6036,N_5978,N_5929);
nand U6037 (N_6037,N_5923,N_5896);
or U6038 (N_6038,N_5965,N_5935);
nor U6039 (N_6039,N_5981,N_5848);
or U6040 (N_6040,N_5911,N_5954);
or U6041 (N_6041,N_5843,N_5891);
or U6042 (N_6042,N_5925,N_5879);
nand U6043 (N_6043,N_5937,N_5906);
nand U6044 (N_6044,N_5811,N_5842);
and U6045 (N_6045,N_5817,N_5973);
nor U6046 (N_6046,N_5999,N_5949);
or U6047 (N_6047,N_5980,N_5998);
or U6048 (N_6048,N_5976,N_5832);
and U6049 (N_6049,N_5885,N_5962);
and U6050 (N_6050,N_5908,N_5849);
or U6051 (N_6051,N_5920,N_5840);
nor U6052 (N_6052,N_5821,N_5801);
nor U6053 (N_6053,N_5869,N_5814);
and U6054 (N_6054,N_5870,N_5812);
and U6055 (N_6055,N_5983,N_5977);
nor U6056 (N_6056,N_5969,N_5877);
and U6057 (N_6057,N_5863,N_5839);
nand U6058 (N_6058,N_5847,N_5867);
xor U6059 (N_6059,N_5942,N_5984);
and U6060 (N_6060,N_5985,N_5893);
nand U6061 (N_6061,N_5963,N_5934);
or U6062 (N_6062,N_5878,N_5947);
nand U6063 (N_6063,N_5813,N_5805);
nor U6064 (N_6064,N_5959,N_5826);
or U6065 (N_6065,N_5948,N_5921);
and U6066 (N_6066,N_5804,N_5995);
or U6067 (N_6067,N_5862,N_5802);
nand U6068 (N_6068,N_5946,N_5907);
nor U6069 (N_6069,N_5874,N_5844);
nand U6070 (N_6070,N_5961,N_5939);
or U6071 (N_6071,N_5970,N_5899);
or U6072 (N_6072,N_5898,N_5957);
and U6073 (N_6073,N_5895,N_5897);
nand U6074 (N_6074,N_5951,N_5838);
and U6075 (N_6075,N_5822,N_5876);
or U6076 (N_6076,N_5890,N_5924);
or U6077 (N_6077,N_5986,N_5902);
nor U6078 (N_6078,N_5883,N_5882);
nor U6079 (N_6079,N_5971,N_5865);
xor U6080 (N_6080,N_5936,N_5853);
or U6081 (N_6081,N_5824,N_5808);
and U6082 (N_6082,N_5829,N_5928);
nor U6083 (N_6083,N_5900,N_5904);
nor U6084 (N_6084,N_5916,N_5856);
and U6085 (N_6085,N_5903,N_5857);
or U6086 (N_6086,N_5905,N_5901);
or U6087 (N_6087,N_5930,N_5866);
and U6088 (N_6088,N_5989,N_5819);
and U6089 (N_6089,N_5835,N_5944);
nor U6090 (N_6090,N_5837,N_5833);
and U6091 (N_6091,N_5818,N_5845);
nand U6092 (N_6092,N_5855,N_5994);
or U6093 (N_6093,N_5953,N_5888);
or U6094 (N_6094,N_5968,N_5933);
and U6095 (N_6095,N_5967,N_5803);
and U6096 (N_6096,N_5886,N_5914);
nor U6097 (N_6097,N_5841,N_5860);
and U6098 (N_6098,N_5919,N_5810);
and U6099 (N_6099,N_5864,N_5831);
nand U6100 (N_6100,N_5826,N_5885);
nand U6101 (N_6101,N_5921,N_5836);
and U6102 (N_6102,N_5980,N_5875);
nor U6103 (N_6103,N_5850,N_5800);
nand U6104 (N_6104,N_5938,N_5990);
or U6105 (N_6105,N_5982,N_5829);
nor U6106 (N_6106,N_5921,N_5995);
and U6107 (N_6107,N_5887,N_5995);
nand U6108 (N_6108,N_5821,N_5891);
nor U6109 (N_6109,N_5982,N_5904);
nor U6110 (N_6110,N_5923,N_5895);
nor U6111 (N_6111,N_5909,N_5904);
nand U6112 (N_6112,N_5840,N_5947);
nor U6113 (N_6113,N_5970,N_5834);
nand U6114 (N_6114,N_5813,N_5999);
xor U6115 (N_6115,N_5865,N_5931);
xor U6116 (N_6116,N_5943,N_5977);
or U6117 (N_6117,N_5860,N_5919);
and U6118 (N_6118,N_5809,N_5812);
nor U6119 (N_6119,N_5879,N_5864);
or U6120 (N_6120,N_5935,N_5838);
or U6121 (N_6121,N_5955,N_5856);
or U6122 (N_6122,N_5898,N_5987);
or U6123 (N_6123,N_5942,N_5925);
nor U6124 (N_6124,N_5867,N_5879);
and U6125 (N_6125,N_5835,N_5811);
and U6126 (N_6126,N_5904,N_5839);
xor U6127 (N_6127,N_5953,N_5832);
and U6128 (N_6128,N_5967,N_5938);
or U6129 (N_6129,N_5810,N_5960);
and U6130 (N_6130,N_5925,N_5921);
or U6131 (N_6131,N_5966,N_5968);
nor U6132 (N_6132,N_5989,N_5867);
or U6133 (N_6133,N_5824,N_5934);
or U6134 (N_6134,N_5883,N_5950);
or U6135 (N_6135,N_5844,N_5936);
nand U6136 (N_6136,N_5951,N_5931);
and U6137 (N_6137,N_5993,N_5977);
and U6138 (N_6138,N_5940,N_5912);
or U6139 (N_6139,N_5936,N_5828);
nand U6140 (N_6140,N_5803,N_5933);
and U6141 (N_6141,N_5812,N_5976);
nor U6142 (N_6142,N_5977,N_5831);
xnor U6143 (N_6143,N_5990,N_5924);
nand U6144 (N_6144,N_5803,N_5890);
xnor U6145 (N_6145,N_5883,N_5832);
xnor U6146 (N_6146,N_5870,N_5917);
nor U6147 (N_6147,N_5966,N_5860);
nand U6148 (N_6148,N_5950,N_5889);
or U6149 (N_6149,N_5965,N_5908);
or U6150 (N_6150,N_5967,N_5821);
and U6151 (N_6151,N_5825,N_5909);
nor U6152 (N_6152,N_5896,N_5989);
nor U6153 (N_6153,N_5898,N_5865);
or U6154 (N_6154,N_5891,N_5920);
and U6155 (N_6155,N_5879,N_5964);
or U6156 (N_6156,N_5883,N_5970);
and U6157 (N_6157,N_5860,N_5906);
nand U6158 (N_6158,N_5831,N_5862);
nor U6159 (N_6159,N_5959,N_5942);
xor U6160 (N_6160,N_5939,N_5886);
or U6161 (N_6161,N_5949,N_5911);
nand U6162 (N_6162,N_5879,N_5842);
nand U6163 (N_6163,N_5995,N_5880);
or U6164 (N_6164,N_5890,N_5918);
or U6165 (N_6165,N_5967,N_5910);
and U6166 (N_6166,N_5835,N_5881);
nand U6167 (N_6167,N_5985,N_5858);
nor U6168 (N_6168,N_5924,N_5979);
nand U6169 (N_6169,N_5857,N_5844);
nor U6170 (N_6170,N_5904,N_5801);
or U6171 (N_6171,N_5959,N_5962);
and U6172 (N_6172,N_5893,N_5881);
nor U6173 (N_6173,N_5924,N_5981);
and U6174 (N_6174,N_5968,N_5804);
nor U6175 (N_6175,N_5822,N_5905);
and U6176 (N_6176,N_5819,N_5914);
or U6177 (N_6177,N_5856,N_5871);
and U6178 (N_6178,N_5966,N_5839);
xor U6179 (N_6179,N_5866,N_5999);
nand U6180 (N_6180,N_5893,N_5999);
nand U6181 (N_6181,N_5973,N_5897);
xor U6182 (N_6182,N_5913,N_5867);
or U6183 (N_6183,N_5900,N_5981);
nor U6184 (N_6184,N_5880,N_5928);
and U6185 (N_6185,N_5990,N_5961);
nor U6186 (N_6186,N_5895,N_5903);
nand U6187 (N_6187,N_5849,N_5873);
or U6188 (N_6188,N_5986,N_5977);
and U6189 (N_6189,N_5904,N_5898);
nor U6190 (N_6190,N_5849,N_5817);
nand U6191 (N_6191,N_5846,N_5842);
and U6192 (N_6192,N_5804,N_5900);
nor U6193 (N_6193,N_5899,N_5885);
or U6194 (N_6194,N_5944,N_5872);
or U6195 (N_6195,N_5904,N_5876);
or U6196 (N_6196,N_5885,N_5868);
or U6197 (N_6197,N_5920,N_5862);
nor U6198 (N_6198,N_5832,N_5868);
nor U6199 (N_6199,N_5936,N_5832);
nand U6200 (N_6200,N_6137,N_6172);
nor U6201 (N_6201,N_6125,N_6184);
nor U6202 (N_6202,N_6199,N_6144);
or U6203 (N_6203,N_6028,N_6074);
or U6204 (N_6204,N_6058,N_6128);
nor U6205 (N_6205,N_6020,N_6011);
nor U6206 (N_6206,N_6046,N_6016);
nor U6207 (N_6207,N_6067,N_6167);
nand U6208 (N_6208,N_6034,N_6130);
nand U6209 (N_6209,N_6084,N_6123);
and U6210 (N_6210,N_6092,N_6036);
xor U6211 (N_6211,N_6080,N_6068);
and U6212 (N_6212,N_6052,N_6169);
and U6213 (N_6213,N_6127,N_6161);
nor U6214 (N_6214,N_6007,N_6004);
nand U6215 (N_6215,N_6042,N_6168);
xor U6216 (N_6216,N_6055,N_6120);
or U6217 (N_6217,N_6145,N_6005);
and U6218 (N_6218,N_6103,N_6090);
xnor U6219 (N_6219,N_6070,N_6158);
or U6220 (N_6220,N_6148,N_6141);
nor U6221 (N_6221,N_6175,N_6176);
or U6222 (N_6222,N_6157,N_6155);
nand U6223 (N_6223,N_6104,N_6050);
nor U6224 (N_6224,N_6194,N_6013);
or U6225 (N_6225,N_6183,N_6159);
nor U6226 (N_6226,N_6027,N_6022);
and U6227 (N_6227,N_6093,N_6160);
nor U6228 (N_6228,N_6069,N_6162);
xor U6229 (N_6229,N_6089,N_6166);
and U6230 (N_6230,N_6056,N_6086);
nand U6231 (N_6231,N_6193,N_6102);
or U6232 (N_6232,N_6047,N_6024);
or U6233 (N_6233,N_6197,N_6195);
xnor U6234 (N_6234,N_6053,N_6048);
or U6235 (N_6235,N_6009,N_6181);
nand U6236 (N_6236,N_6196,N_6015);
nand U6237 (N_6237,N_6190,N_6006);
nor U6238 (N_6238,N_6062,N_6059);
or U6239 (N_6239,N_6087,N_6031);
and U6240 (N_6240,N_6101,N_6091);
and U6241 (N_6241,N_6105,N_6113);
or U6242 (N_6242,N_6170,N_6153);
nor U6243 (N_6243,N_6136,N_6174);
or U6244 (N_6244,N_6094,N_6049);
or U6245 (N_6245,N_6099,N_6187);
or U6246 (N_6246,N_6061,N_6035);
nor U6247 (N_6247,N_6106,N_6021);
or U6248 (N_6248,N_6008,N_6017);
or U6249 (N_6249,N_6147,N_6109);
nand U6250 (N_6250,N_6154,N_6097);
and U6251 (N_6251,N_6057,N_6019);
nor U6252 (N_6252,N_6073,N_6098);
and U6253 (N_6253,N_6060,N_6054);
nand U6254 (N_6254,N_6082,N_6037);
and U6255 (N_6255,N_6085,N_6023);
nor U6256 (N_6256,N_6081,N_6078);
or U6257 (N_6257,N_6156,N_6121);
or U6258 (N_6258,N_6116,N_6143);
nand U6259 (N_6259,N_6150,N_6044);
or U6260 (N_6260,N_6111,N_6151);
nand U6261 (N_6261,N_6002,N_6179);
nor U6262 (N_6262,N_6180,N_6152);
nor U6263 (N_6263,N_6039,N_6177);
nor U6264 (N_6264,N_6076,N_6064);
nor U6265 (N_6265,N_6117,N_6075);
nor U6266 (N_6266,N_6018,N_6112);
and U6267 (N_6267,N_6040,N_6182);
nor U6268 (N_6268,N_6001,N_6186);
and U6269 (N_6269,N_6030,N_6164);
or U6270 (N_6270,N_6140,N_6129);
nor U6271 (N_6271,N_6000,N_6088);
or U6272 (N_6272,N_6051,N_6014);
and U6273 (N_6273,N_6077,N_6146);
nor U6274 (N_6274,N_6110,N_6045);
and U6275 (N_6275,N_6003,N_6100);
nor U6276 (N_6276,N_6188,N_6114);
nand U6277 (N_6277,N_6043,N_6191);
nor U6278 (N_6278,N_6165,N_6010);
or U6279 (N_6279,N_6026,N_6029);
xnor U6280 (N_6280,N_6083,N_6118);
and U6281 (N_6281,N_6072,N_6071);
nor U6282 (N_6282,N_6139,N_6198);
or U6283 (N_6283,N_6107,N_6135);
and U6284 (N_6284,N_6108,N_6132);
nor U6285 (N_6285,N_6096,N_6134);
nor U6286 (N_6286,N_6189,N_6119);
nor U6287 (N_6287,N_6038,N_6173);
or U6288 (N_6288,N_6033,N_6126);
nor U6289 (N_6289,N_6185,N_6178);
and U6290 (N_6290,N_6079,N_6131);
or U6291 (N_6291,N_6065,N_6142);
and U6292 (N_6292,N_6138,N_6122);
nor U6293 (N_6293,N_6041,N_6171);
nor U6294 (N_6294,N_6066,N_6032);
or U6295 (N_6295,N_6115,N_6012);
and U6296 (N_6296,N_6133,N_6124);
and U6297 (N_6297,N_6149,N_6095);
or U6298 (N_6298,N_6025,N_6192);
xnor U6299 (N_6299,N_6163,N_6063);
nand U6300 (N_6300,N_6129,N_6050);
or U6301 (N_6301,N_6129,N_6183);
and U6302 (N_6302,N_6102,N_6099);
nand U6303 (N_6303,N_6168,N_6093);
or U6304 (N_6304,N_6179,N_6036);
and U6305 (N_6305,N_6018,N_6051);
nand U6306 (N_6306,N_6152,N_6010);
nand U6307 (N_6307,N_6114,N_6132);
nand U6308 (N_6308,N_6040,N_6016);
nand U6309 (N_6309,N_6039,N_6066);
or U6310 (N_6310,N_6037,N_6176);
and U6311 (N_6311,N_6057,N_6083);
nand U6312 (N_6312,N_6112,N_6012);
xnor U6313 (N_6313,N_6068,N_6115);
or U6314 (N_6314,N_6185,N_6037);
nor U6315 (N_6315,N_6019,N_6152);
nand U6316 (N_6316,N_6158,N_6115);
xnor U6317 (N_6317,N_6074,N_6182);
nand U6318 (N_6318,N_6179,N_6181);
or U6319 (N_6319,N_6153,N_6086);
nand U6320 (N_6320,N_6141,N_6084);
nand U6321 (N_6321,N_6090,N_6069);
or U6322 (N_6322,N_6118,N_6165);
and U6323 (N_6323,N_6102,N_6170);
or U6324 (N_6324,N_6192,N_6096);
or U6325 (N_6325,N_6110,N_6123);
and U6326 (N_6326,N_6058,N_6112);
nand U6327 (N_6327,N_6085,N_6163);
nand U6328 (N_6328,N_6117,N_6027);
xor U6329 (N_6329,N_6181,N_6051);
xnor U6330 (N_6330,N_6168,N_6151);
and U6331 (N_6331,N_6041,N_6109);
nor U6332 (N_6332,N_6193,N_6107);
and U6333 (N_6333,N_6055,N_6049);
nor U6334 (N_6334,N_6199,N_6083);
nand U6335 (N_6335,N_6115,N_6063);
or U6336 (N_6336,N_6178,N_6055);
or U6337 (N_6337,N_6063,N_6070);
nor U6338 (N_6338,N_6173,N_6014);
nor U6339 (N_6339,N_6082,N_6096);
nor U6340 (N_6340,N_6125,N_6153);
or U6341 (N_6341,N_6081,N_6147);
nor U6342 (N_6342,N_6065,N_6110);
nand U6343 (N_6343,N_6190,N_6099);
nand U6344 (N_6344,N_6001,N_6043);
and U6345 (N_6345,N_6039,N_6166);
and U6346 (N_6346,N_6182,N_6188);
or U6347 (N_6347,N_6042,N_6013);
and U6348 (N_6348,N_6080,N_6002);
nor U6349 (N_6349,N_6043,N_6017);
xnor U6350 (N_6350,N_6199,N_6044);
nand U6351 (N_6351,N_6002,N_6064);
nand U6352 (N_6352,N_6160,N_6054);
or U6353 (N_6353,N_6196,N_6026);
nand U6354 (N_6354,N_6155,N_6096);
and U6355 (N_6355,N_6182,N_6142);
nand U6356 (N_6356,N_6070,N_6039);
nor U6357 (N_6357,N_6074,N_6186);
nor U6358 (N_6358,N_6083,N_6149);
or U6359 (N_6359,N_6023,N_6011);
or U6360 (N_6360,N_6033,N_6160);
nand U6361 (N_6361,N_6023,N_6092);
nor U6362 (N_6362,N_6186,N_6118);
nand U6363 (N_6363,N_6165,N_6099);
or U6364 (N_6364,N_6166,N_6101);
or U6365 (N_6365,N_6010,N_6198);
and U6366 (N_6366,N_6004,N_6079);
nor U6367 (N_6367,N_6134,N_6143);
nor U6368 (N_6368,N_6050,N_6010);
and U6369 (N_6369,N_6059,N_6115);
or U6370 (N_6370,N_6105,N_6083);
nor U6371 (N_6371,N_6190,N_6118);
or U6372 (N_6372,N_6139,N_6167);
and U6373 (N_6373,N_6011,N_6067);
or U6374 (N_6374,N_6000,N_6022);
and U6375 (N_6375,N_6120,N_6167);
and U6376 (N_6376,N_6111,N_6042);
or U6377 (N_6377,N_6104,N_6116);
nand U6378 (N_6378,N_6105,N_6046);
nor U6379 (N_6379,N_6159,N_6031);
nand U6380 (N_6380,N_6180,N_6188);
xnor U6381 (N_6381,N_6130,N_6152);
or U6382 (N_6382,N_6184,N_6157);
xnor U6383 (N_6383,N_6049,N_6043);
or U6384 (N_6384,N_6178,N_6004);
and U6385 (N_6385,N_6148,N_6090);
and U6386 (N_6386,N_6034,N_6062);
nand U6387 (N_6387,N_6035,N_6104);
or U6388 (N_6388,N_6199,N_6061);
and U6389 (N_6389,N_6063,N_6025);
or U6390 (N_6390,N_6034,N_6029);
or U6391 (N_6391,N_6144,N_6093);
nor U6392 (N_6392,N_6087,N_6157);
nand U6393 (N_6393,N_6111,N_6043);
or U6394 (N_6394,N_6024,N_6114);
and U6395 (N_6395,N_6022,N_6019);
and U6396 (N_6396,N_6090,N_6061);
nor U6397 (N_6397,N_6171,N_6025);
or U6398 (N_6398,N_6112,N_6136);
nand U6399 (N_6399,N_6142,N_6080);
nor U6400 (N_6400,N_6362,N_6219);
nor U6401 (N_6401,N_6311,N_6366);
or U6402 (N_6402,N_6201,N_6394);
nor U6403 (N_6403,N_6202,N_6212);
nor U6404 (N_6404,N_6363,N_6251);
nor U6405 (N_6405,N_6364,N_6268);
xnor U6406 (N_6406,N_6389,N_6215);
or U6407 (N_6407,N_6236,N_6309);
and U6408 (N_6408,N_6387,N_6210);
or U6409 (N_6409,N_6242,N_6345);
and U6410 (N_6410,N_6337,N_6207);
or U6411 (N_6411,N_6203,N_6336);
nor U6412 (N_6412,N_6252,N_6205);
xnor U6413 (N_6413,N_6262,N_6237);
xnor U6414 (N_6414,N_6383,N_6399);
and U6415 (N_6415,N_6211,N_6281);
or U6416 (N_6416,N_6370,N_6290);
or U6417 (N_6417,N_6318,N_6302);
nand U6418 (N_6418,N_6379,N_6213);
and U6419 (N_6419,N_6253,N_6323);
nor U6420 (N_6420,N_6289,N_6348);
xnor U6421 (N_6421,N_6308,N_6293);
or U6422 (N_6422,N_6291,N_6288);
xor U6423 (N_6423,N_6378,N_6304);
nor U6424 (N_6424,N_6350,N_6352);
or U6425 (N_6425,N_6238,N_6277);
nor U6426 (N_6426,N_6327,N_6324);
and U6427 (N_6427,N_6388,N_6384);
and U6428 (N_6428,N_6217,N_6260);
or U6429 (N_6429,N_6306,N_6346);
nand U6430 (N_6430,N_6278,N_6249);
nand U6431 (N_6431,N_6221,N_6233);
nand U6432 (N_6432,N_6276,N_6247);
and U6433 (N_6433,N_6232,N_6230);
nor U6434 (N_6434,N_6270,N_6299);
or U6435 (N_6435,N_6358,N_6376);
nor U6436 (N_6436,N_6355,N_6285);
xor U6437 (N_6437,N_6266,N_6282);
or U6438 (N_6438,N_6382,N_6334);
nor U6439 (N_6439,N_6231,N_6244);
nand U6440 (N_6440,N_6367,N_6329);
and U6441 (N_6441,N_6349,N_6279);
and U6442 (N_6442,N_6371,N_6377);
and U6443 (N_6443,N_6374,N_6385);
nor U6444 (N_6444,N_6225,N_6322);
xnor U6445 (N_6445,N_6274,N_6314);
nand U6446 (N_6446,N_6261,N_6258);
and U6447 (N_6447,N_6300,N_6234);
or U6448 (N_6448,N_6326,N_6246);
or U6449 (N_6449,N_6305,N_6287);
xor U6450 (N_6450,N_6360,N_6259);
nor U6451 (N_6451,N_6295,N_6343);
or U6452 (N_6452,N_6235,N_6257);
and U6453 (N_6453,N_6297,N_6245);
and U6454 (N_6454,N_6284,N_6395);
nor U6455 (N_6455,N_6375,N_6208);
nand U6456 (N_6456,N_6333,N_6338);
nor U6457 (N_6457,N_6292,N_6353);
or U6458 (N_6458,N_6316,N_6373);
or U6459 (N_6459,N_6386,N_6397);
nand U6460 (N_6460,N_6301,N_6303);
nor U6461 (N_6461,N_6347,N_6254);
xor U6462 (N_6462,N_6313,N_6393);
and U6463 (N_6463,N_6264,N_6365);
nand U6464 (N_6464,N_6357,N_6200);
or U6465 (N_6465,N_6354,N_6272);
or U6466 (N_6466,N_6241,N_6380);
and U6467 (N_6467,N_6339,N_6325);
nor U6468 (N_6468,N_6312,N_6228);
and U6469 (N_6469,N_6269,N_6271);
or U6470 (N_6470,N_6321,N_6398);
and U6471 (N_6471,N_6229,N_6224);
nand U6472 (N_6472,N_6239,N_6310);
nand U6473 (N_6473,N_6359,N_6361);
nand U6474 (N_6474,N_6250,N_6392);
and U6475 (N_6475,N_6331,N_6280);
nand U6476 (N_6476,N_6390,N_6317);
or U6477 (N_6477,N_6220,N_6256);
or U6478 (N_6478,N_6243,N_6320);
xor U6479 (N_6479,N_6391,N_6344);
nor U6480 (N_6480,N_6283,N_6307);
nor U6481 (N_6481,N_6332,N_6340);
nor U6482 (N_6482,N_6328,N_6204);
xor U6483 (N_6483,N_6319,N_6294);
xnor U6484 (N_6484,N_6222,N_6248);
or U6485 (N_6485,N_6265,N_6315);
nand U6486 (N_6486,N_6296,N_6240);
and U6487 (N_6487,N_6255,N_6351);
nand U6488 (N_6488,N_6335,N_6206);
or U6489 (N_6489,N_6263,N_6227);
nand U6490 (N_6490,N_6286,N_6226);
and U6491 (N_6491,N_6330,N_6369);
and U6492 (N_6492,N_6216,N_6368);
nand U6493 (N_6493,N_6209,N_6298);
nand U6494 (N_6494,N_6342,N_6223);
or U6495 (N_6495,N_6214,N_6218);
xnor U6496 (N_6496,N_6267,N_6341);
or U6497 (N_6497,N_6273,N_6356);
nor U6498 (N_6498,N_6275,N_6381);
nor U6499 (N_6499,N_6372,N_6396);
nor U6500 (N_6500,N_6335,N_6284);
or U6501 (N_6501,N_6234,N_6374);
or U6502 (N_6502,N_6393,N_6219);
or U6503 (N_6503,N_6385,N_6379);
or U6504 (N_6504,N_6312,N_6219);
xor U6505 (N_6505,N_6261,N_6229);
and U6506 (N_6506,N_6338,N_6350);
and U6507 (N_6507,N_6340,N_6344);
or U6508 (N_6508,N_6274,N_6240);
or U6509 (N_6509,N_6279,N_6238);
xnor U6510 (N_6510,N_6392,N_6262);
or U6511 (N_6511,N_6227,N_6391);
or U6512 (N_6512,N_6228,N_6241);
or U6513 (N_6513,N_6271,N_6200);
or U6514 (N_6514,N_6399,N_6342);
nand U6515 (N_6515,N_6215,N_6376);
nor U6516 (N_6516,N_6222,N_6241);
nand U6517 (N_6517,N_6257,N_6299);
nand U6518 (N_6518,N_6218,N_6216);
nor U6519 (N_6519,N_6282,N_6303);
xnor U6520 (N_6520,N_6397,N_6384);
or U6521 (N_6521,N_6380,N_6263);
or U6522 (N_6522,N_6325,N_6396);
or U6523 (N_6523,N_6360,N_6260);
nor U6524 (N_6524,N_6397,N_6311);
nor U6525 (N_6525,N_6287,N_6369);
nand U6526 (N_6526,N_6398,N_6354);
xor U6527 (N_6527,N_6330,N_6270);
nor U6528 (N_6528,N_6356,N_6293);
or U6529 (N_6529,N_6373,N_6246);
and U6530 (N_6530,N_6232,N_6289);
and U6531 (N_6531,N_6342,N_6301);
and U6532 (N_6532,N_6351,N_6201);
nand U6533 (N_6533,N_6329,N_6253);
or U6534 (N_6534,N_6331,N_6307);
or U6535 (N_6535,N_6308,N_6244);
nor U6536 (N_6536,N_6399,N_6279);
nor U6537 (N_6537,N_6355,N_6327);
nand U6538 (N_6538,N_6212,N_6392);
and U6539 (N_6539,N_6237,N_6280);
nor U6540 (N_6540,N_6290,N_6372);
nand U6541 (N_6541,N_6384,N_6240);
and U6542 (N_6542,N_6370,N_6278);
nand U6543 (N_6543,N_6292,N_6332);
or U6544 (N_6544,N_6202,N_6354);
nand U6545 (N_6545,N_6317,N_6289);
nor U6546 (N_6546,N_6248,N_6399);
nand U6547 (N_6547,N_6381,N_6376);
xor U6548 (N_6548,N_6206,N_6352);
xor U6549 (N_6549,N_6270,N_6329);
or U6550 (N_6550,N_6317,N_6250);
nand U6551 (N_6551,N_6266,N_6237);
nand U6552 (N_6552,N_6219,N_6216);
nand U6553 (N_6553,N_6293,N_6315);
and U6554 (N_6554,N_6204,N_6349);
and U6555 (N_6555,N_6225,N_6238);
nor U6556 (N_6556,N_6378,N_6265);
or U6557 (N_6557,N_6307,N_6320);
nand U6558 (N_6558,N_6307,N_6216);
nor U6559 (N_6559,N_6250,N_6225);
or U6560 (N_6560,N_6335,N_6230);
or U6561 (N_6561,N_6313,N_6356);
or U6562 (N_6562,N_6307,N_6254);
xor U6563 (N_6563,N_6294,N_6289);
or U6564 (N_6564,N_6281,N_6319);
nand U6565 (N_6565,N_6318,N_6259);
and U6566 (N_6566,N_6230,N_6256);
or U6567 (N_6567,N_6262,N_6383);
xor U6568 (N_6568,N_6376,N_6303);
and U6569 (N_6569,N_6278,N_6292);
or U6570 (N_6570,N_6210,N_6207);
or U6571 (N_6571,N_6294,N_6215);
and U6572 (N_6572,N_6259,N_6321);
nand U6573 (N_6573,N_6225,N_6340);
nor U6574 (N_6574,N_6257,N_6324);
and U6575 (N_6575,N_6369,N_6280);
or U6576 (N_6576,N_6330,N_6280);
and U6577 (N_6577,N_6255,N_6346);
nor U6578 (N_6578,N_6248,N_6344);
and U6579 (N_6579,N_6378,N_6317);
and U6580 (N_6580,N_6238,N_6325);
nand U6581 (N_6581,N_6381,N_6223);
and U6582 (N_6582,N_6232,N_6282);
or U6583 (N_6583,N_6221,N_6386);
nand U6584 (N_6584,N_6265,N_6322);
or U6585 (N_6585,N_6260,N_6321);
xnor U6586 (N_6586,N_6226,N_6202);
or U6587 (N_6587,N_6245,N_6383);
nor U6588 (N_6588,N_6352,N_6354);
nor U6589 (N_6589,N_6290,N_6269);
nor U6590 (N_6590,N_6218,N_6205);
or U6591 (N_6591,N_6390,N_6302);
and U6592 (N_6592,N_6306,N_6230);
or U6593 (N_6593,N_6272,N_6280);
xor U6594 (N_6594,N_6216,N_6266);
nor U6595 (N_6595,N_6353,N_6241);
or U6596 (N_6596,N_6285,N_6266);
nor U6597 (N_6597,N_6307,N_6341);
nor U6598 (N_6598,N_6275,N_6226);
nor U6599 (N_6599,N_6389,N_6242);
or U6600 (N_6600,N_6556,N_6526);
and U6601 (N_6601,N_6459,N_6546);
nand U6602 (N_6602,N_6478,N_6432);
nand U6603 (N_6603,N_6584,N_6552);
xnor U6604 (N_6604,N_6542,N_6419);
nand U6605 (N_6605,N_6460,N_6588);
xor U6606 (N_6606,N_6498,N_6538);
and U6607 (N_6607,N_6511,N_6487);
or U6608 (N_6608,N_6446,N_6528);
nor U6609 (N_6609,N_6407,N_6456);
and U6610 (N_6610,N_6406,N_6585);
nand U6611 (N_6611,N_6494,N_6566);
and U6612 (N_6612,N_6402,N_6568);
nor U6613 (N_6613,N_6562,N_6499);
and U6614 (N_6614,N_6464,N_6555);
and U6615 (N_6615,N_6586,N_6574);
and U6616 (N_6616,N_6535,N_6417);
nand U6617 (N_6617,N_6537,N_6401);
or U6618 (N_6618,N_6463,N_6548);
nand U6619 (N_6619,N_6523,N_6480);
xor U6620 (N_6620,N_6557,N_6465);
or U6621 (N_6621,N_6529,N_6409);
or U6622 (N_6622,N_6400,N_6495);
nor U6623 (N_6623,N_6579,N_6578);
nand U6624 (N_6624,N_6420,N_6484);
or U6625 (N_6625,N_6413,N_6505);
and U6626 (N_6626,N_6458,N_6519);
nor U6627 (N_6627,N_6411,N_6434);
or U6628 (N_6628,N_6580,N_6508);
nor U6629 (N_6629,N_6506,N_6572);
or U6630 (N_6630,N_6539,N_6437);
and U6631 (N_6631,N_6563,N_6450);
xor U6632 (N_6632,N_6558,N_6534);
or U6633 (N_6633,N_6520,N_6414);
nor U6634 (N_6634,N_6408,N_6521);
or U6635 (N_6635,N_6507,N_6492);
xor U6636 (N_6636,N_6571,N_6531);
or U6637 (N_6637,N_6481,N_6472);
and U6638 (N_6638,N_6451,N_6582);
nand U6639 (N_6639,N_6564,N_6444);
or U6640 (N_6640,N_6559,N_6416);
nand U6641 (N_6641,N_6423,N_6560);
and U6642 (N_6642,N_6470,N_6404);
xnor U6643 (N_6643,N_6425,N_6482);
and U6644 (N_6644,N_6550,N_6599);
or U6645 (N_6645,N_6412,N_6488);
xor U6646 (N_6646,N_6544,N_6501);
nand U6647 (N_6647,N_6491,N_6569);
nor U6648 (N_6648,N_6471,N_6457);
or U6649 (N_6649,N_6510,N_6593);
and U6650 (N_6650,N_6581,N_6403);
and U6651 (N_6651,N_6469,N_6428);
and U6652 (N_6652,N_6441,N_6504);
xnor U6653 (N_6653,N_6527,N_6490);
or U6654 (N_6654,N_6452,N_6536);
and U6655 (N_6655,N_6485,N_6448);
and U6656 (N_6656,N_6594,N_6424);
nand U6657 (N_6657,N_6573,N_6517);
and U6658 (N_6658,N_6554,N_6410);
nand U6659 (N_6659,N_6575,N_6533);
and U6660 (N_6660,N_6476,N_6541);
nand U6661 (N_6661,N_6597,N_6595);
nand U6662 (N_6662,N_6583,N_6454);
nand U6663 (N_6663,N_6496,N_6455);
and U6664 (N_6664,N_6524,N_6418);
nand U6665 (N_6665,N_6462,N_6502);
nor U6666 (N_6666,N_6512,N_6483);
nor U6667 (N_6667,N_6532,N_6525);
or U6668 (N_6668,N_6598,N_6589);
and U6669 (N_6669,N_6430,N_6576);
nand U6670 (N_6670,N_6590,N_6415);
nor U6671 (N_6671,N_6474,N_6587);
and U6672 (N_6672,N_6473,N_6553);
and U6673 (N_6673,N_6468,N_6421);
or U6674 (N_6674,N_6547,N_6503);
and U6675 (N_6675,N_6431,N_6509);
nor U6676 (N_6676,N_6570,N_6477);
or U6677 (N_6677,N_6500,N_6445);
nand U6678 (N_6678,N_6436,N_6543);
nand U6679 (N_6679,N_6493,N_6435);
and U6680 (N_6680,N_6475,N_6479);
nand U6681 (N_6681,N_6518,N_6540);
nand U6682 (N_6682,N_6561,N_6551);
nand U6683 (N_6683,N_6522,N_6447);
or U6684 (N_6684,N_6567,N_6514);
and U6685 (N_6685,N_6405,N_6515);
or U6686 (N_6686,N_6449,N_6549);
and U6687 (N_6687,N_6467,N_6426);
nor U6688 (N_6688,N_6422,N_6530);
nor U6689 (N_6689,N_6433,N_6486);
and U6690 (N_6690,N_6427,N_6443);
nand U6691 (N_6691,N_6461,N_6565);
xor U6692 (N_6692,N_6489,N_6545);
and U6693 (N_6693,N_6438,N_6513);
nor U6694 (N_6694,N_6439,N_6442);
nor U6695 (N_6695,N_6577,N_6596);
nand U6696 (N_6696,N_6592,N_6497);
or U6697 (N_6697,N_6453,N_6466);
and U6698 (N_6698,N_6591,N_6429);
nand U6699 (N_6699,N_6440,N_6516);
nor U6700 (N_6700,N_6592,N_6553);
nor U6701 (N_6701,N_6542,N_6562);
or U6702 (N_6702,N_6458,N_6421);
nor U6703 (N_6703,N_6435,N_6497);
xnor U6704 (N_6704,N_6535,N_6459);
nand U6705 (N_6705,N_6410,N_6548);
nor U6706 (N_6706,N_6551,N_6529);
nor U6707 (N_6707,N_6527,N_6471);
and U6708 (N_6708,N_6524,N_6584);
or U6709 (N_6709,N_6594,N_6531);
xnor U6710 (N_6710,N_6531,N_6458);
nand U6711 (N_6711,N_6401,N_6581);
and U6712 (N_6712,N_6437,N_6453);
or U6713 (N_6713,N_6459,N_6596);
nor U6714 (N_6714,N_6429,N_6489);
or U6715 (N_6715,N_6535,N_6513);
nor U6716 (N_6716,N_6454,N_6419);
nand U6717 (N_6717,N_6515,N_6431);
nand U6718 (N_6718,N_6439,N_6446);
or U6719 (N_6719,N_6420,N_6436);
and U6720 (N_6720,N_6596,N_6401);
or U6721 (N_6721,N_6495,N_6447);
xor U6722 (N_6722,N_6499,N_6502);
or U6723 (N_6723,N_6429,N_6509);
or U6724 (N_6724,N_6418,N_6419);
and U6725 (N_6725,N_6445,N_6511);
and U6726 (N_6726,N_6477,N_6460);
and U6727 (N_6727,N_6427,N_6400);
nor U6728 (N_6728,N_6534,N_6581);
nor U6729 (N_6729,N_6471,N_6445);
xor U6730 (N_6730,N_6506,N_6561);
and U6731 (N_6731,N_6479,N_6497);
nand U6732 (N_6732,N_6599,N_6463);
and U6733 (N_6733,N_6571,N_6540);
and U6734 (N_6734,N_6595,N_6526);
and U6735 (N_6735,N_6459,N_6517);
nand U6736 (N_6736,N_6596,N_6524);
nor U6737 (N_6737,N_6513,N_6516);
or U6738 (N_6738,N_6453,N_6555);
nand U6739 (N_6739,N_6401,N_6554);
or U6740 (N_6740,N_6585,N_6453);
or U6741 (N_6741,N_6498,N_6569);
or U6742 (N_6742,N_6481,N_6467);
xor U6743 (N_6743,N_6466,N_6494);
nor U6744 (N_6744,N_6458,N_6402);
xor U6745 (N_6745,N_6433,N_6412);
or U6746 (N_6746,N_6436,N_6478);
or U6747 (N_6747,N_6516,N_6538);
nand U6748 (N_6748,N_6564,N_6531);
and U6749 (N_6749,N_6405,N_6571);
and U6750 (N_6750,N_6473,N_6432);
nor U6751 (N_6751,N_6585,N_6531);
or U6752 (N_6752,N_6566,N_6480);
and U6753 (N_6753,N_6426,N_6406);
or U6754 (N_6754,N_6454,N_6484);
and U6755 (N_6755,N_6555,N_6419);
nor U6756 (N_6756,N_6506,N_6553);
or U6757 (N_6757,N_6521,N_6543);
or U6758 (N_6758,N_6522,N_6467);
or U6759 (N_6759,N_6410,N_6510);
nand U6760 (N_6760,N_6509,N_6545);
nor U6761 (N_6761,N_6558,N_6574);
nand U6762 (N_6762,N_6520,N_6435);
or U6763 (N_6763,N_6416,N_6500);
and U6764 (N_6764,N_6486,N_6578);
nor U6765 (N_6765,N_6541,N_6552);
nor U6766 (N_6766,N_6441,N_6584);
nor U6767 (N_6767,N_6405,N_6458);
nand U6768 (N_6768,N_6461,N_6546);
nor U6769 (N_6769,N_6402,N_6583);
nor U6770 (N_6770,N_6596,N_6479);
nor U6771 (N_6771,N_6576,N_6591);
nor U6772 (N_6772,N_6588,N_6512);
nor U6773 (N_6773,N_6590,N_6536);
nand U6774 (N_6774,N_6428,N_6522);
nor U6775 (N_6775,N_6514,N_6557);
xnor U6776 (N_6776,N_6557,N_6431);
nand U6777 (N_6777,N_6435,N_6517);
nor U6778 (N_6778,N_6459,N_6522);
nand U6779 (N_6779,N_6426,N_6562);
and U6780 (N_6780,N_6454,N_6462);
or U6781 (N_6781,N_6442,N_6555);
nor U6782 (N_6782,N_6402,N_6575);
and U6783 (N_6783,N_6447,N_6547);
or U6784 (N_6784,N_6451,N_6489);
nand U6785 (N_6785,N_6409,N_6453);
nand U6786 (N_6786,N_6495,N_6432);
or U6787 (N_6787,N_6505,N_6417);
nor U6788 (N_6788,N_6564,N_6591);
or U6789 (N_6789,N_6416,N_6536);
or U6790 (N_6790,N_6476,N_6434);
nor U6791 (N_6791,N_6547,N_6440);
nand U6792 (N_6792,N_6526,N_6590);
nand U6793 (N_6793,N_6580,N_6478);
xnor U6794 (N_6794,N_6568,N_6573);
and U6795 (N_6795,N_6452,N_6472);
nand U6796 (N_6796,N_6467,N_6409);
nand U6797 (N_6797,N_6403,N_6424);
xnor U6798 (N_6798,N_6503,N_6562);
xor U6799 (N_6799,N_6576,N_6529);
xnor U6800 (N_6800,N_6760,N_6735);
or U6801 (N_6801,N_6692,N_6659);
or U6802 (N_6802,N_6645,N_6775);
xnor U6803 (N_6803,N_6747,N_6723);
nand U6804 (N_6804,N_6722,N_6632);
or U6805 (N_6805,N_6633,N_6706);
and U6806 (N_6806,N_6609,N_6619);
and U6807 (N_6807,N_6602,N_6696);
or U6808 (N_6808,N_6674,N_6748);
and U6809 (N_6809,N_6622,N_6648);
or U6810 (N_6810,N_6707,N_6720);
nand U6811 (N_6811,N_6681,N_6612);
nor U6812 (N_6812,N_6667,N_6610);
nor U6813 (N_6813,N_6640,N_6755);
and U6814 (N_6814,N_6733,N_6744);
and U6815 (N_6815,N_6693,N_6763);
and U6816 (N_6816,N_6660,N_6737);
nor U6817 (N_6817,N_6646,N_6690);
nand U6818 (N_6818,N_6757,N_6784);
nor U6819 (N_6819,N_6698,N_6761);
or U6820 (N_6820,N_6656,N_6637);
or U6821 (N_6821,N_6708,N_6756);
or U6822 (N_6822,N_6684,N_6714);
nor U6823 (N_6823,N_6768,N_6686);
nor U6824 (N_6824,N_6751,N_6673);
nor U6825 (N_6825,N_6629,N_6742);
nand U6826 (N_6826,N_6704,N_6616);
or U6827 (N_6827,N_6741,N_6726);
nand U6828 (N_6828,N_6634,N_6750);
nand U6829 (N_6829,N_6730,N_6752);
and U6830 (N_6830,N_6772,N_6653);
or U6831 (N_6831,N_6724,N_6762);
xnor U6832 (N_6832,N_6689,N_6611);
or U6833 (N_6833,N_6666,N_6627);
or U6834 (N_6834,N_6606,N_6786);
nor U6835 (N_6835,N_6700,N_6743);
and U6836 (N_6836,N_6617,N_6652);
or U6837 (N_6837,N_6703,N_6765);
nand U6838 (N_6838,N_6626,N_6663);
nand U6839 (N_6839,N_6635,N_6771);
xnor U6840 (N_6840,N_6620,N_6655);
and U6841 (N_6841,N_6683,N_6740);
nand U6842 (N_6842,N_6644,N_6642);
xor U6843 (N_6843,N_6710,N_6608);
or U6844 (N_6844,N_6783,N_6709);
nand U6845 (N_6845,N_6713,N_6732);
nor U6846 (N_6846,N_6603,N_6764);
and U6847 (N_6847,N_6647,N_6672);
nand U6848 (N_6848,N_6669,N_6725);
nand U6849 (N_6849,N_6787,N_6643);
nand U6850 (N_6850,N_6717,N_6753);
or U6851 (N_6851,N_6651,N_6798);
nand U6852 (N_6852,N_6662,N_6675);
or U6853 (N_6853,N_6604,N_6668);
nor U6854 (N_6854,N_6780,N_6621);
or U6855 (N_6855,N_6715,N_6745);
nor U6856 (N_6856,N_6613,N_6718);
nand U6857 (N_6857,N_6623,N_6661);
and U6858 (N_6858,N_6694,N_6657);
and U6859 (N_6859,N_6770,N_6794);
or U6860 (N_6860,N_6749,N_6776);
nand U6861 (N_6861,N_6679,N_6793);
xnor U6862 (N_6862,N_6614,N_6716);
xor U6863 (N_6863,N_6600,N_6788);
or U6864 (N_6864,N_6671,N_6699);
nand U6865 (N_6865,N_6685,N_6795);
nand U6866 (N_6866,N_6785,N_6624);
or U6867 (N_6867,N_6797,N_6639);
or U6868 (N_6868,N_6781,N_6796);
or U6869 (N_6869,N_6650,N_6658);
nand U6870 (N_6870,N_6777,N_6680);
nand U6871 (N_6871,N_6705,N_6670);
nor U6872 (N_6872,N_6758,N_6782);
or U6873 (N_6873,N_6778,N_6677);
and U6874 (N_6874,N_6701,N_6759);
nand U6875 (N_6875,N_6799,N_6664);
xor U6876 (N_6876,N_6711,N_6607);
nor U6877 (N_6877,N_6736,N_6631);
or U6878 (N_6878,N_6767,N_6638);
xnor U6879 (N_6879,N_6766,N_6636);
xnor U6880 (N_6880,N_6665,N_6721);
and U6881 (N_6881,N_6739,N_6695);
xnor U6882 (N_6882,N_6712,N_6727);
nor U6883 (N_6883,N_6791,N_6702);
xnor U6884 (N_6884,N_6738,N_6734);
nand U6885 (N_6885,N_6687,N_6630);
nor U6886 (N_6886,N_6688,N_6779);
and U6887 (N_6887,N_6789,N_6792);
nor U6888 (N_6888,N_6731,N_6697);
and U6889 (N_6889,N_6601,N_6774);
or U6890 (N_6890,N_6625,N_6605);
or U6891 (N_6891,N_6691,N_6728);
or U6892 (N_6892,N_6676,N_6649);
or U6893 (N_6893,N_6769,N_6746);
xor U6894 (N_6894,N_6682,N_6678);
nor U6895 (N_6895,N_6790,N_6628);
and U6896 (N_6896,N_6719,N_6754);
and U6897 (N_6897,N_6654,N_6641);
and U6898 (N_6898,N_6618,N_6615);
nor U6899 (N_6899,N_6773,N_6729);
nor U6900 (N_6900,N_6613,N_6612);
nand U6901 (N_6901,N_6750,N_6720);
nor U6902 (N_6902,N_6623,N_6626);
and U6903 (N_6903,N_6619,N_6611);
nor U6904 (N_6904,N_6764,N_6656);
xnor U6905 (N_6905,N_6717,N_6689);
nor U6906 (N_6906,N_6699,N_6785);
xor U6907 (N_6907,N_6621,N_6740);
nand U6908 (N_6908,N_6744,N_6750);
or U6909 (N_6909,N_6618,N_6757);
or U6910 (N_6910,N_6635,N_6679);
or U6911 (N_6911,N_6756,N_6753);
or U6912 (N_6912,N_6728,N_6782);
nor U6913 (N_6913,N_6626,N_6624);
and U6914 (N_6914,N_6749,N_6606);
xor U6915 (N_6915,N_6689,N_6696);
xnor U6916 (N_6916,N_6720,N_6785);
nand U6917 (N_6917,N_6651,N_6761);
nand U6918 (N_6918,N_6746,N_6719);
or U6919 (N_6919,N_6635,N_6698);
nand U6920 (N_6920,N_6769,N_6756);
or U6921 (N_6921,N_6647,N_6608);
xor U6922 (N_6922,N_6750,N_6632);
or U6923 (N_6923,N_6620,N_6717);
xor U6924 (N_6924,N_6714,N_6782);
nand U6925 (N_6925,N_6778,N_6758);
nand U6926 (N_6926,N_6681,N_6735);
nor U6927 (N_6927,N_6614,N_6641);
nand U6928 (N_6928,N_6728,N_6648);
nand U6929 (N_6929,N_6795,N_6679);
xnor U6930 (N_6930,N_6727,N_6680);
nand U6931 (N_6931,N_6768,N_6628);
nand U6932 (N_6932,N_6791,N_6721);
nor U6933 (N_6933,N_6688,N_6639);
or U6934 (N_6934,N_6713,N_6602);
nand U6935 (N_6935,N_6642,N_6792);
nor U6936 (N_6936,N_6744,N_6796);
or U6937 (N_6937,N_6613,N_6606);
xor U6938 (N_6938,N_6634,N_6606);
nand U6939 (N_6939,N_6763,N_6676);
nand U6940 (N_6940,N_6710,N_6739);
nand U6941 (N_6941,N_6786,N_6734);
nor U6942 (N_6942,N_6778,N_6746);
xnor U6943 (N_6943,N_6706,N_6767);
nand U6944 (N_6944,N_6751,N_6783);
xnor U6945 (N_6945,N_6643,N_6654);
xnor U6946 (N_6946,N_6655,N_6786);
or U6947 (N_6947,N_6779,N_6628);
and U6948 (N_6948,N_6713,N_6645);
xor U6949 (N_6949,N_6741,N_6607);
xor U6950 (N_6950,N_6745,N_6710);
or U6951 (N_6951,N_6650,N_6735);
nor U6952 (N_6952,N_6601,N_6795);
nor U6953 (N_6953,N_6789,N_6690);
nand U6954 (N_6954,N_6620,N_6647);
and U6955 (N_6955,N_6647,N_6795);
and U6956 (N_6956,N_6641,N_6797);
and U6957 (N_6957,N_6609,N_6709);
nor U6958 (N_6958,N_6641,N_6719);
nor U6959 (N_6959,N_6789,N_6678);
and U6960 (N_6960,N_6663,N_6721);
and U6961 (N_6961,N_6671,N_6675);
or U6962 (N_6962,N_6667,N_6634);
or U6963 (N_6963,N_6724,N_6641);
nor U6964 (N_6964,N_6702,N_6615);
nand U6965 (N_6965,N_6686,N_6775);
and U6966 (N_6966,N_6687,N_6617);
nand U6967 (N_6967,N_6633,N_6728);
nor U6968 (N_6968,N_6741,N_6653);
or U6969 (N_6969,N_6649,N_6764);
or U6970 (N_6970,N_6713,N_6765);
and U6971 (N_6971,N_6797,N_6695);
nand U6972 (N_6972,N_6629,N_6633);
or U6973 (N_6973,N_6660,N_6723);
xor U6974 (N_6974,N_6669,N_6744);
nor U6975 (N_6975,N_6724,N_6775);
xnor U6976 (N_6976,N_6681,N_6668);
or U6977 (N_6977,N_6633,N_6660);
and U6978 (N_6978,N_6709,N_6628);
xnor U6979 (N_6979,N_6739,N_6743);
or U6980 (N_6980,N_6763,N_6718);
nand U6981 (N_6981,N_6717,N_6694);
or U6982 (N_6982,N_6633,N_6744);
or U6983 (N_6983,N_6795,N_6646);
and U6984 (N_6984,N_6660,N_6690);
nor U6985 (N_6985,N_6607,N_6659);
and U6986 (N_6986,N_6755,N_6602);
and U6987 (N_6987,N_6742,N_6779);
and U6988 (N_6988,N_6649,N_6686);
nand U6989 (N_6989,N_6787,N_6616);
nor U6990 (N_6990,N_6673,N_6686);
nand U6991 (N_6991,N_6737,N_6636);
or U6992 (N_6992,N_6773,N_6719);
or U6993 (N_6993,N_6742,N_6715);
or U6994 (N_6994,N_6677,N_6614);
nand U6995 (N_6995,N_6731,N_6627);
nand U6996 (N_6996,N_6686,N_6714);
nor U6997 (N_6997,N_6726,N_6723);
nand U6998 (N_6998,N_6787,N_6686);
nor U6999 (N_6999,N_6724,N_6791);
and U7000 (N_7000,N_6966,N_6842);
nand U7001 (N_7001,N_6886,N_6879);
xnor U7002 (N_7002,N_6999,N_6908);
nand U7003 (N_7003,N_6857,N_6945);
nor U7004 (N_7004,N_6950,N_6812);
or U7005 (N_7005,N_6905,N_6858);
or U7006 (N_7006,N_6820,N_6807);
nand U7007 (N_7007,N_6972,N_6937);
and U7008 (N_7008,N_6801,N_6979);
nor U7009 (N_7009,N_6996,N_6824);
xnor U7010 (N_7010,N_6891,N_6989);
and U7011 (N_7011,N_6822,N_6893);
nand U7012 (N_7012,N_6918,N_6814);
or U7013 (N_7013,N_6867,N_6919);
and U7014 (N_7014,N_6816,N_6895);
and U7015 (N_7015,N_6809,N_6926);
nor U7016 (N_7016,N_6849,N_6994);
nand U7017 (N_7017,N_6903,N_6869);
xnor U7018 (N_7018,N_6952,N_6909);
nand U7019 (N_7019,N_6991,N_6916);
nor U7020 (N_7020,N_6823,N_6990);
xnor U7021 (N_7021,N_6811,N_6936);
or U7022 (N_7022,N_6815,N_6831);
and U7023 (N_7023,N_6957,N_6804);
and U7024 (N_7024,N_6901,N_6912);
nand U7025 (N_7025,N_6803,N_6942);
nand U7026 (N_7026,N_6840,N_6958);
and U7027 (N_7027,N_6921,N_6946);
and U7028 (N_7028,N_6927,N_6922);
and U7029 (N_7029,N_6883,N_6915);
nand U7030 (N_7030,N_6941,N_6907);
or U7031 (N_7031,N_6951,N_6954);
and U7032 (N_7032,N_6988,N_6976);
xor U7033 (N_7033,N_6913,N_6947);
and U7034 (N_7034,N_6889,N_6839);
nand U7035 (N_7035,N_6987,N_6825);
nand U7036 (N_7036,N_6943,N_6948);
and U7037 (N_7037,N_6884,N_6882);
nand U7038 (N_7038,N_6964,N_6828);
or U7039 (N_7039,N_6995,N_6826);
nand U7040 (N_7040,N_6863,N_6920);
nand U7041 (N_7041,N_6961,N_6876);
xor U7042 (N_7042,N_6938,N_6899);
nand U7043 (N_7043,N_6959,N_6844);
or U7044 (N_7044,N_6865,N_6944);
and U7045 (N_7045,N_6859,N_6874);
nand U7046 (N_7046,N_6956,N_6805);
and U7047 (N_7047,N_6911,N_6851);
or U7048 (N_7048,N_6885,N_6892);
xor U7049 (N_7049,N_6845,N_6819);
nor U7050 (N_7050,N_6939,N_6827);
xor U7051 (N_7051,N_6847,N_6977);
nand U7052 (N_7052,N_6971,N_6953);
or U7053 (N_7053,N_6850,N_6860);
or U7054 (N_7054,N_6923,N_6810);
nor U7055 (N_7055,N_6853,N_6968);
nor U7056 (N_7056,N_6978,N_6897);
or U7057 (N_7057,N_6917,N_6981);
and U7058 (N_7058,N_6870,N_6856);
xor U7059 (N_7059,N_6806,N_6838);
nand U7060 (N_7060,N_6837,N_6969);
or U7061 (N_7061,N_6963,N_6962);
nor U7062 (N_7062,N_6877,N_6967);
or U7063 (N_7063,N_6855,N_6925);
nand U7064 (N_7064,N_6843,N_6872);
and U7065 (N_7065,N_6983,N_6894);
or U7066 (N_7066,N_6873,N_6832);
nor U7067 (N_7067,N_6861,N_6984);
or U7068 (N_7068,N_6993,N_6930);
xnor U7069 (N_7069,N_6802,N_6900);
or U7070 (N_7070,N_6833,N_6980);
nor U7071 (N_7071,N_6914,N_6931);
nor U7072 (N_7072,N_6862,N_6848);
or U7073 (N_7073,N_6955,N_6890);
or U7074 (N_7074,N_6854,N_6821);
or U7075 (N_7075,N_6932,N_6906);
or U7076 (N_7076,N_6880,N_6960);
nand U7077 (N_7077,N_6875,N_6949);
xnor U7078 (N_7078,N_6934,N_6997);
or U7079 (N_7079,N_6924,N_6800);
nand U7080 (N_7080,N_6868,N_6986);
and U7081 (N_7081,N_6904,N_6998);
xor U7082 (N_7082,N_6818,N_6898);
or U7083 (N_7083,N_6841,N_6852);
and U7084 (N_7084,N_6813,N_6817);
and U7085 (N_7085,N_6871,N_6965);
and U7086 (N_7086,N_6940,N_6935);
xor U7087 (N_7087,N_6888,N_6910);
or U7088 (N_7088,N_6846,N_6878);
or U7089 (N_7089,N_6836,N_6929);
or U7090 (N_7090,N_6902,N_6970);
or U7091 (N_7091,N_6829,N_6808);
nand U7092 (N_7092,N_6881,N_6834);
nor U7093 (N_7093,N_6928,N_6973);
nor U7094 (N_7094,N_6864,N_6866);
or U7095 (N_7095,N_6992,N_6933);
xnor U7096 (N_7096,N_6830,N_6974);
nand U7097 (N_7097,N_6985,N_6982);
nor U7098 (N_7098,N_6896,N_6887);
and U7099 (N_7099,N_6835,N_6975);
nand U7100 (N_7100,N_6934,N_6814);
nor U7101 (N_7101,N_6815,N_6990);
and U7102 (N_7102,N_6931,N_6854);
nor U7103 (N_7103,N_6869,N_6971);
xor U7104 (N_7104,N_6823,N_6953);
nor U7105 (N_7105,N_6919,N_6925);
and U7106 (N_7106,N_6850,N_6960);
nor U7107 (N_7107,N_6983,N_6913);
xnor U7108 (N_7108,N_6855,N_6952);
nand U7109 (N_7109,N_6810,N_6815);
or U7110 (N_7110,N_6951,N_6925);
or U7111 (N_7111,N_6813,N_6977);
and U7112 (N_7112,N_6994,N_6923);
and U7113 (N_7113,N_6970,N_6921);
nand U7114 (N_7114,N_6923,N_6970);
or U7115 (N_7115,N_6843,N_6973);
xor U7116 (N_7116,N_6936,N_6952);
nand U7117 (N_7117,N_6801,N_6858);
nor U7118 (N_7118,N_6952,N_6803);
xor U7119 (N_7119,N_6906,N_6831);
nor U7120 (N_7120,N_6836,N_6841);
nand U7121 (N_7121,N_6981,N_6873);
nand U7122 (N_7122,N_6865,N_6830);
nor U7123 (N_7123,N_6833,N_6895);
xor U7124 (N_7124,N_6985,N_6934);
nand U7125 (N_7125,N_6809,N_6908);
nand U7126 (N_7126,N_6830,N_6895);
or U7127 (N_7127,N_6831,N_6958);
nor U7128 (N_7128,N_6908,N_6989);
and U7129 (N_7129,N_6830,N_6945);
nand U7130 (N_7130,N_6953,N_6969);
nor U7131 (N_7131,N_6814,N_6890);
xor U7132 (N_7132,N_6877,N_6916);
and U7133 (N_7133,N_6804,N_6817);
xor U7134 (N_7134,N_6913,N_6945);
nand U7135 (N_7135,N_6894,N_6898);
nand U7136 (N_7136,N_6897,N_6844);
or U7137 (N_7137,N_6904,N_6912);
nand U7138 (N_7138,N_6881,N_6963);
and U7139 (N_7139,N_6994,N_6922);
or U7140 (N_7140,N_6994,N_6934);
nor U7141 (N_7141,N_6821,N_6867);
nor U7142 (N_7142,N_6930,N_6861);
nor U7143 (N_7143,N_6867,N_6803);
and U7144 (N_7144,N_6996,N_6977);
nor U7145 (N_7145,N_6887,N_6976);
nand U7146 (N_7146,N_6806,N_6879);
nor U7147 (N_7147,N_6920,N_6873);
and U7148 (N_7148,N_6821,N_6805);
and U7149 (N_7149,N_6993,N_6937);
nand U7150 (N_7150,N_6891,N_6848);
xnor U7151 (N_7151,N_6930,N_6939);
nor U7152 (N_7152,N_6910,N_6832);
nand U7153 (N_7153,N_6942,N_6872);
nand U7154 (N_7154,N_6882,N_6893);
nand U7155 (N_7155,N_6947,N_6956);
nor U7156 (N_7156,N_6890,N_6833);
nand U7157 (N_7157,N_6929,N_6984);
and U7158 (N_7158,N_6820,N_6976);
and U7159 (N_7159,N_6811,N_6801);
nand U7160 (N_7160,N_6908,N_6980);
and U7161 (N_7161,N_6809,N_6840);
or U7162 (N_7162,N_6982,N_6834);
nand U7163 (N_7163,N_6922,N_6962);
nand U7164 (N_7164,N_6945,N_6941);
and U7165 (N_7165,N_6939,N_6870);
nand U7166 (N_7166,N_6898,N_6837);
or U7167 (N_7167,N_6808,N_6992);
nor U7168 (N_7168,N_6982,N_6877);
nand U7169 (N_7169,N_6980,N_6956);
and U7170 (N_7170,N_6809,N_6930);
xor U7171 (N_7171,N_6944,N_6911);
nand U7172 (N_7172,N_6924,N_6865);
nor U7173 (N_7173,N_6847,N_6964);
and U7174 (N_7174,N_6943,N_6855);
nor U7175 (N_7175,N_6898,N_6963);
nor U7176 (N_7176,N_6952,N_6802);
nor U7177 (N_7177,N_6839,N_6863);
nand U7178 (N_7178,N_6912,N_6834);
nand U7179 (N_7179,N_6869,N_6862);
or U7180 (N_7180,N_6994,N_6891);
nand U7181 (N_7181,N_6975,N_6882);
or U7182 (N_7182,N_6965,N_6972);
and U7183 (N_7183,N_6814,N_6935);
xor U7184 (N_7184,N_6939,N_6801);
and U7185 (N_7185,N_6809,N_6914);
nand U7186 (N_7186,N_6891,N_6887);
nor U7187 (N_7187,N_6874,N_6983);
nand U7188 (N_7188,N_6896,N_6988);
nor U7189 (N_7189,N_6837,N_6967);
nor U7190 (N_7190,N_6870,N_6886);
or U7191 (N_7191,N_6850,N_6935);
nand U7192 (N_7192,N_6941,N_6960);
xor U7193 (N_7193,N_6914,N_6991);
nand U7194 (N_7194,N_6964,N_6900);
and U7195 (N_7195,N_6892,N_6883);
nand U7196 (N_7196,N_6841,N_6992);
or U7197 (N_7197,N_6913,N_6842);
nand U7198 (N_7198,N_6944,N_6868);
xnor U7199 (N_7199,N_6960,N_6872);
nor U7200 (N_7200,N_7153,N_7109);
or U7201 (N_7201,N_7150,N_7070);
nand U7202 (N_7202,N_7022,N_7051);
and U7203 (N_7203,N_7014,N_7125);
nand U7204 (N_7204,N_7132,N_7178);
xor U7205 (N_7205,N_7120,N_7044);
or U7206 (N_7206,N_7110,N_7139);
or U7207 (N_7207,N_7112,N_7005);
nand U7208 (N_7208,N_7168,N_7163);
nand U7209 (N_7209,N_7094,N_7177);
and U7210 (N_7210,N_7102,N_7009);
xor U7211 (N_7211,N_7140,N_7117);
nor U7212 (N_7212,N_7195,N_7021);
nand U7213 (N_7213,N_7010,N_7133);
and U7214 (N_7214,N_7188,N_7081);
or U7215 (N_7215,N_7013,N_7037);
or U7216 (N_7216,N_7033,N_7170);
nand U7217 (N_7217,N_7023,N_7045);
nand U7218 (N_7218,N_7025,N_7060);
and U7219 (N_7219,N_7189,N_7054);
or U7220 (N_7220,N_7171,N_7080);
xnor U7221 (N_7221,N_7151,N_7027);
xor U7222 (N_7222,N_7186,N_7018);
or U7223 (N_7223,N_7115,N_7103);
or U7224 (N_7224,N_7059,N_7169);
and U7225 (N_7225,N_7075,N_7032);
nand U7226 (N_7226,N_7087,N_7137);
and U7227 (N_7227,N_7155,N_7058);
or U7228 (N_7228,N_7172,N_7126);
nand U7229 (N_7229,N_7176,N_7089);
or U7230 (N_7230,N_7124,N_7141);
nor U7231 (N_7231,N_7166,N_7064);
and U7232 (N_7232,N_7052,N_7041);
or U7233 (N_7233,N_7198,N_7161);
and U7234 (N_7234,N_7116,N_7156);
nand U7235 (N_7235,N_7020,N_7056);
nand U7236 (N_7236,N_7136,N_7122);
nand U7237 (N_7237,N_7074,N_7144);
xnor U7238 (N_7238,N_7197,N_7131);
nor U7239 (N_7239,N_7187,N_7101);
and U7240 (N_7240,N_7040,N_7024);
or U7241 (N_7241,N_7082,N_7062);
nor U7242 (N_7242,N_7048,N_7008);
nor U7243 (N_7243,N_7049,N_7012);
nand U7244 (N_7244,N_7199,N_7183);
nor U7245 (N_7245,N_7193,N_7002);
and U7246 (N_7246,N_7174,N_7164);
nor U7247 (N_7247,N_7095,N_7162);
or U7248 (N_7248,N_7068,N_7130);
nand U7249 (N_7249,N_7108,N_7028);
or U7250 (N_7250,N_7063,N_7160);
nor U7251 (N_7251,N_7096,N_7107);
nor U7252 (N_7252,N_7053,N_7091);
nand U7253 (N_7253,N_7065,N_7077);
nor U7254 (N_7254,N_7145,N_7083);
or U7255 (N_7255,N_7142,N_7042);
and U7256 (N_7256,N_7090,N_7105);
or U7257 (N_7257,N_7113,N_7179);
and U7258 (N_7258,N_7128,N_7154);
or U7259 (N_7259,N_7026,N_7015);
nor U7260 (N_7260,N_7046,N_7084);
or U7261 (N_7261,N_7067,N_7143);
nand U7262 (N_7262,N_7182,N_7190);
nand U7263 (N_7263,N_7184,N_7165);
nor U7264 (N_7264,N_7098,N_7088);
and U7265 (N_7265,N_7057,N_7055);
nor U7266 (N_7266,N_7001,N_7030);
and U7267 (N_7267,N_7047,N_7016);
and U7268 (N_7268,N_7158,N_7159);
and U7269 (N_7269,N_7181,N_7085);
or U7270 (N_7270,N_7111,N_7138);
nand U7271 (N_7271,N_7034,N_7011);
and U7272 (N_7272,N_7149,N_7071);
nor U7273 (N_7273,N_7104,N_7029);
nor U7274 (N_7274,N_7031,N_7147);
nor U7275 (N_7275,N_7072,N_7114);
or U7276 (N_7276,N_7118,N_7146);
and U7277 (N_7277,N_7019,N_7038);
nand U7278 (N_7278,N_7191,N_7119);
or U7279 (N_7279,N_7017,N_7073);
or U7280 (N_7280,N_7007,N_7097);
nand U7281 (N_7281,N_7036,N_7167);
nor U7282 (N_7282,N_7127,N_7192);
or U7283 (N_7283,N_7129,N_7121);
nand U7284 (N_7284,N_7006,N_7148);
and U7285 (N_7285,N_7099,N_7185);
xor U7286 (N_7286,N_7078,N_7123);
nor U7287 (N_7287,N_7100,N_7093);
nor U7288 (N_7288,N_7152,N_7000);
nand U7289 (N_7289,N_7092,N_7069);
or U7290 (N_7290,N_7076,N_7066);
nor U7291 (N_7291,N_7175,N_7039);
and U7292 (N_7292,N_7043,N_7194);
nand U7293 (N_7293,N_7086,N_7180);
and U7294 (N_7294,N_7035,N_7196);
nor U7295 (N_7295,N_7050,N_7004);
and U7296 (N_7296,N_7173,N_7157);
nor U7297 (N_7297,N_7079,N_7003);
nor U7298 (N_7298,N_7061,N_7106);
and U7299 (N_7299,N_7135,N_7134);
or U7300 (N_7300,N_7039,N_7078);
or U7301 (N_7301,N_7141,N_7153);
nand U7302 (N_7302,N_7083,N_7158);
and U7303 (N_7303,N_7099,N_7035);
xnor U7304 (N_7304,N_7191,N_7126);
nor U7305 (N_7305,N_7048,N_7045);
and U7306 (N_7306,N_7072,N_7021);
nor U7307 (N_7307,N_7015,N_7195);
nand U7308 (N_7308,N_7112,N_7094);
and U7309 (N_7309,N_7053,N_7109);
or U7310 (N_7310,N_7038,N_7002);
nand U7311 (N_7311,N_7045,N_7174);
xnor U7312 (N_7312,N_7023,N_7033);
nand U7313 (N_7313,N_7183,N_7052);
nand U7314 (N_7314,N_7079,N_7024);
nand U7315 (N_7315,N_7187,N_7092);
or U7316 (N_7316,N_7179,N_7064);
and U7317 (N_7317,N_7068,N_7171);
nand U7318 (N_7318,N_7113,N_7015);
nand U7319 (N_7319,N_7129,N_7127);
or U7320 (N_7320,N_7158,N_7145);
and U7321 (N_7321,N_7102,N_7163);
xnor U7322 (N_7322,N_7079,N_7111);
nor U7323 (N_7323,N_7072,N_7006);
or U7324 (N_7324,N_7118,N_7058);
or U7325 (N_7325,N_7052,N_7019);
and U7326 (N_7326,N_7100,N_7054);
and U7327 (N_7327,N_7028,N_7082);
nor U7328 (N_7328,N_7168,N_7068);
and U7329 (N_7329,N_7045,N_7018);
nor U7330 (N_7330,N_7162,N_7025);
nand U7331 (N_7331,N_7098,N_7198);
or U7332 (N_7332,N_7178,N_7014);
and U7333 (N_7333,N_7018,N_7052);
or U7334 (N_7334,N_7147,N_7181);
nor U7335 (N_7335,N_7039,N_7003);
nand U7336 (N_7336,N_7087,N_7093);
nor U7337 (N_7337,N_7103,N_7083);
nand U7338 (N_7338,N_7018,N_7047);
or U7339 (N_7339,N_7035,N_7181);
nand U7340 (N_7340,N_7022,N_7196);
xor U7341 (N_7341,N_7027,N_7101);
nand U7342 (N_7342,N_7120,N_7111);
xor U7343 (N_7343,N_7100,N_7059);
nand U7344 (N_7344,N_7020,N_7053);
and U7345 (N_7345,N_7114,N_7189);
or U7346 (N_7346,N_7174,N_7094);
nor U7347 (N_7347,N_7101,N_7185);
nand U7348 (N_7348,N_7135,N_7013);
nor U7349 (N_7349,N_7079,N_7043);
nand U7350 (N_7350,N_7041,N_7194);
and U7351 (N_7351,N_7094,N_7013);
nand U7352 (N_7352,N_7048,N_7000);
or U7353 (N_7353,N_7062,N_7105);
or U7354 (N_7354,N_7078,N_7011);
or U7355 (N_7355,N_7091,N_7143);
and U7356 (N_7356,N_7131,N_7169);
or U7357 (N_7357,N_7031,N_7108);
nor U7358 (N_7358,N_7157,N_7049);
or U7359 (N_7359,N_7041,N_7071);
nand U7360 (N_7360,N_7178,N_7157);
and U7361 (N_7361,N_7155,N_7198);
nand U7362 (N_7362,N_7017,N_7090);
nor U7363 (N_7363,N_7194,N_7084);
and U7364 (N_7364,N_7038,N_7076);
nor U7365 (N_7365,N_7104,N_7129);
and U7366 (N_7366,N_7122,N_7063);
and U7367 (N_7367,N_7063,N_7018);
xor U7368 (N_7368,N_7002,N_7146);
nand U7369 (N_7369,N_7051,N_7088);
nand U7370 (N_7370,N_7057,N_7026);
or U7371 (N_7371,N_7055,N_7128);
and U7372 (N_7372,N_7167,N_7108);
and U7373 (N_7373,N_7043,N_7112);
and U7374 (N_7374,N_7198,N_7167);
or U7375 (N_7375,N_7124,N_7077);
or U7376 (N_7376,N_7128,N_7063);
nor U7377 (N_7377,N_7053,N_7140);
xnor U7378 (N_7378,N_7194,N_7087);
or U7379 (N_7379,N_7075,N_7122);
nand U7380 (N_7380,N_7101,N_7173);
and U7381 (N_7381,N_7185,N_7039);
nand U7382 (N_7382,N_7067,N_7135);
nand U7383 (N_7383,N_7056,N_7196);
and U7384 (N_7384,N_7140,N_7114);
nand U7385 (N_7385,N_7047,N_7178);
and U7386 (N_7386,N_7198,N_7192);
xor U7387 (N_7387,N_7125,N_7038);
and U7388 (N_7388,N_7038,N_7100);
nor U7389 (N_7389,N_7089,N_7066);
nor U7390 (N_7390,N_7188,N_7198);
nor U7391 (N_7391,N_7071,N_7014);
and U7392 (N_7392,N_7076,N_7053);
nand U7393 (N_7393,N_7158,N_7174);
nor U7394 (N_7394,N_7019,N_7161);
and U7395 (N_7395,N_7159,N_7125);
nand U7396 (N_7396,N_7012,N_7048);
nor U7397 (N_7397,N_7127,N_7146);
nand U7398 (N_7398,N_7149,N_7113);
and U7399 (N_7399,N_7115,N_7072);
and U7400 (N_7400,N_7267,N_7228);
nor U7401 (N_7401,N_7246,N_7234);
nor U7402 (N_7402,N_7237,N_7241);
nand U7403 (N_7403,N_7276,N_7387);
nand U7404 (N_7404,N_7334,N_7347);
nand U7405 (N_7405,N_7208,N_7391);
nor U7406 (N_7406,N_7271,N_7318);
nand U7407 (N_7407,N_7212,N_7346);
nor U7408 (N_7408,N_7225,N_7289);
nand U7409 (N_7409,N_7362,N_7299);
nand U7410 (N_7410,N_7338,N_7217);
nor U7411 (N_7411,N_7221,N_7363);
nor U7412 (N_7412,N_7245,N_7231);
nor U7413 (N_7413,N_7304,N_7303);
nand U7414 (N_7414,N_7287,N_7311);
nand U7415 (N_7415,N_7355,N_7348);
xor U7416 (N_7416,N_7308,N_7224);
xnor U7417 (N_7417,N_7254,N_7295);
or U7418 (N_7418,N_7356,N_7297);
nor U7419 (N_7419,N_7339,N_7331);
xnor U7420 (N_7420,N_7281,N_7310);
nand U7421 (N_7421,N_7230,N_7305);
and U7422 (N_7422,N_7285,N_7314);
and U7423 (N_7423,N_7213,N_7364);
nor U7424 (N_7424,N_7280,N_7286);
and U7425 (N_7425,N_7220,N_7274);
nor U7426 (N_7426,N_7240,N_7204);
or U7427 (N_7427,N_7319,N_7290);
nand U7428 (N_7428,N_7370,N_7309);
nor U7429 (N_7429,N_7379,N_7223);
nor U7430 (N_7430,N_7366,N_7203);
nand U7431 (N_7431,N_7359,N_7343);
nor U7432 (N_7432,N_7385,N_7229);
and U7433 (N_7433,N_7263,N_7380);
nand U7434 (N_7434,N_7389,N_7353);
and U7435 (N_7435,N_7372,N_7215);
nor U7436 (N_7436,N_7253,N_7317);
nand U7437 (N_7437,N_7368,N_7256);
nand U7438 (N_7438,N_7349,N_7272);
and U7439 (N_7439,N_7376,N_7367);
xnor U7440 (N_7440,N_7216,N_7238);
and U7441 (N_7441,N_7313,N_7211);
nand U7442 (N_7442,N_7307,N_7291);
nand U7443 (N_7443,N_7296,N_7351);
and U7444 (N_7444,N_7265,N_7249);
xor U7445 (N_7445,N_7273,N_7374);
and U7446 (N_7446,N_7327,N_7312);
and U7447 (N_7447,N_7259,N_7328);
and U7448 (N_7448,N_7342,N_7336);
nor U7449 (N_7449,N_7269,N_7218);
nor U7450 (N_7450,N_7322,N_7397);
and U7451 (N_7451,N_7323,N_7392);
xnor U7452 (N_7452,N_7396,N_7315);
nor U7453 (N_7453,N_7268,N_7284);
nand U7454 (N_7454,N_7278,N_7357);
nor U7455 (N_7455,N_7205,N_7382);
xnor U7456 (N_7456,N_7332,N_7227);
xnor U7457 (N_7457,N_7360,N_7373);
or U7458 (N_7458,N_7214,N_7242);
nand U7459 (N_7459,N_7361,N_7300);
nand U7460 (N_7460,N_7202,N_7298);
and U7461 (N_7461,N_7399,N_7395);
nor U7462 (N_7462,N_7371,N_7337);
or U7463 (N_7463,N_7264,N_7325);
nand U7464 (N_7464,N_7283,N_7306);
and U7465 (N_7465,N_7384,N_7239);
or U7466 (N_7466,N_7206,N_7209);
or U7467 (N_7467,N_7282,N_7200);
and U7468 (N_7468,N_7383,N_7394);
or U7469 (N_7469,N_7255,N_7262);
or U7470 (N_7470,N_7236,N_7233);
nand U7471 (N_7471,N_7316,N_7354);
xor U7472 (N_7472,N_7329,N_7292);
nand U7473 (N_7473,N_7393,N_7288);
or U7474 (N_7474,N_7275,N_7333);
or U7475 (N_7475,N_7344,N_7335);
nand U7476 (N_7476,N_7252,N_7219);
or U7477 (N_7477,N_7207,N_7244);
nor U7478 (N_7478,N_7369,N_7251);
or U7479 (N_7479,N_7277,N_7294);
and U7480 (N_7480,N_7301,N_7226);
or U7481 (N_7481,N_7260,N_7302);
nor U7482 (N_7482,N_7201,N_7222);
or U7483 (N_7483,N_7270,N_7345);
nor U7484 (N_7484,N_7377,N_7250);
nor U7485 (N_7485,N_7340,N_7358);
or U7486 (N_7486,N_7279,N_7341);
nand U7487 (N_7487,N_7378,N_7210);
and U7488 (N_7488,N_7352,N_7261);
nand U7489 (N_7489,N_7235,N_7365);
or U7490 (N_7490,N_7386,N_7243);
nor U7491 (N_7491,N_7375,N_7390);
nand U7492 (N_7492,N_7324,N_7381);
nor U7493 (N_7493,N_7398,N_7388);
nand U7494 (N_7494,N_7326,N_7258);
xnor U7495 (N_7495,N_7321,N_7266);
nor U7496 (N_7496,N_7232,N_7320);
nand U7497 (N_7497,N_7257,N_7293);
xor U7498 (N_7498,N_7248,N_7247);
and U7499 (N_7499,N_7330,N_7350);
or U7500 (N_7500,N_7284,N_7223);
nand U7501 (N_7501,N_7354,N_7346);
nor U7502 (N_7502,N_7265,N_7343);
and U7503 (N_7503,N_7298,N_7280);
nor U7504 (N_7504,N_7257,N_7233);
or U7505 (N_7505,N_7335,N_7305);
or U7506 (N_7506,N_7275,N_7385);
xor U7507 (N_7507,N_7386,N_7396);
and U7508 (N_7508,N_7345,N_7289);
and U7509 (N_7509,N_7318,N_7379);
nand U7510 (N_7510,N_7391,N_7239);
and U7511 (N_7511,N_7361,N_7389);
and U7512 (N_7512,N_7220,N_7330);
and U7513 (N_7513,N_7292,N_7280);
xnor U7514 (N_7514,N_7242,N_7338);
nand U7515 (N_7515,N_7223,N_7299);
or U7516 (N_7516,N_7339,N_7384);
and U7517 (N_7517,N_7349,N_7261);
nor U7518 (N_7518,N_7215,N_7380);
and U7519 (N_7519,N_7236,N_7327);
nor U7520 (N_7520,N_7286,N_7211);
or U7521 (N_7521,N_7211,N_7377);
and U7522 (N_7522,N_7254,N_7270);
and U7523 (N_7523,N_7246,N_7263);
and U7524 (N_7524,N_7215,N_7331);
nor U7525 (N_7525,N_7209,N_7307);
and U7526 (N_7526,N_7331,N_7321);
and U7527 (N_7527,N_7297,N_7269);
nand U7528 (N_7528,N_7257,N_7240);
xnor U7529 (N_7529,N_7274,N_7316);
and U7530 (N_7530,N_7226,N_7229);
nor U7531 (N_7531,N_7345,N_7381);
and U7532 (N_7532,N_7268,N_7311);
xor U7533 (N_7533,N_7359,N_7277);
nand U7534 (N_7534,N_7373,N_7202);
and U7535 (N_7535,N_7330,N_7308);
nor U7536 (N_7536,N_7303,N_7331);
nor U7537 (N_7537,N_7318,N_7305);
and U7538 (N_7538,N_7281,N_7377);
and U7539 (N_7539,N_7306,N_7206);
or U7540 (N_7540,N_7230,N_7395);
or U7541 (N_7541,N_7277,N_7306);
and U7542 (N_7542,N_7371,N_7358);
or U7543 (N_7543,N_7300,N_7221);
and U7544 (N_7544,N_7200,N_7332);
or U7545 (N_7545,N_7308,N_7392);
and U7546 (N_7546,N_7364,N_7269);
nor U7547 (N_7547,N_7290,N_7232);
and U7548 (N_7548,N_7213,N_7336);
xor U7549 (N_7549,N_7218,N_7392);
xnor U7550 (N_7550,N_7286,N_7205);
and U7551 (N_7551,N_7399,N_7202);
nor U7552 (N_7552,N_7226,N_7294);
nand U7553 (N_7553,N_7334,N_7353);
and U7554 (N_7554,N_7302,N_7351);
xor U7555 (N_7555,N_7326,N_7290);
and U7556 (N_7556,N_7237,N_7279);
nand U7557 (N_7557,N_7200,N_7385);
or U7558 (N_7558,N_7378,N_7256);
nand U7559 (N_7559,N_7309,N_7363);
or U7560 (N_7560,N_7283,N_7393);
nand U7561 (N_7561,N_7397,N_7364);
nand U7562 (N_7562,N_7375,N_7302);
nand U7563 (N_7563,N_7288,N_7272);
and U7564 (N_7564,N_7238,N_7344);
nand U7565 (N_7565,N_7217,N_7213);
or U7566 (N_7566,N_7209,N_7317);
or U7567 (N_7567,N_7354,N_7209);
nor U7568 (N_7568,N_7316,N_7340);
or U7569 (N_7569,N_7274,N_7293);
and U7570 (N_7570,N_7202,N_7207);
nand U7571 (N_7571,N_7295,N_7318);
or U7572 (N_7572,N_7204,N_7337);
or U7573 (N_7573,N_7249,N_7323);
nand U7574 (N_7574,N_7201,N_7225);
nand U7575 (N_7575,N_7290,N_7203);
nor U7576 (N_7576,N_7342,N_7224);
nor U7577 (N_7577,N_7353,N_7263);
nor U7578 (N_7578,N_7364,N_7271);
and U7579 (N_7579,N_7292,N_7272);
nor U7580 (N_7580,N_7266,N_7364);
xor U7581 (N_7581,N_7314,N_7219);
nor U7582 (N_7582,N_7332,N_7350);
nor U7583 (N_7583,N_7282,N_7239);
and U7584 (N_7584,N_7214,N_7307);
and U7585 (N_7585,N_7395,N_7209);
and U7586 (N_7586,N_7388,N_7200);
or U7587 (N_7587,N_7326,N_7393);
nor U7588 (N_7588,N_7236,N_7257);
nor U7589 (N_7589,N_7268,N_7254);
nor U7590 (N_7590,N_7327,N_7240);
nand U7591 (N_7591,N_7362,N_7399);
nand U7592 (N_7592,N_7359,N_7325);
and U7593 (N_7593,N_7301,N_7344);
and U7594 (N_7594,N_7280,N_7328);
or U7595 (N_7595,N_7275,N_7203);
and U7596 (N_7596,N_7373,N_7287);
nand U7597 (N_7597,N_7246,N_7321);
nand U7598 (N_7598,N_7232,N_7314);
nor U7599 (N_7599,N_7310,N_7344);
or U7600 (N_7600,N_7562,N_7429);
xnor U7601 (N_7601,N_7408,N_7435);
or U7602 (N_7602,N_7433,N_7472);
and U7603 (N_7603,N_7478,N_7491);
nor U7604 (N_7604,N_7502,N_7579);
or U7605 (N_7605,N_7409,N_7516);
nor U7606 (N_7606,N_7583,N_7552);
nand U7607 (N_7607,N_7553,N_7437);
or U7608 (N_7608,N_7531,N_7426);
and U7609 (N_7609,N_7450,N_7447);
xnor U7610 (N_7610,N_7507,N_7561);
nand U7611 (N_7611,N_7411,N_7536);
and U7612 (N_7612,N_7467,N_7477);
and U7613 (N_7613,N_7566,N_7572);
nor U7614 (N_7614,N_7508,N_7456);
and U7615 (N_7615,N_7521,N_7453);
or U7616 (N_7616,N_7468,N_7532);
or U7617 (N_7617,N_7405,N_7410);
and U7618 (N_7618,N_7551,N_7458);
nor U7619 (N_7619,N_7485,N_7500);
nand U7620 (N_7620,N_7587,N_7495);
or U7621 (N_7621,N_7591,N_7471);
nand U7622 (N_7622,N_7476,N_7549);
nor U7623 (N_7623,N_7509,N_7525);
nand U7624 (N_7624,N_7506,N_7582);
nor U7625 (N_7625,N_7596,N_7480);
or U7626 (N_7626,N_7479,N_7580);
nor U7627 (N_7627,N_7415,N_7510);
or U7628 (N_7628,N_7436,N_7486);
and U7629 (N_7629,N_7440,N_7565);
nor U7630 (N_7630,N_7545,N_7524);
nand U7631 (N_7631,N_7599,N_7513);
or U7632 (N_7632,N_7519,N_7463);
and U7633 (N_7633,N_7412,N_7403);
nand U7634 (N_7634,N_7539,N_7404);
nor U7635 (N_7635,N_7558,N_7464);
nand U7636 (N_7636,N_7465,N_7444);
or U7637 (N_7637,N_7452,N_7592);
xor U7638 (N_7638,N_7449,N_7446);
xor U7639 (N_7639,N_7497,N_7431);
or U7640 (N_7640,N_7407,N_7504);
or U7641 (N_7641,N_7540,N_7460);
and U7642 (N_7642,N_7578,N_7575);
nor U7643 (N_7643,N_7439,N_7597);
and U7644 (N_7644,N_7454,N_7505);
or U7645 (N_7645,N_7402,N_7424);
xor U7646 (N_7646,N_7533,N_7581);
nor U7647 (N_7647,N_7514,N_7593);
and U7648 (N_7648,N_7498,N_7541);
or U7649 (N_7649,N_7530,N_7470);
or U7650 (N_7650,N_7420,N_7573);
nand U7651 (N_7651,N_7534,N_7434);
or U7652 (N_7652,N_7482,N_7401);
xor U7653 (N_7653,N_7584,N_7515);
nor U7654 (N_7654,N_7569,N_7547);
or U7655 (N_7655,N_7481,N_7438);
and U7656 (N_7656,N_7421,N_7490);
nand U7657 (N_7657,N_7537,N_7511);
or U7658 (N_7658,N_7418,N_7590);
nand U7659 (N_7659,N_7432,N_7496);
xnor U7660 (N_7660,N_7448,N_7589);
and U7661 (N_7661,N_7577,N_7417);
and U7662 (N_7662,N_7441,N_7564);
nand U7663 (N_7663,N_7474,N_7503);
xor U7664 (N_7664,N_7517,N_7554);
and U7665 (N_7665,N_7576,N_7492);
or U7666 (N_7666,N_7488,N_7527);
or U7667 (N_7667,N_7568,N_7487);
or U7668 (N_7668,N_7520,N_7571);
nand U7669 (N_7669,N_7574,N_7425);
or U7670 (N_7670,N_7475,N_7588);
nor U7671 (N_7671,N_7542,N_7543);
xor U7672 (N_7672,N_7489,N_7512);
or U7673 (N_7673,N_7422,N_7570);
nor U7674 (N_7674,N_7550,N_7406);
nor U7675 (N_7675,N_7400,N_7494);
nand U7676 (N_7676,N_7598,N_7428);
and U7677 (N_7677,N_7526,N_7457);
nand U7678 (N_7678,N_7535,N_7501);
nand U7679 (N_7679,N_7556,N_7455);
nor U7680 (N_7680,N_7560,N_7522);
xnor U7681 (N_7681,N_7469,N_7466);
or U7682 (N_7682,N_7461,N_7423);
or U7683 (N_7683,N_7538,N_7595);
or U7684 (N_7684,N_7529,N_7459);
or U7685 (N_7685,N_7473,N_7546);
and U7686 (N_7686,N_7427,N_7414);
nand U7687 (N_7687,N_7548,N_7557);
nor U7688 (N_7688,N_7493,N_7563);
xnor U7689 (N_7689,N_7462,N_7416);
nor U7690 (N_7690,N_7518,N_7544);
nor U7691 (N_7691,N_7445,N_7442);
or U7692 (N_7692,N_7413,N_7528);
or U7693 (N_7693,N_7484,N_7559);
nand U7694 (N_7694,N_7586,N_7585);
xnor U7695 (N_7695,N_7451,N_7419);
and U7696 (N_7696,N_7555,N_7430);
nor U7697 (N_7697,N_7567,N_7523);
xnor U7698 (N_7698,N_7483,N_7499);
nor U7699 (N_7699,N_7443,N_7594);
nor U7700 (N_7700,N_7513,N_7529);
or U7701 (N_7701,N_7583,N_7403);
or U7702 (N_7702,N_7404,N_7443);
or U7703 (N_7703,N_7563,N_7468);
or U7704 (N_7704,N_7491,N_7474);
and U7705 (N_7705,N_7446,N_7498);
and U7706 (N_7706,N_7404,N_7513);
and U7707 (N_7707,N_7426,N_7430);
nand U7708 (N_7708,N_7497,N_7494);
or U7709 (N_7709,N_7541,N_7584);
and U7710 (N_7710,N_7458,N_7590);
nor U7711 (N_7711,N_7404,N_7560);
nor U7712 (N_7712,N_7469,N_7473);
nand U7713 (N_7713,N_7440,N_7538);
nand U7714 (N_7714,N_7480,N_7591);
nor U7715 (N_7715,N_7520,N_7500);
nor U7716 (N_7716,N_7440,N_7450);
nor U7717 (N_7717,N_7420,N_7551);
xor U7718 (N_7718,N_7423,N_7472);
nand U7719 (N_7719,N_7484,N_7521);
nand U7720 (N_7720,N_7546,N_7577);
nor U7721 (N_7721,N_7451,N_7460);
xnor U7722 (N_7722,N_7545,N_7446);
nand U7723 (N_7723,N_7553,N_7517);
nor U7724 (N_7724,N_7478,N_7503);
nand U7725 (N_7725,N_7584,N_7432);
and U7726 (N_7726,N_7477,N_7455);
and U7727 (N_7727,N_7517,N_7588);
or U7728 (N_7728,N_7568,N_7572);
and U7729 (N_7729,N_7548,N_7529);
nand U7730 (N_7730,N_7579,N_7423);
xor U7731 (N_7731,N_7457,N_7538);
or U7732 (N_7732,N_7491,N_7413);
nor U7733 (N_7733,N_7524,N_7425);
or U7734 (N_7734,N_7565,N_7588);
nand U7735 (N_7735,N_7498,N_7470);
nand U7736 (N_7736,N_7470,N_7567);
or U7737 (N_7737,N_7402,N_7519);
or U7738 (N_7738,N_7478,N_7539);
and U7739 (N_7739,N_7424,N_7414);
nand U7740 (N_7740,N_7424,N_7488);
or U7741 (N_7741,N_7457,N_7463);
xnor U7742 (N_7742,N_7578,N_7471);
or U7743 (N_7743,N_7438,N_7598);
nor U7744 (N_7744,N_7480,N_7456);
nor U7745 (N_7745,N_7564,N_7517);
nand U7746 (N_7746,N_7565,N_7577);
or U7747 (N_7747,N_7582,N_7435);
or U7748 (N_7748,N_7535,N_7497);
nand U7749 (N_7749,N_7536,N_7477);
or U7750 (N_7750,N_7563,N_7519);
or U7751 (N_7751,N_7418,N_7413);
or U7752 (N_7752,N_7513,N_7542);
or U7753 (N_7753,N_7526,N_7424);
nor U7754 (N_7754,N_7526,N_7503);
nor U7755 (N_7755,N_7435,N_7407);
or U7756 (N_7756,N_7435,N_7509);
nor U7757 (N_7757,N_7567,N_7572);
and U7758 (N_7758,N_7449,N_7506);
nor U7759 (N_7759,N_7577,N_7596);
or U7760 (N_7760,N_7507,N_7450);
and U7761 (N_7761,N_7527,N_7563);
nor U7762 (N_7762,N_7480,N_7593);
xor U7763 (N_7763,N_7514,N_7531);
nand U7764 (N_7764,N_7586,N_7509);
xnor U7765 (N_7765,N_7420,N_7597);
nor U7766 (N_7766,N_7456,N_7492);
nand U7767 (N_7767,N_7590,N_7508);
or U7768 (N_7768,N_7437,N_7537);
nand U7769 (N_7769,N_7500,N_7529);
nor U7770 (N_7770,N_7476,N_7504);
nand U7771 (N_7771,N_7555,N_7599);
nor U7772 (N_7772,N_7598,N_7407);
nand U7773 (N_7773,N_7515,N_7429);
xnor U7774 (N_7774,N_7412,N_7497);
or U7775 (N_7775,N_7442,N_7489);
and U7776 (N_7776,N_7491,N_7430);
nand U7777 (N_7777,N_7537,N_7574);
nor U7778 (N_7778,N_7460,N_7575);
nor U7779 (N_7779,N_7465,N_7426);
nor U7780 (N_7780,N_7499,N_7447);
or U7781 (N_7781,N_7559,N_7413);
and U7782 (N_7782,N_7450,N_7432);
and U7783 (N_7783,N_7486,N_7494);
or U7784 (N_7784,N_7401,N_7453);
nor U7785 (N_7785,N_7440,N_7439);
nand U7786 (N_7786,N_7485,N_7519);
and U7787 (N_7787,N_7485,N_7511);
nor U7788 (N_7788,N_7491,N_7421);
or U7789 (N_7789,N_7525,N_7409);
or U7790 (N_7790,N_7491,N_7429);
or U7791 (N_7791,N_7448,N_7470);
or U7792 (N_7792,N_7455,N_7502);
xor U7793 (N_7793,N_7551,N_7557);
nand U7794 (N_7794,N_7563,N_7425);
xor U7795 (N_7795,N_7476,N_7427);
or U7796 (N_7796,N_7477,N_7476);
and U7797 (N_7797,N_7556,N_7498);
nand U7798 (N_7798,N_7457,N_7503);
or U7799 (N_7799,N_7467,N_7597);
nand U7800 (N_7800,N_7742,N_7688);
nor U7801 (N_7801,N_7767,N_7694);
nor U7802 (N_7802,N_7781,N_7729);
and U7803 (N_7803,N_7740,N_7621);
or U7804 (N_7804,N_7680,N_7798);
or U7805 (N_7805,N_7747,N_7749);
nor U7806 (N_7806,N_7643,N_7652);
or U7807 (N_7807,N_7610,N_7719);
or U7808 (N_7808,N_7724,N_7698);
and U7809 (N_7809,N_7774,N_7614);
nor U7810 (N_7810,N_7794,N_7615);
and U7811 (N_7811,N_7618,N_7735);
and U7812 (N_7812,N_7780,N_7681);
or U7813 (N_7813,N_7776,N_7671);
nor U7814 (N_7814,N_7653,N_7683);
xor U7815 (N_7815,N_7754,N_7715);
nor U7816 (N_7816,N_7764,N_7649);
or U7817 (N_7817,N_7674,N_7650);
nand U7818 (N_7818,N_7753,N_7668);
or U7819 (N_7819,N_7752,N_7770);
nand U7820 (N_7820,N_7775,N_7795);
and U7821 (N_7821,N_7684,N_7672);
nand U7822 (N_7822,N_7655,N_7631);
or U7823 (N_7823,N_7667,N_7604);
or U7824 (N_7824,N_7759,N_7745);
nand U7825 (N_7825,N_7708,N_7651);
nand U7826 (N_7826,N_7634,N_7760);
and U7827 (N_7827,N_7687,N_7734);
nor U7828 (N_7828,N_7706,N_7716);
nor U7829 (N_7829,N_7785,N_7758);
nor U7830 (N_7830,N_7628,N_7702);
nor U7831 (N_7831,N_7601,N_7658);
nor U7832 (N_7832,N_7721,N_7726);
and U7833 (N_7833,N_7704,N_7765);
or U7834 (N_7834,N_7748,N_7647);
or U7835 (N_7835,N_7731,N_7600);
nor U7836 (N_7836,N_7736,N_7761);
and U7837 (N_7837,N_7763,N_7642);
nand U7838 (N_7838,N_7608,N_7689);
nand U7839 (N_7839,N_7782,N_7746);
and U7840 (N_7840,N_7701,N_7697);
or U7841 (N_7841,N_7728,N_7675);
nor U7842 (N_7842,N_7640,N_7739);
and U7843 (N_7843,N_7793,N_7677);
and U7844 (N_7844,N_7654,N_7605);
and U7845 (N_7845,N_7656,N_7630);
xor U7846 (N_7846,N_7769,N_7626);
and U7847 (N_7847,N_7779,N_7703);
nor U7848 (N_7848,N_7709,N_7778);
nand U7849 (N_7849,N_7696,N_7661);
and U7850 (N_7850,N_7797,N_7788);
or U7851 (N_7851,N_7691,N_7711);
nor U7852 (N_7852,N_7730,N_7723);
nand U7853 (N_7853,N_7771,N_7641);
nand U7854 (N_7854,N_7741,N_7620);
nor U7855 (N_7855,N_7710,N_7659);
and U7856 (N_7856,N_7676,N_7606);
and U7857 (N_7857,N_7766,N_7617);
nor U7858 (N_7858,N_7602,N_7682);
or U7859 (N_7859,N_7743,N_7777);
and U7860 (N_7860,N_7638,N_7679);
nor U7861 (N_7861,N_7796,N_7693);
nand U7862 (N_7862,N_7792,N_7637);
nor U7863 (N_7863,N_7646,N_7662);
nand U7864 (N_7864,N_7648,N_7619);
nand U7865 (N_7865,N_7627,N_7609);
and U7866 (N_7866,N_7712,N_7714);
nor U7867 (N_7867,N_7664,N_7663);
nand U7868 (N_7868,N_7738,N_7612);
and U7869 (N_7869,N_7699,N_7645);
nand U7870 (N_7870,N_7666,N_7657);
or U7871 (N_7871,N_7611,N_7629);
nand U7872 (N_7872,N_7603,N_7707);
or U7873 (N_7873,N_7636,N_7690);
and U7874 (N_7874,N_7613,N_7773);
and U7875 (N_7875,N_7783,N_7633);
and U7876 (N_7876,N_7737,N_7670);
xnor U7877 (N_7877,N_7644,N_7750);
nor U7878 (N_7878,N_7607,N_7673);
nand U7879 (N_7879,N_7678,N_7727);
nand U7880 (N_7880,N_7725,N_7720);
nor U7881 (N_7881,N_7632,N_7624);
xnor U7882 (N_7882,N_7732,N_7772);
nand U7883 (N_7883,N_7660,N_7695);
xnor U7884 (N_7884,N_7705,N_7717);
nor U7885 (N_7885,N_7639,N_7756);
nand U7886 (N_7886,N_7768,N_7733);
nor U7887 (N_7887,N_7635,N_7786);
nand U7888 (N_7888,N_7784,N_7623);
nor U7889 (N_7889,N_7762,N_7789);
or U7890 (N_7890,N_7787,N_7692);
and U7891 (N_7891,N_7625,N_7665);
or U7892 (N_7892,N_7622,N_7791);
and U7893 (N_7893,N_7713,N_7616);
nand U7894 (N_7894,N_7718,N_7685);
nand U7895 (N_7895,N_7751,N_7790);
and U7896 (N_7896,N_7669,N_7722);
nand U7897 (N_7897,N_7755,N_7686);
and U7898 (N_7898,N_7744,N_7700);
or U7899 (N_7899,N_7757,N_7799);
and U7900 (N_7900,N_7707,N_7661);
xor U7901 (N_7901,N_7675,N_7768);
and U7902 (N_7902,N_7726,N_7727);
nor U7903 (N_7903,N_7696,N_7655);
and U7904 (N_7904,N_7735,N_7682);
nand U7905 (N_7905,N_7606,N_7772);
or U7906 (N_7906,N_7657,N_7650);
nor U7907 (N_7907,N_7774,N_7777);
nand U7908 (N_7908,N_7645,N_7776);
nor U7909 (N_7909,N_7715,N_7707);
or U7910 (N_7910,N_7797,N_7729);
and U7911 (N_7911,N_7663,N_7779);
nand U7912 (N_7912,N_7648,N_7731);
xnor U7913 (N_7913,N_7632,N_7637);
and U7914 (N_7914,N_7713,N_7631);
or U7915 (N_7915,N_7667,N_7734);
and U7916 (N_7916,N_7633,N_7700);
or U7917 (N_7917,N_7625,N_7687);
nor U7918 (N_7918,N_7739,N_7781);
nor U7919 (N_7919,N_7781,N_7665);
xor U7920 (N_7920,N_7771,N_7752);
nor U7921 (N_7921,N_7631,N_7626);
or U7922 (N_7922,N_7764,N_7627);
and U7923 (N_7923,N_7619,N_7631);
nand U7924 (N_7924,N_7615,N_7766);
and U7925 (N_7925,N_7650,N_7636);
and U7926 (N_7926,N_7694,N_7712);
nor U7927 (N_7927,N_7756,N_7719);
nor U7928 (N_7928,N_7682,N_7690);
or U7929 (N_7929,N_7648,N_7640);
nor U7930 (N_7930,N_7645,N_7738);
nor U7931 (N_7931,N_7787,N_7665);
and U7932 (N_7932,N_7611,N_7798);
and U7933 (N_7933,N_7639,N_7746);
nand U7934 (N_7934,N_7618,N_7798);
nand U7935 (N_7935,N_7672,N_7637);
nor U7936 (N_7936,N_7780,N_7783);
xor U7937 (N_7937,N_7746,N_7714);
or U7938 (N_7938,N_7706,N_7675);
nand U7939 (N_7939,N_7674,N_7631);
nand U7940 (N_7940,N_7722,N_7628);
nand U7941 (N_7941,N_7659,N_7771);
and U7942 (N_7942,N_7660,N_7714);
nand U7943 (N_7943,N_7691,N_7683);
or U7944 (N_7944,N_7796,N_7758);
nor U7945 (N_7945,N_7793,N_7769);
nor U7946 (N_7946,N_7746,N_7720);
or U7947 (N_7947,N_7636,N_7668);
xor U7948 (N_7948,N_7743,N_7677);
nand U7949 (N_7949,N_7609,N_7764);
nand U7950 (N_7950,N_7726,N_7663);
xor U7951 (N_7951,N_7766,N_7650);
or U7952 (N_7952,N_7662,N_7616);
nand U7953 (N_7953,N_7777,N_7608);
xnor U7954 (N_7954,N_7784,N_7665);
and U7955 (N_7955,N_7783,N_7645);
and U7956 (N_7956,N_7653,N_7716);
and U7957 (N_7957,N_7691,N_7755);
and U7958 (N_7958,N_7690,N_7696);
nor U7959 (N_7959,N_7797,N_7651);
nor U7960 (N_7960,N_7791,N_7681);
and U7961 (N_7961,N_7760,N_7715);
nor U7962 (N_7962,N_7692,N_7668);
nor U7963 (N_7963,N_7787,N_7780);
nor U7964 (N_7964,N_7773,N_7626);
nor U7965 (N_7965,N_7780,N_7669);
nor U7966 (N_7966,N_7614,N_7748);
nand U7967 (N_7967,N_7640,N_7690);
nor U7968 (N_7968,N_7742,N_7732);
and U7969 (N_7969,N_7720,N_7776);
and U7970 (N_7970,N_7737,N_7788);
and U7971 (N_7971,N_7715,N_7793);
nand U7972 (N_7972,N_7653,N_7784);
nand U7973 (N_7973,N_7666,N_7715);
xnor U7974 (N_7974,N_7708,N_7647);
and U7975 (N_7975,N_7713,N_7648);
nor U7976 (N_7976,N_7750,N_7789);
or U7977 (N_7977,N_7783,N_7771);
nor U7978 (N_7978,N_7621,N_7650);
and U7979 (N_7979,N_7641,N_7615);
nor U7980 (N_7980,N_7689,N_7660);
and U7981 (N_7981,N_7668,N_7630);
xnor U7982 (N_7982,N_7601,N_7670);
and U7983 (N_7983,N_7651,N_7727);
and U7984 (N_7984,N_7763,N_7649);
nand U7985 (N_7985,N_7617,N_7710);
and U7986 (N_7986,N_7710,N_7676);
xor U7987 (N_7987,N_7648,N_7786);
nand U7988 (N_7988,N_7671,N_7793);
and U7989 (N_7989,N_7645,N_7779);
nand U7990 (N_7990,N_7729,N_7776);
nor U7991 (N_7991,N_7631,N_7668);
nand U7992 (N_7992,N_7673,N_7747);
xnor U7993 (N_7993,N_7756,N_7606);
nor U7994 (N_7994,N_7601,N_7773);
nor U7995 (N_7995,N_7702,N_7701);
and U7996 (N_7996,N_7677,N_7629);
nor U7997 (N_7997,N_7665,N_7740);
nand U7998 (N_7998,N_7721,N_7660);
nor U7999 (N_7999,N_7785,N_7747);
nand U8000 (N_8000,N_7825,N_7935);
or U8001 (N_8001,N_7894,N_7882);
xor U8002 (N_8002,N_7998,N_7956);
nand U8003 (N_8003,N_7980,N_7858);
nor U8004 (N_8004,N_7888,N_7834);
or U8005 (N_8005,N_7969,N_7806);
and U8006 (N_8006,N_7921,N_7870);
nor U8007 (N_8007,N_7836,N_7982);
nor U8008 (N_8008,N_7846,N_7905);
nand U8009 (N_8009,N_7983,N_7810);
or U8010 (N_8010,N_7831,N_7800);
nand U8011 (N_8011,N_7920,N_7918);
nand U8012 (N_8012,N_7939,N_7829);
nor U8013 (N_8013,N_7867,N_7901);
nor U8014 (N_8014,N_7832,N_7811);
nor U8015 (N_8015,N_7840,N_7860);
or U8016 (N_8016,N_7854,N_7835);
nor U8017 (N_8017,N_7898,N_7814);
nor U8018 (N_8018,N_7885,N_7966);
and U8019 (N_8019,N_7861,N_7917);
nor U8020 (N_8020,N_7987,N_7880);
nand U8021 (N_8021,N_7812,N_7887);
nor U8022 (N_8022,N_7893,N_7927);
and U8023 (N_8023,N_7957,N_7972);
nand U8024 (N_8024,N_7938,N_7878);
xnor U8025 (N_8025,N_7974,N_7965);
nor U8026 (N_8026,N_7943,N_7967);
or U8027 (N_8027,N_7907,N_7815);
xor U8028 (N_8028,N_7890,N_7977);
and U8029 (N_8029,N_7855,N_7841);
or U8030 (N_8030,N_7820,N_7818);
or U8031 (N_8031,N_7857,N_7819);
nand U8032 (N_8032,N_7959,N_7906);
nor U8033 (N_8033,N_7940,N_7899);
nor U8034 (N_8034,N_7911,N_7902);
xor U8035 (N_8035,N_7925,N_7951);
and U8036 (N_8036,N_7884,N_7984);
or U8037 (N_8037,N_7881,N_7872);
and U8038 (N_8038,N_7994,N_7837);
nand U8039 (N_8039,N_7922,N_7838);
or U8040 (N_8040,N_7808,N_7849);
and U8041 (N_8041,N_7823,N_7942);
nand U8042 (N_8042,N_7869,N_7850);
nor U8043 (N_8043,N_7828,N_7986);
and U8044 (N_8044,N_7876,N_7801);
and U8045 (N_8045,N_7950,N_7937);
nor U8046 (N_8046,N_7891,N_7847);
nor U8047 (N_8047,N_7873,N_7991);
or U8048 (N_8048,N_7827,N_7912);
and U8049 (N_8049,N_7992,N_7839);
nor U8050 (N_8050,N_7963,N_7978);
or U8051 (N_8051,N_7822,N_7868);
or U8052 (N_8052,N_7826,N_7916);
nor U8053 (N_8053,N_7817,N_7999);
or U8054 (N_8054,N_7904,N_7923);
and U8055 (N_8055,N_7993,N_7903);
or U8056 (N_8056,N_7961,N_7946);
xnor U8057 (N_8057,N_7866,N_7976);
nor U8058 (N_8058,N_7988,N_7877);
nor U8059 (N_8059,N_7962,N_7845);
or U8060 (N_8060,N_7874,N_7804);
nor U8061 (N_8061,N_7843,N_7886);
nor U8062 (N_8062,N_7973,N_7871);
nor U8063 (N_8063,N_7809,N_7883);
or U8064 (N_8064,N_7915,N_7889);
or U8065 (N_8065,N_7944,N_7865);
nor U8066 (N_8066,N_7931,N_7953);
and U8067 (N_8067,N_7853,N_7896);
nand U8068 (N_8068,N_7919,N_7833);
nand U8069 (N_8069,N_7892,N_7821);
nand U8070 (N_8070,N_7805,N_7954);
and U8071 (N_8071,N_7930,N_7830);
or U8072 (N_8072,N_7897,N_7910);
nor U8073 (N_8073,N_7852,N_7964);
nor U8074 (N_8074,N_7803,N_7879);
nor U8075 (N_8075,N_7941,N_7948);
nor U8076 (N_8076,N_7975,N_7997);
nor U8077 (N_8077,N_7908,N_7945);
and U8078 (N_8078,N_7971,N_7802);
and U8079 (N_8079,N_7844,N_7995);
nand U8080 (N_8080,N_7813,N_7909);
nand U8081 (N_8081,N_7807,N_7932);
and U8082 (N_8082,N_7979,N_7947);
and U8083 (N_8083,N_7924,N_7862);
and U8084 (N_8084,N_7848,N_7929);
nand U8085 (N_8085,N_7816,N_7928);
xnor U8086 (N_8086,N_7842,N_7933);
nand U8087 (N_8087,N_7913,N_7958);
or U8088 (N_8088,N_7981,N_7955);
xor U8089 (N_8089,N_7952,N_7968);
and U8090 (N_8090,N_7985,N_7936);
and U8091 (N_8091,N_7859,N_7895);
or U8092 (N_8092,N_7863,N_7864);
and U8093 (N_8093,N_7856,N_7824);
nand U8094 (N_8094,N_7926,N_7934);
nor U8095 (N_8095,N_7851,N_7990);
nand U8096 (N_8096,N_7949,N_7996);
nor U8097 (N_8097,N_7914,N_7900);
or U8098 (N_8098,N_7960,N_7970);
and U8099 (N_8099,N_7989,N_7875);
xor U8100 (N_8100,N_7913,N_7943);
or U8101 (N_8101,N_7956,N_7885);
or U8102 (N_8102,N_7837,N_7810);
xor U8103 (N_8103,N_7966,N_7880);
or U8104 (N_8104,N_7908,N_7989);
nand U8105 (N_8105,N_7816,N_7801);
nor U8106 (N_8106,N_7865,N_7876);
nor U8107 (N_8107,N_7980,N_7833);
nor U8108 (N_8108,N_7917,N_7848);
xnor U8109 (N_8109,N_7973,N_7961);
nor U8110 (N_8110,N_7838,N_7820);
nor U8111 (N_8111,N_7851,N_7946);
nor U8112 (N_8112,N_7857,N_7946);
and U8113 (N_8113,N_7884,N_7959);
nor U8114 (N_8114,N_7924,N_7991);
nand U8115 (N_8115,N_7832,N_7906);
nor U8116 (N_8116,N_7886,N_7893);
nor U8117 (N_8117,N_7894,N_7840);
and U8118 (N_8118,N_7958,N_7857);
nor U8119 (N_8119,N_7843,N_7999);
nor U8120 (N_8120,N_7863,N_7997);
and U8121 (N_8121,N_7895,N_7948);
and U8122 (N_8122,N_7806,N_7827);
or U8123 (N_8123,N_7930,N_7844);
nor U8124 (N_8124,N_7998,N_7818);
nor U8125 (N_8125,N_7907,N_7859);
nand U8126 (N_8126,N_7898,N_7987);
or U8127 (N_8127,N_7922,N_7820);
nand U8128 (N_8128,N_7853,N_7970);
nand U8129 (N_8129,N_7989,N_7906);
nand U8130 (N_8130,N_7910,N_7837);
and U8131 (N_8131,N_7971,N_7981);
and U8132 (N_8132,N_7911,N_7954);
nand U8133 (N_8133,N_7941,N_7846);
xnor U8134 (N_8134,N_7903,N_7830);
nor U8135 (N_8135,N_7842,N_7817);
nand U8136 (N_8136,N_7884,N_7840);
or U8137 (N_8137,N_7838,N_7827);
nand U8138 (N_8138,N_7852,N_7990);
nand U8139 (N_8139,N_7808,N_7893);
and U8140 (N_8140,N_7847,N_7878);
xor U8141 (N_8141,N_7853,N_7847);
nand U8142 (N_8142,N_7996,N_7927);
nor U8143 (N_8143,N_7971,N_7864);
nand U8144 (N_8144,N_7822,N_7937);
or U8145 (N_8145,N_7882,N_7810);
or U8146 (N_8146,N_7870,N_7816);
nor U8147 (N_8147,N_7853,N_7811);
or U8148 (N_8148,N_7918,N_7831);
xor U8149 (N_8149,N_7904,N_7802);
or U8150 (N_8150,N_7866,N_7969);
nand U8151 (N_8151,N_7970,N_7923);
and U8152 (N_8152,N_7942,N_7979);
or U8153 (N_8153,N_7960,N_7934);
nand U8154 (N_8154,N_7926,N_7810);
nor U8155 (N_8155,N_7824,N_7897);
or U8156 (N_8156,N_7963,N_7961);
nand U8157 (N_8157,N_7931,N_7803);
xor U8158 (N_8158,N_7902,N_7984);
and U8159 (N_8159,N_7818,N_7993);
or U8160 (N_8160,N_7828,N_7911);
nand U8161 (N_8161,N_7832,N_7808);
nand U8162 (N_8162,N_7851,N_7815);
nand U8163 (N_8163,N_7934,N_7928);
nand U8164 (N_8164,N_7970,N_7850);
nor U8165 (N_8165,N_7966,N_7896);
and U8166 (N_8166,N_7990,N_7980);
or U8167 (N_8167,N_7834,N_7815);
and U8168 (N_8168,N_7871,N_7981);
nand U8169 (N_8169,N_7880,N_7860);
or U8170 (N_8170,N_7894,N_7926);
nor U8171 (N_8171,N_7997,N_7912);
nor U8172 (N_8172,N_7847,N_7981);
and U8173 (N_8173,N_7980,N_7805);
and U8174 (N_8174,N_7830,N_7946);
nand U8175 (N_8175,N_7886,N_7940);
nor U8176 (N_8176,N_7957,N_7971);
nand U8177 (N_8177,N_7814,N_7865);
nand U8178 (N_8178,N_7835,N_7907);
nand U8179 (N_8179,N_7963,N_7845);
nand U8180 (N_8180,N_7864,N_7973);
nand U8181 (N_8181,N_7963,N_7874);
or U8182 (N_8182,N_7987,N_7830);
xor U8183 (N_8183,N_7836,N_7940);
xnor U8184 (N_8184,N_7926,N_7973);
and U8185 (N_8185,N_7823,N_7909);
and U8186 (N_8186,N_7825,N_7984);
nand U8187 (N_8187,N_7994,N_7936);
xor U8188 (N_8188,N_7872,N_7941);
and U8189 (N_8189,N_7973,N_7982);
and U8190 (N_8190,N_7904,N_7827);
nor U8191 (N_8191,N_7905,N_7852);
and U8192 (N_8192,N_7835,N_7919);
and U8193 (N_8193,N_7832,N_7879);
nand U8194 (N_8194,N_7805,N_7825);
nand U8195 (N_8195,N_7901,N_7811);
and U8196 (N_8196,N_7835,N_7887);
nand U8197 (N_8197,N_7908,N_7940);
nor U8198 (N_8198,N_7883,N_7841);
nor U8199 (N_8199,N_7925,N_7912);
and U8200 (N_8200,N_8191,N_8181);
or U8201 (N_8201,N_8188,N_8137);
or U8202 (N_8202,N_8141,N_8148);
nor U8203 (N_8203,N_8083,N_8091);
xnor U8204 (N_8204,N_8089,N_8024);
or U8205 (N_8205,N_8062,N_8057);
xor U8206 (N_8206,N_8125,N_8005);
or U8207 (N_8207,N_8014,N_8072);
xnor U8208 (N_8208,N_8053,N_8006);
nand U8209 (N_8209,N_8115,N_8081);
and U8210 (N_8210,N_8047,N_8192);
or U8211 (N_8211,N_8086,N_8159);
xnor U8212 (N_8212,N_8071,N_8170);
nand U8213 (N_8213,N_8025,N_8147);
and U8214 (N_8214,N_8058,N_8002);
nor U8215 (N_8215,N_8186,N_8050);
nor U8216 (N_8216,N_8116,N_8035);
or U8217 (N_8217,N_8044,N_8160);
nor U8218 (N_8218,N_8084,N_8101);
nor U8219 (N_8219,N_8165,N_8105);
and U8220 (N_8220,N_8080,N_8133);
nand U8221 (N_8221,N_8039,N_8010);
or U8222 (N_8222,N_8135,N_8109);
and U8223 (N_8223,N_8028,N_8150);
or U8224 (N_8224,N_8004,N_8193);
nand U8225 (N_8225,N_8008,N_8177);
nor U8226 (N_8226,N_8000,N_8023);
nand U8227 (N_8227,N_8114,N_8016);
nor U8228 (N_8228,N_8164,N_8138);
nand U8229 (N_8229,N_8104,N_8056);
nand U8230 (N_8230,N_8151,N_8111);
xor U8231 (N_8231,N_8167,N_8129);
and U8232 (N_8232,N_8113,N_8027);
xnor U8233 (N_8233,N_8009,N_8187);
or U8234 (N_8234,N_8045,N_8124);
and U8235 (N_8235,N_8117,N_8197);
or U8236 (N_8236,N_8195,N_8054);
nor U8237 (N_8237,N_8065,N_8146);
xnor U8238 (N_8238,N_8041,N_8198);
xor U8239 (N_8239,N_8175,N_8019);
nor U8240 (N_8240,N_8060,N_8103);
or U8241 (N_8241,N_8055,N_8088);
nand U8242 (N_8242,N_8163,N_8048);
nor U8243 (N_8243,N_8171,N_8180);
nand U8244 (N_8244,N_8042,N_8108);
nor U8245 (N_8245,N_8153,N_8040);
nand U8246 (N_8246,N_8092,N_8136);
nand U8247 (N_8247,N_8076,N_8011);
xor U8248 (N_8248,N_8022,N_8017);
nor U8249 (N_8249,N_8095,N_8087);
nor U8250 (N_8250,N_8145,N_8026);
nand U8251 (N_8251,N_8037,N_8029);
or U8252 (N_8252,N_8033,N_8030);
and U8253 (N_8253,N_8007,N_8094);
or U8254 (N_8254,N_8110,N_8106);
nand U8255 (N_8255,N_8018,N_8099);
nor U8256 (N_8256,N_8067,N_8121);
nand U8257 (N_8257,N_8168,N_8155);
nor U8258 (N_8258,N_8070,N_8182);
nor U8259 (N_8259,N_8043,N_8140);
nand U8260 (N_8260,N_8032,N_8199);
or U8261 (N_8261,N_8185,N_8063);
and U8262 (N_8262,N_8157,N_8021);
nand U8263 (N_8263,N_8128,N_8068);
or U8264 (N_8264,N_8064,N_8038);
nand U8265 (N_8265,N_8090,N_8178);
or U8266 (N_8266,N_8196,N_8098);
nand U8267 (N_8267,N_8020,N_8012);
and U8268 (N_8268,N_8190,N_8184);
nor U8269 (N_8269,N_8085,N_8132);
or U8270 (N_8270,N_8096,N_8052);
and U8271 (N_8271,N_8173,N_8183);
nor U8272 (N_8272,N_8144,N_8162);
nand U8273 (N_8273,N_8119,N_8107);
or U8274 (N_8274,N_8066,N_8118);
and U8275 (N_8275,N_8093,N_8051);
or U8276 (N_8276,N_8156,N_8179);
or U8277 (N_8277,N_8174,N_8046);
and U8278 (N_8278,N_8134,N_8100);
xnor U8279 (N_8279,N_8130,N_8077);
or U8280 (N_8280,N_8061,N_8158);
and U8281 (N_8281,N_8127,N_8001);
nor U8282 (N_8282,N_8112,N_8143);
nor U8283 (N_8283,N_8120,N_8169);
nand U8284 (N_8284,N_8075,N_8003);
nand U8285 (N_8285,N_8049,N_8036);
nor U8286 (N_8286,N_8149,N_8069);
nor U8287 (N_8287,N_8073,N_8176);
and U8288 (N_8288,N_8194,N_8189);
and U8289 (N_8289,N_8154,N_8074);
nor U8290 (N_8290,N_8123,N_8082);
or U8291 (N_8291,N_8122,N_8079);
xnor U8292 (N_8292,N_8139,N_8015);
and U8293 (N_8293,N_8126,N_8078);
nor U8294 (N_8294,N_8161,N_8172);
nor U8295 (N_8295,N_8102,N_8034);
xor U8296 (N_8296,N_8031,N_8142);
and U8297 (N_8297,N_8059,N_8097);
nor U8298 (N_8298,N_8152,N_8166);
nor U8299 (N_8299,N_8013,N_8131);
nor U8300 (N_8300,N_8016,N_8044);
nor U8301 (N_8301,N_8029,N_8160);
nand U8302 (N_8302,N_8191,N_8137);
nor U8303 (N_8303,N_8157,N_8046);
xnor U8304 (N_8304,N_8055,N_8144);
nand U8305 (N_8305,N_8155,N_8170);
and U8306 (N_8306,N_8030,N_8123);
xor U8307 (N_8307,N_8103,N_8112);
nand U8308 (N_8308,N_8067,N_8010);
nand U8309 (N_8309,N_8188,N_8013);
and U8310 (N_8310,N_8162,N_8125);
and U8311 (N_8311,N_8059,N_8021);
nor U8312 (N_8312,N_8148,N_8068);
nand U8313 (N_8313,N_8028,N_8165);
nand U8314 (N_8314,N_8148,N_8156);
nand U8315 (N_8315,N_8070,N_8183);
nand U8316 (N_8316,N_8079,N_8163);
and U8317 (N_8317,N_8098,N_8138);
nor U8318 (N_8318,N_8060,N_8190);
or U8319 (N_8319,N_8143,N_8077);
xor U8320 (N_8320,N_8015,N_8154);
or U8321 (N_8321,N_8153,N_8063);
nor U8322 (N_8322,N_8174,N_8062);
xor U8323 (N_8323,N_8088,N_8003);
and U8324 (N_8324,N_8124,N_8154);
and U8325 (N_8325,N_8063,N_8135);
or U8326 (N_8326,N_8147,N_8178);
nor U8327 (N_8327,N_8029,N_8117);
nor U8328 (N_8328,N_8015,N_8007);
nand U8329 (N_8329,N_8180,N_8132);
nor U8330 (N_8330,N_8009,N_8114);
and U8331 (N_8331,N_8064,N_8109);
or U8332 (N_8332,N_8040,N_8058);
and U8333 (N_8333,N_8045,N_8039);
nor U8334 (N_8334,N_8020,N_8178);
nand U8335 (N_8335,N_8102,N_8122);
nor U8336 (N_8336,N_8114,N_8170);
xnor U8337 (N_8337,N_8007,N_8062);
nor U8338 (N_8338,N_8092,N_8143);
and U8339 (N_8339,N_8086,N_8037);
nor U8340 (N_8340,N_8132,N_8044);
nand U8341 (N_8341,N_8080,N_8068);
nor U8342 (N_8342,N_8013,N_8136);
nand U8343 (N_8343,N_8072,N_8037);
nand U8344 (N_8344,N_8145,N_8093);
nand U8345 (N_8345,N_8177,N_8006);
nor U8346 (N_8346,N_8037,N_8096);
and U8347 (N_8347,N_8054,N_8124);
nand U8348 (N_8348,N_8025,N_8079);
or U8349 (N_8349,N_8064,N_8031);
and U8350 (N_8350,N_8018,N_8188);
or U8351 (N_8351,N_8082,N_8041);
and U8352 (N_8352,N_8001,N_8179);
nand U8353 (N_8353,N_8087,N_8022);
and U8354 (N_8354,N_8080,N_8053);
or U8355 (N_8355,N_8097,N_8179);
or U8356 (N_8356,N_8011,N_8106);
nand U8357 (N_8357,N_8090,N_8109);
nor U8358 (N_8358,N_8143,N_8182);
and U8359 (N_8359,N_8033,N_8178);
xnor U8360 (N_8360,N_8029,N_8126);
nand U8361 (N_8361,N_8107,N_8004);
xor U8362 (N_8362,N_8122,N_8167);
nor U8363 (N_8363,N_8026,N_8030);
or U8364 (N_8364,N_8014,N_8107);
and U8365 (N_8365,N_8115,N_8116);
or U8366 (N_8366,N_8089,N_8159);
nand U8367 (N_8367,N_8107,N_8118);
nand U8368 (N_8368,N_8074,N_8016);
nor U8369 (N_8369,N_8029,N_8010);
nor U8370 (N_8370,N_8185,N_8010);
or U8371 (N_8371,N_8014,N_8018);
nand U8372 (N_8372,N_8046,N_8132);
or U8373 (N_8373,N_8180,N_8028);
nand U8374 (N_8374,N_8074,N_8147);
and U8375 (N_8375,N_8171,N_8054);
and U8376 (N_8376,N_8124,N_8014);
or U8377 (N_8377,N_8108,N_8068);
nand U8378 (N_8378,N_8017,N_8175);
nor U8379 (N_8379,N_8025,N_8055);
nand U8380 (N_8380,N_8161,N_8198);
nand U8381 (N_8381,N_8130,N_8175);
and U8382 (N_8382,N_8055,N_8149);
nor U8383 (N_8383,N_8050,N_8017);
and U8384 (N_8384,N_8058,N_8145);
nor U8385 (N_8385,N_8151,N_8065);
or U8386 (N_8386,N_8061,N_8110);
nor U8387 (N_8387,N_8098,N_8059);
or U8388 (N_8388,N_8187,N_8068);
and U8389 (N_8389,N_8078,N_8100);
and U8390 (N_8390,N_8044,N_8147);
or U8391 (N_8391,N_8030,N_8189);
nor U8392 (N_8392,N_8125,N_8038);
nor U8393 (N_8393,N_8003,N_8048);
nand U8394 (N_8394,N_8016,N_8158);
and U8395 (N_8395,N_8030,N_8083);
and U8396 (N_8396,N_8045,N_8151);
nand U8397 (N_8397,N_8172,N_8176);
xnor U8398 (N_8398,N_8034,N_8126);
nor U8399 (N_8399,N_8022,N_8077);
nand U8400 (N_8400,N_8388,N_8276);
nor U8401 (N_8401,N_8362,N_8245);
and U8402 (N_8402,N_8286,N_8299);
xor U8403 (N_8403,N_8216,N_8374);
xor U8404 (N_8404,N_8230,N_8229);
nor U8405 (N_8405,N_8351,N_8312);
xor U8406 (N_8406,N_8342,N_8328);
and U8407 (N_8407,N_8316,N_8205);
nand U8408 (N_8408,N_8244,N_8259);
nor U8409 (N_8409,N_8284,N_8211);
or U8410 (N_8410,N_8266,N_8214);
nand U8411 (N_8411,N_8338,N_8355);
nor U8412 (N_8412,N_8354,N_8203);
and U8413 (N_8413,N_8232,N_8309);
or U8414 (N_8414,N_8201,N_8285);
xor U8415 (N_8415,N_8277,N_8310);
or U8416 (N_8416,N_8369,N_8335);
nor U8417 (N_8417,N_8218,N_8290);
xnor U8418 (N_8418,N_8255,N_8327);
nand U8419 (N_8419,N_8225,N_8297);
nor U8420 (N_8420,N_8340,N_8343);
nand U8421 (N_8421,N_8261,N_8359);
nand U8422 (N_8422,N_8248,N_8206);
nor U8423 (N_8423,N_8293,N_8386);
and U8424 (N_8424,N_8283,N_8372);
and U8425 (N_8425,N_8243,N_8358);
or U8426 (N_8426,N_8300,N_8302);
nor U8427 (N_8427,N_8282,N_8397);
nor U8428 (N_8428,N_8375,N_8376);
and U8429 (N_8429,N_8356,N_8249);
and U8430 (N_8430,N_8365,N_8332);
nor U8431 (N_8431,N_8281,N_8237);
nand U8432 (N_8432,N_8287,N_8242);
nor U8433 (N_8433,N_8220,N_8320);
xor U8434 (N_8434,N_8348,N_8315);
or U8435 (N_8435,N_8268,N_8322);
nor U8436 (N_8436,N_8326,N_8321);
or U8437 (N_8437,N_8208,N_8257);
nor U8438 (N_8438,N_8250,N_8274);
nand U8439 (N_8439,N_8398,N_8391);
nand U8440 (N_8440,N_8384,N_8238);
nand U8441 (N_8441,N_8381,N_8223);
and U8442 (N_8442,N_8380,N_8373);
nor U8443 (N_8443,N_8377,N_8221);
or U8444 (N_8444,N_8331,N_8213);
nor U8445 (N_8445,N_8395,N_8270);
or U8446 (N_8446,N_8260,N_8217);
nand U8447 (N_8447,N_8364,N_8215);
and U8448 (N_8448,N_8334,N_8325);
and U8449 (N_8449,N_8247,N_8361);
and U8450 (N_8450,N_8269,N_8234);
nand U8451 (N_8451,N_8378,N_8280);
and U8452 (N_8452,N_8367,N_8265);
and U8453 (N_8453,N_8289,N_8324);
or U8454 (N_8454,N_8251,N_8212);
nand U8455 (N_8455,N_8313,N_8389);
or U8456 (N_8456,N_8308,N_8288);
or U8457 (N_8457,N_8228,N_8204);
and U8458 (N_8458,N_8279,N_8319);
nand U8459 (N_8459,N_8368,N_8371);
nor U8460 (N_8460,N_8360,N_8379);
nand U8461 (N_8461,N_8239,N_8382);
nand U8462 (N_8462,N_8267,N_8254);
and U8463 (N_8463,N_8291,N_8262);
nor U8464 (N_8464,N_8390,N_8329);
and U8465 (N_8465,N_8207,N_8200);
nor U8466 (N_8466,N_8258,N_8275);
and U8467 (N_8467,N_8305,N_8271);
and U8468 (N_8468,N_8210,N_8311);
or U8469 (N_8469,N_8253,N_8241);
and U8470 (N_8470,N_8346,N_8263);
xor U8471 (N_8471,N_8352,N_8273);
nor U8472 (N_8472,N_8303,N_8256);
and U8473 (N_8473,N_8350,N_8347);
and U8474 (N_8474,N_8240,N_8252);
nor U8475 (N_8475,N_8317,N_8387);
xnor U8476 (N_8476,N_8222,N_8370);
nor U8477 (N_8477,N_8341,N_8383);
nor U8478 (N_8478,N_8344,N_8314);
and U8479 (N_8479,N_8399,N_8323);
nor U8480 (N_8480,N_8219,N_8233);
or U8481 (N_8481,N_8396,N_8294);
nor U8482 (N_8482,N_8278,N_8363);
nor U8483 (N_8483,N_8304,N_8236);
and U8484 (N_8484,N_8209,N_8353);
or U8485 (N_8485,N_8392,N_8337);
and U8486 (N_8486,N_8272,N_8227);
nor U8487 (N_8487,N_8345,N_8296);
or U8488 (N_8488,N_8226,N_8306);
or U8489 (N_8489,N_8246,N_8318);
and U8490 (N_8490,N_8385,N_8292);
or U8491 (N_8491,N_8224,N_8357);
nand U8492 (N_8492,N_8295,N_8330);
and U8493 (N_8493,N_8393,N_8307);
or U8494 (N_8494,N_8264,N_8333);
or U8495 (N_8495,N_8298,N_8231);
nor U8496 (N_8496,N_8394,N_8235);
nand U8497 (N_8497,N_8339,N_8366);
and U8498 (N_8498,N_8349,N_8336);
or U8499 (N_8499,N_8301,N_8202);
xnor U8500 (N_8500,N_8212,N_8360);
and U8501 (N_8501,N_8283,N_8395);
or U8502 (N_8502,N_8273,N_8302);
and U8503 (N_8503,N_8217,N_8239);
and U8504 (N_8504,N_8296,N_8205);
nand U8505 (N_8505,N_8342,N_8324);
or U8506 (N_8506,N_8327,N_8307);
nor U8507 (N_8507,N_8288,N_8269);
and U8508 (N_8508,N_8215,N_8246);
and U8509 (N_8509,N_8346,N_8356);
nor U8510 (N_8510,N_8326,N_8314);
nand U8511 (N_8511,N_8243,N_8368);
xor U8512 (N_8512,N_8264,N_8318);
nand U8513 (N_8513,N_8387,N_8300);
nand U8514 (N_8514,N_8320,N_8205);
xor U8515 (N_8515,N_8305,N_8366);
or U8516 (N_8516,N_8278,N_8247);
and U8517 (N_8517,N_8308,N_8206);
nor U8518 (N_8518,N_8206,N_8205);
and U8519 (N_8519,N_8356,N_8384);
and U8520 (N_8520,N_8279,N_8229);
nor U8521 (N_8521,N_8201,N_8267);
nor U8522 (N_8522,N_8244,N_8333);
xnor U8523 (N_8523,N_8280,N_8248);
nand U8524 (N_8524,N_8306,N_8257);
or U8525 (N_8525,N_8325,N_8393);
nand U8526 (N_8526,N_8211,N_8355);
nor U8527 (N_8527,N_8374,N_8250);
and U8528 (N_8528,N_8290,N_8279);
nor U8529 (N_8529,N_8307,N_8353);
xor U8530 (N_8530,N_8364,N_8338);
xnor U8531 (N_8531,N_8380,N_8342);
nand U8532 (N_8532,N_8347,N_8209);
nor U8533 (N_8533,N_8302,N_8281);
xnor U8534 (N_8534,N_8364,N_8201);
and U8535 (N_8535,N_8283,N_8256);
or U8536 (N_8536,N_8384,N_8304);
xor U8537 (N_8537,N_8322,N_8269);
nor U8538 (N_8538,N_8387,N_8250);
or U8539 (N_8539,N_8284,N_8219);
xor U8540 (N_8540,N_8235,N_8290);
or U8541 (N_8541,N_8385,N_8220);
xnor U8542 (N_8542,N_8232,N_8368);
and U8543 (N_8543,N_8204,N_8351);
or U8544 (N_8544,N_8219,N_8257);
nand U8545 (N_8545,N_8297,N_8336);
xnor U8546 (N_8546,N_8245,N_8208);
or U8547 (N_8547,N_8340,N_8346);
and U8548 (N_8548,N_8356,N_8214);
and U8549 (N_8549,N_8371,N_8229);
or U8550 (N_8550,N_8275,N_8257);
nand U8551 (N_8551,N_8321,N_8304);
nand U8552 (N_8552,N_8216,N_8225);
or U8553 (N_8553,N_8399,N_8306);
nor U8554 (N_8554,N_8270,N_8281);
or U8555 (N_8555,N_8395,N_8223);
nand U8556 (N_8556,N_8354,N_8351);
nor U8557 (N_8557,N_8245,N_8218);
and U8558 (N_8558,N_8260,N_8274);
nand U8559 (N_8559,N_8303,N_8236);
or U8560 (N_8560,N_8258,N_8236);
nor U8561 (N_8561,N_8315,N_8242);
xnor U8562 (N_8562,N_8383,N_8301);
or U8563 (N_8563,N_8334,N_8226);
nor U8564 (N_8564,N_8378,N_8302);
and U8565 (N_8565,N_8270,N_8299);
nand U8566 (N_8566,N_8229,N_8359);
or U8567 (N_8567,N_8245,N_8327);
xnor U8568 (N_8568,N_8277,N_8362);
and U8569 (N_8569,N_8202,N_8286);
and U8570 (N_8570,N_8385,N_8315);
xnor U8571 (N_8571,N_8218,N_8219);
nand U8572 (N_8572,N_8244,N_8201);
and U8573 (N_8573,N_8353,N_8335);
and U8574 (N_8574,N_8260,N_8288);
or U8575 (N_8575,N_8333,N_8367);
nand U8576 (N_8576,N_8354,N_8320);
nor U8577 (N_8577,N_8215,N_8367);
or U8578 (N_8578,N_8325,N_8295);
xor U8579 (N_8579,N_8255,N_8215);
and U8580 (N_8580,N_8262,N_8248);
nand U8581 (N_8581,N_8267,N_8345);
xor U8582 (N_8582,N_8396,N_8267);
nor U8583 (N_8583,N_8221,N_8312);
nor U8584 (N_8584,N_8377,N_8218);
and U8585 (N_8585,N_8274,N_8297);
nand U8586 (N_8586,N_8284,N_8372);
nand U8587 (N_8587,N_8258,N_8398);
or U8588 (N_8588,N_8238,N_8315);
nor U8589 (N_8589,N_8273,N_8366);
nand U8590 (N_8590,N_8301,N_8314);
or U8591 (N_8591,N_8254,N_8219);
xor U8592 (N_8592,N_8221,N_8269);
nor U8593 (N_8593,N_8381,N_8315);
nor U8594 (N_8594,N_8337,N_8388);
and U8595 (N_8595,N_8275,N_8387);
nand U8596 (N_8596,N_8332,N_8355);
or U8597 (N_8597,N_8214,N_8334);
nand U8598 (N_8598,N_8215,N_8358);
nand U8599 (N_8599,N_8291,N_8207);
nor U8600 (N_8600,N_8599,N_8414);
or U8601 (N_8601,N_8401,N_8403);
nand U8602 (N_8602,N_8421,N_8438);
or U8603 (N_8603,N_8475,N_8565);
xor U8604 (N_8604,N_8425,N_8545);
and U8605 (N_8605,N_8494,N_8529);
and U8606 (N_8606,N_8479,N_8544);
or U8607 (N_8607,N_8525,N_8463);
nand U8608 (N_8608,N_8484,N_8568);
nor U8609 (N_8609,N_8464,N_8528);
nand U8610 (N_8610,N_8572,N_8509);
or U8611 (N_8611,N_8555,N_8570);
xnor U8612 (N_8612,N_8411,N_8596);
or U8613 (N_8613,N_8523,N_8473);
nand U8614 (N_8614,N_8504,N_8554);
and U8615 (N_8615,N_8478,N_8448);
xor U8616 (N_8616,N_8583,N_8417);
nor U8617 (N_8617,N_8501,N_8513);
xor U8618 (N_8618,N_8569,N_8502);
nor U8619 (N_8619,N_8433,N_8452);
nand U8620 (N_8620,N_8423,N_8587);
or U8621 (N_8621,N_8576,N_8486);
nor U8622 (N_8622,N_8437,N_8493);
and U8623 (N_8623,N_8500,N_8506);
nor U8624 (N_8624,N_8512,N_8558);
xor U8625 (N_8625,N_8469,N_8434);
or U8626 (N_8626,N_8514,N_8424);
or U8627 (N_8627,N_8520,N_8440);
and U8628 (N_8628,N_8540,N_8499);
nand U8629 (N_8629,N_8563,N_8518);
or U8630 (N_8630,N_8598,N_8496);
nor U8631 (N_8631,N_8562,N_8412);
or U8632 (N_8632,N_8508,N_8553);
and U8633 (N_8633,N_8453,N_8560);
nand U8634 (N_8634,N_8515,N_8455);
nand U8635 (N_8635,N_8483,N_8409);
and U8636 (N_8636,N_8505,N_8461);
nor U8637 (N_8637,N_8591,N_8444);
and U8638 (N_8638,N_8597,N_8435);
nor U8639 (N_8639,N_8441,N_8405);
and U8640 (N_8640,N_8510,N_8533);
or U8641 (N_8641,N_8460,N_8549);
and U8642 (N_8642,N_8428,N_8404);
and U8643 (N_8643,N_8446,N_8431);
nor U8644 (N_8644,N_8419,N_8556);
or U8645 (N_8645,N_8450,N_8491);
nand U8646 (N_8646,N_8482,N_8575);
nor U8647 (N_8647,N_8407,N_8548);
and U8648 (N_8648,N_8402,N_8420);
nor U8649 (N_8649,N_8481,N_8588);
nand U8650 (N_8650,N_8527,N_8586);
nor U8651 (N_8651,N_8443,N_8526);
or U8652 (N_8652,N_8467,N_8517);
and U8653 (N_8653,N_8559,N_8507);
nor U8654 (N_8654,N_8480,N_8427);
or U8655 (N_8655,N_8577,N_8477);
or U8656 (N_8656,N_8538,N_8497);
nor U8657 (N_8657,N_8445,N_8571);
nor U8658 (N_8658,N_8487,N_8524);
and U8659 (N_8659,N_8580,N_8539);
or U8660 (N_8660,N_8485,N_8415);
and U8661 (N_8661,N_8451,N_8408);
nor U8662 (N_8662,N_8418,N_8489);
xor U8663 (N_8663,N_8436,N_8457);
and U8664 (N_8664,N_8537,N_8400);
xnor U8665 (N_8665,N_8456,N_8566);
and U8666 (N_8666,N_8594,N_8578);
and U8667 (N_8667,N_8521,N_8466);
and U8668 (N_8668,N_8536,N_8474);
nor U8669 (N_8669,N_8574,N_8593);
xor U8670 (N_8670,N_8561,N_8582);
or U8671 (N_8671,N_8429,N_8595);
or U8672 (N_8672,N_8552,N_8476);
and U8673 (N_8673,N_8426,N_8532);
nor U8674 (N_8674,N_8488,N_8585);
nand U8675 (N_8675,N_8590,N_8522);
or U8676 (N_8676,N_8542,N_8470);
or U8677 (N_8677,N_8511,N_8458);
or U8678 (N_8678,N_8541,N_8406);
xor U8679 (N_8679,N_8495,N_8432);
and U8680 (N_8680,N_8430,N_8573);
and U8681 (N_8681,N_8592,N_8519);
or U8682 (N_8682,N_8550,N_8547);
nand U8683 (N_8683,N_8449,N_8557);
nor U8684 (N_8684,N_8459,N_8490);
and U8685 (N_8685,N_8471,N_8465);
nand U8686 (N_8686,N_8454,N_8551);
and U8687 (N_8687,N_8564,N_8534);
and U8688 (N_8688,N_8439,N_8498);
or U8689 (N_8689,N_8535,N_8472);
and U8690 (N_8690,N_8422,N_8413);
and U8691 (N_8691,N_8410,N_8567);
nand U8692 (N_8692,N_8584,N_8531);
nand U8693 (N_8693,N_8579,N_8442);
and U8694 (N_8694,N_8416,N_8589);
nand U8695 (N_8695,N_8462,N_8546);
xnor U8696 (N_8696,N_8516,N_8492);
and U8697 (N_8697,N_8543,N_8581);
nor U8698 (N_8698,N_8530,N_8503);
xnor U8699 (N_8699,N_8447,N_8468);
nand U8700 (N_8700,N_8596,N_8425);
nor U8701 (N_8701,N_8495,N_8449);
or U8702 (N_8702,N_8552,N_8461);
xnor U8703 (N_8703,N_8542,N_8477);
nand U8704 (N_8704,N_8430,N_8473);
or U8705 (N_8705,N_8470,N_8458);
and U8706 (N_8706,N_8449,N_8475);
xnor U8707 (N_8707,N_8429,N_8404);
nor U8708 (N_8708,N_8446,N_8574);
nor U8709 (N_8709,N_8554,N_8474);
nor U8710 (N_8710,N_8444,N_8501);
nor U8711 (N_8711,N_8504,N_8460);
nor U8712 (N_8712,N_8547,N_8480);
and U8713 (N_8713,N_8544,N_8524);
xor U8714 (N_8714,N_8409,N_8464);
nand U8715 (N_8715,N_8407,N_8411);
nand U8716 (N_8716,N_8454,N_8564);
nor U8717 (N_8717,N_8529,N_8561);
nand U8718 (N_8718,N_8425,N_8593);
nor U8719 (N_8719,N_8516,N_8478);
and U8720 (N_8720,N_8416,N_8559);
or U8721 (N_8721,N_8442,N_8494);
nor U8722 (N_8722,N_8540,N_8537);
or U8723 (N_8723,N_8584,N_8408);
nor U8724 (N_8724,N_8483,N_8598);
nand U8725 (N_8725,N_8527,N_8512);
nor U8726 (N_8726,N_8553,N_8550);
and U8727 (N_8727,N_8543,N_8461);
and U8728 (N_8728,N_8462,N_8484);
and U8729 (N_8729,N_8599,N_8562);
nor U8730 (N_8730,N_8558,N_8588);
and U8731 (N_8731,N_8403,N_8420);
and U8732 (N_8732,N_8551,N_8582);
and U8733 (N_8733,N_8462,N_8431);
nand U8734 (N_8734,N_8583,N_8406);
and U8735 (N_8735,N_8499,N_8415);
and U8736 (N_8736,N_8453,N_8486);
nor U8737 (N_8737,N_8577,N_8473);
nor U8738 (N_8738,N_8556,N_8596);
or U8739 (N_8739,N_8428,N_8590);
or U8740 (N_8740,N_8588,N_8520);
or U8741 (N_8741,N_8585,N_8550);
or U8742 (N_8742,N_8435,N_8532);
nand U8743 (N_8743,N_8427,N_8488);
nor U8744 (N_8744,N_8514,N_8448);
nor U8745 (N_8745,N_8474,N_8569);
nand U8746 (N_8746,N_8432,N_8581);
nor U8747 (N_8747,N_8542,N_8512);
or U8748 (N_8748,N_8472,N_8538);
or U8749 (N_8749,N_8525,N_8407);
nand U8750 (N_8750,N_8409,N_8530);
nand U8751 (N_8751,N_8403,N_8468);
and U8752 (N_8752,N_8488,N_8524);
xnor U8753 (N_8753,N_8411,N_8552);
nor U8754 (N_8754,N_8413,N_8450);
and U8755 (N_8755,N_8524,N_8448);
nor U8756 (N_8756,N_8463,N_8473);
and U8757 (N_8757,N_8528,N_8453);
nand U8758 (N_8758,N_8457,N_8485);
nor U8759 (N_8759,N_8576,N_8401);
nand U8760 (N_8760,N_8439,N_8538);
and U8761 (N_8761,N_8513,N_8531);
xor U8762 (N_8762,N_8434,N_8476);
and U8763 (N_8763,N_8590,N_8404);
nand U8764 (N_8764,N_8527,N_8545);
xnor U8765 (N_8765,N_8427,N_8589);
xor U8766 (N_8766,N_8500,N_8515);
or U8767 (N_8767,N_8425,N_8503);
xnor U8768 (N_8768,N_8465,N_8435);
xnor U8769 (N_8769,N_8429,N_8457);
and U8770 (N_8770,N_8509,N_8518);
nor U8771 (N_8771,N_8455,N_8492);
and U8772 (N_8772,N_8512,N_8572);
nand U8773 (N_8773,N_8545,N_8407);
nor U8774 (N_8774,N_8574,N_8410);
nor U8775 (N_8775,N_8426,N_8496);
or U8776 (N_8776,N_8461,N_8562);
nand U8777 (N_8777,N_8585,N_8479);
nor U8778 (N_8778,N_8598,N_8424);
or U8779 (N_8779,N_8504,N_8506);
nand U8780 (N_8780,N_8416,N_8455);
or U8781 (N_8781,N_8432,N_8491);
nor U8782 (N_8782,N_8409,N_8412);
and U8783 (N_8783,N_8403,N_8492);
nand U8784 (N_8784,N_8501,N_8489);
or U8785 (N_8785,N_8407,N_8466);
and U8786 (N_8786,N_8517,N_8453);
nand U8787 (N_8787,N_8536,N_8442);
nand U8788 (N_8788,N_8445,N_8401);
xor U8789 (N_8789,N_8590,N_8532);
and U8790 (N_8790,N_8501,N_8427);
nor U8791 (N_8791,N_8430,N_8543);
nand U8792 (N_8792,N_8446,N_8404);
and U8793 (N_8793,N_8456,N_8405);
xor U8794 (N_8794,N_8508,N_8524);
and U8795 (N_8795,N_8552,N_8475);
and U8796 (N_8796,N_8479,N_8517);
and U8797 (N_8797,N_8599,N_8486);
or U8798 (N_8798,N_8465,N_8556);
xnor U8799 (N_8799,N_8590,N_8579);
and U8800 (N_8800,N_8628,N_8668);
nand U8801 (N_8801,N_8649,N_8602);
nand U8802 (N_8802,N_8630,N_8690);
and U8803 (N_8803,N_8691,N_8638);
nand U8804 (N_8804,N_8794,N_8744);
nor U8805 (N_8805,N_8639,N_8656);
or U8806 (N_8806,N_8783,N_8686);
or U8807 (N_8807,N_8688,N_8616);
nand U8808 (N_8808,N_8615,N_8623);
and U8809 (N_8809,N_8696,N_8787);
xnor U8810 (N_8810,N_8746,N_8606);
and U8811 (N_8811,N_8678,N_8663);
xor U8812 (N_8812,N_8689,N_8665);
and U8813 (N_8813,N_8661,N_8728);
and U8814 (N_8814,N_8733,N_8666);
nand U8815 (N_8815,N_8621,N_8693);
nand U8816 (N_8816,N_8618,N_8612);
and U8817 (N_8817,N_8782,N_8667);
xor U8818 (N_8818,N_8731,N_8720);
or U8819 (N_8819,N_8613,N_8799);
or U8820 (N_8820,N_8694,N_8709);
or U8821 (N_8821,N_8756,N_8772);
and U8822 (N_8822,N_8722,N_8626);
nor U8823 (N_8823,N_8672,N_8622);
or U8824 (N_8824,N_8695,N_8673);
or U8825 (N_8825,N_8645,N_8675);
or U8826 (N_8826,N_8614,N_8767);
and U8827 (N_8827,N_8788,N_8635);
nand U8828 (N_8828,N_8797,N_8617);
nand U8829 (N_8829,N_8711,N_8798);
xnor U8830 (N_8830,N_8710,N_8679);
and U8831 (N_8831,N_8732,N_8781);
nor U8832 (N_8832,N_8779,N_8729);
nand U8833 (N_8833,N_8701,N_8723);
nor U8834 (N_8834,N_8726,N_8771);
nor U8835 (N_8835,N_8790,N_8662);
or U8836 (N_8836,N_8766,N_8719);
or U8837 (N_8837,N_8780,N_8743);
and U8838 (N_8838,N_8795,N_8727);
nand U8839 (N_8839,N_8741,N_8785);
xor U8840 (N_8840,N_8793,N_8611);
and U8841 (N_8841,N_8627,N_8759);
or U8842 (N_8842,N_8633,N_8708);
nor U8843 (N_8843,N_8704,N_8637);
nor U8844 (N_8844,N_8601,N_8674);
nand U8845 (N_8845,N_8715,N_8653);
xnor U8846 (N_8846,N_8684,N_8629);
nor U8847 (N_8847,N_8681,N_8713);
xor U8848 (N_8848,N_8647,N_8640);
or U8849 (N_8849,N_8625,N_8761);
or U8850 (N_8850,N_8754,N_8676);
and U8851 (N_8851,N_8700,N_8740);
nand U8852 (N_8852,N_8654,N_8610);
or U8853 (N_8853,N_8739,N_8671);
nor U8854 (N_8854,N_8619,N_8725);
nor U8855 (N_8855,N_8669,N_8774);
and U8856 (N_8856,N_8692,N_8760);
nor U8857 (N_8857,N_8636,N_8791);
xnor U8858 (N_8858,N_8605,N_8765);
nand U8859 (N_8859,N_8670,N_8603);
nand U8860 (N_8860,N_8737,N_8757);
and U8861 (N_8861,N_8697,N_8677);
and U8862 (N_8862,N_8792,N_8604);
or U8863 (N_8863,N_8648,N_8655);
or U8864 (N_8864,N_8748,N_8770);
or U8865 (N_8865,N_8706,N_8718);
nor U8866 (N_8866,N_8776,N_8769);
and U8867 (N_8867,N_8724,N_8608);
nand U8868 (N_8868,N_8784,N_8751);
and U8869 (N_8869,N_8753,N_8607);
nor U8870 (N_8870,N_8703,N_8763);
or U8871 (N_8871,N_8721,N_8735);
and U8872 (N_8872,N_8624,N_8600);
or U8873 (N_8873,N_8683,N_8747);
and U8874 (N_8874,N_8702,N_8699);
or U8875 (N_8875,N_8762,N_8730);
nand U8876 (N_8876,N_8657,N_8644);
nor U8877 (N_8877,N_8752,N_8712);
nor U8878 (N_8878,N_8789,N_8717);
and U8879 (N_8879,N_8750,N_8716);
nand U8880 (N_8880,N_8609,N_8632);
and U8881 (N_8881,N_8734,N_8664);
nand U8882 (N_8882,N_8778,N_8659);
or U8883 (N_8883,N_8738,N_8651);
or U8884 (N_8884,N_8742,N_8641);
and U8885 (N_8885,N_8773,N_8643);
nor U8886 (N_8886,N_8687,N_8685);
nor U8887 (N_8887,N_8777,N_8646);
and U8888 (N_8888,N_8745,N_8642);
or U8889 (N_8889,N_8620,N_8658);
nand U8890 (N_8890,N_8768,N_8758);
nand U8891 (N_8891,N_8749,N_8652);
nor U8892 (N_8892,N_8705,N_8634);
nand U8893 (N_8893,N_8714,N_8755);
nand U8894 (N_8894,N_8736,N_8786);
and U8895 (N_8895,N_8796,N_8764);
or U8896 (N_8896,N_8775,N_8650);
nand U8897 (N_8897,N_8682,N_8707);
and U8898 (N_8898,N_8680,N_8698);
nand U8899 (N_8899,N_8660,N_8631);
nor U8900 (N_8900,N_8741,N_8682);
nor U8901 (N_8901,N_8698,N_8795);
nand U8902 (N_8902,N_8719,N_8640);
or U8903 (N_8903,N_8670,N_8649);
nand U8904 (N_8904,N_8764,N_8799);
nand U8905 (N_8905,N_8669,N_8798);
xnor U8906 (N_8906,N_8785,N_8706);
nor U8907 (N_8907,N_8691,N_8672);
and U8908 (N_8908,N_8697,N_8629);
nor U8909 (N_8909,N_8658,N_8681);
or U8910 (N_8910,N_8760,N_8650);
and U8911 (N_8911,N_8775,N_8762);
nand U8912 (N_8912,N_8725,N_8747);
or U8913 (N_8913,N_8691,N_8701);
nand U8914 (N_8914,N_8654,N_8755);
nand U8915 (N_8915,N_8610,N_8797);
nand U8916 (N_8916,N_8614,N_8650);
nand U8917 (N_8917,N_8658,N_8715);
nor U8918 (N_8918,N_8655,N_8741);
nor U8919 (N_8919,N_8701,N_8634);
and U8920 (N_8920,N_8746,N_8739);
nand U8921 (N_8921,N_8707,N_8696);
and U8922 (N_8922,N_8600,N_8673);
or U8923 (N_8923,N_8744,N_8644);
xor U8924 (N_8924,N_8696,N_8739);
nand U8925 (N_8925,N_8624,N_8691);
or U8926 (N_8926,N_8661,N_8795);
nand U8927 (N_8927,N_8601,N_8766);
nand U8928 (N_8928,N_8649,N_8677);
nor U8929 (N_8929,N_8715,N_8762);
nor U8930 (N_8930,N_8769,N_8709);
nand U8931 (N_8931,N_8767,N_8600);
and U8932 (N_8932,N_8676,N_8684);
xnor U8933 (N_8933,N_8778,N_8668);
and U8934 (N_8934,N_8672,N_8642);
nor U8935 (N_8935,N_8790,N_8615);
or U8936 (N_8936,N_8782,N_8642);
or U8937 (N_8937,N_8762,N_8663);
or U8938 (N_8938,N_8722,N_8792);
and U8939 (N_8939,N_8662,N_8754);
nand U8940 (N_8940,N_8681,N_8778);
and U8941 (N_8941,N_8608,N_8747);
and U8942 (N_8942,N_8603,N_8755);
nand U8943 (N_8943,N_8770,N_8653);
or U8944 (N_8944,N_8647,N_8770);
or U8945 (N_8945,N_8667,N_8608);
xnor U8946 (N_8946,N_8690,N_8732);
nand U8947 (N_8947,N_8647,N_8793);
or U8948 (N_8948,N_8629,N_8751);
nor U8949 (N_8949,N_8650,N_8712);
and U8950 (N_8950,N_8625,N_8769);
nor U8951 (N_8951,N_8789,N_8708);
nand U8952 (N_8952,N_8642,N_8641);
nand U8953 (N_8953,N_8745,N_8687);
nand U8954 (N_8954,N_8711,N_8750);
and U8955 (N_8955,N_8697,N_8610);
and U8956 (N_8956,N_8603,N_8749);
xor U8957 (N_8957,N_8674,N_8721);
nand U8958 (N_8958,N_8652,N_8758);
xnor U8959 (N_8959,N_8656,N_8732);
or U8960 (N_8960,N_8781,N_8637);
and U8961 (N_8961,N_8682,N_8718);
and U8962 (N_8962,N_8651,N_8670);
nor U8963 (N_8963,N_8688,N_8673);
nand U8964 (N_8964,N_8678,N_8708);
or U8965 (N_8965,N_8740,N_8656);
xor U8966 (N_8966,N_8751,N_8754);
nor U8967 (N_8967,N_8667,N_8750);
xor U8968 (N_8968,N_8721,N_8680);
xnor U8969 (N_8969,N_8787,N_8663);
nor U8970 (N_8970,N_8721,N_8619);
nor U8971 (N_8971,N_8769,N_8740);
and U8972 (N_8972,N_8758,N_8670);
nand U8973 (N_8973,N_8649,N_8732);
nand U8974 (N_8974,N_8630,N_8736);
nor U8975 (N_8975,N_8776,N_8687);
nor U8976 (N_8976,N_8650,N_8678);
nor U8977 (N_8977,N_8636,N_8617);
nor U8978 (N_8978,N_8662,N_8697);
or U8979 (N_8979,N_8723,N_8793);
nor U8980 (N_8980,N_8646,N_8651);
nor U8981 (N_8981,N_8770,N_8696);
nor U8982 (N_8982,N_8758,N_8641);
or U8983 (N_8983,N_8711,N_8752);
nand U8984 (N_8984,N_8637,N_8638);
or U8985 (N_8985,N_8699,N_8691);
nand U8986 (N_8986,N_8652,N_8717);
or U8987 (N_8987,N_8784,N_8687);
nand U8988 (N_8988,N_8757,N_8767);
xor U8989 (N_8989,N_8638,N_8750);
nand U8990 (N_8990,N_8706,N_8604);
or U8991 (N_8991,N_8784,N_8686);
or U8992 (N_8992,N_8750,N_8799);
nor U8993 (N_8993,N_8612,N_8722);
and U8994 (N_8994,N_8698,N_8692);
nand U8995 (N_8995,N_8797,N_8615);
nand U8996 (N_8996,N_8635,N_8735);
nand U8997 (N_8997,N_8746,N_8770);
nor U8998 (N_8998,N_8798,N_8792);
or U8999 (N_8999,N_8659,N_8625);
nand U9000 (N_9000,N_8897,N_8990);
nand U9001 (N_9001,N_8846,N_8913);
or U9002 (N_9002,N_8865,N_8839);
nor U9003 (N_9003,N_8847,N_8822);
or U9004 (N_9004,N_8817,N_8981);
or U9005 (N_9005,N_8992,N_8952);
and U9006 (N_9006,N_8963,N_8842);
or U9007 (N_9007,N_8920,N_8820);
and U9008 (N_9008,N_8994,N_8856);
nor U9009 (N_9009,N_8840,N_8806);
and U9010 (N_9010,N_8801,N_8943);
nand U9011 (N_9011,N_8815,N_8991);
or U9012 (N_9012,N_8829,N_8821);
nand U9013 (N_9013,N_8802,N_8930);
xor U9014 (N_9014,N_8838,N_8964);
nor U9015 (N_9015,N_8880,N_8888);
or U9016 (N_9016,N_8939,N_8833);
xor U9017 (N_9017,N_8858,N_8905);
or U9018 (N_9018,N_8844,N_8906);
nand U9019 (N_9019,N_8947,N_8974);
or U9020 (N_9020,N_8879,N_8898);
and U9021 (N_9021,N_8861,N_8935);
nand U9022 (N_9022,N_8966,N_8910);
nand U9023 (N_9023,N_8800,N_8851);
or U9024 (N_9024,N_8883,N_8908);
and U9025 (N_9025,N_8911,N_8958);
and U9026 (N_9026,N_8859,N_8954);
nand U9027 (N_9027,N_8933,N_8909);
xor U9028 (N_9028,N_8985,N_8887);
nor U9029 (N_9029,N_8921,N_8946);
nand U9030 (N_9030,N_8987,N_8929);
and U9031 (N_9031,N_8843,N_8890);
and U9032 (N_9032,N_8926,N_8896);
and U9033 (N_9033,N_8928,N_8993);
and U9034 (N_9034,N_8894,N_8891);
nor U9035 (N_9035,N_8996,N_8830);
nor U9036 (N_9036,N_8919,N_8874);
nor U9037 (N_9037,N_8807,N_8810);
nor U9038 (N_9038,N_8892,N_8828);
and U9039 (N_9039,N_8968,N_8824);
and U9040 (N_9040,N_8977,N_8812);
nor U9041 (N_9041,N_8850,N_8826);
nor U9042 (N_9042,N_8982,N_8834);
nand U9043 (N_9043,N_8823,N_8848);
and U9044 (N_9044,N_8827,N_8961);
or U9045 (N_9045,N_8957,N_8857);
or U9046 (N_9046,N_8855,N_8931);
nand U9047 (N_9047,N_8927,N_8860);
nor U9048 (N_9048,N_8932,N_8899);
nand U9049 (N_9049,N_8978,N_8983);
and U9050 (N_9050,N_8944,N_8889);
nand U9051 (N_9051,N_8813,N_8837);
xnor U9052 (N_9052,N_8832,N_8962);
nor U9053 (N_9053,N_8852,N_8818);
xnor U9054 (N_9054,N_8904,N_8971);
nor U9055 (N_9055,N_8975,N_8989);
nor U9056 (N_9056,N_8979,N_8959);
nor U9057 (N_9057,N_8853,N_8901);
nor U9058 (N_9058,N_8809,N_8804);
nor U9059 (N_9059,N_8972,N_8845);
xor U9060 (N_9060,N_8814,N_8862);
nor U9061 (N_9061,N_8941,N_8849);
or U9062 (N_9062,N_8956,N_8882);
nor U9063 (N_9063,N_8980,N_8937);
xor U9064 (N_9064,N_8872,N_8886);
nor U9065 (N_9065,N_8999,N_8923);
or U9066 (N_9066,N_8973,N_8922);
and U9067 (N_9067,N_8903,N_8918);
and U9068 (N_9068,N_8831,N_8976);
or U9069 (N_9069,N_8967,N_8942);
nor U9070 (N_9070,N_8825,N_8819);
or U9071 (N_9071,N_8938,N_8969);
or U9072 (N_9072,N_8816,N_8876);
nor U9073 (N_9073,N_8893,N_8912);
or U9074 (N_9074,N_8936,N_8986);
or U9075 (N_9075,N_8878,N_8866);
nor U9076 (N_9076,N_8948,N_8869);
nand U9077 (N_9077,N_8895,N_8864);
nand U9078 (N_9078,N_8988,N_8873);
or U9079 (N_9079,N_8949,N_8940);
and U9080 (N_9080,N_8871,N_8914);
and U9081 (N_9081,N_8868,N_8997);
nand U9082 (N_9082,N_8877,N_8835);
or U9083 (N_9083,N_8916,N_8955);
or U9084 (N_9084,N_8950,N_8970);
nand U9085 (N_9085,N_8924,N_8960);
nand U9086 (N_9086,N_8915,N_8808);
or U9087 (N_9087,N_8907,N_8925);
or U9088 (N_9088,N_8854,N_8945);
xnor U9089 (N_9089,N_8870,N_8875);
nand U9090 (N_9090,N_8917,N_8867);
and U9091 (N_9091,N_8934,N_8900);
nor U9092 (N_9092,N_8836,N_8984);
nor U9093 (N_9093,N_8881,N_8805);
or U9094 (N_9094,N_8841,N_8884);
and U9095 (N_9095,N_8902,N_8951);
xor U9096 (N_9096,N_8965,N_8803);
nor U9097 (N_9097,N_8995,N_8953);
and U9098 (N_9098,N_8811,N_8863);
or U9099 (N_9099,N_8885,N_8998);
and U9100 (N_9100,N_8811,N_8849);
nor U9101 (N_9101,N_8878,N_8810);
nor U9102 (N_9102,N_8898,N_8864);
nor U9103 (N_9103,N_8915,N_8965);
and U9104 (N_9104,N_8809,N_8805);
nand U9105 (N_9105,N_8901,N_8961);
and U9106 (N_9106,N_8804,N_8892);
nor U9107 (N_9107,N_8924,N_8891);
nor U9108 (N_9108,N_8976,N_8986);
and U9109 (N_9109,N_8913,N_8970);
and U9110 (N_9110,N_8970,N_8918);
nor U9111 (N_9111,N_8909,N_8820);
or U9112 (N_9112,N_8946,N_8857);
nor U9113 (N_9113,N_8917,N_8845);
or U9114 (N_9114,N_8997,N_8938);
xnor U9115 (N_9115,N_8807,N_8834);
or U9116 (N_9116,N_8914,N_8952);
nand U9117 (N_9117,N_8857,N_8958);
nand U9118 (N_9118,N_8886,N_8871);
or U9119 (N_9119,N_8999,N_8874);
or U9120 (N_9120,N_8912,N_8898);
or U9121 (N_9121,N_8845,N_8862);
nand U9122 (N_9122,N_8817,N_8964);
nand U9123 (N_9123,N_8924,N_8966);
or U9124 (N_9124,N_8990,N_8871);
and U9125 (N_9125,N_8934,N_8812);
nand U9126 (N_9126,N_8848,N_8959);
or U9127 (N_9127,N_8949,N_8926);
nand U9128 (N_9128,N_8960,N_8831);
and U9129 (N_9129,N_8865,N_8894);
or U9130 (N_9130,N_8899,N_8905);
and U9131 (N_9131,N_8879,N_8961);
or U9132 (N_9132,N_8911,N_8873);
nand U9133 (N_9133,N_8970,N_8985);
nor U9134 (N_9134,N_8813,N_8820);
and U9135 (N_9135,N_8853,N_8960);
or U9136 (N_9136,N_8984,N_8915);
and U9137 (N_9137,N_8976,N_8848);
xor U9138 (N_9138,N_8915,N_8930);
xnor U9139 (N_9139,N_8866,N_8812);
and U9140 (N_9140,N_8952,N_8904);
and U9141 (N_9141,N_8901,N_8963);
and U9142 (N_9142,N_8819,N_8911);
and U9143 (N_9143,N_8969,N_8863);
nand U9144 (N_9144,N_8859,N_8946);
and U9145 (N_9145,N_8997,N_8857);
nor U9146 (N_9146,N_8911,N_8900);
nor U9147 (N_9147,N_8967,N_8811);
nor U9148 (N_9148,N_8995,N_8866);
xnor U9149 (N_9149,N_8810,N_8895);
and U9150 (N_9150,N_8930,N_8896);
xnor U9151 (N_9151,N_8870,N_8916);
or U9152 (N_9152,N_8904,N_8965);
and U9153 (N_9153,N_8813,N_8869);
xor U9154 (N_9154,N_8966,N_8933);
nor U9155 (N_9155,N_8938,N_8862);
nand U9156 (N_9156,N_8874,N_8912);
and U9157 (N_9157,N_8899,N_8934);
nor U9158 (N_9158,N_8886,N_8829);
or U9159 (N_9159,N_8982,N_8910);
or U9160 (N_9160,N_8892,N_8841);
and U9161 (N_9161,N_8911,N_8907);
nand U9162 (N_9162,N_8805,N_8900);
and U9163 (N_9163,N_8903,N_8813);
nand U9164 (N_9164,N_8853,N_8891);
and U9165 (N_9165,N_8842,N_8881);
xnor U9166 (N_9166,N_8992,N_8928);
or U9167 (N_9167,N_8994,N_8903);
nor U9168 (N_9168,N_8978,N_8864);
nand U9169 (N_9169,N_8889,N_8812);
nand U9170 (N_9170,N_8998,N_8954);
or U9171 (N_9171,N_8806,N_8983);
and U9172 (N_9172,N_8813,N_8892);
or U9173 (N_9173,N_8933,N_8803);
and U9174 (N_9174,N_8991,N_8912);
or U9175 (N_9175,N_8981,N_8967);
xor U9176 (N_9176,N_8896,N_8922);
and U9177 (N_9177,N_8985,N_8881);
or U9178 (N_9178,N_8804,N_8945);
nor U9179 (N_9179,N_8928,N_8913);
nor U9180 (N_9180,N_8975,N_8999);
nor U9181 (N_9181,N_8986,N_8853);
or U9182 (N_9182,N_8947,N_8807);
nand U9183 (N_9183,N_8977,N_8957);
or U9184 (N_9184,N_8812,N_8968);
and U9185 (N_9185,N_8856,N_8892);
xor U9186 (N_9186,N_8938,N_8976);
nor U9187 (N_9187,N_8933,N_8937);
or U9188 (N_9188,N_8836,N_8843);
nand U9189 (N_9189,N_8892,N_8988);
nand U9190 (N_9190,N_8843,N_8917);
nand U9191 (N_9191,N_8828,N_8918);
nor U9192 (N_9192,N_8815,N_8834);
and U9193 (N_9193,N_8938,N_8952);
or U9194 (N_9194,N_8830,N_8932);
nor U9195 (N_9195,N_8821,N_8818);
nor U9196 (N_9196,N_8815,N_8896);
and U9197 (N_9197,N_8949,N_8983);
nor U9198 (N_9198,N_8934,N_8967);
or U9199 (N_9199,N_8846,N_8893);
nor U9200 (N_9200,N_9161,N_9071);
and U9201 (N_9201,N_9081,N_9057);
nand U9202 (N_9202,N_9035,N_9117);
nor U9203 (N_9203,N_9136,N_9198);
nand U9204 (N_9204,N_9024,N_9116);
and U9205 (N_9205,N_9171,N_9154);
nor U9206 (N_9206,N_9138,N_9001);
or U9207 (N_9207,N_9034,N_9056);
or U9208 (N_9208,N_9009,N_9137);
and U9209 (N_9209,N_9011,N_9195);
or U9210 (N_9210,N_9189,N_9048);
nor U9211 (N_9211,N_9096,N_9092);
and U9212 (N_9212,N_9043,N_9039);
nor U9213 (N_9213,N_9126,N_9067);
nand U9214 (N_9214,N_9021,N_9124);
nand U9215 (N_9215,N_9014,N_9055);
or U9216 (N_9216,N_9132,N_9064);
xor U9217 (N_9217,N_9032,N_9181);
or U9218 (N_9218,N_9058,N_9089);
nand U9219 (N_9219,N_9157,N_9075);
and U9220 (N_9220,N_9162,N_9063);
or U9221 (N_9221,N_9179,N_9106);
nor U9222 (N_9222,N_9140,N_9040);
or U9223 (N_9223,N_9004,N_9142);
and U9224 (N_9224,N_9192,N_9196);
xor U9225 (N_9225,N_9012,N_9165);
or U9226 (N_9226,N_9033,N_9079);
and U9227 (N_9227,N_9070,N_9152);
or U9228 (N_9228,N_9003,N_9194);
or U9229 (N_9229,N_9010,N_9186);
and U9230 (N_9230,N_9098,N_9121);
and U9231 (N_9231,N_9135,N_9066);
nand U9232 (N_9232,N_9190,N_9150);
and U9233 (N_9233,N_9041,N_9019);
xnor U9234 (N_9234,N_9065,N_9008);
and U9235 (N_9235,N_9013,N_9061);
and U9236 (N_9236,N_9097,N_9146);
and U9237 (N_9237,N_9185,N_9080);
nand U9238 (N_9238,N_9184,N_9174);
xnor U9239 (N_9239,N_9122,N_9053);
and U9240 (N_9240,N_9006,N_9088);
nor U9241 (N_9241,N_9119,N_9112);
or U9242 (N_9242,N_9148,N_9193);
and U9243 (N_9243,N_9158,N_9160);
and U9244 (N_9244,N_9046,N_9159);
nand U9245 (N_9245,N_9077,N_9020);
or U9246 (N_9246,N_9128,N_9005);
or U9247 (N_9247,N_9129,N_9100);
nand U9248 (N_9248,N_9018,N_9076);
or U9249 (N_9249,N_9147,N_9108);
nand U9250 (N_9250,N_9094,N_9101);
nand U9251 (N_9251,N_9180,N_9175);
nand U9252 (N_9252,N_9115,N_9107);
or U9253 (N_9253,N_9172,N_9037);
nand U9254 (N_9254,N_9141,N_9191);
and U9255 (N_9255,N_9168,N_9016);
or U9256 (N_9256,N_9052,N_9105);
nand U9257 (N_9257,N_9002,N_9095);
nor U9258 (N_9258,N_9111,N_9143);
nor U9259 (N_9259,N_9023,N_9173);
nor U9260 (N_9260,N_9027,N_9166);
nand U9261 (N_9261,N_9029,N_9155);
and U9262 (N_9262,N_9176,N_9178);
nand U9263 (N_9263,N_9127,N_9050);
nor U9264 (N_9264,N_9025,N_9078);
nor U9265 (N_9265,N_9118,N_9091);
and U9266 (N_9266,N_9099,N_9133);
xnor U9267 (N_9267,N_9169,N_9139);
and U9268 (N_9268,N_9036,N_9028);
or U9269 (N_9269,N_9163,N_9054);
or U9270 (N_9270,N_9060,N_9059);
and U9271 (N_9271,N_9104,N_9197);
nor U9272 (N_9272,N_9110,N_9015);
and U9273 (N_9273,N_9145,N_9167);
and U9274 (N_9274,N_9051,N_9102);
nand U9275 (N_9275,N_9022,N_9085);
nand U9276 (N_9276,N_9030,N_9183);
and U9277 (N_9277,N_9082,N_9130);
nor U9278 (N_9278,N_9087,N_9187);
xor U9279 (N_9279,N_9045,N_9114);
nand U9280 (N_9280,N_9199,N_9090);
nor U9281 (N_9281,N_9093,N_9083);
nand U9282 (N_9282,N_9042,N_9017);
xnor U9283 (N_9283,N_9103,N_9123);
nor U9284 (N_9284,N_9153,N_9188);
and U9285 (N_9285,N_9007,N_9182);
nor U9286 (N_9286,N_9156,N_9177);
nor U9287 (N_9287,N_9068,N_9072);
or U9288 (N_9288,N_9038,N_9164);
and U9289 (N_9289,N_9049,N_9000);
or U9290 (N_9290,N_9062,N_9151);
nor U9291 (N_9291,N_9120,N_9134);
or U9292 (N_9292,N_9144,N_9044);
nand U9293 (N_9293,N_9026,N_9113);
nor U9294 (N_9294,N_9131,N_9073);
xnor U9295 (N_9295,N_9125,N_9031);
nor U9296 (N_9296,N_9170,N_9149);
or U9297 (N_9297,N_9086,N_9047);
and U9298 (N_9298,N_9109,N_9069);
and U9299 (N_9299,N_9074,N_9084);
nand U9300 (N_9300,N_9048,N_9149);
nor U9301 (N_9301,N_9075,N_9091);
and U9302 (N_9302,N_9032,N_9028);
nand U9303 (N_9303,N_9083,N_9018);
or U9304 (N_9304,N_9193,N_9042);
and U9305 (N_9305,N_9000,N_9047);
nor U9306 (N_9306,N_9176,N_9198);
xor U9307 (N_9307,N_9011,N_9135);
or U9308 (N_9308,N_9115,N_9080);
nor U9309 (N_9309,N_9114,N_9157);
nand U9310 (N_9310,N_9062,N_9119);
and U9311 (N_9311,N_9125,N_9150);
and U9312 (N_9312,N_9003,N_9045);
or U9313 (N_9313,N_9161,N_9026);
and U9314 (N_9314,N_9097,N_9137);
nand U9315 (N_9315,N_9147,N_9185);
nor U9316 (N_9316,N_9194,N_9074);
or U9317 (N_9317,N_9192,N_9095);
and U9318 (N_9318,N_9073,N_9024);
or U9319 (N_9319,N_9111,N_9087);
xnor U9320 (N_9320,N_9195,N_9050);
xor U9321 (N_9321,N_9093,N_9124);
and U9322 (N_9322,N_9023,N_9075);
xor U9323 (N_9323,N_9110,N_9072);
nor U9324 (N_9324,N_9063,N_9004);
nand U9325 (N_9325,N_9033,N_9164);
nor U9326 (N_9326,N_9083,N_9070);
or U9327 (N_9327,N_9199,N_9113);
nand U9328 (N_9328,N_9143,N_9073);
or U9329 (N_9329,N_9025,N_9067);
nand U9330 (N_9330,N_9055,N_9084);
xnor U9331 (N_9331,N_9098,N_9167);
nor U9332 (N_9332,N_9182,N_9121);
and U9333 (N_9333,N_9116,N_9030);
and U9334 (N_9334,N_9121,N_9141);
nor U9335 (N_9335,N_9035,N_9096);
or U9336 (N_9336,N_9131,N_9011);
nand U9337 (N_9337,N_9041,N_9036);
xnor U9338 (N_9338,N_9120,N_9086);
or U9339 (N_9339,N_9086,N_9064);
nor U9340 (N_9340,N_9043,N_9194);
nand U9341 (N_9341,N_9165,N_9027);
nand U9342 (N_9342,N_9184,N_9017);
or U9343 (N_9343,N_9164,N_9149);
nand U9344 (N_9344,N_9161,N_9023);
nand U9345 (N_9345,N_9072,N_9038);
nand U9346 (N_9346,N_9034,N_9068);
or U9347 (N_9347,N_9151,N_9198);
xor U9348 (N_9348,N_9007,N_9153);
nand U9349 (N_9349,N_9194,N_9120);
xnor U9350 (N_9350,N_9199,N_9052);
nor U9351 (N_9351,N_9123,N_9065);
or U9352 (N_9352,N_9170,N_9172);
nand U9353 (N_9353,N_9064,N_9190);
or U9354 (N_9354,N_9183,N_9059);
xnor U9355 (N_9355,N_9144,N_9081);
nor U9356 (N_9356,N_9141,N_9041);
nor U9357 (N_9357,N_9106,N_9158);
and U9358 (N_9358,N_9008,N_9182);
nand U9359 (N_9359,N_9183,N_9026);
xnor U9360 (N_9360,N_9000,N_9195);
nand U9361 (N_9361,N_9025,N_9148);
or U9362 (N_9362,N_9086,N_9016);
and U9363 (N_9363,N_9167,N_9038);
or U9364 (N_9364,N_9157,N_9125);
and U9365 (N_9365,N_9138,N_9017);
or U9366 (N_9366,N_9114,N_9137);
nor U9367 (N_9367,N_9005,N_9008);
nand U9368 (N_9368,N_9081,N_9186);
and U9369 (N_9369,N_9106,N_9071);
nand U9370 (N_9370,N_9164,N_9185);
nor U9371 (N_9371,N_9089,N_9119);
and U9372 (N_9372,N_9067,N_9008);
nand U9373 (N_9373,N_9047,N_9168);
nand U9374 (N_9374,N_9039,N_9014);
nor U9375 (N_9375,N_9144,N_9152);
xnor U9376 (N_9376,N_9167,N_9003);
nand U9377 (N_9377,N_9134,N_9127);
or U9378 (N_9378,N_9180,N_9082);
and U9379 (N_9379,N_9067,N_9114);
nand U9380 (N_9380,N_9024,N_9196);
and U9381 (N_9381,N_9006,N_9184);
nand U9382 (N_9382,N_9155,N_9001);
or U9383 (N_9383,N_9116,N_9106);
and U9384 (N_9384,N_9181,N_9021);
xor U9385 (N_9385,N_9022,N_9009);
or U9386 (N_9386,N_9182,N_9111);
or U9387 (N_9387,N_9073,N_9188);
xnor U9388 (N_9388,N_9185,N_9136);
nand U9389 (N_9389,N_9176,N_9002);
or U9390 (N_9390,N_9198,N_9034);
nor U9391 (N_9391,N_9148,N_9034);
and U9392 (N_9392,N_9086,N_9121);
and U9393 (N_9393,N_9040,N_9131);
or U9394 (N_9394,N_9147,N_9072);
and U9395 (N_9395,N_9038,N_9035);
nand U9396 (N_9396,N_9021,N_9178);
and U9397 (N_9397,N_9098,N_9172);
and U9398 (N_9398,N_9180,N_9102);
nor U9399 (N_9399,N_9098,N_9081);
or U9400 (N_9400,N_9259,N_9220);
or U9401 (N_9401,N_9323,N_9237);
or U9402 (N_9402,N_9389,N_9284);
nand U9403 (N_9403,N_9383,N_9260);
and U9404 (N_9404,N_9262,N_9392);
or U9405 (N_9405,N_9363,N_9351);
nand U9406 (N_9406,N_9293,N_9341);
nand U9407 (N_9407,N_9344,N_9331);
xnor U9408 (N_9408,N_9391,N_9345);
nand U9409 (N_9409,N_9305,N_9209);
and U9410 (N_9410,N_9210,N_9332);
nand U9411 (N_9411,N_9206,N_9273);
nand U9412 (N_9412,N_9352,N_9204);
nor U9413 (N_9413,N_9384,N_9368);
or U9414 (N_9414,N_9295,N_9288);
or U9415 (N_9415,N_9286,N_9285);
xor U9416 (N_9416,N_9283,N_9378);
nor U9417 (N_9417,N_9361,N_9251);
nand U9418 (N_9418,N_9207,N_9304);
or U9419 (N_9419,N_9313,N_9329);
and U9420 (N_9420,N_9356,N_9269);
nand U9421 (N_9421,N_9264,N_9231);
nand U9422 (N_9422,N_9221,N_9303);
or U9423 (N_9423,N_9245,N_9333);
and U9424 (N_9424,N_9244,N_9297);
and U9425 (N_9425,N_9203,N_9340);
or U9426 (N_9426,N_9364,N_9240);
nand U9427 (N_9427,N_9353,N_9228);
nor U9428 (N_9428,N_9395,N_9242);
nand U9429 (N_9429,N_9214,N_9372);
nand U9430 (N_9430,N_9370,N_9230);
nor U9431 (N_9431,N_9385,N_9294);
and U9432 (N_9432,N_9249,N_9274);
nand U9433 (N_9433,N_9390,N_9238);
and U9434 (N_9434,N_9365,N_9299);
and U9435 (N_9435,N_9387,N_9217);
or U9436 (N_9436,N_9307,N_9239);
nor U9437 (N_9437,N_9316,N_9394);
and U9438 (N_9438,N_9263,N_9362);
nand U9439 (N_9439,N_9243,N_9218);
or U9440 (N_9440,N_9257,N_9398);
or U9441 (N_9441,N_9290,N_9334);
nor U9442 (N_9442,N_9270,N_9219);
nor U9443 (N_9443,N_9298,N_9376);
nor U9444 (N_9444,N_9254,N_9236);
or U9445 (N_9445,N_9234,N_9222);
or U9446 (N_9446,N_9275,N_9324);
xor U9447 (N_9447,N_9250,N_9346);
nor U9448 (N_9448,N_9322,N_9278);
and U9449 (N_9449,N_9227,N_9213);
and U9450 (N_9450,N_9287,N_9399);
nand U9451 (N_9451,N_9267,N_9319);
or U9452 (N_9452,N_9380,N_9225);
nor U9453 (N_9453,N_9276,N_9311);
nand U9454 (N_9454,N_9235,N_9349);
or U9455 (N_9455,N_9241,N_9347);
and U9456 (N_9456,N_9261,N_9358);
xnor U9457 (N_9457,N_9318,N_9296);
nor U9458 (N_9458,N_9335,N_9246);
nand U9459 (N_9459,N_9374,N_9224);
or U9460 (N_9460,N_9337,N_9382);
nor U9461 (N_9461,N_9381,N_9310);
nand U9462 (N_9462,N_9336,N_9301);
nand U9463 (N_9463,N_9312,N_9367);
and U9464 (N_9464,N_9354,N_9253);
nor U9465 (N_9465,N_9359,N_9282);
nand U9466 (N_9466,N_9377,N_9388);
nand U9467 (N_9467,N_9309,N_9371);
nand U9468 (N_9468,N_9281,N_9386);
nand U9469 (N_9469,N_9321,N_9338);
nor U9470 (N_9470,N_9397,N_9306);
nor U9471 (N_9471,N_9226,N_9320);
nand U9472 (N_9472,N_9326,N_9317);
or U9473 (N_9473,N_9212,N_9202);
nand U9474 (N_9474,N_9208,N_9265);
or U9475 (N_9475,N_9205,N_9255);
nor U9476 (N_9476,N_9355,N_9280);
and U9477 (N_9477,N_9369,N_9302);
or U9478 (N_9478,N_9258,N_9211);
nand U9479 (N_9479,N_9271,N_9216);
nor U9480 (N_9480,N_9291,N_9232);
and U9481 (N_9481,N_9252,N_9200);
and U9482 (N_9482,N_9229,N_9289);
and U9483 (N_9483,N_9373,N_9396);
or U9484 (N_9484,N_9330,N_9327);
nand U9485 (N_9485,N_9342,N_9256);
and U9486 (N_9486,N_9233,N_9308);
xnor U9487 (N_9487,N_9300,N_9325);
and U9488 (N_9488,N_9379,N_9277);
nand U9489 (N_9489,N_9201,N_9266);
nor U9490 (N_9490,N_9215,N_9328);
nand U9491 (N_9491,N_9247,N_9350);
nor U9492 (N_9492,N_9366,N_9375);
and U9493 (N_9493,N_9360,N_9314);
xnor U9494 (N_9494,N_9393,N_9279);
nand U9495 (N_9495,N_9223,N_9268);
and U9496 (N_9496,N_9343,N_9315);
nand U9497 (N_9497,N_9292,N_9248);
or U9498 (N_9498,N_9348,N_9272);
xnor U9499 (N_9499,N_9339,N_9357);
xnor U9500 (N_9500,N_9310,N_9252);
xnor U9501 (N_9501,N_9299,N_9393);
or U9502 (N_9502,N_9256,N_9243);
or U9503 (N_9503,N_9295,N_9346);
or U9504 (N_9504,N_9365,N_9379);
nor U9505 (N_9505,N_9320,N_9207);
nand U9506 (N_9506,N_9347,N_9319);
or U9507 (N_9507,N_9289,N_9220);
nand U9508 (N_9508,N_9361,N_9281);
nand U9509 (N_9509,N_9262,N_9245);
nor U9510 (N_9510,N_9311,N_9218);
nor U9511 (N_9511,N_9328,N_9350);
nor U9512 (N_9512,N_9386,N_9208);
and U9513 (N_9513,N_9294,N_9310);
nand U9514 (N_9514,N_9322,N_9207);
and U9515 (N_9515,N_9223,N_9309);
nand U9516 (N_9516,N_9348,N_9286);
and U9517 (N_9517,N_9227,N_9329);
nor U9518 (N_9518,N_9303,N_9326);
nand U9519 (N_9519,N_9231,N_9268);
nor U9520 (N_9520,N_9210,N_9242);
or U9521 (N_9521,N_9306,N_9241);
xor U9522 (N_9522,N_9351,N_9275);
or U9523 (N_9523,N_9346,N_9366);
nand U9524 (N_9524,N_9288,N_9238);
nor U9525 (N_9525,N_9249,N_9303);
nand U9526 (N_9526,N_9342,N_9279);
nor U9527 (N_9527,N_9387,N_9285);
or U9528 (N_9528,N_9385,N_9248);
and U9529 (N_9529,N_9249,N_9380);
and U9530 (N_9530,N_9393,N_9309);
xnor U9531 (N_9531,N_9290,N_9215);
nor U9532 (N_9532,N_9343,N_9325);
and U9533 (N_9533,N_9386,N_9384);
nor U9534 (N_9534,N_9329,N_9226);
nor U9535 (N_9535,N_9326,N_9358);
and U9536 (N_9536,N_9343,N_9395);
nand U9537 (N_9537,N_9232,N_9264);
and U9538 (N_9538,N_9228,N_9390);
and U9539 (N_9539,N_9235,N_9287);
xor U9540 (N_9540,N_9373,N_9310);
and U9541 (N_9541,N_9279,N_9221);
nand U9542 (N_9542,N_9323,N_9286);
nand U9543 (N_9543,N_9398,N_9247);
and U9544 (N_9544,N_9303,N_9293);
nor U9545 (N_9545,N_9367,N_9351);
nand U9546 (N_9546,N_9388,N_9338);
nand U9547 (N_9547,N_9331,N_9359);
and U9548 (N_9548,N_9311,N_9220);
and U9549 (N_9549,N_9227,N_9287);
nand U9550 (N_9550,N_9343,N_9210);
or U9551 (N_9551,N_9302,N_9394);
nand U9552 (N_9552,N_9225,N_9279);
and U9553 (N_9553,N_9381,N_9274);
nor U9554 (N_9554,N_9388,N_9389);
or U9555 (N_9555,N_9277,N_9373);
xor U9556 (N_9556,N_9326,N_9300);
nand U9557 (N_9557,N_9228,N_9227);
nand U9558 (N_9558,N_9364,N_9307);
or U9559 (N_9559,N_9304,N_9399);
or U9560 (N_9560,N_9293,N_9345);
or U9561 (N_9561,N_9370,N_9354);
nand U9562 (N_9562,N_9232,N_9299);
nand U9563 (N_9563,N_9228,N_9358);
or U9564 (N_9564,N_9245,N_9233);
or U9565 (N_9565,N_9284,N_9265);
and U9566 (N_9566,N_9248,N_9202);
nor U9567 (N_9567,N_9372,N_9308);
or U9568 (N_9568,N_9291,N_9337);
nor U9569 (N_9569,N_9339,N_9280);
or U9570 (N_9570,N_9381,N_9356);
and U9571 (N_9571,N_9347,N_9320);
or U9572 (N_9572,N_9263,N_9307);
nand U9573 (N_9573,N_9346,N_9277);
nand U9574 (N_9574,N_9341,N_9392);
xnor U9575 (N_9575,N_9296,N_9389);
nand U9576 (N_9576,N_9206,N_9307);
and U9577 (N_9577,N_9206,N_9336);
nor U9578 (N_9578,N_9259,N_9290);
xor U9579 (N_9579,N_9228,N_9357);
or U9580 (N_9580,N_9399,N_9259);
or U9581 (N_9581,N_9349,N_9262);
nand U9582 (N_9582,N_9326,N_9221);
and U9583 (N_9583,N_9255,N_9320);
or U9584 (N_9584,N_9329,N_9338);
or U9585 (N_9585,N_9291,N_9394);
nand U9586 (N_9586,N_9296,N_9254);
and U9587 (N_9587,N_9264,N_9394);
nand U9588 (N_9588,N_9284,N_9244);
and U9589 (N_9589,N_9232,N_9318);
xor U9590 (N_9590,N_9208,N_9251);
and U9591 (N_9591,N_9239,N_9394);
nand U9592 (N_9592,N_9329,N_9237);
and U9593 (N_9593,N_9314,N_9227);
nor U9594 (N_9594,N_9276,N_9344);
nand U9595 (N_9595,N_9293,N_9231);
xor U9596 (N_9596,N_9331,N_9219);
nor U9597 (N_9597,N_9260,N_9226);
and U9598 (N_9598,N_9330,N_9292);
or U9599 (N_9599,N_9255,N_9230);
and U9600 (N_9600,N_9550,N_9404);
nand U9601 (N_9601,N_9568,N_9402);
nand U9602 (N_9602,N_9436,N_9499);
and U9603 (N_9603,N_9566,N_9470);
nor U9604 (N_9604,N_9555,N_9488);
or U9605 (N_9605,N_9526,N_9539);
nand U9606 (N_9606,N_9595,N_9548);
and U9607 (N_9607,N_9569,N_9554);
nor U9608 (N_9608,N_9545,N_9508);
xnor U9609 (N_9609,N_9558,N_9557);
nor U9610 (N_9610,N_9537,N_9471);
xor U9611 (N_9611,N_9407,N_9424);
and U9612 (N_9612,N_9408,N_9547);
and U9613 (N_9613,N_9438,N_9431);
and U9614 (N_9614,N_9523,N_9587);
or U9615 (N_9615,N_9417,N_9449);
nor U9616 (N_9616,N_9597,N_9519);
nand U9617 (N_9617,N_9511,N_9462);
or U9618 (N_9618,N_9446,N_9452);
nor U9619 (N_9619,N_9529,N_9453);
nor U9620 (N_9620,N_9428,N_9559);
nand U9621 (N_9621,N_9564,N_9457);
xor U9622 (N_9622,N_9484,N_9433);
nand U9623 (N_9623,N_9472,N_9426);
and U9624 (N_9624,N_9464,N_9582);
nand U9625 (N_9625,N_9584,N_9429);
and U9626 (N_9626,N_9580,N_9401);
nor U9627 (N_9627,N_9542,N_9549);
nand U9628 (N_9628,N_9482,N_9466);
nand U9629 (N_9629,N_9562,N_9563);
xor U9630 (N_9630,N_9496,N_9535);
xor U9631 (N_9631,N_9487,N_9593);
or U9632 (N_9632,N_9536,N_9413);
nor U9633 (N_9633,N_9430,N_9509);
or U9634 (N_9634,N_9543,N_9479);
or U9635 (N_9635,N_9448,N_9571);
nand U9636 (N_9636,N_9515,N_9418);
or U9637 (N_9637,N_9522,N_9551);
nor U9638 (N_9638,N_9492,N_9406);
nor U9639 (N_9639,N_9596,N_9503);
nand U9640 (N_9640,N_9437,N_9514);
and U9641 (N_9641,N_9530,N_9560);
or U9642 (N_9642,N_9588,N_9507);
or U9643 (N_9643,N_9546,N_9544);
or U9644 (N_9644,N_9454,N_9458);
nand U9645 (N_9645,N_9456,N_9502);
nand U9646 (N_9646,N_9411,N_9415);
nor U9647 (N_9647,N_9441,N_9494);
or U9648 (N_9648,N_9516,N_9495);
and U9649 (N_9649,N_9463,N_9591);
nor U9650 (N_9650,N_9517,N_9577);
nor U9651 (N_9651,N_9491,N_9512);
and U9652 (N_9652,N_9592,N_9541);
xor U9653 (N_9653,N_9581,N_9423);
and U9654 (N_9654,N_9506,N_9510);
or U9655 (N_9655,N_9497,N_9403);
or U9656 (N_9656,N_9578,N_9478);
or U9657 (N_9657,N_9585,N_9435);
nand U9658 (N_9658,N_9434,N_9533);
xor U9659 (N_9659,N_9443,N_9410);
or U9660 (N_9660,N_9493,N_9440);
nor U9661 (N_9661,N_9476,N_9474);
nand U9662 (N_9662,N_9486,N_9467);
and U9663 (N_9663,N_9570,N_9485);
xor U9664 (N_9664,N_9459,N_9576);
or U9665 (N_9665,N_9594,N_9501);
nand U9666 (N_9666,N_9527,N_9412);
nand U9667 (N_9667,N_9468,N_9445);
nand U9668 (N_9668,N_9481,N_9531);
and U9669 (N_9669,N_9575,N_9534);
or U9670 (N_9670,N_9590,N_9556);
and U9671 (N_9671,N_9469,N_9419);
or U9672 (N_9672,N_9572,N_9565);
or U9673 (N_9673,N_9409,N_9477);
nand U9674 (N_9674,N_9420,N_9505);
nand U9675 (N_9675,N_9483,N_9432);
or U9676 (N_9676,N_9528,N_9520);
and U9677 (N_9677,N_9567,N_9422);
nand U9678 (N_9678,N_9425,N_9538);
nor U9679 (N_9679,N_9405,N_9427);
nand U9680 (N_9680,N_9447,N_9518);
nand U9681 (N_9681,N_9461,N_9421);
and U9682 (N_9682,N_9540,N_9573);
xor U9683 (N_9683,N_9586,N_9598);
nor U9684 (N_9684,N_9442,N_9451);
nor U9685 (N_9685,N_9589,N_9473);
nand U9686 (N_9686,N_9455,N_9553);
nand U9687 (N_9687,N_9500,N_9552);
nand U9688 (N_9688,N_9532,N_9498);
and U9689 (N_9689,N_9599,N_9489);
or U9690 (N_9690,N_9416,N_9524);
or U9691 (N_9691,N_9579,N_9521);
or U9692 (N_9692,N_9460,N_9439);
or U9693 (N_9693,N_9574,N_9525);
nor U9694 (N_9694,N_9414,N_9400);
or U9695 (N_9695,N_9450,N_9444);
or U9696 (N_9696,N_9561,N_9513);
or U9697 (N_9697,N_9465,N_9504);
nand U9698 (N_9698,N_9480,N_9583);
and U9699 (N_9699,N_9475,N_9490);
or U9700 (N_9700,N_9584,N_9587);
or U9701 (N_9701,N_9484,N_9537);
and U9702 (N_9702,N_9485,N_9574);
nor U9703 (N_9703,N_9501,N_9406);
or U9704 (N_9704,N_9438,N_9516);
nor U9705 (N_9705,N_9528,N_9534);
nor U9706 (N_9706,N_9589,N_9499);
or U9707 (N_9707,N_9442,N_9573);
or U9708 (N_9708,N_9450,N_9401);
nand U9709 (N_9709,N_9554,N_9489);
nor U9710 (N_9710,N_9546,N_9525);
or U9711 (N_9711,N_9479,N_9491);
xnor U9712 (N_9712,N_9546,N_9548);
nand U9713 (N_9713,N_9414,N_9490);
or U9714 (N_9714,N_9543,N_9596);
and U9715 (N_9715,N_9493,N_9556);
or U9716 (N_9716,N_9536,N_9537);
nand U9717 (N_9717,N_9491,N_9541);
nand U9718 (N_9718,N_9548,N_9538);
or U9719 (N_9719,N_9518,N_9506);
and U9720 (N_9720,N_9517,N_9525);
or U9721 (N_9721,N_9463,N_9509);
or U9722 (N_9722,N_9583,N_9458);
xnor U9723 (N_9723,N_9569,N_9431);
and U9724 (N_9724,N_9438,N_9463);
and U9725 (N_9725,N_9422,N_9575);
nand U9726 (N_9726,N_9506,N_9466);
and U9727 (N_9727,N_9535,N_9591);
xor U9728 (N_9728,N_9477,N_9446);
nand U9729 (N_9729,N_9525,N_9551);
nand U9730 (N_9730,N_9432,N_9507);
and U9731 (N_9731,N_9521,N_9599);
or U9732 (N_9732,N_9419,N_9411);
nand U9733 (N_9733,N_9548,N_9521);
nor U9734 (N_9734,N_9429,N_9594);
xnor U9735 (N_9735,N_9538,N_9596);
and U9736 (N_9736,N_9496,N_9552);
or U9737 (N_9737,N_9525,N_9448);
nor U9738 (N_9738,N_9578,N_9420);
and U9739 (N_9739,N_9435,N_9423);
or U9740 (N_9740,N_9523,N_9569);
nor U9741 (N_9741,N_9452,N_9572);
xor U9742 (N_9742,N_9507,N_9594);
nor U9743 (N_9743,N_9489,N_9485);
and U9744 (N_9744,N_9416,N_9548);
and U9745 (N_9745,N_9501,N_9506);
or U9746 (N_9746,N_9469,N_9555);
or U9747 (N_9747,N_9425,N_9524);
xnor U9748 (N_9748,N_9534,N_9465);
nor U9749 (N_9749,N_9468,N_9565);
and U9750 (N_9750,N_9438,N_9491);
nand U9751 (N_9751,N_9451,N_9552);
and U9752 (N_9752,N_9596,N_9445);
and U9753 (N_9753,N_9474,N_9593);
nand U9754 (N_9754,N_9432,N_9551);
and U9755 (N_9755,N_9468,N_9472);
nor U9756 (N_9756,N_9578,N_9540);
or U9757 (N_9757,N_9556,N_9480);
or U9758 (N_9758,N_9565,N_9457);
or U9759 (N_9759,N_9580,N_9407);
nor U9760 (N_9760,N_9540,N_9569);
or U9761 (N_9761,N_9408,N_9599);
or U9762 (N_9762,N_9461,N_9445);
and U9763 (N_9763,N_9489,N_9570);
xor U9764 (N_9764,N_9492,N_9468);
nor U9765 (N_9765,N_9572,N_9477);
nor U9766 (N_9766,N_9592,N_9510);
nor U9767 (N_9767,N_9503,N_9411);
and U9768 (N_9768,N_9468,N_9524);
and U9769 (N_9769,N_9447,N_9527);
nor U9770 (N_9770,N_9475,N_9521);
or U9771 (N_9771,N_9522,N_9402);
nor U9772 (N_9772,N_9562,N_9432);
nor U9773 (N_9773,N_9480,N_9432);
or U9774 (N_9774,N_9544,N_9499);
and U9775 (N_9775,N_9432,N_9409);
and U9776 (N_9776,N_9589,N_9498);
and U9777 (N_9777,N_9530,N_9552);
nor U9778 (N_9778,N_9588,N_9514);
nand U9779 (N_9779,N_9455,N_9545);
nand U9780 (N_9780,N_9468,N_9576);
nor U9781 (N_9781,N_9551,N_9508);
and U9782 (N_9782,N_9455,N_9565);
and U9783 (N_9783,N_9491,N_9599);
and U9784 (N_9784,N_9551,N_9529);
and U9785 (N_9785,N_9527,N_9431);
and U9786 (N_9786,N_9498,N_9533);
nor U9787 (N_9787,N_9561,N_9472);
nor U9788 (N_9788,N_9403,N_9591);
xnor U9789 (N_9789,N_9490,N_9433);
or U9790 (N_9790,N_9404,N_9415);
nor U9791 (N_9791,N_9582,N_9549);
or U9792 (N_9792,N_9425,N_9445);
nand U9793 (N_9793,N_9489,N_9497);
nor U9794 (N_9794,N_9436,N_9437);
nor U9795 (N_9795,N_9491,N_9418);
nor U9796 (N_9796,N_9513,N_9448);
or U9797 (N_9797,N_9561,N_9459);
and U9798 (N_9798,N_9431,N_9418);
and U9799 (N_9799,N_9522,N_9429);
or U9800 (N_9800,N_9684,N_9717);
or U9801 (N_9801,N_9672,N_9693);
nand U9802 (N_9802,N_9749,N_9644);
xnor U9803 (N_9803,N_9762,N_9638);
or U9804 (N_9804,N_9615,N_9635);
nor U9805 (N_9805,N_9776,N_9695);
nor U9806 (N_9806,N_9738,N_9649);
nor U9807 (N_9807,N_9793,N_9788);
or U9808 (N_9808,N_9613,N_9732);
or U9809 (N_9809,N_9711,N_9702);
nand U9810 (N_9810,N_9643,N_9608);
or U9811 (N_9811,N_9761,N_9757);
or U9812 (N_9812,N_9659,N_9634);
or U9813 (N_9813,N_9715,N_9718);
or U9814 (N_9814,N_9748,N_9754);
nand U9815 (N_9815,N_9646,N_9650);
nand U9816 (N_9816,N_9614,N_9605);
and U9817 (N_9817,N_9791,N_9642);
nor U9818 (N_9818,N_9792,N_9799);
and U9819 (N_9819,N_9699,N_9733);
and U9820 (N_9820,N_9758,N_9723);
nand U9821 (N_9821,N_9679,N_9780);
nand U9822 (N_9822,N_9728,N_9618);
nand U9823 (N_9823,N_9633,N_9662);
and U9824 (N_9824,N_9736,N_9674);
or U9825 (N_9825,N_9645,N_9683);
nor U9826 (N_9826,N_9706,N_9726);
and U9827 (N_9827,N_9669,N_9685);
nor U9828 (N_9828,N_9787,N_9677);
nor U9829 (N_9829,N_9774,N_9730);
or U9830 (N_9830,N_9713,N_9790);
or U9831 (N_9831,N_9766,N_9627);
or U9832 (N_9832,N_9745,N_9640);
nor U9833 (N_9833,N_9625,N_9668);
or U9834 (N_9834,N_9676,N_9783);
or U9835 (N_9835,N_9789,N_9781);
xor U9836 (N_9836,N_9734,N_9630);
nand U9837 (N_9837,N_9691,N_9637);
nand U9838 (N_9838,N_9655,N_9652);
nand U9839 (N_9839,N_9688,N_9663);
nor U9840 (N_9840,N_9664,N_9768);
nor U9841 (N_9841,N_9641,N_9671);
nand U9842 (N_9842,N_9798,N_9705);
nor U9843 (N_9843,N_9721,N_9657);
nor U9844 (N_9844,N_9670,N_9740);
and U9845 (N_9845,N_9786,N_9604);
nand U9846 (N_9846,N_9620,N_9704);
or U9847 (N_9847,N_9744,N_9617);
or U9848 (N_9848,N_9743,N_9739);
nand U9849 (N_9849,N_9722,N_9742);
and U9850 (N_9850,N_9779,N_9607);
and U9851 (N_9851,N_9796,N_9612);
nor U9852 (N_9852,N_9770,N_9753);
nor U9853 (N_9853,N_9755,N_9785);
xor U9854 (N_9854,N_9665,N_9678);
or U9855 (N_9855,N_9716,N_9775);
and U9856 (N_9856,N_9603,N_9623);
nand U9857 (N_9857,N_9741,N_9621);
or U9858 (N_9858,N_9794,N_9756);
nor U9859 (N_9859,N_9606,N_9700);
nor U9860 (N_9860,N_9760,N_9656);
xnor U9861 (N_9861,N_9619,N_9720);
or U9862 (N_9862,N_9658,N_9639);
or U9863 (N_9863,N_9600,N_9751);
nand U9864 (N_9864,N_9767,N_9759);
nor U9865 (N_9865,N_9752,N_9769);
nand U9866 (N_9866,N_9661,N_9631);
or U9867 (N_9867,N_9681,N_9710);
and U9868 (N_9868,N_9727,N_9647);
or U9869 (N_9869,N_9601,N_9777);
and U9870 (N_9870,N_9765,N_9689);
and U9871 (N_9871,N_9686,N_9773);
or U9872 (N_9872,N_9632,N_9750);
or U9873 (N_9873,N_9666,N_9714);
and U9874 (N_9874,N_9707,N_9636);
nor U9875 (N_9875,N_9763,N_9622);
and U9876 (N_9876,N_9667,N_9737);
or U9877 (N_9877,N_9602,N_9690);
or U9878 (N_9878,N_9651,N_9682);
nand U9879 (N_9879,N_9611,N_9719);
nor U9880 (N_9880,N_9696,N_9697);
or U9881 (N_9881,N_9747,N_9675);
and U9882 (N_9882,N_9660,N_9729);
or U9883 (N_9883,N_9708,N_9687);
or U9884 (N_9884,N_9694,N_9784);
or U9885 (N_9885,N_9654,N_9624);
nand U9886 (N_9886,N_9709,N_9782);
nand U9887 (N_9887,N_9648,N_9609);
xnor U9888 (N_9888,N_9692,N_9698);
and U9889 (N_9889,N_9712,N_9701);
nand U9890 (N_9890,N_9629,N_9771);
nor U9891 (N_9891,N_9724,N_9653);
nand U9892 (N_9892,N_9610,N_9703);
and U9893 (N_9893,N_9735,N_9626);
or U9894 (N_9894,N_9725,N_9778);
and U9895 (N_9895,N_9795,N_9731);
nor U9896 (N_9896,N_9673,N_9764);
or U9897 (N_9897,N_9680,N_9746);
or U9898 (N_9898,N_9772,N_9797);
or U9899 (N_9899,N_9616,N_9628);
nand U9900 (N_9900,N_9669,N_9716);
and U9901 (N_9901,N_9757,N_9707);
nor U9902 (N_9902,N_9642,N_9767);
nor U9903 (N_9903,N_9614,N_9719);
or U9904 (N_9904,N_9686,N_9648);
nor U9905 (N_9905,N_9718,N_9738);
or U9906 (N_9906,N_9641,N_9728);
nand U9907 (N_9907,N_9728,N_9653);
nor U9908 (N_9908,N_9712,N_9673);
nand U9909 (N_9909,N_9646,N_9736);
or U9910 (N_9910,N_9645,N_9768);
and U9911 (N_9911,N_9701,N_9639);
or U9912 (N_9912,N_9606,N_9634);
xnor U9913 (N_9913,N_9633,N_9773);
xor U9914 (N_9914,N_9685,N_9717);
nand U9915 (N_9915,N_9781,N_9653);
nand U9916 (N_9916,N_9729,N_9609);
nor U9917 (N_9917,N_9704,N_9642);
nand U9918 (N_9918,N_9649,N_9662);
or U9919 (N_9919,N_9677,N_9795);
or U9920 (N_9920,N_9748,N_9703);
nor U9921 (N_9921,N_9611,N_9703);
and U9922 (N_9922,N_9713,N_9701);
and U9923 (N_9923,N_9684,N_9732);
nor U9924 (N_9924,N_9603,N_9741);
nand U9925 (N_9925,N_9643,N_9645);
nand U9926 (N_9926,N_9738,N_9679);
nand U9927 (N_9927,N_9798,N_9692);
nand U9928 (N_9928,N_9642,N_9664);
or U9929 (N_9929,N_9603,N_9781);
and U9930 (N_9930,N_9703,N_9734);
and U9931 (N_9931,N_9631,N_9615);
nand U9932 (N_9932,N_9753,N_9755);
and U9933 (N_9933,N_9734,N_9774);
or U9934 (N_9934,N_9634,N_9633);
or U9935 (N_9935,N_9698,N_9693);
xnor U9936 (N_9936,N_9711,N_9664);
or U9937 (N_9937,N_9675,N_9711);
nand U9938 (N_9938,N_9743,N_9707);
or U9939 (N_9939,N_9624,N_9641);
or U9940 (N_9940,N_9676,N_9626);
and U9941 (N_9941,N_9622,N_9616);
nor U9942 (N_9942,N_9708,N_9788);
nand U9943 (N_9943,N_9617,N_9745);
or U9944 (N_9944,N_9656,N_9744);
or U9945 (N_9945,N_9633,N_9658);
and U9946 (N_9946,N_9737,N_9635);
xor U9947 (N_9947,N_9764,N_9606);
nor U9948 (N_9948,N_9612,N_9681);
and U9949 (N_9949,N_9600,N_9717);
and U9950 (N_9950,N_9682,N_9620);
or U9951 (N_9951,N_9791,N_9789);
or U9952 (N_9952,N_9771,N_9774);
and U9953 (N_9953,N_9686,N_9635);
nor U9954 (N_9954,N_9655,N_9690);
and U9955 (N_9955,N_9689,N_9603);
or U9956 (N_9956,N_9632,N_9762);
nor U9957 (N_9957,N_9726,N_9730);
nor U9958 (N_9958,N_9722,N_9652);
xnor U9959 (N_9959,N_9655,N_9686);
or U9960 (N_9960,N_9780,N_9704);
nand U9961 (N_9961,N_9646,N_9732);
nand U9962 (N_9962,N_9743,N_9790);
or U9963 (N_9963,N_9659,N_9615);
or U9964 (N_9964,N_9651,N_9626);
and U9965 (N_9965,N_9792,N_9785);
and U9966 (N_9966,N_9638,N_9712);
nand U9967 (N_9967,N_9680,N_9776);
nand U9968 (N_9968,N_9763,N_9792);
nor U9969 (N_9969,N_9618,N_9790);
nand U9970 (N_9970,N_9692,N_9651);
nor U9971 (N_9971,N_9645,N_9629);
and U9972 (N_9972,N_9657,N_9672);
xor U9973 (N_9973,N_9646,N_9692);
nand U9974 (N_9974,N_9689,N_9634);
xor U9975 (N_9975,N_9631,N_9611);
xnor U9976 (N_9976,N_9766,N_9747);
nand U9977 (N_9977,N_9651,N_9640);
xnor U9978 (N_9978,N_9606,N_9673);
nand U9979 (N_9979,N_9782,N_9672);
nor U9980 (N_9980,N_9696,N_9686);
and U9981 (N_9981,N_9752,N_9734);
or U9982 (N_9982,N_9651,N_9747);
nand U9983 (N_9983,N_9786,N_9691);
and U9984 (N_9984,N_9609,N_9655);
and U9985 (N_9985,N_9674,N_9754);
and U9986 (N_9986,N_9608,N_9711);
nor U9987 (N_9987,N_9682,N_9779);
nand U9988 (N_9988,N_9629,N_9754);
nand U9989 (N_9989,N_9674,N_9646);
or U9990 (N_9990,N_9602,N_9794);
and U9991 (N_9991,N_9741,N_9700);
nor U9992 (N_9992,N_9600,N_9654);
or U9993 (N_9993,N_9641,N_9696);
nand U9994 (N_9994,N_9706,N_9743);
nand U9995 (N_9995,N_9659,N_9641);
or U9996 (N_9996,N_9792,N_9777);
nand U9997 (N_9997,N_9658,N_9776);
and U9998 (N_9998,N_9764,N_9701);
xor U9999 (N_9999,N_9698,N_9618);
and U10000 (N_10000,N_9812,N_9884);
and U10001 (N_10001,N_9874,N_9817);
nand U10002 (N_10002,N_9842,N_9808);
or U10003 (N_10003,N_9848,N_9905);
or U10004 (N_10004,N_9939,N_9959);
nor U10005 (N_10005,N_9908,N_9953);
nand U10006 (N_10006,N_9846,N_9837);
nand U10007 (N_10007,N_9913,N_9919);
and U10008 (N_10008,N_9920,N_9886);
nand U10009 (N_10009,N_9967,N_9902);
nor U10010 (N_10010,N_9809,N_9963);
and U10011 (N_10011,N_9910,N_9966);
nor U10012 (N_10012,N_9945,N_9960);
nand U10013 (N_10013,N_9813,N_9841);
and U10014 (N_10014,N_9906,N_9972);
and U10015 (N_10015,N_9896,N_9801);
and U10016 (N_10016,N_9830,N_9851);
nand U10017 (N_10017,N_9974,N_9880);
nand U10018 (N_10018,N_9980,N_9968);
nor U10019 (N_10019,N_9863,N_9868);
or U10020 (N_10020,N_9958,N_9975);
and U10021 (N_10021,N_9956,N_9893);
or U10022 (N_10022,N_9971,N_9864);
or U10023 (N_10023,N_9836,N_9997);
and U10024 (N_10024,N_9933,N_9844);
nand U10025 (N_10025,N_9877,N_9954);
nor U10026 (N_10026,N_9934,N_9810);
or U10027 (N_10027,N_9938,N_9860);
nor U10028 (N_10028,N_9949,N_9914);
nand U10029 (N_10029,N_9951,N_9823);
and U10030 (N_10030,N_9940,N_9927);
nand U10031 (N_10031,N_9845,N_9921);
nand U10032 (N_10032,N_9881,N_9917);
nand U10033 (N_10033,N_9982,N_9947);
or U10034 (N_10034,N_9964,N_9878);
or U10035 (N_10035,N_9911,N_9818);
and U10036 (N_10036,N_9916,N_9936);
and U10037 (N_10037,N_9876,N_9998);
and U10038 (N_10038,N_9932,N_9983);
nor U10039 (N_10039,N_9888,N_9946);
and U10040 (N_10040,N_9981,N_9875);
nor U10041 (N_10041,N_9929,N_9814);
or U10042 (N_10042,N_9977,N_9885);
nand U10043 (N_10043,N_9843,N_9952);
nand U10044 (N_10044,N_9850,N_9832);
or U10045 (N_10045,N_9866,N_9918);
or U10046 (N_10046,N_9827,N_9811);
and U10047 (N_10047,N_9815,N_9990);
and U10048 (N_10048,N_9838,N_9804);
nand U10049 (N_10049,N_9870,N_9904);
or U10050 (N_10050,N_9834,N_9943);
or U10051 (N_10051,N_9969,N_9987);
or U10052 (N_10052,N_9907,N_9852);
and U10053 (N_10053,N_9992,N_9829);
or U10054 (N_10054,N_9805,N_9819);
and U10055 (N_10055,N_9923,N_9995);
or U10056 (N_10056,N_9942,N_9991);
and U10057 (N_10057,N_9894,N_9857);
and U10058 (N_10058,N_9999,N_9883);
and U10059 (N_10059,N_9873,N_9891);
or U10060 (N_10060,N_9901,N_9978);
and U10061 (N_10061,N_9835,N_9803);
or U10062 (N_10062,N_9993,N_9909);
nand U10063 (N_10063,N_9900,N_9915);
and U10064 (N_10064,N_9965,N_9869);
or U10065 (N_10065,N_9824,N_9825);
and U10066 (N_10066,N_9985,N_9853);
and U10067 (N_10067,N_9897,N_9833);
nor U10068 (N_10068,N_9889,N_9944);
and U10069 (N_10069,N_9859,N_9890);
or U10070 (N_10070,N_9849,N_9950);
nand U10071 (N_10071,N_9957,N_9899);
nor U10072 (N_10072,N_9872,N_9882);
nor U10073 (N_10073,N_9931,N_9831);
and U10074 (N_10074,N_9986,N_9800);
or U10075 (N_10075,N_9979,N_9925);
and U10076 (N_10076,N_9822,N_9996);
nor U10077 (N_10077,N_9924,N_9955);
nor U10078 (N_10078,N_9816,N_9922);
nand U10079 (N_10079,N_9984,N_9970);
nand U10080 (N_10080,N_9898,N_9926);
nand U10081 (N_10081,N_9976,N_9903);
and U10082 (N_10082,N_9871,N_9840);
and U10083 (N_10083,N_9821,N_9892);
nand U10084 (N_10084,N_9895,N_9826);
or U10085 (N_10085,N_9855,N_9941);
or U10086 (N_10086,N_9928,N_9839);
xor U10087 (N_10087,N_9973,N_9807);
or U10088 (N_10088,N_9865,N_9937);
nor U10089 (N_10089,N_9994,N_9962);
nor U10090 (N_10090,N_9989,N_9854);
nor U10091 (N_10091,N_9867,N_9820);
and U10092 (N_10092,N_9935,N_9847);
and U10093 (N_10093,N_9856,N_9861);
nand U10094 (N_10094,N_9802,N_9887);
nor U10095 (N_10095,N_9988,N_9912);
and U10096 (N_10096,N_9806,N_9879);
nand U10097 (N_10097,N_9858,N_9862);
nor U10098 (N_10098,N_9828,N_9961);
nor U10099 (N_10099,N_9948,N_9930);
nor U10100 (N_10100,N_9874,N_9983);
nand U10101 (N_10101,N_9856,N_9927);
and U10102 (N_10102,N_9816,N_9979);
nand U10103 (N_10103,N_9817,N_9802);
nor U10104 (N_10104,N_9811,N_9918);
nor U10105 (N_10105,N_9938,N_9884);
nor U10106 (N_10106,N_9924,N_9882);
nand U10107 (N_10107,N_9992,N_9916);
nand U10108 (N_10108,N_9806,N_9989);
and U10109 (N_10109,N_9911,N_9863);
nor U10110 (N_10110,N_9976,N_9959);
nand U10111 (N_10111,N_9949,N_9818);
and U10112 (N_10112,N_9869,N_9899);
and U10113 (N_10113,N_9925,N_9809);
or U10114 (N_10114,N_9938,N_9967);
nor U10115 (N_10115,N_9911,N_9982);
and U10116 (N_10116,N_9914,N_9963);
nand U10117 (N_10117,N_9957,N_9939);
or U10118 (N_10118,N_9982,N_9887);
xor U10119 (N_10119,N_9991,N_9906);
or U10120 (N_10120,N_9961,N_9831);
nand U10121 (N_10121,N_9818,N_9804);
nor U10122 (N_10122,N_9892,N_9835);
nand U10123 (N_10123,N_9833,N_9857);
nor U10124 (N_10124,N_9870,N_9922);
nand U10125 (N_10125,N_9833,N_9920);
nor U10126 (N_10126,N_9808,N_9881);
xor U10127 (N_10127,N_9870,N_9990);
and U10128 (N_10128,N_9916,N_9805);
and U10129 (N_10129,N_9848,N_9992);
nand U10130 (N_10130,N_9986,N_9836);
and U10131 (N_10131,N_9985,N_9847);
nor U10132 (N_10132,N_9814,N_9909);
and U10133 (N_10133,N_9951,N_9924);
and U10134 (N_10134,N_9821,N_9836);
or U10135 (N_10135,N_9985,N_9818);
or U10136 (N_10136,N_9941,N_9862);
and U10137 (N_10137,N_9892,N_9875);
or U10138 (N_10138,N_9890,N_9955);
nand U10139 (N_10139,N_9976,N_9859);
or U10140 (N_10140,N_9981,N_9994);
nor U10141 (N_10141,N_9810,N_9868);
nor U10142 (N_10142,N_9873,N_9860);
and U10143 (N_10143,N_9807,N_9833);
nand U10144 (N_10144,N_9897,N_9998);
nand U10145 (N_10145,N_9920,N_9938);
or U10146 (N_10146,N_9848,N_9907);
nand U10147 (N_10147,N_9988,N_9813);
nand U10148 (N_10148,N_9877,N_9994);
and U10149 (N_10149,N_9994,N_9840);
nand U10150 (N_10150,N_9846,N_9901);
or U10151 (N_10151,N_9969,N_9835);
nor U10152 (N_10152,N_9922,N_9952);
or U10153 (N_10153,N_9910,N_9896);
nand U10154 (N_10154,N_9901,N_9916);
and U10155 (N_10155,N_9879,N_9890);
or U10156 (N_10156,N_9866,N_9831);
nand U10157 (N_10157,N_9802,N_9860);
nor U10158 (N_10158,N_9858,N_9996);
xor U10159 (N_10159,N_9806,N_9869);
nand U10160 (N_10160,N_9800,N_9880);
xnor U10161 (N_10161,N_9838,N_9958);
nor U10162 (N_10162,N_9948,N_9839);
nand U10163 (N_10163,N_9972,N_9814);
or U10164 (N_10164,N_9863,N_9974);
nand U10165 (N_10165,N_9943,N_9893);
nand U10166 (N_10166,N_9951,N_9808);
or U10167 (N_10167,N_9927,N_9883);
nand U10168 (N_10168,N_9818,N_9921);
and U10169 (N_10169,N_9903,N_9877);
nand U10170 (N_10170,N_9959,N_9837);
nor U10171 (N_10171,N_9945,N_9878);
and U10172 (N_10172,N_9936,N_9933);
or U10173 (N_10173,N_9857,N_9925);
nand U10174 (N_10174,N_9856,N_9819);
or U10175 (N_10175,N_9939,N_9838);
nand U10176 (N_10176,N_9890,N_9963);
nor U10177 (N_10177,N_9955,N_9819);
and U10178 (N_10178,N_9981,N_9978);
nor U10179 (N_10179,N_9992,N_9823);
nand U10180 (N_10180,N_9821,N_9883);
and U10181 (N_10181,N_9892,N_9996);
nor U10182 (N_10182,N_9877,N_9895);
nand U10183 (N_10183,N_9847,N_9974);
or U10184 (N_10184,N_9929,N_9946);
and U10185 (N_10185,N_9927,N_9963);
and U10186 (N_10186,N_9836,N_9893);
nand U10187 (N_10187,N_9921,N_9963);
or U10188 (N_10188,N_9828,N_9824);
and U10189 (N_10189,N_9848,N_9858);
or U10190 (N_10190,N_9867,N_9928);
nand U10191 (N_10191,N_9923,N_9934);
and U10192 (N_10192,N_9975,N_9871);
nand U10193 (N_10193,N_9814,N_9870);
and U10194 (N_10194,N_9810,N_9943);
and U10195 (N_10195,N_9800,N_9908);
nor U10196 (N_10196,N_9842,N_9996);
xor U10197 (N_10197,N_9941,N_9926);
nor U10198 (N_10198,N_9929,N_9820);
nor U10199 (N_10199,N_9877,N_9929);
nand U10200 (N_10200,N_10063,N_10162);
nand U10201 (N_10201,N_10061,N_10176);
nor U10202 (N_10202,N_10066,N_10044);
and U10203 (N_10203,N_10177,N_10160);
or U10204 (N_10204,N_10083,N_10191);
and U10205 (N_10205,N_10134,N_10064);
nor U10206 (N_10206,N_10067,N_10185);
nand U10207 (N_10207,N_10169,N_10183);
xor U10208 (N_10208,N_10079,N_10068);
xor U10209 (N_10209,N_10156,N_10190);
nand U10210 (N_10210,N_10195,N_10171);
or U10211 (N_10211,N_10010,N_10000);
nor U10212 (N_10212,N_10126,N_10172);
or U10213 (N_10213,N_10035,N_10046);
or U10214 (N_10214,N_10076,N_10019);
nor U10215 (N_10215,N_10097,N_10138);
nand U10216 (N_10216,N_10008,N_10105);
or U10217 (N_10217,N_10065,N_10011);
xor U10218 (N_10218,N_10012,N_10121);
or U10219 (N_10219,N_10143,N_10056);
nor U10220 (N_10220,N_10043,N_10086);
xnor U10221 (N_10221,N_10047,N_10096);
nand U10222 (N_10222,N_10193,N_10118);
and U10223 (N_10223,N_10139,N_10005);
or U10224 (N_10224,N_10125,N_10040);
or U10225 (N_10225,N_10137,N_10114);
or U10226 (N_10226,N_10099,N_10130);
and U10227 (N_10227,N_10009,N_10145);
nor U10228 (N_10228,N_10036,N_10020);
xnor U10229 (N_10229,N_10117,N_10164);
nor U10230 (N_10230,N_10165,N_10007);
xnor U10231 (N_10231,N_10136,N_10075);
and U10232 (N_10232,N_10186,N_10030);
xor U10233 (N_10233,N_10053,N_10018);
and U10234 (N_10234,N_10052,N_10017);
and U10235 (N_10235,N_10074,N_10198);
nand U10236 (N_10236,N_10022,N_10051);
or U10237 (N_10237,N_10016,N_10108);
or U10238 (N_10238,N_10199,N_10116);
nor U10239 (N_10239,N_10194,N_10098);
xor U10240 (N_10240,N_10102,N_10111);
and U10241 (N_10241,N_10129,N_10034);
nand U10242 (N_10242,N_10015,N_10140);
nand U10243 (N_10243,N_10039,N_10158);
nand U10244 (N_10244,N_10178,N_10101);
nor U10245 (N_10245,N_10014,N_10123);
and U10246 (N_10246,N_10106,N_10104);
or U10247 (N_10247,N_10084,N_10153);
and U10248 (N_10248,N_10163,N_10023);
and U10249 (N_10249,N_10058,N_10112);
or U10250 (N_10250,N_10124,N_10002);
and U10251 (N_10251,N_10045,N_10090);
or U10252 (N_10252,N_10071,N_10166);
and U10253 (N_10253,N_10080,N_10003);
nor U10254 (N_10254,N_10155,N_10196);
and U10255 (N_10255,N_10062,N_10154);
nor U10256 (N_10256,N_10142,N_10006);
nor U10257 (N_10257,N_10146,N_10001);
and U10258 (N_10258,N_10069,N_10004);
nand U10259 (N_10259,N_10159,N_10100);
or U10260 (N_10260,N_10149,N_10024);
nor U10261 (N_10261,N_10152,N_10060);
and U10262 (N_10262,N_10093,N_10073);
nor U10263 (N_10263,N_10048,N_10025);
nand U10264 (N_10264,N_10141,N_10148);
nand U10265 (N_10265,N_10031,N_10187);
nand U10266 (N_10266,N_10147,N_10050);
or U10267 (N_10267,N_10055,N_10122);
nand U10268 (N_10268,N_10042,N_10110);
xnor U10269 (N_10269,N_10192,N_10085);
nor U10270 (N_10270,N_10174,N_10188);
and U10271 (N_10271,N_10131,N_10173);
nor U10272 (N_10272,N_10095,N_10054);
or U10273 (N_10273,N_10120,N_10197);
and U10274 (N_10274,N_10021,N_10113);
nand U10275 (N_10275,N_10115,N_10170);
or U10276 (N_10276,N_10092,N_10167);
xor U10277 (N_10277,N_10070,N_10027);
nor U10278 (N_10278,N_10026,N_10189);
nor U10279 (N_10279,N_10144,N_10057);
and U10280 (N_10280,N_10059,N_10119);
and U10281 (N_10281,N_10161,N_10088);
or U10282 (N_10282,N_10082,N_10091);
nand U10283 (N_10283,N_10151,N_10135);
nand U10284 (N_10284,N_10109,N_10081);
nor U10285 (N_10285,N_10182,N_10038);
nand U10286 (N_10286,N_10127,N_10078);
and U10287 (N_10287,N_10077,N_10175);
or U10288 (N_10288,N_10157,N_10089);
and U10289 (N_10289,N_10028,N_10133);
or U10290 (N_10290,N_10184,N_10168);
xor U10291 (N_10291,N_10132,N_10049);
or U10292 (N_10292,N_10029,N_10032);
and U10293 (N_10293,N_10033,N_10103);
nand U10294 (N_10294,N_10087,N_10128);
nor U10295 (N_10295,N_10094,N_10107);
nor U10296 (N_10296,N_10041,N_10181);
nor U10297 (N_10297,N_10037,N_10150);
and U10298 (N_10298,N_10013,N_10180);
nor U10299 (N_10299,N_10179,N_10072);
nand U10300 (N_10300,N_10001,N_10111);
xor U10301 (N_10301,N_10037,N_10189);
nor U10302 (N_10302,N_10117,N_10096);
nor U10303 (N_10303,N_10133,N_10074);
nor U10304 (N_10304,N_10059,N_10096);
or U10305 (N_10305,N_10148,N_10164);
or U10306 (N_10306,N_10134,N_10017);
nor U10307 (N_10307,N_10008,N_10161);
nand U10308 (N_10308,N_10013,N_10073);
nand U10309 (N_10309,N_10038,N_10053);
and U10310 (N_10310,N_10039,N_10075);
nand U10311 (N_10311,N_10065,N_10094);
or U10312 (N_10312,N_10160,N_10080);
xnor U10313 (N_10313,N_10108,N_10018);
nand U10314 (N_10314,N_10008,N_10037);
and U10315 (N_10315,N_10139,N_10145);
nand U10316 (N_10316,N_10141,N_10080);
or U10317 (N_10317,N_10173,N_10012);
or U10318 (N_10318,N_10076,N_10045);
and U10319 (N_10319,N_10063,N_10019);
or U10320 (N_10320,N_10172,N_10104);
or U10321 (N_10321,N_10001,N_10190);
and U10322 (N_10322,N_10071,N_10084);
and U10323 (N_10323,N_10159,N_10016);
xor U10324 (N_10324,N_10095,N_10037);
nand U10325 (N_10325,N_10195,N_10026);
and U10326 (N_10326,N_10051,N_10046);
or U10327 (N_10327,N_10055,N_10023);
or U10328 (N_10328,N_10075,N_10153);
or U10329 (N_10329,N_10129,N_10110);
or U10330 (N_10330,N_10060,N_10037);
nor U10331 (N_10331,N_10116,N_10128);
nand U10332 (N_10332,N_10010,N_10185);
xor U10333 (N_10333,N_10022,N_10159);
nand U10334 (N_10334,N_10148,N_10000);
nor U10335 (N_10335,N_10022,N_10143);
nor U10336 (N_10336,N_10058,N_10048);
or U10337 (N_10337,N_10047,N_10182);
or U10338 (N_10338,N_10058,N_10145);
nor U10339 (N_10339,N_10000,N_10054);
and U10340 (N_10340,N_10004,N_10157);
nand U10341 (N_10341,N_10023,N_10123);
or U10342 (N_10342,N_10070,N_10043);
and U10343 (N_10343,N_10180,N_10023);
or U10344 (N_10344,N_10036,N_10136);
nor U10345 (N_10345,N_10083,N_10025);
nand U10346 (N_10346,N_10102,N_10091);
and U10347 (N_10347,N_10045,N_10010);
or U10348 (N_10348,N_10000,N_10172);
xor U10349 (N_10349,N_10030,N_10003);
nand U10350 (N_10350,N_10135,N_10085);
xor U10351 (N_10351,N_10119,N_10047);
and U10352 (N_10352,N_10080,N_10159);
nor U10353 (N_10353,N_10087,N_10152);
or U10354 (N_10354,N_10028,N_10113);
or U10355 (N_10355,N_10116,N_10148);
and U10356 (N_10356,N_10162,N_10191);
and U10357 (N_10357,N_10058,N_10158);
xor U10358 (N_10358,N_10100,N_10161);
or U10359 (N_10359,N_10064,N_10079);
nor U10360 (N_10360,N_10121,N_10148);
or U10361 (N_10361,N_10032,N_10127);
nor U10362 (N_10362,N_10030,N_10036);
or U10363 (N_10363,N_10058,N_10000);
and U10364 (N_10364,N_10004,N_10091);
or U10365 (N_10365,N_10068,N_10020);
or U10366 (N_10366,N_10141,N_10047);
nand U10367 (N_10367,N_10174,N_10181);
xnor U10368 (N_10368,N_10105,N_10098);
and U10369 (N_10369,N_10001,N_10158);
nand U10370 (N_10370,N_10080,N_10149);
or U10371 (N_10371,N_10131,N_10179);
or U10372 (N_10372,N_10026,N_10134);
nor U10373 (N_10373,N_10195,N_10022);
nor U10374 (N_10374,N_10158,N_10003);
nand U10375 (N_10375,N_10092,N_10152);
nand U10376 (N_10376,N_10132,N_10121);
nand U10377 (N_10377,N_10056,N_10064);
xnor U10378 (N_10378,N_10143,N_10100);
nor U10379 (N_10379,N_10132,N_10013);
nand U10380 (N_10380,N_10073,N_10157);
and U10381 (N_10381,N_10188,N_10189);
and U10382 (N_10382,N_10046,N_10136);
and U10383 (N_10383,N_10157,N_10146);
and U10384 (N_10384,N_10151,N_10077);
and U10385 (N_10385,N_10061,N_10146);
nor U10386 (N_10386,N_10084,N_10041);
or U10387 (N_10387,N_10149,N_10031);
nand U10388 (N_10388,N_10119,N_10148);
and U10389 (N_10389,N_10062,N_10075);
or U10390 (N_10390,N_10057,N_10021);
nand U10391 (N_10391,N_10100,N_10002);
nor U10392 (N_10392,N_10098,N_10127);
and U10393 (N_10393,N_10015,N_10087);
nand U10394 (N_10394,N_10091,N_10058);
nor U10395 (N_10395,N_10077,N_10138);
nor U10396 (N_10396,N_10185,N_10150);
nand U10397 (N_10397,N_10016,N_10190);
nor U10398 (N_10398,N_10188,N_10180);
and U10399 (N_10399,N_10191,N_10047);
nand U10400 (N_10400,N_10298,N_10280);
xnor U10401 (N_10401,N_10394,N_10284);
and U10402 (N_10402,N_10219,N_10238);
and U10403 (N_10403,N_10385,N_10222);
nand U10404 (N_10404,N_10216,N_10335);
nor U10405 (N_10405,N_10362,N_10371);
and U10406 (N_10406,N_10381,N_10380);
nor U10407 (N_10407,N_10249,N_10342);
nand U10408 (N_10408,N_10339,N_10225);
nor U10409 (N_10409,N_10289,N_10368);
and U10410 (N_10410,N_10291,N_10200);
nand U10411 (N_10411,N_10207,N_10276);
xor U10412 (N_10412,N_10217,N_10221);
nand U10413 (N_10413,N_10377,N_10234);
or U10414 (N_10414,N_10333,N_10312);
or U10415 (N_10415,N_10345,N_10245);
or U10416 (N_10416,N_10259,N_10265);
nor U10417 (N_10417,N_10272,N_10290);
and U10418 (N_10418,N_10391,N_10205);
or U10419 (N_10419,N_10375,N_10322);
and U10420 (N_10420,N_10330,N_10305);
xor U10421 (N_10421,N_10328,N_10384);
nor U10422 (N_10422,N_10390,N_10370);
or U10423 (N_10423,N_10315,N_10373);
and U10424 (N_10424,N_10354,N_10310);
and U10425 (N_10425,N_10376,N_10383);
and U10426 (N_10426,N_10331,N_10395);
xnor U10427 (N_10427,N_10239,N_10283);
xor U10428 (N_10428,N_10348,N_10223);
xor U10429 (N_10429,N_10299,N_10211);
and U10430 (N_10430,N_10268,N_10338);
nand U10431 (N_10431,N_10267,N_10303);
or U10432 (N_10432,N_10227,N_10347);
nand U10433 (N_10433,N_10241,N_10349);
and U10434 (N_10434,N_10285,N_10398);
nor U10435 (N_10435,N_10336,N_10256);
nand U10436 (N_10436,N_10230,N_10316);
nand U10437 (N_10437,N_10296,N_10286);
nor U10438 (N_10438,N_10212,N_10399);
xnor U10439 (N_10439,N_10369,N_10271);
or U10440 (N_10440,N_10360,N_10334);
nor U10441 (N_10441,N_10387,N_10287);
xnor U10442 (N_10442,N_10246,N_10317);
or U10443 (N_10443,N_10357,N_10204);
and U10444 (N_10444,N_10228,N_10242);
or U10445 (N_10445,N_10311,N_10302);
nor U10446 (N_10446,N_10243,N_10215);
and U10447 (N_10447,N_10306,N_10363);
and U10448 (N_10448,N_10294,N_10300);
or U10449 (N_10449,N_10254,N_10233);
and U10450 (N_10450,N_10232,N_10214);
nor U10451 (N_10451,N_10277,N_10313);
nor U10452 (N_10452,N_10253,N_10206);
and U10453 (N_10453,N_10327,N_10393);
nor U10454 (N_10454,N_10237,N_10367);
nand U10455 (N_10455,N_10372,N_10351);
or U10456 (N_10456,N_10386,N_10374);
nor U10457 (N_10457,N_10364,N_10378);
or U10458 (N_10458,N_10325,N_10392);
and U10459 (N_10459,N_10355,N_10275);
nand U10460 (N_10460,N_10266,N_10208);
and U10461 (N_10461,N_10213,N_10274);
or U10462 (N_10462,N_10350,N_10292);
and U10463 (N_10463,N_10324,N_10320);
or U10464 (N_10464,N_10257,N_10252);
xor U10465 (N_10465,N_10201,N_10353);
xor U10466 (N_10466,N_10304,N_10326);
nor U10467 (N_10467,N_10341,N_10389);
nor U10468 (N_10468,N_10358,N_10321);
and U10469 (N_10469,N_10329,N_10282);
or U10470 (N_10470,N_10279,N_10361);
nor U10471 (N_10471,N_10301,N_10264);
nor U10472 (N_10472,N_10202,N_10220);
or U10473 (N_10473,N_10224,N_10382);
and U10474 (N_10474,N_10278,N_10270);
xnor U10475 (N_10475,N_10269,N_10247);
nor U10476 (N_10476,N_10293,N_10260);
nor U10477 (N_10477,N_10344,N_10295);
and U10478 (N_10478,N_10262,N_10343);
nor U10479 (N_10479,N_10346,N_10314);
or U10480 (N_10480,N_10337,N_10203);
nor U10481 (N_10481,N_10226,N_10288);
nand U10482 (N_10482,N_10359,N_10235);
and U10483 (N_10483,N_10210,N_10308);
or U10484 (N_10484,N_10240,N_10229);
or U10485 (N_10485,N_10388,N_10396);
and U10486 (N_10486,N_10319,N_10356);
or U10487 (N_10487,N_10258,N_10250);
and U10488 (N_10488,N_10281,N_10352);
and U10489 (N_10489,N_10379,N_10248);
and U10490 (N_10490,N_10323,N_10366);
nor U10491 (N_10491,N_10332,N_10340);
or U10492 (N_10492,N_10307,N_10261);
and U10493 (N_10493,N_10397,N_10263);
nand U10494 (N_10494,N_10209,N_10318);
or U10495 (N_10495,N_10273,N_10309);
or U10496 (N_10496,N_10236,N_10231);
nor U10497 (N_10497,N_10297,N_10218);
xnor U10498 (N_10498,N_10244,N_10251);
nand U10499 (N_10499,N_10365,N_10255);
and U10500 (N_10500,N_10241,N_10237);
or U10501 (N_10501,N_10234,N_10380);
nor U10502 (N_10502,N_10240,N_10237);
nand U10503 (N_10503,N_10281,N_10304);
nand U10504 (N_10504,N_10344,N_10305);
xor U10505 (N_10505,N_10399,N_10255);
and U10506 (N_10506,N_10319,N_10210);
or U10507 (N_10507,N_10345,N_10347);
xor U10508 (N_10508,N_10241,N_10385);
nand U10509 (N_10509,N_10203,N_10346);
nor U10510 (N_10510,N_10225,N_10210);
or U10511 (N_10511,N_10324,N_10341);
nor U10512 (N_10512,N_10290,N_10208);
and U10513 (N_10513,N_10311,N_10227);
nor U10514 (N_10514,N_10262,N_10314);
nor U10515 (N_10515,N_10298,N_10349);
and U10516 (N_10516,N_10377,N_10297);
and U10517 (N_10517,N_10229,N_10317);
nor U10518 (N_10518,N_10295,N_10247);
nor U10519 (N_10519,N_10234,N_10222);
or U10520 (N_10520,N_10369,N_10342);
nand U10521 (N_10521,N_10386,N_10347);
and U10522 (N_10522,N_10247,N_10296);
nand U10523 (N_10523,N_10347,N_10228);
and U10524 (N_10524,N_10378,N_10397);
nor U10525 (N_10525,N_10325,N_10381);
nor U10526 (N_10526,N_10296,N_10317);
or U10527 (N_10527,N_10356,N_10254);
and U10528 (N_10528,N_10321,N_10218);
nor U10529 (N_10529,N_10379,N_10398);
nand U10530 (N_10530,N_10345,N_10308);
nor U10531 (N_10531,N_10206,N_10305);
and U10532 (N_10532,N_10257,N_10369);
or U10533 (N_10533,N_10294,N_10302);
xnor U10534 (N_10534,N_10330,N_10378);
or U10535 (N_10535,N_10201,N_10337);
nor U10536 (N_10536,N_10209,N_10298);
nand U10537 (N_10537,N_10255,N_10243);
or U10538 (N_10538,N_10310,N_10240);
or U10539 (N_10539,N_10351,N_10263);
nor U10540 (N_10540,N_10386,N_10266);
or U10541 (N_10541,N_10277,N_10358);
nand U10542 (N_10542,N_10267,N_10309);
or U10543 (N_10543,N_10243,N_10225);
xor U10544 (N_10544,N_10355,N_10264);
and U10545 (N_10545,N_10391,N_10200);
or U10546 (N_10546,N_10377,N_10319);
or U10547 (N_10547,N_10215,N_10298);
nor U10548 (N_10548,N_10329,N_10270);
nor U10549 (N_10549,N_10293,N_10284);
nand U10550 (N_10550,N_10349,N_10293);
or U10551 (N_10551,N_10387,N_10274);
nor U10552 (N_10552,N_10261,N_10215);
or U10553 (N_10553,N_10219,N_10337);
xnor U10554 (N_10554,N_10376,N_10236);
xnor U10555 (N_10555,N_10292,N_10200);
nor U10556 (N_10556,N_10229,N_10227);
or U10557 (N_10557,N_10234,N_10207);
and U10558 (N_10558,N_10351,N_10302);
nor U10559 (N_10559,N_10206,N_10323);
nand U10560 (N_10560,N_10336,N_10289);
nand U10561 (N_10561,N_10217,N_10295);
xnor U10562 (N_10562,N_10246,N_10376);
xor U10563 (N_10563,N_10226,N_10399);
or U10564 (N_10564,N_10270,N_10206);
nand U10565 (N_10565,N_10329,N_10253);
nor U10566 (N_10566,N_10364,N_10310);
xor U10567 (N_10567,N_10337,N_10276);
nand U10568 (N_10568,N_10243,N_10283);
xor U10569 (N_10569,N_10358,N_10327);
xnor U10570 (N_10570,N_10243,N_10248);
nor U10571 (N_10571,N_10393,N_10259);
or U10572 (N_10572,N_10214,N_10394);
nand U10573 (N_10573,N_10347,N_10313);
xor U10574 (N_10574,N_10251,N_10262);
nand U10575 (N_10575,N_10336,N_10282);
and U10576 (N_10576,N_10269,N_10398);
and U10577 (N_10577,N_10293,N_10335);
nor U10578 (N_10578,N_10261,N_10394);
nand U10579 (N_10579,N_10230,N_10269);
nor U10580 (N_10580,N_10250,N_10351);
or U10581 (N_10581,N_10217,N_10386);
or U10582 (N_10582,N_10274,N_10376);
nor U10583 (N_10583,N_10340,N_10322);
nand U10584 (N_10584,N_10312,N_10304);
or U10585 (N_10585,N_10273,N_10265);
or U10586 (N_10586,N_10340,N_10244);
or U10587 (N_10587,N_10369,N_10252);
and U10588 (N_10588,N_10234,N_10370);
nand U10589 (N_10589,N_10306,N_10316);
and U10590 (N_10590,N_10247,N_10306);
nand U10591 (N_10591,N_10362,N_10363);
and U10592 (N_10592,N_10292,N_10331);
or U10593 (N_10593,N_10230,N_10264);
or U10594 (N_10594,N_10228,N_10206);
nor U10595 (N_10595,N_10201,N_10394);
or U10596 (N_10596,N_10279,N_10258);
nand U10597 (N_10597,N_10211,N_10278);
and U10598 (N_10598,N_10373,N_10235);
and U10599 (N_10599,N_10326,N_10203);
or U10600 (N_10600,N_10497,N_10422);
xor U10601 (N_10601,N_10565,N_10571);
and U10602 (N_10602,N_10404,N_10572);
nor U10603 (N_10603,N_10593,N_10455);
nand U10604 (N_10604,N_10413,N_10482);
nand U10605 (N_10605,N_10471,N_10436);
nand U10606 (N_10606,N_10530,N_10539);
nand U10607 (N_10607,N_10598,N_10420);
nor U10608 (N_10608,N_10462,N_10474);
nor U10609 (N_10609,N_10515,N_10480);
or U10610 (N_10610,N_10586,N_10536);
nor U10611 (N_10611,N_10492,N_10503);
and U10612 (N_10612,N_10564,N_10538);
xor U10613 (N_10613,N_10496,N_10444);
or U10614 (N_10614,N_10549,N_10533);
nand U10615 (N_10615,N_10412,N_10439);
and U10616 (N_10616,N_10575,N_10542);
or U10617 (N_10617,N_10518,N_10573);
or U10618 (N_10618,N_10451,N_10450);
nor U10619 (N_10619,N_10406,N_10464);
or U10620 (N_10620,N_10400,N_10402);
nand U10621 (N_10621,N_10475,N_10421);
nand U10622 (N_10622,N_10456,N_10485);
and U10623 (N_10623,N_10561,N_10558);
and U10624 (N_10624,N_10563,N_10448);
nand U10625 (N_10625,N_10452,N_10589);
or U10626 (N_10626,N_10559,N_10529);
nand U10627 (N_10627,N_10437,N_10591);
or U10628 (N_10628,N_10407,N_10583);
xor U10629 (N_10629,N_10554,N_10570);
nor U10630 (N_10630,N_10528,N_10423);
xnor U10631 (N_10631,N_10581,N_10524);
or U10632 (N_10632,N_10599,N_10434);
nor U10633 (N_10633,N_10576,N_10507);
and U10634 (N_10634,N_10535,N_10495);
nand U10635 (N_10635,N_10553,N_10499);
and U10636 (N_10636,N_10419,N_10425);
nor U10637 (N_10637,N_10566,N_10479);
and U10638 (N_10638,N_10458,N_10521);
xor U10639 (N_10639,N_10597,N_10476);
nand U10640 (N_10640,N_10552,N_10588);
nor U10641 (N_10641,N_10459,N_10442);
nand U10642 (N_10642,N_10494,N_10555);
or U10643 (N_10643,N_10433,N_10534);
and U10644 (N_10644,N_10526,N_10544);
nor U10645 (N_10645,N_10467,N_10537);
nand U10646 (N_10646,N_10473,N_10513);
or U10647 (N_10647,N_10424,N_10416);
xor U10648 (N_10648,N_10440,N_10584);
or U10649 (N_10649,N_10441,N_10569);
nor U10650 (N_10650,N_10405,N_10595);
and U10651 (N_10651,N_10582,N_10468);
or U10652 (N_10652,N_10527,N_10580);
or U10653 (N_10653,N_10415,N_10501);
or U10654 (N_10654,N_10532,N_10505);
nor U10655 (N_10655,N_10432,N_10506);
xor U10656 (N_10656,N_10401,N_10519);
nor U10657 (N_10657,N_10568,N_10435);
nand U10658 (N_10658,N_10484,N_10478);
and U10659 (N_10659,N_10548,N_10508);
xor U10660 (N_10660,N_10585,N_10556);
nor U10661 (N_10661,N_10483,N_10523);
and U10662 (N_10662,N_10410,N_10500);
nor U10663 (N_10663,N_10481,N_10562);
or U10664 (N_10664,N_10531,N_10460);
nor U10665 (N_10665,N_10541,N_10461);
nand U10666 (N_10666,N_10417,N_10594);
or U10667 (N_10667,N_10550,N_10587);
or U10668 (N_10668,N_10486,N_10428);
or U10669 (N_10669,N_10574,N_10487);
nand U10670 (N_10670,N_10511,N_10414);
and U10671 (N_10671,N_10517,N_10463);
and U10672 (N_10672,N_10466,N_10430);
nor U10673 (N_10673,N_10446,N_10431);
or U10674 (N_10674,N_10509,N_10590);
or U10675 (N_10675,N_10438,N_10545);
nor U10676 (N_10676,N_10477,N_10514);
or U10677 (N_10677,N_10411,N_10596);
nand U10678 (N_10678,N_10488,N_10578);
nor U10679 (N_10679,N_10546,N_10510);
nor U10680 (N_10680,N_10470,N_10427);
nand U10681 (N_10681,N_10445,N_10490);
and U10682 (N_10682,N_10512,N_10469);
and U10683 (N_10683,N_10498,N_10560);
or U10684 (N_10684,N_10465,N_10567);
or U10685 (N_10685,N_10449,N_10429);
or U10686 (N_10686,N_10547,N_10403);
xor U10687 (N_10687,N_10525,N_10489);
xnor U10688 (N_10688,N_10408,N_10516);
nor U10689 (N_10689,N_10577,N_10543);
nand U10690 (N_10690,N_10453,N_10520);
nor U10691 (N_10691,N_10540,N_10502);
nand U10692 (N_10692,N_10454,N_10557);
nand U10693 (N_10693,N_10579,N_10443);
or U10694 (N_10694,N_10551,N_10418);
or U10695 (N_10695,N_10493,N_10426);
and U10696 (N_10696,N_10522,N_10409);
nor U10697 (N_10697,N_10457,N_10504);
nor U10698 (N_10698,N_10491,N_10472);
nor U10699 (N_10699,N_10592,N_10447);
or U10700 (N_10700,N_10546,N_10520);
or U10701 (N_10701,N_10578,N_10509);
xor U10702 (N_10702,N_10550,N_10492);
or U10703 (N_10703,N_10523,N_10413);
and U10704 (N_10704,N_10490,N_10431);
xor U10705 (N_10705,N_10572,N_10533);
xor U10706 (N_10706,N_10501,N_10512);
nor U10707 (N_10707,N_10595,N_10458);
nor U10708 (N_10708,N_10429,N_10539);
xor U10709 (N_10709,N_10520,N_10458);
nand U10710 (N_10710,N_10422,N_10555);
nand U10711 (N_10711,N_10526,N_10432);
nor U10712 (N_10712,N_10531,N_10512);
or U10713 (N_10713,N_10405,N_10466);
nand U10714 (N_10714,N_10498,N_10447);
and U10715 (N_10715,N_10486,N_10514);
nor U10716 (N_10716,N_10451,N_10555);
xnor U10717 (N_10717,N_10554,N_10563);
nor U10718 (N_10718,N_10517,N_10577);
and U10719 (N_10719,N_10474,N_10545);
nor U10720 (N_10720,N_10421,N_10509);
or U10721 (N_10721,N_10556,N_10564);
nor U10722 (N_10722,N_10510,N_10584);
nor U10723 (N_10723,N_10496,N_10449);
or U10724 (N_10724,N_10508,N_10595);
nand U10725 (N_10725,N_10462,N_10578);
nor U10726 (N_10726,N_10586,N_10450);
nand U10727 (N_10727,N_10418,N_10597);
nor U10728 (N_10728,N_10472,N_10418);
nor U10729 (N_10729,N_10461,N_10474);
xor U10730 (N_10730,N_10458,N_10561);
and U10731 (N_10731,N_10404,N_10450);
nand U10732 (N_10732,N_10514,N_10560);
and U10733 (N_10733,N_10515,N_10452);
or U10734 (N_10734,N_10526,N_10581);
and U10735 (N_10735,N_10460,N_10474);
xor U10736 (N_10736,N_10487,N_10599);
and U10737 (N_10737,N_10422,N_10419);
or U10738 (N_10738,N_10401,N_10568);
or U10739 (N_10739,N_10453,N_10525);
or U10740 (N_10740,N_10489,N_10418);
nor U10741 (N_10741,N_10454,N_10416);
xor U10742 (N_10742,N_10599,N_10582);
nor U10743 (N_10743,N_10461,N_10565);
xor U10744 (N_10744,N_10488,N_10428);
nor U10745 (N_10745,N_10584,N_10420);
nand U10746 (N_10746,N_10521,N_10543);
nor U10747 (N_10747,N_10446,N_10547);
or U10748 (N_10748,N_10415,N_10599);
or U10749 (N_10749,N_10584,N_10598);
nor U10750 (N_10750,N_10447,N_10412);
or U10751 (N_10751,N_10567,N_10488);
nor U10752 (N_10752,N_10417,N_10435);
and U10753 (N_10753,N_10475,N_10452);
nand U10754 (N_10754,N_10474,N_10576);
nor U10755 (N_10755,N_10591,N_10491);
and U10756 (N_10756,N_10514,N_10425);
xor U10757 (N_10757,N_10536,N_10457);
nand U10758 (N_10758,N_10581,N_10530);
xnor U10759 (N_10759,N_10540,N_10411);
and U10760 (N_10760,N_10497,N_10500);
nand U10761 (N_10761,N_10486,N_10410);
nand U10762 (N_10762,N_10502,N_10555);
nor U10763 (N_10763,N_10591,N_10582);
or U10764 (N_10764,N_10424,N_10436);
or U10765 (N_10765,N_10429,N_10574);
xnor U10766 (N_10766,N_10518,N_10416);
nand U10767 (N_10767,N_10530,N_10426);
nand U10768 (N_10768,N_10538,N_10590);
and U10769 (N_10769,N_10568,N_10412);
or U10770 (N_10770,N_10450,N_10543);
or U10771 (N_10771,N_10431,N_10503);
nand U10772 (N_10772,N_10457,N_10426);
and U10773 (N_10773,N_10513,N_10509);
nor U10774 (N_10774,N_10442,N_10497);
nand U10775 (N_10775,N_10458,N_10465);
nand U10776 (N_10776,N_10481,N_10572);
nand U10777 (N_10777,N_10416,N_10412);
nand U10778 (N_10778,N_10478,N_10532);
or U10779 (N_10779,N_10495,N_10415);
or U10780 (N_10780,N_10444,N_10475);
nor U10781 (N_10781,N_10496,N_10499);
and U10782 (N_10782,N_10563,N_10539);
and U10783 (N_10783,N_10479,N_10435);
nor U10784 (N_10784,N_10455,N_10551);
and U10785 (N_10785,N_10553,N_10548);
and U10786 (N_10786,N_10595,N_10407);
xor U10787 (N_10787,N_10448,N_10494);
or U10788 (N_10788,N_10534,N_10528);
or U10789 (N_10789,N_10490,N_10494);
nand U10790 (N_10790,N_10561,N_10591);
nor U10791 (N_10791,N_10585,N_10506);
and U10792 (N_10792,N_10574,N_10534);
or U10793 (N_10793,N_10414,N_10512);
nor U10794 (N_10794,N_10530,N_10439);
or U10795 (N_10795,N_10505,N_10427);
or U10796 (N_10796,N_10559,N_10548);
nor U10797 (N_10797,N_10530,N_10551);
xnor U10798 (N_10798,N_10485,N_10559);
and U10799 (N_10799,N_10571,N_10576);
nor U10800 (N_10800,N_10688,N_10754);
nand U10801 (N_10801,N_10682,N_10609);
or U10802 (N_10802,N_10710,N_10641);
and U10803 (N_10803,N_10716,N_10666);
and U10804 (N_10804,N_10635,N_10736);
and U10805 (N_10805,N_10735,N_10612);
or U10806 (N_10806,N_10604,N_10606);
xnor U10807 (N_10807,N_10611,N_10762);
or U10808 (N_10808,N_10698,N_10605);
and U10809 (N_10809,N_10654,N_10773);
nand U10810 (N_10810,N_10610,N_10625);
nor U10811 (N_10811,N_10731,N_10700);
nand U10812 (N_10812,N_10781,N_10768);
nand U10813 (N_10813,N_10628,N_10653);
nand U10814 (N_10814,N_10633,N_10697);
and U10815 (N_10815,N_10739,N_10744);
nor U10816 (N_10816,N_10786,N_10657);
or U10817 (N_10817,N_10707,N_10656);
or U10818 (N_10818,N_10699,N_10780);
nand U10819 (N_10819,N_10703,N_10619);
and U10820 (N_10820,N_10718,N_10752);
nor U10821 (N_10821,N_10730,N_10713);
and U10822 (N_10822,N_10791,N_10749);
and U10823 (N_10823,N_10663,N_10681);
or U10824 (N_10824,N_10759,N_10709);
or U10825 (N_10825,N_10689,N_10651);
nor U10826 (N_10826,N_10683,N_10799);
nand U10827 (N_10827,N_10690,N_10636);
nor U10828 (N_10828,N_10643,N_10722);
or U10829 (N_10829,N_10797,N_10741);
nand U10830 (N_10830,N_10670,N_10783);
nand U10831 (N_10831,N_10669,N_10665);
nor U10832 (N_10832,N_10715,N_10789);
and U10833 (N_10833,N_10765,N_10694);
nor U10834 (N_10834,N_10672,N_10761);
or U10835 (N_10835,N_10734,N_10705);
or U10836 (N_10836,N_10602,N_10687);
or U10837 (N_10837,N_10766,N_10649);
and U10838 (N_10838,N_10652,N_10679);
nand U10839 (N_10839,N_10720,N_10678);
nor U10840 (N_10840,N_10695,N_10756);
nand U10841 (N_10841,N_10757,N_10711);
or U10842 (N_10842,N_10684,N_10647);
or U10843 (N_10843,N_10737,N_10769);
and U10844 (N_10844,N_10701,N_10732);
or U10845 (N_10845,N_10753,N_10637);
nand U10846 (N_10846,N_10788,N_10717);
and U10847 (N_10847,N_10616,N_10618);
or U10848 (N_10848,N_10747,N_10660);
and U10849 (N_10849,N_10659,N_10621);
or U10850 (N_10850,N_10620,N_10685);
nand U10851 (N_10851,N_10726,N_10784);
nor U10852 (N_10852,N_10631,N_10764);
or U10853 (N_10853,N_10686,N_10646);
nor U10854 (N_10854,N_10740,N_10785);
nor U10855 (N_10855,N_10738,N_10680);
and U10856 (N_10856,N_10622,N_10630);
and U10857 (N_10857,N_10742,N_10648);
nand U10858 (N_10858,N_10640,N_10650);
or U10859 (N_10859,N_10658,N_10794);
nor U10860 (N_10860,N_10692,N_10645);
nand U10861 (N_10861,N_10607,N_10760);
nor U10862 (N_10862,N_10626,N_10639);
nand U10863 (N_10863,N_10728,N_10704);
and U10864 (N_10864,N_10706,N_10774);
or U10865 (N_10865,N_10623,N_10721);
nor U10866 (N_10866,N_10798,N_10746);
and U10867 (N_10867,N_10733,N_10796);
nand U10868 (N_10868,N_10615,N_10727);
nor U10869 (N_10869,N_10763,N_10696);
xnor U10870 (N_10870,N_10714,N_10787);
or U10871 (N_10871,N_10691,N_10674);
and U10872 (N_10872,N_10632,N_10603);
nor U10873 (N_10873,N_10751,N_10677);
or U10874 (N_10874,N_10624,N_10771);
xnor U10875 (N_10875,N_10702,N_10782);
and U10876 (N_10876,N_10613,N_10675);
and U10877 (N_10877,N_10617,N_10790);
nor U10878 (N_10878,N_10776,N_10725);
nor U10879 (N_10879,N_10664,N_10792);
xor U10880 (N_10880,N_10661,N_10608);
nor U10881 (N_10881,N_10668,N_10748);
nor U10882 (N_10882,N_10712,N_10758);
and U10883 (N_10883,N_10601,N_10745);
nand U10884 (N_10884,N_10655,N_10723);
or U10885 (N_10885,N_10767,N_10662);
nor U10886 (N_10886,N_10778,N_10693);
nor U10887 (N_10887,N_10775,N_10779);
nor U10888 (N_10888,N_10642,N_10724);
nand U10889 (N_10889,N_10638,N_10772);
nand U10890 (N_10890,N_10750,N_10793);
xnor U10891 (N_10891,N_10770,N_10671);
and U10892 (N_10892,N_10627,N_10708);
nand U10893 (N_10893,N_10600,N_10629);
nor U10894 (N_10894,N_10676,N_10719);
and U10895 (N_10895,N_10777,N_10634);
nand U10896 (N_10896,N_10743,N_10755);
or U10897 (N_10897,N_10795,N_10614);
or U10898 (N_10898,N_10644,N_10729);
nand U10899 (N_10899,N_10667,N_10673);
nor U10900 (N_10900,N_10633,N_10661);
or U10901 (N_10901,N_10650,N_10664);
and U10902 (N_10902,N_10722,N_10626);
and U10903 (N_10903,N_10761,N_10748);
nor U10904 (N_10904,N_10785,N_10604);
or U10905 (N_10905,N_10718,N_10753);
xor U10906 (N_10906,N_10656,N_10791);
nand U10907 (N_10907,N_10647,N_10749);
xor U10908 (N_10908,N_10753,N_10686);
or U10909 (N_10909,N_10678,N_10710);
or U10910 (N_10910,N_10719,N_10718);
or U10911 (N_10911,N_10691,N_10734);
and U10912 (N_10912,N_10792,N_10746);
nand U10913 (N_10913,N_10750,N_10787);
and U10914 (N_10914,N_10661,N_10718);
nand U10915 (N_10915,N_10738,N_10656);
nor U10916 (N_10916,N_10784,N_10608);
nor U10917 (N_10917,N_10748,N_10651);
nor U10918 (N_10918,N_10608,N_10610);
and U10919 (N_10919,N_10676,N_10792);
xnor U10920 (N_10920,N_10751,N_10774);
nand U10921 (N_10921,N_10654,N_10644);
and U10922 (N_10922,N_10739,N_10711);
and U10923 (N_10923,N_10770,N_10629);
nand U10924 (N_10924,N_10784,N_10738);
and U10925 (N_10925,N_10771,N_10748);
and U10926 (N_10926,N_10752,N_10753);
or U10927 (N_10927,N_10696,N_10759);
nor U10928 (N_10928,N_10767,N_10616);
or U10929 (N_10929,N_10744,N_10786);
and U10930 (N_10930,N_10743,N_10715);
nor U10931 (N_10931,N_10663,N_10682);
nor U10932 (N_10932,N_10652,N_10637);
or U10933 (N_10933,N_10688,N_10609);
or U10934 (N_10934,N_10649,N_10627);
nand U10935 (N_10935,N_10681,N_10721);
xor U10936 (N_10936,N_10726,N_10705);
or U10937 (N_10937,N_10604,N_10660);
and U10938 (N_10938,N_10635,N_10707);
and U10939 (N_10939,N_10723,N_10792);
and U10940 (N_10940,N_10637,N_10641);
and U10941 (N_10941,N_10762,N_10719);
or U10942 (N_10942,N_10651,N_10652);
xnor U10943 (N_10943,N_10648,N_10766);
and U10944 (N_10944,N_10653,N_10649);
xor U10945 (N_10945,N_10723,N_10712);
and U10946 (N_10946,N_10617,N_10669);
nor U10947 (N_10947,N_10757,N_10632);
xnor U10948 (N_10948,N_10604,N_10688);
or U10949 (N_10949,N_10767,N_10657);
and U10950 (N_10950,N_10711,N_10716);
nand U10951 (N_10951,N_10612,N_10615);
or U10952 (N_10952,N_10653,N_10660);
nand U10953 (N_10953,N_10665,N_10791);
xor U10954 (N_10954,N_10695,N_10787);
nand U10955 (N_10955,N_10641,N_10634);
xor U10956 (N_10956,N_10610,N_10630);
nand U10957 (N_10957,N_10651,N_10681);
nor U10958 (N_10958,N_10634,N_10741);
nand U10959 (N_10959,N_10756,N_10694);
nor U10960 (N_10960,N_10771,N_10686);
and U10961 (N_10961,N_10737,N_10732);
nor U10962 (N_10962,N_10623,N_10705);
xor U10963 (N_10963,N_10779,N_10615);
or U10964 (N_10964,N_10685,N_10774);
nand U10965 (N_10965,N_10636,N_10603);
nand U10966 (N_10966,N_10629,N_10764);
nand U10967 (N_10967,N_10604,N_10781);
xor U10968 (N_10968,N_10749,N_10623);
and U10969 (N_10969,N_10710,N_10750);
nor U10970 (N_10970,N_10642,N_10657);
or U10971 (N_10971,N_10730,N_10620);
and U10972 (N_10972,N_10637,N_10700);
nand U10973 (N_10973,N_10778,N_10634);
xnor U10974 (N_10974,N_10742,N_10651);
nand U10975 (N_10975,N_10616,N_10660);
or U10976 (N_10976,N_10653,N_10777);
and U10977 (N_10977,N_10758,N_10659);
nor U10978 (N_10978,N_10761,N_10726);
nor U10979 (N_10979,N_10652,N_10770);
nor U10980 (N_10980,N_10652,N_10754);
and U10981 (N_10981,N_10707,N_10790);
and U10982 (N_10982,N_10626,N_10787);
nand U10983 (N_10983,N_10613,N_10602);
nor U10984 (N_10984,N_10663,N_10606);
nor U10985 (N_10985,N_10624,N_10797);
or U10986 (N_10986,N_10702,N_10741);
nand U10987 (N_10987,N_10707,N_10785);
or U10988 (N_10988,N_10632,N_10675);
and U10989 (N_10989,N_10648,N_10629);
xor U10990 (N_10990,N_10727,N_10748);
or U10991 (N_10991,N_10715,N_10659);
nor U10992 (N_10992,N_10685,N_10777);
and U10993 (N_10993,N_10717,N_10666);
and U10994 (N_10994,N_10710,N_10722);
or U10995 (N_10995,N_10716,N_10634);
and U10996 (N_10996,N_10614,N_10745);
or U10997 (N_10997,N_10608,N_10633);
nor U10998 (N_10998,N_10793,N_10682);
nand U10999 (N_10999,N_10731,N_10639);
xor U11000 (N_11000,N_10856,N_10826);
or U11001 (N_11001,N_10984,N_10904);
nor U11002 (N_11002,N_10941,N_10897);
nor U11003 (N_11003,N_10968,N_10867);
and U11004 (N_11004,N_10926,N_10976);
or U11005 (N_11005,N_10900,N_10927);
and U11006 (N_11006,N_10969,N_10951);
or U11007 (N_11007,N_10866,N_10993);
nand U11008 (N_11008,N_10880,N_10874);
nor U11009 (N_11009,N_10872,N_10813);
xnor U11010 (N_11010,N_10978,N_10985);
and U11011 (N_11011,N_10935,N_10944);
nor U11012 (N_11012,N_10830,N_10922);
nand U11013 (N_11013,N_10939,N_10934);
nor U11014 (N_11014,N_10859,N_10977);
or U11015 (N_11015,N_10947,N_10851);
or U11016 (N_11016,N_10950,N_10848);
nor U11017 (N_11017,N_10907,N_10920);
and U11018 (N_11018,N_10917,N_10995);
or U11019 (N_11019,N_10852,N_10827);
or U11020 (N_11020,N_10801,N_10837);
and U11021 (N_11021,N_10955,N_10850);
nor U11022 (N_11022,N_10916,N_10835);
nand U11023 (N_11023,N_10975,N_10819);
and U11024 (N_11024,N_10967,N_10865);
or U11025 (N_11025,N_10890,N_10805);
nand U11026 (N_11026,N_10930,N_10943);
nand U11027 (N_11027,N_10909,N_10962);
nand U11028 (N_11028,N_10808,N_10949);
and U11029 (N_11029,N_10822,N_10844);
and U11030 (N_11030,N_10841,N_10855);
nand U11031 (N_11031,N_10946,N_10983);
and U11032 (N_11032,N_10936,N_10942);
and U11033 (N_11033,N_10845,N_10817);
and U11034 (N_11034,N_10986,N_10875);
nand U11035 (N_11035,N_10883,N_10901);
and U11036 (N_11036,N_10965,N_10931);
or U11037 (N_11037,N_10878,N_10997);
xor U11038 (N_11038,N_10903,N_10994);
nor U11039 (N_11039,N_10893,N_10840);
or U11040 (N_11040,N_10802,N_10892);
nor U11041 (N_11041,N_10823,N_10910);
or U11042 (N_11042,N_10873,N_10973);
nor U11043 (N_11043,N_10996,N_10990);
or U11044 (N_11044,N_10906,N_10863);
nor U11045 (N_11045,N_10843,N_10902);
nand U11046 (N_11046,N_10921,N_10891);
nor U11047 (N_11047,N_10895,N_10948);
nand U11048 (N_11048,N_10894,N_10957);
nand U11049 (N_11049,N_10882,N_10876);
nand U11050 (N_11050,N_10846,N_10924);
nand U11051 (N_11051,N_10989,N_10980);
xor U11052 (N_11052,N_10862,N_10963);
or U11053 (N_11053,N_10816,N_10858);
nor U11054 (N_11054,N_10871,N_10981);
and U11055 (N_11055,N_10861,N_10815);
and U11056 (N_11056,N_10982,N_10905);
or U11057 (N_11057,N_10864,N_10810);
nor U11058 (N_11058,N_10800,N_10914);
nor U11059 (N_11059,N_10869,N_10836);
and U11060 (N_11060,N_10825,N_10896);
or U11061 (N_11061,N_10821,N_10912);
nand U11062 (N_11062,N_10877,N_10829);
and U11063 (N_11063,N_10807,N_10834);
and U11064 (N_11064,N_10919,N_10960);
xor U11065 (N_11065,N_10913,N_10945);
or U11066 (N_11066,N_10887,N_10879);
and U11067 (N_11067,N_10959,N_10987);
xnor U11068 (N_11068,N_10838,N_10999);
nand U11069 (N_11069,N_10970,N_10979);
or U11070 (N_11070,N_10812,N_10886);
or U11071 (N_11071,N_10911,N_10958);
nor U11072 (N_11072,N_10888,N_10937);
nand U11073 (N_11073,N_10961,N_10933);
and U11074 (N_11074,N_10938,N_10899);
nor U11075 (N_11075,N_10828,N_10854);
nand U11076 (N_11076,N_10923,N_10940);
nand U11077 (N_11077,N_10842,N_10918);
or U11078 (N_11078,N_10908,N_10929);
nand U11079 (N_11079,N_10928,N_10972);
or U11080 (N_11080,N_10849,N_10925);
or U11081 (N_11081,N_10952,N_10814);
nand U11082 (N_11082,N_10806,N_10870);
and U11083 (N_11083,N_10832,N_10847);
nor U11084 (N_11084,N_10831,N_10833);
nand U11085 (N_11085,N_10998,N_10974);
or U11086 (N_11086,N_10992,N_10804);
xnor U11087 (N_11087,N_10956,N_10811);
and U11088 (N_11088,N_10809,N_10889);
nor U11089 (N_11089,N_10818,N_10971);
and U11090 (N_11090,N_10839,N_10953);
nand U11091 (N_11091,N_10860,N_10898);
nor U11092 (N_11092,N_10991,N_10881);
or U11093 (N_11093,N_10932,N_10884);
and U11094 (N_11094,N_10966,N_10820);
nand U11095 (N_11095,N_10857,N_10868);
and U11096 (N_11096,N_10964,N_10824);
nor U11097 (N_11097,N_10853,N_10885);
or U11098 (N_11098,N_10803,N_10954);
or U11099 (N_11099,N_10988,N_10915);
nand U11100 (N_11100,N_10924,N_10850);
or U11101 (N_11101,N_10883,N_10991);
nand U11102 (N_11102,N_10859,N_10891);
and U11103 (N_11103,N_10861,N_10920);
nand U11104 (N_11104,N_10969,N_10930);
nand U11105 (N_11105,N_10887,N_10852);
nor U11106 (N_11106,N_10958,N_10898);
nand U11107 (N_11107,N_10993,N_10944);
xor U11108 (N_11108,N_10872,N_10821);
and U11109 (N_11109,N_10914,N_10957);
or U11110 (N_11110,N_10913,N_10810);
or U11111 (N_11111,N_10852,N_10809);
nand U11112 (N_11112,N_10941,N_10955);
xor U11113 (N_11113,N_10846,N_10807);
or U11114 (N_11114,N_10856,N_10949);
or U11115 (N_11115,N_10984,N_10813);
and U11116 (N_11116,N_10966,N_10957);
nor U11117 (N_11117,N_10851,N_10922);
xnor U11118 (N_11118,N_10875,N_10922);
nor U11119 (N_11119,N_10908,N_10952);
nor U11120 (N_11120,N_10860,N_10844);
xnor U11121 (N_11121,N_10845,N_10807);
nand U11122 (N_11122,N_10953,N_10883);
or U11123 (N_11123,N_10845,N_10825);
or U11124 (N_11124,N_10988,N_10928);
nor U11125 (N_11125,N_10972,N_10806);
and U11126 (N_11126,N_10874,N_10890);
or U11127 (N_11127,N_10888,N_10927);
nor U11128 (N_11128,N_10844,N_10940);
or U11129 (N_11129,N_10898,N_10832);
or U11130 (N_11130,N_10801,N_10920);
and U11131 (N_11131,N_10997,N_10809);
nand U11132 (N_11132,N_10859,N_10974);
nand U11133 (N_11133,N_10825,N_10853);
and U11134 (N_11134,N_10892,N_10882);
nand U11135 (N_11135,N_10877,N_10849);
and U11136 (N_11136,N_10907,N_10813);
xnor U11137 (N_11137,N_10926,N_10951);
nand U11138 (N_11138,N_10880,N_10923);
and U11139 (N_11139,N_10967,N_10955);
and U11140 (N_11140,N_10810,N_10938);
or U11141 (N_11141,N_10969,N_10901);
or U11142 (N_11142,N_10847,N_10951);
and U11143 (N_11143,N_10860,N_10848);
nor U11144 (N_11144,N_10870,N_10829);
and U11145 (N_11145,N_10951,N_10965);
nor U11146 (N_11146,N_10961,N_10889);
and U11147 (N_11147,N_10840,N_10907);
nand U11148 (N_11148,N_10997,N_10803);
or U11149 (N_11149,N_10818,N_10871);
nand U11150 (N_11150,N_10960,N_10935);
nor U11151 (N_11151,N_10874,N_10940);
or U11152 (N_11152,N_10883,N_10825);
or U11153 (N_11153,N_10988,N_10967);
and U11154 (N_11154,N_10997,N_10826);
and U11155 (N_11155,N_10928,N_10863);
or U11156 (N_11156,N_10868,N_10844);
nor U11157 (N_11157,N_10932,N_10957);
or U11158 (N_11158,N_10832,N_10810);
or U11159 (N_11159,N_10827,N_10913);
nor U11160 (N_11160,N_10807,N_10968);
nand U11161 (N_11161,N_10916,N_10942);
nand U11162 (N_11162,N_10985,N_10938);
nor U11163 (N_11163,N_10897,N_10892);
xor U11164 (N_11164,N_10987,N_10860);
or U11165 (N_11165,N_10919,N_10916);
nand U11166 (N_11166,N_10833,N_10970);
nand U11167 (N_11167,N_10836,N_10963);
and U11168 (N_11168,N_10935,N_10886);
nand U11169 (N_11169,N_10802,N_10979);
or U11170 (N_11170,N_10826,N_10909);
and U11171 (N_11171,N_10855,N_10993);
nor U11172 (N_11172,N_10917,N_10902);
nand U11173 (N_11173,N_10980,N_10933);
and U11174 (N_11174,N_10929,N_10813);
nor U11175 (N_11175,N_10941,N_10893);
or U11176 (N_11176,N_10971,N_10941);
or U11177 (N_11177,N_10999,N_10937);
or U11178 (N_11178,N_10816,N_10887);
xor U11179 (N_11179,N_10856,N_10915);
and U11180 (N_11180,N_10901,N_10965);
nor U11181 (N_11181,N_10868,N_10992);
nand U11182 (N_11182,N_10861,N_10906);
and U11183 (N_11183,N_10886,N_10960);
nor U11184 (N_11184,N_10968,N_10844);
xnor U11185 (N_11185,N_10917,N_10898);
xnor U11186 (N_11186,N_10853,N_10824);
or U11187 (N_11187,N_10989,N_10829);
nor U11188 (N_11188,N_10873,N_10994);
and U11189 (N_11189,N_10955,N_10951);
nand U11190 (N_11190,N_10811,N_10922);
or U11191 (N_11191,N_10986,N_10924);
nand U11192 (N_11192,N_10827,N_10929);
nor U11193 (N_11193,N_10900,N_10996);
or U11194 (N_11194,N_10870,N_10927);
or U11195 (N_11195,N_10848,N_10887);
or U11196 (N_11196,N_10894,N_10855);
and U11197 (N_11197,N_10858,N_10861);
and U11198 (N_11198,N_10871,N_10884);
xnor U11199 (N_11199,N_10886,N_10880);
nand U11200 (N_11200,N_11142,N_11195);
xor U11201 (N_11201,N_11032,N_11073);
nand U11202 (N_11202,N_11038,N_11099);
xnor U11203 (N_11203,N_11008,N_11117);
or U11204 (N_11204,N_11051,N_11186);
and U11205 (N_11205,N_11034,N_11044);
or U11206 (N_11206,N_11130,N_11095);
or U11207 (N_11207,N_11190,N_11163);
or U11208 (N_11208,N_11052,N_11134);
or U11209 (N_11209,N_11193,N_11176);
nor U11210 (N_11210,N_11063,N_11159);
or U11211 (N_11211,N_11045,N_11167);
and U11212 (N_11212,N_11065,N_11165);
nand U11213 (N_11213,N_11067,N_11157);
and U11214 (N_11214,N_11000,N_11018);
xnor U11215 (N_11215,N_11006,N_11162);
xor U11216 (N_11216,N_11143,N_11055);
nor U11217 (N_11217,N_11048,N_11027);
or U11218 (N_11218,N_11182,N_11128);
xnor U11219 (N_11219,N_11087,N_11080);
and U11220 (N_11220,N_11039,N_11188);
xor U11221 (N_11221,N_11075,N_11156);
xor U11222 (N_11222,N_11185,N_11196);
and U11223 (N_11223,N_11140,N_11171);
nor U11224 (N_11224,N_11031,N_11060);
and U11225 (N_11225,N_11106,N_11124);
or U11226 (N_11226,N_11037,N_11041);
and U11227 (N_11227,N_11043,N_11197);
xor U11228 (N_11228,N_11126,N_11184);
nand U11229 (N_11229,N_11139,N_11105);
nand U11230 (N_11230,N_11078,N_11173);
or U11231 (N_11231,N_11169,N_11191);
or U11232 (N_11232,N_11179,N_11042);
nand U11233 (N_11233,N_11110,N_11172);
nand U11234 (N_11234,N_11146,N_11009);
nand U11235 (N_11235,N_11153,N_11181);
xnor U11236 (N_11236,N_11001,N_11144);
and U11237 (N_11237,N_11025,N_11118);
or U11238 (N_11238,N_11069,N_11115);
nand U11239 (N_11239,N_11109,N_11024);
nor U11240 (N_11240,N_11168,N_11022);
xor U11241 (N_11241,N_11108,N_11077);
and U11242 (N_11242,N_11189,N_11132);
nor U11243 (N_11243,N_11053,N_11135);
or U11244 (N_11244,N_11133,N_11033);
xor U11245 (N_11245,N_11129,N_11005);
nor U11246 (N_11246,N_11103,N_11097);
nor U11247 (N_11247,N_11056,N_11183);
or U11248 (N_11248,N_11054,N_11023);
and U11249 (N_11249,N_11068,N_11137);
or U11250 (N_11250,N_11064,N_11145);
nor U11251 (N_11251,N_11035,N_11199);
or U11252 (N_11252,N_11046,N_11026);
nor U11253 (N_11253,N_11158,N_11013);
and U11254 (N_11254,N_11076,N_11071);
xor U11255 (N_11255,N_11177,N_11072);
or U11256 (N_11256,N_11082,N_11058);
nor U11257 (N_11257,N_11094,N_11123);
nand U11258 (N_11258,N_11047,N_11125);
or U11259 (N_11259,N_11180,N_11114);
and U11260 (N_11260,N_11170,N_11020);
and U11261 (N_11261,N_11083,N_11017);
nand U11262 (N_11262,N_11113,N_11175);
or U11263 (N_11263,N_11015,N_11019);
or U11264 (N_11264,N_11007,N_11092);
nor U11265 (N_11265,N_11147,N_11002);
nor U11266 (N_11266,N_11174,N_11194);
and U11267 (N_11267,N_11122,N_11079);
xnor U11268 (N_11268,N_11119,N_11116);
nand U11269 (N_11269,N_11091,N_11011);
nand U11270 (N_11270,N_11003,N_11086);
nor U11271 (N_11271,N_11016,N_11059);
xnor U11272 (N_11272,N_11198,N_11049);
xnor U11273 (N_11273,N_11036,N_11166);
nand U11274 (N_11274,N_11155,N_11178);
or U11275 (N_11275,N_11107,N_11030);
nand U11276 (N_11276,N_11100,N_11062);
or U11277 (N_11277,N_11029,N_11161);
nand U11278 (N_11278,N_11120,N_11187);
nor U11279 (N_11279,N_11085,N_11012);
or U11280 (N_11280,N_11070,N_11096);
or U11281 (N_11281,N_11121,N_11112);
nand U11282 (N_11282,N_11160,N_11148);
nor U11283 (N_11283,N_11154,N_11104);
nand U11284 (N_11284,N_11040,N_11074);
xor U11285 (N_11285,N_11084,N_11150);
or U11286 (N_11286,N_11136,N_11152);
nor U11287 (N_11287,N_11066,N_11138);
or U11288 (N_11288,N_11098,N_11149);
xnor U11289 (N_11289,N_11004,N_11102);
xor U11290 (N_11290,N_11057,N_11061);
nand U11291 (N_11291,N_11141,N_11014);
nor U11292 (N_11292,N_11101,N_11050);
nor U11293 (N_11293,N_11028,N_11151);
nand U11294 (N_11294,N_11192,N_11088);
nand U11295 (N_11295,N_11131,N_11089);
and U11296 (N_11296,N_11090,N_11093);
nand U11297 (N_11297,N_11081,N_11111);
nor U11298 (N_11298,N_11127,N_11021);
nor U11299 (N_11299,N_11164,N_11010);
or U11300 (N_11300,N_11134,N_11137);
and U11301 (N_11301,N_11085,N_11176);
and U11302 (N_11302,N_11100,N_11032);
and U11303 (N_11303,N_11038,N_11171);
or U11304 (N_11304,N_11041,N_11142);
nand U11305 (N_11305,N_11183,N_11153);
nor U11306 (N_11306,N_11020,N_11143);
and U11307 (N_11307,N_11141,N_11137);
nor U11308 (N_11308,N_11025,N_11013);
or U11309 (N_11309,N_11042,N_11168);
nor U11310 (N_11310,N_11126,N_11099);
nor U11311 (N_11311,N_11135,N_11072);
nand U11312 (N_11312,N_11047,N_11096);
nand U11313 (N_11313,N_11101,N_11123);
and U11314 (N_11314,N_11158,N_11101);
and U11315 (N_11315,N_11065,N_11028);
or U11316 (N_11316,N_11124,N_11119);
xnor U11317 (N_11317,N_11152,N_11003);
or U11318 (N_11318,N_11005,N_11035);
nand U11319 (N_11319,N_11026,N_11151);
nand U11320 (N_11320,N_11180,N_11035);
and U11321 (N_11321,N_11039,N_11007);
and U11322 (N_11322,N_11177,N_11076);
or U11323 (N_11323,N_11190,N_11037);
nand U11324 (N_11324,N_11027,N_11132);
or U11325 (N_11325,N_11003,N_11051);
nor U11326 (N_11326,N_11171,N_11199);
nand U11327 (N_11327,N_11004,N_11002);
and U11328 (N_11328,N_11090,N_11050);
xor U11329 (N_11329,N_11026,N_11139);
nor U11330 (N_11330,N_11179,N_11016);
nand U11331 (N_11331,N_11181,N_11042);
nor U11332 (N_11332,N_11069,N_11043);
nand U11333 (N_11333,N_11089,N_11008);
nor U11334 (N_11334,N_11087,N_11073);
nor U11335 (N_11335,N_11154,N_11192);
nand U11336 (N_11336,N_11163,N_11082);
nand U11337 (N_11337,N_11188,N_11182);
or U11338 (N_11338,N_11024,N_11110);
and U11339 (N_11339,N_11043,N_11189);
or U11340 (N_11340,N_11106,N_11052);
nor U11341 (N_11341,N_11037,N_11022);
or U11342 (N_11342,N_11087,N_11054);
or U11343 (N_11343,N_11028,N_11000);
nand U11344 (N_11344,N_11193,N_11149);
nor U11345 (N_11345,N_11108,N_11138);
or U11346 (N_11346,N_11191,N_11106);
or U11347 (N_11347,N_11099,N_11042);
or U11348 (N_11348,N_11069,N_11073);
nand U11349 (N_11349,N_11067,N_11141);
or U11350 (N_11350,N_11176,N_11104);
xnor U11351 (N_11351,N_11057,N_11099);
and U11352 (N_11352,N_11179,N_11183);
xor U11353 (N_11353,N_11088,N_11118);
nor U11354 (N_11354,N_11046,N_11023);
nand U11355 (N_11355,N_11033,N_11125);
and U11356 (N_11356,N_11153,N_11103);
xnor U11357 (N_11357,N_11019,N_11052);
nand U11358 (N_11358,N_11104,N_11135);
nor U11359 (N_11359,N_11172,N_11145);
xnor U11360 (N_11360,N_11020,N_11026);
nand U11361 (N_11361,N_11164,N_11181);
nor U11362 (N_11362,N_11061,N_11146);
nor U11363 (N_11363,N_11153,N_11117);
nand U11364 (N_11364,N_11049,N_11024);
xor U11365 (N_11365,N_11199,N_11111);
nand U11366 (N_11366,N_11115,N_11141);
nand U11367 (N_11367,N_11080,N_11033);
nor U11368 (N_11368,N_11033,N_11102);
nand U11369 (N_11369,N_11105,N_11189);
and U11370 (N_11370,N_11033,N_11191);
and U11371 (N_11371,N_11086,N_11184);
or U11372 (N_11372,N_11064,N_11177);
nand U11373 (N_11373,N_11022,N_11097);
and U11374 (N_11374,N_11144,N_11013);
nor U11375 (N_11375,N_11186,N_11071);
nor U11376 (N_11376,N_11067,N_11182);
and U11377 (N_11377,N_11113,N_11116);
nand U11378 (N_11378,N_11174,N_11056);
and U11379 (N_11379,N_11011,N_11121);
or U11380 (N_11380,N_11151,N_11183);
nor U11381 (N_11381,N_11169,N_11188);
nand U11382 (N_11382,N_11196,N_11162);
nand U11383 (N_11383,N_11131,N_11087);
or U11384 (N_11384,N_11128,N_11076);
or U11385 (N_11385,N_11104,N_11121);
and U11386 (N_11386,N_11000,N_11152);
or U11387 (N_11387,N_11145,N_11027);
nand U11388 (N_11388,N_11134,N_11155);
or U11389 (N_11389,N_11181,N_11159);
xor U11390 (N_11390,N_11026,N_11149);
nor U11391 (N_11391,N_11055,N_11111);
xor U11392 (N_11392,N_11004,N_11194);
and U11393 (N_11393,N_11008,N_11052);
or U11394 (N_11394,N_11050,N_11133);
or U11395 (N_11395,N_11124,N_11127);
nand U11396 (N_11396,N_11115,N_11098);
nor U11397 (N_11397,N_11183,N_11143);
and U11398 (N_11398,N_11010,N_11134);
or U11399 (N_11399,N_11199,N_11183);
nand U11400 (N_11400,N_11294,N_11209);
xnor U11401 (N_11401,N_11311,N_11369);
nor U11402 (N_11402,N_11212,N_11367);
nor U11403 (N_11403,N_11360,N_11343);
and U11404 (N_11404,N_11250,N_11393);
or U11405 (N_11405,N_11264,N_11262);
and U11406 (N_11406,N_11266,N_11247);
nor U11407 (N_11407,N_11399,N_11340);
nor U11408 (N_11408,N_11238,N_11361);
and U11409 (N_11409,N_11297,N_11332);
nand U11410 (N_11410,N_11253,N_11259);
and U11411 (N_11411,N_11375,N_11338);
or U11412 (N_11412,N_11215,N_11208);
or U11413 (N_11413,N_11305,N_11252);
nor U11414 (N_11414,N_11378,N_11346);
or U11415 (N_11415,N_11279,N_11224);
or U11416 (N_11416,N_11239,N_11296);
and U11417 (N_11417,N_11372,N_11363);
and U11418 (N_11418,N_11366,N_11324);
or U11419 (N_11419,N_11321,N_11287);
or U11420 (N_11420,N_11202,N_11293);
xnor U11421 (N_11421,N_11274,N_11267);
and U11422 (N_11422,N_11258,N_11242);
nand U11423 (N_11423,N_11398,N_11244);
or U11424 (N_11424,N_11211,N_11391);
nand U11425 (N_11425,N_11243,N_11235);
and U11426 (N_11426,N_11320,N_11381);
nor U11427 (N_11427,N_11308,N_11268);
nand U11428 (N_11428,N_11388,N_11335);
or U11429 (N_11429,N_11248,N_11219);
nor U11430 (N_11430,N_11336,N_11263);
nor U11431 (N_11431,N_11328,N_11218);
or U11432 (N_11432,N_11387,N_11384);
nand U11433 (N_11433,N_11281,N_11379);
or U11434 (N_11434,N_11396,N_11260);
xor U11435 (N_11435,N_11233,N_11241);
xor U11436 (N_11436,N_11226,N_11350);
nor U11437 (N_11437,N_11345,N_11344);
and U11438 (N_11438,N_11280,N_11323);
and U11439 (N_11439,N_11327,N_11245);
or U11440 (N_11440,N_11277,N_11236);
and U11441 (N_11441,N_11374,N_11357);
nor U11442 (N_11442,N_11213,N_11255);
and U11443 (N_11443,N_11307,N_11394);
or U11444 (N_11444,N_11317,N_11225);
nor U11445 (N_11445,N_11330,N_11214);
or U11446 (N_11446,N_11256,N_11355);
or U11447 (N_11447,N_11397,N_11284);
xor U11448 (N_11448,N_11298,N_11356);
xor U11449 (N_11449,N_11318,N_11276);
nor U11450 (N_11450,N_11333,N_11270);
or U11451 (N_11451,N_11354,N_11295);
or U11452 (N_11452,N_11269,N_11373);
or U11453 (N_11453,N_11313,N_11288);
nand U11454 (N_11454,N_11392,N_11286);
nand U11455 (N_11455,N_11207,N_11231);
nand U11456 (N_11456,N_11386,N_11221);
nand U11457 (N_11457,N_11303,N_11201);
and U11458 (N_11458,N_11364,N_11319);
or U11459 (N_11459,N_11203,N_11230);
nor U11460 (N_11460,N_11223,N_11380);
and U11461 (N_11461,N_11275,N_11206);
nand U11462 (N_11462,N_11358,N_11261);
nand U11463 (N_11463,N_11389,N_11342);
or U11464 (N_11464,N_11217,N_11227);
nand U11465 (N_11465,N_11368,N_11222);
and U11466 (N_11466,N_11301,N_11290);
xor U11467 (N_11467,N_11246,N_11334);
or U11468 (N_11468,N_11383,N_11370);
and U11469 (N_11469,N_11265,N_11272);
or U11470 (N_11470,N_11309,N_11302);
nor U11471 (N_11471,N_11306,N_11310);
and U11472 (N_11472,N_11341,N_11339);
xnor U11473 (N_11473,N_11312,N_11292);
xnor U11474 (N_11474,N_11316,N_11337);
xnor U11475 (N_11475,N_11395,N_11348);
or U11476 (N_11476,N_11200,N_11362);
nor U11477 (N_11477,N_11314,N_11220);
and U11478 (N_11478,N_11237,N_11390);
and U11479 (N_11479,N_11347,N_11216);
nor U11480 (N_11480,N_11285,N_11249);
xor U11481 (N_11481,N_11353,N_11359);
nand U11482 (N_11482,N_11322,N_11352);
and U11483 (N_11483,N_11365,N_11205);
nand U11484 (N_11484,N_11385,N_11382);
nor U11485 (N_11485,N_11251,N_11254);
nor U11486 (N_11486,N_11315,N_11351);
nand U11487 (N_11487,N_11257,N_11329);
xnor U11488 (N_11488,N_11331,N_11278);
nand U11489 (N_11489,N_11376,N_11349);
nor U11490 (N_11490,N_11377,N_11325);
and U11491 (N_11491,N_11229,N_11234);
nand U11492 (N_11492,N_11289,N_11371);
nor U11493 (N_11493,N_11204,N_11299);
and U11494 (N_11494,N_11240,N_11232);
or U11495 (N_11495,N_11283,N_11304);
xor U11496 (N_11496,N_11300,N_11273);
nor U11497 (N_11497,N_11282,N_11271);
nor U11498 (N_11498,N_11291,N_11326);
or U11499 (N_11499,N_11228,N_11210);
xor U11500 (N_11500,N_11385,N_11246);
and U11501 (N_11501,N_11253,N_11260);
nor U11502 (N_11502,N_11313,N_11226);
and U11503 (N_11503,N_11360,N_11244);
and U11504 (N_11504,N_11350,N_11384);
and U11505 (N_11505,N_11317,N_11208);
and U11506 (N_11506,N_11373,N_11200);
nand U11507 (N_11507,N_11287,N_11361);
and U11508 (N_11508,N_11318,N_11292);
or U11509 (N_11509,N_11314,N_11346);
or U11510 (N_11510,N_11348,N_11225);
xor U11511 (N_11511,N_11380,N_11343);
and U11512 (N_11512,N_11371,N_11336);
and U11513 (N_11513,N_11298,N_11250);
or U11514 (N_11514,N_11266,N_11376);
nand U11515 (N_11515,N_11397,N_11277);
nor U11516 (N_11516,N_11356,N_11368);
or U11517 (N_11517,N_11280,N_11202);
nor U11518 (N_11518,N_11279,N_11374);
or U11519 (N_11519,N_11348,N_11221);
and U11520 (N_11520,N_11296,N_11382);
nand U11521 (N_11521,N_11316,N_11259);
or U11522 (N_11522,N_11223,N_11262);
nand U11523 (N_11523,N_11326,N_11296);
nor U11524 (N_11524,N_11255,N_11236);
and U11525 (N_11525,N_11390,N_11394);
nand U11526 (N_11526,N_11315,N_11395);
nor U11527 (N_11527,N_11250,N_11316);
nand U11528 (N_11528,N_11353,N_11387);
or U11529 (N_11529,N_11257,N_11215);
nor U11530 (N_11530,N_11334,N_11228);
and U11531 (N_11531,N_11391,N_11359);
or U11532 (N_11532,N_11331,N_11328);
and U11533 (N_11533,N_11249,N_11271);
or U11534 (N_11534,N_11240,N_11325);
or U11535 (N_11535,N_11275,N_11339);
nand U11536 (N_11536,N_11325,N_11261);
and U11537 (N_11537,N_11329,N_11214);
or U11538 (N_11538,N_11396,N_11264);
nand U11539 (N_11539,N_11344,N_11326);
and U11540 (N_11540,N_11352,N_11382);
or U11541 (N_11541,N_11393,N_11208);
nand U11542 (N_11542,N_11358,N_11259);
nor U11543 (N_11543,N_11241,N_11287);
nor U11544 (N_11544,N_11261,N_11296);
nand U11545 (N_11545,N_11294,N_11371);
and U11546 (N_11546,N_11237,N_11371);
and U11547 (N_11547,N_11350,N_11396);
nor U11548 (N_11548,N_11347,N_11205);
and U11549 (N_11549,N_11247,N_11282);
nand U11550 (N_11550,N_11212,N_11369);
nor U11551 (N_11551,N_11345,N_11207);
and U11552 (N_11552,N_11252,N_11213);
nor U11553 (N_11553,N_11276,N_11225);
and U11554 (N_11554,N_11266,N_11391);
and U11555 (N_11555,N_11375,N_11385);
nor U11556 (N_11556,N_11275,N_11250);
and U11557 (N_11557,N_11216,N_11337);
nand U11558 (N_11558,N_11262,N_11253);
and U11559 (N_11559,N_11262,N_11315);
or U11560 (N_11560,N_11292,N_11393);
or U11561 (N_11561,N_11326,N_11270);
and U11562 (N_11562,N_11282,N_11237);
or U11563 (N_11563,N_11306,N_11366);
or U11564 (N_11564,N_11347,N_11331);
nor U11565 (N_11565,N_11232,N_11265);
nand U11566 (N_11566,N_11337,N_11378);
nand U11567 (N_11567,N_11211,N_11252);
nand U11568 (N_11568,N_11296,N_11330);
or U11569 (N_11569,N_11391,N_11298);
or U11570 (N_11570,N_11244,N_11269);
and U11571 (N_11571,N_11213,N_11309);
or U11572 (N_11572,N_11361,N_11351);
nand U11573 (N_11573,N_11329,N_11305);
or U11574 (N_11574,N_11310,N_11276);
nor U11575 (N_11575,N_11338,N_11263);
nand U11576 (N_11576,N_11393,N_11321);
nand U11577 (N_11577,N_11331,N_11234);
nand U11578 (N_11578,N_11339,N_11289);
and U11579 (N_11579,N_11208,N_11307);
nor U11580 (N_11580,N_11252,N_11261);
xor U11581 (N_11581,N_11284,N_11262);
and U11582 (N_11582,N_11293,N_11378);
nor U11583 (N_11583,N_11334,N_11279);
nor U11584 (N_11584,N_11248,N_11213);
nor U11585 (N_11585,N_11264,N_11398);
or U11586 (N_11586,N_11326,N_11266);
or U11587 (N_11587,N_11223,N_11233);
nor U11588 (N_11588,N_11366,N_11248);
or U11589 (N_11589,N_11355,N_11230);
and U11590 (N_11590,N_11247,N_11321);
nor U11591 (N_11591,N_11281,N_11341);
and U11592 (N_11592,N_11383,N_11228);
and U11593 (N_11593,N_11305,N_11253);
nor U11594 (N_11594,N_11290,N_11359);
nor U11595 (N_11595,N_11384,N_11263);
xnor U11596 (N_11596,N_11349,N_11211);
nor U11597 (N_11597,N_11318,N_11213);
and U11598 (N_11598,N_11385,N_11244);
xor U11599 (N_11599,N_11248,N_11369);
xor U11600 (N_11600,N_11534,N_11434);
nand U11601 (N_11601,N_11527,N_11404);
nand U11602 (N_11602,N_11448,N_11403);
or U11603 (N_11603,N_11426,N_11455);
and U11604 (N_11604,N_11595,N_11485);
and U11605 (N_11605,N_11511,N_11585);
nor U11606 (N_11606,N_11552,N_11532);
or U11607 (N_11607,N_11437,N_11420);
or U11608 (N_11608,N_11576,N_11423);
nand U11609 (N_11609,N_11590,N_11495);
or U11610 (N_11610,N_11531,N_11407);
nor U11611 (N_11611,N_11571,N_11451);
xor U11612 (N_11612,N_11529,N_11476);
and U11613 (N_11613,N_11596,N_11486);
nor U11614 (N_11614,N_11543,N_11540);
or U11615 (N_11615,N_11414,N_11447);
nor U11616 (N_11616,N_11450,N_11412);
nand U11617 (N_11617,N_11424,N_11578);
nand U11618 (N_11618,N_11598,N_11453);
nor U11619 (N_11619,N_11435,N_11508);
nor U11620 (N_11620,N_11494,N_11583);
and U11621 (N_11621,N_11521,N_11402);
or U11622 (N_11622,N_11557,N_11410);
nand U11623 (N_11623,N_11483,N_11409);
nor U11624 (N_11624,N_11489,N_11575);
nand U11625 (N_11625,N_11501,N_11482);
nand U11626 (N_11626,N_11528,N_11425);
and U11627 (N_11627,N_11471,N_11572);
nand U11628 (N_11628,N_11490,N_11523);
or U11629 (N_11629,N_11481,N_11497);
or U11630 (N_11630,N_11454,N_11446);
and U11631 (N_11631,N_11550,N_11445);
and U11632 (N_11632,N_11522,N_11473);
or U11633 (N_11633,N_11415,N_11460);
or U11634 (N_11634,N_11584,N_11456);
nand U11635 (N_11635,N_11479,N_11480);
and U11636 (N_11636,N_11477,N_11568);
nand U11637 (N_11637,N_11440,N_11505);
or U11638 (N_11638,N_11565,N_11589);
or U11639 (N_11639,N_11563,N_11520);
nand U11640 (N_11640,N_11530,N_11566);
nor U11641 (N_11641,N_11587,N_11558);
and U11642 (N_11642,N_11555,N_11496);
or U11643 (N_11643,N_11500,N_11549);
or U11644 (N_11644,N_11551,N_11444);
nand U11645 (N_11645,N_11561,N_11400);
xor U11646 (N_11646,N_11577,N_11449);
nor U11647 (N_11647,N_11567,N_11544);
and U11648 (N_11648,N_11436,N_11488);
nor U11649 (N_11649,N_11417,N_11581);
or U11650 (N_11650,N_11533,N_11580);
nor U11651 (N_11651,N_11510,N_11433);
or U11652 (N_11652,N_11452,N_11470);
xnor U11653 (N_11653,N_11457,N_11512);
and U11654 (N_11654,N_11594,N_11487);
nor U11655 (N_11655,N_11579,N_11593);
or U11656 (N_11656,N_11562,N_11465);
xor U11657 (N_11657,N_11504,N_11492);
nor U11658 (N_11658,N_11411,N_11459);
or U11659 (N_11659,N_11443,N_11597);
or U11660 (N_11660,N_11439,N_11537);
xnor U11661 (N_11661,N_11401,N_11545);
nand U11662 (N_11662,N_11462,N_11586);
nor U11663 (N_11663,N_11467,N_11428);
and U11664 (N_11664,N_11484,N_11431);
and U11665 (N_11665,N_11466,N_11542);
nand U11666 (N_11666,N_11419,N_11556);
nor U11667 (N_11667,N_11502,N_11475);
and U11668 (N_11668,N_11503,N_11499);
xor U11669 (N_11669,N_11441,N_11588);
xnor U11670 (N_11670,N_11559,N_11599);
nand U11671 (N_11671,N_11413,N_11461);
and U11672 (N_11672,N_11546,N_11422);
or U11673 (N_11673,N_11516,N_11574);
nand U11674 (N_11674,N_11570,N_11514);
nor U11675 (N_11675,N_11469,N_11582);
xnor U11676 (N_11676,N_11538,N_11541);
or U11677 (N_11677,N_11432,N_11519);
and U11678 (N_11678,N_11464,N_11408);
nor U11679 (N_11679,N_11526,N_11554);
nor U11680 (N_11680,N_11468,N_11569);
xnor U11681 (N_11681,N_11573,N_11458);
nor U11682 (N_11682,N_11405,N_11474);
nand U11683 (N_11683,N_11463,N_11524);
or U11684 (N_11684,N_11498,N_11547);
and U11685 (N_11685,N_11513,N_11518);
nand U11686 (N_11686,N_11416,N_11553);
nor U11687 (N_11687,N_11427,N_11430);
and U11688 (N_11688,N_11591,N_11535);
xor U11689 (N_11689,N_11418,N_11491);
or U11690 (N_11690,N_11506,N_11525);
nor U11691 (N_11691,N_11517,N_11406);
or U11692 (N_11692,N_11438,N_11421);
xnor U11693 (N_11693,N_11548,N_11564);
and U11694 (N_11694,N_11560,N_11429);
nand U11695 (N_11695,N_11509,N_11478);
xnor U11696 (N_11696,N_11592,N_11472);
nor U11697 (N_11697,N_11515,N_11442);
nor U11698 (N_11698,N_11539,N_11507);
nand U11699 (N_11699,N_11536,N_11493);
nor U11700 (N_11700,N_11555,N_11549);
and U11701 (N_11701,N_11472,N_11561);
nand U11702 (N_11702,N_11552,N_11480);
xor U11703 (N_11703,N_11468,N_11546);
or U11704 (N_11704,N_11464,N_11581);
nor U11705 (N_11705,N_11482,N_11440);
or U11706 (N_11706,N_11488,N_11465);
or U11707 (N_11707,N_11530,N_11469);
and U11708 (N_11708,N_11555,N_11444);
and U11709 (N_11709,N_11481,N_11546);
nor U11710 (N_11710,N_11557,N_11453);
and U11711 (N_11711,N_11501,N_11568);
or U11712 (N_11712,N_11555,N_11558);
and U11713 (N_11713,N_11480,N_11471);
and U11714 (N_11714,N_11470,N_11459);
or U11715 (N_11715,N_11460,N_11579);
or U11716 (N_11716,N_11573,N_11596);
or U11717 (N_11717,N_11500,N_11402);
or U11718 (N_11718,N_11515,N_11423);
nand U11719 (N_11719,N_11566,N_11477);
and U11720 (N_11720,N_11417,N_11473);
and U11721 (N_11721,N_11540,N_11442);
nand U11722 (N_11722,N_11419,N_11529);
xor U11723 (N_11723,N_11483,N_11459);
or U11724 (N_11724,N_11549,N_11431);
nor U11725 (N_11725,N_11498,N_11528);
xor U11726 (N_11726,N_11590,N_11415);
nor U11727 (N_11727,N_11459,N_11474);
or U11728 (N_11728,N_11524,N_11455);
or U11729 (N_11729,N_11520,N_11439);
nand U11730 (N_11730,N_11502,N_11526);
and U11731 (N_11731,N_11496,N_11474);
nand U11732 (N_11732,N_11527,N_11506);
nor U11733 (N_11733,N_11448,N_11573);
and U11734 (N_11734,N_11469,N_11493);
or U11735 (N_11735,N_11541,N_11416);
or U11736 (N_11736,N_11416,N_11577);
and U11737 (N_11737,N_11565,N_11496);
and U11738 (N_11738,N_11566,N_11433);
or U11739 (N_11739,N_11458,N_11528);
and U11740 (N_11740,N_11497,N_11427);
xor U11741 (N_11741,N_11512,N_11598);
or U11742 (N_11742,N_11583,N_11516);
or U11743 (N_11743,N_11554,N_11424);
and U11744 (N_11744,N_11427,N_11460);
and U11745 (N_11745,N_11591,N_11586);
and U11746 (N_11746,N_11513,N_11546);
xor U11747 (N_11747,N_11497,N_11466);
or U11748 (N_11748,N_11542,N_11581);
or U11749 (N_11749,N_11450,N_11551);
and U11750 (N_11750,N_11599,N_11577);
xor U11751 (N_11751,N_11484,N_11421);
and U11752 (N_11752,N_11547,N_11497);
nand U11753 (N_11753,N_11583,N_11570);
or U11754 (N_11754,N_11554,N_11558);
xor U11755 (N_11755,N_11485,N_11566);
or U11756 (N_11756,N_11491,N_11471);
or U11757 (N_11757,N_11428,N_11411);
and U11758 (N_11758,N_11503,N_11556);
or U11759 (N_11759,N_11523,N_11572);
nor U11760 (N_11760,N_11549,N_11595);
nand U11761 (N_11761,N_11545,N_11420);
and U11762 (N_11762,N_11458,N_11560);
and U11763 (N_11763,N_11578,N_11594);
or U11764 (N_11764,N_11418,N_11549);
or U11765 (N_11765,N_11578,N_11410);
or U11766 (N_11766,N_11574,N_11440);
and U11767 (N_11767,N_11501,N_11444);
and U11768 (N_11768,N_11559,N_11458);
or U11769 (N_11769,N_11493,N_11591);
nor U11770 (N_11770,N_11493,N_11511);
nand U11771 (N_11771,N_11481,N_11545);
and U11772 (N_11772,N_11564,N_11419);
or U11773 (N_11773,N_11469,N_11417);
nor U11774 (N_11774,N_11551,N_11553);
nand U11775 (N_11775,N_11464,N_11587);
or U11776 (N_11776,N_11549,N_11514);
nor U11777 (N_11777,N_11540,N_11502);
or U11778 (N_11778,N_11580,N_11535);
or U11779 (N_11779,N_11472,N_11481);
xor U11780 (N_11780,N_11464,N_11599);
or U11781 (N_11781,N_11461,N_11537);
and U11782 (N_11782,N_11419,N_11537);
or U11783 (N_11783,N_11506,N_11547);
xor U11784 (N_11784,N_11557,N_11531);
nor U11785 (N_11785,N_11505,N_11400);
xor U11786 (N_11786,N_11506,N_11499);
nand U11787 (N_11787,N_11471,N_11487);
and U11788 (N_11788,N_11435,N_11568);
or U11789 (N_11789,N_11464,N_11531);
or U11790 (N_11790,N_11599,N_11590);
xor U11791 (N_11791,N_11473,N_11496);
and U11792 (N_11792,N_11482,N_11432);
nor U11793 (N_11793,N_11485,N_11511);
or U11794 (N_11794,N_11538,N_11571);
and U11795 (N_11795,N_11533,N_11571);
and U11796 (N_11796,N_11420,N_11483);
and U11797 (N_11797,N_11542,N_11463);
xnor U11798 (N_11798,N_11417,N_11423);
xor U11799 (N_11799,N_11451,N_11461);
or U11800 (N_11800,N_11795,N_11622);
or U11801 (N_11801,N_11608,N_11626);
and U11802 (N_11802,N_11620,N_11659);
or U11803 (N_11803,N_11640,N_11733);
or U11804 (N_11804,N_11706,N_11782);
nand U11805 (N_11805,N_11762,N_11704);
nand U11806 (N_11806,N_11787,N_11628);
nor U11807 (N_11807,N_11788,N_11666);
xnor U11808 (N_11808,N_11764,N_11645);
nor U11809 (N_11809,N_11636,N_11698);
nor U11810 (N_11810,N_11778,N_11798);
or U11811 (N_11811,N_11703,N_11618);
and U11812 (N_11812,N_11757,N_11669);
nor U11813 (N_11813,N_11665,N_11758);
or U11814 (N_11814,N_11710,N_11724);
nand U11815 (N_11815,N_11716,N_11745);
nand U11816 (N_11816,N_11775,N_11797);
and U11817 (N_11817,N_11756,N_11684);
nor U11818 (N_11818,N_11779,N_11751);
nand U11819 (N_11819,N_11726,N_11654);
nor U11820 (N_11820,N_11789,N_11790);
or U11821 (N_11821,N_11765,N_11613);
nor U11822 (N_11822,N_11708,N_11721);
xnor U11823 (N_11823,N_11695,N_11760);
nand U11824 (N_11824,N_11784,N_11794);
and U11825 (N_11825,N_11754,N_11651);
nand U11826 (N_11826,N_11799,N_11689);
nor U11827 (N_11827,N_11650,N_11639);
or U11828 (N_11828,N_11702,N_11773);
or U11829 (N_11829,N_11786,N_11648);
or U11830 (N_11830,N_11612,N_11673);
nor U11831 (N_11831,N_11675,N_11731);
xor U11832 (N_11832,N_11683,N_11619);
or U11833 (N_11833,N_11727,N_11667);
or U11834 (N_11834,N_11652,N_11714);
nor U11835 (N_11835,N_11709,N_11769);
and U11836 (N_11836,N_11723,N_11615);
nand U11837 (N_11837,N_11604,N_11602);
or U11838 (N_11838,N_11725,N_11771);
and U11839 (N_11839,N_11658,N_11693);
nor U11840 (N_11840,N_11629,N_11768);
nand U11841 (N_11841,N_11774,N_11661);
nand U11842 (N_11842,N_11711,N_11780);
or U11843 (N_11843,N_11627,N_11719);
or U11844 (N_11844,N_11690,N_11718);
and U11845 (N_11845,N_11749,N_11776);
nand U11846 (N_11846,N_11647,N_11793);
nand U11847 (N_11847,N_11777,N_11740);
or U11848 (N_11848,N_11696,N_11672);
nand U11849 (N_11849,N_11717,N_11734);
nor U11850 (N_11850,N_11638,N_11720);
nand U11851 (N_11851,N_11748,N_11692);
nor U11852 (N_11852,N_11635,N_11722);
or U11853 (N_11853,N_11741,N_11678);
nor U11854 (N_11854,N_11633,N_11701);
or U11855 (N_11855,N_11713,N_11674);
xor U11856 (N_11856,N_11770,N_11603);
and U11857 (N_11857,N_11670,N_11705);
nand U11858 (N_11858,N_11697,N_11796);
nor U11859 (N_11859,N_11737,N_11655);
or U11860 (N_11860,N_11643,N_11671);
and U11861 (N_11861,N_11606,N_11792);
and U11862 (N_11862,N_11759,N_11766);
and U11863 (N_11863,N_11657,N_11767);
nor U11864 (N_11864,N_11610,N_11663);
nand U11865 (N_11865,N_11712,N_11682);
or U11866 (N_11866,N_11742,N_11743);
nand U11867 (N_11867,N_11746,N_11681);
nor U11868 (N_11868,N_11614,N_11644);
nor U11869 (N_11869,N_11611,N_11755);
or U11870 (N_11870,N_11616,N_11607);
nand U11871 (N_11871,N_11686,N_11730);
nand U11872 (N_11872,N_11634,N_11738);
xor U11873 (N_11873,N_11783,N_11600);
and U11874 (N_11874,N_11676,N_11617);
nor U11875 (N_11875,N_11700,N_11752);
nor U11876 (N_11876,N_11699,N_11688);
and U11877 (N_11877,N_11668,N_11631);
and U11878 (N_11878,N_11642,N_11624);
nand U11879 (N_11879,N_11736,N_11656);
nand U11880 (N_11880,N_11653,N_11729);
nand U11881 (N_11881,N_11785,N_11625);
nand U11882 (N_11882,N_11687,N_11735);
and U11883 (N_11883,N_11691,N_11739);
nand U11884 (N_11884,N_11632,N_11750);
xnor U11885 (N_11885,N_11662,N_11623);
or U11886 (N_11886,N_11791,N_11744);
nand U11887 (N_11887,N_11664,N_11772);
nand U11888 (N_11888,N_11753,N_11646);
xor U11889 (N_11889,N_11601,N_11732);
or U11890 (N_11890,N_11660,N_11685);
nand U11891 (N_11891,N_11677,N_11763);
nand U11892 (N_11892,N_11649,N_11680);
or U11893 (N_11893,N_11707,N_11679);
and U11894 (N_11894,N_11781,N_11621);
xor U11895 (N_11895,N_11609,N_11605);
and U11896 (N_11896,N_11728,N_11630);
nor U11897 (N_11897,N_11694,N_11761);
or U11898 (N_11898,N_11641,N_11715);
nand U11899 (N_11899,N_11637,N_11747);
or U11900 (N_11900,N_11670,N_11791);
nor U11901 (N_11901,N_11653,N_11636);
or U11902 (N_11902,N_11766,N_11731);
and U11903 (N_11903,N_11646,N_11620);
and U11904 (N_11904,N_11672,N_11728);
and U11905 (N_11905,N_11697,N_11729);
nor U11906 (N_11906,N_11697,N_11630);
nand U11907 (N_11907,N_11660,N_11677);
nand U11908 (N_11908,N_11785,N_11787);
nor U11909 (N_11909,N_11727,N_11674);
nor U11910 (N_11910,N_11696,N_11717);
and U11911 (N_11911,N_11682,N_11612);
and U11912 (N_11912,N_11683,N_11794);
nor U11913 (N_11913,N_11625,N_11600);
or U11914 (N_11914,N_11620,N_11681);
or U11915 (N_11915,N_11675,N_11649);
nor U11916 (N_11916,N_11766,N_11768);
and U11917 (N_11917,N_11666,N_11725);
nor U11918 (N_11918,N_11741,N_11708);
or U11919 (N_11919,N_11746,N_11718);
nor U11920 (N_11920,N_11751,N_11797);
nor U11921 (N_11921,N_11740,N_11774);
nand U11922 (N_11922,N_11702,N_11639);
nor U11923 (N_11923,N_11721,N_11710);
nor U11924 (N_11924,N_11626,N_11600);
and U11925 (N_11925,N_11671,N_11725);
nor U11926 (N_11926,N_11601,N_11605);
nor U11927 (N_11927,N_11789,N_11656);
xor U11928 (N_11928,N_11691,N_11716);
or U11929 (N_11929,N_11773,N_11752);
or U11930 (N_11930,N_11747,N_11744);
or U11931 (N_11931,N_11745,N_11734);
or U11932 (N_11932,N_11762,N_11734);
or U11933 (N_11933,N_11766,N_11695);
or U11934 (N_11934,N_11685,N_11709);
and U11935 (N_11935,N_11639,N_11619);
nor U11936 (N_11936,N_11666,N_11773);
and U11937 (N_11937,N_11731,N_11605);
nand U11938 (N_11938,N_11663,N_11659);
nand U11939 (N_11939,N_11640,N_11787);
and U11940 (N_11940,N_11688,N_11769);
xor U11941 (N_11941,N_11630,N_11753);
nand U11942 (N_11942,N_11754,N_11722);
or U11943 (N_11943,N_11732,N_11718);
or U11944 (N_11944,N_11712,N_11707);
and U11945 (N_11945,N_11654,N_11714);
or U11946 (N_11946,N_11756,N_11702);
nand U11947 (N_11947,N_11630,N_11781);
nor U11948 (N_11948,N_11607,N_11717);
nand U11949 (N_11949,N_11632,N_11659);
nand U11950 (N_11950,N_11703,N_11635);
nand U11951 (N_11951,N_11620,N_11742);
or U11952 (N_11952,N_11790,N_11685);
nor U11953 (N_11953,N_11681,N_11616);
nand U11954 (N_11954,N_11703,N_11689);
and U11955 (N_11955,N_11725,N_11674);
and U11956 (N_11956,N_11787,N_11606);
xor U11957 (N_11957,N_11684,N_11702);
nand U11958 (N_11958,N_11775,N_11744);
nor U11959 (N_11959,N_11740,N_11609);
or U11960 (N_11960,N_11672,N_11769);
and U11961 (N_11961,N_11637,N_11792);
nor U11962 (N_11962,N_11684,N_11723);
nor U11963 (N_11963,N_11787,N_11745);
xor U11964 (N_11964,N_11743,N_11768);
nand U11965 (N_11965,N_11628,N_11795);
nor U11966 (N_11966,N_11631,N_11614);
or U11967 (N_11967,N_11705,N_11761);
and U11968 (N_11968,N_11690,N_11763);
nand U11969 (N_11969,N_11769,N_11735);
or U11970 (N_11970,N_11767,N_11661);
or U11971 (N_11971,N_11783,N_11611);
nor U11972 (N_11972,N_11711,N_11650);
nor U11973 (N_11973,N_11777,N_11628);
and U11974 (N_11974,N_11662,N_11600);
and U11975 (N_11975,N_11613,N_11670);
nor U11976 (N_11976,N_11729,N_11724);
and U11977 (N_11977,N_11738,N_11749);
nand U11978 (N_11978,N_11743,N_11733);
nand U11979 (N_11979,N_11783,N_11705);
nand U11980 (N_11980,N_11653,N_11682);
nor U11981 (N_11981,N_11673,N_11760);
and U11982 (N_11982,N_11748,N_11787);
xor U11983 (N_11983,N_11734,N_11673);
nor U11984 (N_11984,N_11754,N_11674);
and U11985 (N_11985,N_11747,N_11614);
or U11986 (N_11986,N_11735,N_11698);
and U11987 (N_11987,N_11768,N_11664);
and U11988 (N_11988,N_11616,N_11779);
nand U11989 (N_11989,N_11660,N_11624);
or U11990 (N_11990,N_11708,N_11651);
or U11991 (N_11991,N_11621,N_11797);
and U11992 (N_11992,N_11625,N_11739);
nor U11993 (N_11993,N_11740,N_11622);
and U11994 (N_11994,N_11761,N_11735);
nand U11995 (N_11995,N_11690,N_11733);
nor U11996 (N_11996,N_11613,N_11726);
nor U11997 (N_11997,N_11742,N_11707);
nand U11998 (N_11998,N_11734,N_11624);
nor U11999 (N_11999,N_11640,N_11719);
and U12000 (N_12000,N_11922,N_11966);
or U12001 (N_12001,N_11880,N_11907);
nand U12002 (N_12002,N_11823,N_11834);
or U12003 (N_12003,N_11835,N_11949);
and U12004 (N_12004,N_11873,N_11985);
and U12005 (N_12005,N_11871,N_11831);
or U12006 (N_12006,N_11973,N_11964);
nand U12007 (N_12007,N_11923,N_11867);
or U12008 (N_12008,N_11970,N_11839);
nand U12009 (N_12009,N_11926,N_11953);
and U12010 (N_12010,N_11908,N_11899);
and U12011 (N_12011,N_11905,N_11897);
nand U12012 (N_12012,N_11844,N_11960);
or U12013 (N_12013,N_11884,N_11824);
nor U12014 (N_12014,N_11843,N_11801);
xor U12015 (N_12015,N_11861,N_11991);
nor U12016 (N_12016,N_11877,N_11963);
nand U12017 (N_12017,N_11993,N_11814);
nor U12018 (N_12018,N_11918,N_11864);
xnor U12019 (N_12019,N_11817,N_11948);
xnor U12020 (N_12020,N_11984,N_11950);
or U12021 (N_12021,N_11957,N_11933);
or U12022 (N_12022,N_11946,N_11997);
or U12023 (N_12023,N_11856,N_11828);
and U12024 (N_12024,N_11974,N_11837);
and U12025 (N_12025,N_11826,N_11800);
nand U12026 (N_12026,N_11872,N_11893);
or U12027 (N_12027,N_11958,N_11888);
nor U12028 (N_12028,N_11878,N_11956);
nor U12029 (N_12029,N_11804,N_11924);
nor U12030 (N_12030,N_11846,N_11821);
and U12031 (N_12031,N_11827,N_11981);
or U12032 (N_12032,N_11930,N_11935);
nor U12033 (N_12033,N_11860,N_11915);
and U12034 (N_12034,N_11862,N_11809);
xor U12035 (N_12035,N_11857,N_11932);
and U12036 (N_12036,N_11829,N_11876);
xor U12037 (N_12037,N_11977,N_11921);
or U12038 (N_12038,N_11845,N_11945);
or U12039 (N_12039,N_11965,N_11886);
or U12040 (N_12040,N_11810,N_11961);
and U12041 (N_12041,N_11927,N_11901);
nand U12042 (N_12042,N_11863,N_11943);
xnor U12043 (N_12043,N_11870,N_11937);
nand U12044 (N_12044,N_11836,N_11902);
nand U12045 (N_12045,N_11986,N_11978);
xor U12046 (N_12046,N_11842,N_11920);
and U12047 (N_12047,N_11904,N_11941);
nand U12048 (N_12048,N_11975,N_11962);
xor U12049 (N_12049,N_11995,N_11822);
nand U12050 (N_12050,N_11881,N_11840);
nand U12051 (N_12051,N_11979,N_11811);
or U12052 (N_12052,N_11925,N_11896);
nand U12053 (N_12053,N_11802,N_11833);
nand U12054 (N_12054,N_11882,N_11971);
xor U12055 (N_12055,N_11848,N_11955);
xnor U12056 (N_12056,N_11853,N_11883);
xor U12057 (N_12057,N_11994,N_11969);
nor U12058 (N_12058,N_11989,N_11940);
nor U12059 (N_12059,N_11976,N_11917);
nor U12060 (N_12060,N_11938,N_11890);
and U12061 (N_12061,N_11990,N_11913);
and U12062 (N_12062,N_11911,N_11912);
and U12063 (N_12063,N_11929,N_11931);
nand U12064 (N_12064,N_11869,N_11858);
and U12065 (N_12065,N_11952,N_11874);
xnor U12066 (N_12066,N_11898,N_11852);
nand U12067 (N_12067,N_11954,N_11847);
xnor U12068 (N_12068,N_11889,N_11914);
and U12069 (N_12069,N_11919,N_11859);
and U12070 (N_12070,N_11875,N_11999);
xnor U12071 (N_12071,N_11818,N_11895);
or U12072 (N_12072,N_11936,N_11832);
xnor U12073 (N_12073,N_11815,N_11934);
xor U12074 (N_12074,N_11996,N_11998);
or U12075 (N_12075,N_11825,N_11959);
or U12076 (N_12076,N_11806,N_11928);
xor U12077 (N_12077,N_11900,N_11944);
xnor U12078 (N_12078,N_11866,N_11803);
xor U12079 (N_12079,N_11807,N_11980);
or U12080 (N_12080,N_11850,N_11951);
or U12081 (N_12081,N_11988,N_11854);
nand U12082 (N_12082,N_11916,N_11865);
or U12083 (N_12083,N_11868,N_11987);
or U12084 (N_12084,N_11830,N_11983);
nor U12085 (N_12085,N_11942,N_11819);
nand U12086 (N_12086,N_11906,N_11813);
or U12087 (N_12087,N_11939,N_11855);
or U12088 (N_12088,N_11816,N_11909);
or U12089 (N_12089,N_11805,N_11838);
nor U12090 (N_12090,N_11968,N_11812);
nor U12091 (N_12091,N_11992,N_11841);
and U12092 (N_12092,N_11891,N_11892);
and U12093 (N_12093,N_11967,N_11947);
nand U12094 (N_12094,N_11903,N_11972);
and U12095 (N_12095,N_11879,N_11820);
xnor U12096 (N_12096,N_11851,N_11982);
xnor U12097 (N_12097,N_11910,N_11808);
nand U12098 (N_12098,N_11887,N_11894);
and U12099 (N_12099,N_11849,N_11885);
nand U12100 (N_12100,N_11859,N_11910);
and U12101 (N_12101,N_11941,N_11997);
nand U12102 (N_12102,N_11969,N_11956);
nand U12103 (N_12103,N_11817,N_11984);
nor U12104 (N_12104,N_11995,N_11913);
nor U12105 (N_12105,N_11880,N_11849);
nor U12106 (N_12106,N_11902,N_11959);
nand U12107 (N_12107,N_11962,N_11974);
nor U12108 (N_12108,N_11935,N_11841);
nor U12109 (N_12109,N_11909,N_11811);
or U12110 (N_12110,N_11903,N_11816);
and U12111 (N_12111,N_11913,N_11997);
or U12112 (N_12112,N_11928,N_11965);
nand U12113 (N_12113,N_11968,N_11961);
nor U12114 (N_12114,N_11980,N_11904);
xnor U12115 (N_12115,N_11914,N_11966);
xnor U12116 (N_12116,N_11821,N_11818);
xnor U12117 (N_12117,N_11852,N_11932);
and U12118 (N_12118,N_11839,N_11977);
xor U12119 (N_12119,N_11806,N_11841);
nor U12120 (N_12120,N_11952,N_11892);
and U12121 (N_12121,N_11868,N_11961);
xnor U12122 (N_12122,N_11869,N_11900);
nand U12123 (N_12123,N_11873,N_11887);
nand U12124 (N_12124,N_11843,N_11952);
and U12125 (N_12125,N_11916,N_11810);
nand U12126 (N_12126,N_11955,N_11828);
or U12127 (N_12127,N_11800,N_11982);
and U12128 (N_12128,N_11909,N_11966);
nand U12129 (N_12129,N_11858,N_11850);
or U12130 (N_12130,N_11801,N_11802);
nand U12131 (N_12131,N_11977,N_11889);
xor U12132 (N_12132,N_11915,N_11813);
nand U12133 (N_12133,N_11899,N_11957);
or U12134 (N_12134,N_11819,N_11821);
xor U12135 (N_12135,N_11834,N_11839);
and U12136 (N_12136,N_11837,N_11961);
xor U12137 (N_12137,N_11916,N_11872);
nor U12138 (N_12138,N_11914,N_11911);
nor U12139 (N_12139,N_11855,N_11927);
nand U12140 (N_12140,N_11823,N_11800);
nand U12141 (N_12141,N_11925,N_11824);
or U12142 (N_12142,N_11833,N_11880);
and U12143 (N_12143,N_11827,N_11931);
nand U12144 (N_12144,N_11820,N_11916);
nor U12145 (N_12145,N_11862,N_11814);
and U12146 (N_12146,N_11831,N_11836);
or U12147 (N_12147,N_11919,N_11889);
nand U12148 (N_12148,N_11828,N_11834);
nand U12149 (N_12149,N_11894,N_11802);
nand U12150 (N_12150,N_11844,N_11896);
and U12151 (N_12151,N_11822,N_11985);
or U12152 (N_12152,N_11924,N_11943);
or U12153 (N_12153,N_11961,N_11886);
or U12154 (N_12154,N_11926,N_11846);
and U12155 (N_12155,N_11950,N_11994);
and U12156 (N_12156,N_11902,N_11857);
and U12157 (N_12157,N_11808,N_11872);
nor U12158 (N_12158,N_11808,N_11840);
nand U12159 (N_12159,N_11813,N_11961);
nand U12160 (N_12160,N_11923,N_11912);
xnor U12161 (N_12161,N_11836,N_11927);
and U12162 (N_12162,N_11930,N_11874);
or U12163 (N_12163,N_11882,N_11817);
nor U12164 (N_12164,N_11875,N_11854);
nor U12165 (N_12165,N_11858,N_11972);
and U12166 (N_12166,N_11903,N_11964);
xnor U12167 (N_12167,N_11871,N_11834);
nand U12168 (N_12168,N_11811,N_11913);
and U12169 (N_12169,N_11900,N_11875);
nor U12170 (N_12170,N_11946,N_11949);
xnor U12171 (N_12171,N_11855,N_11902);
nor U12172 (N_12172,N_11815,N_11920);
or U12173 (N_12173,N_11946,N_11830);
nor U12174 (N_12174,N_11901,N_11862);
xnor U12175 (N_12175,N_11913,N_11904);
or U12176 (N_12176,N_11905,N_11871);
and U12177 (N_12177,N_11970,N_11963);
and U12178 (N_12178,N_11898,N_11945);
xor U12179 (N_12179,N_11826,N_11870);
nor U12180 (N_12180,N_11875,N_11907);
or U12181 (N_12181,N_11844,N_11916);
or U12182 (N_12182,N_11937,N_11954);
and U12183 (N_12183,N_11919,N_11877);
nor U12184 (N_12184,N_11938,N_11912);
nor U12185 (N_12185,N_11888,N_11843);
or U12186 (N_12186,N_11829,N_11925);
xnor U12187 (N_12187,N_11862,N_11873);
nand U12188 (N_12188,N_11872,N_11871);
xnor U12189 (N_12189,N_11883,N_11907);
and U12190 (N_12190,N_11882,N_11888);
nand U12191 (N_12191,N_11821,N_11919);
nand U12192 (N_12192,N_11911,N_11929);
and U12193 (N_12193,N_11823,N_11828);
nor U12194 (N_12194,N_11968,N_11941);
nor U12195 (N_12195,N_11948,N_11814);
nand U12196 (N_12196,N_11845,N_11882);
or U12197 (N_12197,N_11887,N_11879);
nand U12198 (N_12198,N_11874,N_11892);
xnor U12199 (N_12199,N_11913,N_11840);
or U12200 (N_12200,N_12174,N_12126);
nor U12201 (N_12201,N_12018,N_12020);
or U12202 (N_12202,N_12140,N_12038);
xnor U12203 (N_12203,N_12099,N_12109);
or U12204 (N_12204,N_12035,N_12139);
or U12205 (N_12205,N_12125,N_12007);
nand U12206 (N_12206,N_12144,N_12155);
or U12207 (N_12207,N_12012,N_12003);
nand U12208 (N_12208,N_12179,N_12138);
nor U12209 (N_12209,N_12188,N_12096);
and U12210 (N_12210,N_12192,N_12122);
nand U12211 (N_12211,N_12142,N_12197);
and U12212 (N_12212,N_12199,N_12068);
nor U12213 (N_12213,N_12130,N_12158);
nor U12214 (N_12214,N_12061,N_12101);
nor U12215 (N_12215,N_12047,N_12127);
nand U12216 (N_12216,N_12031,N_12080);
or U12217 (N_12217,N_12186,N_12041);
or U12218 (N_12218,N_12062,N_12052);
or U12219 (N_12219,N_12073,N_12180);
nor U12220 (N_12220,N_12048,N_12094);
and U12221 (N_12221,N_12100,N_12193);
xor U12222 (N_12222,N_12009,N_12059);
and U12223 (N_12223,N_12161,N_12055);
and U12224 (N_12224,N_12065,N_12103);
and U12225 (N_12225,N_12106,N_12071);
nor U12226 (N_12226,N_12115,N_12011);
or U12227 (N_12227,N_12028,N_12133);
nor U12228 (N_12228,N_12019,N_12163);
nor U12229 (N_12229,N_12078,N_12081);
nor U12230 (N_12230,N_12150,N_12086);
nor U12231 (N_12231,N_12119,N_12146);
or U12232 (N_12232,N_12016,N_12051);
or U12233 (N_12233,N_12176,N_12175);
or U12234 (N_12234,N_12151,N_12191);
xnor U12235 (N_12235,N_12006,N_12136);
nand U12236 (N_12236,N_12043,N_12025);
nor U12237 (N_12237,N_12046,N_12069);
or U12238 (N_12238,N_12110,N_12024);
nand U12239 (N_12239,N_12195,N_12004);
nand U12240 (N_12240,N_12160,N_12148);
or U12241 (N_12241,N_12084,N_12105);
nor U12242 (N_12242,N_12164,N_12107);
nor U12243 (N_12243,N_12167,N_12137);
or U12244 (N_12244,N_12097,N_12085);
nor U12245 (N_12245,N_12005,N_12091);
nand U12246 (N_12246,N_12066,N_12087);
nand U12247 (N_12247,N_12014,N_12098);
and U12248 (N_12248,N_12143,N_12172);
and U12249 (N_12249,N_12108,N_12056);
nand U12250 (N_12250,N_12153,N_12002);
nor U12251 (N_12251,N_12134,N_12162);
nand U12252 (N_12252,N_12022,N_12183);
or U12253 (N_12253,N_12178,N_12112);
and U12254 (N_12254,N_12171,N_12154);
or U12255 (N_12255,N_12039,N_12045);
nand U12256 (N_12256,N_12187,N_12182);
and U12257 (N_12257,N_12030,N_12181);
or U12258 (N_12258,N_12128,N_12000);
nor U12259 (N_12259,N_12185,N_12170);
and U12260 (N_12260,N_12189,N_12060);
or U12261 (N_12261,N_12147,N_12013);
and U12262 (N_12262,N_12169,N_12082);
and U12263 (N_12263,N_12194,N_12102);
and U12264 (N_12264,N_12015,N_12032);
and U12265 (N_12265,N_12053,N_12177);
or U12266 (N_12266,N_12117,N_12074);
xor U12267 (N_12267,N_12124,N_12064);
and U12268 (N_12268,N_12121,N_12077);
nor U12269 (N_12269,N_12168,N_12029);
and U12270 (N_12270,N_12131,N_12040);
xnor U12271 (N_12271,N_12196,N_12149);
and U12272 (N_12272,N_12076,N_12063);
nor U12273 (N_12273,N_12054,N_12072);
nor U12274 (N_12274,N_12118,N_12044);
nor U12275 (N_12275,N_12008,N_12027);
nor U12276 (N_12276,N_12157,N_12089);
or U12277 (N_12277,N_12104,N_12116);
nor U12278 (N_12278,N_12114,N_12049);
or U12279 (N_12279,N_12058,N_12132);
and U12280 (N_12280,N_12090,N_12034);
or U12281 (N_12281,N_12159,N_12057);
nor U12282 (N_12282,N_12070,N_12037);
and U12283 (N_12283,N_12042,N_12088);
or U12284 (N_12284,N_12152,N_12165);
or U12285 (N_12285,N_12092,N_12123);
and U12286 (N_12286,N_12190,N_12129);
or U12287 (N_12287,N_12075,N_12093);
nor U12288 (N_12288,N_12141,N_12184);
nand U12289 (N_12289,N_12145,N_12173);
nor U12290 (N_12290,N_12067,N_12079);
nor U12291 (N_12291,N_12198,N_12036);
and U12292 (N_12292,N_12050,N_12113);
xnor U12293 (N_12293,N_12001,N_12095);
nand U12294 (N_12294,N_12033,N_12026);
nor U12295 (N_12295,N_12111,N_12010);
nor U12296 (N_12296,N_12156,N_12017);
or U12297 (N_12297,N_12135,N_12120);
or U12298 (N_12298,N_12023,N_12166);
or U12299 (N_12299,N_12083,N_12021);
nand U12300 (N_12300,N_12148,N_12063);
nand U12301 (N_12301,N_12008,N_12046);
nand U12302 (N_12302,N_12000,N_12165);
and U12303 (N_12303,N_12091,N_12145);
nand U12304 (N_12304,N_12070,N_12033);
and U12305 (N_12305,N_12097,N_12042);
nand U12306 (N_12306,N_12167,N_12164);
xnor U12307 (N_12307,N_12120,N_12157);
nor U12308 (N_12308,N_12014,N_12111);
and U12309 (N_12309,N_12167,N_12196);
nor U12310 (N_12310,N_12040,N_12168);
or U12311 (N_12311,N_12044,N_12097);
xnor U12312 (N_12312,N_12051,N_12030);
and U12313 (N_12313,N_12099,N_12033);
or U12314 (N_12314,N_12114,N_12095);
nand U12315 (N_12315,N_12100,N_12045);
nand U12316 (N_12316,N_12084,N_12110);
nand U12317 (N_12317,N_12134,N_12124);
nand U12318 (N_12318,N_12079,N_12043);
or U12319 (N_12319,N_12191,N_12051);
nand U12320 (N_12320,N_12157,N_12167);
or U12321 (N_12321,N_12027,N_12063);
or U12322 (N_12322,N_12148,N_12153);
and U12323 (N_12323,N_12198,N_12015);
or U12324 (N_12324,N_12148,N_12017);
nor U12325 (N_12325,N_12011,N_12124);
and U12326 (N_12326,N_12181,N_12196);
nor U12327 (N_12327,N_12090,N_12124);
or U12328 (N_12328,N_12148,N_12009);
nor U12329 (N_12329,N_12006,N_12094);
nor U12330 (N_12330,N_12187,N_12158);
nor U12331 (N_12331,N_12009,N_12076);
or U12332 (N_12332,N_12054,N_12099);
and U12333 (N_12333,N_12057,N_12056);
or U12334 (N_12334,N_12066,N_12110);
nor U12335 (N_12335,N_12127,N_12038);
nor U12336 (N_12336,N_12071,N_12064);
nor U12337 (N_12337,N_12068,N_12056);
and U12338 (N_12338,N_12070,N_12071);
and U12339 (N_12339,N_12090,N_12188);
xnor U12340 (N_12340,N_12024,N_12055);
and U12341 (N_12341,N_12132,N_12015);
and U12342 (N_12342,N_12033,N_12161);
nand U12343 (N_12343,N_12052,N_12032);
nor U12344 (N_12344,N_12112,N_12154);
nand U12345 (N_12345,N_12124,N_12149);
and U12346 (N_12346,N_12171,N_12108);
or U12347 (N_12347,N_12194,N_12086);
nand U12348 (N_12348,N_12055,N_12056);
nor U12349 (N_12349,N_12133,N_12121);
nand U12350 (N_12350,N_12108,N_12107);
nor U12351 (N_12351,N_12118,N_12137);
or U12352 (N_12352,N_12114,N_12072);
nor U12353 (N_12353,N_12014,N_12072);
xor U12354 (N_12354,N_12121,N_12170);
or U12355 (N_12355,N_12185,N_12133);
or U12356 (N_12356,N_12003,N_12028);
or U12357 (N_12357,N_12075,N_12056);
and U12358 (N_12358,N_12060,N_12112);
xor U12359 (N_12359,N_12012,N_12162);
or U12360 (N_12360,N_12030,N_12149);
nor U12361 (N_12361,N_12193,N_12053);
and U12362 (N_12362,N_12134,N_12145);
or U12363 (N_12363,N_12131,N_12137);
and U12364 (N_12364,N_12053,N_12160);
or U12365 (N_12365,N_12107,N_12028);
nor U12366 (N_12366,N_12081,N_12025);
nor U12367 (N_12367,N_12143,N_12159);
nand U12368 (N_12368,N_12008,N_12166);
nor U12369 (N_12369,N_12050,N_12044);
nand U12370 (N_12370,N_12193,N_12068);
nor U12371 (N_12371,N_12172,N_12060);
nor U12372 (N_12372,N_12001,N_12195);
nor U12373 (N_12373,N_12002,N_12113);
nor U12374 (N_12374,N_12173,N_12112);
nor U12375 (N_12375,N_12031,N_12165);
and U12376 (N_12376,N_12090,N_12078);
or U12377 (N_12377,N_12112,N_12035);
nor U12378 (N_12378,N_12001,N_12154);
or U12379 (N_12379,N_12122,N_12146);
and U12380 (N_12380,N_12115,N_12122);
or U12381 (N_12381,N_12043,N_12063);
and U12382 (N_12382,N_12078,N_12006);
nor U12383 (N_12383,N_12173,N_12155);
nor U12384 (N_12384,N_12159,N_12192);
or U12385 (N_12385,N_12171,N_12188);
or U12386 (N_12386,N_12094,N_12192);
nor U12387 (N_12387,N_12080,N_12172);
nor U12388 (N_12388,N_12045,N_12098);
and U12389 (N_12389,N_12116,N_12182);
nor U12390 (N_12390,N_12112,N_12080);
and U12391 (N_12391,N_12062,N_12082);
or U12392 (N_12392,N_12110,N_12139);
or U12393 (N_12393,N_12010,N_12149);
nor U12394 (N_12394,N_12118,N_12026);
nand U12395 (N_12395,N_12000,N_12192);
and U12396 (N_12396,N_12013,N_12090);
nor U12397 (N_12397,N_12003,N_12147);
or U12398 (N_12398,N_12155,N_12058);
nor U12399 (N_12399,N_12015,N_12149);
nor U12400 (N_12400,N_12287,N_12288);
and U12401 (N_12401,N_12239,N_12341);
or U12402 (N_12402,N_12221,N_12370);
xor U12403 (N_12403,N_12213,N_12353);
or U12404 (N_12404,N_12336,N_12329);
nand U12405 (N_12405,N_12318,N_12202);
nor U12406 (N_12406,N_12248,N_12223);
xnor U12407 (N_12407,N_12256,N_12286);
or U12408 (N_12408,N_12343,N_12242);
and U12409 (N_12409,N_12381,N_12290);
nor U12410 (N_12410,N_12241,N_12210);
and U12411 (N_12411,N_12280,N_12283);
and U12412 (N_12412,N_12293,N_12279);
nand U12413 (N_12413,N_12332,N_12383);
and U12414 (N_12414,N_12333,N_12229);
nand U12415 (N_12415,N_12396,N_12384);
or U12416 (N_12416,N_12296,N_12399);
xor U12417 (N_12417,N_12390,N_12207);
or U12418 (N_12418,N_12310,N_12204);
and U12419 (N_12419,N_12216,N_12226);
and U12420 (N_12420,N_12214,N_12386);
xor U12421 (N_12421,N_12316,N_12355);
xnor U12422 (N_12422,N_12259,N_12325);
nand U12423 (N_12423,N_12376,N_12361);
nor U12424 (N_12424,N_12227,N_12299);
nand U12425 (N_12425,N_12208,N_12366);
xor U12426 (N_12426,N_12393,N_12245);
nand U12427 (N_12427,N_12362,N_12275);
nand U12428 (N_12428,N_12206,N_12368);
or U12429 (N_12429,N_12235,N_12262);
and U12430 (N_12430,N_12250,N_12268);
or U12431 (N_12431,N_12385,N_12311);
and U12432 (N_12432,N_12301,N_12252);
nand U12433 (N_12433,N_12367,N_12211);
or U12434 (N_12434,N_12265,N_12369);
and U12435 (N_12435,N_12324,N_12326);
nand U12436 (N_12436,N_12398,N_12261);
and U12437 (N_12437,N_12269,N_12371);
and U12438 (N_12438,N_12349,N_12345);
nand U12439 (N_12439,N_12321,N_12330);
nor U12440 (N_12440,N_12328,N_12388);
and U12441 (N_12441,N_12323,N_12304);
nand U12442 (N_12442,N_12253,N_12247);
or U12443 (N_12443,N_12334,N_12379);
and U12444 (N_12444,N_12307,N_12317);
xnor U12445 (N_12445,N_12305,N_12258);
or U12446 (N_12446,N_12295,N_12282);
and U12447 (N_12447,N_12201,N_12277);
and U12448 (N_12448,N_12205,N_12387);
xnor U12449 (N_12449,N_12392,N_12342);
xnor U12450 (N_12450,N_12270,N_12374);
and U12451 (N_12451,N_12327,N_12292);
and U12452 (N_12452,N_12306,N_12313);
or U12453 (N_12453,N_12224,N_12237);
nor U12454 (N_12454,N_12243,N_12234);
and U12455 (N_12455,N_12364,N_12281);
nor U12456 (N_12456,N_12373,N_12391);
or U12457 (N_12457,N_12260,N_12320);
and U12458 (N_12458,N_12359,N_12338);
nor U12459 (N_12459,N_12394,N_12322);
nand U12460 (N_12460,N_12382,N_12244);
xor U12461 (N_12461,N_12284,N_12230);
xnor U12462 (N_12462,N_12222,N_12218);
and U12463 (N_12463,N_12215,N_12231);
nand U12464 (N_12464,N_12238,N_12251);
nor U12465 (N_12465,N_12337,N_12236);
and U12466 (N_12466,N_12200,N_12397);
xor U12467 (N_12467,N_12340,N_12240);
nand U12468 (N_12468,N_12255,N_12285);
or U12469 (N_12469,N_12389,N_12346);
nor U12470 (N_12470,N_12257,N_12273);
xnor U12471 (N_12471,N_12302,N_12267);
nor U12472 (N_12472,N_12380,N_12350);
nand U12473 (N_12473,N_12395,N_12378);
and U12474 (N_12474,N_12203,N_12246);
or U12475 (N_12475,N_12348,N_12263);
nand U12476 (N_12476,N_12264,N_12358);
or U12477 (N_12477,N_12219,N_12266);
nor U12478 (N_12478,N_12254,N_12309);
nand U12479 (N_12479,N_12274,N_12249);
and U12480 (N_12480,N_12272,N_12351);
nand U12481 (N_12481,N_12303,N_12291);
and U12482 (N_12482,N_12276,N_12352);
nor U12483 (N_12483,N_12217,N_12339);
or U12484 (N_12484,N_12297,N_12314);
xnor U12485 (N_12485,N_12335,N_12356);
or U12486 (N_12486,N_12360,N_12331);
nand U12487 (N_12487,N_12289,N_12375);
nand U12488 (N_12488,N_12344,N_12372);
xnor U12489 (N_12489,N_12357,N_12294);
or U12490 (N_12490,N_12354,N_12298);
and U12491 (N_12491,N_12365,N_12233);
and U12492 (N_12492,N_12363,N_12212);
nand U12493 (N_12493,N_12278,N_12209);
nor U12494 (N_12494,N_12271,N_12228);
nor U12495 (N_12495,N_12300,N_12308);
nor U12496 (N_12496,N_12315,N_12319);
xnor U12497 (N_12497,N_12220,N_12225);
and U12498 (N_12498,N_12312,N_12377);
and U12499 (N_12499,N_12347,N_12232);
and U12500 (N_12500,N_12312,N_12232);
nor U12501 (N_12501,N_12384,N_12317);
or U12502 (N_12502,N_12277,N_12290);
or U12503 (N_12503,N_12228,N_12260);
nor U12504 (N_12504,N_12396,N_12226);
nor U12505 (N_12505,N_12211,N_12342);
xor U12506 (N_12506,N_12252,N_12248);
and U12507 (N_12507,N_12338,N_12236);
nor U12508 (N_12508,N_12269,N_12326);
nand U12509 (N_12509,N_12223,N_12310);
and U12510 (N_12510,N_12246,N_12360);
or U12511 (N_12511,N_12356,N_12297);
or U12512 (N_12512,N_12225,N_12223);
or U12513 (N_12513,N_12354,N_12340);
xnor U12514 (N_12514,N_12383,N_12205);
xor U12515 (N_12515,N_12371,N_12308);
or U12516 (N_12516,N_12394,N_12220);
and U12517 (N_12517,N_12317,N_12231);
nand U12518 (N_12518,N_12228,N_12345);
nor U12519 (N_12519,N_12353,N_12221);
nor U12520 (N_12520,N_12283,N_12233);
nand U12521 (N_12521,N_12311,N_12362);
or U12522 (N_12522,N_12221,N_12360);
xor U12523 (N_12523,N_12356,N_12282);
or U12524 (N_12524,N_12214,N_12266);
or U12525 (N_12525,N_12255,N_12296);
and U12526 (N_12526,N_12362,N_12241);
or U12527 (N_12527,N_12371,N_12275);
and U12528 (N_12528,N_12327,N_12261);
nand U12529 (N_12529,N_12306,N_12223);
xnor U12530 (N_12530,N_12326,N_12365);
or U12531 (N_12531,N_12269,N_12325);
and U12532 (N_12532,N_12347,N_12318);
nand U12533 (N_12533,N_12247,N_12266);
nor U12534 (N_12534,N_12276,N_12263);
or U12535 (N_12535,N_12229,N_12342);
or U12536 (N_12536,N_12363,N_12267);
or U12537 (N_12537,N_12250,N_12397);
or U12538 (N_12538,N_12237,N_12311);
and U12539 (N_12539,N_12306,N_12216);
and U12540 (N_12540,N_12386,N_12217);
or U12541 (N_12541,N_12207,N_12295);
or U12542 (N_12542,N_12263,N_12283);
and U12543 (N_12543,N_12281,N_12211);
and U12544 (N_12544,N_12252,N_12343);
or U12545 (N_12545,N_12242,N_12336);
and U12546 (N_12546,N_12257,N_12358);
nand U12547 (N_12547,N_12298,N_12381);
or U12548 (N_12548,N_12375,N_12234);
nand U12549 (N_12549,N_12264,N_12286);
nor U12550 (N_12550,N_12229,N_12295);
or U12551 (N_12551,N_12304,N_12288);
nor U12552 (N_12552,N_12398,N_12323);
nand U12553 (N_12553,N_12394,N_12315);
or U12554 (N_12554,N_12336,N_12209);
or U12555 (N_12555,N_12205,N_12329);
and U12556 (N_12556,N_12329,N_12293);
nor U12557 (N_12557,N_12378,N_12234);
xnor U12558 (N_12558,N_12294,N_12386);
nor U12559 (N_12559,N_12204,N_12356);
xor U12560 (N_12560,N_12317,N_12291);
and U12561 (N_12561,N_12376,N_12395);
and U12562 (N_12562,N_12387,N_12243);
nor U12563 (N_12563,N_12303,N_12376);
or U12564 (N_12564,N_12314,N_12278);
nor U12565 (N_12565,N_12384,N_12211);
nor U12566 (N_12566,N_12325,N_12338);
nand U12567 (N_12567,N_12365,N_12213);
and U12568 (N_12568,N_12347,N_12359);
and U12569 (N_12569,N_12223,N_12350);
xnor U12570 (N_12570,N_12370,N_12365);
nor U12571 (N_12571,N_12359,N_12371);
nand U12572 (N_12572,N_12247,N_12207);
nor U12573 (N_12573,N_12304,N_12298);
xor U12574 (N_12574,N_12248,N_12295);
nor U12575 (N_12575,N_12395,N_12277);
or U12576 (N_12576,N_12224,N_12281);
and U12577 (N_12577,N_12218,N_12200);
nand U12578 (N_12578,N_12391,N_12243);
or U12579 (N_12579,N_12324,N_12355);
xnor U12580 (N_12580,N_12245,N_12383);
nor U12581 (N_12581,N_12273,N_12360);
and U12582 (N_12582,N_12213,N_12356);
and U12583 (N_12583,N_12393,N_12257);
and U12584 (N_12584,N_12218,N_12267);
nand U12585 (N_12585,N_12386,N_12234);
xor U12586 (N_12586,N_12377,N_12376);
nor U12587 (N_12587,N_12359,N_12333);
nor U12588 (N_12588,N_12301,N_12211);
nor U12589 (N_12589,N_12265,N_12331);
nand U12590 (N_12590,N_12245,N_12311);
nand U12591 (N_12591,N_12205,N_12263);
nor U12592 (N_12592,N_12336,N_12279);
nor U12593 (N_12593,N_12266,N_12254);
nor U12594 (N_12594,N_12354,N_12349);
nor U12595 (N_12595,N_12229,N_12247);
nand U12596 (N_12596,N_12223,N_12316);
nand U12597 (N_12597,N_12371,N_12216);
nor U12598 (N_12598,N_12305,N_12249);
nor U12599 (N_12599,N_12249,N_12205);
and U12600 (N_12600,N_12526,N_12492);
nand U12601 (N_12601,N_12562,N_12591);
or U12602 (N_12602,N_12453,N_12411);
or U12603 (N_12603,N_12582,N_12487);
xor U12604 (N_12604,N_12572,N_12468);
nor U12605 (N_12605,N_12529,N_12538);
or U12606 (N_12606,N_12420,N_12508);
and U12607 (N_12607,N_12449,N_12592);
nand U12608 (N_12608,N_12481,N_12563);
nand U12609 (N_12609,N_12458,N_12524);
xor U12610 (N_12610,N_12541,N_12558);
or U12611 (N_12611,N_12535,N_12551);
and U12612 (N_12612,N_12555,N_12596);
or U12613 (N_12613,N_12403,N_12486);
and U12614 (N_12614,N_12514,N_12435);
or U12615 (N_12615,N_12471,N_12595);
and U12616 (N_12616,N_12495,N_12525);
nor U12617 (N_12617,N_12578,N_12440);
and U12618 (N_12618,N_12587,N_12569);
or U12619 (N_12619,N_12549,N_12465);
nand U12620 (N_12620,N_12427,N_12410);
nand U12621 (N_12621,N_12405,N_12447);
nor U12622 (N_12622,N_12527,N_12590);
nor U12623 (N_12623,N_12476,N_12485);
and U12624 (N_12624,N_12452,N_12546);
or U12625 (N_12625,N_12533,N_12478);
nor U12626 (N_12626,N_12509,N_12571);
and U12627 (N_12627,N_12483,N_12424);
or U12628 (N_12628,N_12581,N_12473);
nand U12629 (N_12629,N_12488,N_12474);
xnor U12630 (N_12630,N_12461,N_12414);
and U12631 (N_12631,N_12413,N_12537);
nand U12632 (N_12632,N_12511,N_12441);
nand U12633 (N_12633,N_12536,N_12497);
nand U12634 (N_12634,N_12520,N_12530);
and U12635 (N_12635,N_12517,N_12598);
and U12636 (N_12636,N_12489,N_12510);
or U12637 (N_12637,N_12532,N_12460);
nor U12638 (N_12638,N_12574,N_12498);
nand U12639 (N_12639,N_12432,N_12428);
and U12640 (N_12640,N_12426,N_12505);
and U12641 (N_12641,N_12470,N_12576);
xnor U12642 (N_12642,N_12518,N_12455);
or U12643 (N_12643,N_12528,N_12573);
nand U12644 (N_12644,N_12456,N_12431);
or U12645 (N_12645,N_12545,N_12457);
nor U12646 (N_12646,N_12547,N_12519);
nand U12647 (N_12647,N_12503,N_12531);
xnor U12648 (N_12648,N_12448,N_12513);
or U12649 (N_12649,N_12472,N_12522);
and U12650 (N_12650,N_12521,N_12542);
and U12651 (N_12651,N_12480,N_12477);
nor U12652 (N_12652,N_12442,N_12425);
nand U12653 (N_12653,N_12512,N_12479);
and U12654 (N_12654,N_12422,N_12500);
or U12655 (N_12655,N_12543,N_12561);
and U12656 (N_12656,N_12534,N_12554);
nor U12657 (N_12657,N_12567,N_12516);
nor U12658 (N_12658,N_12482,N_12484);
nand U12659 (N_12659,N_12586,N_12423);
and U12660 (N_12660,N_12557,N_12540);
or U12661 (N_12661,N_12443,N_12594);
and U12662 (N_12662,N_12406,N_12560);
or U12663 (N_12663,N_12417,N_12589);
nand U12664 (N_12664,N_12407,N_12467);
nor U12665 (N_12665,N_12416,N_12409);
xor U12666 (N_12666,N_12577,N_12491);
and U12667 (N_12667,N_12466,N_12418);
or U12668 (N_12668,N_12493,N_12553);
nor U12669 (N_12669,N_12515,N_12463);
or U12670 (N_12670,N_12436,N_12499);
nand U12671 (N_12671,N_12597,N_12496);
nand U12672 (N_12672,N_12575,N_12579);
nand U12673 (N_12673,N_12494,N_12550);
nor U12674 (N_12674,N_12593,N_12556);
nand U12675 (N_12675,N_12568,N_12408);
nor U12676 (N_12676,N_12565,N_12459);
or U12677 (N_12677,N_12599,N_12490);
or U12678 (N_12678,N_12444,N_12415);
or U12679 (N_12679,N_12412,N_12451);
and U12680 (N_12680,N_12507,N_12539);
and U12681 (N_12681,N_12438,N_12437);
or U12682 (N_12682,N_12429,N_12523);
or U12683 (N_12683,N_12504,N_12433);
or U12684 (N_12684,N_12462,N_12450);
or U12685 (N_12685,N_12566,N_12464);
nor U12686 (N_12686,N_12502,N_12400);
nand U12687 (N_12687,N_12419,N_12454);
nand U12688 (N_12688,N_12401,N_12430);
and U12689 (N_12689,N_12434,N_12570);
or U12690 (N_12690,N_12580,N_12475);
or U12691 (N_12691,N_12584,N_12588);
or U12692 (N_12692,N_12552,N_12439);
nand U12693 (N_12693,N_12548,N_12544);
nand U12694 (N_12694,N_12421,N_12585);
nand U12695 (N_12695,N_12404,N_12564);
nor U12696 (N_12696,N_12583,N_12559);
and U12697 (N_12697,N_12501,N_12469);
nor U12698 (N_12698,N_12445,N_12402);
nand U12699 (N_12699,N_12506,N_12446);
nor U12700 (N_12700,N_12422,N_12479);
or U12701 (N_12701,N_12500,N_12471);
nand U12702 (N_12702,N_12548,N_12408);
and U12703 (N_12703,N_12410,N_12431);
xor U12704 (N_12704,N_12552,N_12489);
nand U12705 (N_12705,N_12514,N_12461);
xor U12706 (N_12706,N_12427,N_12405);
nor U12707 (N_12707,N_12533,N_12439);
and U12708 (N_12708,N_12457,N_12454);
or U12709 (N_12709,N_12549,N_12548);
nor U12710 (N_12710,N_12544,N_12430);
or U12711 (N_12711,N_12460,N_12430);
and U12712 (N_12712,N_12494,N_12506);
nor U12713 (N_12713,N_12487,N_12410);
xor U12714 (N_12714,N_12521,N_12426);
or U12715 (N_12715,N_12453,N_12525);
and U12716 (N_12716,N_12430,N_12482);
and U12717 (N_12717,N_12479,N_12576);
nand U12718 (N_12718,N_12533,N_12594);
nor U12719 (N_12719,N_12407,N_12509);
and U12720 (N_12720,N_12477,N_12425);
xor U12721 (N_12721,N_12520,N_12454);
or U12722 (N_12722,N_12515,N_12545);
or U12723 (N_12723,N_12411,N_12465);
or U12724 (N_12724,N_12440,N_12411);
nor U12725 (N_12725,N_12468,N_12589);
nor U12726 (N_12726,N_12574,N_12507);
xor U12727 (N_12727,N_12587,N_12570);
nand U12728 (N_12728,N_12561,N_12490);
nand U12729 (N_12729,N_12445,N_12581);
xor U12730 (N_12730,N_12403,N_12534);
xor U12731 (N_12731,N_12447,N_12502);
and U12732 (N_12732,N_12401,N_12571);
nor U12733 (N_12733,N_12599,N_12451);
nor U12734 (N_12734,N_12400,N_12559);
nor U12735 (N_12735,N_12528,N_12495);
nor U12736 (N_12736,N_12517,N_12571);
and U12737 (N_12737,N_12445,N_12532);
nand U12738 (N_12738,N_12589,N_12439);
xor U12739 (N_12739,N_12591,N_12563);
xor U12740 (N_12740,N_12456,N_12534);
and U12741 (N_12741,N_12560,N_12508);
nor U12742 (N_12742,N_12539,N_12404);
nand U12743 (N_12743,N_12415,N_12498);
nor U12744 (N_12744,N_12570,N_12579);
or U12745 (N_12745,N_12414,N_12560);
nand U12746 (N_12746,N_12514,N_12501);
nor U12747 (N_12747,N_12411,N_12507);
or U12748 (N_12748,N_12411,N_12423);
and U12749 (N_12749,N_12494,N_12518);
or U12750 (N_12750,N_12583,N_12525);
and U12751 (N_12751,N_12555,N_12450);
and U12752 (N_12752,N_12493,N_12441);
and U12753 (N_12753,N_12411,N_12485);
nor U12754 (N_12754,N_12507,N_12470);
nand U12755 (N_12755,N_12548,N_12572);
and U12756 (N_12756,N_12455,N_12573);
and U12757 (N_12757,N_12571,N_12559);
nand U12758 (N_12758,N_12432,N_12487);
and U12759 (N_12759,N_12553,N_12454);
nand U12760 (N_12760,N_12499,N_12492);
or U12761 (N_12761,N_12574,N_12563);
and U12762 (N_12762,N_12411,N_12515);
nor U12763 (N_12763,N_12510,N_12499);
or U12764 (N_12764,N_12585,N_12594);
or U12765 (N_12765,N_12454,N_12417);
or U12766 (N_12766,N_12509,N_12547);
nand U12767 (N_12767,N_12448,N_12590);
and U12768 (N_12768,N_12418,N_12523);
and U12769 (N_12769,N_12489,N_12571);
nand U12770 (N_12770,N_12430,N_12585);
or U12771 (N_12771,N_12485,N_12528);
or U12772 (N_12772,N_12484,N_12510);
nand U12773 (N_12773,N_12443,N_12454);
and U12774 (N_12774,N_12541,N_12525);
nand U12775 (N_12775,N_12524,N_12501);
nand U12776 (N_12776,N_12477,N_12485);
and U12777 (N_12777,N_12414,N_12415);
nand U12778 (N_12778,N_12430,N_12525);
or U12779 (N_12779,N_12590,N_12425);
or U12780 (N_12780,N_12479,N_12529);
nand U12781 (N_12781,N_12401,N_12532);
nor U12782 (N_12782,N_12536,N_12418);
xnor U12783 (N_12783,N_12486,N_12487);
or U12784 (N_12784,N_12554,N_12570);
and U12785 (N_12785,N_12414,N_12515);
nor U12786 (N_12786,N_12545,N_12596);
nor U12787 (N_12787,N_12568,N_12551);
nor U12788 (N_12788,N_12465,N_12526);
nand U12789 (N_12789,N_12425,N_12481);
or U12790 (N_12790,N_12575,N_12592);
or U12791 (N_12791,N_12538,N_12526);
or U12792 (N_12792,N_12424,N_12401);
or U12793 (N_12793,N_12415,N_12550);
nor U12794 (N_12794,N_12591,N_12441);
or U12795 (N_12795,N_12523,N_12463);
and U12796 (N_12796,N_12485,N_12475);
or U12797 (N_12797,N_12452,N_12454);
nor U12798 (N_12798,N_12442,N_12456);
and U12799 (N_12799,N_12575,N_12451);
or U12800 (N_12800,N_12660,N_12695);
and U12801 (N_12801,N_12664,N_12772);
and U12802 (N_12802,N_12701,N_12662);
or U12803 (N_12803,N_12793,N_12670);
and U12804 (N_12804,N_12746,N_12623);
and U12805 (N_12805,N_12784,N_12744);
or U12806 (N_12806,N_12680,N_12779);
or U12807 (N_12807,N_12745,N_12794);
or U12808 (N_12808,N_12697,N_12602);
xor U12809 (N_12809,N_12667,N_12731);
and U12810 (N_12810,N_12618,N_12620);
or U12811 (N_12811,N_12790,N_12669);
or U12812 (N_12812,N_12704,N_12648);
nand U12813 (N_12813,N_12675,N_12696);
nor U12814 (N_12814,N_12707,N_12785);
and U12815 (N_12815,N_12754,N_12774);
nor U12816 (N_12816,N_12681,N_12751);
nor U12817 (N_12817,N_12655,N_12674);
or U12818 (N_12818,N_12762,N_12702);
and U12819 (N_12819,N_12716,N_12605);
nand U12820 (N_12820,N_12758,N_12649);
or U12821 (N_12821,N_12725,N_12703);
nor U12822 (N_12822,N_12719,N_12760);
and U12823 (N_12823,N_12636,N_12615);
nor U12824 (N_12824,N_12690,N_12632);
and U12825 (N_12825,N_12673,N_12633);
nor U12826 (N_12826,N_12663,N_12645);
and U12827 (N_12827,N_12775,N_12752);
or U12828 (N_12828,N_12603,N_12611);
nand U12829 (N_12829,N_12728,N_12726);
xor U12830 (N_12830,N_12727,N_12708);
nand U12831 (N_12831,N_12769,N_12768);
or U12832 (N_12832,N_12627,N_12694);
and U12833 (N_12833,N_12640,N_12734);
nand U12834 (N_12834,N_12748,N_12770);
or U12835 (N_12835,N_12687,N_12736);
or U12836 (N_12836,N_12720,N_12616);
or U12837 (N_12837,N_12604,N_12685);
or U12838 (N_12838,N_12749,N_12786);
and U12839 (N_12839,N_12722,N_12705);
or U12840 (N_12840,N_12622,N_12607);
and U12841 (N_12841,N_12766,N_12757);
nor U12842 (N_12842,N_12796,N_12709);
nand U12843 (N_12843,N_12647,N_12672);
nor U12844 (N_12844,N_12631,N_12756);
nand U12845 (N_12845,N_12635,N_12763);
nor U12846 (N_12846,N_12706,N_12610);
nand U12847 (N_12847,N_12679,N_12630);
nor U12848 (N_12848,N_12693,N_12651);
nor U12849 (N_12849,N_12628,N_12713);
or U12850 (N_12850,N_12733,N_12743);
nor U12851 (N_12851,N_12755,N_12729);
and U12852 (N_12852,N_12776,N_12724);
and U12853 (N_12853,N_12637,N_12765);
nand U12854 (N_12854,N_12735,N_12747);
xnor U12855 (N_12855,N_12712,N_12710);
or U12856 (N_12856,N_12659,N_12606);
nor U12857 (N_12857,N_12799,N_12661);
nand U12858 (N_12858,N_12778,N_12641);
nor U12859 (N_12859,N_12617,N_12782);
xor U12860 (N_12860,N_12783,N_12797);
nand U12861 (N_12861,N_12666,N_12718);
nand U12862 (N_12862,N_12739,N_12624);
nor U12863 (N_12863,N_12759,N_12798);
xor U12864 (N_12864,N_12740,N_12665);
and U12865 (N_12865,N_12643,N_12642);
or U12866 (N_12866,N_12644,N_12625);
xnor U12867 (N_12867,N_12781,N_12717);
xor U12868 (N_12868,N_12761,N_12653);
and U12869 (N_12869,N_12609,N_12780);
nand U12870 (N_12870,N_12629,N_12753);
xor U12871 (N_12871,N_12737,N_12677);
and U12872 (N_12872,N_12683,N_12676);
nor U12873 (N_12873,N_12684,N_12771);
and U12874 (N_12874,N_12764,N_12692);
and U12875 (N_12875,N_12795,N_12721);
nor U12876 (N_12876,N_12767,N_12714);
nor U12877 (N_12877,N_12656,N_12682);
and U12878 (N_12878,N_12612,N_12671);
nand U12879 (N_12879,N_12691,N_12686);
nand U12880 (N_12880,N_12614,N_12634);
nand U12881 (N_12881,N_12698,N_12600);
xor U12882 (N_12882,N_12638,N_12613);
nor U12883 (N_12883,N_12689,N_12773);
and U12884 (N_12884,N_12668,N_12639);
or U12885 (N_12885,N_12787,N_12741);
and U12886 (N_12886,N_12715,N_12738);
nor U12887 (N_12887,N_12646,N_12723);
nand U12888 (N_12888,N_12688,N_12788);
and U12889 (N_12889,N_12608,N_12789);
nor U12890 (N_12890,N_12742,N_12654);
nand U12891 (N_12891,N_12650,N_12619);
and U12892 (N_12892,N_12791,N_12750);
nand U12893 (N_12893,N_12626,N_12652);
and U12894 (N_12894,N_12657,N_12792);
and U12895 (N_12895,N_12700,N_12711);
nor U12896 (N_12896,N_12732,N_12678);
and U12897 (N_12897,N_12621,N_12730);
nor U12898 (N_12898,N_12777,N_12601);
and U12899 (N_12899,N_12699,N_12658);
nand U12900 (N_12900,N_12667,N_12797);
or U12901 (N_12901,N_12654,N_12745);
and U12902 (N_12902,N_12791,N_12701);
nor U12903 (N_12903,N_12670,N_12791);
and U12904 (N_12904,N_12772,N_12749);
or U12905 (N_12905,N_12602,N_12705);
nand U12906 (N_12906,N_12749,N_12630);
nand U12907 (N_12907,N_12638,N_12617);
and U12908 (N_12908,N_12649,N_12738);
or U12909 (N_12909,N_12763,N_12688);
nand U12910 (N_12910,N_12616,N_12756);
nor U12911 (N_12911,N_12777,N_12739);
or U12912 (N_12912,N_12702,N_12691);
or U12913 (N_12913,N_12774,N_12683);
nor U12914 (N_12914,N_12667,N_12745);
nand U12915 (N_12915,N_12726,N_12645);
and U12916 (N_12916,N_12689,N_12730);
nand U12917 (N_12917,N_12723,N_12608);
nor U12918 (N_12918,N_12624,N_12670);
nand U12919 (N_12919,N_12788,N_12767);
xor U12920 (N_12920,N_12654,N_12705);
xnor U12921 (N_12921,N_12653,N_12639);
nor U12922 (N_12922,N_12697,N_12660);
nor U12923 (N_12923,N_12742,N_12630);
or U12924 (N_12924,N_12607,N_12796);
nor U12925 (N_12925,N_12708,N_12731);
and U12926 (N_12926,N_12663,N_12789);
and U12927 (N_12927,N_12608,N_12695);
or U12928 (N_12928,N_12648,N_12651);
nor U12929 (N_12929,N_12622,N_12710);
xor U12930 (N_12930,N_12742,N_12789);
nor U12931 (N_12931,N_12668,N_12723);
and U12932 (N_12932,N_12694,N_12685);
nand U12933 (N_12933,N_12612,N_12605);
nor U12934 (N_12934,N_12784,N_12614);
or U12935 (N_12935,N_12676,N_12687);
and U12936 (N_12936,N_12640,N_12762);
nand U12937 (N_12937,N_12790,N_12767);
and U12938 (N_12938,N_12723,N_12730);
and U12939 (N_12939,N_12716,N_12743);
nand U12940 (N_12940,N_12621,N_12627);
nor U12941 (N_12941,N_12630,N_12600);
xor U12942 (N_12942,N_12689,N_12789);
nor U12943 (N_12943,N_12677,N_12725);
nor U12944 (N_12944,N_12603,N_12766);
or U12945 (N_12945,N_12799,N_12654);
or U12946 (N_12946,N_12621,N_12789);
nand U12947 (N_12947,N_12728,N_12747);
or U12948 (N_12948,N_12621,N_12769);
and U12949 (N_12949,N_12695,N_12605);
or U12950 (N_12950,N_12652,N_12616);
nand U12951 (N_12951,N_12680,N_12653);
nor U12952 (N_12952,N_12755,N_12769);
and U12953 (N_12953,N_12638,N_12722);
and U12954 (N_12954,N_12782,N_12778);
nor U12955 (N_12955,N_12637,N_12688);
nand U12956 (N_12956,N_12769,N_12676);
nor U12957 (N_12957,N_12641,N_12625);
or U12958 (N_12958,N_12617,N_12756);
nand U12959 (N_12959,N_12666,N_12610);
and U12960 (N_12960,N_12792,N_12687);
and U12961 (N_12961,N_12728,N_12664);
or U12962 (N_12962,N_12717,N_12606);
or U12963 (N_12963,N_12609,N_12781);
xnor U12964 (N_12964,N_12604,N_12765);
nor U12965 (N_12965,N_12735,N_12648);
nand U12966 (N_12966,N_12711,N_12771);
or U12967 (N_12967,N_12695,N_12777);
or U12968 (N_12968,N_12720,N_12697);
and U12969 (N_12969,N_12665,N_12624);
or U12970 (N_12970,N_12701,N_12611);
and U12971 (N_12971,N_12726,N_12752);
or U12972 (N_12972,N_12780,N_12649);
and U12973 (N_12973,N_12762,N_12759);
xor U12974 (N_12974,N_12719,N_12619);
nor U12975 (N_12975,N_12650,N_12796);
and U12976 (N_12976,N_12772,N_12660);
nor U12977 (N_12977,N_12757,N_12796);
nand U12978 (N_12978,N_12783,N_12688);
or U12979 (N_12979,N_12711,N_12657);
and U12980 (N_12980,N_12673,N_12753);
xnor U12981 (N_12981,N_12741,N_12734);
and U12982 (N_12982,N_12733,N_12695);
and U12983 (N_12983,N_12607,N_12762);
nor U12984 (N_12984,N_12647,N_12606);
nand U12985 (N_12985,N_12701,N_12643);
nand U12986 (N_12986,N_12684,N_12615);
nor U12987 (N_12987,N_12604,N_12706);
nand U12988 (N_12988,N_12717,N_12777);
and U12989 (N_12989,N_12703,N_12701);
nand U12990 (N_12990,N_12696,N_12739);
or U12991 (N_12991,N_12791,N_12685);
and U12992 (N_12992,N_12690,N_12672);
and U12993 (N_12993,N_12672,N_12664);
nand U12994 (N_12994,N_12723,N_12712);
nor U12995 (N_12995,N_12709,N_12622);
or U12996 (N_12996,N_12700,N_12671);
nand U12997 (N_12997,N_12747,N_12650);
nor U12998 (N_12998,N_12623,N_12730);
nor U12999 (N_12999,N_12706,N_12791);
nor U13000 (N_13000,N_12826,N_12810);
nor U13001 (N_13001,N_12925,N_12914);
and U13002 (N_13002,N_12905,N_12968);
or U13003 (N_13003,N_12845,N_12937);
nor U13004 (N_13004,N_12900,N_12913);
and U13005 (N_13005,N_12917,N_12827);
or U13006 (N_13006,N_12870,N_12805);
xnor U13007 (N_13007,N_12950,N_12813);
nand U13008 (N_13008,N_12976,N_12971);
nand U13009 (N_13009,N_12985,N_12880);
xnor U13010 (N_13010,N_12938,N_12876);
and U13011 (N_13011,N_12801,N_12850);
xnor U13012 (N_13012,N_12919,N_12903);
and U13013 (N_13013,N_12871,N_12918);
or U13014 (N_13014,N_12869,N_12910);
or U13015 (N_13015,N_12947,N_12970);
and U13016 (N_13016,N_12853,N_12811);
xor U13017 (N_13017,N_12906,N_12885);
nand U13018 (N_13018,N_12806,N_12819);
xor U13019 (N_13019,N_12888,N_12804);
and U13020 (N_13020,N_12974,N_12941);
or U13021 (N_13021,N_12933,N_12896);
nand U13022 (N_13022,N_12955,N_12998);
nand U13023 (N_13023,N_12835,N_12808);
or U13024 (N_13024,N_12832,N_12883);
and U13025 (N_13025,N_12908,N_12857);
nor U13026 (N_13026,N_12829,N_12833);
and U13027 (N_13027,N_12861,N_12856);
nand U13028 (N_13028,N_12800,N_12996);
nand U13029 (N_13029,N_12915,N_12864);
or U13030 (N_13030,N_12939,N_12866);
nor U13031 (N_13031,N_12989,N_12958);
or U13032 (N_13032,N_12803,N_12844);
nor U13033 (N_13033,N_12959,N_12840);
or U13034 (N_13034,N_12993,N_12886);
nand U13035 (N_13035,N_12843,N_12821);
or U13036 (N_13036,N_12868,N_12863);
and U13037 (N_13037,N_12994,N_12949);
nor U13038 (N_13038,N_12975,N_12940);
nor U13039 (N_13039,N_12930,N_12807);
and U13040 (N_13040,N_12839,N_12894);
or U13041 (N_13041,N_12922,N_12890);
nand U13042 (N_13042,N_12904,N_12924);
nor U13043 (N_13043,N_12809,N_12892);
and U13044 (N_13044,N_12935,N_12847);
and U13045 (N_13045,N_12846,N_12838);
xnor U13046 (N_13046,N_12928,N_12972);
nor U13047 (N_13047,N_12872,N_12875);
and U13048 (N_13048,N_12934,N_12945);
and U13049 (N_13049,N_12952,N_12860);
and U13050 (N_13050,N_12884,N_12907);
nor U13051 (N_13051,N_12966,N_12814);
nor U13052 (N_13052,N_12921,N_12891);
or U13053 (N_13053,N_12957,N_12862);
or U13054 (N_13054,N_12902,N_12920);
nor U13055 (N_13055,N_12916,N_12977);
nand U13056 (N_13056,N_12817,N_12927);
nand U13057 (N_13057,N_12995,N_12983);
or U13058 (N_13058,N_12901,N_12893);
nor U13059 (N_13059,N_12967,N_12960);
nor U13060 (N_13060,N_12987,N_12963);
nand U13061 (N_13061,N_12887,N_12858);
nor U13062 (N_13062,N_12943,N_12848);
or U13063 (N_13063,N_12841,N_12831);
xor U13064 (N_13064,N_12836,N_12988);
or U13065 (N_13065,N_12978,N_12823);
and U13066 (N_13066,N_12951,N_12855);
nor U13067 (N_13067,N_12881,N_12992);
nand U13068 (N_13068,N_12877,N_12997);
nand U13069 (N_13069,N_12873,N_12944);
and U13070 (N_13070,N_12911,N_12936);
nor U13071 (N_13071,N_12802,N_12874);
and U13072 (N_13072,N_12969,N_12820);
xor U13073 (N_13073,N_12953,N_12825);
or U13074 (N_13074,N_12984,N_12912);
xor U13075 (N_13075,N_12923,N_12946);
nand U13076 (N_13076,N_12942,N_12956);
and U13077 (N_13077,N_12834,N_12859);
nand U13078 (N_13078,N_12982,N_12898);
nand U13079 (N_13079,N_12929,N_12954);
xor U13080 (N_13080,N_12986,N_12981);
nand U13081 (N_13081,N_12897,N_12849);
nand U13082 (N_13082,N_12879,N_12909);
and U13083 (N_13083,N_12822,N_12815);
or U13084 (N_13084,N_12948,N_12889);
nor U13085 (N_13085,N_12818,N_12999);
nand U13086 (N_13086,N_12965,N_12842);
and U13087 (N_13087,N_12812,N_12854);
and U13088 (N_13088,N_12878,N_12932);
nand U13089 (N_13089,N_12931,N_12979);
or U13090 (N_13090,N_12828,N_12980);
nand U13091 (N_13091,N_12824,N_12962);
nor U13092 (N_13092,N_12961,N_12991);
and U13093 (N_13093,N_12964,N_12899);
or U13094 (N_13094,N_12990,N_12867);
or U13095 (N_13095,N_12926,N_12816);
nand U13096 (N_13096,N_12837,N_12830);
nand U13097 (N_13097,N_12973,N_12852);
nand U13098 (N_13098,N_12851,N_12882);
and U13099 (N_13099,N_12895,N_12865);
and U13100 (N_13100,N_12960,N_12835);
or U13101 (N_13101,N_12874,N_12885);
nor U13102 (N_13102,N_12992,N_12988);
nand U13103 (N_13103,N_12948,N_12885);
nand U13104 (N_13104,N_12966,N_12897);
and U13105 (N_13105,N_12835,N_12814);
xnor U13106 (N_13106,N_12847,N_12853);
and U13107 (N_13107,N_12863,N_12838);
xnor U13108 (N_13108,N_12881,N_12962);
or U13109 (N_13109,N_12870,N_12900);
nor U13110 (N_13110,N_12975,N_12841);
or U13111 (N_13111,N_12867,N_12969);
or U13112 (N_13112,N_12854,N_12800);
nor U13113 (N_13113,N_12975,N_12812);
or U13114 (N_13114,N_12961,N_12850);
or U13115 (N_13115,N_12956,N_12941);
or U13116 (N_13116,N_12997,N_12975);
and U13117 (N_13117,N_12966,N_12939);
or U13118 (N_13118,N_12961,N_12951);
nand U13119 (N_13119,N_12851,N_12855);
or U13120 (N_13120,N_12819,N_12970);
and U13121 (N_13121,N_12855,N_12813);
xnor U13122 (N_13122,N_12939,N_12945);
and U13123 (N_13123,N_12857,N_12995);
and U13124 (N_13124,N_12977,N_12831);
and U13125 (N_13125,N_12856,N_12831);
nand U13126 (N_13126,N_12827,N_12806);
nand U13127 (N_13127,N_12875,N_12957);
and U13128 (N_13128,N_12988,N_12814);
or U13129 (N_13129,N_12925,N_12878);
or U13130 (N_13130,N_12956,N_12931);
or U13131 (N_13131,N_12942,N_12802);
or U13132 (N_13132,N_12990,N_12807);
nor U13133 (N_13133,N_12814,N_12934);
nor U13134 (N_13134,N_12833,N_12998);
nor U13135 (N_13135,N_12856,N_12898);
xnor U13136 (N_13136,N_12889,N_12809);
nor U13137 (N_13137,N_12824,N_12879);
and U13138 (N_13138,N_12883,N_12971);
and U13139 (N_13139,N_12819,N_12992);
xor U13140 (N_13140,N_12992,N_12925);
nor U13141 (N_13141,N_12967,N_12856);
nand U13142 (N_13142,N_12934,N_12835);
and U13143 (N_13143,N_12936,N_12855);
or U13144 (N_13144,N_12897,N_12808);
nor U13145 (N_13145,N_12816,N_12823);
and U13146 (N_13146,N_12896,N_12891);
xor U13147 (N_13147,N_12831,N_12917);
or U13148 (N_13148,N_12837,N_12865);
nor U13149 (N_13149,N_12870,N_12841);
nand U13150 (N_13150,N_12814,N_12847);
and U13151 (N_13151,N_12841,N_12912);
nor U13152 (N_13152,N_12864,N_12943);
xor U13153 (N_13153,N_12824,N_12942);
or U13154 (N_13154,N_12821,N_12950);
or U13155 (N_13155,N_12934,N_12844);
nand U13156 (N_13156,N_12978,N_12848);
and U13157 (N_13157,N_12922,N_12867);
or U13158 (N_13158,N_12916,N_12998);
nand U13159 (N_13159,N_12984,N_12800);
xnor U13160 (N_13160,N_12884,N_12888);
and U13161 (N_13161,N_12877,N_12889);
and U13162 (N_13162,N_12879,N_12939);
nand U13163 (N_13163,N_12824,N_12834);
nand U13164 (N_13164,N_12863,N_12913);
and U13165 (N_13165,N_12960,N_12819);
nand U13166 (N_13166,N_12895,N_12959);
nor U13167 (N_13167,N_12800,N_12915);
xor U13168 (N_13168,N_12805,N_12997);
nor U13169 (N_13169,N_12941,N_12981);
nor U13170 (N_13170,N_12999,N_12814);
nand U13171 (N_13171,N_12960,N_12933);
and U13172 (N_13172,N_12888,N_12941);
nor U13173 (N_13173,N_12922,N_12985);
xnor U13174 (N_13174,N_12956,N_12977);
nand U13175 (N_13175,N_12946,N_12907);
or U13176 (N_13176,N_12889,N_12899);
xor U13177 (N_13177,N_12936,N_12853);
or U13178 (N_13178,N_12888,N_12909);
nor U13179 (N_13179,N_12943,N_12891);
and U13180 (N_13180,N_12800,N_12863);
xnor U13181 (N_13181,N_12979,N_12959);
nor U13182 (N_13182,N_12989,N_12860);
nand U13183 (N_13183,N_12972,N_12957);
and U13184 (N_13184,N_12823,N_12831);
nor U13185 (N_13185,N_12932,N_12832);
nand U13186 (N_13186,N_12877,N_12837);
xor U13187 (N_13187,N_12940,N_12914);
and U13188 (N_13188,N_12944,N_12865);
and U13189 (N_13189,N_12858,N_12862);
nand U13190 (N_13190,N_12896,N_12860);
or U13191 (N_13191,N_12885,N_12922);
or U13192 (N_13192,N_12804,N_12966);
nor U13193 (N_13193,N_12955,N_12819);
and U13194 (N_13194,N_12842,N_12959);
nand U13195 (N_13195,N_12821,N_12966);
nor U13196 (N_13196,N_12976,N_12944);
nor U13197 (N_13197,N_12913,N_12931);
nand U13198 (N_13198,N_12895,N_12844);
and U13199 (N_13199,N_12987,N_12919);
and U13200 (N_13200,N_13193,N_13124);
and U13201 (N_13201,N_13049,N_13003);
nand U13202 (N_13202,N_13079,N_13121);
and U13203 (N_13203,N_13103,N_13132);
xnor U13204 (N_13204,N_13141,N_13192);
nand U13205 (N_13205,N_13001,N_13101);
and U13206 (N_13206,N_13061,N_13034);
and U13207 (N_13207,N_13028,N_13188);
xor U13208 (N_13208,N_13063,N_13070);
nor U13209 (N_13209,N_13097,N_13140);
nor U13210 (N_13210,N_13168,N_13176);
or U13211 (N_13211,N_13081,N_13004);
nand U13212 (N_13212,N_13156,N_13020);
nand U13213 (N_13213,N_13045,N_13091);
nor U13214 (N_13214,N_13119,N_13096);
xor U13215 (N_13215,N_13105,N_13137);
or U13216 (N_13216,N_13163,N_13051);
xnor U13217 (N_13217,N_13050,N_13012);
or U13218 (N_13218,N_13133,N_13185);
nand U13219 (N_13219,N_13148,N_13073);
xnor U13220 (N_13220,N_13026,N_13112);
or U13221 (N_13221,N_13082,N_13042);
nand U13222 (N_13222,N_13074,N_13167);
and U13223 (N_13223,N_13136,N_13144);
nand U13224 (N_13224,N_13077,N_13066);
or U13225 (N_13225,N_13002,N_13175);
and U13226 (N_13226,N_13009,N_13098);
nand U13227 (N_13227,N_13099,N_13019);
nand U13228 (N_13228,N_13169,N_13102);
xnor U13229 (N_13229,N_13094,N_13014);
and U13230 (N_13230,N_13198,N_13147);
nand U13231 (N_13231,N_13106,N_13052);
xor U13232 (N_13232,N_13111,N_13044);
or U13233 (N_13233,N_13040,N_13037);
xnor U13234 (N_13234,N_13100,N_13021);
and U13235 (N_13235,N_13115,N_13065);
nor U13236 (N_13236,N_13010,N_13158);
and U13237 (N_13237,N_13022,N_13161);
nor U13238 (N_13238,N_13143,N_13076);
or U13239 (N_13239,N_13181,N_13125);
and U13240 (N_13240,N_13157,N_13071);
nor U13241 (N_13241,N_13183,N_13129);
xnor U13242 (N_13242,N_13197,N_13109);
nand U13243 (N_13243,N_13131,N_13114);
nand U13244 (N_13244,N_13007,N_13038);
nand U13245 (N_13245,N_13023,N_13146);
nand U13246 (N_13246,N_13060,N_13083);
xnor U13247 (N_13247,N_13011,N_13152);
or U13248 (N_13248,N_13191,N_13172);
nand U13249 (N_13249,N_13015,N_13027);
or U13250 (N_13250,N_13118,N_13090);
nand U13251 (N_13251,N_13180,N_13159);
xor U13252 (N_13252,N_13029,N_13033);
or U13253 (N_13253,N_13024,N_13128);
nor U13254 (N_13254,N_13092,N_13174);
nand U13255 (N_13255,N_13043,N_13187);
or U13256 (N_13256,N_13107,N_13178);
nor U13257 (N_13257,N_13093,N_13186);
nand U13258 (N_13258,N_13108,N_13134);
nand U13259 (N_13259,N_13113,N_13046);
and U13260 (N_13260,N_13095,N_13057);
nor U13261 (N_13261,N_13032,N_13030);
nand U13262 (N_13262,N_13122,N_13075);
or U13263 (N_13263,N_13058,N_13005);
or U13264 (N_13264,N_13035,N_13155);
or U13265 (N_13265,N_13055,N_13126);
and U13266 (N_13266,N_13160,N_13116);
xor U13267 (N_13267,N_13054,N_13170);
or U13268 (N_13268,N_13138,N_13025);
and U13269 (N_13269,N_13031,N_13120);
and U13270 (N_13270,N_13036,N_13072);
and U13271 (N_13271,N_13067,N_13130);
nor U13272 (N_13272,N_13069,N_13041);
nand U13273 (N_13273,N_13123,N_13047);
xor U13274 (N_13274,N_13048,N_13062);
nand U13275 (N_13275,N_13056,N_13086);
and U13276 (N_13276,N_13196,N_13078);
nand U13277 (N_13277,N_13135,N_13087);
and U13278 (N_13278,N_13127,N_13084);
nand U13279 (N_13279,N_13199,N_13165);
nand U13280 (N_13280,N_13142,N_13166);
and U13281 (N_13281,N_13064,N_13184);
and U13282 (N_13282,N_13190,N_13117);
or U13283 (N_13283,N_13189,N_13177);
nand U13284 (N_13284,N_13059,N_13089);
nor U13285 (N_13285,N_13194,N_13018);
or U13286 (N_13286,N_13173,N_13039);
or U13287 (N_13287,N_13013,N_13080);
or U13288 (N_13288,N_13179,N_13139);
nand U13289 (N_13289,N_13164,N_13171);
xor U13290 (N_13290,N_13068,N_13053);
nor U13291 (N_13291,N_13182,N_13016);
nand U13292 (N_13292,N_13104,N_13088);
nand U13293 (N_13293,N_13195,N_13085);
nor U13294 (N_13294,N_13008,N_13006);
or U13295 (N_13295,N_13145,N_13110);
nand U13296 (N_13296,N_13154,N_13000);
nand U13297 (N_13297,N_13162,N_13149);
nor U13298 (N_13298,N_13151,N_13153);
or U13299 (N_13299,N_13150,N_13017);
nand U13300 (N_13300,N_13062,N_13033);
and U13301 (N_13301,N_13021,N_13067);
xnor U13302 (N_13302,N_13031,N_13100);
nor U13303 (N_13303,N_13035,N_13024);
nor U13304 (N_13304,N_13082,N_13159);
and U13305 (N_13305,N_13041,N_13193);
and U13306 (N_13306,N_13006,N_13130);
and U13307 (N_13307,N_13150,N_13108);
and U13308 (N_13308,N_13182,N_13164);
xnor U13309 (N_13309,N_13181,N_13197);
nand U13310 (N_13310,N_13002,N_13130);
nor U13311 (N_13311,N_13027,N_13090);
and U13312 (N_13312,N_13091,N_13134);
nor U13313 (N_13313,N_13120,N_13189);
nand U13314 (N_13314,N_13188,N_13186);
and U13315 (N_13315,N_13014,N_13056);
or U13316 (N_13316,N_13096,N_13125);
or U13317 (N_13317,N_13087,N_13079);
nand U13318 (N_13318,N_13165,N_13033);
or U13319 (N_13319,N_13007,N_13103);
and U13320 (N_13320,N_13124,N_13194);
nand U13321 (N_13321,N_13084,N_13090);
xnor U13322 (N_13322,N_13197,N_13152);
nor U13323 (N_13323,N_13115,N_13166);
nor U13324 (N_13324,N_13123,N_13043);
and U13325 (N_13325,N_13083,N_13119);
and U13326 (N_13326,N_13160,N_13114);
or U13327 (N_13327,N_13180,N_13114);
nor U13328 (N_13328,N_13018,N_13094);
xor U13329 (N_13329,N_13088,N_13159);
xnor U13330 (N_13330,N_13075,N_13147);
or U13331 (N_13331,N_13135,N_13076);
nand U13332 (N_13332,N_13119,N_13134);
nand U13333 (N_13333,N_13086,N_13043);
or U13334 (N_13334,N_13103,N_13015);
nand U13335 (N_13335,N_13168,N_13146);
xnor U13336 (N_13336,N_13047,N_13131);
nor U13337 (N_13337,N_13115,N_13124);
nand U13338 (N_13338,N_13111,N_13039);
nor U13339 (N_13339,N_13046,N_13129);
xor U13340 (N_13340,N_13123,N_13112);
nor U13341 (N_13341,N_13048,N_13112);
nand U13342 (N_13342,N_13020,N_13083);
and U13343 (N_13343,N_13192,N_13080);
or U13344 (N_13344,N_13076,N_13139);
nor U13345 (N_13345,N_13107,N_13118);
nor U13346 (N_13346,N_13037,N_13029);
nand U13347 (N_13347,N_13114,N_13164);
xor U13348 (N_13348,N_13009,N_13167);
nor U13349 (N_13349,N_13027,N_13127);
nand U13350 (N_13350,N_13175,N_13125);
nor U13351 (N_13351,N_13003,N_13112);
nor U13352 (N_13352,N_13143,N_13065);
or U13353 (N_13353,N_13152,N_13160);
nand U13354 (N_13354,N_13102,N_13017);
and U13355 (N_13355,N_13112,N_13152);
and U13356 (N_13356,N_13183,N_13142);
or U13357 (N_13357,N_13182,N_13028);
or U13358 (N_13358,N_13131,N_13092);
nor U13359 (N_13359,N_13117,N_13173);
nor U13360 (N_13360,N_13075,N_13080);
xnor U13361 (N_13361,N_13159,N_13127);
nand U13362 (N_13362,N_13121,N_13187);
nand U13363 (N_13363,N_13141,N_13171);
nand U13364 (N_13364,N_13084,N_13188);
or U13365 (N_13365,N_13144,N_13171);
nor U13366 (N_13366,N_13168,N_13117);
xnor U13367 (N_13367,N_13054,N_13107);
nand U13368 (N_13368,N_13149,N_13119);
or U13369 (N_13369,N_13105,N_13164);
or U13370 (N_13370,N_13090,N_13059);
or U13371 (N_13371,N_13077,N_13018);
nor U13372 (N_13372,N_13005,N_13186);
xnor U13373 (N_13373,N_13035,N_13159);
or U13374 (N_13374,N_13017,N_13090);
and U13375 (N_13375,N_13045,N_13030);
nor U13376 (N_13376,N_13188,N_13101);
nor U13377 (N_13377,N_13055,N_13031);
xor U13378 (N_13378,N_13173,N_13186);
nor U13379 (N_13379,N_13163,N_13153);
nor U13380 (N_13380,N_13158,N_13063);
and U13381 (N_13381,N_13046,N_13146);
or U13382 (N_13382,N_13198,N_13077);
xnor U13383 (N_13383,N_13157,N_13115);
or U13384 (N_13384,N_13049,N_13160);
xor U13385 (N_13385,N_13107,N_13132);
and U13386 (N_13386,N_13043,N_13176);
nand U13387 (N_13387,N_13099,N_13098);
or U13388 (N_13388,N_13131,N_13178);
nand U13389 (N_13389,N_13052,N_13030);
nand U13390 (N_13390,N_13071,N_13042);
or U13391 (N_13391,N_13141,N_13183);
or U13392 (N_13392,N_13131,N_13080);
nor U13393 (N_13393,N_13061,N_13012);
xnor U13394 (N_13394,N_13017,N_13182);
nand U13395 (N_13395,N_13103,N_13183);
and U13396 (N_13396,N_13040,N_13020);
nor U13397 (N_13397,N_13139,N_13157);
nor U13398 (N_13398,N_13155,N_13199);
and U13399 (N_13399,N_13186,N_13135);
nand U13400 (N_13400,N_13310,N_13223);
xnor U13401 (N_13401,N_13317,N_13233);
and U13402 (N_13402,N_13354,N_13361);
nand U13403 (N_13403,N_13259,N_13242);
or U13404 (N_13404,N_13371,N_13243);
nor U13405 (N_13405,N_13398,N_13325);
or U13406 (N_13406,N_13397,N_13230);
xor U13407 (N_13407,N_13318,N_13357);
xnor U13408 (N_13408,N_13258,N_13239);
nand U13409 (N_13409,N_13313,N_13200);
and U13410 (N_13410,N_13294,N_13399);
and U13411 (N_13411,N_13215,N_13329);
and U13412 (N_13412,N_13382,N_13358);
nor U13413 (N_13413,N_13342,N_13207);
nand U13414 (N_13414,N_13285,N_13348);
xor U13415 (N_13415,N_13331,N_13302);
or U13416 (N_13416,N_13349,N_13224);
or U13417 (N_13417,N_13336,N_13221);
nand U13418 (N_13418,N_13332,N_13216);
and U13419 (N_13419,N_13250,N_13328);
nor U13420 (N_13420,N_13205,N_13312);
or U13421 (N_13421,N_13376,N_13295);
nand U13422 (N_13422,N_13375,N_13365);
xnor U13423 (N_13423,N_13235,N_13238);
and U13424 (N_13424,N_13248,N_13340);
nor U13425 (N_13425,N_13395,N_13222);
nand U13426 (N_13426,N_13229,N_13268);
and U13427 (N_13427,N_13262,N_13299);
nand U13428 (N_13428,N_13347,N_13300);
or U13429 (N_13429,N_13290,N_13335);
nand U13430 (N_13430,N_13297,N_13373);
xor U13431 (N_13431,N_13351,N_13372);
nor U13432 (N_13432,N_13355,N_13341);
or U13433 (N_13433,N_13293,N_13392);
or U13434 (N_13434,N_13324,N_13280);
and U13435 (N_13435,N_13385,N_13226);
nor U13436 (N_13436,N_13284,N_13287);
or U13437 (N_13437,N_13319,N_13209);
or U13438 (N_13438,N_13327,N_13273);
nor U13439 (N_13439,N_13288,N_13366);
nor U13440 (N_13440,N_13247,N_13265);
xor U13441 (N_13441,N_13387,N_13277);
and U13442 (N_13442,N_13256,N_13345);
nand U13443 (N_13443,N_13218,N_13343);
nor U13444 (N_13444,N_13263,N_13374);
xor U13445 (N_13445,N_13260,N_13278);
xnor U13446 (N_13446,N_13307,N_13379);
and U13447 (N_13447,N_13234,N_13369);
and U13448 (N_13448,N_13384,N_13344);
and U13449 (N_13449,N_13305,N_13241);
nand U13450 (N_13450,N_13314,N_13252);
nor U13451 (N_13451,N_13326,N_13352);
xnor U13452 (N_13452,N_13396,N_13338);
nand U13453 (N_13453,N_13362,N_13270);
nor U13454 (N_13454,N_13323,N_13311);
nand U13455 (N_13455,N_13289,N_13266);
and U13456 (N_13456,N_13237,N_13292);
or U13457 (N_13457,N_13279,N_13272);
and U13458 (N_13458,N_13322,N_13334);
or U13459 (N_13459,N_13367,N_13274);
nor U13460 (N_13460,N_13206,N_13346);
nand U13461 (N_13461,N_13308,N_13208);
nand U13462 (N_13462,N_13315,N_13388);
and U13463 (N_13463,N_13244,N_13219);
nor U13464 (N_13464,N_13304,N_13390);
and U13465 (N_13465,N_13282,N_13225);
xor U13466 (N_13466,N_13231,N_13381);
nand U13467 (N_13467,N_13283,N_13337);
nor U13468 (N_13468,N_13202,N_13303);
or U13469 (N_13469,N_13321,N_13394);
and U13470 (N_13470,N_13261,N_13350);
nor U13471 (N_13471,N_13320,N_13201);
nor U13472 (N_13472,N_13377,N_13333);
nor U13473 (N_13473,N_13217,N_13236);
xnor U13474 (N_13474,N_13214,N_13378);
and U13475 (N_13475,N_13301,N_13339);
nor U13476 (N_13476,N_13253,N_13356);
xnor U13477 (N_13477,N_13276,N_13353);
and U13478 (N_13478,N_13271,N_13255);
nand U13479 (N_13479,N_13227,N_13240);
nor U13480 (N_13480,N_13264,N_13286);
or U13481 (N_13481,N_13281,N_13296);
nor U13482 (N_13482,N_13386,N_13275);
nor U13483 (N_13483,N_13306,N_13212);
and U13484 (N_13484,N_13210,N_13211);
nor U13485 (N_13485,N_13368,N_13359);
or U13486 (N_13486,N_13393,N_13298);
or U13487 (N_13487,N_13232,N_13257);
nand U13488 (N_13488,N_13391,N_13251);
or U13489 (N_13489,N_13383,N_13254);
and U13490 (N_13490,N_13245,N_13364);
or U13491 (N_13491,N_13269,N_13316);
nor U13492 (N_13492,N_13360,N_13228);
or U13493 (N_13493,N_13246,N_13363);
and U13494 (N_13494,N_13203,N_13267);
nand U13495 (N_13495,N_13291,N_13309);
nand U13496 (N_13496,N_13389,N_13370);
and U13497 (N_13497,N_13380,N_13249);
nor U13498 (N_13498,N_13330,N_13213);
and U13499 (N_13499,N_13220,N_13204);
or U13500 (N_13500,N_13397,N_13358);
and U13501 (N_13501,N_13208,N_13219);
nor U13502 (N_13502,N_13200,N_13357);
nor U13503 (N_13503,N_13204,N_13239);
nor U13504 (N_13504,N_13262,N_13210);
xnor U13505 (N_13505,N_13376,N_13226);
nor U13506 (N_13506,N_13242,N_13299);
and U13507 (N_13507,N_13311,N_13224);
nand U13508 (N_13508,N_13336,N_13360);
or U13509 (N_13509,N_13326,N_13341);
and U13510 (N_13510,N_13212,N_13238);
nor U13511 (N_13511,N_13322,N_13332);
or U13512 (N_13512,N_13224,N_13203);
nand U13513 (N_13513,N_13241,N_13251);
and U13514 (N_13514,N_13330,N_13223);
nor U13515 (N_13515,N_13381,N_13326);
and U13516 (N_13516,N_13238,N_13305);
and U13517 (N_13517,N_13389,N_13387);
xor U13518 (N_13518,N_13239,N_13379);
nor U13519 (N_13519,N_13390,N_13381);
nand U13520 (N_13520,N_13360,N_13306);
xor U13521 (N_13521,N_13362,N_13250);
and U13522 (N_13522,N_13354,N_13252);
or U13523 (N_13523,N_13200,N_13327);
nand U13524 (N_13524,N_13363,N_13236);
and U13525 (N_13525,N_13327,N_13250);
nor U13526 (N_13526,N_13212,N_13357);
xnor U13527 (N_13527,N_13209,N_13346);
nand U13528 (N_13528,N_13298,N_13216);
nand U13529 (N_13529,N_13211,N_13295);
and U13530 (N_13530,N_13355,N_13255);
and U13531 (N_13531,N_13231,N_13262);
nand U13532 (N_13532,N_13251,N_13216);
xor U13533 (N_13533,N_13210,N_13369);
nand U13534 (N_13534,N_13311,N_13274);
and U13535 (N_13535,N_13374,N_13370);
nor U13536 (N_13536,N_13228,N_13369);
and U13537 (N_13537,N_13210,N_13206);
nand U13538 (N_13538,N_13310,N_13358);
nor U13539 (N_13539,N_13237,N_13305);
nor U13540 (N_13540,N_13326,N_13208);
or U13541 (N_13541,N_13350,N_13338);
and U13542 (N_13542,N_13217,N_13368);
or U13543 (N_13543,N_13201,N_13251);
or U13544 (N_13544,N_13237,N_13218);
nor U13545 (N_13545,N_13299,N_13388);
and U13546 (N_13546,N_13216,N_13367);
or U13547 (N_13547,N_13285,N_13230);
nor U13548 (N_13548,N_13359,N_13224);
xor U13549 (N_13549,N_13226,N_13290);
or U13550 (N_13550,N_13278,N_13378);
nor U13551 (N_13551,N_13295,N_13207);
and U13552 (N_13552,N_13253,N_13368);
or U13553 (N_13553,N_13330,N_13338);
nand U13554 (N_13554,N_13397,N_13282);
nand U13555 (N_13555,N_13240,N_13314);
nand U13556 (N_13556,N_13281,N_13386);
nor U13557 (N_13557,N_13370,N_13292);
nand U13558 (N_13558,N_13330,N_13391);
nand U13559 (N_13559,N_13226,N_13341);
or U13560 (N_13560,N_13302,N_13285);
nor U13561 (N_13561,N_13208,N_13293);
nand U13562 (N_13562,N_13213,N_13277);
and U13563 (N_13563,N_13367,N_13353);
and U13564 (N_13564,N_13216,N_13312);
or U13565 (N_13565,N_13277,N_13214);
and U13566 (N_13566,N_13258,N_13224);
and U13567 (N_13567,N_13302,N_13374);
or U13568 (N_13568,N_13313,N_13269);
or U13569 (N_13569,N_13345,N_13229);
and U13570 (N_13570,N_13318,N_13323);
and U13571 (N_13571,N_13236,N_13344);
xor U13572 (N_13572,N_13293,N_13204);
or U13573 (N_13573,N_13378,N_13339);
nor U13574 (N_13574,N_13278,N_13389);
nand U13575 (N_13575,N_13347,N_13340);
and U13576 (N_13576,N_13252,N_13375);
xnor U13577 (N_13577,N_13364,N_13278);
nand U13578 (N_13578,N_13258,N_13223);
xnor U13579 (N_13579,N_13382,N_13335);
xnor U13580 (N_13580,N_13338,N_13270);
or U13581 (N_13581,N_13311,N_13371);
or U13582 (N_13582,N_13312,N_13239);
nand U13583 (N_13583,N_13224,N_13264);
or U13584 (N_13584,N_13338,N_13300);
nor U13585 (N_13585,N_13366,N_13226);
xor U13586 (N_13586,N_13203,N_13336);
xor U13587 (N_13587,N_13302,N_13268);
or U13588 (N_13588,N_13251,N_13323);
or U13589 (N_13589,N_13389,N_13305);
nand U13590 (N_13590,N_13333,N_13375);
xor U13591 (N_13591,N_13369,N_13286);
nand U13592 (N_13592,N_13399,N_13381);
or U13593 (N_13593,N_13358,N_13355);
or U13594 (N_13594,N_13298,N_13232);
and U13595 (N_13595,N_13302,N_13259);
or U13596 (N_13596,N_13342,N_13383);
and U13597 (N_13597,N_13217,N_13230);
nor U13598 (N_13598,N_13220,N_13322);
nand U13599 (N_13599,N_13310,N_13287);
or U13600 (N_13600,N_13438,N_13505);
or U13601 (N_13601,N_13516,N_13409);
nor U13602 (N_13602,N_13506,N_13496);
and U13603 (N_13603,N_13486,N_13418);
and U13604 (N_13604,N_13469,N_13594);
or U13605 (N_13605,N_13568,N_13540);
and U13606 (N_13606,N_13487,N_13404);
nor U13607 (N_13607,N_13500,N_13453);
nor U13608 (N_13608,N_13546,N_13435);
nand U13609 (N_13609,N_13517,N_13544);
nor U13610 (N_13610,N_13592,N_13455);
and U13611 (N_13611,N_13530,N_13518);
and U13612 (N_13612,N_13548,N_13482);
or U13613 (N_13613,N_13556,N_13541);
nand U13614 (N_13614,N_13531,N_13470);
nor U13615 (N_13615,N_13533,N_13590);
or U13616 (N_13616,N_13429,N_13471);
or U13617 (N_13617,N_13468,N_13412);
nand U13618 (N_13618,N_13492,N_13450);
or U13619 (N_13619,N_13581,N_13422);
and U13620 (N_13620,N_13465,N_13423);
nor U13621 (N_13621,N_13413,N_13573);
nor U13622 (N_13622,N_13431,N_13575);
nand U13623 (N_13623,N_13499,N_13428);
xor U13624 (N_13624,N_13558,N_13561);
nand U13625 (N_13625,N_13459,N_13443);
nor U13626 (N_13626,N_13447,N_13501);
or U13627 (N_13627,N_13521,N_13572);
nand U13628 (N_13628,N_13585,N_13439);
nor U13629 (N_13629,N_13485,N_13483);
xnor U13630 (N_13630,N_13513,N_13508);
or U13631 (N_13631,N_13547,N_13400);
nor U13632 (N_13632,N_13491,N_13557);
nor U13633 (N_13633,N_13444,N_13597);
or U13634 (N_13634,N_13526,N_13466);
nand U13635 (N_13635,N_13522,N_13566);
nand U13636 (N_13636,N_13514,N_13420);
nand U13637 (N_13637,N_13542,N_13570);
or U13638 (N_13638,N_13454,N_13552);
or U13639 (N_13639,N_13523,N_13583);
nor U13640 (N_13640,N_13574,N_13586);
and U13641 (N_13641,N_13416,N_13555);
xor U13642 (N_13642,N_13445,N_13545);
and U13643 (N_13643,N_13562,N_13576);
nor U13644 (N_13644,N_13419,N_13587);
nor U13645 (N_13645,N_13589,N_13451);
or U13646 (N_13646,N_13503,N_13571);
and U13647 (N_13647,N_13569,N_13509);
nor U13648 (N_13648,N_13473,N_13430);
nand U13649 (N_13649,N_13560,N_13515);
and U13650 (N_13650,N_13593,N_13577);
or U13651 (N_13651,N_13414,N_13563);
nor U13652 (N_13652,N_13446,N_13584);
xor U13653 (N_13653,N_13474,N_13528);
and U13654 (N_13654,N_13452,N_13421);
or U13655 (N_13655,N_13426,N_13478);
and U13656 (N_13656,N_13539,N_13488);
and U13657 (N_13657,N_13417,N_13472);
and U13658 (N_13658,N_13489,N_13565);
and U13659 (N_13659,N_13549,N_13437);
nor U13660 (N_13660,N_13507,N_13424);
nand U13661 (N_13661,N_13525,N_13476);
nor U13662 (N_13662,N_13405,N_13462);
or U13663 (N_13663,N_13534,N_13588);
xnor U13664 (N_13664,N_13432,N_13407);
and U13665 (N_13665,N_13564,N_13578);
nor U13666 (N_13666,N_13463,N_13458);
nor U13667 (N_13667,N_13553,N_13519);
nor U13668 (N_13668,N_13442,N_13490);
or U13669 (N_13669,N_13464,N_13480);
or U13670 (N_13670,N_13411,N_13406);
and U13671 (N_13671,N_13498,N_13538);
nand U13672 (N_13672,N_13477,N_13520);
nand U13673 (N_13673,N_13402,N_13559);
nand U13674 (N_13674,N_13427,N_13497);
xnor U13675 (N_13675,N_13460,N_13536);
xnor U13676 (N_13676,N_13479,N_13410);
nor U13677 (N_13677,N_13449,N_13448);
or U13678 (N_13678,N_13403,N_13510);
and U13679 (N_13679,N_13512,N_13524);
and U13680 (N_13680,N_13537,N_13425);
and U13681 (N_13681,N_13495,N_13433);
nor U13682 (N_13682,N_13551,N_13527);
or U13683 (N_13683,N_13582,N_13461);
nor U13684 (N_13684,N_13554,N_13596);
nor U13685 (N_13685,N_13599,N_13401);
nor U13686 (N_13686,N_13467,N_13550);
or U13687 (N_13687,N_13502,N_13493);
and U13688 (N_13688,N_13504,N_13595);
or U13689 (N_13689,N_13580,N_13567);
nand U13690 (N_13690,N_13543,N_13484);
nor U13691 (N_13691,N_13535,N_13441);
and U13692 (N_13692,N_13591,N_13494);
nand U13693 (N_13693,N_13457,N_13579);
nand U13694 (N_13694,N_13532,N_13475);
xnor U13695 (N_13695,N_13436,N_13456);
nor U13696 (N_13696,N_13440,N_13529);
and U13697 (N_13697,N_13481,N_13434);
nor U13698 (N_13698,N_13415,N_13408);
nor U13699 (N_13699,N_13511,N_13598);
nand U13700 (N_13700,N_13529,N_13562);
and U13701 (N_13701,N_13573,N_13475);
nor U13702 (N_13702,N_13479,N_13482);
nor U13703 (N_13703,N_13426,N_13472);
xor U13704 (N_13704,N_13425,N_13436);
and U13705 (N_13705,N_13557,N_13587);
nor U13706 (N_13706,N_13495,N_13487);
nand U13707 (N_13707,N_13401,N_13494);
and U13708 (N_13708,N_13425,N_13533);
nor U13709 (N_13709,N_13551,N_13454);
nand U13710 (N_13710,N_13560,N_13492);
and U13711 (N_13711,N_13472,N_13464);
or U13712 (N_13712,N_13558,N_13559);
nand U13713 (N_13713,N_13515,N_13595);
and U13714 (N_13714,N_13452,N_13459);
and U13715 (N_13715,N_13440,N_13464);
and U13716 (N_13716,N_13591,N_13477);
nor U13717 (N_13717,N_13507,N_13552);
nand U13718 (N_13718,N_13429,N_13458);
nor U13719 (N_13719,N_13541,N_13416);
or U13720 (N_13720,N_13582,N_13534);
xnor U13721 (N_13721,N_13563,N_13561);
nand U13722 (N_13722,N_13513,N_13569);
and U13723 (N_13723,N_13569,N_13486);
nand U13724 (N_13724,N_13577,N_13446);
and U13725 (N_13725,N_13411,N_13421);
nor U13726 (N_13726,N_13563,N_13498);
nor U13727 (N_13727,N_13427,N_13465);
and U13728 (N_13728,N_13492,N_13520);
xnor U13729 (N_13729,N_13486,N_13402);
nand U13730 (N_13730,N_13508,N_13584);
and U13731 (N_13731,N_13559,N_13485);
or U13732 (N_13732,N_13530,N_13523);
nand U13733 (N_13733,N_13401,N_13504);
or U13734 (N_13734,N_13462,N_13427);
nand U13735 (N_13735,N_13587,N_13420);
or U13736 (N_13736,N_13460,N_13526);
or U13737 (N_13737,N_13495,N_13448);
and U13738 (N_13738,N_13444,N_13534);
or U13739 (N_13739,N_13578,N_13544);
xor U13740 (N_13740,N_13510,N_13464);
nand U13741 (N_13741,N_13572,N_13493);
or U13742 (N_13742,N_13414,N_13428);
xnor U13743 (N_13743,N_13580,N_13550);
nand U13744 (N_13744,N_13525,N_13591);
nor U13745 (N_13745,N_13448,N_13461);
nor U13746 (N_13746,N_13526,N_13473);
or U13747 (N_13747,N_13499,N_13517);
nor U13748 (N_13748,N_13456,N_13552);
and U13749 (N_13749,N_13459,N_13585);
nor U13750 (N_13750,N_13565,N_13562);
nor U13751 (N_13751,N_13436,N_13495);
nor U13752 (N_13752,N_13564,N_13581);
and U13753 (N_13753,N_13409,N_13440);
or U13754 (N_13754,N_13499,N_13504);
or U13755 (N_13755,N_13547,N_13582);
nor U13756 (N_13756,N_13546,N_13404);
nand U13757 (N_13757,N_13523,N_13495);
nor U13758 (N_13758,N_13486,N_13450);
and U13759 (N_13759,N_13427,N_13535);
nand U13760 (N_13760,N_13458,N_13449);
nand U13761 (N_13761,N_13519,N_13509);
nor U13762 (N_13762,N_13464,N_13413);
and U13763 (N_13763,N_13435,N_13472);
nor U13764 (N_13764,N_13531,N_13422);
or U13765 (N_13765,N_13551,N_13425);
or U13766 (N_13766,N_13409,N_13507);
nand U13767 (N_13767,N_13501,N_13449);
xor U13768 (N_13768,N_13435,N_13421);
nand U13769 (N_13769,N_13490,N_13448);
nand U13770 (N_13770,N_13503,N_13461);
nor U13771 (N_13771,N_13488,N_13425);
or U13772 (N_13772,N_13466,N_13431);
or U13773 (N_13773,N_13401,N_13564);
or U13774 (N_13774,N_13521,N_13440);
and U13775 (N_13775,N_13590,N_13451);
and U13776 (N_13776,N_13558,N_13576);
nand U13777 (N_13777,N_13418,N_13516);
or U13778 (N_13778,N_13513,N_13524);
xor U13779 (N_13779,N_13565,N_13524);
or U13780 (N_13780,N_13474,N_13402);
and U13781 (N_13781,N_13417,N_13402);
nand U13782 (N_13782,N_13409,N_13432);
and U13783 (N_13783,N_13565,N_13529);
or U13784 (N_13784,N_13554,N_13454);
nand U13785 (N_13785,N_13509,N_13566);
and U13786 (N_13786,N_13584,N_13447);
or U13787 (N_13787,N_13540,N_13485);
nor U13788 (N_13788,N_13480,N_13408);
nor U13789 (N_13789,N_13576,N_13520);
and U13790 (N_13790,N_13568,N_13498);
nand U13791 (N_13791,N_13566,N_13469);
nand U13792 (N_13792,N_13447,N_13577);
nor U13793 (N_13793,N_13439,N_13521);
nor U13794 (N_13794,N_13511,N_13442);
nor U13795 (N_13795,N_13560,N_13481);
nand U13796 (N_13796,N_13532,N_13564);
nand U13797 (N_13797,N_13485,N_13403);
and U13798 (N_13798,N_13491,N_13550);
or U13799 (N_13799,N_13507,N_13458);
and U13800 (N_13800,N_13743,N_13768);
nor U13801 (N_13801,N_13697,N_13717);
nand U13802 (N_13802,N_13617,N_13691);
nor U13803 (N_13803,N_13765,N_13660);
nand U13804 (N_13804,N_13781,N_13608);
nor U13805 (N_13805,N_13622,N_13642);
nand U13806 (N_13806,N_13764,N_13686);
or U13807 (N_13807,N_13737,N_13751);
and U13808 (N_13808,N_13723,N_13650);
and U13809 (N_13809,N_13710,N_13770);
xor U13810 (N_13810,N_13644,N_13756);
and U13811 (N_13811,N_13782,N_13614);
xor U13812 (N_13812,N_13610,N_13663);
or U13813 (N_13813,N_13706,N_13783);
xnor U13814 (N_13814,N_13739,N_13772);
or U13815 (N_13815,N_13613,N_13602);
nand U13816 (N_13816,N_13604,N_13621);
and U13817 (N_13817,N_13678,N_13605);
nand U13818 (N_13818,N_13734,N_13716);
and U13819 (N_13819,N_13626,N_13759);
and U13820 (N_13820,N_13679,N_13667);
xor U13821 (N_13821,N_13703,N_13777);
or U13822 (N_13822,N_13636,N_13714);
nand U13823 (N_13823,N_13767,N_13701);
or U13824 (N_13824,N_13646,N_13662);
nand U13825 (N_13825,N_13790,N_13740);
nor U13826 (N_13826,N_13769,N_13713);
xnor U13827 (N_13827,N_13784,N_13623);
or U13828 (N_13828,N_13773,N_13688);
and U13829 (N_13829,N_13631,N_13612);
nor U13830 (N_13830,N_13653,N_13632);
nor U13831 (N_13831,N_13661,N_13620);
or U13832 (N_13832,N_13752,N_13685);
xnor U13833 (N_13833,N_13648,N_13721);
and U13834 (N_13834,N_13651,N_13793);
xor U13835 (N_13835,N_13615,N_13635);
nor U13836 (N_13836,N_13624,N_13641);
nand U13837 (N_13837,N_13733,N_13600);
and U13838 (N_13838,N_13744,N_13758);
or U13839 (N_13839,N_13796,N_13746);
nand U13840 (N_13840,N_13687,N_13748);
nand U13841 (N_13841,N_13698,N_13780);
or U13842 (N_13842,N_13702,N_13666);
or U13843 (N_13843,N_13729,N_13724);
nor U13844 (N_13844,N_13647,N_13619);
nor U13845 (N_13845,N_13634,N_13618);
xnor U13846 (N_13846,N_13616,N_13704);
and U13847 (N_13847,N_13637,N_13794);
nand U13848 (N_13848,N_13774,N_13639);
and U13849 (N_13849,N_13673,N_13786);
or U13850 (N_13850,N_13779,N_13690);
nor U13851 (N_13851,N_13699,N_13700);
and U13852 (N_13852,N_13655,N_13625);
or U13853 (N_13853,N_13730,N_13665);
or U13854 (N_13854,N_13692,N_13785);
or U13855 (N_13855,N_13749,N_13657);
or U13856 (N_13856,N_13681,N_13775);
and U13857 (N_13857,N_13683,N_13771);
and U13858 (N_13858,N_13638,N_13603);
nor U13859 (N_13859,N_13719,N_13671);
and U13860 (N_13860,N_13684,N_13672);
nand U13861 (N_13861,N_13761,N_13643);
xor U13862 (N_13862,N_13725,N_13720);
nor U13863 (N_13863,N_13736,N_13694);
or U13864 (N_13864,N_13726,N_13633);
nor U13865 (N_13865,N_13664,N_13677);
or U13866 (N_13866,N_13670,N_13652);
or U13867 (N_13867,N_13735,N_13680);
and U13868 (N_13868,N_13718,N_13727);
or U13869 (N_13869,N_13715,N_13728);
nor U13870 (N_13870,N_13731,N_13674);
and U13871 (N_13871,N_13762,N_13747);
nand U13872 (N_13872,N_13776,N_13745);
or U13873 (N_13873,N_13629,N_13755);
and U13874 (N_13874,N_13792,N_13709);
and U13875 (N_13875,N_13738,N_13675);
nand U13876 (N_13876,N_13787,N_13645);
xor U13877 (N_13877,N_13695,N_13753);
xnor U13878 (N_13878,N_13696,N_13611);
nand U13879 (N_13879,N_13640,N_13750);
nand U13880 (N_13880,N_13705,N_13654);
nand U13881 (N_13881,N_13627,N_13742);
xor U13882 (N_13882,N_13693,N_13760);
and U13883 (N_13883,N_13682,N_13630);
and U13884 (N_13884,N_13668,N_13656);
or U13885 (N_13885,N_13708,N_13711);
xnor U13886 (N_13886,N_13795,N_13766);
or U13887 (N_13887,N_13676,N_13788);
or U13888 (N_13888,N_13669,N_13628);
xor U13889 (N_13889,N_13799,N_13658);
nor U13890 (N_13890,N_13757,N_13754);
nor U13891 (N_13891,N_13659,N_13689);
nand U13892 (N_13892,N_13732,N_13712);
nand U13893 (N_13893,N_13722,N_13791);
nor U13894 (N_13894,N_13798,N_13778);
nor U13895 (N_13895,N_13601,N_13763);
and U13896 (N_13896,N_13789,N_13741);
and U13897 (N_13897,N_13649,N_13707);
and U13898 (N_13898,N_13609,N_13607);
or U13899 (N_13899,N_13797,N_13606);
nand U13900 (N_13900,N_13630,N_13776);
nand U13901 (N_13901,N_13695,N_13701);
xor U13902 (N_13902,N_13763,N_13778);
or U13903 (N_13903,N_13683,N_13702);
nand U13904 (N_13904,N_13641,N_13794);
or U13905 (N_13905,N_13743,N_13698);
nand U13906 (N_13906,N_13642,N_13746);
and U13907 (N_13907,N_13796,N_13734);
and U13908 (N_13908,N_13763,N_13797);
and U13909 (N_13909,N_13631,N_13680);
and U13910 (N_13910,N_13789,N_13673);
nand U13911 (N_13911,N_13784,N_13633);
and U13912 (N_13912,N_13776,N_13705);
nand U13913 (N_13913,N_13772,N_13734);
xor U13914 (N_13914,N_13674,N_13772);
nor U13915 (N_13915,N_13652,N_13660);
nand U13916 (N_13916,N_13710,N_13776);
nor U13917 (N_13917,N_13741,N_13793);
or U13918 (N_13918,N_13696,N_13751);
or U13919 (N_13919,N_13729,N_13787);
and U13920 (N_13920,N_13639,N_13699);
nor U13921 (N_13921,N_13794,N_13625);
and U13922 (N_13922,N_13604,N_13719);
and U13923 (N_13923,N_13799,N_13772);
nand U13924 (N_13924,N_13698,N_13694);
nor U13925 (N_13925,N_13765,N_13729);
nand U13926 (N_13926,N_13650,N_13670);
and U13927 (N_13927,N_13658,N_13738);
or U13928 (N_13928,N_13749,N_13717);
nor U13929 (N_13929,N_13638,N_13657);
nor U13930 (N_13930,N_13749,N_13625);
nor U13931 (N_13931,N_13799,N_13627);
or U13932 (N_13932,N_13772,N_13764);
nor U13933 (N_13933,N_13620,N_13785);
xor U13934 (N_13934,N_13688,N_13633);
or U13935 (N_13935,N_13600,N_13744);
or U13936 (N_13936,N_13793,N_13780);
or U13937 (N_13937,N_13757,N_13689);
nor U13938 (N_13938,N_13745,N_13733);
nor U13939 (N_13939,N_13770,N_13641);
xnor U13940 (N_13940,N_13604,N_13794);
or U13941 (N_13941,N_13763,N_13757);
nor U13942 (N_13942,N_13787,N_13604);
nor U13943 (N_13943,N_13795,N_13784);
nand U13944 (N_13944,N_13692,N_13626);
nand U13945 (N_13945,N_13756,N_13648);
nand U13946 (N_13946,N_13718,N_13761);
nand U13947 (N_13947,N_13651,N_13678);
nor U13948 (N_13948,N_13604,N_13622);
or U13949 (N_13949,N_13650,N_13688);
nor U13950 (N_13950,N_13762,N_13772);
nor U13951 (N_13951,N_13766,N_13698);
nand U13952 (N_13952,N_13680,N_13697);
or U13953 (N_13953,N_13636,N_13791);
or U13954 (N_13954,N_13752,N_13636);
or U13955 (N_13955,N_13790,N_13744);
and U13956 (N_13956,N_13725,N_13721);
or U13957 (N_13957,N_13786,N_13663);
nand U13958 (N_13958,N_13744,N_13666);
and U13959 (N_13959,N_13682,N_13688);
nor U13960 (N_13960,N_13638,N_13769);
xor U13961 (N_13961,N_13668,N_13619);
nor U13962 (N_13962,N_13729,N_13763);
nand U13963 (N_13963,N_13679,N_13639);
and U13964 (N_13964,N_13737,N_13620);
nand U13965 (N_13965,N_13734,N_13754);
nor U13966 (N_13966,N_13625,N_13720);
and U13967 (N_13967,N_13737,N_13789);
nor U13968 (N_13968,N_13606,N_13687);
nor U13969 (N_13969,N_13678,N_13765);
or U13970 (N_13970,N_13708,N_13778);
or U13971 (N_13971,N_13611,N_13762);
and U13972 (N_13972,N_13710,N_13735);
nor U13973 (N_13973,N_13718,N_13701);
and U13974 (N_13974,N_13756,N_13799);
nor U13975 (N_13975,N_13687,N_13647);
nor U13976 (N_13976,N_13759,N_13779);
nand U13977 (N_13977,N_13741,N_13636);
nand U13978 (N_13978,N_13714,N_13653);
and U13979 (N_13979,N_13739,N_13653);
nand U13980 (N_13980,N_13792,N_13725);
nand U13981 (N_13981,N_13790,N_13742);
and U13982 (N_13982,N_13772,N_13735);
nor U13983 (N_13983,N_13756,N_13638);
and U13984 (N_13984,N_13738,N_13712);
nand U13985 (N_13985,N_13713,N_13665);
and U13986 (N_13986,N_13787,N_13733);
nor U13987 (N_13987,N_13674,N_13736);
nand U13988 (N_13988,N_13664,N_13652);
and U13989 (N_13989,N_13729,N_13726);
xnor U13990 (N_13990,N_13734,N_13700);
and U13991 (N_13991,N_13648,N_13711);
and U13992 (N_13992,N_13749,N_13771);
or U13993 (N_13993,N_13651,N_13650);
or U13994 (N_13994,N_13766,N_13739);
nand U13995 (N_13995,N_13774,N_13730);
and U13996 (N_13996,N_13627,N_13673);
nor U13997 (N_13997,N_13656,N_13754);
nand U13998 (N_13998,N_13752,N_13719);
or U13999 (N_13999,N_13770,N_13667);
nand U14000 (N_14000,N_13940,N_13947);
or U14001 (N_14001,N_13876,N_13815);
or U14002 (N_14002,N_13859,N_13971);
nor U14003 (N_14003,N_13908,N_13872);
and U14004 (N_14004,N_13902,N_13897);
and U14005 (N_14005,N_13893,N_13868);
xnor U14006 (N_14006,N_13853,N_13927);
or U14007 (N_14007,N_13914,N_13923);
or U14008 (N_14008,N_13874,N_13968);
nand U14009 (N_14009,N_13836,N_13953);
nand U14010 (N_14010,N_13888,N_13926);
nor U14011 (N_14011,N_13941,N_13986);
xor U14012 (N_14012,N_13809,N_13921);
and U14013 (N_14013,N_13974,N_13913);
nand U14014 (N_14014,N_13866,N_13989);
nand U14015 (N_14015,N_13826,N_13991);
nor U14016 (N_14016,N_13831,N_13969);
and U14017 (N_14017,N_13845,N_13867);
nand U14018 (N_14018,N_13945,N_13892);
or U14019 (N_14019,N_13808,N_13838);
and U14020 (N_14020,N_13988,N_13973);
and U14021 (N_14021,N_13822,N_13857);
or U14022 (N_14022,N_13871,N_13824);
nand U14023 (N_14023,N_13807,N_13967);
or U14024 (N_14024,N_13832,N_13855);
and U14025 (N_14025,N_13978,N_13932);
and U14026 (N_14026,N_13950,N_13802);
nand U14027 (N_14027,N_13865,N_13919);
or U14028 (N_14028,N_13964,N_13870);
and U14029 (N_14029,N_13999,N_13825);
or U14030 (N_14030,N_13891,N_13957);
or U14031 (N_14031,N_13970,N_13886);
and U14032 (N_14032,N_13800,N_13931);
nand U14033 (N_14033,N_13849,N_13814);
or U14034 (N_14034,N_13875,N_13883);
or U14035 (N_14035,N_13905,N_13909);
nand U14036 (N_14036,N_13803,N_13965);
nor U14037 (N_14037,N_13985,N_13984);
xor U14038 (N_14038,N_13930,N_13918);
xor U14039 (N_14039,N_13920,N_13887);
and U14040 (N_14040,N_13976,N_13804);
nor U14041 (N_14041,N_13966,N_13995);
nand U14042 (N_14042,N_13858,N_13860);
nand U14043 (N_14043,N_13980,N_13917);
nand U14044 (N_14044,N_13959,N_13934);
nor U14045 (N_14045,N_13882,N_13951);
nand U14046 (N_14046,N_13958,N_13827);
and U14047 (N_14047,N_13801,N_13901);
nor U14048 (N_14048,N_13904,N_13990);
and U14049 (N_14049,N_13937,N_13873);
nand U14050 (N_14050,N_13847,N_13933);
xor U14051 (N_14051,N_13850,N_13906);
xnor U14052 (N_14052,N_13811,N_13963);
nand U14053 (N_14053,N_13997,N_13936);
nand U14054 (N_14054,N_13916,N_13810);
nand U14055 (N_14055,N_13813,N_13885);
nor U14056 (N_14056,N_13992,N_13983);
and U14057 (N_14057,N_13907,N_13977);
or U14058 (N_14058,N_13856,N_13818);
or U14059 (N_14059,N_13928,N_13828);
nor U14060 (N_14060,N_13924,N_13946);
or U14061 (N_14061,N_13929,N_13889);
nand U14062 (N_14062,N_13880,N_13829);
and U14063 (N_14063,N_13846,N_13837);
and U14064 (N_14064,N_13996,N_13962);
nand U14065 (N_14065,N_13839,N_13993);
or U14066 (N_14066,N_13833,N_13884);
or U14067 (N_14067,N_13938,N_13806);
nor U14068 (N_14068,N_13981,N_13841);
nor U14069 (N_14069,N_13915,N_13979);
nand U14070 (N_14070,N_13954,N_13942);
nor U14071 (N_14071,N_13840,N_13817);
xor U14072 (N_14072,N_13948,N_13987);
nor U14073 (N_14073,N_13943,N_13949);
or U14074 (N_14074,N_13972,N_13898);
or U14075 (N_14075,N_13844,N_13922);
nand U14076 (N_14076,N_13820,N_13812);
or U14077 (N_14077,N_13869,N_13834);
and U14078 (N_14078,N_13955,N_13911);
nand U14079 (N_14079,N_13903,N_13994);
xor U14080 (N_14080,N_13935,N_13896);
and U14081 (N_14081,N_13830,N_13819);
or U14082 (N_14082,N_13881,N_13961);
or U14083 (N_14083,N_13900,N_13952);
nand U14084 (N_14084,N_13877,N_13848);
and U14085 (N_14085,N_13899,N_13852);
and U14086 (N_14086,N_13925,N_13975);
nor U14087 (N_14087,N_13956,N_13960);
xnor U14088 (N_14088,N_13861,N_13998);
nand U14089 (N_14089,N_13851,N_13912);
nand U14090 (N_14090,N_13879,N_13842);
nor U14091 (N_14091,N_13805,N_13878);
nor U14092 (N_14092,N_13982,N_13843);
and U14093 (N_14093,N_13939,N_13835);
and U14094 (N_14094,N_13863,N_13895);
nand U14095 (N_14095,N_13816,N_13944);
nand U14096 (N_14096,N_13821,N_13910);
and U14097 (N_14097,N_13823,N_13862);
or U14098 (N_14098,N_13854,N_13894);
or U14099 (N_14099,N_13864,N_13890);
and U14100 (N_14100,N_13942,N_13849);
and U14101 (N_14101,N_13829,N_13989);
xor U14102 (N_14102,N_13840,N_13998);
and U14103 (N_14103,N_13938,N_13819);
nor U14104 (N_14104,N_13825,N_13918);
nand U14105 (N_14105,N_13901,N_13963);
nand U14106 (N_14106,N_13955,N_13870);
or U14107 (N_14107,N_13934,N_13984);
and U14108 (N_14108,N_13899,N_13814);
nand U14109 (N_14109,N_13921,N_13817);
and U14110 (N_14110,N_13807,N_13879);
nand U14111 (N_14111,N_13915,N_13949);
and U14112 (N_14112,N_13918,N_13824);
and U14113 (N_14113,N_13959,N_13994);
nor U14114 (N_14114,N_13814,N_13852);
xnor U14115 (N_14115,N_13932,N_13895);
nand U14116 (N_14116,N_13963,N_13945);
xnor U14117 (N_14117,N_13936,N_13972);
and U14118 (N_14118,N_13871,N_13957);
or U14119 (N_14119,N_13960,N_13936);
nor U14120 (N_14120,N_13821,N_13859);
nand U14121 (N_14121,N_13825,N_13949);
or U14122 (N_14122,N_13914,N_13992);
or U14123 (N_14123,N_13814,N_13920);
nor U14124 (N_14124,N_13855,N_13953);
and U14125 (N_14125,N_13855,N_13999);
nand U14126 (N_14126,N_13839,N_13862);
nor U14127 (N_14127,N_13950,N_13966);
nand U14128 (N_14128,N_13870,N_13927);
nor U14129 (N_14129,N_13995,N_13881);
and U14130 (N_14130,N_13945,N_13815);
nand U14131 (N_14131,N_13916,N_13971);
or U14132 (N_14132,N_13944,N_13945);
nor U14133 (N_14133,N_13970,N_13871);
xnor U14134 (N_14134,N_13990,N_13932);
and U14135 (N_14135,N_13967,N_13869);
nand U14136 (N_14136,N_13819,N_13927);
nor U14137 (N_14137,N_13960,N_13884);
nor U14138 (N_14138,N_13896,N_13938);
or U14139 (N_14139,N_13933,N_13945);
xor U14140 (N_14140,N_13866,N_13865);
nand U14141 (N_14141,N_13896,N_13937);
nand U14142 (N_14142,N_13965,N_13958);
and U14143 (N_14143,N_13970,N_13881);
and U14144 (N_14144,N_13931,N_13965);
and U14145 (N_14145,N_13993,N_13863);
and U14146 (N_14146,N_13956,N_13839);
and U14147 (N_14147,N_13960,N_13969);
nand U14148 (N_14148,N_13873,N_13823);
xnor U14149 (N_14149,N_13987,N_13908);
and U14150 (N_14150,N_13942,N_13903);
or U14151 (N_14151,N_13924,N_13893);
and U14152 (N_14152,N_13840,N_13802);
nor U14153 (N_14153,N_13963,N_13919);
nand U14154 (N_14154,N_13866,N_13877);
nand U14155 (N_14155,N_13930,N_13801);
xor U14156 (N_14156,N_13979,N_13810);
xor U14157 (N_14157,N_13800,N_13914);
and U14158 (N_14158,N_13936,N_13925);
xor U14159 (N_14159,N_13919,N_13888);
nand U14160 (N_14160,N_13998,N_13891);
nor U14161 (N_14161,N_13976,N_13999);
nor U14162 (N_14162,N_13958,N_13890);
or U14163 (N_14163,N_13850,N_13848);
or U14164 (N_14164,N_13845,N_13898);
or U14165 (N_14165,N_13859,N_13989);
and U14166 (N_14166,N_13874,N_13994);
nor U14167 (N_14167,N_13932,N_13925);
nand U14168 (N_14168,N_13940,N_13989);
nand U14169 (N_14169,N_13968,N_13848);
nand U14170 (N_14170,N_13862,N_13832);
and U14171 (N_14171,N_13891,N_13945);
xor U14172 (N_14172,N_13963,N_13809);
nand U14173 (N_14173,N_13995,N_13917);
or U14174 (N_14174,N_13993,N_13974);
nor U14175 (N_14175,N_13974,N_13971);
or U14176 (N_14176,N_13971,N_13980);
xor U14177 (N_14177,N_13850,N_13933);
or U14178 (N_14178,N_13980,N_13895);
or U14179 (N_14179,N_13837,N_13835);
or U14180 (N_14180,N_13907,N_13866);
and U14181 (N_14181,N_13946,N_13983);
nor U14182 (N_14182,N_13888,N_13869);
and U14183 (N_14183,N_13858,N_13953);
nand U14184 (N_14184,N_13892,N_13881);
or U14185 (N_14185,N_13853,N_13900);
nand U14186 (N_14186,N_13899,N_13905);
nor U14187 (N_14187,N_13920,N_13931);
xor U14188 (N_14188,N_13892,N_13862);
nor U14189 (N_14189,N_13923,N_13979);
nand U14190 (N_14190,N_13943,N_13802);
or U14191 (N_14191,N_13809,N_13827);
or U14192 (N_14192,N_13917,N_13894);
nand U14193 (N_14193,N_13894,N_13922);
and U14194 (N_14194,N_13994,N_13901);
nand U14195 (N_14195,N_13856,N_13872);
and U14196 (N_14196,N_13818,N_13842);
nand U14197 (N_14197,N_13843,N_13845);
or U14198 (N_14198,N_13923,N_13910);
nand U14199 (N_14199,N_13926,N_13863);
and U14200 (N_14200,N_14149,N_14014);
and U14201 (N_14201,N_14167,N_14151);
nand U14202 (N_14202,N_14063,N_14035);
nand U14203 (N_14203,N_14124,N_14138);
nand U14204 (N_14204,N_14017,N_14182);
and U14205 (N_14205,N_14085,N_14026);
nand U14206 (N_14206,N_14199,N_14005);
or U14207 (N_14207,N_14052,N_14039);
nand U14208 (N_14208,N_14018,N_14171);
nor U14209 (N_14209,N_14133,N_14053);
xnor U14210 (N_14210,N_14075,N_14148);
or U14211 (N_14211,N_14033,N_14082);
or U14212 (N_14212,N_14008,N_14094);
or U14213 (N_14213,N_14025,N_14143);
xor U14214 (N_14214,N_14144,N_14037);
nor U14215 (N_14215,N_14046,N_14131);
or U14216 (N_14216,N_14040,N_14066);
or U14217 (N_14217,N_14024,N_14150);
nand U14218 (N_14218,N_14006,N_14166);
nor U14219 (N_14219,N_14173,N_14176);
and U14220 (N_14220,N_14194,N_14095);
nand U14221 (N_14221,N_14165,N_14136);
and U14222 (N_14222,N_14177,N_14135);
or U14223 (N_14223,N_14071,N_14047);
nor U14224 (N_14224,N_14129,N_14105);
nand U14225 (N_14225,N_14057,N_14032);
nor U14226 (N_14226,N_14019,N_14116);
nor U14227 (N_14227,N_14020,N_14043);
nand U14228 (N_14228,N_14181,N_14141);
and U14229 (N_14229,N_14193,N_14098);
nand U14230 (N_14230,N_14108,N_14041);
and U14231 (N_14231,N_14190,N_14107);
and U14232 (N_14232,N_14048,N_14086);
nor U14233 (N_14233,N_14178,N_14013);
and U14234 (N_14234,N_14023,N_14139);
nor U14235 (N_14235,N_14186,N_14092);
nor U14236 (N_14236,N_14076,N_14004);
nand U14237 (N_14237,N_14029,N_14187);
and U14238 (N_14238,N_14134,N_14093);
or U14239 (N_14239,N_14100,N_14115);
xnor U14240 (N_14240,N_14189,N_14103);
xor U14241 (N_14241,N_14049,N_14123);
xnor U14242 (N_14242,N_14090,N_14036);
or U14243 (N_14243,N_14003,N_14021);
and U14244 (N_14244,N_14045,N_14031);
nor U14245 (N_14245,N_14120,N_14101);
or U14246 (N_14246,N_14169,N_14089);
and U14247 (N_14247,N_14059,N_14130);
nor U14248 (N_14248,N_14154,N_14172);
and U14249 (N_14249,N_14081,N_14099);
and U14250 (N_14250,N_14077,N_14125);
nand U14251 (N_14251,N_14027,N_14113);
nor U14252 (N_14252,N_14011,N_14002);
or U14253 (N_14253,N_14001,N_14010);
and U14254 (N_14254,N_14067,N_14126);
or U14255 (N_14255,N_14028,N_14104);
and U14256 (N_14256,N_14112,N_14078);
and U14257 (N_14257,N_14137,N_14000);
or U14258 (N_14258,N_14110,N_14069);
or U14259 (N_14259,N_14087,N_14161);
nand U14260 (N_14260,N_14064,N_14160);
or U14261 (N_14261,N_14097,N_14163);
nor U14262 (N_14262,N_14157,N_14179);
and U14263 (N_14263,N_14196,N_14128);
or U14264 (N_14264,N_14073,N_14121);
and U14265 (N_14265,N_14184,N_14195);
xnor U14266 (N_14266,N_14061,N_14088);
nand U14267 (N_14267,N_14117,N_14058);
nor U14268 (N_14268,N_14192,N_14170);
or U14269 (N_14269,N_14106,N_14044);
nor U14270 (N_14270,N_14091,N_14162);
xor U14271 (N_14271,N_14015,N_14072);
and U14272 (N_14272,N_14152,N_14083);
nand U14273 (N_14273,N_14198,N_14132);
or U14274 (N_14274,N_14175,N_14142);
and U14275 (N_14275,N_14119,N_14188);
xor U14276 (N_14276,N_14185,N_14109);
nor U14277 (N_14277,N_14146,N_14158);
nor U14278 (N_14278,N_14096,N_14145);
nand U14279 (N_14279,N_14016,N_14084);
xor U14280 (N_14280,N_14012,N_14114);
xnor U14281 (N_14281,N_14156,N_14168);
nand U14282 (N_14282,N_14007,N_14056);
xnor U14283 (N_14283,N_14065,N_14155);
and U14284 (N_14284,N_14060,N_14127);
nor U14285 (N_14285,N_14111,N_14055);
or U14286 (N_14286,N_14034,N_14054);
or U14287 (N_14287,N_14180,N_14118);
and U14288 (N_14288,N_14050,N_14042);
nand U14289 (N_14289,N_14038,N_14197);
and U14290 (N_14290,N_14122,N_14147);
and U14291 (N_14291,N_14079,N_14164);
or U14292 (N_14292,N_14030,N_14074);
or U14293 (N_14293,N_14051,N_14009);
xnor U14294 (N_14294,N_14062,N_14140);
nand U14295 (N_14295,N_14068,N_14102);
or U14296 (N_14296,N_14174,N_14022);
nand U14297 (N_14297,N_14183,N_14080);
or U14298 (N_14298,N_14191,N_14070);
and U14299 (N_14299,N_14153,N_14159);
nand U14300 (N_14300,N_14186,N_14045);
nand U14301 (N_14301,N_14022,N_14027);
or U14302 (N_14302,N_14132,N_14119);
nand U14303 (N_14303,N_14197,N_14057);
or U14304 (N_14304,N_14038,N_14040);
or U14305 (N_14305,N_14071,N_14129);
or U14306 (N_14306,N_14018,N_14006);
and U14307 (N_14307,N_14032,N_14080);
and U14308 (N_14308,N_14042,N_14061);
or U14309 (N_14309,N_14093,N_14084);
nor U14310 (N_14310,N_14134,N_14124);
nand U14311 (N_14311,N_14063,N_14184);
nand U14312 (N_14312,N_14112,N_14074);
nor U14313 (N_14313,N_14033,N_14086);
nand U14314 (N_14314,N_14101,N_14127);
and U14315 (N_14315,N_14117,N_14142);
nand U14316 (N_14316,N_14044,N_14108);
nand U14317 (N_14317,N_14117,N_14054);
and U14318 (N_14318,N_14009,N_14160);
nor U14319 (N_14319,N_14124,N_14033);
and U14320 (N_14320,N_14041,N_14006);
and U14321 (N_14321,N_14184,N_14175);
or U14322 (N_14322,N_14175,N_14162);
or U14323 (N_14323,N_14191,N_14118);
nor U14324 (N_14324,N_14124,N_14010);
or U14325 (N_14325,N_14172,N_14058);
and U14326 (N_14326,N_14177,N_14161);
nand U14327 (N_14327,N_14106,N_14083);
or U14328 (N_14328,N_14184,N_14012);
nand U14329 (N_14329,N_14005,N_14186);
nor U14330 (N_14330,N_14198,N_14054);
xnor U14331 (N_14331,N_14083,N_14197);
or U14332 (N_14332,N_14176,N_14083);
nand U14333 (N_14333,N_14052,N_14183);
or U14334 (N_14334,N_14090,N_14133);
or U14335 (N_14335,N_14109,N_14112);
nand U14336 (N_14336,N_14127,N_14169);
nor U14337 (N_14337,N_14117,N_14065);
nand U14338 (N_14338,N_14118,N_14123);
xnor U14339 (N_14339,N_14156,N_14049);
nand U14340 (N_14340,N_14138,N_14183);
nand U14341 (N_14341,N_14065,N_14079);
and U14342 (N_14342,N_14089,N_14175);
and U14343 (N_14343,N_14082,N_14132);
and U14344 (N_14344,N_14105,N_14101);
and U14345 (N_14345,N_14051,N_14136);
and U14346 (N_14346,N_14170,N_14077);
or U14347 (N_14347,N_14006,N_14181);
nand U14348 (N_14348,N_14023,N_14077);
and U14349 (N_14349,N_14071,N_14078);
and U14350 (N_14350,N_14084,N_14190);
nor U14351 (N_14351,N_14171,N_14099);
nand U14352 (N_14352,N_14151,N_14153);
nand U14353 (N_14353,N_14060,N_14182);
and U14354 (N_14354,N_14114,N_14157);
nor U14355 (N_14355,N_14140,N_14036);
or U14356 (N_14356,N_14183,N_14168);
xor U14357 (N_14357,N_14185,N_14044);
xor U14358 (N_14358,N_14064,N_14111);
and U14359 (N_14359,N_14007,N_14173);
or U14360 (N_14360,N_14067,N_14018);
nor U14361 (N_14361,N_14180,N_14133);
and U14362 (N_14362,N_14088,N_14166);
nand U14363 (N_14363,N_14136,N_14042);
nor U14364 (N_14364,N_14168,N_14021);
and U14365 (N_14365,N_14043,N_14132);
nand U14366 (N_14366,N_14025,N_14067);
or U14367 (N_14367,N_14166,N_14156);
and U14368 (N_14368,N_14120,N_14094);
or U14369 (N_14369,N_14096,N_14034);
and U14370 (N_14370,N_14183,N_14116);
nor U14371 (N_14371,N_14185,N_14113);
or U14372 (N_14372,N_14095,N_14010);
nand U14373 (N_14373,N_14123,N_14150);
xnor U14374 (N_14374,N_14195,N_14137);
and U14375 (N_14375,N_14076,N_14139);
nor U14376 (N_14376,N_14186,N_14178);
and U14377 (N_14377,N_14082,N_14191);
nand U14378 (N_14378,N_14170,N_14193);
xnor U14379 (N_14379,N_14046,N_14108);
xnor U14380 (N_14380,N_14019,N_14152);
nand U14381 (N_14381,N_14003,N_14093);
xnor U14382 (N_14382,N_14136,N_14154);
nand U14383 (N_14383,N_14188,N_14108);
and U14384 (N_14384,N_14035,N_14049);
nand U14385 (N_14385,N_14014,N_14037);
and U14386 (N_14386,N_14092,N_14045);
or U14387 (N_14387,N_14069,N_14018);
or U14388 (N_14388,N_14187,N_14128);
xor U14389 (N_14389,N_14045,N_14138);
nand U14390 (N_14390,N_14078,N_14115);
and U14391 (N_14391,N_14077,N_14076);
nor U14392 (N_14392,N_14106,N_14053);
and U14393 (N_14393,N_14195,N_14173);
or U14394 (N_14394,N_14064,N_14128);
nand U14395 (N_14395,N_14095,N_14001);
nor U14396 (N_14396,N_14068,N_14085);
nor U14397 (N_14397,N_14096,N_14106);
nand U14398 (N_14398,N_14009,N_14069);
xor U14399 (N_14399,N_14007,N_14027);
nor U14400 (N_14400,N_14255,N_14275);
and U14401 (N_14401,N_14387,N_14323);
nand U14402 (N_14402,N_14308,N_14210);
xor U14403 (N_14403,N_14230,N_14373);
or U14404 (N_14404,N_14270,N_14268);
nand U14405 (N_14405,N_14245,N_14340);
or U14406 (N_14406,N_14292,N_14372);
nand U14407 (N_14407,N_14360,N_14249);
nand U14408 (N_14408,N_14286,N_14223);
and U14409 (N_14409,N_14229,N_14246);
nor U14410 (N_14410,N_14259,N_14336);
nor U14411 (N_14411,N_14321,N_14374);
or U14412 (N_14412,N_14218,N_14297);
and U14413 (N_14413,N_14322,N_14234);
nand U14414 (N_14414,N_14248,N_14225);
and U14415 (N_14415,N_14277,N_14231);
nand U14416 (N_14416,N_14381,N_14228);
nand U14417 (N_14417,N_14298,N_14201);
nor U14418 (N_14418,N_14314,N_14318);
nand U14419 (N_14419,N_14385,N_14200);
xnor U14420 (N_14420,N_14261,N_14222);
xnor U14421 (N_14421,N_14273,N_14398);
xnor U14422 (N_14422,N_14371,N_14219);
nor U14423 (N_14423,N_14383,N_14291);
xor U14424 (N_14424,N_14312,N_14379);
nand U14425 (N_14425,N_14376,N_14296);
and U14426 (N_14426,N_14339,N_14317);
nand U14427 (N_14427,N_14375,N_14370);
nor U14428 (N_14428,N_14206,N_14350);
nor U14429 (N_14429,N_14203,N_14325);
nor U14430 (N_14430,N_14331,N_14282);
and U14431 (N_14431,N_14319,N_14324);
and U14432 (N_14432,N_14356,N_14204);
nor U14433 (N_14433,N_14377,N_14217);
xnor U14434 (N_14434,N_14279,N_14236);
nor U14435 (N_14435,N_14252,N_14281);
nand U14436 (N_14436,N_14304,N_14239);
nor U14437 (N_14437,N_14258,N_14250);
nor U14438 (N_14438,N_14251,N_14399);
or U14439 (N_14439,N_14278,N_14263);
nor U14440 (N_14440,N_14346,N_14320);
or U14441 (N_14441,N_14396,N_14334);
and U14442 (N_14442,N_14299,N_14240);
and U14443 (N_14443,N_14216,N_14352);
or U14444 (N_14444,N_14215,N_14333);
nand U14445 (N_14445,N_14305,N_14253);
nand U14446 (N_14446,N_14208,N_14311);
nand U14447 (N_14447,N_14302,N_14232);
and U14448 (N_14448,N_14337,N_14280);
or U14449 (N_14449,N_14369,N_14345);
xnor U14450 (N_14450,N_14362,N_14256);
nor U14451 (N_14451,N_14207,N_14392);
and U14452 (N_14452,N_14205,N_14264);
xor U14453 (N_14453,N_14288,N_14202);
nand U14454 (N_14454,N_14332,N_14390);
or U14455 (N_14455,N_14303,N_14307);
and U14456 (N_14456,N_14348,N_14238);
and U14457 (N_14457,N_14294,N_14293);
nor U14458 (N_14458,N_14310,N_14326);
xor U14459 (N_14459,N_14241,N_14358);
nor U14460 (N_14460,N_14226,N_14342);
nor U14461 (N_14461,N_14368,N_14316);
or U14462 (N_14462,N_14393,N_14284);
nand U14463 (N_14463,N_14367,N_14397);
and U14464 (N_14464,N_14287,N_14295);
or U14465 (N_14465,N_14366,N_14313);
nand U14466 (N_14466,N_14355,N_14365);
nand U14467 (N_14467,N_14388,N_14354);
nand U14468 (N_14468,N_14391,N_14220);
nor U14469 (N_14469,N_14254,N_14233);
or U14470 (N_14470,N_14224,N_14260);
nand U14471 (N_14471,N_14309,N_14235);
or U14472 (N_14472,N_14244,N_14283);
and U14473 (N_14473,N_14386,N_14384);
nand U14474 (N_14474,N_14214,N_14327);
nor U14475 (N_14475,N_14243,N_14209);
nand U14476 (N_14476,N_14301,N_14394);
nand U14477 (N_14477,N_14213,N_14289);
and U14478 (N_14478,N_14227,N_14272);
or U14479 (N_14479,N_14285,N_14242);
nand U14480 (N_14480,N_14290,N_14343);
or U14481 (N_14481,N_14344,N_14364);
nor U14482 (N_14482,N_14349,N_14382);
or U14483 (N_14483,N_14257,N_14271);
or U14484 (N_14484,N_14211,N_14274);
and U14485 (N_14485,N_14265,N_14335);
or U14486 (N_14486,N_14353,N_14262);
and U14487 (N_14487,N_14276,N_14237);
or U14488 (N_14488,N_14266,N_14267);
nand U14489 (N_14489,N_14315,N_14380);
nand U14490 (N_14490,N_14330,N_14378);
or U14491 (N_14491,N_14212,N_14347);
xnor U14492 (N_14492,N_14351,N_14329);
and U14493 (N_14493,N_14357,N_14328);
and U14494 (N_14494,N_14306,N_14247);
and U14495 (N_14495,N_14389,N_14361);
nand U14496 (N_14496,N_14363,N_14395);
and U14497 (N_14497,N_14300,N_14221);
or U14498 (N_14498,N_14269,N_14341);
or U14499 (N_14499,N_14359,N_14338);
nand U14500 (N_14500,N_14361,N_14211);
and U14501 (N_14501,N_14363,N_14397);
xor U14502 (N_14502,N_14240,N_14371);
nand U14503 (N_14503,N_14367,N_14387);
nor U14504 (N_14504,N_14355,N_14207);
and U14505 (N_14505,N_14271,N_14337);
and U14506 (N_14506,N_14340,N_14218);
nor U14507 (N_14507,N_14366,N_14266);
and U14508 (N_14508,N_14237,N_14317);
xnor U14509 (N_14509,N_14329,N_14233);
or U14510 (N_14510,N_14391,N_14350);
or U14511 (N_14511,N_14370,N_14388);
nor U14512 (N_14512,N_14256,N_14323);
nor U14513 (N_14513,N_14311,N_14398);
nand U14514 (N_14514,N_14281,N_14346);
nand U14515 (N_14515,N_14236,N_14241);
or U14516 (N_14516,N_14294,N_14324);
nand U14517 (N_14517,N_14384,N_14292);
nand U14518 (N_14518,N_14276,N_14351);
and U14519 (N_14519,N_14234,N_14265);
nor U14520 (N_14520,N_14221,N_14362);
and U14521 (N_14521,N_14330,N_14281);
and U14522 (N_14522,N_14312,N_14310);
and U14523 (N_14523,N_14310,N_14305);
nand U14524 (N_14524,N_14309,N_14234);
and U14525 (N_14525,N_14341,N_14346);
and U14526 (N_14526,N_14215,N_14341);
nor U14527 (N_14527,N_14223,N_14361);
xnor U14528 (N_14528,N_14291,N_14315);
or U14529 (N_14529,N_14323,N_14203);
nor U14530 (N_14530,N_14349,N_14296);
nor U14531 (N_14531,N_14356,N_14371);
nand U14532 (N_14532,N_14395,N_14228);
or U14533 (N_14533,N_14306,N_14214);
and U14534 (N_14534,N_14372,N_14248);
and U14535 (N_14535,N_14379,N_14253);
or U14536 (N_14536,N_14399,N_14250);
xor U14537 (N_14537,N_14282,N_14229);
and U14538 (N_14538,N_14319,N_14333);
or U14539 (N_14539,N_14236,N_14262);
and U14540 (N_14540,N_14303,N_14395);
nand U14541 (N_14541,N_14296,N_14289);
nand U14542 (N_14542,N_14306,N_14381);
nor U14543 (N_14543,N_14208,N_14369);
and U14544 (N_14544,N_14319,N_14228);
and U14545 (N_14545,N_14336,N_14385);
nand U14546 (N_14546,N_14320,N_14235);
or U14547 (N_14547,N_14283,N_14205);
or U14548 (N_14548,N_14235,N_14391);
nor U14549 (N_14549,N_14329,N_14222);
xor U14550 (N_14550,N_14224,N_14201);
and U14551 (N_14551,N_14200,N_14284);
and U14552 (N_14552,N_14319,N_14387);
and U14553 (N_14553,N_14233,N_14321);
nor U14554 (N_14554,N_14344,N_14274);
nor U14555 (N_14555,N_14370,N_14221);
nor U14556 (N_14556,N_14316,N_14367);
nand U14557 (N_14557,N_14364,N_14373);
or U14558 (N_14558,N_14350,N_14274);
or U14559 (N_14559,N_14213,N_14292);
or U14560 (N_14560,N_14227,N_14393);
and U14561 (N_14561,N_14203,N_14339);
or U14562 (N_14562,N_14367,N_14285);
nor U14563 (N_14563,N_14309,N_14239);
nand U14564 (N_14564,N_14266,N_14385);
and U14565 (N_14565,N_14212,N_14281);
nor U14566 (N_14566,N_14276,N_14291);
xnor U14567 (N_14567,N_14209,N_14394);
or U14568 (N_14568,N_14341,N_14360);
or U14569 (N_14569,N_14202,N_14348);
nor U14570 (N_14570,N_14257,N_14397);
and U14571 (N_14571,N_14380,N_14349);
or U14572 (N_14572,N_14322,N_14366);
nor U14573 (N_14573,N_14333,N_14236);
nand U14574 (N_14574,N_14355,N_14270);
and U14575 (N_14575,N_14238,N_14322);
or U14576 (N_14576,N_14370,N_14365);
nand U14577 (N_14577,N_14342,N_14228);
or U14578 (N_14578,N_14372,N_14223);
and U14579 (N_14579,N_14309,N_14253);
nand U14580 (N_14580,N_14306,N_14391);
and U14581 (N_14581,N_14230,N_14201);
nor U14582 (N_14582,N_14332,N_14377);
nand U14583 (N_14583,N_14327,N_14330);
nor U14584 (N_14584,N_14329,N_14334);
xnor U14585 (N_14585,N_14322,N_14203);
and U14586 (N_14586,N_14310,N_14295);
nor U14587 (N_14587,N_14311,N_14245);
and U14588 (N_14588,N_14238,N_14291);
nand U14589 (N_14589,N_14284,N_14341);
and U14590 (N_14590,N_14289,N_14227);
nand U14591 (N_14591,N_14203,N_14359);
nand U14592 (N_14592,N_14355,N_14376);
xnor U14593 (N_14593,N_14254,N_14307);
or U14594 (N_14594,N_14213,N_14322);
xnor U14595 (N_14595,N_14284,N_14343);
nand U14596 (N_14596,N_14263,N_14355);
xnor U14597 (N_14597,N_14323,N_14347);
nor U14598 (N_14598,N_14209,N_14356);
nor U14599 (N_14599,N_14201,N_14294);
xor U14600 (N_14600,N_14573,N_14494);
or U14601 (N_14601,N_14425,N_14515);
or U14602 (N_14602,N_14520,N_14480);
or U14603 (N_14603,N_14489,N_14579);
nor U14604 (N_14604,N_14427,N_14432);
or U14605 (N_14605,N_14424,N_14485);
and U14606 (N_14606,N_14500,N_14445);
or U14607 (N_14607,N_14576,N_14598);
nand U14608 (N_14608,N_14479,N_14434);
or U14609 (N_14609,N_14521,N_14501);
nor U14610 (N_14610,N_14530,N_14556);
xnor U14611 (N_14611,N_14478,N_14514);
nand U14612 (N_14612,N_14509,N_14451);
nand U14613 (N_14613,N_14578,N_14420);
nand U14614 (N_14614,N_14512,N_14558);
nand U14615 (N_14615,N_14452,N_14547);
nand U14616 (N_14616,N_14462,N_14562);
nor U14617 (N_14617,N_14542,N_14511);
or U14618 (N_14618,N_14444,N_14519);
nor U14619 (N_14619,N_14475,N_14402);
nand U14620 (N_14620,N_14412,N_14477);
nand U14621 (N_14621,N_14551,N_14554);
and U14622 (N_14622,N_14414,N_14454);
and U14623 (N_14623,N_14580,N_14570);
and U14624 (N_14624,N_14428,N_14599);
nand U14625 (N_14625,N_14552,N_14563);
nand U14626 (N_14626,N_14539,N_14585);
nand U14627 (N_14627,N_14429,N_14410);
nand U14628 (N_14628,N_14442,N_14491);
nand U14629 (N_14629,N_14474,N_14409);
nor U14630 (N_14630,N_14415,N_14437);
or U14631 (N_14631,N_14400,N_14565);
nor U14632 (N_14632,N_14470,N_14411);
nor U14633 (N_14633,N_14418,N_14543);
nor U14634 (N_14634,N_14495,N_14527);
nor U14635 (N_14635,N_14533,N_14589);
nor U14636 (N_14636,N_14540,N_14545);
nand U14637 (N_14637,N_14564,N_14404);
nor U14638 (N_14638,N_14522,N_14526);
or U14639 (N_14639,N_14513,N_14464);
xor U14640 (N_14640,N_14468,N_14488);
nor U14641 (N_14641,N_14476,N_14504);
nor U14642 (N_14642,N_14557,N_14426);
and U14643 (N_14643,N_14571,N_14456);
or U14644 (N_14644,N_14498,N_14487);
nor U14645 (N_14645,N_14593,N_14532);
xor U14646 (N_14646,N_14518,N_14484);
or U14647 (N_14647,N_14544,N_14506);
xor U14648 (N_14648,N_14496,N_14531);
and U14649 (N_14649,N_14457,N_14465);
and U14650 (N_14650,N_14566,N_14471);
or U14651 (N_14651,N_14463,N_14422);
nand U14652 (N_14652,N_14455,N_14523);
or U14653 (N_14653,N_14441,N_14555);
nand U14654 (N_14654,N_14583,N_14569);
nand U14655 (N_14655,N_14560,N_14449);
and U14656 (N_14656,N_14586,N_14472);
nand U14657 (N_14657,N_14417,N_14597);
and U14658 (N_14658,N_14440,N_14546);
or U14659 (N_14659,N_14497,N_14436);
or U14660 (N_14660,N_14469,N_14447);
nor U14661 (N_14661,N_14406,N_14507);
or U14662 (N_14662,N_14482,N_14505);
nand U14663 (N_14663,N_14458,N_14433);
nand U14664 (N_14664,N_14517,N_14516);
nand U14665 (N_14665,N_14446,N_14588);
nor U14666 (N_14666,N_14439,N_14508);
nor U14667 (N_14667,N_14535,N_14407);
nor U14668 (N_14668,N_14419,N_14460);
nand U14669 (N_14669,N_14575,N_14524);
xor U14670 (N_14670,N_14423,N_14537);
nor U14671 (N_14671,N_14525,N_14592);
nor U14672 (N_14672,N_14541,N_14403);
xnor U14673 (N_14673,N_14408,N_14550);
xnor U14674 (N_14674,N_14450,N_14572);
or U14675 (N_14675,N_14529,N_14559);
nor U14676 (N_14676,N_14453,N_14549);
nor U14677 (N_14677,N_14461,N_14581);
or U14678 (N_14678,N_14584,N_14413);
or U14679 (N_14679,N_14536,N_14421);
or U14680 (N_14680,N_14538,N_14405);
or U14681 (N_14681,N_14561,N_14448);
or U14682 (N_14682,N_14568,N_14567);
nor U14683 (N_14683,N_14577,N_14459);
or U14684 (N_14684,N_14574,N_14486);
nand U14685 (N_14685,N_14467,N_14595);
or U14686 (N_14686,N_14499,N_14466);
or U14687 (N_14687,N_14431,N_14591);
nor U14688 (N_14688,N_14490,N_14582);
or U14689 (N_14689,N_14435,N_14553);
nand U14690 (N_14690,N_14587,N_14493);
nand U14691 (N_14691,N_14594,N_14590);
nand U14692 (N_14692,N_14481,N_14502);
nand U14693 (N_14693,N_14438,N_14528);
nor U14694 (N_14694,N_14416,N_14596);
or U14695 (N_14695,N_14548,N_14534);
nand U14696 (N_14696,N_14492,N_14510);
nand U14697 (N_14697,N_14503,N_14473);
or U14698 (N_14698,N_14443,N_14483);
nand U14699 (N_14699,N_14401,N_14430);
and U14700 (N_14700,N_14462,N_14490);
or U14701 (N_14701,N_14402,N_14526);
nand U14702 (N_14702,N_14592,N_14561);
nand U14703 (N_14703,N_14402,N_14581);
and U14704 (N_14704,N_14495,N_14509);
and U14705 (N_14705,N_14501,N_14434);
nor U14706 (N_14706,N_14511,N_14429);
and U14707 (N_14707,N_14514,N_14508);
xnor U14708 (N_14708,N_14514,N_14579);
nor U14709 (N_14709,N_14536,N_14496);
nand U14710 (N_14710,N_14500,N_14546);
nand U14711 (N_14711,N_14450,N_14411);
nor U14712 (N_14712,N_14446,N_14436);
nand U14713 (N_14713,N_14513,N_14565);
nand U14714 (N_14714,N_14481,N_14548);
nor U14715 (N_14715,N_14417,N_14411);
and U14716 (N_14716,N_14462,N_14426);
or U14717 (N_14717,N_14523,N_14457);
or U14718 (N_14718,N_14414,N_14402);
nand U14719 (N_14719,N_14459,N_14401);
nor U14720 (N_14720,N_14432,N_14436);
nand U14721 (N_14721,N_14471,N_14473);
nor U14722 (N_14722,N_14508,N_14577);
nor U14723 (N_14723,N_14474,N_14540);
nand U14724 (N_14724,N_14508,N_14418);
nand U14725 (N_14725,N_14495,N_14414);
xor U14726 (N_14726,N_14449,N_14531);
or U14727 (N_14727,N_14528,N_14580);
nor U14728 (N_14728,N_14589,N_14448);
xor U14729 (N_14729,N_14471,N_14588);
xor U14730 (N_14730,N_14584,N_14536);
nand U14731 (N_14731,N_14533,N_14529);
and U14732 (N_14732,N_14459,N_14599);
nor U14733 (N_14733,N_14421,N_14407);
nor U14734 (N_14734,N_14495,N_14413);
and U14735 (N_14735,N_14573,N_14489);
or U14736 (N_14736,N_14596,N_14514);
nand U14737 (N_14737,N_14467,N_14576);
nor U14738 (N_14738,N_14510,N_14572);
nand U14739 (N_14739,N_14547,N_14403);
nand U14740 (N_14740,N_14598,N_14539);
or U14741 (N_14741,N_14515,N_14421);
xnor U14742 (N_14742,N_14510,N_14429);
nand U14743 (N_14743,N_14446,N_14491);
nor U14744 (N_14744,N_14464,N_14434);
or U14745 (N_14745,N_14495,N_14580);
nand U14746 (N_14746,N_14529,N_14413);
nand U14747 (N_14747,N_14562,N_14420);
nand U14748 (N_14748,N_14475,N_14534);
or U14749 (N_14749,N_14577,N_14551);
nand U14750 (N_14750,N_14442,N_14404);
or U14751 (N_14751,N_14527,N_14557);
nand U14752 (N_14752,N_14532,N_14468);
xnor U14753 (N_14753,N_14440,N_14536);
and U14754 (N_14754,N_14406,N_14464);
and U14755 (N_14755,N_14405,N_14511);
xor U14756 (N_14756,N_14547,N_14537);
xnor U14757 (N_14757,N_14551,N_14449);
or U14758 (N_14758,N_14580,N_14571);
nand U14759 (N_14759,N_14530,N_14422);
or U14760 (N_14760,N_14552,N_14426);
nand U14761 (N_14761,N_14489,N_14436);
nand U14762 (N_14762,N_14429,N_14599);
nor U14763 (N_14763,N_14561,N_14590);
or U14764 (N_14764,N_14407,N_14548);
nand U14765 (N_14765,N_14462,N_14459);
nor U14766 (N_14766,N_14449,N_14514);
and U14767 (N_14767,N_14563,N_14406);
nand U14768 (N_14768,N_14546,N_14594);
nand U14769 (N_14769,N_14542,N_14497);
nor U14770 (N_14770,N_14504,N_14487);
nand U14771 (N_14771,N_14591,N_14486);
nor U14772 (N_14772,N_14558,N_14525);
xor U14773 (N_14773,N_14582,N_14495);
nor U14774 (N_14774,N_14566,N_14413);
nor U14775 (N_14775,N_14456,N_14436);
or U14776 (N_14776,N_14531,N_14497);
nor U14777 (N_14777,N_14493,N_14590);
and U14778 (N_14778,N_14436,N_14400);
or U14779 (N_14779,N_14590,N_14579);
or U14780 (N_14780,N_14564,N_14451);
nand U14781 (N_14781,N_14573,N_14515);
xnor U14782 (N_14782,N_14552,N_14572);
and U14783 (N_14783,N_14513,N_14500);
nor U14784 (N_14784,N_14530,N_14453);
nor U14785 (N_14785,N_14433,N_14533);
or U14786 (N_14786,N_14536,N_14476);
xor U14787 (N_14787,N_14411,N_14439);
or U14788 (N_14788,N_14429,N_14497);
and U14789 (N_14789,N_14424,N_14561);
nand U14790 (N_14790,N_14401,N_14417);
nand U14791 (N_14791,N_14404,N_14518);
or U14792 (N_14792,N_14431,N_14559);
nor U14793 (N_14793,N_14593,N_14427);
and U14794 (N_14794,N_14557,N_14523);
nand U14795 (N_14795,N_14475,N_14487);
or U14796 (N_14796,N_14424,N_14448);
nand U14797 (N_14797,N_14449,N_14414);
nor U14798 (N_14798,N_14522,N_14513);
nand U14799 (N_14799,N_14595,N_14517);
nand U14800 (N_14800,N_14729,N_14610);
nor U14801 (N_14801,N_14749,N_14792);
and U14802 (N_14802,N_14731,N_14691);
and U14803 (N_14803,N_14611,N_14743);
xnor U14804 (N_14804,N_14655,N_14783);
xnor U14805 (N_14805,N_14780,N_14794);
and U14806 (N_14806,N_14720,N_14609);
and U14807 (N_14807,N_14651,N_14796);
nor U14808 (N_14808,N_14613,N_14640);
nor U14809 (N_14809,N_14678,N_14671);
and U14810 (N_14810,N_14774,N_14701);
and U14811 (N_14811,N_14681,N_14776);
nand U14812 (N_14812,N_14733,N_14706);
nand U14813 (N_14813,N_14646,N_14614);
nand U14814 (N_14814,N_14675,N_14739);
nor U14815 (N_14815,N_14652,N_14732);
nor U14816 (N_14816,N_14659,N_14735);
or U14817 (N_14817,N_14782,N_14606);
and U14818 (N_14818,N_14661,N_14742);
and U14819 (N_14819,N_14694,N_14789);
and U14820 (N_14820,N_14638,N_14639);
and U14821 (N_14821,N_14654,N_14762);
nand U14822 (N_14822,N_14622,N_14664);
or U14823 (N_14823,N_14764,N_14605);
nand U14824 (N_14824,N_14628,N_14790);
and U14825 (N_14825,N_14663,N_14788);
nor U14826 (N_14826,N_14620,N_14756);
xnor U14827 (N_14827,N_14647,N_14696);
and U14828 (N_14828,N_14786,N_14630);
xnor U14829 (N_14829,N_14777,N_14693);
nand U14830 (N_14830,N_14744,N_14722);
nand U14831 (N_14831,N_14616,N_14716);
nand U14832 (N_14832,N_14715,N_14726);
nand U14833 (N_14833,N_14632,N_14684);
nand U14834 (N_14834,N_14736,N_14757);
and U14835 (N_14835,N_14626,N_14673);
xnor U14836 (N_14836,N_14703,N_14644);
nor U14837 (N_14837,N_14688,N_14772);
or U14838 (N_14838,N_14636,N_14650);
or U14839 (N_14839,N_14666,N_14773);
nor U14840 (N_14840,N_14665,N_14676);
or U14841 (N_14841,N_14752,N_14761);
nor U14842 (N_14842,N_14692,N_14689);
nor U14843 (N_14843,N_14766,N_14769);
nand U14844 (N_14844,N_14759,N_14635);
xnor U14845 (N_14845,N_14658,N_14799);
or U14846 (N_14846,N_14771,N_14698);
nand U14847 (N_14847,N_14791,N_14699);
nand U14848 (N_14848,N_14704,N_14784);
and U14849 (N_14849,N_14719,N_14708);
or U14850 (N_14850,N_14672,N_14755);
or U14851 (N_14851,N_14770,N_14741);
or U14852 (N_14852,N_14656,N_14730);
nand U14853 (N_14853,N_14685,N_14760);
or U14854 (N_14854,N_14767,N_14662);
nand U14855 (N_14855,N_14738,N_14718);
nand U14856 (N_14856,N_14723,N_14748);
nor U14857 (N_14857,N_14642,N_14618);
nand U14858 (N_14858,N_14612,N_14680);
and U14859 (N_14859,N_14674,N_14600);
nor U14860 (N_14860,N_14607,N_14763);
and U14861 (N_14861,N_14781,N_14751);
or U14862 (N_14862,N_14617,N_14737);
nand U14863 (N_14863,N_14787,N_14670);
nor U14864 (N_14864,N_14793,N_14734);
or U14865 (N_14865,N_14775,N_14746);
xnor U14866 (N_14866,N_14725,N_14697);
xor U14867 (N_14867,N_14623,N_14687);
nand U14868 (N_14868,N_14619,N_14669);
nand U14869 (N_14869,N_14603,N_14634);
nand U14870 (N_14870,N_14690,N_14702);
nor U14871 (N_14871,N_14682,N_14768);
nand U14872 (N_14872,N_14785,N_14795);
or U14873 (N_14873,N_14683,N_14625);
xnor U14874 (N_14874,N_14710,N_14627);
nand U14875 (N_14875,N_14645,N_14717);
nand U14876 (N_14876,N_14705,N_14667);
nand U14877 (N_14877,N_14754,N_14637);
and U14878 (N_14878,N_14633,N_14712);
or U14879 (N_14879,N_14601,N_14753);
nand U14880 (N_14880,N_14657,N_14714);
and U14881 (N_14881,N_14747,N_14649);
nand U14882 (N_14882,N_14629,N_14713);
nor U14883 (N_14883,N_14624,N_14631);
nand U14884 (N_14884,N_14608,N_14679);
nand U14885 (N_14885,N_14695,N_14653);
nand U14886 (N_14886,N_14707,N_14648);
and U14887 (N_14887,N_14711,N_14643);
and U14888 (N_14888,N_14778,N_14745);
nand U14889 (N_14889,N_14615,N_14709);
or U14890 (N_14890,N_14797,N_14700);
nand U14891 (N_14891,N_14765,N_14798);
and U14892 (N_14892,N_14740,N_14641);
and U14893 (N_14893,N_14660,N_14758);
nand U14894 (N_14894,N_14728,N_14779);
or U14895 (N_14895,N_14621,N_14750);
nor U14896 (N_14896,N_14668,N_14604);
or U14897 (N_14897,N_14721,N_14727);
and U14898 (N_14898,N_14724,N_14686);
nor U14899 (N_14899,N_14677,N_14602);
nand U14900 (N_14900,N_14732,N_14717);
nand U14901 (N_14901,N_14739,N_14730);
nor U14902 (N_14902,N_14705,N_14620);
and U14903 (N_14903,N_14736,N_14688);
xnor U14904 (N_14904,N_14627,N_14770);
nor U14905 (N_14905,N_14783,N_14624);
or U14906 (N_14906,N_14771,N_14606);
nor U14907 (N_14907,N_14717,N_14706);
nor U14908 (N_14908,N_14689,N_14705);
or U14909 (N_14909,N_14665,N_14700);
nand U14910 (N_14910,N_14785,N_14648);
nand U14911 (N_14911,N_14651,N_14783);
and U14912 (N_14912,N_14712,N_14683);
or U14913 (N_14913,N_14779,N_14783);
nand U14914 (N_14914,N_14632,N_14763);
nand U14915 (N_14915,N_14677,N_14692);
or U14916 (N_14916,N_14676,N_14682);
nor U14917 (N_14917,N_14678,N_14730);
nand U14918 (N_14918,N_14764,N_14709);
and U14919 (N_14919,N_14631,N_14740);
nand U14920 (N_14920,N_14766,N_14763);
nand U14921 (N_14921,N_14711,N_14772);
nor U14922 (N_14922,N_14682,N_14754);
and U14923 (N_14923,N_14629,N_14720);
and U14924 (N_14924,N_14743,N_14624);
xor U14925 (N_14925,N_14650,N_14673);
nand U14926 (N_14926,N_14679,N_14699);
xor U14927 (N_14927,N_14648,N_14615);
xor U14928 (N_14928,N_14789,N_14615);
nand U14929 (N_14929,N_14691,N_14654);
or U14930 (N_14930,N_14663,N_14799);
nand U14931 (N_14931,N_14683,N_14662);
and U14932 (N_14932,N_14613,N_14614);
nor U14933 (N_14933,N_14682,N_14660);
xnor U14934 (N_14934,N_14736,N_14658);
nor U14935 (N_14935,N_14691,N_14606);
nor U14936 (N_14936,N_14788,N_14618);
nand U14937 (N_14937,N_14734,N_14718);
nand U14938 (N_14938,N_14621,N_14763);
nor U14939 (N_14939,N_14629,N_14777);
nand U14940 (N_14940,N_14749,N_14710);
nand U14941 (N_14941,N_14604,N_14669);
or U14942 (N_14942,N_14623,N_14678);
nand U14943 (N_14943,N_14782,N_14684);
and U14944 (N_14944,N_14730,N_14702);
nor U14945 (N_14945,N_14602,N_14603);
nor U14946 (N_14946,N_14721,N_14657);
nand U14947 (N_14947,N_14636,N_14706);
nor U14948 (N_14948,N_14739,N_14757);
nand U14949 (N_14949,N_14702,N_14695);
nor U14950 (N_14950,N_14790,N_14648);
and U14951 (N_14951,N_14796,N_14775);
and U14952 (N_14952,N_14710,N_14648);
xnor U14953 (N_14953,N_14654,N_14666);
nand U14954 (N_14954,N_14759,N_14697);
nor U14955 (N_14955,N_14731,N_14793);
or U14956 (N_14956,N_14767,N_14669);
nand U14957 (N_14957,N_14735,N_14618);
nor U14958 (N_14958,N_14663,N_14652);
and U14959 (N_14959,N_14753,N_14757);
and U14960 (N_14960,N_14799,N_14749);
nand U14961 (N_14961,N_14620,N_14684);
nor U14962 (N_14962,N_14748,N_14730);
and U14963 (N_14963,N_14616,N_14636);
or U14964 (N_14964,N_14652,N_14771);
or U14965 (N_14965,N_14774,N_14772);
and U14966 (N_14966,N_14733,N_14643);
nand U14967 (N_14967,N_14718,N_14794);
or U14968 (N_14968,N_14676,N_14679);
nor U14969 (N_14969,N_14745,N_14743);
nor U14970 (N_14970,N_14625,N_14759);
or U14971 (N_14971,N_14662,N_14724);
xor U14972 (N_14972,N_14689,N_14750);
nor U14973 (N_14973,N_14731,N_14628);
and U14974 (N_14974,N_14625,N_14774);
and U14975 (N_14975,N_14668,N_14770);
and U14976 (N_14976,N_14770,N_14631);
and U14977 (N_14977,N_14799,N_14677);
and U14978 (N_14978,N_14685,N_14627);
and U14979 (N_14979,N_14661,N_14721);
nand U14980 (N_14980,N_14766,N_14606);
nand U14981 (N_14981,N_14616,N_14722);
nand U14982 (N_14982,N_14643,N_14650);
nand U14983 (N_14983,N_14761,N_14626);
nor U14984 (N_14984,N_14693,N_14763);
or U14985 (N_14985,N_14762,N_14733);
nor U14986 (N_14986,N_14614,N_14619);
nand U14987 (N_14987,N_14713,N_14770);
xnor U14988 (N_14988,N_14623,N_14610);
nor U14989 (N_14989,N_14789,N_14798);
and U14990 (N_14990,N_14742,N_14669);
xor U14991 (N_14991,N_14715,N_14686);
xor U14992 (N_14992,N_14600,N_14639);
xor U14993 (N_14993,N_14606,N_14628);
nor U14994 (N_14994,N_14647,N_14658);
or U14995 (N_14995,N_14766,N_14693);
and U14996 (N_14996,N_14607,N_14612);
nor U14997 (N_14997,N_14623,N_14637);
nor U14998 (N_14998,N_14674,N_14762);
nand U14999 (N_14999,N_14777,N_14753);
and UO_0 (O_0,N_14899,N_14851);
nor UO_1 (O_1,N_14809,N_14859);
and UO_2 (O_2,N_14912,N_14925);
or UO_3 (O_3,N_14961,N_14864);
nor UO_4 (O_4,N_14897,N_14824);
xor UO_5 (O_5,N_14835,N_14936);
nand UO_6 (O_6,N_14834,N_14847);
or UO_7 (O_7,N_14874,N_14911);
and UO_8 (O_8,N_14916,N_14901);
xor UO_9 (O_9,N_14976,N_14883);
xor UO_10 (O_10,N_14826,N_14960);
nor UO_11 (O_11,N_14998,N_14831);
nand UO_12 (O_12,N_14969,N_14999);
and UO_13 (O_13,N_14931,N_14879);
nand UO_14 (O_14,N_14853,N_14904);
and UO_15 (O_15,N_14873,N_14946);
nand UO_16 (O_16,N_14935,N_14881);
nor UO_17 (O_17,N_14804,N_14808);
or UO_18 (O_18,N_14948,N_14829);
nor UO_19 (O_19,N_14842,N_14887);
or UO_20 (O_20,N_14856,N_14855);
and UO_21 (O_21,N_14869,N_14983);
nand UO_22 (O_22,N_14813,N_14937);
nor UO_23 (O_23,N_14920,N_14955);
and UO_24 (O_24,N_14979,N_14862);
xnor UO_25 (O_25,N_14845,N_14885);
and UO_26 (O_26,N_14801,N_14872);
or UO_27 (O_27,N_14972,N_14819);
or UO_28 (O_28,N_14910,N_14923);
nand UO_29 (O_29,N_14918,N_14876);
xnor UO_30 (O_30,N_14858,N_14861);
or UO_31 (O_31,N_14933,N_14956);
nor UO_32 (O_32,N_14970,N_14803);
nand UO_33 (O_33,N_14909,N_14841);
nand UO_34 (O_34,N_14940,N_14894);
or UO_35 (O_35,N_14973,N_14882);
and UO_36 (O_36,N_14898,N_14815);
nand UO_37 (O_37,N_14832,N_14914);
nor UO_38 (O_38,N_14891,N_14958);
nand UO_39 (O_39,N_14828,N_14896);
or UO_40 (O_40,N_14850,N_14836);
nor UO_41 (O_41,N_14848,N_14963);
nor UO_42 (O_42,N_14895,N_14844);
or UO_43 (O_43,N_14886,N_14945);
nand UO_44 (O_44,N_14964,N_14857);
and UO_45 (O_45,N_14852,N_14839);
nor UO_46 (O_46,N_14990,N_14843);
and UO_47 (O_47,N_14978,N_14965);
and UO_48 (O_48,N_14866,N_14989);
xnor UO_49 (O_49,N_14902,N_14967);
nand UO_50 (O_50,N_14928,N_14878);
xor UO_51 (O_51,N_14868,N_14849);
nand UO_52 (O_52,N_14917,N_14877);
nand UO_53 (O_53,N_14957,N_14988);
or UO_54 (O_54,N_14870,N_14997);
nor UO_55 (O_55,N_14949,N_14837);
xor UO_56 (O_56,N_14977,N_14943);
xnor UO_57 (O_57,N_14986,N_14906);
or UO_58 (O_58,N_14980,N_14867);
and UO_59 (O_59,N_14814,N_14954);
nor UO_60 (O_60,N_14995,N_14982);
nor UO_61 (O_61,N_14822,N_14825);
or UO_62 (O_62,N_14875,N_14929);
nand UO_63 (O_63,N_14806,N_14975);
or UO_64 (O_64,N_14865,N_14846);
and UO_65 (O_65,N_14830,N_14924);
or UO_66 (O_66,N_14854,N_14952);
or UO_67 (O_67,N_14922,N_14971);
xnor UO_68 (O_68,N_14932,N_14903);
and UO_69 (O_69,N_14817,N_14941);
or UO_70 (O_70,N_14900,N_14816);
nand UO_71 (O_71,N_14863,N_14993);
xnor UO_72 (O_72,N_14893,N_14939);
and UO_73 (O_73,N_14892,N_14915);
or UO_74 (O_74,N_14938,N_14944);
xor UO_75 (O_75,N_14913,N_14820);
nor UO_76 (O_76,N_14919,N_14947);
and UO_77 (O_77,N_14818,N_14884);
nor UO_78 (O_78,N_14927,N_14802);
or UO_79 (O_79,N_14908,N_14921);
or UO_80 (O_80,N_14833,N_14805);
and UO_81 (O_81,N_14984,N_14907);
nand UO_82 (O_82,N_14926,N_14840);
xnor UO_83 (O_83,N_14959,N_14966);
or UO_84 (O_84,N_14953,N_14985);
and UO_85 (O_85,N_14994,N_14974);
and UO_86 (O_86,N_14827,N_14890);
nand UO_87 (O_87,N_14821,N_14871);
xnor UO_88 (O_88,N_14951,N_14962);
and UO_89 (O_89,N_14934,N_14968);
or UO_90 (O_90,N_14991,N_14860);
and UO_91 (O_91,N_14889,N_14810);
nand UO_92 (O_92,N_14992,N_14823);
and UO_93 (O_93,N_14942,N_14987);
nand UO_94 (O_94,N_14930,N_14838);
nor UO_95 (O_95,N_14888,N_14981);
nand UO_96 (O_96,N_14811,N_14800);
nand UO_97 (O_97,N_14996,N_14905);
or UO_98 (O_98,N_14950,N_14807);
nand UO_99 (O_99,N_14812,N_14880);
and UO_100 (O_100,N_14823,N_14834);
nor UO_101 (O_101,N_14914,N_14909);
and UO_102 (O_102,N_14889,N_14803);
or UO_103 (O_103,N_14953,N_14867);
nor UO_104 (O_104,N_14831,N_14976);
nor UO_105 (O_105,N_14897,N_14875);
nor UO_106 (O_106,N_14882,N_14939);
and UO_107 (O_107,N_14936,N_14892);
xor UO_108 (O_108,N_14964,N_14924);
and UO_109 (O_109,N_14992,N_14951);
xor UO_110 (O_110,N_14826,N_14959);
nand UO_111 (O_111,N_14947,N_14810);
nor UO_112 (O_112,N_14982,N_14993);
nor UO_113 (O_113,N_14895,N_14887);
or UO_114 (O_114,N_14859,N_14973);
xor UO_115 (O_115,N_14901,N_14962);
nor UO_116 (O_116,N_14866,N_14833);
and UO_117 (O_117,N_14816,N_14950);
or UO_118 (O_118,N_14837,N_14858);
nand UO_119 (O_119,N_14944,N_14891);
and UO_120 (O_120,N_14913,N_14862);
nand UO_121 (O_121,N_14936,N_14935);
and UO_122 (O_122,N_14898,N_14910);
nand UO_123 (O_123,N_14896,N_14920);
and UO_124 (O_124,N_14820,N_14814);
xnor UO_125 (O_125,N_14997,N_14864);
and UO_126 (O_126,N_14865,N_14864);
or UO_127 (O_127,N_14997,N_14915);
nor UO_128 (O_128,N_14810,N_14854);
xnor UO_129 (O_129,N_14970,N_14932);
nor UO_130 (O_130,N_14918,N_14899);
nand UO_131 (O_131,N_14918,N_14916);
and UO_132 (O_132,N_14879,N_14989);
nand UO_133 (O_133,N_14819,N_14929);
nand UO_134 (O_134,N_14827,N_14852);
and UO_135 (O_135,N_14937,N_14931);
nor UO_136 (O_136,N_14964,N_14830);
nor UO_137 (O_137,N_14881,N_14895);
nand UO_138 (O_138,N_14966,N_14943);
and UO_139 (O_139,N_14917,N_14813);
nor UO_140 (O_140,N_14923,N_14823);
or UO_141 (O_141,N_14859,N_14857);
or UO_142 (O_142,N_14986,N_14953);
nor UO_143 (O_143,N_14966,N_14909);
nand UO_144 (O_144,N_14853,N_14980);
and UO_145 (O_145,N_14918,N_14982);
nand UO_146 (O_146,N_14852,N_14923);
nor UO_147 (O_147,N_14826,N_14970);
and UO_148 (O_148,N_14907,N_14873);
or UO_149 (O_149,N_14802,N_14948);
nand UO_150 (O_150,N_14880,N_14894);
nor UO_151 (O_151,N_14973,N_14910);
or UO_152 (O_152,N_14920,N_14979);
or UO_153 (O_153,N_14813,N_14966);
or UO_154 (O_154,N_14813,N_14913);
nand UO_155 (O_155,N_14939,N_14934);
nor UO_156 (O_156,N_14857,N_14903);
xnor UO_157 (O_157,N_14864,N_14807);
nand UO_158 (O_158,N_14883,N_14916);
nor UO_159 (O_159,N_14839,N_14854);
or UO_160 (O_160,N_14839,N_14848);
or UO_161 (O_161,N_14989,N_14833);
or UO_162 (O_162,N_14831,N_14810);
nor UO_163 (O_163,N_14850,N_14982);
nand UO_164 (O_164,N_14810,N_14897);
xnor UO_165 (O_165,N_14887,N_14902);
nand UO_166 (O_166,N_14933,N_14919);
nand UO_167 (O_167,N_14870,N_14822);
or UO_168 (O_168,N_14952,N_14887);
or UO_169 (O_169,N_14844,N_14925);
and UO_170 (O_170,N_14935,N_14865);
nand UO_171 (O_171,N_14949,N_14963);
or UO_172 (O_172,N_14970,N_14819);
nand UO_173 (O_173,N_14951,N_14944);
xnor UO_174 (O_174,N_14982,N_14805);
and UO_175 (O_175,N_14886,N_14879);
xor UO_176 (O_176,N_14856,N_14881);
nand UO_177 (O_177,N_14876,N_14864);
and UO_178 (O_178,N_14981,N_14849);
nand UO_179 (O_179,N_14827,N_14837);
and UO_180 (O_180,N_14910,N_14860);
or UO_181 (O_181,N_14971,N_14921);
nand UO_182 (O_182,N_14853,N_14993);
nand UO_183 (O_183,N_14924,N_14900);
xnor UO_184 (O_184,N_14987,N_14968);
and UO_185 (O_185,N_14961,N_14970);
xnor UO_186 (O_186,N_14957,N_14862);
or UO_187 (O_187,N_14932,N_14893);
and UO_188 (O_188,N_14869,N_14850);
or UO_189 (O_189,N_14986,N_14811);
nand UO_190 (O_190,N_14897,N_14988);
nand UO_191 (O_191,N_14995,N_14988);
nor UO_192 (O_192,N_14840,N_14935);
or UO_193 (O_193,N_14873,N_14878);
nand UO_194 (O_194,N_14994,N_14939);
nand UO_195 (O_195,N_14953,N_14875);
or UO_196 (O_196,N_14845,N_14893);
nor UO_197 (O_197,N_14889,N_14858);
nand UO_198 (O_198,N_14946,N_14856);
and UO_199 (O_199,N_14834,N_14917);
xnor UO_200 (O_200,N_14995,N_14944);
nand UO_201 (O_201,N_14956,N_14994);
or UO_202 (O_202,N_14959,N_14875);
nor UO_203 (O_203,N_14891,N_14976);
and UO_204 (O_204,N_14905,N_14849);
nand UO_205 (O_205,N_14879,N_14836);
nor UO_206 (O_206,N_14978,N_14875);
xnor UO_207 (O_207,N_14917,N_14903);
nor UO_208 (O_208,N_14989,N_14995);
nor UO_209 (O_209,N_14890,N_14918);
and UO_210 (O_210,N_14864,N_14996);
xor UO_211 (O_211,N_14883,N_14829);
and UO_212 (O_212,N_14937,N_14852);
nand UO_213 (O_213,N_14917,N_14963);
nor UO_214 (O_214,N_14829,N_14943);
or UO_215 (O_215,N_14973,N_14921);
nand UO_216 (O_216,N_14907,N_14978);
nor UO_217 (O_217,N_14842,N_14937);
nor UO_218 (O_218,N_14980,N_14839);
nor UO_219 (O_219,N_14948,N_14827);
or UO_220 (O_220,N_14860,N_14938);
nand UO_221 (O_221,N_14900,N_14872);
nor UO_222 (O_222,N_14815,N_14959);
or UO_223 (O_223,N_14861,N_14850);
nor UO_224 (O_224,N_14895,N_14825);
nand UO_225 (O_225,N_14916,N_14838);
xnor UO_226 (O_226,N_14981,N_14877);
and UO_227 (O_227,N_14929,N_14909);
or UO_228 (O_228,N_14892,N_14932);
and UO_229 (O_229,N_14910,N_14911);
nand UO_230 (O_230,N_14872,N_14888);
nor UO_231 (O_231,N_14877,N_14907);
or UO_232 (O_232,N_14802,N_14817);
and UO_233 (O_233,N_14852,N_14833);
xor UO_234 (O_234,N_14946,N_14881);
or UO_235 (O_235,N_14983,N_14960);
nor UO_236 (O_236,N_14877,N_14849);
nand UO_237 (O_237,N_14918,N_14898);
xnor UO_238 (O_238,N_14912,N_14918);
nor UO_239 (O_239,N_14869,N_14865);
nor UO_240 (O_240,N_14830,N_14966);
or UO_241 (O_241,N_14913,N_14818);
or UO_242 (O_242,N_14977,N_14819);
or UO_243 (O_243,N_14899,N_14870);
and UO_244 (O_244,N_14841,N_14940);
or UO_245 (O_245,N_14987,N_14930);
or UO_246 (O_246,N_14843,N_14915);
and UO_247 (O_247,N_14977,N_14828);
nor UO_248 (O_248,N_14918,N_14942);
or UO_249 (O_249,N_14997,N_14903);
xor UO_250 (O_250,N_14806,N_14846);
nor UO_251 (O_251,N_14888,N_14868);
or UO_252 (O_252,N_14917,N_14821);
nor UO_253 (O_253,N_14852,N_14828);
or UO_254 (O_254,N_14874,N_14927);
nor UO_255 (O_255,N_14829,N_14866);
and UO_256 (O_256,N_14894,N_14996);
nand UO_257 (O_257,N_14910,N_14998);
nor UO_258 (O_258,N_14966,N_14803);
and UO_259 (O_259,N_14902,N_14974);
or UO_260 (O_260,N_14991,N_14844);
nand UO_261 (O_261,N_14930,N_14831);
and UO_262 (O_262,N_14875,N_14950);
or UO_263 (O_263,N_14979,N_14850);
and UO_264 (O_264,N_14845,N_14984);
nand UO_265 (O_265,N_14901,N_14855);
and UO_266 (O_266,N_14916,N_14957);
and UO_267 (O_267,N_14856,N_14925);
and UO_268 (O_268,N_14861,N_14841);
nand UO_269 (O_269,N_14862,N_14978);
nand UO_270 (O_270,N_14819,N_14957);
or UO_271 (O_271,N_14826,N_14842);
and UO_272 (O_272,N_14862,N_14973);
and UO_273 (O_273,N_14836,N_14807);
nor UO_274 (O_274,N_14897,N_14932);
nand UO_275 (O_275,N_14881,N_14910);
nor UO_276 (O_276,N_14999,N_14879);
nor UO_277 (O_277,N_14850,N_14987);
nand UO_278 (O_278,N_14868,N_14930);
nand UO_279 (O_279,N_14914,N_14945);
or UO_280 (O_280,N_14882,N_14944);
and UO_281 (O_281,N_14900,N_14841);
xor UO_282 (O_282,N_14821,N_14977);
nor UO_283 (O_283,N_14888,N_14804);
xor UO_284 (O_284,N_14998,N_14965);
nand UO_285 (O_285,N_14963,N_14985);
nor UO_286 (O_286,N_14932,N_14817);
and UO_287 (O_287,N_14897,N_14960);
nor UO_288 (O_288,N_14927,N_14973);
and UO_289 (O_289,N_14855,N_14994);
or UO_290 (O_290,N_14932,N_14840);
or UO_291 (O_291,N_14992,N_14828);
nor UO_292 (O_292,N_14962,N_14887);
nor UO_293 (O_293,N_14981,N_14935);
and UO_294 (O_294,N_14974,N_14820);
and UO_295 (O_295,N_14939,N_14983);
xor UO_296 (O_296,N_14968,N_14983);
nor UO_297 (O_297,N_14806,N_14903);
nor UO_298 (O_298,N_14901,N_14804);
and UO_299 (O_299,N_14890,N_14853);
nor UO_300 (O_300,N_14903,N_14888);
nor UO_301 (O_301,N_14821,N_14909);
and UO_302 (O_302,N_14879,N_14917);
nand UO_303 (O_303,N_14825,N_14943);
or UO_304 (O_304,N_14917,N_14987);
nand UO_305 (O_305,N_14959,N_14910);
xor UO_306 (O_306,N_14903,N_14863);
nand UO_307 (O_307,N_14811,N_14993);
nor UO_308 (O_308,N_14846,N_14871);
or UO_309 (O_309,N_14866,N_14869);
and UO_310 (O_310,N_14887,N_14890);
xnor UO_311 (O_311,N_14939,N_14890);
and UO_312 (O_312,N_14876,N_14839);
and UO_313 (O_313,N_14825,N_14862);
and UO_314 (O_314,N_14898,N_14949);
or UO_315 (O_315,N_14989,N_14847);
or UO_316 (O_316,N_14973,N_14923);
and UO_317 (O_317,N_14936,N_14982);
nor UO_318 (O_318,N_14811,N_14850);
nor UO_319 (O_319,N_14935,N_14820);
nor UO_320 (O_320,N_14910,N_14821);
nand UO_321 (O_321,N_14879,N_14863);
and UO_322 (O_322,N_14961,N_14821);
and UO_323 (O_323,N_14845,N_14847);
nand UO_324 (O_324,N_14973,N_14872);
nand UO_325 (O_325,N_14960,N_14962);
nand UO_326 (O_326,N_14914,N_14880);
and UO_327 (O_327,N_14926,N_14934);
and UO_328 (O_328,N_14885,N_14877);
and UO_329 (O_329,N_14885,N_14961);
nand UO_330 (O_330,N_14968,N_14919);
nor UO_331 (O_331,N_14916,N_14949);
nor UO_332 (O_332,N_14934,N_14952);
nand UO_333 (O_333,N_14853,N_14823);
nor UO_334 (O_334,N_14897,N_14839);
xnor UO_335 (O_335,N_14937,N_14841);
nand UO_336 (O_336,N_14920,N_14879);
nor UO_337 (O_337,N_14944,N_14996);
and UO_338 (O_338,N_14878,N_14973);
nor UO_339 (O_339,N_14876,N_14829);
or UO_340 (O_340,N_14900,N_14972);
xor UO_341 (O_341,N_14898,N_14922);
nor UO_342 (O_342,N_14934,N_14883);
nand UO_343 (O_343,N_14837,N_14960);
or UO_344 (O_344,N_14869,N_14981);
nand UO_345 (O_345,N_14825,N_14853);
and UO_346 (O_346,N_14830,N_14996);
or UO_347 (O_347,N_14933,N_14895);
and UO_348 (O_348,N_14960,N_14814);
or UO_349 (O_349,N_14920,N_14801);
nand UO_350 (O_350,N_14852,N_14947);
nor UO_351 (O_351,N_14909,N_14891);
nor UO_352 (O_352,N_14952,N_14888);
and UO_353 (O_353,N_14936,N_14851);
nand UO_354 (O_354,N_14959,N_14823);
nand UO_355 (O_355,N_14801,N_14928);
and UO_356 (O_356,N_14926,N_14903);
nand UO_357 (O_357,N_14841,N_14859);
or UO_358 (O_358,N_14824,N_14916);
nor UO_359 (O_359,N_14822,N_14917);
and UO_360 (O_360,N_14931,N_14932);
nand UO_361 (O_361,N_14906,N_14894);
nand UO_362 (O_362,N_14899,N_14939);
nand UO_363 (O_363,N_14976,N_14943);
nor UO_364 (O_364,N_14818,N_14910);
nor UO_365 (O_365,N_14918,N_14840);
nand UO_366 (O_366,N_14873,N_14849);
nor UO_367 (O_367,N_14818,N_14981);
nor UO_368 (O_368,N_14816,N_14930);
and UO_369 (O_369,N_14836,N_14809);
nor UO_370 (O_370,N_14959,N_14962);
and UO_371 (O_371,N_14886,N_14862);
and UO_372 (O_372,N_14889,N_14925);
xor UO_373 (O_373,N_14813,N_14824);
or UO_374 (O_374,N_14807,N_14941);
nand UO_375 (O_375,N_14894,N_14819);
and UO_376 (O_376,N_14903,N_14817);
or UO_377 (O_377,N_14857,N_14817);
and UO_378 (O_378,N_14850,N_14865);
nand UO_379 (O_379,N_14833,N_14909);
nor UO_380 (O_380,N_14872,N_14927);
nor UO_381 (O_381,N_14900,N_14913);
xor UO_382 (O_382,N_14938,N_14882);
and UO_383 (O_383,N_14912,N_14887);
nor UO_384 (O_384,N_14992,N_14931);
and UO_385 (O_385,N_14978,N_14837);
nand UO_386 (O_386,N_14818,N_14927);
nand UO_387 (O_387,N_14913,N_14974);
xor UO_388 (O_388,N_14879,N_14927);
nor UO_389 (O_389,N_14965,N_14842);
nor UO_390 (O_390,N_14975,N_14910);
and UO_391 (O_391,N_14838,N_14886);
and UO_392 (O_392,N_14881,N_14964);
or UO_393 (O_393,N_14965,N_14983);
and UO_394 (O_394,N_14802,N_14985);
nand UO_395 (O_395,N_14948,N_14992);
nor UO_396 (O_396,N_14994,N_14851);
and UO_397 (O_397,N_14878,N_14961);
nand UO_398 (O_398,N_14880,N_14834);
xnor UO_399 (O_399,N_14827,N_14952);
nand UO_400 (O_400,N_14827,N_14812);
nor UO_401 (O_401,N_14980,N_14938);
nand UO_402 (O_402,N_14821,N_14823);
and UO_403 (O_403,N_14899,N_14844);
nor UO_404 (O_404,N_14845,N_14854);
nor UO_405 (O_405,N_14850,N_14872);
nand UO_406 (O_406,N_14869,N_14915);
or UO_407 (O_407,N_14820,N_14875);
and UO_408 (O_408,N_14939,N_14835);
and UO_409 (O_409,N_14970,N_14929);
nand UO_410 (O_410,N_14801,N_14873);
nand UO_411 (O_411,N_14960,N_14980);
xor UO_412 (O_412,N_14811,N_14869);
xnor UO_413 (O_413,N_14919,N_14951);
nor UO_414 (O_414,N_14853,N_14926);
nand UO_415 (O_415,N_14902,N_14957);
or UO_416 (O_416,N_14802,N_14906);
nor UO_417 (O_417,N_14806,N_14937);
nand UO_418 (O_418,N_14873,N_14953);
and UO_419 (O_419,N_14985,N_14828);
or UO_420 (O_420,N_14822,N_14926);
or UO_421 (O_421,N_14894,N_14813);
and UO_422 (O_422,N_14972,N_14911);
or UO_423 (O_423,N_14830,N_14928);
nor UO_424 (O_424,N_14973,N_14802);
xnor UO_425 (O_425,N_14894,N_14915);
or UO_426 (O_426,N_14975,N_14998);
nand UO_427 (O_427,N_14873,N_14851);
xnor UO_428 (O_428,N_14874,N_14869);
nor UO_429 (O_429,N_14894,N_14907);
or UO_430 (O_430,N_14872,N_14964);
nor UO_431 (O_431,N_14982,N_14991);
nand UO_432 (O_432,N_14992,N_14999);
nand UO_433 (O_433,N_14970,N_14810);
and UO_434 (O_434,N_14846,N_14983);
or UO_435 (O_435,N_14955,N_14800);
nand UO_436 (O_436,N_14856,N_14913);
nor UO_437 (O_437,N_14933,N_14857);
or UO_438 (O_438,N_14851,N_14935);
or UO_439 (O_439,N_14808,N_14875);
and UO_440 (O_440,N_14875,N_14836);
nor UO_441 (O_441,N_14822,N_14967);
xnor UO_442 (O_442,N_14903,N_14808);
nor UO_443 (O_443,N_14940,N_14835);
or UO_444 (O_444,N_14888,N_14974);
and UO_445 (O_445,N_14828,N_14966);
xnor UO_446 (O_446,N_14927,N_14943);
nor UO_447 (O_447,N_14832,N_14823);
xnor UO_448 (O_448,N_14819,N_14906);
or UO_449 (O_449,N_14909,N_14917);
nand UO_450 (O_450,N_14934,N_14862);
or UO_451 (O_451,N_14928,N_14875);
xor UO_452 (O_452,N_14809,N_14900);
or UO_453 (O_453,N_14898,N_14805);
or UO_454 (O_454,N_14871,N_14839);
or UO_455 (O_455,N_14940,N_14895);
and UO_456 (O_456,N_14902,N_14925);
and UO_457 (O_457,N_14851,N_14981);
and UO_458 (O_458,N_14952,N_14985);
nor UO_459 (O_459,N_14839,N_14878);
nand UO_460 (O_460,N_14801,N_14931);
nor UO_461 (O_461,N_14966,N_14809);
nand UO_462 (O_462,N_14878,N_14882);
and UO_463 (O_463,N_14974,N_14813);
xor UO_464 (O_464,N_14893,N_14909);
nor UO_465 (O_465,N_14820,N_14940);
nor UO_466 (O_466,N_14906,N_14865);
and UO_467 (O_467,N_14810,N_14862);
or UO_468 (O_468,N_14994,N_14879);
nor UO_469 (O_469,N_14902,N_14845);
or UO_470 (O_470,N_14930,N_14910);
nand UO_471 (O_471,N_14876,N_14865);
nand UO_472 (O_472,N_14970,N_14973);
and UO_473 (O_473,N_14804,N_14970);
nand UO_474 (O_474,N_14852,N_14803);
and UO_475 (O_475,N_14866,N_14923);
nand UO_476 (O_476,N_14840,N_14848);
and UO_477 (O_477,N_14922,N_14877);
nand UO_478 (O_478,N_14830,N_14884);
nand UO_479 (O_479,N_14843,N_14994);
nor UO_480 (O_480,N_14999,N_14868);
or UO_481 (O_481,N_14849,N_14800);
or UO_482 (O_482,N_14985,N_14976);
nand UO_483 (O_483,N_14914,N_14881);
and UO_484 (O_484,N_14920,N_14916);
nor UO_485 (O_485,N_14967,N_14881);
and UO_486 (O_486,N_14972,N_14901);
xnor UO_487 (O_487,N_14995,N_14948);
nor UO_488 (O_488,N_14971,N_14872);
nand UO_489 (O_489,N_14983,N_14810);
nor UO_490 (O_490,N_14977,N_14945);
nor UO_491 (O_491,N_14816,N_14892);
nand UO_492 (O_492,N_14869,N_14940);
nor UO_493 (O_493,N_14811,N_14802);
xor UO_494 (O_494,N_14944,N_14855);
or UO_495 (O_495,N_14899,N_14831);
xnor UO_496 (O_496,N_14883,N_14936);
nand UO_497 (O_497,N_14921,N_14900);
xnor UO_498 (O_498,N_14847,N_14910);
or UO_499 (O_499,N_14858,N_14956);
nand UO_500 (O_500,N_14988,N_14821);
nor UO_501 (O_501,N_14805,N_14908);
xor UO_502 (O_502,N_14805,N_14858);
nand UO_503 (O_503,N_14821,N_14852);
nor UO_504 (O_504,N_14907,N_14960);
nor UO_505 (O_505,N_14973,N_14808);
nor UO_506 (O_506,N_14951,N_14846);
nand UO_507 (O_507,N_14971,N_14873);
or UO_508 (O_508,N_14965,N_14956);
nand UO_509 (O_509,N_14876,N_14982);
or UO_510 (O_510,N_14942,N_14951);
or UO_511 (O_511,N_14832,N_14933);
or UO_512 (O_512,N_14930,N_14850);
nand UO_513 (O_513,N_14849,N_14832);
xnor UO_514 (O_514,N_14961,N_14820);
nand UO_515 (O_515,N_14926,N_14826);
nand UO_516 (O_516,N_14959,N_14827);
and UO_517 (O_517,N_14812,N_14989);
or UO_518 (O_518,N_14816,N_14959);
or UO_519 (O_519,N_14942,N_14814);
nor UO_520 (O_520,N_14803,N_14918);
nor UO_521 (O_521,N_14880,N_14937);
and UO_522 (O_522,N_14878,N_14967);
nor UO_523 (O_523,N_14801,N_14912);
xor UO_524 (O_524,N_14860,N_14822);
nor UO_525 (O_525,N_14972,N_14921);
xnor UO_526 (O_526,N_14877,N_14838);
and UO_527 (O_527,N_14834,N_14806);
nor UO_528 (O_528,N_14814,N_14930);
xnor UO_529 (O_529,N_14890,N_14822);
xnor UO_530 (O_530,N_14816,N_14972);
or UO_531 (O_531,N_14987,N_14975);
or UO_532 (O_532,N_14889,N_14973);
or UO_533 (O_533,N_14882,N_14964);
nor UO_534 (O_534,N_14913,N_14885);
and UO_535 (O_535,N_14812,N_14801);
and UO_536 (O_536,N_14984,N_14858);
nand UO_537 (O_537,N_14973,N_14894);
and UO_538 (O_538,N_14956,N_14982);
xor UO_539 (O_539,N_14888,N_14824);
nor UO_540 (O_540,N_14861,N_14842);
or UO_541 (O_541,N_14948,N_14996);
and UO_542 (O_542,N_14873,N_14822);
or UO_543 (O_543,N_14850,N_14887);
nand UO_544 (O_544,N_14872,N_14947);
or UO_545 (O_545,N_14806,N_14875);
nand UO_546 (O_546,N_14827,N_14976);
nor UO_547 (O_547,N_14867,N_14952);
nand UO_548 (O_548,N_14921,N_14907);
and UO_549 (O_549,N_14874,N_14842);
nor UO_550 (O_550,N_14864,N_14808);
or UO_551 (O_551,N_14989,N_14988);
xor UO_552 (O_552,N_14829,N_14907);
and UO_553 (O_553,N_14944,N_14864);
and UO_554 (O_554,N_14852,N_14942);
xnor UO_555 (O_555,N_14983,N_14936);
nand UO_556 (O_556,N_14832,N_14890);
nand UO_557 (O_557,N_14962,N_14920);
or UO_558 (O_558,N_14833,N_14916);
and UO_559 (O_559,N_14954,N_14869);
nor UO_560 (O_560,N_14834,N_14918);
or UO_561 (O_561,N_14832,N_14847);
nand UO_562 (O_562,N_14843,N_14927);
and UO_563 (O_563,N_14933,N_14943);
and UO_564 (O_564,N_14946,N_14943);
or UO_565 (O_565,N_14977,N_14846);
and UO_566 (O_566,N_14939,N_14884);
and UO_567 (O_567,N_14842,N_14864);
and UO_568 (O_568,N_14908,N_14855);
and UO_569 (O_569,N_14894,N_14991);
and UO_570 (O_570,N_14919,N_14895);
and UO_571 (O_571,N_14991,N_14990);
or UO_572 (O_572,N_14967,N_14897);
nand UO_573 (O_573,N_14992,N_14942);
nand UO_574 (O_574,N_14881,N_14878);
or UO_575 (O_575,N_14915,N_14973);
nor UO_576 (O_576,N_14955,N_14892);
and UO_577 (O_577,N_14937,N_14952);
or UO_578 (O_578,N_14857,N_14828);
nor UO_579 (O_579,N_14892,N_14978);
nand UO_580 (O_580,N_14852,N_14892);
or UO_581 (O_581,N_14848,N_14872);
nand UO_582 (O_582,N_14937,N_14901);
nand UO_583 (O_583,N_14979,N_14885);
nor UO_584 (O_584,N_14923,N_14817);
xor UO_585 (O_585,N_14907,N_14821);
xnor UO_586 (O_586,N_14967,N_14935);
and UO_587 (O_587,N_14800,N_14993);
nor UO_588 (O_588,N_14886,N_14954);
nand UO_589 (O_589,N_14895,N_14837);
and UO_590 (O_590,N_14844,N_14831);
or UO_591 (O_591,N_14998,N_14992);
or UO_592 (O_592,N_14934,N_14946);
nand UO_593 (O_593,N_14892,N_14967);
nor UO_594 (O_594,N_14974,N_14968);
nor UO_595 (O_595,N_14896,N_14949);
nor UO_596 (O_596,N_14832,N_14910);
and UO_597 (O_597,N_14858,N_14901);
xnor UO_598 (O_598,N_14873,N_14820);
nand UO_599 (O_599,N_14947,N_14961);
and UO_600 (O_600,N_14955,N_14918);
nor UO_601 (O_601,N_14829,N_14998);
nor UO_602 (O_602,N_14967,N_14901);
or UO_603 (O_603,N_14847,N_14929);
xnor UO_604 (O_604,N_14871,N_14955);
nor UO_605 (O_605,N_14911,N_14971);
nor UO_606 (O_606,N_14970,N_14852);
nor UO_607 (O_607,N_14972,N_14894);
nor UO_608 (O_608,N_14859,N_14844);
or UO_609 (O_609,N_14900,N_14937);
nand UO_610 (O_610,N_14818,N_14974);
nor UO_611 (O_611,N_14871,N_14850);
nor UO_612 (O_612,N_14945,N_14935);
nand UO_613 (O_613,N_14904,N_14920);
or UO_614 (O_614,N_14948,N_14892);
nand UO_615 (O_615,N_14973,N_14982);
nor UO_616 (O_616,N_14910,N_14994);
or UO_617 (O_617,N_14960,N_14900);
nor UO_618 (O_618,N_14864,N_14800);
nor UO_619 (O_619,N_14869,N_14999);
nand UO_620 (O_620,N_14970,N_14942);
xor UO_621 (O_621,N_14940,N_14897);
nand UO_622 (O_622,N_14851,N_14830);
nand UO_623 (O_623,N_14846,N_14992);
nand UO_624 (O_624,N_14835,N_14805);
xnor UO_625 (O_625,N_14941,N_14882);
nand UO_626 (O_626,N_14994,N_14902);
and UO_627 (O_627,N_14978,N_14941);
nand UO_628 (O_628,N_14968,N_14847);
and UO_629 (O_629,N_14872,N_14857);
and UO_630 (O_630,N_14911,N_14895);
and UO_631 (O_631,N_14860,N_14887);
or UO_632 (O_632,N_14916,N_14938);
nand UO_633 (O_633,N_14997,N_14994);
or UO_634 (O_634,N_14817,N_14937);
xnor UO_635 (O_635,N_14900,N_14831);
nor UO_636 (O_636,N_14876,N_14984);
or UO_637 (O_637,N_14858,N_14983);
nand UO_638 (O_638,N_14886,N_14865);
nor UO_639 (O_639,N_14975,N_14913);
nor UO_640 (O_640,N_14807,N_14841);
and UO_641 (O_641,N_14900,N_14962);
or UO_642 (O_642,N_14800,N_14984);
xor UO_643 (O_643,N_14928,N_14904);
and UO_644 (O_644,N_14992,N_14981);
or UO_645 (O_645,N_14955,N_14886);
and UO_646 (O_646,N_14870,N_14918);
and UO_647 (O_647,N_14915,N_14956);
nand UO_648 (O_648,N_14990,N_14955);
nand UO_649 (O_649,N_14948,N_14943);
nor UO_650 (O_650,N_14810,N_14828);
nand UO_651 (O_651,N_14808,N_14910);
nand UO_652 (O_652,N_14958,N_14978);
nor UO_653 (O_653,N_14863,N_14938);
or UO_654 (O_654,N_14813,N_14995);
and UO_655 (O_655,N_14979,N_14953);
nor UO_656 (O_656,N_14914,N_14857);
or UO_657 (O_657,N_14951,N_14890);
and UO_658 (O_658,N_14945,N_14823);
nor UO_659 (O_659,N_14804,N_14803);
nor UO_660 (O_660,N_14809,N_14802);
and UO_661 (O_661,N_14901,N_14936);
or UO_662 (O_662,N_14880,N_14964);
or UO_663 (O_663,N_14839,N_14873);
nor UO_664 (O_664,N_14845,N_14939);
nand UO_665 (O_665,N_14979,N_14935);
nor UO_666 (O_666,N_14955,N_14865);
and UO_667 (O_667,N_14948,N_14824);
or UO_668 (O_668,N_14904,N_14901);
or UO_669 (O_669,N_14880,N_14841);
or UO_670 (O_670,N_14859,N_14977);
and UO_671 (O_671,N_14958,N_14810);
xnor UO_672 (O_672,N_14974,N_14830);
and UO_673 (O_673,N_14990,N_14903);
xnor UO_674 (O_674,N_14886,N_14859);
or UO_675 (O_675,N_14861,N_14839);
and UO_676 (O_676,N_14912,N_14967);
nor UO_677 (O_677,N_14861,N_14922);
nor UO_678 (O_678,N_14985,N_14913);
or UO_679 (O_679,N_14863,N_14833);
and UO_680 (O_680,N_14938,N_14826);
or UO_681 (O_681,N_14830,N_14813);
nor UO_682 (O_682,N_14984,N_14881);
and UO_683 (O_683,N_14829,N_14863);
and UO_684 (O_684,N_14929,N_14992);
or UO_685 (O_685,N_14850,N_14876);
and UO_686 (O_686,N_14819,N_14841);
and UO_687 (O_687,N_14974,N_14814);
nor UO_688 (O_688,N_14800,N_14945);
and UO_689 (O_689,N_14827,N_14970);
or UO_690 (O_690,N_14807,N_14817);
nor UO_691 (O_691,N_14885,N_14872);
nor UO_692 (O_692,N_14884,N_14852);
xnor UO_693 (O_693,N_14883,N_14941);
and UO_694 (O_694,N_14801,N_14829);
nor UO_695 (O_695,N_14813,N_14893);
or UO_696 (O_696,N_14881,N_14833);
and UO_697 (O_697,N_14898,N_14884);
nor UO_698 (O_698,N_14816,N_14933);
nor UO_699 (O_699,N_14928,N_14923);
and UO_700 (O_700,N_14966,N_14857);
or UO_701 (O_701,N_14821,N_14941);
and UO_702 (O_702,N_14960,N_14912);
nand UO_703 (O_703,N_14896,N_14846);
and UO_704 (O_704,N_14888,N_14985);
nor UO_705 (O_705,N_14824,N_14843);
or UO_706 (O_706,N_14958,N_14996);
or UO_707 (O_707,N_14862,N_14931);
nand UO_708 (O_708,N_14821,N_14965);
and UO_709 (O_709,N_14862,N_14983);
and UO_710 (O_710,N_14863,N_14843);
nor UO_711 (O_711,N_14976,N_14856);
and UO_712 (O_712,N_14920,N_14808);
xnor UO_713 (O_713,N_14926,N_14824);
nor UO_714 (O_714,N_14865,N_14949);
nor UO_715 (O_715,N_14834,N_14882);
or UO_716 (O_716,N_14951,N_14852);
and UO_717 (O_717,N_14816,N_14840);
or UO_718 (O_718,N_14859,N_14820);
nand UO_719 (O_719,N_14920,N_14811);
nand UO_720 (O_720,N_14841,N_14944);
or UO_721 (O_721,N_14863,N_14876);
or UO_722 (O_722,N_14852,N_14979);
nand UO_723 (O_723,N_14907,N_14892);
nand UO_724 (O_724,N_14874,N_14864);
or UO_725 (O_725,N_14971,N_14952);
or UO_726 (O_726,N_14811,N_14884);
nand UO_727 (O_727,N_14885,N_14804);
nand UO_728 (O_728,N_14941,N_14836);
nand UO_729 (O_729,N_14929,N_14878);
or UO_730 (O_730,N_14882,N_14896);
nor UO_731 (O_731,N_14870,N_14891);
nand UO_732 (O_732,N_14839,N_14930);
and UO_733 (O_733,N_14811,N_14881);
and UO_734 (O_734,N_14899,N_14856);
nor UO_735 (O_735,N_14979,N_14983);
nand UO_736 (O_736,N_14952,N_14955);
nand UO_737 (O_737,N_14835,N_14928);
and UO_738 (O_738,N_14835,N_14969);
xnor UO_739 (O_739,N_14934,N_14814);
and UO_740 (O_740,N_14918,N_14915);
xor UO_741 (O_741,N_14826,N_14819);
nor UO_742 (O_742,N_14808,N_14851);
nand UO_743 (O_743,N_14950,N_14897);
or UO_744 (O_744,N_14854,N_14846);
nor UO_745 (O_745,N_14957,N_14829);
or UO_746 (O_746,N_14982,N_14803);
nand UO_747 (O_747,N_14901,N_14929);
or UO_748 (O_748,N_14893,N_14888);
nand UO_749 (O_749,N_14900,N_14882);
nor UO_750 (O_750,N_14952,N_14860);
nor UO_751 (O_751,N_14836,N_14889);
or UO_752 (O_752,N_14886,N_14982);
nand UO_753 (O_753,N_14833,N_14889);
nor UO_754 (O_754,N_14975,N_14894);
nand UO_755 (O_755,N_14946,N_14833);
and UO_756 (O_756,N_14810,N_14937);
nand UO_757 (O_757,N_14949,N_14864);
or UO_758 (O_758,N_14925,N_14967);
and UO_759 (O_759,N_14924,N_14926);
nand UO_760 (O_760,N_14886,N_14958);
xnor UO_761 (O_761,N_14834,N_14937);
nand UO_762 (O_762,N_14933,N_14968);
xnor UO_763 (O_763,N_14877,N_14987);
or UO_764 (O_764,N_14800,N_14916);
xor UO_765 (O_765,N_14952,N_14950);
or UO_766 (O_766,N_14951,N_14994);
and UO_767 (O_767,N_14855,N_14805);
or UO_768 (O_768,N_14858,N_14887);
nand UO_769 (O_769,N_14847,N_14867);
and UO_770 (O_770,N_14826,N_14987);
nor UO_771 (O_771,N_14820,N_14983);
nor UO_772 (O_772,N_14885,N_14892);
xor UO_773 (O_773,N_14896,N_14847);
nor UO_774 (O_774,N_14801,N_14845);
and UO_775 (O_775,N_14861,N_14936);
xnor UO_776 (O_776,N_14991,N_14865);
nand UO_777 (O_777,N_14975,N_14917);
nand UO_778 (O_778,N_14833,N_14800);
nand UO_779 (O_779,N_14997,N_14998);
or UO_780 (O_780,N_14962,N_14992);
nor UO_781 (O_781,N_14829,N_14936);
nor UO_782 (O_782,N_14966,N_14884);
and UO_783 (O_783,N_14933,N_14913);
nor UO_784 (O_784,N_14937,N_14991);
or UO_785 (O_785,N_14888,N_14835);
xor UO_786 (O_786,N_14816,N_14969);
nand UO_787 (O_787,N_14884,N_14977);
and UO_788 (O_788,N_14899,N_14874);
and UO_789 (O_789,N_14998,N_14866);
and UO_790 (O_790,N_14903,N_14913);
nand UO_791 (O_791,N_14827,N_14842);
and UO_792 (O_792,N_14818,N_14973);
nand UO_793 (O_793,N_14814,N_14947);
nand UO_794 (O_794,N_14929,N_14998);
and UO_795 (O_795,N_14842,N_14939);
nor UO_796 (O_796,N_14855,N_14928);
or UO_797 (O_797,N_14900,N_14869);
and UO_798 (O_798,N_14994,N_14865);
or UO_799 (O_799,N_14925,N_14899);
and UO_800 (O_800,N_14903,N_14849);
nand UO_801 (O_801,N_14801,N_14886);
nand UO_802 (O_802,N_14826,N_14983);
nand UO_803 (O_803,N_14862,N_14880);
nor UO_804 (O_804,N_14979,N_14952);
and UO_805 (O_805,N_14856,N_14919);
or UO_806 (O_806,N_14905,N_14809);
nor UO_807 (O_807,N_14898,N_14811);
nand UO_808 (O_808,N_14903,N_14886);
nor UO_809 (O_809,N_14841,N_14856);
nand UO_810 (O_810,N_14926,N_14959);
xnor UO_811 (O_811,N_14853,N_14971);
xor UO_812 (O_812,N_14950,N_14986);
nor UO_813 (O_813,N_14982,N_14836);
xor UO_814 (O_814,N_14850,N_14841);
nor UO_815 (O_815,N_14937,N_14800);
nand UO_816 (O_816,N_14981,N_14908);
nand UO_817 (O_817,N_14899,N_14903);
nor UO_818 (O_818,N_14944,N_14820);
nor UO_819 (O_819,N_14890,N_14841);
and UO_820 (O_820,N_14916,N_14847);
and UO_821 (O_821,N_14919,N_14887);
nor UO_822 (O_822,N_14940,N_14998);
and UO_823 (O_823,N_14848,N_14906);
and UO_824 (O_824,N_14958,N_14801);
nand UO_825 (O_825,N_14819,N_14825);
nor UO_826 (O_826,N_14864,N_14915);
and UO_827 (O_827,N_14884,N_14923);
or UO_828 (O_828,N_14892,N_14959);
xnor UO_829 (O_829,N_14879,N_14830);
nor UO_830 (O_830,N_14861,N_14881);
or UO_831 (O_831,N_14890,N_14844);
and UO_832 (O_832,N_14952,N_14978);
xor UO_833 (O_833,N_14979,N_14940);
nand UO_834 (O_834,N_14953,N_14915);
xnor UO_835 (O_835,N_14972,N_14815);
or UO_836 (O_836,N_14994,N_14947);
nand UO_837 (O_837,N_14912,N_14800);
or UO_838 (O_838,N_14873,N_14867);
nor UO_839 (O_839,N_14813,N_14967);
xor UO_840 (O_840,N_14954,N_14925);
and UO_841 (O_841,N_14875,N_14815);
nand UO_842 (O_842,N_14914,N_14837);
or UO_843 (O_843,N_14913,N_14896);
xor UO_844 (O_844,N_14835,N_14867);
nand UO_845 (O_845,N_14992,N_14987);
nor UO_846 (O_846,N_14963,N_14915);
nand UO_847 (O_847,N_14967,N_14844);
nand UO_848 (O_848,N_14843,N_14917);
xnor UO_849 (O_849,N_14878,N_14801);
nand UO_850 (O_850,N_14986,N_14973);
or UO_851 (O_851,N_14813,N_14899);
and UO_852 (O_852,N_14924,N_14979);
and UO_853 (O_853,N_14885,N_14822);
nor UO_854 (O_854,N_14850,N_14943);
or UO_855 (O_855,N_14857,N_14996);
and UO_856 (O_856,N_14856,N_14985);
nor UO_857 (O_857,N_14801,N_14948);
or UO_858 (O_858,N_14815,N_14920);
or UO_859 (O_859,N_14898,N_14850);
xor UO_860 (O_860,N_14887,N_14953);
and UO_861 (O_861,N_14957,N_14915);
nand UO_862 (O_862,N_14927,N_14856);
xnor UO_863 (O_863,N_14970,N_14850);
and UO_864 (O_864,N_14961,N_14883);
nor UO_865 (O_865,N_14989,N_14961);
and UO_866 (O_866,N_14803,N_14858);
or UO_867 (O_867,N_14885,N_14999);
nor UO_868 (O_868,N_14903,N_14988);
or UO_869 (O_869,N_14948,N_14886);
and UO_870 (O_870,N_14931,N_14982);
or UO_871 (O_871,N_14805,N_14938);
and UO_872 (O_872,N_14902,N_14968);
nand UO_873 (O_873,N_14934,N_14944);
nand UO_874 (O_874,N_14926,N_14865);
and UO_875 (O_875,N_14846,N_14885);
and UO_876 (O_876,N_14891,N_14960);
or UO_877 (O_877,N_14857,N_14984);
nand UO_878 (O_878,N_14876,N_14809);
and UO_879 (O_879,N_14886,N_14943);
nor UO_880 (O_880,N_14836,N_14930);
or UO_881 (O_881,N_14895,N_14920);
nor UO_882 (O_882,N_14971,N_14846);
and UO_883 (O_883,N_14837,N_14918);
or UO_884 (O_884,N_14858,N_14949);
and UO_885 (O_885,N_14967,N_14928);
nor UO_886 (O_886,N_14852,N_14929);
xor UO_887 (O_887,N_14887,N_14957);
nand UO_888 (O_888,N_14887,N_14898);
nor UO_889 (O_889,N_14942,N_14936);
or UO_890 (O_890,N_14961,N_14905);
and UO_891 (O_891,N_14821,N_14951);
and UO_892 (O_892,N_14935,N_14838);
and UO_893 (O_893,N_14900,N_14893);
or UO_894 (O_894,N_14864,N_14973);
or UO_895 (O_895,N_14810,N_14894);
xor UO_896 (O_896,N_14832,N_14846);
or UO_897 (O_897,N_14930,N_14976);
xnor UO_898 (O_898,N_14830,N_14950);
and UO_899 (O_899,N_14942,N_14967);
nand UO_900 (O_900,N_14911,N_14938);
nand UO_901 (O_901,N_14935,N_14859);
or UO_902 (O_902,N_14808,N_14955);
nand UO_903 (O_903,N_14955,N_14927);
or UO_904 (O_904,N_14857,N_14943);
or UO_905 (O_905,N_14960,N_14959);
xnor UO_906 (O_906,N_14940,N_14852);
or UO_907 (O_907,N_14914,N_14808);
nand UO_908 (O_908,N_14923,N_14803);
nand UO_909 (O_909,N_14954,N_14974);
nor UO_910 (O_910,N_14893,N_14981);
and UO_911 (O_911,N_14879,N_14838);
nor UO_912 (O_912,N_14826,N_14910);
or UO_913 (O_913,N_14955,N_14994);
and UO_914 (O_914,N_14856,N_14884);
or UO_915 (O_915,N_14836,N_14909);
and UO_916 (O_916,N_14854,N_14961);
nor UO_917 (O_917,N_14894,N_14969);
nor UO_918 (O_918,N_14966,N_14907);
nand UO_919 (O_919,N_14958,N_14868);
and UO_920 (O_920,N_14801,N_14911);
nor UO_921 (O_921,N_14941,N_14951);
or UO_922 (O_922,N_14929,N_14884);
nor UO_923 (O_923,N_14915,N_14809);
and UO_924 (O_924,N_14800,N_14932);
nand UO_925 (O_925,N_14827,N_14805);
or UO_926 (O_926,N_14824,N_14907);
nor UO_927 (O_927,N_14811,N_14926);
or UO_928 (O_928,N_14987,N_14897);
and UO_929 (O_929,N_14993,N_14852);
and UO_930 (O_930,N_14917,N_14964);
or UO_931 (O_931,N_14991,N_14954);
and UO_932 (O_932,N_14946,N_14915);
nand UO_933 (O_933,N_14992,N_14888);
and UO_934 (O_934,N_14974,N_14943);
or UO_935 (O_935,N_14888,N_14949);
nor UO_936 (O_936,N_14953,N_14960);
and UO_937 (O_937,N_14820,N_14867);
nand UO_938 (O_938,N_14822,N_14832);
and UO_939 (O_939,N_14999,N_14846);
nand UO_940 (O_940,N_14979,N_14925);
nor UO_941 (O_941,N_14973,N_14929);
xnor UO_942 (O_942,N_14972,N_14949);
and UO_943 (O_943,N_14973,N_14985);
or UO_944 (O_944,N_14888,N_14928);
nand UO_945 (O_945,N_14969,N_14945);
and UO_946 (O_946,N_14959,N_14915);
nand UO_947 (O_947,N_14911,N_14956);
xor UO_948 (O_948,N_14981,N_14963);
nor UO_949 (O_949,N_14920,N_14954);
nor UO_950 (O_950,N_14883,N_14972);
nor UO_951 (O_951,N_14927,N_14976);
xnor UO_952 (O_952,N_14860,N_14812);
xor UO_953 (O_953,N_14865,N_14838);
and UO_954 (O_954,N_14817,N_14827);
and UO_955 (O_955,N_14884,N_14930);
or UO_956 (O_956,N_14954,N_14862);
nor UO_957 (O_957,N_14844,N_14829);
nor UO_958 (O_958,N_14935,N_14887);
nor UO_959 (O_959,N_14926,N_14897);
nand UO_960 (O_960,N_14890,N_14843);
and UO_961 (O_961,N_14891,N_14894);
nor UO_962 (O_962,N_14964,N_14811);
or UO_963 (O_963,N_14917,N_14876);
or UO_964 (O_964,N_14969,N_14958);
xnor UO_965 (O_965,N_14984,N_14829);
and UO_966 (O_966,N_14850,N_14915);
or UO_967 (O_967,N_14853,N_14954);
nor UO_968 (O_968,N_14857,N_14963);
nand UO_969 (O_969,N_14826,N_14889);
and UO_970 (O_970,N_14986,N_14808);
and UO_971 (O_971,N_14840,N_14875);
xor UO_972 (O_972,N_14939,N_14856);
or UO_973 (O_973,N_14851,N_14953);
nor UO_974 (O_974,N_14928,N_14978);
and UO_975 (O_975,N_14882,N_14961);
nand UO_976 (O_976,N_14877,N_14928);
nand UO_977 (O_977,N_14890,N_14829);
nor UO_978 (O_978,N_14990,N_14998);
nand UO_979 (O_979,N_14871,N_14804);
or UO_980 (O_980,N_14858,N_14966);
nor UO_981 (O_981,N_14876,N_14873);
nand UO_982 (O_982,N_14892,N_14981);
nand UO_983 (O_983,N_14843,N_14822);
xnor UO_984 (O_984,N_14900,N_14862);
xor UO_985 (O_985,N_14980,N_14973);
and UO_986 (O_986,N_14861,N_14949);
nand UO_987 (O_987,N_14972,N_14964);
and UO_988 (O_988,N_14870,N_14838);
and UO_989 (O_989,N_14942,N_14999);
and UO_990 (O_990,N_14955,N_14872);
nand UO_991 (O_991,N_14946,N_14966);
nor UO_992 (O_992,N_14974,N_14878);
nand UO_993 (O_993,N_14969,N_14952);
nor UO_994 (O_994,N_14888,N_14918);
nor UO_995 (O_995,N_14929,N_14999);
nor UO_996 (O_996,N_14969,N_14859);
or UO_997 (O_997,N_14934,N_14851);
nand UO_998 (O_998,N_14843,N_14858);
or UO_999 (O_999,N_14997,N_14968);
nand UO_1000 (O_1000,N_14979,N_14875);
and UO_1001 (O_1001,N_14806,N_14941);
nor UO_1002 (O_1002,N_14954,N_14906);
or UO_1003 (O_1003,N_14871,N_14941);
or UO_1004 (O_1004,N_14838,N_14868);
nand UO_1005 (O_1005,N_14849,N_14806);
and UO_1006 (O_1006,N_14841,N_14921);
or UO_1007 (O_1007,N_14871,N_14970);
xnor UO_1008 (O_1008,N_14836,N_14912);
or UO_1009 (O_1009,N_14926,N_14928);
and UO_1010 (O_1010,N_14966,N_14832);
nand UO_1011 (O_1011,N_14887,N_14855);
or UO_1012 (O_1012,N_14968,N_14908);
nand UO_1013 (O_1013,N_14808,N_14844);
nor UO_1014 (O_1014,N_14947,N_14996);
or UO_1015 (O_1015,N_14988,N_14888);
xnor UO_1016 (O_1016,N_14906,N_14835);
nand UO_1017 (O_1017,N_14928,N_14996);
or UO_1018 (O_1018,N_14848,N_14957);
nand UO_1019 (O_1019,N_14936,N_14932);
and UO_1020 (O_1020,N_14993,N_14887);
nor UO_1021 (O_1021,N_14847,N_14814);
nor UO_1022 (O_1022,N_14917,N_14888);
and UO_1023 (O_1023,N_14854,N_14815);
or UO_1024 (O_1024,N_14907,N_14983);
and UO_1025 (O_1025,N_14888,N_14857);
nand UO_1026 (O_1026,N_14870,N_14977);
and UO_1027 (O_1027,N_14941,N_14904);
or UO_1028 (O_1028,N_14867,N_14866);
and UO_1029 (O_1029,N_14832,N_14956);
nor UO_1030 (O_1030,N_14988,N_14920);
and UO_1031 (O_1031,N_14925,N_14832);
or UO_1032 (O_1032,N_14954,N_14826);
nor UO_1033 (O_1033,N_14927,N_14864);
or UO_1034 (O_1034,N_14838,N_14921);
nand UO_1035 (O_1035,N_14864,N_14821);
and UO_1036 (O_1036,N_14856,N_14852);
or UO_1037 (O_1037,N_14989,N_14864);
or UO_1038 (O_1038,N_14967,N_14946);
or UO_1039 (O_1039,N_14836,N_14867);
nor UO_1040 (O_1040,N_14854,N_14865);
and UO_1041 (O_1041,N_14982,N_14812);
nor UO_1042 (O_1042,N_14957,N_14964);
nor UO_1043 (O_1043,N_14962,N_14803);
nand UO_1044 (O_1044,N_14959,N_14802);
xnor UO_1045 (O_1045,N_14921,N_14815);
nor UO_1046 (O_1046,N_14948,N_14927);
nor UO_1047 (O_1047,N_14998,N_14971);
and UO_1048 (O_1048,N_14809,N_14825);
nand UO_1049 (O_1049,N_14995,N_14849);
nand UO_1050 (O_1050,N_14958,N_14841);
nand UO_1051 (O_1051,N_14989,N_14870);
and UO_1052 (O_1052,N_14956,N_14960);
nand UO_1053 (O_1053,N_14825,N_14841);
nor UO_1054 (O_1054,N_14948,N_14859);
and UO_1055 (O_1055,N_14911,N_14951);
nor UO_1056 (O_1056,N_14856,N_14930);
nor UO_1057 (O_1057,N_14872,N_14997);
xor UO_1058 (O_1058,N_14867,N_14852);
nand UO_1059 (O_1059,N_14809,N_14816);
and UO_1060 (O_1060,N_14959,N_14981);
nor UO_1061 (O_1061,N_14856,N_14901);
or UO_1062 (O_1062,N_14814,N_14980);
or UO_1063 (O_1063,N_14920,N_14969);
and UO_1064 (O_1064,N_14974,N_14846);
xor UO_1065 (O_1065,N_14967,N_14970);
nand UO_1066 (O_1066,N_14842,N_14948);
or UO_1067 (O_1067,N_14925,N_14851);
nand UO_1068 (O_1068,N_14980,N_14895);
and UO_1069 (O_1069,N_14888,N_14966);
xnor UO_1070 (O_1070,N_14939,N_14860);
nor UO_1071 (O_1071,N_14880,N_14971);
and UO_1072 (O_1072,N_14912,N_14943);
and UO_1073 (O_1073,N_14994,N_14820);
nand UO_1074 (O_1074,N_14810,N_14913);
and UO_1075 (O_1075,N_14881,N_14901);
xnor UO_1076 (O_1076,N_14816,N_14905);
and UO_1077 (O_1077,N_14994,N_14831);
nor UO_1078 (O_1078,N_14992,N_14840);
or UO_1079 (O_1079,N_14909,N_14826);
or UO_1080 (O_1080,N_14804,N_14845);
or UO_1081 (O_1081,N_14920,N_14884);
nor UO_1082 (O_1082,N_14996,N_14953);
xor UO_1083 (O_1083,N_14880,N_14897);
nor UO_1084 (O_1084,N_14887,N_14974);
nand UO_1085 (O_1085,N_14812,N_14840);
nand UO_1086 (O_1086,N_14822,N_14806);
nor UO_1087 (O_1087,N_14857,N_14822);
nand UO_1088 (O_1088,N_14862,N_14840);
nand UO_1089 (O_1089,N_14893,N_14976);
nor UO_1090 (O_1090,N_14804,N_14995);
nand UO_1091 (O_1091,N_14825,N_14897);
nor UO_1092 (O_1092,N_14880,N_14932);
nor UO_1093 (O_1093,N_14984,N_14938);
or UO_1094 (O_1094,N_14941,N_14837);
xnor UO_1095 (O_1095,N_14970,N_14935);
and UO_1096 (O_1096,N_14830,N_14978);
nand UO_1097 (O_1097,N_14988,N_14886);
xnor UO_1098 (O_1098,N_14937,N_14850);
nor UO_1099 (O_1099,N_14883,N_14854);
and UO_1100 (O_1100,N_14867,N_14999);
or UO_1101 (O_1101,N_14842,N_14858);
nand UO_1102 (O_1102,N_14859,N_14896);
nor UO_1103 (O_1103,N_14962,N_14918);
nor UO_1104 (O_1104,N_14931,N_14811);
nand UO_1105 (O_1105,N_14904,N_14836);
or UO_1106 (O_1106,N_14954,N_14823);
nor UO_1107 (O_1107,N_14865,N_14914);
and UO_1108 (O_1108,N_14952,N_14847);
and UO_1109 (O_1109,N_14982,N_14823);
nor UO_1110 (O_1110,N_14900,N_14836);
or UO_1111 (O_1111,N_14850,N_14917);
nor UO_1112 (O_1112,N_14811,N_14911);
nand UO_1113 (O_1113,N_14958,N_14931);
and UO_1114 (O_1114,N_14844,N_14923);
and UO_1115 (O_1115,N_14999,N_14890);
and UO_1116 (O_1116,N_14997,N_14844);
nor UO_1117 (O_1117,N_14804,N_14924);
nor UO_1118 (O_1118,N_14831,N_14830);
xor UO_1119 (O_1119,N_14804,N_14963);
and UO_1120 (O_1120,N_14989,N_14976);
or UO_1121 (O_1121,N_14855,N_14834);
xnor UO_1122 (O_1122,N_14931,N_14996);
or UO_1123 (O_1123,N_14895,N_14806);
nand UO_1124 (O_1124,N_14807,N_14949);
nor UO_1125 (O_1125,N_14880,N_14813);
and UO_1126 (O_1126,N_14825,N_14973);
or UO_1127 (O_1127,N_14980,N_14989);
and UO_1128 (O_1128,N_14862,N_14992);
nand UO_1129 (O_1129,N_14961,N_14997);
nor UO_1130 (O_1130,N_14997,N_14895);
nor UO_1131 (O_1131,N_14918,N_14826);
or UO_1132 (O_1132,N_14954,N_14995);
nor UO_1133 (O_1133,N_14993,N_14963);
nand UO_1134 (O_1134,N_14856,N_14961);
nand UO_1135 (O_1135,N_14976,N_14865);
nor UO_1136 (O_1136,N_14875,N_14865);
and UO_1137 (O_1137,N_14873,N_14872);
nor UO_1138 (O_1138,N_14934,N_14913);
and UO_1139 (O_1139,N_14829,N_14854);
nor UO_1140 (O_1140,N_14815,N_14998);
or UO_1141 (O_1141,N_14913,N_14841);
and UO_1142 (O_1142,N_14930,N_14893);
nand UO_1143 (O_1143,N_14984,N_14847);
nor UO_1144 (O_1144,N_14866,N_14815);
nor UO_1145 (O_1145,N_14812,N_14822);
nand UO_1146 (O_1146,N_14867,N_14998);
nand UO_1147 (O_1147,N_14971,N_14805);
or UO_1148 (O_1148,N_14876,N_14815);
and UO_1149 (O_1149,N_14956,N_14818);
or UO_1150 (O_1150,N_14820,N_14816);
or UO_1151 (O_1151,N_14918,N_14924);
or UO_1152 (O_1152,N_14906,N_14974);
or UO_1153 (O_1153,N_14974,N_14869);
nand UO_1154 (O_1154,N_14823,N_14830);
or UO_1155 (O_1155,N_14821,N_14847);
nand UO_1156 (O_1156,N_14882,N_14934);
or UO_1157 (O_1157,N_14923,N_14921);
xor UO_1158 (O_1158,N_14800,N_14918);
and UO_1159 (O_1159,N_14989,N_14857);
or UO_1160 (O_1160,N_14877,N_14817);
nand UO_1161 (O_1161,N_14813,N_14852);
and UO_1162 (O_1162,N_14864,N_14831);
nor UO_1163 (O_1163,N_14963,N_14839);
or UO_1164 (O_1164,N_14961,N_14873);
or UO_1165 (O_1165,N_14911,N_14865);
nand UO_1166 (O_1166,N_14851,N_14883);
nor UO_1167 (O_1167,N_14892,N_14827);
xor UO_1168 (O_1168,N_14889,N_14998);
nor UO_1169 (O_1169,N_14969,N_14989);
xnor UO_1170 (O_1170,N_14929,N_14879);
nand UO_1171 (O_1171,N_14826,N_14948);
nand UO_1172 (O_1172,N_14949,N_14957);
and UO_1173 (O_1173,N_14971,N_14967);
and UO_1174 (O_1174,N_14918,N_14860);
nor UO_1175 (O_1175,N_14842,N_14896);
or UO_1176 (O_1176,N_14991,N_14919);
nand UO_1177 (O_1177,N_14820,N_14868);
nand UO_1178 (O_1178,N_14942,N_14822);
or UO_1179 (O_1179,N_14973,N_14855);
and UO_1180 (O_1180,N_14851,N_14840);
or UO_1181 (O_1181,N_14872,N_14942);
or UO_1182 (O_1182,N_14927,N_14986);
or UO_1183 (O_1183,N_14967,N_14958);
nand UO_1184 (O_1184,N_14861,N_14811);
nor UO_1185 (O_1185,N_14981,N_14803);
nand UO_1186 (O_1186,N_14946,N_14991);
xor UO_1187 (O_1187,N_14832,N_14919);
nor UO_1188 (O_1188,N_14890,N_14933);
or UO_1189 (O_1189,N_14817,N_14865);
or UO_1190 (O_1190,N_14834,N_14859);
nor UO_1191 (O_1191,N_14924,N_14991);
nor UO_1192 (O_1192,N_14877,N_14898);
and UO_1193 (O_1193,N_14839,N_14949);
nand UO_1194 (O_1194,N_14897,N_14903);
and UO_1195 (O_1195,N_14966,N_14919);
nand UO_1196 (O_1196,N_14842,N_14876);
nand UO_1197 (O_1197,N_14963,N_14979);
xor UO_1198 (O_1198,N_14992,N_14895);
or UO_1199 (O_1199,N_14932,N_14967);
nand UO_1200 (O_1200,N_14905,N_14834);
and UO_1201 (O_1201,N_14884,N_14960);
nor UO_1202 (O_1202,N_14954,N_14828);
or UO_1203 (O_1203,N_14889,N_14875);
or UO_1204 (O_1204,N_14909,N_14880);
or UO_1205 (O_1205,N_14802,N_14950);
xnor UO_1206 (O_1206,N_14930,N_14928);
nor UO_1207 (O_1207,N_14961,N_14805);
or UO_1208 (O_1208,N_14857,N_14897);
and UO_1209 (O_1209,N_14909,N_14872);
nand UO_1210 (O_1210,N_14843,N_14806);
or UO_1211 (O_1211,N_14824,N_14804);
and UO_1212 (O_1212,N_14976,N_14965);
nand UO_1213 (O_1213,N_14835,N_14950);
or UO_1214 (O_1214,N_14964,N_14933);
and UO_1215 (O_1215,N_14873,N_14890);
or UO_1216 (O_1216,N_14888,N_14821);
nor UO_1217 (O_1217,N_14869,N_14895);
and UO_1218 (O_1218,N_14988,N_14991);
or UO_1219 (O_1219,N_14850,N_14800);
and UO_1220 (O_1220,N_14962,N_14991);
nor UO_1221 (O_1221,N_14995,N_14873);
and UO_1222 (O_1222,N_14886,N_14816);
nor UO_1223 (O_1223,N_14862,N_14822);
or UO_1224 (O_1224,N_14847,N_14861);
and UO_1225 (O_1225,N_14943,N_14909);
and UO_1226 (O_1226,N_14800,N_14922);
nand UO_1227 (O_1227,N_14929,N_14954);
and UO_1228 (O_1228,N_14978,N_14853);
xnor UO_1229 (O_1229,N_14854,N_14925);
nand UO_1230 (O_1230,N_14860,N_14890);
xor UO_1231 (O_1231,N_14998,N_14923);
nand UO_1232 (O_1232,N_14993,N_14846);
nand UO_1233 (O_1233,N_14912,N_14842);
and UO_1234 (O_1234,N_14803,N_14864);
and UO_1235 (O_1235,N_14966,N_14999);
xor UO_1236 (O_1236,N_14831,N_14927);
nor UO_1237 (O_1237,N_14883,N_14951);
nand UO_1238 (O_1238,N_14985,N_14948);
and UO_1239 (O_1239,N_14838,N_14962);
or UO_1240 (O_1240,N_14937,N_14885);
and UO_1241 (O_1241,N_14917,N_14849);
nand UO_1242 (O_1242,N_14903,N_14896);
or UO_1243 (O_1243,N_14831,N_14983);
nor UO_1244 (O_1244,N_14852,N_14882);
or UO_1245 (O_1245,N_14904,N_14915);
or UO_1246 (O_1246,N_14853,N_14916);
nand UO_1247 (O_1247,N_14846,N_14826);
and UO_1248 (O_1248,N_14800,N_14892);
nand UO_1249 (O_1249,N_14976,N_14826);
nand UO_1250 (O_1250,N_14836,N_14871);
nor UO_1251 (O_1251,N_14903,N_14975);
nand UO_1252 (O_1252,N_14971,N_14918);
or UO_1253 (O_1253,N_14837,N_14992);
nor UO_1254 (O_1254,N_14965,N_14823);
or UO_1255 (O_1255,N_14931,N_14843);
and UO_1256 (O_1256,N_14815,N_14944);
nor UO_1257 (O_1257,N_14828,N_14860);
nor UO_1258 (O_1258,N_14815,N_14814);
or UO_1259 (O_1259,N_14806,N_14925);
nor UO_1260 (O_1260,N_14926,N_14938);
or UO_1261 (O_1261,N_14961,N_14849);
xor UO_1262 (O_1262,N_14982,N_14896);
nor UO_1263 (O_1263,N_14920,N_14881);
or UO_1264 (O_1264,N_14973,N_14841);
nand UO_1265 (O_1265,N_14881,N_14886);
and UO_1266 (O_1266,N_14854,N_14834);
or UO_1267 (O_1267,N_14937,N_14978);
and UO_1268 (O_1268,N_14898,N_14890);
or UO_1269 (O_1269,N_14961,N_14826);
nor UO_1270 (O_1270,N_14924,N_14942);
nand UO_1271 (O_1271,N_14883,N_14895);
xnor UO_1272 (O_1272,N_14984,N_14934);
nor UO_1273 (O_1273,N_14925,N_14860);
or UO_1274 (O_1274,N_14918,N_14941);
nand UO_1275 (O_1275,N_14939,N_14825);
nor UO_1276 (O_1276,N_14864,N_14965);
nor UO_1277 (O_1277,N_14917,N_14880);
or UO_1278 (O_1278,N_14983,N_14879);
nand UO_1279 (O_1279,N_14899,N_14811);
or UO_1280 (O_1280,N_14940,N_14876);
nand UO_1281 (O_1281,N_14834,N_14809);
nor UO_1282 (O_1282,N_14967,N_14816);
nand UO_1283 (O_1283,N_14919,N_14974);
nor UO_1284 (O_1284,N_14865,N_14902);
nor UO_1285 (O_1285,N_14962,N_14852);
nor UO_1286 (O_1286,N_14889,N_14950);
nand UO_1287 (O_1287,N_14869,N_14853);
and UO_1288 (O_1288,N_14981,N_14858);
nor UO_1289 (O_1289,N_14900,N_14892);
and UO_1290 (O_1290,N_14893,N_14984);
nor UO_1291 (O_1291,N_14988,N_14817);
nor UO_1292 (O_1292,N_14844,N_14909);
or UO_1293 (O_1293,N_14800,N_14831);
nand UO_1294 (O_1294,N_14884,N_14871);
and UO_1295 (O_1295,N_14831,N_14984);
or UO_1296 (O_1296,N_14951,N_14836);
nor UO_1297 (O_1297,N_14829,N_14928);
and UO_1298 (O_1298,N_14870,N_14894);
or UO_1299 (O_1299,N_14845,N_14889);
or UO_1300 (O_1300,N_14815,N_14922);
nand UO_1301 (O_1301,N_14813,N_14915);
nand UO_1302 (O_1302,N_14887,N_14914);
or UO_1303 (O_1303,N_14948,N_14983);
nand UO_1304 (O_1304,N_14979,N_14914);
or UO_1305 (O_1305,N_14969,N_14908);
and UO_1306 (O_1306,N_14860,N_14900);
and UO_1307 (O_1307,N_14879,N_14845);
nand UO_1308 (O_1308,N_14887,N_14844);
xnor UO_1309 (O_1309,N_14929,N_14848);
and UO_1310 (O_1310,N_14813,N_14961);
nand UO_1311 (O_1311,N_14996,N_14979);
or UO_1312 (O_1312,N_14982,N_14817);
and UO_1313 (O_1313,N_14898,N_14999);
and UO_1314 (O_1314,N_14951,N_14869);
and UO_1315 (O_1315,N_14939,N_14907);
and UO_1316 (O_1316,N_14987,N_14953);
and UO_1317 (O_1317,N_14869,N_14908);
nand UO_1318 (O_1318,N_14978,N_14802);
and UO_1319 (O_1319,N_14918,N_14950);
or UO_1320 (O_1320,N_14849,N_14969);
nand UO_1321 (O_1321,N_14929,N_14933);
nand UO_1322 (O_1322,N_14977,N_14902);
and UO_1323 (O_1323,N_14824,N_14855);
nand UO_1324 (O_1324,N_14999,N_14921);
or UO_1325 (O_1325,N_14893,N_14827);
nand UO_1326 (O_1326,N_14810,N_14832);
or UO_1327 (O_1327,N_14895,N_14924);
nor UO_1328 (O_1328,N_14903,N_14818);
nor UO_1329 (O_1329,N_14968,N_14946);
or UO_1330 (O_1330,N_14823,N_14811);
or UO_1331 (O_1331,N_14980,N_14800);
xnor UO_1332 (O_1332,N_14910,N_14917);
or UO_1333 (O_1333,N_14974,N_14858);
nor UO_1334 (O_1334,N_14837,N_14924);
and UO_1335 (O_1335,N_14812,N_14829);
nor UO_1336 (O_1336,N_14876,N_14968);
or UO_1337 (O_1337,N_14886,N_14896);
nor UO_1338 (O_1338,N_14854,N_14814);
and UO_1339 (O_1339,N_14856,N_14909);
nor UO_1340 (O_1340,N_14935,N_14983);
nor UO_1341 (O_1341,N_14952,N_14821);
and UO_1342 (O_1342,N_14826,N_14936);
or UO_1343 (O_1343,N_14912,N_14901);
or UO_1344 (O_1344,N_14886,N_14938);
nor UO_1345 (O_1345,N_14844,N_14966);
or UO_1346 (O_1346,N_14894,N_14983);
or UO_1347 (O_1347,N_14938,N_14941);
nor UO_1348 (O_1348,N_14854,N_14843);
and UO_1349 (O_1349,N_14926,N_14972);
and UO_1350 (O_1350,N_14951,N_14811);
nand UO_1351 (O_1351,N_14803,N_14904);
and UO_1352 (O_1352,N_14997,N_14829);
or UO_1353 (O_1353,N_14923,N_14859);
nor UO_1354 (O_1354,N_14861,N_14941);
or UO_1355 (O_1355,N_14937,N_14910);
or UO_1356 (O_1356,N_14937,N_14959);
nand UO_1357 (O_1357,N_14911,N_14831);
nand UO_1358 (O_1358,N_14838,N_14888);
xor UO_1359 (O_1359,N_14806,N_14897);
and UO_1360 (O_1360,N_14915,N_14845);
nor UO_1361 (O_1361,N_14809,N_14847);
nor UO_1362 (O_1362,N_14872,N_14928);
or UO_1363 (O_1363,N_14869,N_14956);
nand UO_1364 (O_1364,N_14918,N_14881);
and UO_1365 (O_1365,N_14858,N_14878);
nor UO_1366 (O_1366,N_14962,N_14931);
and UO_1367 (O_1367,N_14990,N_14850);
or UO_1368 (O_1368,N_14822,N_14867);
nor UO_1369 (O_1369,N_14813,N_14989);
nor UO_1370 (O_1370,N_14878,N_14850);
nor UO_1371 (O_1371,N_14909,N_14992);
or UO_1372 (O_1372,N_14924,N_14813);
or UO_1373 (O_1373,N_14802,N_14964);
nor UO_1374 (O_1374,N_14843,N_14988);
nand UO_1375 (O_1375,N_14835,N_14960);
or UO_1376 (O_1376,N_14939,N_14896);
nand UO_1377 (O_1377,N_14840,N_14876);
nand UO_1378 (O_1378,N_14830,N_14969);
or UO_1379 (O_1379,N_14879,N_14905);
and UO_1380 (O_1380,N_14989,N_14871);
and UO_1381 (O_1381,N_14867,N_14884);
or UO_1382 (O_1382,N_14816,N_14802);
and UO_1383 (O_1383,N_14968,N_14829);
nor UO_1384 (O_1384,N_14816,N_14835);
xnor UO_1385 (O_1385,N_14967,N_14830);
or UO_1386 (O_1386,N_14841,N_14804);
nor UO_1387 (O_1387,N_14931,N_14940);
nor UO_1388 (O_1388,N_14995,N_14833);
nand UO_1389 (O_1389,N_14887,N_14875);
nor UO_1390 (O_1390,N_14966,N_14826);
and UO_1391 (O_1391,N_14945,N_14811);
and UO_1392 (O_1392,N_14922,N_14842);
nand UO_1393 (O_1393,N_14924,N_14889);
nor UO_1394 (O_1394,N_14851,N_14967);
nand UO_1395 (O_1395,N_14894,N_14806);
and UO_1396 (O_1396,N_14913,N_14977);
xor UO_1397 (O_1397,N_14816,N_14819);
and UO_1398 (O_1398,N_14820,N_14876);
and UO_1399 (O_1399,N_14933,N_14824);
or UO_1400 (O_1400,N_14919,N_14880);
nor UO_1401 (O_1401,N_14849,N_14988);
or UO_1402 (O_1402,N_14880,N_14938);
nand UO_1403 (O_1403,N_14984,N_14946);
nand UO_1404 (O_1404,N_14996,N_14978);
nand UO_1405 (O_1405,N_14899,N_14960);
and UO_1406 (O_1406,N_14885,N_14964);
nand UO_1407 (O_1407,N_14986,N_14897);
nand UO_1408 (O_1408,N_14967,N_14907);
and UO_1409 (O_1409,N_14839,N_14951);
or UO_1410 (O_1410,N_14834,N_14959);
and UO_1411 (O_1411,N_14860,N_14937);
or UO_1412 (O_1412,N_14816,N_14869);
nor UO_1413 (O_1413,N_14895,N_14983);
and UO_1414 (O_1414,N_14822,N_14978);
nor UO_1415 (O_1415,N_14881,N_14897);
or UO_1416 (O_1416,N_14984,N_14803);
nor UO_1417 (O_1417,N_14825,N_14961);
nor UO_1418 (O_1418,N_14905,N_14805);
nand UO_1419 (O_1419,N_14812,N_14986);
or UO_1420 (O_1420,N_14967,N_14916);
nand UO_1421 (O_1421,N_14973,N_14817);
nor UO_1422 (O_1422,N_14833,N_14965);
nand UO_1423 (O_1423,N_14804,N_14860);
and UO_1424 (O_1424,N_14986,N_14874);
nor UO_1425 (O_1425,N_14966,N_14953);
nand UO_1426 (O_1426,N_14849,N_14944);
nand UO_1427 (O_1427,N_14997,N_14894);
and UO_1428 (O_1428,N_14842,N_14969);
and UO_1429 (O_1429,N_14954,N_14919);
nand UO_1430 (O_1430,N_14883,N_14902);
or UO_1431 (O_1431,N_14860,N_14859);
nand UO_1432 (O_1432,N_14810,N_14861);
nor UO_1433 (O_1433,N_14900,N_14954);
or UO_1434 (O_1434,N_14987,N_14867);
nand UO_1435 (O_1435,N_14969,N_14938);
xnor UO_1436 (O_1436,N_14976,N_14990);
nand UO_1437 (O_1437,N_14873,N_14970);
nor UO_1438 (O_1438,N_14981,N_14883);
nand UO_1439 (O_1439,N_14953,N_14976);
or UO_1440 (O_1440,N_14947,N_14890);
and UO_1441 (O_1441,N_14978,N_14890);
and UO_1442 (O_1442,N_14977,N_14983);
nor UO_1443 (O_1443,N_14899,N_14809);
nand UO_1444 (O_1444,N_14996,N_14999);
or UO_1445 (O_1445,N_14984,N_14911);
and UO_1446 (O_1446,N_14943,N_14989);
and UO_1447 (O_1447,N_14912,N_14802);
nor UO_1448 (O_1448,N_14920,N_14987);
and UO_1449 (O_1449,N_14803,N_14828);
nand UO_1450 (O_1450,N_14983,N_14809);
nor UO_1451 (O_1451,N_14857,N_14877);
or UO_1452 (O_1452,N_14996,N_14838);
nor UO_1453 (O_1453,N_14981,N_14825);
nor UO_1454 (O_1454,N_14957,N_14867);
nand UO_1455 (O_1455,N_14834,N_14845);
or UO_1456 (O_1456,N_14989,N_14842);
nor UO_1457 (O_1457,N_14970,N_14903);
and UO_1458 (O_1458,N_14819,N_14857);
or UO_1459 (O_1459,N_14943,N_14832);
and UO_1460 (O_1460,N_14804,N_14928);
nand UO_1461 (O_1461,N_14967,N_14857);
and UO_1462 (O_1462,N_14995,N_14956);
nor UO_1463 (O_1463,N_14860,N_14915);
nor UO_1464 (O_1464,N_14850,N_14918);
or UO_1465 (O_1465,N_14966,N_14994);
nand UO_1466 (O_1466,N_14904,N_14842);
or UO_1467 (O_1467,N_14962,N_14903);
nor UO_1468 (O_1468,N_14891,N_14814);
or UO_1469 (O_1469,N_14800,N_14887);
or UO_1470 (O_1470,N_14929,N_14877);
nand UO_1471 (O_1471,N_14961,N_14843);
nand UO_1472 (O_1472,N_14993,N_14879);
or UO_1473 (O_1473,N_14867,N_14918);
xnor UO_1474 (O_1474,N_14835,N_14965);
or UO_1475 (O_1475,N_14807,N_14849);
and UO_1476 (O_1476,N_14901,N_14958);
nor UO_1477 (O_1477,N_14813,N_14925);
and UO_1478 (O_1478,N_14816,N_14818);
nand UO_1479 (O_1479,N_14804,N_14869);
or UO_1480 (O_1480,N_14805,N_14987);
nand UO_1481 (O_1481,N_14947,N_14913);
nor UO_1482 (O_1482,N_14915,N_14986);
nand UO_1483 (O_1483,N_14932,N_14828);
nor UO_1484 (O_1484,N_14856,N_14874);
nand UO_1485 (O_1485,N_14818,N_14963);
xnor UO_1486 (O_1486,N_14818,N_14811);
nand UO_1487 (O_1487,N_14996,N_14895);
nor UO_1488 (O_1488,N_14908,N_14830);
or UO_1489 (O_1489,N_14943,N_14944);
or UO_1490 (O_1490,N_14818,N_14945);
nor UO_1491 (O_1491,N_14978,N_14931);
nor UO_1492 (O_1492,N_14882,N_14930);
nand UO_1493 (O_1493,N_14849,N_14908);
nand UO_1494 (O_1494,N_14916,N_14975);
and UO_1495 (O_1495,N_14834,N_14888);
nor UO_1496 (O_1496,N_14925,N_14991);
and UO_1497 (O_1497,N_14810,N_14887);
or UO_1498 (O_1498,N_14869,N_14831);
nor UO_1499 (O_1499,N_14843,N_14829);
or UO_1500 (O_1500,N_14910,N_14915);
and UO_1501 (O_1501,N_14991,N_14805);
or UO_1502 (O_1502,N_14938,N_14986);
nand UO_1503 (O_1503,N_14888,N_14815);
and UO_1504 (O_1504,N_14983,N_14807);
nor UO_1505 (O_1505,N_14927,N_14919);
nand UO_1506 (O_1506,N_14895,N_14901);
or UO_1507 (O_1507,N_14954,N_14815);
nand UO_1508 (O_1508,N_14901,N_14987);
nand UO_1509 (O_1509,N_14909,N_14875);
and UO_1510 (O_1510,N_14913,N_14921);
or UO_1511 (O_1511,N_14954,N_14822);
and UO_1512 (O_1512,N_14832,N_14865);
and UO_1513 (O_1513,N_14912,N_14885);
and UO_1514 (O_1514,N_14979,N_14841);
and UO_1515 (O_1515,N_14963,N_14902);
or UO_1516 (O_1516,N_14846,N_14938);
nor UO_1517 (O_1517,N_14800,N_14823);
and UO_1518 (O_1518,N_14971,N_14815);
or UO_1519 (O_1519,N_14951,N_14921);
nand UO_1520 (O_1520,N_14971,N_14980);
or UO_1521 (O_1521,N_14832,N_14987);
and UO_1522 (O_1522,N_14896,N_14902);
and UO_1523 (O_1523,N_14816,N_14832);
nand UO_1524 (O_1524,N_14836,N_14801);
nor UO_1525 (O_1525,N_14872,N_14908);
or UO_1526 (O_1526,N_14931,N_14941);
xor UO_1527 (O_1527,N_14868,N_14923);
nand UO_1528 (O_1528,N_14933,N_14950);
nor UO_1529 (O_1529,N_14848,N_14968);
xor UO_1530 (O_1530,N_14850,N_14975);
and UO_1531 (O_1531,N_14861,N_14880);
xnor UO_1532 (O_1532,N_14843,N_14982);
or UO_1533 (O_1533,N_14936,N_14854);
nor UO_1534 (O_1534,N_14946,N_14971);
nor UO_1535 (O_1535,N_14876,N_14837);
and UO_1536 (O_1536,N_14900,N_14857);
nand UO_1537 (O_1537,N_14944,N_14899);
or UO_1538 (O_1538,N_14947,N_14959);
and UO_1539 (O_1539,N_14884,N_14829);
or UO_1540 (O_1540,N_14986,N_14830);
nand UO_1541 (O_1541,N_14930,N_14806);
or UO_1542 (O_1542,N_14921,N_14920);
nand UO_1543 (O_1543,N_14814,N_14871);
xor UO_1544 (O_1544,N_14810,N_14997);
or UO_1545 (O_1545,N_14975,N_14886);
and UO_1546 (O_1546,N_14953,N_14897);
nand UO_1547 (O_1547,N_14805,N_14882);
and UO_1548 (O_1548,N_14903,N_14879);
or UO_1549 (O_1549,N_14811,N_14909);
and UO_1550 (O_1550,N_14836,N_14803);
nor UO_1551 (O_1551,N_14954,N_14813);
nand UO_1552 (O_1552,N_14816,N_14924);
nor UO_1553 (O_1553,N_14828,N_14941);
and UO_1554 (O_1554,N_14924,N_14969);
or UO_1555 (O_1555,N_14905,N_14821);
nor UO_1556 (O_1556,N_14813,N_14905);
and UO_1557 (O_1557,N_14970,N_14857);
and UO_1558 (O_1558,N_14843,N_14871);
nor UO_1559 (O_1559,N_14923,N_14962);
and UO_1560 (O_1560,N_14858,N_14822);
nand UO_1561 (O_1561,N_14899,N_14883);
and UO_1562 (O_1562,N_14969,N_14904);
nor UO_1563 (O_1563,N_14905,N_14911);
xnor UO_1564 (O_1564,N_14888,N_14876);
or UO_1565 (O_1565,N_14834,N_14998);
nor UO_1566 (O_1566,N_14877,N_14834);
nor UO_1567 (O_1567,N_14998,N_14966);
and UO_1568 (O_1568,N_14883,N_14938);
nor UO_1569 (O_1569,N_14897,N_14905);
xnor UO_1570 (O_1570,N_14911,N_14855);
xnor UO_1571 (O_1571,N_14910,N_14801);
and UO_1572 (O_1572,N_14973,N_14857);
xnor UO_1573 (O_1573,N_14850,N_14843);
and UO_1574 (O_1574,N_14990,N_14887);
nor UO_1575 (O_1575,N_14803,N_14821);
nand UO_1576 (O_1576,N_14891,N_14921);
nand UO_1577 (O_1577,N_14902,N_14858);
nor UO_1578 (O_1578,N_14820,N_14957);
nand UO_1579 (O_1579,N_14994,N_14818);
and UO_1580 (O_1580,N_14812,N_14987);
nand UO_1581 (O_1581,N_14812,N_14834);
nor UO_1582 (O_1582,N_14919,N_14848);
or UO_1583 (O_1583,N_14907,N_14918);
nor UO_1584 (O_1584,N_14930,N_14979);
xnor UO_1585 (O_1585,N_14950,N_14927);
nand UO_1586 (O_1586,N_14849,N_14974);
or UO_1587 (O_1587,N_14829,N_14963);
nand UO_1588 (O_1588,N_14985,N_14958);
and UO_1589 (O_1589,N_14892,N_14999);
or UO_1590 (O_1590,N_14970,N_14802);
and UO_1591 (O_1591,N_14820,N_14911);
xor UO_1592 (O_1592,N_14825,N_14849);
nand UO_1593 (O_1593,N_14801,N_14975);
or UO_1594 (O_1594,N_14895,N_14907);
nor UO_1595 (O_1595,N_14989,N_14818);
nand UO_1596 (O_1596,N_14838,N_14825);
and UO_1597 (O_1597,N_14936,N_14896);
nand UO_1598 (O_1598,N_14946,N_14955);
nor UO_1599 (O_1599,N_14890,N_14940);
xnor UO_1600 (O_1600,N_14903,N_14901);
nand UO_1601 (O_1601,N_14975,N_14860);
nand UO_1602 (O_1602,N_14935,N_14839);
xor UO_1603 (O_1603,N_14834,N_14979);
nand UO_1604 (O_1604,N_14955,N_14802);
or UO_1605 (O_1605,N_14953,N_14807);
nand UO_1606 (O_1606,N_14900,N_14815);
or UO_1607 (O_1607,N_14823,N_14927);
xnor UO_1608 (O_1608,N_14836,N_14974);
nand UO_1609 (O_1609,N_14976,N_14969);
nor UO_1610 (O_1610,N_14934,N_14932);
and UO_1611 (O_1611,N_14827,N_14901);
nor UO_1612 (O_1612,N_14894,N_14837);
or UO_1613 (O_1613,N_14937,N_14954);
nor UO_1614 (O_1614,N_14932,N_14860);
xnor UO_1615 (O_1615,N_14823,N_14876);
nand UO_1616 (O_1616,N_14971,N_14802);
nand UO_1617 (O_1617,N_14983,N_14808);
and UO_1618 (O_1618,N_14994,N_14884);
or UO_1619 (O_1619,N_14938,N_14832);
nand UO_1620 (O_1620,N_14946,N_14974);
nor UO_1621 (O_1621,N_14850,N_14954);
and UO_1622 (O_1622,N_14842,N_14810);
xnor UO_1623 (O_1623,N_14886,N_14923);
nor UO_1624 (O_1624,N_14879,N_14818);
nor UO_1625 (O_1625,N_14912,N_14991);
nor UO_1626 (O_1626,N_14882,N_14919);
nor UO_1627 (O_1627,N_14860,N_14959);
nor UO_1628 (O_1628,N_14949,N_14915);
or UO_1629 (O_1629,N_14925,N_14872);
xor UO_1630 (O_1630,N_14951,N_14961);
nand UO_1631 (O_1631,N_14855,N_14990);
nand UO_1632 (O_1632,N_14930,N_14859);
xor UO_1633 (O_1633,N_14927,N_14884);
nand UO_1634 (O_1634,N_14872,N_14854);
xor UO_1635 (O_1635,N_14802,N_14859);
nor UO_1636 (O_1636,N_14953,N_14999);
or UO_1637 (O_1637,N_14911,N_14963);
and UO_1638 (O_1638,N_14861,N_14802);
or UO_1639 (O_1639,N_14962,N_14987);
or UO_1640 (O_1640,N_14825,N_14917);
nand UO_1641 (O_1641,N_14903,N_14956);
and UO_1642 (O_1642,N_14907,N_14959);
or UO_1643 (O_1643,N_14849,N_14838);
nand UO_1644 (O_1644,N_14863,N_14858);
nand UO_1645 (O_1645,N_14908,N_14889);
and UO_1646 (O_1646,N_14822,N_14839);
nor UO_1647 (O_1647,N_14808,N_14916);
and UO_1648 (O_1648,N_14804,N_14984);
nand UO_1649 (O_1649,N_14999,N_14911);
nand UO_1650 (O_1650,N_14820,N_14888);
nand UO_1651 (O_1651,N_14987,N_14967);
or UO_1652 (O_1652,N_14934,N_14942);
xor UO_1653 (O_1653,N_14895,N_14982);
nand UO_1654 (O_1654,N_14941,N_14907);
nor UO_1655 (O_1655,N_14962,N_14976);
or UO_1656 (O_1656,N_14988,N_14828);
nand UO_1657 (O_1657,N_14951,N_14832);
nor UO_1658 (O_1658,N_14824,N_14895);
xnor UO_1659 (O_1659,N_14962,N_14830);
or UO_1660 (O_1660,N_14927,N_14939);
nand UO_1661 (O_1661,N_14928,N_14983);
nand UO_1662 (O_1662,N_14927,N_14926);
and UO_1663 (O_1663,N_14846,N_14898);
or UO_1664 (O_1664,N_14994,N_14856);
or UO_1665 (O_1665,N_14824,N_14920);
nand UO_1666 (O_1666,N_14942,N_14959);
xnor UO_1667 (O_1667,N_14969,N_14934);
nor UO_1668 (O_1668,N_14829,N_14946);
or UO_1669 (O_1669,N_14902,N_14909);
and UO_1670 (O_1670,N_14977,N_14930);
nor UO_1671 (O_1671,N_14836,N_14876);
nor UO_1672 (O_1672,N_14982,N_14987);
xor UO_1673 (O_1673,N_14986,N_14870);
nor UO_1674 (O_1674,N_14955,N_14860);
and UO_1675 (O_1675,N_14995,N_14802);
xnor UO_1676 (O_1676,N_14951,N_14899);
xnor UO_1677 (O_1677,N_14876,N_14905);
and UO_1678 (O_1678,N_14830,N_14959);
and UO_1679 (O_1679,N_14804,N_14975);
xnor UO_1680 (O_1680,N_14812,N_14835);
nor UO_1681 (O_1681,N_14978,N_14845);
nor UO_1682 (O_1682,N_14951,N_14833);
or UO_1683 (O_1683,N_14931,N_14874);
nor UO_1684 (O_1684,N_14957,N_14875);
and UO_1685 (O_1685,N_14974,N_14984);
or UO_1686 (O_1686,N_14817,N_14868);
or UO_1687 (O_1687,N_14817,N_14816);
or UO_1688 (O_1688,N_14998,N_14962);
xnor UO_1689 (O_1689,N_14823,N_14985);
nand UO_1690 (O_1690,N_14812,N_14910);
nor UO_1691 (O_1691,N_14932,N_14975);
nand UO_1692 (O_1692,N_14857,N_14868);
nor UO_1693 (O_1693,N_14871,N_14882);
or UO_1694 (O_1694,N_14879,N_14866);
or UO_1695 (O_1695,N_14892,N_14995);
nand UO_1696 (O_1696,N_14844,N_14847);
nor UO_1697 (O_1697,N_14937,N_14943);
nor UO_1698 (O_1698,N_14841,N_14985);
xnor UO_1699 (O_1699,N_14938,N_14873);
and UO_1700 (O_1700,N_14884,N_14995);
and UO_1701 (O_1701,N_14992,N_14905);
nand UO_1702 (O_1702,N_14800,N_14935);
nand UO_1703 (O_1703,N_14992,N_14897);
and UO_1704 (O_1704,N_14884,N_14973);
or UO_1705 (O_1705,N_14982,N_14898);
nand UO_1706 (O_1706,N_14966,N_14993);
nand UO_1707 (O_1707,N_14946,N_14864);
or UO_1708 (O_1708,N_14899,N_14920);
and UO_1709 (O_1709,N_14910,N_14904);
and UO_1710 (O_1710,N_14942,N_14897);
xor UO_1711 (O_1711,N_14982,N_14871);
nand UO_1712 (O_1712,N_14896,N_14951);
nand UO_1713 (O_1713,N_14906,N_14919);
nand UO_1714 (O_1714,N_14950,N_14887);
nand UO_1715 (O_1715,N_14911,N_14891);
nor UO_1716 (O_1716,N_14841,N_14811);
or UO_1717 (O_1717,N_14834,N_14872);
or UO_1718 (O_1718,N_14859,N_14850);
nor UO_1719 (O_1719,N_14953,N_14989);
or UO_1720 (O_1720,N_14877,N_14824);
or UO_1721 (O_1721,N_14876,N_14980);
xnor UO_1722 (O_1722,N_14937,N_14968);
or UO_1723 (O_1723,N_14805,N_14974);
nand UO_1724 (O_1724,N_14815,N_14861);
xnor UO_1725 (O_1725,N_14970,N_14860);
nor UO_1726 (O_1726,N_14843,N_14987);
nand UO_1727 (O_1727,N_14836,N_14927);
xor UO_1728 (O_1728,N_14934,N_14918);
or UO_1729 (O_1729,N_14844,N_14951);
nor UO_1730 (O_1730,N_14886,N_14981);
nand UO_1731 (O_1731,N_14853,N_14934);
or UO_1732 (O_1732,N_14837,N_14917);
nand UO_1733 (O_1733,N_14870,N_14914);
nand UO_1734 (O_1734,N_14925,N_14963);
nand UO_1735 (O_1735,N_14893,N_14927);
nand UO_1736 (O_1736,N_14885,N_14914);
and UO_1737 (O_1737,N_14924,N_14808);
or UO_1738 (O_1738,N_14984,N_14852);
or UO_1739 (O_1739,N_14971,N_14888);
and UO_1740 (O_1740,N_14849,N_14947);
and UO_1741 (O_1741,N_14886,N_14874);
and UO_1742 (O_1742,N_14903,N_14959);
and UO_1743 (O_1743,N_14932,N_14816);
nor UO_1744 (O_1744,N_14817,N_14987);
and UO_1745 (O_1745,N_14840,N_14961);
nand UO_1746 (O_1746,N_14959,N_14891);
nor UO_1747 (O_1747,N_14806,N_14805);
or UO_1748 (O_1748,N_14827,N_14845);
nor UO_1749 (O_1749,N_14844,N_14901);
nand UO_1750 (O_1750,N_14964,N_14849);
or UO_1751 (O_1751,N_14821,N_14900);
nor UO_1752 (O_1752,N_14925,N_14931);
or UO_1753 (O_1753,N_14827,N_14804);
or UO_1754 (O_1754,N_14896,N_14915);
xnor UO_1755 (O_1755,N_14803,N_14883);
or UO_1756 (O_1756,N_14986,N_14896);
and UO_1757 (O_1757,N_14937,N_14989);
nand UO_1758 (O_1758,N_14974,N_14864);
and UO_1759 (O_1759,N_14854,N_14868);
and UO_1760 (O_1760,N_14897,N_14854);
or UO_1761 (O_1761,N_14876,N_14814);
xor UO_1762 (O_1762,N_14812,N_14865);
nor UO_1763 (O_1763,N_14997,N_14935);
nand UO_1764 (O_1764,N_14913,N_14828);
nand UO_1765 (O_1765,N_14896,N_14885);
nand UO_1766 (O_1766,N_14957,N_14837);
nor UO_1767 (O_1767,N_14832,N_14959);
nand UO_1768 (O_1768,N_14927,N_14863);
nand UO_1769 (O_1769,N_14934,N_14829);
nor UO_1770 (O_1770,N_14922,N_14923);
and UO_1771 (O_1771,N_14833,N_14826);
nand UO_1772 (O_1772,N_14959,N_14809);
nor UO_1773 (O_1773,N_14851,N_14879);
and UO_1774 (O_1774,N_14917,N_14970);
nand UO_1775 (O_1775,N_14950,N_14823);
nand UO_1776 (O_1776,N_14876,N_14965);
nand UO_1777 (O_1777,N_14840,N_14880);
xor UO_1778 (O_1778,N_14990,N_14865);
xor UO_1779 (O_1779,N_14864,N_14887);
nor UO_1780 (O_1780,N_14910,N_14926);
nor UO_1781 (O_1781,N_14827,N_14990);
nand UO_1782 (O_1782,N_14858,N_14852);
and UO_1783 (O_1783,N_14900,N_14927);
xor UO_1784 (O_1784,N_14941,N_14970);
xnor UO_1785 (O_1785,N_14831,N_14949);
xnor UO_1786 (O_1786,N_14900,N_14801);
and UO_1787 (O_1787,N_14828,N_14914);
or UO_1788 (O_1788,N_14877,N_14810);
xor UO_1789 (O_1789,N_14892,N_14898);
nand UO_1790 (O_1790,N_14980,N_14907);
nand UO_1791 (O_1791,N_14819,N_14989);
nand UO_1792 (O_1792,N_14890,N_14960);
nand UO_1793 (O_1793,N_14855,N_14953);
nand UO_1794 (O_1794,N_14981,N_14921);
and UO_1795 (O_1795,N_14860,N_14866);
or UO_1796 (O_1796,N_14863,N_14907);
nor UO_1797 (O_1797,N_14870,N_14820);
and UO_1798 (O_1798,N_14981,N_14991);
nand UO_1799 (O_1799,N_14930,N_14834);
or UO_1800 (O_1800,N_14908,N_14960);
nand UO_1801 (O_1801,N_14949,N_14884);
nor UO_1802 (O_1802,N_14813,N_14977);
nand UO_1803 (O_1803,N_14912,N_14859);
or UO_1804 (O_1804,N_14864,N_14818);
nand UO_1805 (O_1805,N_14867,N_14885);
and UO_1806 (O_1806,N_14994,N_14834);
or UO_1807 (O_1807,N_14915,N_14980);
nor UO_1808 (O_1808,N_14844,N_14955);
nand UO_1809 (O_1809,N_14894,N_14988);
nor UO_1810 (O_1810,N_14804,N_14918);
nand UO_1811 (O_1811,N_14830,N_14936);
or UO_1812 (O_1812,N_14909,N_14822);
nand UO_1813 (O_1813,N_14958,N_14981);
nand UO_1814 (O_1814,N_14874,N_14863);
nor UO_1815 (O_1815,N_14872,N_14943);
or UO_1816 (O_1816,N_14853,N_14866);
or UO_1817 (O_1817,N_14843,N_14923);
and UO_1818 (O_1818,N_14945,N_14894);
or UO_1819 (O_1819,N_14940,N_14971);
nor UO_1820 (O_1820,N_14889,N_14882);
or UO_1821 (O_1821,N_14864,N_14890);
or UO_1822 (O_1822,N_14969,N_14836);
nand UO_1823 (O_1823,N_14857,N_14896);
nand UO_1824 (O_1824,N_14885,N_14902);
nor UO_1825 (O_1825,N_14800,N_14992);
and UO_1826 (O_1826,N_14904,N_14897);
nand UO_1827 (O_1827,N_14843,N_14840);
nor UO_1828 (O_1828,N_14968,N_14990);
xor UO_1829 (O_1829,N_14948,N_14990);
or UO_1830 (O_1830,N_14918,N_14894);
or UO_1831 (O_1831,N_14876,N_14976);
or UO_1832 (O_1832,N_14870,N_14910);
nor UO_1833 (O_1833,N_14823,N_14976);
nand UO_1834 (O_1834,N_14875,N_14921);
xor UO_1835 (O_1835,N_14873,N_14826);
and UO_1836 (O_1836,N_14964,N_14895);
nor UO_1837 (O_1837,N_14966,N_14914);
and UO_1838 (O_1838,N_14907,N_14998);
or UO_1839 (O_1839,N_14895,N_14915);
or UO_1840 (O_1840,N_14913,N_14967);
nor UO_1841 (O_1841,N_14871,N_14830);
nor UO_1842 (O_1842,N_14887,N_14926);
and UO_1843 (O_1843,N_14831,N_14974);
or UO_1844 (O_1844,N_14803,N_14931);
or UO_1845 (O_1845,N_14812,N_14897);
nand UO_1846 (O_1846,N_14846,N_14813);
nand UO_1847 (O_1847,N_14977,N_14907);
or UO_1848 (O_1848,N_14882,N_14825);
nand UO_1849 (O_1849,N_14990,N_14881);
nor UO_1850 (O_1850,N_14910,N_14802);
nand UO_1851 (O_1851,N_14837,N_14985);
xnor UO_1852 (O_1852,N_14842,N_14911);
and UO_1853 (O_1853,N_14977,N_14955);
nor UO_1854 (O_1854,N_14844,N_14996);
and UO_1855 (O_1855,N_14992,N_14857);
xor UO_1856 (O_1856,N_14924,N_14954);
nor UO_1857 (O_1857,N_14990,N_14943);
and UO_1858 (O_1858,N_14893,N_14879);
or UO_1859 (O_1859,N_14854,N_14875);
and UO_1860 (O_1860,N_14848,N_14902);
or UO_1861 (O_1861,N_14974,N_14935);
and UO_1862 (O_1862,N_14964,N_14963);
nor UO_1863 (O_1863,N_14934,N_14892);
nand UO_1864 (O_1864,N_14894,N_14867);
and UO_1865 (O_1865,N_14963,N_14879);
or UO_1866 (O_1866,N_14979,N_14865);
nor UO_1867 (O_1867,N_14942,N_14989);
and UO_1868 (O_1868,N_14875,N_14997);
xor UO_1869 (O_1869,N_14863,N_14908);
nor UO_1870 (O_1870,N_14966,N_14958);
nor UO_1871 (O_1871,N_14861,N_14965);
nand UO_1872 (O_1872,N_14897,N_14956);
nor UO_1873 (O_1873,N_14983,N_14964);
or UO_1874 (O_1874,N_14847,N_14942);
and UO_1875 (O_1875,N_14961,N_14803);
and UO_1876 (O_1876,N_14974,N_14995);
or UO_1877 (O_1877,N_14856,N_14867);
and UO_1878 (O_1878,N_14944,N_14854);
nand UO_1879 (O_1879,N_14913,N_14888);
xor UO_1880 (O_1880,N_14854,N_14899);
nor UO_1881 (O_1881,N_14908,N_14843);
or UO_1882 (O_1882,N_14918,N_14875);
nor UO_1883 (O_1883,N_14888,N_14965);
and UO_1884 (O_1884,N_14955,N_14978);
or UO_1885 (O_1885,N_14848,N_14844);
or UO_1886 (O_1886,N_14957,N_14868);
or UO_1887 (O_1887,N_14806,N_14931);
nand UO_1888 (O_1888,N_14903,N_14960);
or UO_1889 (O_1889,N_14983,N_14860);
xor UO_1890 (O_1890,N_14800,N_14966);
nor UO_1891 (O_1891,N_14830,N_14958);
or UO_1892 (O_1892,N_14893,N_14818);
and UO_1893 (O_1893,N_14953,N_14859);
and UO_1894 (O_1894,N_14922,N_14848);
or UO_1895 (O_1895,N_14853,N_14969);
nor UO_1896 (O_1896,N_14850,N_14870);
nand UO_1897 (O_1897,N_14996,N_14966);
and UO_1898 (O_1898,N_14822,N_14892);
or UO_1899 (O_1899,N_14913,N_14959);
and UO_1900 (O_1900,N_14891,N_14847);
nor UO_1901 (O_1901,N_14972,N_14918);
or UO_1902 (O_1902,N_14908,N_14910);
and UO_1903 (O_1903,N_14814,N_14958);
nand UO_1904 (O_1904,N_14802,N_14988);
and UO_1905 (O_1905,N_14994,N_14949);
nand UO_1906 (O_1906,N_14886,N_14969);
or UO_1907 (O_1907,N_14890,N_14904);
or UO_1908 (O_1908,N_14830,N_14824);
or UO_1909 (O_1909,N_14916,N_14954);
xnor UO_1910 (O_1910,N_14921,N_14812);
xnor UO_1911 (O_1911,N_14983,N_14986);
nand UO_1912 (O_1912,N_14869,N_14980);
and UO_1913 (O_1913,N_14889,N_14905);
nand UO_1914 (O_1914,N_14819,N_14838);
and UO_1915 (O_1915,N_14994,N_14900);
or UO_1916 (O_1916,N_14866,N_14988);
and UO_1917 (O_1917,N_14942,N_14846);
or UO_1918 (O_1918,N_14947,N_14817);
nand UO_1919 (O_1919,N_14933,N_14880);
nand UO_1920 (O_1920,N_14833,N_14919);
or UO_1921 (O_1921,N_14952,N_14956);
and UO_1922 (O_1922,N_14889,N_14841);
xor UO_1923 (O_1923,N_14988,N_14937);
or UO_1924 (O_1924,N_14811,N_14849);
nor UO_1925 (O_1925,N_14968,N_14923);
nor UO_1926 (O_1926,N_14942,N_14828);
and UO_1927 (O_1927,N_14893,N_14858);
nor UO_1928 (O_1928,N_14986,N_14813);
and UO_1929 (O_1929,N_14958,N_14951);
xnor UO_1930 (O_1930,N_14986,N_14819);
nor UO_1931 (O_1931,N_14881,N_14844);
and UO_1932 (O_1932,N_14887,N_14824);
or UO_1933 (O_1933,N_14967,N_14871);
nor UO_1934 (O_1934,N_14830,N_14878);
xor UO_1935 (O_1935,N_14806,N_14896);
nor UO_1936 (O_1936,N_14996,N_14862);
nand UO_1937 (O_1937,N_14968,N_14992);
or UO_1938 (O_1938,N_14825,N_14861);
or UO_1939 (O_1939,N_14804,N_14894);
nor UO_1940 (O_1940,N_14887,N_14848);
nor UO_1941 (O_1941,N_14830,N_14968);
or UO_1942 (O_1942,N_14936,N_14843);
and UO_1943 (O_1943,N_14835,N_14946);
or UO_1944 (O_1944,N_14942,N_14932);
nand UO_1945 (O_1945,N_14982,N_14966);
and UO_1946 (O_1946,N_14805,N_14836);
nor UO_1947 (O_1947,N_14959,N_14905);
nand UO_1948 (O_1948,N_14865,N_14951);
nor UO_1949 (O_1949,N_14962,N_14876);
or UO_1950 (O_1950,N_14800,N_14803);
or UO_1951 (O_1951,N_14954,N_14835);
nor UO_1952 (O_1952,N_14947,N_14975);
nand UO_1953 (O_1953,N_14998,N_14859);
nand UO_1954 (O_1954,N_14969,N_14819);
or UO_1955 (O_1955,N_14838,N_14801);
nor UO_1956 (O_1956,N_14991,N_14921);
or UO_1957 (O_1957,N_14841,N_14935);
nand UO_1958 (O_1958,N_14892,N_14924);
nor UO_1959 (O_1959,N_14909,N_14953);
nand UO_1960 (O_1960,N_14967,N_14841);
nand UO_1961 (O_1961,N_14822,N_14835);
and UO_1962 (O_1962,N_14900,N_14883);
and UO_1963 (O_1963,N_14923,N_14856);
or UO_1964 (O_1964,N_14920,N_14873);
nand UO_1965 (O_1965,N_14929,N_14876);
and UO_1966 (O_1966,N_14903,N_14902);
xor UO_1967 (O_1967,N_14890,N_14903);
and UO_1968 (O_1968,N_14886,N_14830);
or UO_1969 (O_1969,N_14804,N_14934);
nand UO_1970 (O_1970,N_14846,N_14841);
nor UO_1971 (O_1971,N_14800,N_14970);
or UO_1972 (O_1972,N_14881,N_14900);
xnor UO_1973 (O_1973,N_14905,N_14921);
xnor UO_1974 (O_1974,N_14912,N_14882);
or UO_1975 (O_1975,N_14995,N_14975);
nor UO_1976 (O_1976,N_14981,N_14856);
nand UO_1977 (O_1977,N_14992,N_14973);
and UO_1978 (O_1978,N_14932,N_14999);
nor UO_1979 (O_1979,N_14957,N_14884);
nand UO_1980 (O_1980,N_14991,N_14976);
nor UO_1981 (O_1981,N_14880,N_14803);
or UO_1982 (O_1982,N_14871,N_14951);
and UO_1983 (O_1983,N_14883,N_14898);
nand UO_1984 (O_1984,N_14848,N_14889);
nor UO_1985 (O_1985,N_14925,N_14933);
or UO_1986 (O_1986,N_14822,N_14903);
nor UO_1987 (O_1987,N_14875,N_14943);
or UO_1988 (O_1988,N_14956,N_14871);
nand UO_1989 (O_1989,N_14993,N_14873);
nand UO_1990 (O_1990,N_14957,N_14983);
or UO_1991 (O_1991,N_14863,N_14964);
and UO_1992 (O_1992,N_14814,N_14949);
or UO_1993 (O_1993,N_14856,N_14883);
nand UO_1994 (O_1994,N_14892,N_14973);
nand UO_1995 (O_1995,N_14996,N_14914);
nand UO_1996 (O_1996,N_14953,N_14994);
xor UO_1997 (O_1997,N_14849,N_14935);
nor UO_1998 (O_1998,N_14975,N_14870);
nor UO_1999 (O_1999,N_14831,N_14816);
endmodule