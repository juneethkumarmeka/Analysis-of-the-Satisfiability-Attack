module basic_3000_30000_3500_30_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nor U0 (N_0,In_1960,In_707);
nor U1 (N_1,In_2465,In_964);
xor U2 (N_2,In_2632,In_242);
or U3 (N_3,In_2319,In_673);
and U4 (N_4,In_2005,In_2886);
nor U5 (N_5,In_2111,In_2671);
nor U6 (N_6,In_1111,In_2483);
or U7 (N_7,In_2722,In_920);
nor U8 (N_8,In_762,In_1181);
or U9 (N_9,In_80,In_869);
or U10 (N_10,In_825,In_2244);
nand U11 (N_11,In_2265,In_957);
nor U12 (N_12,In_314,In_803);
nor U13 (N_13,In_922,In_1120);
xor U14 (N_14,In_1085,In_2270);
and U15 (N_15,In_1571,In_206);
xnor U16 (N_16,In_1376,In_2078);
xnor U17 (N_17,In_1909,In_1456);
nand U18 (N_18,In_1790,In_230);
or U19 (N_19,In_172,In_749);
nor U20 (N_20,In_1044,In_2582);
and U21 (N_21,In_2906,In_226);
nand U22 (N_22,In_1440,In_2364);
and U23 (N_23,In_1795,In_822);
xor U24 (N_24,In_567,In_321);
nand U25 (N_25,In_1600,In_1706);
and U26 (N_26,In_1236,In_175);
nor U27 (N_27,In_45,In_1404);
or U28 (N_28,In_743,In_1531);
nor U29 (N_29,In_2378,In_910);
nand U30 (N_30,In_335,In_1483);
nor U31 (N_31,In_1895,In_2994);
xnor U32 (N_32,In_682,In_287);
and U33 (N_33,In_2362,In_1294);
and U34 (N_34,In_633,In_1827);
nand U35 (N_35,In_1653,In_245);
nor U36 (N_36,In_561,In_1919);
xnor U37 (N_37,In_2814,In_1175);
and U38 (N_38,In_831,In_2278);
or U39 (N_39,In_902,In_1857);
nand U40 (N_40,In_595,In_1921);
nor U41 (N_41,In_110,In_979);
xnor U42 (N_42,In_1545,In_1247);
xor U43 (N_43,In_446,In_1133);
and U44 (N_44,In_2074,In_804);
or U45 (N_45,In_2822,In_50);
xnor U46 (N_46,In_1353,In_860);
and U47 (N_47,In_2885,In_2639);
nor U48 (N_48,In_1580,In_2797);
or U49 (N_49,In_2589,In_480);
xor U50 (N_50,In_2602,In_153);
nor U51 (N_51,In_334,In_2531);
or U52 (N_52,In_2854,In_481);
and U53 (N_53,In_2916,In_1265);
and U54 (N_54,In_1289,In_438);
nand U55 (N_55,In_987,In_1386);
and U56 (N_56,In_1500,In_165);
xnor U57 (N_57,In_2039,In_2380);
nor U58 (N_58,In_2734,In_2291);
and U59 (N_59,In_366,In_2143);
xor U60 (N_60,In_64,In_2847);
or U61 (N_61,In_969,In_2201);
xor U62 (N_62,In_346,In_182);
xor U63 (N_63,In_476,In_1949);
nand U64 (N_64,In_662,In_85);
or U65 (N_65,In_520,In_1620);
nand U66 (N_66,In_1388,In_968);
or U67 (N_67,In_1499,In_2293);
and U68 (N_68,In_1613,In_847);
nand U69 (N_69,In_1665,In_2764);
xor U70 (N_70,In_83,In_247);
or U71 (N_71,In_1764,In_2177);
nor U72 (N_72,In_1801,In_1532);
nor U73 (N_73,In_477,In_1806);
and U74 (N_74,In_2209,In_871);
nand U75 (N_75,In_1660,In_621);
nor U76 (N_76,In_2899,In_1402);
xnor U77 (N_77,In_1584,In_255);
nor U78 (N_78,In_529,In_2996);
nor U79 (N_79,In_781,In_48);
xnor U80 (N_80,In_888,In_1437);
nand U81 (N_81,In_38,In_2644);
and U82 (N_82,In_833,In_2837);
nand U83 (N_83,In_1115,In_2840);
nand U84 (N_84,In_2423,In_2988);
xor U85 (N_85,In_1064,In_722);
xnor U86 (N_86,In_2215,In_311);
xor U87 (N_87,In_1639,In_2615);
nand U88 (N_88,In_1868,In_756);
nor U89 (N_89,In_2190,In_1113);
xor U90 (N_90,In_700,In_1497);
nor U91 (N_91,In_1479,In_292);
nand U92 (N_92,In_2732,In_2684);
xnor U93 (N_93,In_1931,In_194);
nand U94 (N_94,In_0,In_2943);
or U95 (N_95,In_302,In_889);
nand U96 (N_96,In_2813,In_2607);
xnor U97 (N_97,In_768,In_2875);
nor U98 (N_98,In_148,In_386);
nand U99 (N_99,In_53,In_445);
xor U100 (N_100,In_179,In_1271);
xor U101 (N_101,In_1775,In_609);
xor U102 (N_102,In_1876,In_2281);
or U103 (N_103,In_2989,In_1991);
or U104 (N_104,In_1235,In_1715);
nor U105 (N_105,In_2972,In_1918);
nand U106 (N_106,In_128,In_101);
nor U107 (N_107,In_1306,In_272);
and U108 (N_108,In_2805,In_909);
and U109 (N_109,In_991,In_1615);
nor U110 (N_110,In_1482,In_1618);
nor U111 (N_111,In_2577,In_1155);
nor U112 (N_112,In_2913,In_2451);
xor U113 (N_113,In_1952,In_1209);
and U114 (N_114,In_2772,In_1623);
nand U115 (N_115,In_2739,In_2975);
or U116 (N_116,In_2486,In_170);
nand U117 (N_117,In_1215,In_1834);
nor U118 (N_118,In_2012,In_1872);
and U119 (N_119,In_916,In_21);
xnor U120 (N_120,In_903,In_2651);
xnor U121 (N_121,In_687,In_1858);
or U122 (N_122,In_1776,In_1561);
and U123 (N_123,In_345,In_2882);
nand U124 (N_124,In_924,In_706);
and U125 (N_125,In_2763,In_623);
xor U126 (N_126,In_2250,In_1896);
and U127 (N_127,In_2321,In_2016);
nor U128 (N_128,In_2112,In_1645);
and U129 (N_129,In_350,In_2510);
nand U130 (N_130,In_695,In_1212);
xnor U131 (N_131,In_2502,In_1826);
xor U132 (N_132,In_2981,In_378);
nand U133 (N_133,In_2402,In_1956);
xnor U134 (N_134,In_197,In_130);
and U135 (N_135,In_1824,In_1039);
xnor U136 (N_136,In_2650,In_2898);
nand U137 (N_137,In_1264,In_1902);
nor U138 (N_138,In_881,In_2371);
nor U139 (N_139,In_241,In_1225);
xor U140 (N_140,In_2939,In_2528);
or U141 (N_141,In_995,In_2731);
nand U142 (N_142,In_2770,In_2817);
or U143 (N_143,In_2273,In_138);
nand U144 (N_144,In_1446,In_2450);
or U145 (N_145,In_2153,In_2300);
and U146 (N_146,In_407,In_2663);
nor U147 (N_147,In_1784,In_2280);
nand U148 (N_148,In_1309,In_2066);
nor U149 (N_149,In_2211,In_519);
xor U150 (N_150,In_1177,In_1537);
and U151 (N_151,In_1380,In_1298);
xnor U152 (N_152,In_405,In_629);
or U153 (N_153,In_689,In_2150);
or U154 (N_154,In_2833,In_901);
nor U155 (N_155,In_329,In_631);
nor U156 (N_156,In_2944,In_2193);
nor U157 (N_157,In_872,In_598);
or U158 (N_158,In_843,In_1903);
or U159 (N_159,In_1518,In_2263);
and U160 (N_160,In_2735,In_2277);
or U161 (N_161,In_1074,In_167);
or U162 (N_162,In_611,In_389);
nand U163 (N_163,In_1760,In_792);
nand U164 (N_164,In_2396,In_2079);
xor U165 (N_165,In_1159,In_2747);
or U166 (N_166,In_813,In_1677);
nand U167 (N_167,In_2969,In_1278);
xnor U168 (N_168,In_2477,In_2010);
nor U169 (N_169,In_12,In_2626);
nand U170 (N_170,In_1932,In_625);
nand U171 (N_171,In_2680,In_1578);
nand U172 (N_172,In_2141,In_739);
xor U173 (N_173,In_2545,In_258);
nor U174 (N_174,In_2264,In_271);
or U175 (N_175,In_1805,In_2745);
nor U176 (N_176,In_887,In_2068);
nor U177 (N_177,In_2285,In_1812);
xor U178 (N_178,In_712,In_2120);
xor U179 (N_179,In_1375,In_2606);
or U180 (N_180,In_720,In_267);
nand U181 (N_181,In_2771,In_1714);
or U182 (N_182,In_2258,In_2021);
xnor U183 (N_183,In_2977,In_1988);
xor U184 (N_184,In_1308,In_2260);
nand U185 (N_185,In_1414,In_2729);
or U186 (N_186,In_2821,In_1399);
nor U187 (N_187,In_261,In_2248);
and U188 (N_188,In_2432,In_1652);
xor U189 (N_189,In_2816,In_1658);
or U190 (N_190,In_2839,In_2521);
nand U191 (N_191,In_440,In_2419);
nor U192 (N_192,In_1527,In_1598);
xnor U193 (N_193,In_677,In_933);
or U194 (N_194,In_1444,In_2634);
and U195 (N_195,In_2155,In_2983);
nor U196 (N_196,In_2812,In_2748);
and U197 (N_197,In_1293,In_94);
or U198 (N_198,In_355,In_2304);
or U199 (N_199,In_448,In_1324);
nand U200 (N_200,In_1110,In_1643);
and U201 (N_201,In_2147,In_2914);
nor U202 (N_202,In_671,In_2896);
and U203 (N_203,In_1281,In_826);
nand U204 (N_204,In_1152,In_502);
nand U205 (N_205,In_1505,In_744);
nor U206 (N_206,In_528,In_1621);
nor U207 (N_207,In_2004,In_2517);
xor U208 (N_208,In_1705,In_2256);
nor U209 (N_209,In_5,In_562);
and U210 (N_210,In_542,In_2391);
and U211 (N_211,In_1441,In_681);
xnor U212 (N_212,In_1053,In_2974);
nor U213 (N_213,In_1086,In_1469);
nor U214 (N_214,In_760,In_602);
xor U215 (N_215,In_1761,In_316);
nor U216 (N_216,In_2455,In_1741);
nand U217 (N_217,In_1649,In_391);
nor U218 (N_218,In_2071,In_1369);
xnor U219 (N_219,In_435,In_118);
or U220 (N_220,In_2668,In_473);
nor U221 (N_221,In_1690,In_1245);
or U222 (N_222,In_2709,In_1205);
nand U223 (N_223,In_61,In_2593);
and U224 (N_224,In_2538,In_2493);
xor U225 (N_225,In_1214,In_2034);
nor U226 (N_226,In_1725,In_2340);
xor U227 (N_227,In_2296,In_1165);
or U228 (N_228,In_1738,In_1641);
or U229 (N_229,In_766,In_2229);
or U230 (N_230,In_2730,In_2931);
or U231 (N_231,In_1221,In_790);
or U232 (N_232,In_2469,In_2773);
nand U233 (N_233,In_158,In_2238);
nor U234 (N_234,In_2951,In_1562);
xor U235 (N_235,In_2056,In_1077);
and U236 (N_236,In_1171,In_2154);
or U237 (N_237,In_593,In_451);
and U238 (N_238,In_147,In_1233);
nor U239 (N_239,In_2165,In_533);
and U240 (N_240,In_758,In_754);
and U241 (N_241,In_317,In_2971);
and U242 (N_242,In_2113,In_1471);
or U243 (N_243,In_1395,In_1928);
nand U244 (N_244,In_734,In_151);
nand U245 (N_245,In_2893,In_1299);
nand U246 (N_246,In_1357,In_775);
xnor U247 (N_247,In_2716,In_256);
xor U248 (N_248,In_1758,In_1130);
xor U249 (N_249,In_646,In_1279);
and U250 (N_250,In_2923,In_2098);
or U251 (N_251,In_390,In_372);
xnor U252 (N_252,In_667,In_2343);
nand U253 (N_253,In_127,In_1914);
nor U254 (N_254,In_235,In_2576);
xor U255 (N_255,In_1145,In_2261);
and U256 (N_256,In_263,In_437);
and U257 (N_257,In_87,In_469);
nor U258 (N_258,In_2895,In_210);
and U259 (N_259,In_1009,In_35);
and U260 (N_260,In_534,In_2213);
and U261 (N_261,In_193,In_458);
xnor U262 (N_262,In_1657,In_1682);
and U263 (N_263,In_2578,In_2308);
xor U264 (N_264,In_369,In_1144);
nand U265 (N_265,In_1798,In_2503);
or U266 (N_266,In_726,In_1157);
nand U267 (N_267,In_2504,In_2834);
nand U268 (N_268,In_717,In_1119);
and U269 (N_269,In_844,In_2013);
nand U270 (N_270,In_1457,In_1884);
nand U271 (N_271,In_2443,In_1109);
nor U272 (N_272,In_1892,In_2214);
or U273 (N_273,In_2656,In_1701);
nand U274 (N_274,In_731,In_2746);
or U275 (N_275,In_925,In_1929);
nor U276 (N_276,In_2637,In_891);
nor U277 (N_277,In_615,In_763);
nor U278 (N_278,In_1581,In_377);
and U279 (N_279,In_636,In_966);
nand U280 (N_280,In_2591,In_1439);
xor U281 (N_281,In_363,In_99);
nand U282 (N_282,In_159,In_2888);
or U283 (N_283,In_794,In_2126);
xor U284 (N_284,In_718,In_2274);
xor U285 (N_285,In_1977,In_2524);
nor U286 (N_286,In_212,In_97);
xor U287 (N_287,In_2024,In_432);
and U288 (N_288,In_475,In_140);
nor U289 (N_289,In_1739,In_1953);
and U290 (N_290,In_2791,In_293);
and U291 (N_291,In_1765,In_2176);
xor U292 (N_292,In_1727,In_1670);
or U293 (N_293,In_1153,In_2184);
or U294 (N_294,In_382,In_1049);
xor U295 (N_295,In_1882,In_1382);
nand U296 (N_296,In_806,In_1925);
and U297 (N_297,In_1924,In_1023);
or U298 (N_298,In_2043,In_1847);
and U299 (N_299,In_37,In_2017);
nor U300 (N_300,In_639,In_2767);
and U301 (N_301,In_2090,In_156);
nand U302 (N_302,In_2870,In_1276);
nand U303 (N_303,In_632,In_1755);
or U304 (N_304,In_74,In_526);
or U305 (N_305,In_285,In_1092);
nand U306 (N_306,In_2614,In_2623);
xnor U307 (N_307,In_1129,In_2349);
nand U308 (N_308,In_2221,In_985);
or U309 (N_309,In_1204,In_1344);
or U310 (N_310,In_367,In_2492);
and U311 (N_311,In_142,In_234);
and U312 (N_312,In_2353,In_977);
xnor U313 (N_313,In_2733,In_2064);
nand U314 (N_314,In_341,In_630);
or U315 (N_315,In_2720,In_2581);
xnor U316 (N_316,In_2041,In_333);
xnor U317 (N_317,In_1038,In_88);
nor U318 (N_318,In_2920,In_2332);
xor U319 (N_319,In_1788,In_2356);
nand U320 (N_320,In_586,In_1253);
nor U321 (N_321,In_55,In_205);
nor U322 (N_322,In_2104,In_414);
or U323 (N_323,In_1073,In_2782);
or U324 (N_324,In_296,In_2358);
and U325 (N_325,In_2890,In_155);
nand U326 (N_326,In_1061,In_647);
nand U327 (N_327,In_2092,In_1651);
and U328 (N_328,In_1223,In_954);
or U329 (N_329,In_2014,In_2131);
nor U330 (N_330,In_2219,In_2123);
nand U331 (N_331,In_2796,In_297);
nand U332 (N_332,In_1771,In_149);
xnor U333 (N_333,In_536,In_2516);
or U334 (N_334,In_552,In_2310);
or U335 (N_335,In_1272,In_820);
or U336 (N_336,In_2490,In_782);
xor U337 (N_337,In_2506,In_1906);
nand U338 (N_338,In_1029,In_2670);
or U339 (N_339,In_26,In_2233);
and U340 (N_340,In_2167,In_2156);
nand U341 (N_341,In_1314,In_2438);
xor U342 (N_342,In_1975,In_2509);
and U343 (N_343,In_1096,In_430);
nand U344 (N_344,In_2231,In_39);
xor U345 (N_345,In_1604,In_220);
nand U346 (N_346,In_436,In_1605);
xnor U347 (N_347,In_1057,In_1787);
and U348 (N_348,In_15,In_324);
nand U349 (N_349,In_1548,In_523);
nand U350 (N_350,In_679,In_343);
nand U351 (N_351,In_859,In_578);
or U352 (N_352,In_1890,In_1521);
nor U353 (N_353,In_1268,In_2006);
nand U354 (N_354,In_2871,In_1180);
or U355 (N_355,In_2379,In_340);
or U356 (N_356,In_1808,In_1090);
or U357 (N_357,In_1331,In_347);
or U358 (N_358,In_2072,In_2845);
and U359 (N_359,In_264,In_81);
and U360 (N_360,In_1297,In_1939);
and U361 (N_361,In_1712,In_2125);
nand U362 (N_362,In_651,In_119);
nor U363 (N_363,In_810,In_2393);
or U364 (N_364,In_1249,In_455);
nand U365 (N_365,In_2413,In_1391);
nand U366 (N_366,In_2317,In_2178);
nor U367 (N_367,In_1724,In_2355);
and U368 (N_368,In_2462,In_2312);
nor U369 (N_369,In_1546,In_236);
or U370 (N_370,In_8,In_184);
xnor U371 (N_371,In_482,In_1782);
or U372 (N_372,In_248,In_716);
nor U373 (N_373,In_1286,In_1523);
xor U374 (N_374,In_1478,In_1128);
nor U375 (N_375,In_2338,In_2133);
or U376 (N_376,In_2376,In_1789);
nor U377 (N_377,In_2491,In_307);
nand U378 (N_378,In_2030,In_1859);
and U379 (N_379,In_1709,In_2370);
nor U380 (N_380,In_2548,In_2991);
or U381 (N_381,In_305,In_1003);
nor U382 (N_382,In_2117,In_114);
xor U383 (N_383,In_1080,In_2927);
nand U384 (N_384,In_976,In_1586);
xor U385 (N_385,In_2019,In_928);
and U386 (N_386,In_1200,In_898);
xor U387 (N_387,In_2086,In_1908);
and U388 (N_388,In_2987,In_67);
nor U389 (N_389,In_1594,In_1726);
nor U390 (N_390,In_2526,In_2853);
and U391 (N_391,In_2683,In_2048);
nand U392 (N_392,In_885,In_51);
nand U393 (N_393,In_2653,In_2533);
and U394 (N_394,In_2753,In_6);
or U395 (N_395,In_215,In_2254);
nand U396 (N_396,In_753,In_2067);
xor U397 (N_397,In_2811,In_488);
or U398 (N_398,In_2130,In_524);
and U399 (N_399,In_2962,In_2103);
nor U400 (N_400,In_2032,In_1802);
xor U401 (N_401,In_259,In_1517);
xor U402 (N_402,In_698,In_2959);
and U403 (N_403,In_522,In_2554);
nor U404 (N_404,In_1560,In_972);
xnor U405 (N_405,In_2011,In_76);
nor U406 (N_406,In_664,In_2046);
or U407 (N_407,In_1487,In_789);
nand U408 (N_408,In_589,In_2081);
xor U409 (N_409,In_322,In_2286);
and U410 (N_410,In_597,In_2170);
or U411 (N_411,In_678,In_942);
or U412 (N_412,In_2808,In_905);
and U413 (N_413,In_2679,In_1210);
nand U414 (N_414,In_2205,In_498);
and U415 (N_415,In_1713,In_1224);
nand U416 (N_416,In_616,In_2879);
nor U417 (N_417,In_456,In_802);
and U418 (N_418,In_486,In_2793);
nand U419 (N_419,In_1550,In_2210);
or U420 (N_420,In_1504,In_463);
xnor U421 (N_421,In_1352,In_2894);
or U422 (N_422,In_1032,In_2995);
xnor U423 (N_423,In_431,In_897);
or U424 (N_424,In_644,In_2535);
and U425 (N_425,In_1316,In_1099);
and U426 (N_426,In_2873,In_2139);
nand U427 (N_427,In_709,In_1759);
and U428 (N_428,In_1830,In_1365);
and U429 (N_429,In_2693,In_2999);
and U430 (N_430,In_1252,In_1442);
nand U431 (N_431,In_2189,In_2571);
and U432 (N_432,In_610,In_1492);
xnor U433 (N_433,In_2194,In_801);
or U434 (N_434,In_1480,In_1511);
nor U435 (N_435,In_2829,In_2963);
nand U436 (N_436,In_332,In_69);
nand U437 (N_437,In_2558,In_1933);
and U438 (N_438,In_2059,In_850);
nor U439 (N_439,In_2351,In_1415);
nand U440 (N_440,In_2512,In_166);
and U441 (N_441,In_1364,In_2889);
nand U442 (N_442,In_1283,In_239);
nand U443 (N_443,In_2106,In_2587);
xor U444 (N_444,In_1559,In_2915);
xor U445 (N_445,In_1869,In_1410);
nor U446 (N_446,In_997,In_2698);
nand U447 (N_447,In_2386,In_331);
or U448 (N_448,In_1476,In_2108);
and U449 (N_449,In_2287,In_361);
nor U450 (N_450,In_2941,In_113);
nand U451 (N_451,In_2819,In_2594);
xnor U452 (N_452,In_2444,In_656);
nor U453 (N_453,In_2118,In_2279);
nor U454 (N_454,In_1799,In_1257);
and U455 (N_455,In_2099,In_946);
nand U456 (N_456,In_32,In_1100);
xor U457 (N_457,In_1676,In_1856);
nor U458 (N_458,In_66,In_2776);
and U459 (N_459,In_2183,In_2831);
and U460 (N_460,In_1347,In_2792);
nor U461 (N_461,In_2481,In_2905);
and U462 (N_462,In_2617,In_1603);
and U463 (N_463,In_2741,In_125);
xor U464 (N_464,In_452,In_460);
nor U465 (N_465,In_2008,In_2586);
or U466 (N_466,In_1672,In_1007);
xor U467 (N_467,In_1547,In_2001);
xor U468 (N_468,In_188,In_851);
xnor U469 (N_469,In_1528,In_2737);
nand U470 (N_470,In_2669,In_2269);
and U471 (N_471,In_1089,In_1138);
or U472 (N_472,In_873,In_809);
nor U473 (N_473,In_2749,In_2240);
or U474 (N_474,In_112,In_2409);
or U475 (N_475,In_1301,In_1034);
and U476 (N_476,In_1526,In_1587);
and U477 (N_477,In_1238,In_1066);
xnor U478 (N_478,In_1718,In_2625);
nor U479 (N_479,In_2197,In_853);
and U480 (N_480,In_2612,In_1026);
nor U481 (N_481,In_2777,In_1794);
xnor U482 (N_482,In_1702,In_886);
nor U483 (N_483,In_1087,In_786);
xor U484 (N_484,In_740,In_103);
or U485 (N_485,In_2416,In_2804);
or U486 (N_486,In_1014,In_2407);
or U487 (N_487,In_62,In_397);
and U488 (N_488,In_2058,In_783);
nand U489 (N_489,In_1585,In_1230);
nand U490 (N_490,In_2036,In_2224);
xor U491 (N_491,In_1768,In_1883);
nor U492 (N_492,In_2692,In_2984);
or U493 (N_493,In_1810,In_2251);
and U494 (N_494,In_501,In_981);
and U495 (N_495,In_423,In_1378);
xnor U496 (N_496,In_1704,In_2945);
nor U497 (N_497,In_1126,In_1982);
or U498 (N_498,In_1757,In_2620);
and U499 (N_499,In_2149,In_666);
or U500 (N_500,In_1028,In_429);
or U501 (N_501,In_1339,In_2466);
nand U502 (N_502,In_1095,In_2);
nor U503 (N_503,In_1819,In_2225);
xnor U504 (N_504,In_1467,In_2627);
or U505 (N_505,In_2523,In_1748);
xor U506 (N_506,In_819,In_592);
and U507 (N_507,In_2360,In_986);
nand U508 (N_508,In_1901,In_2665);
nand U509 (N_509,In_1970,In_1965);
xnor U510 (N_510,In_1078,In_273);
xnor U511 (N_511,In_2755,In_560);
nor U512 (N_512,In_1891,In_34);
nor U513 (N_513,In_2662,In_750);
nor U514 (N_514,In_1121,In_2025);
nand U515 (N_515,In_745,In_2779);
or U516 (N_516,In_531,In_2922);
nor U517 (N_517,In_1635,In_1081);
nand U518 (N_518,In_461,In_1284);
or U519 (N_519,In_2609,In_2333);
nor U520 (N_520,In_2101,In_2426);
nand U521 (N_521,In_2433,In_186);
or U522 (N_522,In_1978,In_2476);
xor U523 (N_523,In_1027,In_715);
xor U524 (N_524,In_548,In_1393);
and U525 (N_525,In_485,In_827);
xnor U526 (N_526,In_1893,In_1179);
nand U527 (N_527,In_2347,In_1194);
and U528 (N_528,In_1072,In_738);
nor U529 (N_529,In_1024,In_1088);
and U530 (N_530,In_2187,In_1127);
or U531 (N_531,In_1590,In_92);
or U532 (N_532,In_2168,In_1433);
nand U533 (N_533,In_856,In_741);
and U534 (N_534,In_1195,In_1610);
nand U535 (N_535,In_2806,In_900);
xor U536 (N_536,In_1963,In_2629);
nand U537 (N_537,In_778,In_1607);
or U538 (N_538,In_1132,In_1803);
or U539 (N_539,In_1992,In_2239);
or U540 (N_540,In_2208,In_2410);
nor U541 (N_541,In_2060,In_1728);
xor U542 (N_542,In_1310,In_30);
xnor U543 (N_543,In_295,In_2175);
nand U544 (N_544,In_2740,In_613);
nand U545 (N_545,In_1011,In_2307);
nor U546 (N_546,In_2784,In_2392);
and U547 (N_547,In_796,In_600);
xnor U548 (N_548,In_919,In_318);
nand U549 (N_549,In_1240,In_415);
nand U550 (N_550,In_283,In_1779);
xor U551 (N_551,In_143,In_1837);
nand U552 (N_552,In_952,In_433);
nor U553 (N_553,In_1720,In_990);
or U554 (N_554,In_2799,In_899);
nor U555 (N_555,In_337,In_1990);
nand U556 (N_556,In_1664,In_1067);
nor U557 (N_557,In_2956,In_1816);
and U558 (N_558,In_814,In_863);
nor U559 (N_559,In_1060,In_730);
nand U560 (N_560,In_2191,In_573);
and U561 (N_561,In_2658,In_1358);
nand U562 (N_562,In_2373,In_1418);
xnor U563 (N_563,In_932,In_2638);
xor U564 (N_564,In_154,In_262);
and U565 (N_565,In_2714,In_1448);
nand U566 (N_566,In_2841,In_1582);
and U567 (N_567,In_1269,In_815);
or U568 (N_568,In_2903,In_596);
nand U569 (N_569,In_1629,In_1821);
nand U570 (N_570,In_1599,In_688);
nand U571 (N_571,In_465,In_2116);
or U572 (N_572,In_978,In_1466);
or U573 (N_573,In_1899,In_1838);
nor U574 (N_574,In_2331,In_729);
xnor U575 (N_575,In_828,In_2434);
nor U576 (N_576,In_1967,In_1166);
and U577 (N_577,In_2507,In_2171);
nor U578 (N_578,In_43,In_180);
nand U579 (N_579,In_1687,In_1655);
nor U580 (N_580,In_225,In_1260);
xor U581 (N_581,In_2940,In_1141);
nand U582 (N_582,In_319,In_2076);
nand U583 (N_583,In_521,In_2910);
or U584 (N_584,In_1552,In_457);
nand U585 (N_585,In_2057,In_617);
and U586 (N_586,In_1509,In_2785);
xor U587 (N_587,In_2850,In_1054);
or U588 (N_588,In_2823,In_422);
xnor U589 (N_589,In_1533,In_565);
nor U590 (N_590,In_858,In_2848);
xor U591 (N_591,In_998,In_288);
xor U592 (N_592,In_2345,In_2673);
nor U593 (N_593,In_1342,In_2574);
nor U594 (N_594,In_1070,In_2990);
nor U595 (N_595,In_1140,In_1611);
or U596 (N_596,In_654,In_1076);
and U597 (N_597,In_191,In_684);
nand U598 (N_598,In_2424,In_683);
nor U599 (N_599,In_1619,In_309);
nor U600 (N_600,In_2633,In_2157);
nor U601 (N_601,In_2884,In_1453);
or U602 (N_602,In_443,In_1507);
and U603 (N_603,In_474,In_980);
nand U604 (N_604,In_2738,In_2474);
nor U605 (N_605,In_2326,In_1661);
or U606 (N_606,In_1841,In_459);
xor U607 (N_607,In_2563,In_2070);
nand U608 (N_608,In_2203,In_211);
nor U609 (N_609,In_428,In_808);
nand U610 (N_610,In_2192,In_2717);
nand U611 (N_611,In_2824,In_2162);
or U612 (N_612,In_1716,In_104);
and U613 (N_613,In_2235,In_1345);
nand U614 (N_614,In_2958,In_2798);
nor U615 (N_615,In_219,In_791);
nand U616 (N_616,In_780,In_770);
nand U617 (N_617,In_874,In_2754);
and U618 (N_618,In_748,In_1688);
nand U619 (N_619,In_2565,In_1013);
nor U620 (N_620,In_2721,In_672);
xnor U621 (N_621,In_450,In_2769);
xnor U622 (N_622,In_56,In_832);
and U623 (N_623,In_11,In_963);
xnor U624 (N_624,In_574,In_237);
or U625 (N_625,In_2654,In_1553);
or U626 (N_626,In_1350,In_1829);
or U627 (N_627,In_2037,In_1368);
nand U628 (N_628,In_2095,In_2275);
xor U629 (N_629,In_2247,In_1403);
nor U630 (N_630,In_1207,In_371);
or U631 (N_631,In_582,In_419);
nand U632 (N_632,In_72,In_425);
or U633 (N_633,In_1524,In_2202);
or U634 (N_634,In_2454,In_2635);
or U635 (N_635,In_1747,In_2309);
and U636 (N_636,In_1846,In_2374);
or U637 (N_637,In_1822,In_1468);
and U638 (N_638,In_1588,In_879);
nor U639 (N_639,In_676,In_1118);
nand U640 (N_640,In_2327,In_2114);
nand U641 (N_641,In_1885,In_1421);
and U642 (N_642,In_277,In_2146);
and U643 (N_643,In_1424,In_587);
and U644 (N_644,In_1583,In_250);
nand U645 (N_645,In_1852,In_765);
or U646 (N_646,In_2765,In_1778);
or U647 (N_647,In_984,In_2044);
or U648 (N_648,In_665,In_1387);
xor U649 (N_649,In_2907,In_352);
nand U650 (N_650,In_2119,In_503);
nor U651 (N_651,In_1295,In_2953);
and U652 (N_652,In_1719,In_1266);
xor U653 (N_653,In_1693,In_1340);
nand U654 (N_654,In_2727,In_1999);
nand U655 (N_655,In_829,In_2458);
and U656 (N_656,In_2200,In_1363);
or U657 (N_657,In_1501,In_325);
nand U658 (N_658,In_824,In_2967);
nor U659 (N_659,In_1750,In_1142);
or U660 (N_660,In_2027,In_1356);
xnor U661 (N_661,In_1258,In_2846);
nor U662 (N_662,In_1556,In_2585);
xnor U663 (N_663,In_2948,In_1381);
nand U664 (N_664,In_608,In_807);
nand U665 (N_665,In_2619,In_409);
nand U666 (N_666,In_2313,In_2616);
or U667 (N_667,In_2180,In_1259);
nand U668 (N_668,In_1069,In_1536);
and U669 (N_669,In_2936,In_1707);
and U670 (N_670,In_1644,In_1409);
or U671 (N_671,In_1139,In_196);
nand U672 (N_672,In_2007,In_516);
xor U673 (N_673,In_1818,In_2613);
and U674 (N_674,In_2061,In_2880);
or U675 (N_675,In_2783,In_1680);
nor U676 (N_676,In_694,In_1346);
nor U677 (N_677,In_19,In_152);
or U678 (N_678,In_2314,In_2713);
nand U679 (N_679,In_550,In_20);
nand U680 (N_680,In_1871,In_1622);
nor U681 (N_681,In_618,In_1513);
or U682 (N_682,In_2825,In_1542);
or U683 (N_683,In_2937,In_1261);
or U684 (N_684,In_268,In_2700);
nand U685 (N_685,In_1831,In_1274);
nor U686 (N_686,In_732,In_2311);
or U687 (N_687,In_845,In_870);
nor U688 (N_688,In_416,In_1804);
nand U689 (N_689,In_2595,In_2390);
xor U690 (N_690,In_579,In_2028);
and U691 (N_691,In_1946,In_1878);
xor U692 (N_692,In_837,In_157);
nand U693 (N_693,In_1068,In_736);
nand U694 (N_694,In_190,In_547);
xnor U695 (N_695,In_2802,In_1408);
and U696 (N_696,In_2836,In_2473);
and U697 (N_697,In_2584,In_2412);
xor U698 (N_698,In_1167,In_2774);
nand U699 (N_699,In_2461,In_1723);
and U700 (N_700,In_1995,In_2026);
nand U701 (N_701,In_784,In_1923);
and U702 (N_702,In_2404,In_95);
xnor U703 (N_703,In_622,In_1484);
nor U704 (N_704,In_540,In_1313);
or U705 (N_705,In_2350,In_1842);
and U706 (N_706,In_2328,In_274);
and U707 (N_707,In_733,In_2590);
nor U708 (N_708,In_1873,In_1282);
nand U709 (N_709,In_208,In_2664);
or U710 (N_710,In_1777,In_2497);
or U711 (N_711,In_1633,In_1881);
xnor U712 (N_712,In_2852,In_2878);
nand U713 (N_713,In_1422,In_1979);
xor U714 (N_714,In_1116,In_1287);
or U715 (N_715,In_1192,In_2357);
or U716 (N_716,In_751,In_2780);
xor U717 (N_717,In_971,In_747);
xnor U718 (N_718,In_249,In_1406);
xor U719 (N_719,In_2138,In_2844);
nand U720 (N_720,In_1811,In_1472);
nand U721 (N_721,In_1174,In_1052);
and U722 (N_722,In_1372,In_1244);
nor U723 (N_723,In_1855,In_797);
nand U724 (N_724,In_129,In_1887);
xor U725 (N_725,In_1936,In_2372);
nor U726 (N_726,In_1564,In_2339);
xor U727 (N_727,In_2430,In_1496);
xor U728 (N_728,In_955,In_171);
nor U729 (N_729,In_1569,In_2144);
xor U730 (N_730,In_2704,In_2723);
nor U731 (N_731,In_1001,In_468);
nor U732 (N_732,In_2909,In_1835);
nand U733 (N_733,In_2472,In_1123);
and U734 (N_734,In_2135,In_992);
xor U735 (N_735,In_2323,In_269);
nor U736 (N_736,In_349,In_1529);
nand U737 (N_737,In_1217,In_705);
xor U738 (N_738,In_1920,In_178);
xor U739 (N_739,In_675,In_2957);
and U740 (N_740,In_2708,In_116);
or U741 (N_741,In_921,In_2666);
or U742 (N_742,In_1551,In_576);
and U743 (N_743,In_895,In_948);
or U744 (N_744,In_447,In_894);
or U745 (N_745,In_1460,In_2513);
or U746 (N_746,In_2908,In_2494);
and U747 (N_747,In_1998,In_2227);
xor U748 (N_748,In_2341,In_1966);
nor U749 (N_749,In_1749,In_2508);
nand U750 (N_750,In_1915,In_1213);
nand U751 (N_751,In_1035,In_2883);
xor U752 (N_752,In_2398,In_1597);
xor U753 (N_753,In_1362,In_120);
nor U754 (N_754,In_1572,In_98);
and U755 (N_755,In_491,In_2257);
and U756 (N_756,In_2266,In_376);
nor U757 (N_757,In_1291,In_17);
nor U758 (N_758,In_338,In_1732);
nand U759 (N_759,In_1734,In_1737);
xor U760 (N_760,In_515,In_506);
nand U761 (N_761,In_505,In_1490);
or U762 (N_762,In_1543,In_63);
and U763 (N_763,In_1377,In_1447);
or U764 (N_764,In_1733,In_424);
nand U765 (N_765,In_1993,In_908);
nor U766 (N_766,In_581,In_1698);
nand U767 (N_767,In_965,In_2301);
or U768 (N_768,In_1865,In_1385);
nor U769 (N_769,In_931,In_2659);
and U770 (N_770,In_2437,In_742);
nand U771 (N_771,In_2610,In_779);
or U772 (N_772,In_1338,In_421);
or U773 (N_773,In_2942,In_927);
and U774 (N_774,In_2352,In_2368);
and U775 (N_775,In_728,In_320);
nand U776 (N_776,In_1678,In_1135);
or U777 (N_777,In_2621,In_1486);
nor U778 (N_778,In_2298,In_2050);
xor U779 (N_779,In_2842,In_1197);
nand U780 (N_780,In_1793,In_18);
nand U781 (N_781,In_940,In_299);
nor U782 (N_782,In_1018,In_1575);
or U783 (N_783,In_442,In_31);
xnor U784 (N_784,In_1304,In_1740);
or U785 (N_785,In_752,In_1796);
or U786 (N_786,In_2134,In_1315);
xor U787 (N_787,In_169,In_1669);
xnor U788 (N_788,In_1898,In_1191);
nand U789 (N_789,In_2366,In_308);
nand U790 (N_790,In_2478,In_65);
nor U791 (N_791,In_1292,In_1183);
nor U792 (N_792,In_470,In_2682);
or U793 (N_793,In_911,In_1341);
xnor U794 (N_794,In_812,In_2807);
or U795 (N_795,In_663,In_40);
nand U796 (N_796,In_1648,In_841);
xnor U797 (N_797,In_2789,In_357);
or U798 (N_798,In_2725,In_203);
nor U799 (N_799,In_988,In_2961);
nor U800 (N_800,In_1394,In_1104);
nand U801 (N_801,In_1190,In_2132);
xor U802 (N_802,In_983,In_2515);
and U803 (N_803,In_1379,In_1392);
or U804 (N_804,In_2950,In_1158);
and U805 (N_805,In_73,In_2566);
nor U806 (N_806,In_2768,In_585);
and U807 (N_807,In_1616,In_2973);
nor U808 (N_808,In_144,In_44);
or U809 (N_809,In_176,In_2759);
nor U810 (N_810,In_499,In_2955);
or U811 (N_811,In_60,In_9);
nand U812 (N_812,In_555,In_2342);
or U813 (N_813,In_1875,In_1972);
nor U814 (N_814,In_1211,In_1671);
or U815 (N_815,In_1996,In_1530);
nand U816 (N_816,In_1206,In_1425);
nor U817 (N_817,In_231,In_1625);
xor U818 (N_818,In_2553,In_1493);
xnor U819 (N_819,In_2367,In_168);
xor U820 (N_820,In_737,In_1506);
nand U821 (N_821,In_2750,In_556);
nor U822 (N_822,In_2863,In_217);
or U823 (N_823,In_685,In_2843);
or U824 (N_824,In_2681,In_2919);
or U825 (N_825,In_2152,In_2965);
nand U826 (N_826,In_2697,In_1189);
or U827 (N_827,In_27,In_1429);
and U828 (N_828,In_2949,In_896);
nor U829 (N_829,In_136,In_883);
nand U830 (N_830,In_2868,In_1934);
or U831 (N_831,In_500,In_146);
nor U832 (N_832,In_1102,In_260);
and U833 (N_833,In_1862,In_373);
nand U834 (N_834,In_2655,In_1763);
nor U835 (N_835,In_187,In_1419);
nand U836 (N_836,In_2369,In_1606);
xnor U837 (N_837,In_1700,In_2976);
xnor U838 (N_838,In_2383,In_838);
nand U839 (N_839,In_1520,In_2087);
and U840 (N_840,In_286,In_994);
xnor U841 (N_841,In_1407,In_1880);
xnor U842 (N_842,In_1951,In_2501);
or U843 (N_843,In_936,In_2459);
nor U844 (N_844,In_1823,In_945);
nand U845 (N_845,In_2421,In_2022);
nand U846 (N_846,In_289,In_2246);
nand U847 (N_847,In_970,In_1888);
xor U848 (N_848,In_2163,In_2912);
and U849 (N_849,In_122,In_2094);
nand U850 (N_850,In_535,In_2464);
and U851 (N_851,In_2009,In_2904);
or U852 (N_852,In_484,In_1815);
xor U853 (N_853,In_1012,In_601);
and U854 (N_854,In_2042,In_266);
or U855 (N_855,In_1813,In_1400);
and U856 (N_856,In_358,In_398);
nand U857 (N_857,In_2415,In_2601);
or U858 (N_858,In_2294,In_1866);
xnor U859 (N_859,In_2015,In_25);
or U860 (N_860,In_253,In_2182);
or U861 (N_861,In_2901,In_1986);
and U862 (N_862,In_1557,In_1262);
nor U863 (N_863,In_2827,In_1722);
nor U864 (N_864,In_1608,In_400);
xnor U865 (N_865,In_2394,In_892);
or U866 (N_866,In_2489,In_590);
nand U867 (N_867,In_2063,In_2268);
or U868 (N_868,In_200,In_1851);
nand U869 (N_869,In_1383,In_568);
xor U870 (N_870,In_2195,In_721);
xnor U871 (N_871,In_854,In_29);
nand U872 (N_872,In_1742,In_2766);
and U873 (N_873,In_137,In_2174);
nand U874 (N_874,In_2220,In_2440);
xnor U875 (N_875,In_202,In_1874);
and U876 (N_876,In_652,In_1864);
or U877 (N_877,In_2762,In_401);
or U878 (N_878,In_2911,In_2929);
xor U879 (N_879,In_222,In_2859);
xor U880 (N_880,In_588,In_1828);
nor U881 (N_881,In_2828,In_2223);
and U882 (N_882,In_1198,In_852);
xnor U883 (N_883,In_2986,In_2245);
or U884 (N_884,In_699,In_865);
or U885 (N_885,In_691,In_2678);
or U886 (N_886,In_2158,In_2334);
and U887 (N_887,In_947,In_2532);
and U888 (N_888,In_2232,In_2514);
xnor U889 (N_889,In_270,In_2530);
nand U890 (N_890,In_426,In_2567);
nor U891 (N_891,In_2775,In_1143);
xnor U892 (N_892,In_1485,In_275);
xor U893 (N_893,In_1079,In_1436);
nand U894 (N_894,In_2877,In_354);
xnor U895 (N_895,In_2105,In_2701);
xor U896 (N_896,In_727,In_2348);
xnor U897 (N_897,In_306,In_1968);
and U898 (N_898,In_195,In_1498);
or U899 (N_899,In_1435,In_513);
nor U900 (N_900,In_79,In_280);
or U901 (N_901,In_392,In_2073);
nor U902 (N_902,In_91,In_2542);
xnor U903 (N_903,In_1201,In_105);
and U904 (N_904,In_1508,In_2605);
xnor U905 (N_905,In_1638,In_1774);
nor U906 (N_906,In_1721,In_1020);
nand U907 (N_907,In_300,In_959);
and U908 (N_908,In_1045,In_680);
and U909 (N_909,In_746,In_1343);
xor U910 (N_910,In_2234,In_1515);
nor U911 (N_911,In_2970,In_1663);
or U912 (N_912,In_1954,In_855);
or U913 (N_913,In_866,In_934);
nor U914 (N_914,In_1222,In_2705);
and U915 (N_915,In_2325,In_2414);
nand U916 (N_916,In_882,In_1427);
nor U917 (N_917,In_868,In_1861);
and U918 (N_918,In_1296,In_1417);
nor U919 (N_919,In_635,In_1334);
xnor U920 (N_920,In_1010,In_2696);
xnor U921 (N_921,In_2411,In_1867);
and U922 (N_922,In_243,In_941);
nor U923 (N_923,In_767,In_558);
nand U924 (N_924,In_189,In_619);
or U925 (N_925,In_1411,In_42);
nor U926 (N_926,In_1989,In_1534);
xnor U927 (N_927,In_1900,In_22);
nand U928 (N_928,In_1563,In_2856);
nand U929 (N_929,In_915,In_173);
or U930 (N_930,In_290,In_388);
and U931 (N_931,In_2040,In_387);
xnor U932 (N_932,In_692,In_2926);
nand U933 (N_933,In_1367,In_1691);
xnor U934 (N_934,In_327,In_2966);
or U935 (N_935,In_410,In_1082);
nand U936 (N_936,In_1146,In_757);
and U937 (N_937,In_1154,In_875);
nor U938 (N_938,In_1666,In_1136);
xnor U939 (N_939,In_2336,In_359);
xnor U940 (N_940,In_2069,In_232);
nand U941 (N_941,In_2787,In_133);
nor U942 (N_942,In_2643,In_958);
nand U943 (N_943,In_1318,In_711);
or U944 (N_944,In_2818,In_1636);
nor U945 (N_945,In_1103,In_1030);
nand U946 (N_946,In_1320,In_857);
nor U947 (N_947,In_1071,In_557);
nand U948 (N_948,In_1637,In_1137);
nand U949 (N_949,In_2687,In_1786);
or U950 (N_950,In_2097,In_1849);
or U951 (N_951,In_2389,In_41);
nor U952 (N_952,In_420,In_2085);
xnor U953 (N_953,In_2935,In_554);
or U954 (N_954,In_2236,In_1772);
xor U955 (N_955,In_28,In_150);
nor U956 (N_956,In_312,In_1031);
nor U957 (N_957,In_1814,In_1943);
and U958 (N_958,In_2284,In_472);
or U959 (N_959,In_2810,In_653);
nor U960 (N_960,In_1489,In_1770);
and U961 (N_961,In_2522,In_890);
xor U962 (N_962,In_1570,In_2160);
or U963 (N_963,In_2688,In_1964);
nor U964 (N_964,In_1927,In_1519);
nor U965 (N_965,In_2573,In_1904);
xnor U966 (N_966,In_109,In_2124);
or U967 (N_967,In_861,In_1654);
xnor U968 (N_968,In_566,In_36);
xor U969 (N_969,In_2065,In_303);
or U970 (N_970,In_1050,In_1940);
and U971 (N_971,In_2420,In_2667);
and U972 (N_972,In_2137,In_487);
nand U973 (N_973,In_661,In_1397);
and U974 (N_974,In_834,In_394);
xnor U975 (N_975,In_2425,In_2049);
nor U976 (N_976,In_2122,In_1330);
nor U977 (N_977,In_1327,In_201);
or U978 (N_978,In_2599,In_2600);
nand U979 (N_979,In_2363,In_1);
xnor U980 (N_980,In_117,In_1361);
nor U981 (N_981,In_70,In_1232);
and U982 (N_982,In_1033,In_2159);
and U983 (N_983,In_2982,In_52);
nor U984 (N_984,In_2661,In_2743);
nor U985 (N_985,In_1917,In_1863);
and U986 (N_986,In_417,In_1075);
and U987 (N_987,In_279,In_1889);
nand U988 (N_988,In_223,In_1783);
and U989 (N_989,In_412,In_2527);
nor U990 (N_990,In_759,In_1659);
nor U991 (N_991,In_1820,In_1208);
and U992 (N_992,In_1097,In_1961);
nand U993 (N_993,In_68,In_2543);
nor U994 (N_994,In_1942,In_2228);
and U995 (N_995,In_1065,In_974);
xnor U996 (N_996,In_1962,In_701);
or U997 (N_997,In_49,In_2255);
and U998 (N_998,In_2109,In_2169);
nand U999 (N_999,In_2790,In_2892);
or U1000 (N_1000,In_2082,In_427);
nor U1001 (N_1001,N_300,N_161);
xor U1002 (N_1002,In_1384,N_629);
nand U1003 (N_1003,N_944,In_1756);
or U1004 (N_1004,In_1040,N_518);
or U1005 (N_1005,In_4,N_475);
or U1006 (N_1006,In_467,N_26);
and U1007 (N_1007,N_516,N_922);
nand U1008 (N_1008,In_2559,In_1945);
and U1009 (N_1009,In_124,N_73);
xor U1010 (N_1010,In_849,In_2290);
or U1011 (N_1011,In_2498,N_815);
nand U1012 (N_1012,N_643,N_728);
or U1013 (N_1013,In_2173,In_1695);
or U1014 (N_1014,N_184,N_362);
xor U1015 (N_1015,In_1450,N_896);
nand U1016 (N_1016,N_119,N_524);
xor U1017 (N_1017,In_1836,In_2077);
nand U1018 (N_1018,N_221,In_2204);
nor U1019 (N_1019,In_1091,N_128);
nor U1020 (N_1020,N_256,In_2329);
and U1021 (N_1021,N_808,In_2630);
or U1022 (N_1022,N_91,N_881);
xor U1023 (N_1023,N_575,In_1193);
or U1024 (N_1024,In_704,In_2872);
nor U1025 (N_1025,N_953,N_608);
nor U1026 (N_1026,N_250,In_637);
nand U1027 (N_1027,N_64,N_705);
nor U1028 (N_1028,In_612,N_359);
nor U1029 (N_1029,In_192,In_1609);
nor U1030 (N_1030,N_695,N_657);
xnor U1031 (N_1031,In_1270,N_955);
and U1032 (N_1032,N_548,N_282);
nor U1033 (N_1033,In_1870,In_642);
and U1034 (N_1034,N_938,N_770);
nor U1035 (N_1035,N_81,In_2475);
nor U1036 (N_1036,In_2865,In_2306);
xnor U1037 (N_1037,In_1300,N_644);
nand U1038 (N_1038,In_2075,N_794);
and U1039 (N_1039,N_685,In_368);
xnor U1040 (N_1040,N_950,In_982);
nand U1041 (N_1041,N_569,N_928);
nand U1042 (N_1042,N_649,In_1634);
or U1043 (N_1043,In_773,In_710);
nand U1044 (N_1044,N_840,N_980);
or U1045 (N_1045,In_2964,In_2703);
or U1046 (N_1046,In_2128,N_420);
nor U1047 (N_1047,In_257,In_708);
or U1048 (N_1048,N_176,In_884);
nor U1049 (N_1049,N_838,N_985);
and U1050 (N_1050,In_2196,N_552);
xnor U1051 (N_1051,N_61,N_777);
or U1052 (N_1052,In_1017,In_54);
nor U1053 (N_1053,N_156,N_688);
nand U1054 (N_1054,N_199,N_220);
nand U1055 (N_1055,In_1973,In_2580);
nor U1056 (N_1056,In_1366,N_913);
nor U1057 (N_1057,In_658,N_215);
nor U1058 (N_1058,N_973,N_212);
nand U1059 (N_1059,N_790,In_1131);
and U1060 (N_1060,N_178,N_7);
xnor U1061 (N_1061,N_1,N_145);
and U1062 (N_1062,In_1767,N_496);
or U1063 (N_1063,N_874,N_756);
nor U1064 (N_1064,N_563,In_464);
and U1065 (N_1065,In_2045,N_721);
or U1066 (N_1066,In_1277,In_224);
xor U1067 (N_1067,N_375,N_761);
nor U1068 (N_1068,N_138,In_627);
nor U1069 (N_1069,N_978,N_449);
xor U1070 (N_1070,In_2575,In_1840);
nand U1071 (N_1071,In_479,N_902);
nor U1072 (N_1072,In_23,N_718);
nor U1073 (N_1073,In_2445,N_851);
xnor U1074 (N_1074,N_646,N_886);
and U1075 (N_1075,N_338,In_365);
and U1076 (N_1076,In_1151,In_1817);
or U1077 (N_1077,N_807,In_504);
nand U1078 (N_1078,N_885,N_912);
xnor U1079 (N_1079,In_2598,In_1423);
and U1080 (N_1080,N_933,N_610);
nor U1081 (N_1081,In_1311,N_366);
nand U1082 (N_1082,N_899,N_605);
nor U1083 (N_1083,N_574,In_2603);
or U1084 (N_1084,N_943,N_847);
and U1085 (N_1085,N_484,N_15);
or U1086 (N_1086,N_547,N_196);
nand U1087 (N_1087,In_2417,In_917);
and U1088 (N_1088,N_759,N_787);
xor U1089 (N_1089,In_2858,In_1107);
nand U1090 (N_1090,N_426,N_941);
nand U1091 (N_1091,In_2038,In_569);
and U1092 (N_1092,In_408,N_455);
or U1093 (N_1093,In_1938,N_616);
or U1094 (N_1094,In_2918,In_1974);
nor U1095 (N_1095,N_755,N_782);
xnor U1096 (N_1096,In_2408,In_395);
and U1097 (N_1097,N_488,In_2544);
and U1098 (N_1098,N_668,In_115);
or U1099 (N_1099,In_1037,N_683);
or U1100 (N_1100,N_504,In_2496);
and U1101 (N_1101,In_2053,N_429);
or U1102 (N_1102,In_2242,N_419);
nand U1103 (N_1103,N_459,N_954);
and U1104 (N_1104,N_614,N_47);
xor U1105 (N_1105,In_537,In_620);
nor U1106 (N_1106,N_502,N_725);
nor U1107 (N_1107,N_799,N_820);
nor U1108 (N_1108,In_1922,In_2488);
nor U1109 (N_1109,In_549,N_193);
and U1110 (N_1110,N_141,N_478);
nand U1111 (N_1111,In_2864,N_869);
xnor U1112 (N_1112,In_1169,In_2691);
nor U1113 (N_1113,In_577,In_572);
or U1114 (N_1114,N_336,In_956);
or U1115 (N_1115,In_199,N_930);
and U1116 (N_1116,N_805,N_473);
or U1117 (N_1117,In_2020,In_2172);
xor U1118 (N_1118,In_1879,N_318);
and U1119 (N_1119,N_121,In_774);
nand U1120 (N_1120,In_584,N_587);
xor U1121 (N_1121,In_2835,In_2292);
nand U1122 (N_1122,In_1220,N_636);
or U1123 (N_1123,In_1650,N_696);
or U1124 (N_1124,N_771,In_1336);
and U1125 (N_1125,In_1016,In_13);
xnor U1126 (N_1126,N_890,In_326);
nor U1127 (N_1127,In_2736,N_783);
or U1128 (N_1128,In_2932,In_489);
xor U1129 (N_1129,In_1178,N_775);
xnor U1130 (N_1130,In_2891,In_2401);
nand U1131 (N_1131,N_158,In_2002);
or U1132 (N_1132,N_28,In_216);
nor U1133 (N_1133,In_2760,N_554);
xnor U1134 (N_1134,N_804,In_518);
nand U1135 (N_1135,N_897,In_1371);
or U1136 (N_1136,In_2384,In_670);
xnor U1137 (N_1137,In_2467,In_1539);
nand U1138 (N_1138,N_861,N_270);
and U1139 (N_1139,N_909,In_1675);
nor U1140 (N_1140,N_17,In_2318);
nand U1141 (N_1141,N_400,In_1251);
or U1142 (N_1142,N_261,In_532);
or U1143 (N_1143,In_1640,In_1464);
nor U1144 (N_1144,In_1243,N_549);
and U1145 (N_1145,N_583,N_381);
and U1146 (N_1146,N_450,In_1984);
nor U1147 (N_1147,In_1673,N_186);
or U1148 (N_1148,N_124,N_3);
nor U1149 (N_1149,N_120,In_135);
nand U1150 (N_1150,N_910,In_967);
xnor U1151 (N_1151,In_607,N_273);
nand U1152 (N_1152,N_527,N_892);
xor U1153 (N_1153,In_2427,In_2267);
nor U1154 (N_1154,N_126,N_54);
nand U1155 (N_1155,In_1807,N_50);
xor U1156 (N_1156,N_507,In_1273);
nor U1157 (N_1157,In_2096,In_406);
xnor U1158 (N_1158,In_643,N_650);
nor U1159 (N_1159,In_1481,N_530);
and U1160 (N_1160,N_829,In_1510);
or U1161 (N_1161,N_468,In_2830);
xor U1162 (N_1162,N_613,In_2346);
and U1163 (N_1163,N_264,In_3);
xor U1164 (N_1164,In_659,In_1237);
nor U1165 (N_1165,In_2695,N_285);
and U1166 (N_1166,N_424,N_894);
nor U1167 (N_1167,N_316,N_606);
and U1168 (N_1168,N_251,N_41);
xnor U1169 (N_1169,N_324,N_494);
nand U1170 (N_1170,N_914,In_2539);
nor U1171 (N_1171,In_214,In_1199);
or U1172 (N_1172,N_265,N_170);
nand U1173 (N_1173,In_929,In_2902);
nand U1174 (N_1174,N_255,N_862);
nor U1175 (N_1175,N_414,N_681);
or U1176 (N_1176,In_846,In_2786);
or U1177 (N_1177,N_809,In_1046);
nor U1178 (N_1178,N_287,In_1226);
and U1179 (N_1179,In_240,In_494);
nor U1180 (N_1180,N_952,In_800);
nand U1181 (N_1181,In_1877,N_200);
and U1182 (N_1182,N_591,In_2604);
and U1183 (N_1183,N_32,In_1997);
and U1184 (N_1184,N_908,N_505);
xnor U1185 (N_1185,N_403,In_1912);
and U1186 (N_1186,N_694,N_389);
or U1187 (N_1187,N_738,In_1098);
xor U1188 (N_1188,In_252,In_1312);
xor U1189 (N_1189,In_2518,N_497);
nand U1190 (N_1190,N_715,N_611);
nand U1191 (N_1191,N_96,In_2724);
xor U1192 (N_1192,N_364,In_1241);
xnor U1193 (N_1193,In_1349,N_879);
nand U1194 (N_1194,In_2140,In_204);
nor U1195 (N_1195,In_949,In_690);
nand U1196 (N_1196,In_1248,N_736);
and U1197 (N_1197,N_187,N_931);
or U1198 (N_1198,In_218,N_489);
xor U1199 (N_1199,N_873,N_626);
and U1200 (N_1200,N_871,N_163);
nor U1201 (N_1201,N_240,In_2869);
nor U1202 (N_1202,N_93,N_986);
and U1203 (N_1203,In_402,In_374);
nand U1204 (N_1204,N_561,N_385);
xnor U1205 (N_1205,In_1969,N_546);
nand U1206 (N_1206,N_198,In_75);
nand U1207 (N_1207,In_1614,In_1219);
and U1208 (N_1208,N_737,N_335);
and U1209 (N_1209,N_355,N_560);
xnor U1210 (N_1210,In_570,N_461);
xor U1211 (N_1211,N_956,N_172);
or U1212 (N_1212,In_714,N_483);
nor U1213 (N_1213,In_1558,In_2218);
nor U1214 (N_1214,N_144,In_1048);
nand U1215 (N_1215,N_571,N_208);
nor U1216 (N_1216,In_944,In_1628);
nand U1217 (N_1217,N_700,N_801);
and U1218 (N_1218,In_2047,In_1910);
and U1219 (N_1219,In_1360,N_916);
or U1220 (N_1220,N_149,N_729);
nand U1221 (N_1221,N_904,In_1971);
nor U1222 (N_1222,N_465,In_2711);
xor U1223 (N_1223,In_877,N_368);
or U1224 (N_1224,In_906,N_889);
or U1225 (N_1225,N_578,N_593);
or U1226 (N_1226,In_2998,N_108);
nand U1227 (N_1227,N_898,In_89);
and U1228 (N_1228,In_953,N_380);
and U1229 (N_1229,N_29,N_993);
or U1230 (N_1230,N_577,N_964);
or U1231 (N_1231,In_2933,N_276);
xnor U1232 (N_1232,N_620,In_2003);
xnor U1233 (N_1233,In_2324,In_1025);
or U1234 (N_1234,In_2744,N_445);
or U1235 (N_1235,N_321,N_490);
nand U1236 (N_1236,N_295,In_1043);
xor U1237 (N_1237,N_470,N_31);
nand U1238 (N_1238,N_181,N_989);
or U1239 (N_1239,N_592,N_749);
nand U1240 (N_1240,In_2608,N_105);
xnor U1241 (N_1241,N_747,N_699);
nand U1242 (N_1242,In_674,In_546);
nor U1243 (N_1243,N_900,N_325);
nand U1244 (N_1244,In_867,In_2645);
and U1245 (N_1245,In_393,In_1105);
nor U1246 (N_1246,In_2388,In_228);
nand U1247 (N_1247,In_2320,N_495);
nor U1248 (N_1248,N_183,In_46);
or U1249 (N_1249,N_523,N_987);
xnor U1250 (N_1250,In_2568,N_343);
and U1251 (N_1251,N_697,In_2718);
nor U1252 (N_1252,N_59,N_409);
nand U1253 (N_1253,N_383,In_1591);
nor U1254 (N_1254,In_1839,In_1461);
and U1255 (N_1255,In_640,N_34);
nand U1256 (N_1256,In_2690,In_492);
xor U1257 (N_1257,In_33,In_580);
and U1258 (N_1258,In_2689,N_297);
and U1259 (N_1259,N_618,In_660);
xor U1260 (N_1260,In_564,In_2952);
xor U1261 (N_1261,N_827,In_2917);
nor U1262 (N_1262,N_195,N_717);
nor U1263 (N_1263,In_553,N_788);
and U1264 (N_1264,In_2676,In_1305);
or U1265 (N_1265,N_224,N_106);
or U1266 (N_1266,In_1708,In_938);
or U1267 (N_1267,In_1449,In_1579);
nand U1268 (N_1268,In_1229,In_2924);
and U1269 (N_1269,In_1022,In_1792);
or U1270 (N_1270,In_1256,In_2921);
xor U1271 (N_1271,In_703,N_735);
nor U1272 (N_1272,In_1454,N_289);
nand U1273 (N_1273,N_152,In_1015);
and U1274 (N_1274,In_1051,In_497);
or U1275 (N_1275,N_337,In_817);
or U1276 (N_1276,In_490,N_525);
nand U1277 (N_1277,N_957,N_71);
nand U1278 (N_1278,In_2406,In_1711);
and U1279 (N_1279,In_2758,In_2778);
and U1280 (N_1280,N_966,N_111);
xor U1281 (N_1281,N_457,In_2452);
xor U1282 (N_1282,N_68,In_2110);
nand U1283 (N_1283,N_937,In_2288);
and U1284 (N_1284,In_1307,N_863);
and U1285 (N_1285,In_1589,In_1656);
xor U1286 (N_1286,N_217,N_607);
xnor U1287 (N_1287,N_617,N_849);
and U1288 (N_1288,In_772,In_1250);
or U1289 (N_1289,In_1843,In_2861);
nor U1290 (N_1290,In_2198,In_2359);
xnor U1291 (N_1291,In_1631,In_2534);
xnor U1292 (N_1292,In_2564,N_396);
nor U1293 (N_1293,N_806,In_82);
or U1294 (N_1294,N_216,N_584);
nand U1295 (N_1295,In_1290,In_2186);
and U1296 (N_1296,N_551,N_286);
nor U1297 (N_1297,N_222,In_2826);
nor U1298 (N_1298,N_982,In_771);
xnor U1299 (N_1299,N_655,N_57);
and U1300 (N_1300,N_180,N_349);
or U1301 (N_1301,N_627,N_155);
xor U1302 (N_1302,In_914,In_2446);
nand U1303 (N_1303,In_1686,N_392);
and U1304 (N_1304,N_162,N_731);
xor U1305 (N_1305,In_2289,In_1443);
nand U1306 (N_1306,In_198,N_786);
and U1307 (N_1307,In_2660,In_304);
nand U1308 (N_1308,N_487,N_875);
nor U1309 (N_1309,In_1729,N_13);
and U1310 (N_1310,N_544,In_1860);
xnor U1311 (N_1311,N_10,In_1326);
and U1312 (N_1312,In_1983,In_1994);
or U1313 (N_1313,In_2387,N_745);
xnor U1314 (N_1314,In_1170,N_893);
nand U1315 (N_1315,N_159,In_2980);
or U1316 (N_1316,In_645,N_792);
nor U1317 (N_1317,N_726,N_153);
xor U1318 (N_1318,In_1463,In_962);
nand U1319 (N_1319,In_2874,N_188);
and U1320 (N_1320,In_697,N_174);
xnor U1321 (N_1321,N_723,In_755);
nand U1322 (N_1322,In_1203,N_654);
or U1323 (N_1323,In_2249,N_290);
nor U1324 (N_1324,N_776,N_245);
and U1325 (N_1325,N_171,N_878);
nor U1326 (N_1326,In_1458,N_369);
nand U1327 (N_1327,In_1359,In_943);
or U1328 (N_1328,N_556,N_540);
xor U1329 (N_1329,N_559,N_880);
xnor U1330 (N_1330,N_907,In_58);
nand U1331 (N_1331,In_84,N_867);
nand U1332 (N_1332,N_422,In_2800);
and U1333 (N_1333,N_148,N_70);
xor U1334 (N_1334,N_82,In_1106);
or U1335 (N_1335,N_818,In_2583);
xor U1336 (N_1336,N_567,N_843);
nand U1337 (N_1337,In_880,In_2712);
nor U1338 (N_1338,In_2505,In_1176);
xor U1339 (N_1339,N_753,N_296);
nand U1340 (N_1340,In_1689,In_973);
and U1341 (N_1341,N_249,In_2795);
or U1342 (N_1342,In_16,In_2985);
and U1343 (N_1343,In_2418,N_440);
and U1344 (N_1344,N_582,N_272);
and U1345 (N_1345,In_2335,N_992);
xnor U1346 (N_1346,In_835,In_1325);
xnor U1347 (N_1347,N_929,N_493);
nor U1348 (N_1348,In_2354,N_711);
nor U1349 (N_1349,N_684,N_65);
xor U1350 (N_1350,N_305,In_836);
and U1351 (N_1351,N_326,In_1462);
nand U1352 (N_1352,In_2084,N_599);
nand U1353 (N_1353,In_1162,In_1329);
and U1354 (N_1354,N_994,In_2851);
nand U1355 (N_1355,In_209,In_1752);
or U1356 (N_1356,N_421,In_348);
nor U1357 (N_1357,In_1267,In_1322);
nand U1358 (N_1358,In_2622,In_1646);
or U1359 (N_1359,N_946,In_2262);
xor U1360 (N_1360,N_704,In_545);
xor U1361 (N_1361,N_959,In_926);
and U1362 (N_1362,N_485,N_298);
xnor U1363 (N_1363,N_205,N_781);
xor U1364 (N_1364,N_513,N_515);
and U1365 (N_1365,In_655,In_2429);
nor U1366 (N_1366,N_58,N_84);
or U1367 (N_1367,In_2897,In_413);
xnor U1368 (N_1368,In_1495,In_923);
xor U1369 (N_1369,In_2597,In_527);
and U1370 (N_1370,N_652,N_391);
and U1371 (N_1371,N_53,N_469);
xor U1372 (N_1372,N_750,In_816);
nand U1373 (N_1373,N_74,In_2675);
xnor U1374 (N_1374,In_539,N_204);
and U1375 (N_1375,In_1218,In_123);
or U1376 (N_1376,N_398,N_638);
xor U1377 (N_1377,In_842,N_9);
and U1378 (N_1378,In_2525,In_1063);
and U1379 (N_1379,In_1565,In_2271);
or U1380 (N_1380,N_977,In_541);
or U1381 (N_1381,N_23,In_1255);
nand U1382 (N_1382,In_1703,In_1164);
xor U1383 (N_1383,In_2129,In_2794);
or U1384 (N_1384,In_2649,In_2089);
xor U1385 (N_1385,In_2495,N_503);
or U1386 (N_1386,In_2303,In_471);
and U1387 (N_1387,In_2900,N_532);
or U1388 (N_1388,In_278,N_89);
or U1389 (N_1389,In_1632,N_565);
and U1390 (N_1390,In_233,In_989);
and U1391 (N_1391,In_244,N_207);
and U1392 (N_1392,In_2480,In_950);
and U1393 (N_1393,N_479,N_958);
and U1394 (N_1394,In_2549,N_519);
nand U1395 (N_1395,N_353,N_631);
or U1396 (N_1396,In_496,In_1502);
and U1397 (N_1397,In_614,In_725);
and U1398 (N_1398,N_659,N_203);
nand U1399 (N_1399,N_680,In_160);
and U1400 (N_1400,N_936,In_1913);
nor U1401 (N_1401,N_462,N_474);
xnor U1402 (N_1402,In_1853,N_888);
or U1403 (N_1403,N_660,N_79);
xnor U1404 (N_1404,N_137,N_573);
or U1405 (N_1405,In_1455,N_51);
xnor U1406 (N_1406,In_493,In_1668);
or U1407 (N_1407,N_939,In_1475);
xor U1408 (N_1408,In_2302,N_926);
nand U1409 (N_1409,N_363,In_604);
xor U1410 (N_1410,In_1809,N_118);
and U1411 (N_1411,N_127,In_265);
nor U1412 (N_1412,N_995,N_209);
and U1413 (N_1413,In_2282,In_1184);
nor U1414 (N_1414,N_595,In_2127);
and U1415 (N_1415,N_520,In_2272);
xnor U1416 (N_1416,In_1751,N_136);
nor U1417 (N_1417,In_2297,N_16);
nor U1418 (N_1418,N_114,In_1405);
or U1419 (N_1419,In_78,In_2499);
or U1420 (N_1420,N_860,N_246);
or U1421 (N_1421,N_866,N_63);
xnor U1422 (N_1422,In_787,N_101);
xor U1423 (N_1423,In_1431,N_390);
nand U1424 (N_1424,N_312,In_478);
or U1425 (N_1425,N_55,N_537);
xnor U1426 (N_1426,N_113,In_735);
or U1427 (N_1427,In_59,In_2091);
nand U1428 (N_1428,N_317,N_206);
xor U1429 (N_1429,N_2,In_2485);
and U1430 (N_1430,In_1566,In_1434);
or U1431 (N_1431,In_2439,In_1000);
or U1432 (N_1432,N_35,N_779);
nand U1433 (N_1433,N_87,In_2631);
nor U1434 (N_1434,In_2102,In_538);
xor U1435 (N_1435,In_1897,N_724);
xnor U1436 (N_1436,In_1684,In_1187);
nor U1437 (N_1437,N_664,In_1950);
nand U1438 (N_1438,In_591,In_2947);
xor U1439 (N_1439,In_229,In_2395);
nand U1440 (N_1440,In_1710,In_1959);
xor U1441 (N_1441,In_47,In_2431);
or U1442 (N_1442,In_811,In_2946);
and U1443 (N_1443,In_2449,N_331);
xnor U1444 (N_1444,In_2855,N_612);
nand U1445 (N_1445,N_437,N_466);
xnor U1446 (N_1446,N_601,N_883);
nor U1447 (N_1447,In_384,N_319);
nand U1448 (N_1448,N_315,N_395);
and U1449 (N_1449,N_39,In_719);
and U1450 (N_1450,N_30,In_1503);
and U1451 (N_1451,In_2618,In_483);
nor U1452 (N_1452,In_284,In_2672);
xor U1453 (N_1453,In_2377,N_734);
or U1454 (N_1454,N_232,N_5);
and U1455 (N_1455,N_826,In_1263);
xor U1456 (N_1456,In_2000,N_269);
nor U1457 (N_1457,In_93,N_634);
and U1458 (N_1458,In_818,In_1985);
nand U1459 (N_1459,N_247,In_559);
xor U1460 (N_1460,In_396,N_784);
and U1461 (N_1461,N_971,In_2642);
and U1462 (N_1462,In_121,N_238);
xor U1463 (N_1463,N_313,In_2397);
nor U1464 (N_1464,In_2442,In_2500);
xor U1465 (N_1465,N_11,In_1833);
xor U1466 (N_1466,N_746,In_1101);
nor U1467 (N_1467,In_1160,In_1055);
nand U1468 (N_1468,In_2742,N_134);
xor U1469 (N_1469,N_774,In_1980);
xnor U1470 (N_1470,N_670,In_2299);
nor U1471 (N_1471,In_1525,N_553);
nand U1472 (N_1472,N_828,N_895);
nand U1473 (N_1473,In_1491,In_2997);
or U1474 (N_1474,In_380,N_974);
or U1475 (N_1475,In_2080,N_763);
xnor U1476 (N_1476,N_686,N_408);
xor U1477 (N_1477,In_2018,In_2428);
nand U1478 (N_1478,N_687,N_906);
or U1479 (N_1479,In_2699,N_202);
xnor U1480 (N_1480,In_2088,In_163);
and U1481 (N_1481,N_72,N_999);
nand U1482 (N_1482,N_486,N_304);
and U1483 (N_1483,N_564,N_963);
xor U1484 (N_1484,In_913,N_865);
nor U1485 (N_1485,In_525,N_447);
and U1486 (N_1486,N_536,In_724);
xnor U1487 (N_1487,In_1370,In_1150);
xnor U1488 (N_1488,N_712,In_1047);
nand U1489 (N_1489,N_24,N_92);
nor U1490 (N_1490,N_190,In_1593);
nand U1491 (N_1491,In_2199,In_2054);
and U1492 (N_1492,In_2978,In_2756);
nor U1493 (N_1493,In_2726,In_454);
or U1494 (N_1494,N_334,In_1624);
or U1495 (N_1495,N_780,N_40);
nor U1496 (N_1496,In_918,In_723);
or U1497 (N_1497,In_1185,In_1905);
nor U1498 (N_1498,N_378,In_100);
and U1499 (N_1499,N_236,In_821);
nor U1500 (N_1500,N_472,N_842);
nand U1501 (N_1501,In_1321,In_207);
or U1502 (N_1502,In_1717,In_2993);
and U1503 (N_1503,N_291,In_1781);
nor U1504 (N_1504,N_541,N_361);
nor U1505 (N_1505,In_1667,N_965);
or U1506 (N_1506,N_323,N_557);
nand U1507 (N_1507,N_590,In_1516);
xor U1508 (N_1508,In_2857,In_111);
nor U1509 (N_1509,In_2375,N_214);
nor U1510 (N_1510,In_1554,N_675);
or U1511 (N_1511,In_2148,In_2968);
nand U1512 (N_1512,N_165,N_822);
and U1513 (N_1513,N_279,In_2142);
or U1514 (N_1514,N_500,In_1538);
xor U1515 (N_1515,N_911,In_339);
or U1516 (N_1516,N_481,In_2230);
nand U1517 (N_1517,In_788,In_1685);
nand U1518 (N_1518,In_2706,In_2052);
or U1519 (N_1519,N_676,N_360);
xnor U1520 (N_1520,N_918,N_95);
nand U1521 (N_1521,N_309,N_589);
xnor U1522 (N_1522,In_2557,In_1916);
or U1523 (N_1523,In_805,N_624);
xor U1524 (N_1524,N_168,N_18);
or U1525 (N_1525,In_939,In_221);
or U1526 (N_1526,N_327,N_751);
xor U1527 (N_1527,In_1935,In_174);
xor U1528 (N_1528,N_189,N_133);
nand U1529 (N_1529,N_585,N_115);
nor U1530 (N_1530,N_333,In_848);
and U1531 (N_1531,In_86,N_416);
or U1532 (N_1532,In_2463,In_878);
or U1533 (N_1533,In_1059,N_278);
or U1534 (N_1534,In_2181,N_522);
nor U1535 (N_1535,In_2241,N_901);
xor U1536 (N_1536,In_626,N_44);
xnor U1537 (N_1537,N_477,In_2259);
nand U1538 (N_1538,N_482,N_823);
nand U1539 (N_1539,In_1926,N_824);
nor U1540 (N_1540,In_1004,In_551);
or U1541 (N_1541,In_1743,In_1094);
xnor U1542 (N_1542,N_579,In_1627);
nand U1543 (N_1543,N_693,N_810);
nand U1544 (N_1544,N_678,In_1172);
or U1545 (N_1545,N_615,N_839);
or U1546 (N_1546,In_935,In_323);
xor U1547 (N_1547,N_748,N_830);
and U1548 (N_1548,N_243,In_2405);
and U1549 (N_1549,In_2226,In_77);
nand U1550 (N_1550,In_793,In_1848);
nand U1551 (N_1551,N_703,In_404);
nor U1552 (N_1552,In_2487,In_1348);
and U1553 (N_1553,N_46,N_371);
and U1554 (N_1554,N_399,N_185);
xnor U1555 (N_1555,N_555,In_381);
xor U1556 (N_1556,N_464,In_624);
or U1557 (N_1557,N_374,N_920);
or U1558 (N_1558,N_637,N_550);
xnor U1559 (N_1559,N_850,N_534);
xnor U1560 (N_1560,N_379,N_714);
nand U1561 (N_1561,In_2468,N_130);
and U1562 (N_1562,N_692,In_2136);
nand U1563 (N_1563,In_2316,N_940);
or U1564 (N_1564,In_583,N_354);
nand U1565 (N_1565,In_2801,In_1390);
nand U1566 (N_1566,N_597,N_672);
nand U1567 (N_1567,N_713,N_14);
nor U1568 (N_1568,In_603,N_98);
nand U1569 (N_1569,N_800,In_1907);
nand U1570 (N_1570,In_276,In_313);
nor U1571 (N_1571,In_2456,In_1254);
xnor U1572 (N_1572,In_2820,In_362);
nand U1573 (N_1573,In_785,N_979);
or U1574 (N_1574,In_2960,N_173);
and U1575 (N_1575,N_259,In_1911);
nand U1576 (N_1576,N_129,In_510);
and U1577 (N_1577,N_658,In_1413);
or U1578 (N_1578,In_370,N_262);
nand U1579 (N_1579,In_1736,N_757);
and U1580 (N_1580,N_811,In_2322);
and U1581 (N_1581,In_543,N_102);
nand U1582 (N_1582,In_669,N_976);
xnor U1583 (N_1583,In_1937,N_373);
or U1584 (N_1584,N_813,In_90);
nand U1585 (N_1585,N_635,In_1188);
nor U1586 (N_1586,N_441,In_1445);
nand U1587 (N_1587,N_509,N_132);
xnor U1588 (N_1588,N_848,N_142);
or U1589 (N_1589,In_7,In_1791);
xnor U1590 (N_1590,N_125,In_2033);
nand U1591 (N_1591,N_283,In_2164);
and U1592 (N_1592,In_1280,N_708);
or U1593 (N_1593,In_2083,N_365);
or U1594 (N_1594,N_0,In_2023);
nor U1595 (N_1595,N_179,In_2628);
nand U1596 (N_1596,N_90,In_2938);
and U1597 (N_1597,N_802,In_2579);
nand U1598 (N_1598,In_1494,N_785);
or U1599 (N_1599,In_1540,N_322);
nor U1600 (N_1600,N_175,N_339);
xor U1601 (N_1601,In_1845,In_1420);
nand U1602 (N_1602,N_38,N_531);
nand U1603 (N_1603,In_2283,N_689);
nor U1604 (N_1604,In_2403,In_1398);
or U1605 (N_1605,N_160,N_566);
or U1606 (N_1606,N_435,N_454);
or U1607 (N_1607,N_558,In_1337);
nand U1608 (N_1608,N_598,N_960);
or U1609 (N_1609,N_415,In_1535);
xnor U1610 (N_1610,N_945,N_857);
nand U1611 (N_1611,In_2179,In_1642);
nor U1612 (N_1612,In_668,N_33);
nand U1613 (N_1613,N_268,In_2728);
or U1614 (N_1614,N_20,In_364);
and U1615 (N_1615,N_417,In_1948);
and U1616 (N_1616,In_1302,N_275);
and U1617 (N_1617,N_760,N_213);
nor U1618 (N_1618,N_767,N_868);
nand U1619 (N_1619,In_2100,N_436);
nor U1620 (N_1620,In_2887,N_384);
nand U1621 (N_1621,N_506,N_854);
or U1622 (N_1622,In_439,N_164);
or U1623 (N_1623,In_1428,N_653);
nor U1624 (N_1624,In_2399,N_471);
or U1625 (N_1625,In_10,N_342);
xor U1626 (N_1626,N_766,N_405);
and U1627 (N_1627,In_2867,N_968);
or U1628 (N_1628,In_2161,N_988);
nor U1629 (N_1629,N_769,N_443);
and U1630 (N_1630,In_145,N_244);
and U1631 (N_1631,N_197,N_284);
and U1632 (N_1632,N_266,N_112);
nand U1633 (N_1633,N_817,In_2866);
xor U1634 (N_1634,N_109,N_798);
xnor U1635 (N_1635,In_1832,N_816);
nand U1636 (N_1636,In_1596,In_183);
nand U1637 (N_1637,N_308,N_228);
nand U1638 (N_1638,In_606,In_2685);
xor U1639 (N_1639,N_758,In_1005);
and U1640 (N_1640,N_242,In_2815);
nor U1641 (N_1641,In_177,N_147);
nor U1642 (N_1642,In_777,In_1769);
nor U1643 (N_1643,N_456,N_97);
or U1644 (N_1644,N_621,In_2788);
xor U1645 (N_1645,In_1744,In_2276);
or U1646 (N_1646,In_2781,In_385);
nand U1647 (N_1647,N_491,In_1694);
xnor U1648 (N_1648,N_43,In_1574);
nor U1649 (N_1649,In_864,In_1239);
nor U1650 (N_1650,In_2151,In_2646);
nand U1651 (N_1651,N_56,In_1459);
nand U1652 (N_1652,N_656,N_404);
nor U1653 (N_1653,In_2400,In_2206);
nand U1654 (N_1654,In_1647,N_80);
or U1655 (N_1655,In_2385,In_2536);
or U1656 (N_1656,In_342,N_921);
nor U1657 (N_1657,N_154,N_604);
nand U1658 (N_1658,N_86,In_960);
nor U1659 (N_1659,N_812,N_397);
or U1660 (N_1660,N_975,In_1335);
nand U1661 (N_1661,N_819,N_140);
and U1662 (N_1662,In_514,In_1156);
and U1663 (N_1663,N_844,In_686);
nand U1664 (N_1664,N_855,N_122);
nand U1665 (N_1665,In_1285,In_131);
and U1666 (N_1666,N_690,N_628);
nor U1667 (N_1667,N_293,N_633);
nand U1668 (N_1668,In_418,N_345);
xnor U1669 (N_1669,In_2107,N_237);
or U1670 (N_1670,In_2207,N_372);
nor U1671 (N_1671,N_254,In_2216);
nand U1672 (N_1672,N_393,In_1083);
or U1673 (N_1673,In_1474,In_2588);
xor U1674 (N_1674,N_600,N_727);
and U1675 (N_1675,In_1735,N_350);
xnor U1676 (N_1676,N_248,N_852);
or U1677 (N_1677,N_411,N_4);
nor U1678 (N_1678,N_406,In_108);
xor U1679 (N_1679,In_2556,In_1987);
and U1680 (N_1680,N_281,N_996);
xor U1681 (N_1681,In_2707,In_1412);
nand U1682 (N_1682,N_716,N_778);
nor U1683 (N_1683,N_451,In_1355);
nor U1684 (N_1684,N_528,N_970);
nor U1685 (N_1685,N_984,N_253);
nand U1686 (N_1686,N_732,In_1196);
and U1687 (N_1687,N_37,In_2448);
or U1688 (N_1688,N_42,N_722);
and U1689 (N_1689,N_241,N_691);
nor U1690 (N_1690,In_375,N_302);
and U1691 (N_1691,In_134,N_418);
and U1692 (N_1692,In_2555,In_1850);
nor U1693 (N_1693,In_310,In_227);
nand U1694 (N_1694,In_2860,In_1058);
and U1695 (N_1695,In_1396,N_791);
nor U1696 (N_1696,In_2145,N_382);
and U1697 (N_1697,In_907,N_632);
nand U1698 (N_1698,N_6,In_379);
xnor U1699 (N_1699,N_710,In_599);
nor U1700 (N_1700,In_1696,N_432);
nor U1701 (N_1701,N_882,In_1947);
xor U1702 (N_1702,In_799,In_1275);
or U1703 (N_1703,N_740,N_169);
nor U1704 (N_1704,In_1389,N_831);
or U1705 (N_1705,In_641,In_1958);
or U1706 (N_1706,N_427,N_677);
nor U1707 (N_1707,N_651,In_509);
nand U1708 (N_1708,N_167,In_2243);
and U1709 (N_1709,In_2832,N_903);
or U1710 (N_1710,N_218,N_762);
xnor U1711 (N_1711,In_1544,N_768);
nand U1712 (N_1712,N_60,In_383);
and U1713 (N_1713,N_110,In_634);
or U1714 (N_1714,In_2457,N_12);
xnor U1715 (N_1715,N_586,In_840);
or U1716 (N_1716,In_2636,In_2093);
xnor U1717 (N_1717,N_733,N_77);
nand U1718 (N_1718,In_2757,N_117);
xor U1719 (N_1719,In_2849,N_666);
or U1720 (N_1720,N_499,N_870);
nor U1721 (N_1721,N_49,In_141);
nand U1722 (N_1722,N_679,In_1328);
and U1723 (N_1723,N_367,In_961);
or U1724 (N_1724,N_271,In_1006);
nor U1725 (N_1725,In_2552,N_85);
nand U1726 (N_1726,In_517,N_630);
nor U1727 (N_1727,In_441,In_96);
nor U1728 (N_1728,N_22,In_2751);
nor U1729 (N_1729,In_2561,In_449);
nor U1730 (N_1730,N_625,N_352);
nor U1731 (N_1731,In_2166,In_2305);
xnor U1732 (N_1732,In_1432,N_177);
nor U1733 (N_1733,In_1754,In_507);
xor U1734 (N_1734,In_2838,In_594);
nor U1735 (N_1735,In_2876,N_292);
nand U1736 (N_1736,In_951,N_116);
nand U1737 (N_1737,In_2212,In_2624);
or U1738 (N_1738,In_1008,N_226);
nand U1739 (N_1739,In_650,In_2570);
or U1740 (N_1740,In_2572,N_310);
nand U1741 (N_1741,N_467,N_358);
xnor U1742 (N_1742,In_2435,N_301);
xor U1743 (N_1743,N_448,In_71);
nor U1744 (N_1744,N_192,N_562);
nor U1745 (N_1745,N_991,In_434);
and U1746 (N_1746,N_94,In_1084);
xor U1747 (N_1747,In_328,N_386);
xnor U1748 (N_1748,In_930,N_961);
nand U1749 (N_1749,N_837,In_1512);
nor U1750 (N_1750,N_876,In_1679);
xor U1751 (N_1751,In_776,N_884);
and U1752 (N_1752,In_1470,N_949);
and U1753 (N_1753,N_835,In_161);
or U1754 (N_1754,N_62,In_1595);
nand U1755 (N_1755,N_239,N_925);
nor U1756 (N_1756,N_853,In_1746);
or U1757 (N_1757,In_1955,In_2803);
nand U1758 (N_1758,N_796,N_229);
or U1759 (N_1759,In_1149,N_856);
nor U1760 (N_1760,In_254,In_1117);
nand U1761 (N_1761,In_904,In_2330);
xnor U1762 (N_1762,In_511,N_545);
nor U1763 (N_1763,N_674,In_57);
nor U1764 (N_1764,In_713,In_795);
and U1765 (N_1765,N_538,In_2361);
nor U1766 (N_1766,In_1785,In_24);
nand U1767 (N_1767,N_231,In_2529);
nor U1768 (N_1768,N_764,In_1957);
nor U1769 (N_1769,N_887,N_307);
or U1770 (N_1770,In_351,In_1108);
nor U1771 (N_1771,N_75,N_641);
nor U1772 (N_1772,N_48,In_1894);
nor U1773 (N_1773,In_1114,N_428);
xor U1774 (N_1774,In_530,In_1147);
xor U1775 (N_1775,In_164,In_1567);
or U1776 (N_1776,In_2640,In_2547);
and U1777 (N_1777,In_1573,N_446);
nand U1778 (N_1778,In_403,N_76);
or U1779 (N_1779,N_83,N_702);
nor U1780 (N_1780,N_260,N_648);
xnor U1781 (N_1781,In_1374,N_743);
xor U1782 (N_1782,In_2537,N_320);
nand U1783 (N_1783,In_1288,In_648);
nor U1784 (N_1784,In_2031,N_442);
xnor U1785 (N_1785,In_1042,In_1662);
nor U1786 (N_1786,N_795,N_69);
or U1787 (N_1787,In_975,In_628);
nor U1788 (N_1788,N_423,In_2441);
or U1789 (N_1789,N_845,In_862);
nand U1790 (N_1790,N_480,N_492);
xor U1791 (N_1791,N_603,In_2029);
nand U1792 (N_1792,N_438,N_430);
or U1793 (N_1793,In_1041,N_917);
nor U1794 (N_1794,In_2560,N_347);
and U1795 (N_1795,In_1426,In_1465);
or U1796 (N_1796,In_1941,In_1161);
nand U1797 (N_1797,N_219,N_439);
nor U1798 (N_1798,In_1697,In_1430);
xnor U1799 (N_1799,In_2710,In_2551);
nor U1800 (N_1800,N_52,In_132);
nor U1801 (N_1801,In_575,N_619);
nor U1802 (N_1802,N_210,In_2520);
xor U1803 (N_1803,In_2295,N_915);
and U1804 (N_1804,In_1332,N_789);
xor U1805 (N_1805,In_1730,N_410);
nor U1806 (N_1806,In_139,N_663);
nor U1807 (N_1807,N_967,N_139);
xor U1808 (N_1808,N_533,N_36);
nand U1809 (N_1809,N_433,In_411);
nor U1810 (N_1810,N_773,In_999);
or U1811 (N_1811,N_182,N_942);
xor U1812 (N_1812,In_2222,N_194);
or U1813 (N_1813,In_466,In_353);
xnor U1814 (N_1814,In_2954,In_693);
or U1815 (N_1815,N_463,In_761);
and U1816 (N_1816,In_294,In_893);
and U1817 (N_1817,In_1766,In_1630);
nand U1818 (N_1818,N_647,In_563);
or U1819 (N_1819,In_453,In_2809);
or U1820 (N_1820,N_25,In_1577);
and U1821 (N_1821,N_990,N_576);
and U1822 (N_1822,N_104,In_1351);
and U1823 (N_1823,In_1844,In_2471);
nor U1824 (N_1824,In_1186,N_927);
or U1825 (N_1825,In_1617,In_1093);
nor U1826 (N_1826,N_526,N_905);
nor U1827 (N_1827,In_1753,In_1674);
xor U1828 (N_1828,In_336,N_252);
and U1829 (N_1829,In_1626,In_1056);
and U1830 (N_1830,In_2881,In_2188);
nand U1831 (N_1831,In_1452,In_1323);
nand U1832 (N_1832,N_263,In_1731);
nor U1833 (N_1833,In_1612,In_444);
or U1834 (N_1834,N_356,N_510);
nand U1835 (N_1835,N_517,In_2562);
nor U1836 (N_1836,N_639,N_444);
nand U1837 (N_1837,In_2422,In_1522);
nand U1838 (N_1838,N_594,N_623);
xor U1839 (N_1839,In_764,N_394);
xor U1840 (N_1840,In_1122,In_1124);
nor U1841 (N_1841,In_181,N_754);
nand U1842 (N_1842,In_2686,In_1602);
or U1843 (N_1843,In_356,In_769);
or U1844 (N_1844,N_387,In_1036);
nand U1845 (N_1845,N_88,N_431);
or U1846 (N_1846,N_832,N_230);
nor U1847 (N_1847,N_720,In_657);
nor U1848 (N_1848,In_1401,In_2253);
nor U1849 (N_1849,In_1800,In_2569);
nor U1850 (N_1850,In_2436,N_661);
or U1851 (N_1851,In_2217,In_1976);
or U1852 (N_1852,In_1930,N_143);
or U1853 (N_1853,In_2185,N_157);
xnor U1854 (N_1854,In_1319,N_306);
nor U1855 (N_1855,In_298,In_1825);
xnor U1856 (N_1856,N_453,N_267);
or U1857 (N_1857,N_924,N_609);
nand U1858 (N_1858,In_2365,N_998);
and U1859 (N_1859,In_996,In_830);
nand U1860 (N_1860,In_281,N_413);
or U1861 (N_1861,N_45,In_2550);
or U1862 (N_1862,N_458,In_1549);
xnor U1863 (N_1863,N_752,In_2121);
xnor U1864 (N_1864,In_649,In_2051);
nor U1865 (N_1865,N_580,In_2719);
nor U1866 (N_1866,N_288,In_1473);
and U1867 (N_1867,N_201,In_2979);
nor U1868 (N_1868,In_2657,N_223);
nor U1869 (N_1869,In_1317,N_67);
xnor U1870 (N_1870,In_1021,N_225);
xor U1871 (N_1871,In_1333,In_1592);
nand U1872 (N_1872,In_512,In_2592);
xor U1873 (N_1873,In_1854,N_299);
xor U1874 (N_1874,N_836,N_707);
nor U1875 (N_1875,In_544,In_1246);
and U1876 (N_1876,N_682,N_376);
nand U1877 (N_1877,In_213,N_66);
nand U1878 (N_1878,In_107,N_997);
nand U1879 (N_1879,N_739,In_2237);
and U1880 (N_1880,In_102,In_2460);
nand U1881 (N_1881,N_872,In_462);
and U1882 (N_1882,In_301,In_2381);
nand U1883 (N_1883,In_571,In_1797);
or U1884 (N_1884,N_671,In_1148);
and U1885 (N_1885,N_514,In_2694);
nand U1886 (N_1886,N_935,N_100);
and U1887 (N_1887,N_511,N_401);
xor U1888 (N_1888,N_460,In_1168);
or U1889 (N_1889,N_765,In_1699);
and U1890 (N_1890,In_1601,N_572);
xnor U1891 (N_1891,N_340,N_972);
nor U1892 (N_1892,In_1981,N_642);
nand U1893 (N_1893,In_1488,N_825);
and U1894 (N_1894,In_2382,In_330);
xor U1895 (N_1895,In_2541,N_741);
nand U1896 (N_1896,In_2315,In_495);
xnor U1897 (N_1897,In_246,N_772);
and U1898 (N_1898,N_146,In_1202);
or U1899 (N_1899,N_529,In_2992);
and U1900 (N_1900,N_19,In_2862);
or U1901 (N_1901,In_162,N_257);
or U1902 (N_1902,In_1681,In_2641);
or U1903 (N_1903,In_1242,In_1683);
or U1904 (N_1904,N_211,N_542);
and U1905 (N_1905,In_251,N_407);
nand U1906 (N_1906,N_962,In_1173);
nor U1907 (N_1907,N_508,N_932);
nor U1908 (N_1908,N_235,In_1062);
and U1909 (N_1909,N_227,N_602);
and U1910 (N_1910,N_698,In_937);
xor U1911 (N_1911,In_1216,In_2652);
nand U1912 (N_1912,In_2546,In_2674);
xor U1913 (N_1913,In_2252,In_2648);
nor U1914 (N_1914,N_166,N_412);
or U1915 (N_1915,N_640,In_1231);
nand U1916 (N_1916,N_258,In_2470);
or U1917 (N_1917,N_332,N_294);
xor U1918 (N_1918,In_2611,N_645);
and U1919 (N_1919,N_135,N_969);
nand U1920 (N_1920,N_8,In_2934);
or U1921 (N_1921,N_919,N_107);
nand U1922 (N_1922,N_859,N_314);
nand U1923 (N_1923,N_370,In_291);
or U1924 (N_1924,In_1773,In_1568);
and U1925 (N_1925,In_2925,N_665);
nand U1926 (N_1926,In_2055,N_701);
xor U1927 (N_1927,In_1354,In_2062);
xnor U1928 (N_1928,In_1227,N_388);
and U1929 (N_1929,N_21,N_498);
or U1930 (N_1930,N_864,In_1780);
nor U1931 (N_1931,In_282,In_1886);
and U1932 (N_1932,N_730,N_150);
and U1933 (N_1933,In_2596,In_2482);
and U1934 (N_1934,N_803,In_2453);
or U1935 (N_1935,In_839,In_2930);
or U1936 (N_1936,N_673,N_709);
nor U1937 (N_1937,In_1576,In_1303);
or U1938 (N_1938,In_823,N_841);
xnor U1939 (N_1939,In_2511,N_234);
nor U1940 (N_1940,N_151,In_1163);
xnor U1941 (N_1941,In_315,In_1134);
nor U1942 (N_1942,N_233,In_238);
or U1943 (N_1943,In_344,In_2702);
nor U1944 (N_1944,In_1944,N_951);
xnor U1945 (N_1945,N_662,N_539);
nor U1946 (N_1946,N_581,N_706);
or U1947 (N_1947,In_508,N_981);
or U1948 (N_1948,N_669,N_742);
nor U1949 (N_1949,N_596,In_1002);
xnor U1950 (N_1950,In_1125,In_1514);
nor U1951 (N_1951,N_948,N_814);
and U1952 (N_1952,In_2484,In_106);
nor U1953 (N_1953,In_399,In_1182);
and U1954 (N_1954,In_1019,In_2540);
or U1955 (N_1955,N_78,In_1234);
nor U1956 (N_1956,N_452,In_2479);
xnor U1957 (N_1957,N_744,In_2344);
and U1958 (N_1958,In_2447,In_2715);
nand U1959 (N_1959,In_1373,In_605);
xor U1960 (N_1960,In_696,N_123);
xor U1961 (N_1961,N_329,In_14);
nor U1962 (N_1962,N_535,In_1416);
or U1963 (N_1963,In_1692,In_2761);
xnor U1964 (N_1964,In_126,N_277);
or U1965 (N_1965,In_2928,N_797);
and U1966 (N_1966,N_99,In_1112);
and U1967 (N_1967,N_821,In_2519);
nor U1968 (N_1968,N_344,In_1477);
nor U1969 (N_1969,N_719,In_1745);
nor U1970 (N_1970,In_1555,N_280);
nor U1971 (N_1971,N_793,N_357);
xor U1972 (N_1972,In_993,N_425);
xnor U1973 (N_1973,N_588,N_131);
and U1974 (N_1974,N_330,N_351);
nor U1975 (N_1975,In_2752,N_891);
xnor U1976 (N_1976,In_360,N_947);
or U1977 (N_1977,N_103,N_521);
or U1978 (N_1978,N_622,N_303);
and U1979 (N_1979,N_834,In_798);
and U1980 (N_1980,N_934,N_377);
nor U1981 (N_1981,N_570,In_1762);
or U1982 (N_1982,N_833,In_1438);
nor U1983 (N_1983,In_185,In_702);
and U1984 (N_1984,In_1451,N_346);
nor U1985 (N_1985,N_846,N_348);
and U1986 (N_1986,In_1541,N_434);
and U1987 (N_1987,N_328,In_638);
nand U1988 (N_1988,N_543,N_476);
and U1989 (N_1989,N_667,In_2677);
nor U1990 (N_1990,N_402,In_1228);
nand U1991 (N_1991,In_2647,In_2337);
nor U1992 (N_1992,N_341,In_876);
and U1993 (N_1993,N_501,N_983);
nor U1994 (N_1994,In_2115,N_311);
nor U1995 (N_1995,N_191,N_512);
xnor U1996 (N_1996,In_2035,N_27);
xor U1997 (N_1997,In_912,N_274);
nand U1998 (N_1998,N_923,N_877);
nand U1999 (N_1999,N_568,N_858);
and U2000 (N_2000,N_1333,N_1328);
nand U2001 (N_2001,N_1065,N_1007);
nand U2002 (N_2002,N_1754,N_1508);
nor U2003 (N_2003,N_1512,N_1395);
and U2004 (N_2004,N_1952,N_1177);
xnor U2005 (N_2005,N_1751,N_1803);
nand U2006 (N_2006,N_1971,N_1975);
or U2007 (N_2007,N_1965,N_1604);
nor U2008 (N_2008,N_1516,N_1721);
nor U2009 (N_2009,N_1723,N_1213);
nor U2010 (N_2010,N_1098,N_1112);
or U2011 (N_2011,N_1635,N_1317);
xnor U2012 (N_2012,N_1248,N_1661);
nor U2013 (N_2013,N_1160,N_1392);
xor U2014 (N_2014,N_1294,N_1659);
xor U2015 (N_2015,N_1057,N_1077);
or U2016 (N_2016,N_1288,N_1176);
or U2017 (N_2017,N_1787,N_1851);
or U2018 (N_2018,N_1562,N_1470);
nor U2019 (N_2019,N_1329,N_1406);
or U2020 (N_2020,N_1890,N_1599);
and U2021 (N_2021,N_1886,N_1617);
or U2022 (N_2022,N_1338,N_1815);
xor U2023 (N_2023,N_1633,N_1427);
nand U2024 (N_2024,N_1296,N_1589);
and U2025 (N_2025,N_1367,N_1286);
and U2026 (N_2026,N_1842,N_1602);
nor U2027 (N_2027,N_1862,N_1685);
nor U2028 (N_2028,N_1527,N_1228);
nand U2029 (N_2029,N_1327,N_1033);
and U2030 (N_2030,N_1740,N_1504);
and U2031 (N_2031,N_1872,N_1239);
xor U2032 (N_2032,N_1896,N_1559);
nand U2033 (N_2033,N_1179,N_1678);
or U2034 (N_2034,N_1380,N_1986);
nand U2035 (N_2035,N_1823,N_1467);
and U2036 (N_2036,N_1864,N_1905);
nand U2037 (N_2037,N_1637,N_1558);
or U2038 (N_2038,N_1246,N_1394);
or U2039 (N_2039,N_1170,N_1901);
or U2040 (N_2040,N_1045,N_1163);
nand U2041 (N_2041,N_1197,N_1948);
and U2042 (N_2042,N_1199,N_1192);
or U2043 (N_2043,N_1004,N_1839);
nand U2044 (N_2044,N_1417,N_1686);
or U2045 (N_2045,N_1315,N_1924);
nand U2046 (N_2046,N_1486,N_1258);
xor U2047 (N_2047,N_1549,N_1505);
nand U2048 (N_2048,N_1591,N_1982);
nor U2049 (N_2049,N_1461,N_1001);
nor U2050 (N_2050,N_1365,N_1237);
nand U2051 (N_2051,N_1989,N_1411);
or U2052 (N_2052,N_1533,N_1820);
nor U2053 (N_2053,N_1696,N_1312);
and U2054 (N_2054,N_1645,N_1804);
and U2055 (N_2055,N_1072,N_1961);
xor U2056 (N_2056,N_1988,N_1852);
and U2057 (N_2057,N_1281,N_1233);
xor U2058 (N_2058,N_1929,N_1204);
nor U2059 (N_2059,N_1746,N_1026);
nand U2060 (N_2060,N_1238,N_1430);
xor U2061 (N_2061,N_1169,N_1959);
nand U2062 (N_2062,N_1222,N_1390);
nor U2063 (N_2063,N_1476,N_1621);
nor U2064 (N_2064,N_1916,N_1231);
or U2065 (N_2065,N_1172,N_1881);
nand U2066 (N_2066,N_1330,N_1434);
nor U2067 (N_2067,N_1437,N_1361);
nand U2068 (N_2068,N_1291,N_1831);
xor U2069 (N_2069,N_1818,N_1601);
nand U2070 (N_2070,N_1927,N_1784);
or U2071 (N_2071,N_1311,N_1126);
nand U2072 (N_2072,N_1907,N_1774);
and U2073 (N_2073,N_1290,N_1373);
nand U2074 (N_2074,N_1347,N_1770);
nor U2075 (N_2075,N_1344,N_1646);
and U2076 (N_2076,N_1984,N_1150);
nor U2077 (N_2077,N_1410,N_1154);
xnor U2078 (N_2078,N_1837,N_1008);
and U2079 (N_2079,N_1935,N_1107);
nand U2080 (N_2080,N_1183,N_1522);
or U2081 (N_2081,N_1594,N_1265);
xnor U2082 (N_2082,N_1649,N_1087);
nor U2083 (N_2083,N_1409,N_1489);
nand U2084 (N_2084,N_1651,N_1156);
nand U2085 (N_2085,N_1991,N_1980);
or U2086 (N_2086,N_1453,N_1071);
or U2087 (N_2087,N_1232,N_1300);
and U2088 (N_2088,N_1938,N_1456);
xnor U2089 (N_2089,N_1573,N_1490);
nor U2090 (N_2090,N_1268,N_1962);
nand U2091 (N_2091,N_1796,N_1114);
nand U2092 (N_2092,N_1700,N_1316);
or U2093 (N_2093,N_1543,N_1359);
nand U2094 (N_2094,N_1657,N_1349);
or U2095 (N_2095,N_1485,N_1612);
nor U2096 (N_2096,N_1352,N_1733);
and U2097 (N_2097,N_1526,N_1292);
xor U2098 (N_2098,N_1499,N_1790);
nor U2099 (N_2099,N_1495,N_1990);
or U2100 (N_2100,N_1750,N_1642);
xnor U2101 (N_2101,N_1285,N_1031);
or U2102 (N_2102,N_1581,N_1983);
nor U2103 (N_2103,N_1335,N_1734);
xnor U2104 (N_2104,N_1301,N_1236);
xnor U2105 (N_2105,N_1458,N_1575);
and U2106 (N_2106,N_1446,N_1964);
and U2107 (N_2107,N_1511,N_1542);
xnor U2108 (N_2108,N_1776,N_1429);
or U2109 (N_2109,N_1920,N_1608);
or U2110 (N_2110,N_1849,N_1203);
nor U2111 (N_2111,N_1000,N_1584);
xnor U2112 (N_2112,N_1110,N_1817);
or U2113 (N_2113,N_1977,N_1912);
nor U2114 (N_2114,N_1436,N_1550);
or U2115 (N_2115,N_1171,N_1838);
and U2116 (N_2116,N_1019,N_1752);
nor U2117 (N_2117,N_1123,N_1827);
nand U2118 (N_2118,N_1759,N_1951);
and U2119 (N_2119,N_1524,N_1810);
nand U2120 (N_2120,N_1566,N_1215);
or U2121 (N_2121,N_1547,N_1539);
nand U2122 (N_2122,N_1477,N_1652);
or U2123 (N_2123,N_1371,N_1819);
xnor U2124 (N_2124,N_1946,N_1133);
xor U2125 (N_2125,N_1287,N_1016);
and U2126 (N_2126,N_1155,N_1705);
nand U2127 (N_2127,N_1168,N_1162);
nand U2128 (N_2128,N_1643,N_1273);
nand U2129 (N_2129,N_1432,N_1888);
nand U2130 (N_2130,N_1710,N_1509);
and U2131 (N_2131,N_1707,N_1264);
xor U2132 (N_2132,N_1868,N_1899);
nor U2133 (N_2133,N_1857,N_1419);
xor U2134 (N_2134,N_1761,N_1363);
nor U2135 (N_2135,N_1497,N_1465);
nand U2136 (N_2136,N_1694,N_1947);
xor U2137 (N_2137,N_1995,N_1629);
and U2138 (N_2138,N_1501,N_1867);
or U2139 (N_2139,N_1537,N_1067);
nand U2140 (N_2140,N_1234,N_1611);
or U2141 (N_2141,N_1944,N_1431);
or U2142 (N_2142,N_1846,N_1459);
or U2143 (N_2143,N_1771,N_1978);
nor U2144 (N_2144,N_1998,N_1828);
xor U2145 (N_2145,N_1841,N_1496);
xnor U2146 (N_2146,N_1923,N_1407);
and U2147 (N_2147,N_1925,N_1731);
or U2148 (N_2148,N_1993,N_1348);
nand U2149 (N_2149,N_1873,N_1047);
nor U2150 (N_2150,N_1758,N_1243);
nand U2151 (N_2151,N_1424,N_1985);
nand U2152 (N_2152,N_1314,N_1362);
or U2153 (N_2153,N_1085,N_1387);
or U2154 (N_2154,N_1099,N_1095);
and U2155 (N_2155,N_1976,N_1120);
nand U2156 (N_2156,N_1519,N_1915);
xnor U2157 (N_2157,N_1032,N_1582);
or U2158 (N_2158,N_1051,N_1748);
nor U2159 (N_2159,N_1523,N_1598);
or U2160 (N_2160,N_1942,N_1850);
xor U2161 (N_2161,N_1339,N_1684);
and U2162 (N_2162,N_1229,N_1420);
or U2163 (N_2163,N_1403,N_1531);
or U2164 (N_2164,N_1809,N_1185);
nor U2165 (N_2165,N_1049,N_1251);
xnor U2166 (N_2166,N_1663,N_1536);
or U2167 (N_2167,N_1615,N_1950);
nand U2168 (N_2168,N_1021,N_1227);
and U2169 (N_2169,N_1833,N_1704);
and U2170 (N_2170,N_1195,N_1194);
nand U2171 (N_2171,N_1764,N_1435);
nor U2172 (N_2172,N_1464,N_1167);
nand U2173 (N_2173,N_1307,N_1036);
and U2174 (N_2174,N_1304,N_1037);
and U2175 (N_2175,N_1792,N_1520);
xnor U2176 (N_2176,N_1673,N_1449);
nor U2177 (N_2177,N_1015,N_1128);
and U2178 (N_2178,N_1366,N_1216);
xor U2179 (N_2179,N_1540,N_1046);
and U2180 (N_2180,N_1949,N_1917);
nand U2181 (N_2181,N_1321,N_1921);
and U2182 (N_2182,N_1058,N_1393);
or U2183 (N_2183,N_1463,N_1870);
nand U2184 (N_2184,N_1018,N_1957);
nor U2185 (N_2185,N_1207,N_1887);
xnor U2186 (N_2186,N_1368,N_1024);
nand U2187 (N_2187,N_1252,N_1681);
nor U2188 (N_2188,N_1571,N_1860);
xnor U2189 (N_2189,N_1040,N_1739);
nor U2190 (N_2190,N_1438,N_1386);
nor U2191 (N_2191,N_1009,N_1127);
or U2192 (N_2192,N_1175,N_1506);
nor U2193 (N_2193,N_1340,N_1412);
nor U2194 (N_2194,N_1389,N_1242);
xor U2195 (N_2195,N_1596,N_1667);
nand U2196 (N_2196,N_1877,N_1484);
nor U2197 (N_2197,N_1580,N_1726);
or U2198 (N_2198,N_1454,N_1769);
xor U2199 (N_2199,N_1378,N_1690);
nor U2200 (N_2200,N_1055,N_1963);
nand U2201 (N_2201,N_1401,N_1421);
xnor U2202 (N_2202,N_1426,N_1697);
or U2203 (N_2203,N_1360,N_1934);
and U2204 (N_2204,N_1910,N_1834);
and U2205 (N_2205,N_1966,N_1060);
or U2206 (N_2206,N_1277,N_1967);
xnor U2207 (N_2207,N_1457,N_1545);
or U2208 (N_2208,N_1137,N_1679);
or U2209 (N_2209,N_1786,N_1318);
xor U2210 (N_2210,N_1138,N_1174);
nand U2211 (N_2211,N_1274,N_1830);
xnor U2212 (N_2212,N_1093,N_1866);
or U2213 (N_2213,N_1498,N_1567);
xnor U2214 (N_2214,N_1152,N_1078);
nor U2215 (N_2215,N_1295,N_1541);
nand U2216 (N_2216,N_1554,N_1006);
nor U2217 (N_2217,N_1034,N_1379);
xor U2218 (N_2218,N_1655,N_1943);
or U2219 (N_2219,N_1848,N_1481);
and U2220 (N_2220,N_1630,N_1780);
xnor U2221 (N_2221,N_1255,N_1263);
xnor U2222 (N_2222,N_1262,N_1074);
nor U2223 (N_2223,N_1743,N_1219);
xor U2224 (N_2224,N_1483,N_1102);
xor U2225 (N_2225,N_1088,N_1022);
and U2226 (N_2226,N_1364,N_1147);
and U2227 (N_2227,N_1718,N_1121);
nor U2228 (N_2228,N_1119,N_1382);
nor U2229 (N_2229,N_1134,N_1092);
nand U2230 (N_2230,N_1105,N_1297);
xnor U2231 (N_2231,N_1418,N_1835);
nor U2232 (N_2232,N_1682,N_1149);
and U2233 (N_2233,N_1788,N_1135);
and U2234 (N_2234,N_1717,N_1053);
and U2235 (N_2235,N_1603,N_1182);
and U2236 (N_2236,N_1413,N_1441);
and U2237 (N_2237,N_1061,N_1094);
or U2238 (N_2238,N_1345,N_1666);
nor U2239 (N_2239,N_1038,N_1878);
and U2240 (N_2240,N_1342,N_1551);
xor U2241 (N_2241,N_1145,N_1936);
nor U2242 (N_2242,N_1257,N_1702);
and U2243 (N_2243,N_1709,N_1423);
and U2244 (N_2244,N_1115,N_1600);
nor U2245 (N_2245,N_1730,N_1958);
and U2246 (N_2246,N_1466,N_1513);
nor U2247 (N_2247,N_1798,N_1336);
xnor U2248 (N_2248,N_1178,N_1478);
or U2249 (N_2249,N_1735,N_1606);
or U2250 (N_2250,N_1668,N_1510);
and U2251 (N_2251,N_1108,N_1416);
nand U2252 (N_2252,N_1869,N_1131);
and U2253 (N_2253,N_1889,N_1043);
nor U2254 (N_2254,N_1535,N_1260);
or U2255 (N_2255,N_1309,N_1742);
nand U2256 (N_2256,N_1028,N_1703);
xor U2257 (N_2257,N_1578,N_1708);
and U2258 (N_2258,N_1247,N_1066);
or U2259 (N_2259,N_1030,N_1906);
nor U2260 (N_2260,N_1737,N_1829);
and U2261 (N_2261,N_1414,N_1142);
xnor U2262 (N_2262,N_1794,N_1245);
or U2263 (N_2263,N_1445,N_1002);
or U2264 (N_2264,N_1760,N_1272);
and U2265 (N_2265,N_1727,N_1041);
and U2266 (N_2266,N_1104,N_1276);
and U2267 (N_2267,N_1744,N_1560);
xor U2268 (N_2268,N_1398,N_1911);
nor U2269 (N_2269,N_1141,N_1614);
and U2270 (N_2270,N_1845,N_1230);
or U2271 (N_2271,N_1676,N_1202);
or U2272 (N_2272,N_1772,N_1455);
xor U2273 (N_2273,N_1100,N_1218);
nand U2274 (N_2274,N_1221,N_1408);
and U2275 (N_2275,N_1191,N_1278);
xnor U2276 (N_2276,N_1383,N_1641);
or U2277 (N_2277,N_1198,N_1208);
xor U2278 (N_2278,N_1415,N_1597);
xor U2279 (N_2279,N_1565,N_1903);
or U2280 (N_2280,N_1847,N_1672);
nand U2281 (N_2281,N_1013,N_1143);
and U2282 (N_2282,N_1576,N_1370);
or U2283 (N_2283,N_1940,N_1280);
or U2284 (N_2284,N_1855,N_1164);
or U2285 (N_2285,N_1157,N_1357);
nor U2286 (N_2286,N_1158,N_1812);
and U2287 (N_2287,N_1166,N_1671);
nand U2288 (N_2288,N_1206,N_1574);
and U2289 (N_2289,N_1048,N_1399);
or U2290 (N_2290,N_1201,N_1561);
nor U2291 (N_2291,N_1969,N_1588);
nor U2292 (N_2292,N_1900,N_1763);
xor U2293 (N_2293,N_1289,N_1186);
nor U2294 (N_2294,N_1473,N_1724);
or U2295 (N_2295,N_1332,N_1083);
and U2296 (N_2296,N_1824,N_1691);
nand U2297 (N_2297,N_1070,N_1665);
and U2298 (N_2298,N_1491,N_1425);
or U2299 (N_2299,N_1023,N_1184);
xnor U2300 (N_2300,N_1544,N_1973);
or U2301 (N_2301,N_1397,N_1354);
nand U2302 (N_2302,N_1548,N_1244);
xnor U2303 (N_2303,N_1711,N_1811);
nor U2304 (N_2304,N_1534,N_1235);
nand U2305 (N_2305,N_1306,N_1475);
nand U2306 (N_2306,N_1660,N_1625);
and U2307 (N_2307,N_1634,N_1586);
nor U2308 (N_2308,N_1358,N_1271);
or U2309 (N_2309,N_1909,N_1836);
and U2310 (N_2310,N_1714,N_1503);
and U2311 (N_2311,N_1897,N_1253);
nand U2312 (N_2312,N_1583,N_1091);
or U2313 (N_2313,N_1747,N_1644);
and U2314 (N_2314,N_1640,N_1632);
nor U2315 (N_2315,N_1139,N_1720);
xnor U2316 (N_2316,N_1122,N_1241);
nor U2317 (N_2317,N_1624,N_1482);
or U2318 (N_2318,N_1814,N_1778);
nand U2319 (N_2319,N_1933,N_1189);
xnor U2320 (N_2320,N_1609,N_1356);
nor U2321 (N_2321,N_1090,N_1715);
nor U2322 (N_2322,N_1775,N_1313);
nand U2323 (N_2323,N_1636,N_1487);
and U2324 (N_2324,N_1885,N_1595);
nand U2325 (N_2325,N_1689,N_1987);
nor U2326 (N_2326,N_1220,N_1181);
nand U2327 (N_2327,N_1736,N_1791);
nand U2328 (N_2328,N_1749,N_1293);
or U2329 (N_2329,N_1256,N_1444);
or U2330 (N_2330,N_1553,N_1658);
xor U2331 (N_2331,N_1259,N_1557);
nand U2332 (N_2332,N_1200,N_1391);
and U2333 (N_2333,N_1904,N_1626);
nor U2334 (N_2334,N_1518,N_1161);
nor U2335 (N_2335,N_1351,N_1261);
nor U2336 (N_2336,N_1479,N_1223);
nand U2337 (N_2337,N_1118,N_1728);
and U2338 (N_2338,N_1765,N_1068);
or U2339 (N_2339,N_1687,N_1337);
nand U2340 (N_2340,N_1546,N_1353);
nand U2341 (N_2341,N_1240,N_1664);
and U2342 (N_2342,N_1190,N_1572);
and U2343 (N_2343,N_1979,N_1879);
or U2344 (N_2344,N_1372,N_1593);
and U2345 (N_2345,N_1129,N_1768);
nor U2346 (N_2346,N_1494,N_1302);
or U2347 (N_2347,N_1439,N_1999);
or U2348 (N_2348,N_1310,N_1688);
or U2349 (N_2349,N_1500,N_1692);
and U2350 (N_2350,N_1738,N_1517);
or U2351 (N_2351,N_1876,N_1622);
and U2352 (N_2352,N_1981,N_1492);
and U2353 (N_2353,N_1620,N_1822);
nand U2354 (N_2354,N_1875,N_1422);
xnor U2355 (N_2355,N_1111,N_1474);
nor U2356 (N_2356,N_1180,N_1767);
nor U2357 (N_2357,N_1521,N_1140);
and U2358 (N_2358,N_1400,N_1270);
nor U2359 (N_2359,N_1913,N_1056);
nand U2360 (N_2360,N_1832,N_1701);
xnor U2361 (N_2361,N_1662,N_1376);
nor U2362 (N_2362,N_1713,N_1225);
or U2363 (N_2363,N_1613,N_1610);
and U2364 (N_2364,N_1196,N_1159);
xor U2365 (N_2365,N_1954,N_1472);
nor U2366 (N_2366,N_1428,N_1050);
nand U2367 (N_2367,N_1089,N_1618);
or U2368 (N_2368,N_1283,N_1590);
xor U2369 (N_2369,N_1029,N_1891);
nor U2370 (N_2370,N_1103,N_1529);
xor U2371 (N_2371,N_1334,N_1840);
xnor U2372 (N_2372,N_1797,N_1569);
xor U2373 (N_2373,N_1874,N_1005);
nor U2374 (N_2374,N_1442,N_1585);
or U2375 (N_2375,N_1165,N_1806);
or U2376 (N_2376,N_1974,N_1124);
xnor U2377 (N_2377,N_1081,N_1109);
and U2378 (N_2378,N_1440,N_1343);
nand U2379 (N_2379,N_1777,N_1076);
and U2380 (N_2380,N_1282,N_1217);
nand U2381 (N_2381,N_1863,N_1698);
nand U2382 (N_2382,N_1807,N_1173);
or U2383 (N_2383,N_1062,N_1308);
nor U2384 (N_2384,N_1011,N_1355);
or U2385 (N_2385,N_1385,N_1579);
or U2386 (N_2386,N_1319,N_1299);
xnor U2387 (N_2387,N_1941,N_1254);
and U2388 (N_2388,N_1577,N_1502);
nand U2389 (N_2389,N_1059,N_1706);
xnor U2390 (N_2390,N_1779,N_1939);
or U2391 (N_2391,N_1930,N_1211);
xnor U2392 (N_2392,N_1825,N_1269);
nand U2393 (N_2393,N_1012,N_1331);
nand U2394 (N_2394,N_1802,N_1783);
xor U2395 (N_2395,N_1858,N_1799);
nor U2396 (N_2396,N_1782,N_1205);
nor U2397 (N_2397,N_1451,N_1918);
nor U2398 (N_2398,N_1042,N_1097);
nor U2399 (N_2399,N_1493,N_1374);
xnor U2400 (N_2400,N_1801,N_1994);
and U2401 (N_2401,N_1341,N_1719);
xor U2402 (N_2402,N_1322,N_1674);
or U2403 (N_2403,N_1369,N_1405);
nor U2404 (N_2404,N_1805,N_1448);
and U2405 (N_2405,N_1388,N_1861);
nand U2406 (N_2406,N_1082,N_1532);
or U2407 (N_2407,N_1214,N_1017);
nand U2408 (N_2408,N_1249,N_1997);
xnor U2409 (N_2409,N_1928,N_1267);
xor U2410 (N_2410,N_1396,N_1992);
nor U2411 (N_2411,N_1808,N_1895);
nand U2412 (N_2412,N_1117,N_1151);
or U2413 (N_2413,N_1148,N_1755);
nor U2414 (N_2414,N_1039,N_1628);
xor U2415 (N_2415,N_1756,N_1266);
xnor U2416 (N_2416,N_1669,N_1027);
or U2417 (N_2417,N_1616,N_1722);
xnor U2418 (N_2418,N_1781,N_1003);
and U2419 (N_2419,N_1144,N_1773);
xor U2420 (N_2420,N_1069,N_1677);
nor U2421 (N_2421,N_1712,N_1813);
nand U2422 (N_2422,N_1648,N_1044);
or U2423 (N_2423,N_1865,N_1675);
xor U2424 (N_2424,N_1462,N_1224);
and U2425 (N_2425,N_1153,N_1384);
or U2426 (N_2426,N_1639,N_1250);
nor U2427 (N_2427,N_1741,N_1279);
and U2428 (N_2428,N_1654,N_1695);
and U2429 (N_2429,N_1563,N_1745);
and U2430 (N_2430,N_1080,N_1960);
and U2431 (N_2431,N_1132,N_1193);
nor U2432 (N_2432,N_1883,N_1375);
xor U2433 (N_2433,N_1035,N_1101);
and U2434 (N_2434,N_1766,N_1647);
xnor U2435 (N_2435,N_1086,N_1785);
nand U2436 (N_2436,N_1871,N_1212);
nor U2437 (N_2437,N_1471,N_1996);
nor U2438 (N_2438,N_1893,N_1075);
nor U2439 (N_2439,N_1753,N_1795);
nand U2440 (N_2440,N_1079,N_1680);
nand U2441 (N_2441,N_1507,N_1209);
xor U2442 (N_2442,N_1125,N_1324);
nand U2443 (N_2443,N_1693,N_1762);
nor U2444 (N_2444,N_1063,N_1619);
nand U2445 (N_2445,N_1631,N_1844);
or U2446 (N_2446,N_1096,N_1605);
or U2447 (N_2447,N_1488,N_1210);
and U2448 (N_2448,N_1607,N_1298);
or U2449 (N_2449,N_1020,N_1638);
nand U2450 (N_2450,N_1014,N_1381);
xor U2451 (N_2451,N_1025,N_1010);
xnor U2452 (N_2452,N_1650,N_1443);
nor U2453 (N_2453,N_1656,N_1555);
and U2454 (N_2454,N_1908,N_1880);
nor U2455 (N_2455,N_1084,N_1926);
nand U2456 (N_2456,N_1130,N_1113);
nand U2457 (N_2457,N_1816,N_1623);
and U2458 (N_2458,N_1305,N_1460);
or U2459 (N_2459,N_1882,N_1528);
nand U2460 (N_2460,N_1116,N_1793);
and U2461 (N_2461,N_1968,N_1146);
and U2462 (N_2462,N_1568,N_1725);
and U2463 (N_2463,N_1323,N_1325);
and U2464 (N_2464,N_1956,N_1932);
nor U2465 (N_2465,N_1592,N_1450);
nor U2466 (N_2466,N_1469,N_1530);
xor U2467 (N_2467,N_1226,N_1902);
xor U2468 (N_2468,N_1729,N_1757);
or U2469 (N_2469,N_1919,N_1188);
nand U2470 (N_2470,N_1570,N_1187);
nand U2471 (N_2471,N_1884,N_1922);
xnor U2472 (N_2472,N_1073,N_1955);
nand U2473 (N_2473,N_1052,N_1350);
and U2474 (N_2474,N_1136,N_1538);
and U2475 (N_2475,N_1821,N_1843);
and U2476 (N_2476,N_1859,N_1402);
nand U2477 (N_2477,N_1468,N_1800);
xor U2478 (N_2478,N_1856,N_1433);
nor U2479 (N_2479,N_1064,N_1826);
nand U2480 (N_2480,N_1452,N_1447);
or U2481 (N_2481,N_1683,N_1346);
nor U2482 (N_2482,N_1404,N_1854);
nor U2483 (N_2483,N_1627,N_1892);
xnor U2484 (N_2484,N_1480,N_1894);
nand U2485 (N_2485,N_1898,N_1552);
and U2486 (N_2486,N_1275,N_1970);
xor U2487 (N_2487,N_1320,N_1525);
xnor U2488 (N_2488,N_1945,N_1914);
or U2489 (N_2489,N_1699,N_1514);
xnor U2490 (N_2490,N_1564,N_1789);
xor U2491 (N_2491,N_1953,N_1931);
xor U2492 (N_2492,N_1054,N_1972);
nor U2493 (N_2493,N_1587,N_1326);
nand U2494 (N_2494,N_1303,N_1716);
xor U2495 (N_2495,N_1670,N_1556);
and U2496 (N_2496,N_1937,N_1853);
or U2497 (N_2497,N_1653,N_1732);
or U2498 (N_2498,N_1284,N_1377);
and U2499 (N_2499,N_1106,N_1515);
or U2500 (N_2500,N_1543,N_1430);
and U2501 (N_2501,N_1070,N_1579);
nor U2502 (N_2502,N_1859,N_1561);
xnor U2503 (N_2503,N_1374,N_1497);
or U2504 (N_2504,N_1050,N_1613);
xnor U2505 (N_2505,N_1429,N_1092);
or U2506 (N_2506,N_1593,N_1955);
nor U2507 (N_2507,N_1709,N_1133);
nand U2508 (N_2508,N_1581,N_1964);
nand U2509 (N_2509,N_1418,N_1337);
or U2510 (N_2510,N_1524,N_1486);
nand U2511 (N_2511,N_1286,N_1882);
nand U2512 (N_2512,N_1899,N_1460);
and U2513 (N_2513,N_1429,N_1382);
xor U2514 (N_2514,N_1148,N_1768);
nand U2515 (N_2515,N_1749,N_1997);
nand U2516 (N_2516,N_1016,N_1819);
nand U2517 (N_2517,N_1420,N_1300);
xor U2518 (N_2518,N_1470,N_1362);
xor U2519 (N_2519,N_1644,N_1274);
and U2520 (N_2520,N_1014,N_1983);
nand U2521 (N_2521,N_1235,N_1943);
nor U2522 (N_2522,N_1707,N_1080);
nand U2523 (N_2523,N_1504,N_1013);
nor U2524 (N_2524,N_1308,N_1858);
and U2525 (N_2525,N_1112,N_1772);
nor U2526 (N_2526,N_1438,N_1832);
nor U2527 (N_2527,N_1819,N_1289);
or U2528 (N_2528,N_1434,N_1753);
nor U2529 (N_2529,N_1271,N_1221);
nand U2530 (N_2530,N_1865,N_1399);
nand U2531 (N_2531,N_1560,N_1970);
nor U2532 (N_2532,N_1704,N_1433);
nand U2533 (N_2533,N_1738,N_1628);
and U2534 (N_2534,N_1675,N_1159);
and U2535 (N_2535,N_1650,N_1876);
or U2536 (N_2536,N_1459,N_1641);
or U2537 (N_2537,N_1490,N_1672);
and U2538 (N_2538,N_1158,N_1464);
nand U2539 (N_2539,N_1287,N_1517);
nand U2540 (N_2540,N_1094,N_1405);
and U2541 (N_2541,N_1855,N_1257);
nand U2542 (N_2542,N_1724,N_1830);
xnor U2543 (N_2543,N_1388,N_1384);
and U2544 (N_2544,N_1752,N_1193);
xnor U2545 (N_2545,N_1873,N_1654);
nor U2546 (N_2546,N_1992,N_1761);
nand U2547 (N_2547,N_1894,N_1818);
or U2548 (N_2548,N_1577,N_1547);
nand U2549 (N_2549,N_1288,N_1810);
nand U2550 (N_2550,N_1108,N_1115);
and U2551 (N_2551,N_1494,N_1493);
nand U2552 (N_2552,N_1997,N_1476);
nor U2553 (N_2553,N_1303,N_1684);
and U2554 (N_2554,N_1480,N_1421);
xnor U2555 (N_2555,N_1576,N_1654);
nand U2556 (N_2556,N_1959,N_1554);
xor U2557 (N_2557,N_1443,N_1400);
xnor U2558 (N_2558,N_1924,N_1367);
or U2559 (N_2559,N_1651,N_1266);
nor U2560 (N_2560,N_1000,N_1052);
xor U2561 (N_2561,N_1648,N_1050);
or U2562 (N_2562,N_1074,N_1918);
nand U2563 (N_2563,N_1978,N_1293);
xor U2564 (N_2564,N_1250,N_1784);
nor U2565 (N_2565,N_1051,N_1052);
nor U2566 (N_2566,N_1939,N_1094);
nand U2567 (N_2567,N_1562,N_1026);
or U2568 (N_2568,N_1643,N_1947);
xnor U2569 (N_2569,N_1896,N_1546);
xnor U2570 (N_2570,N_1998,N_1902);
xnor U2571 (N_2571,N_1829,N_1607);
xor U2572 (N_2572,N_1091,N_1796);
xor U2573 (N_2573,N_1313,N_1562);
and U2574 (N_2574,N_1878,N_1972);
or U2575 (N_2575,N_1572,N_1226);
nor U2576 (N_2576,N_1980,N_1981);
nand U2577 (N_2577,N_1008,N_1809);
nand U2578 (N_2578,N_1304,N_1389);
xnor U2579 (N_2579,N_1435,N_1885);
nor U2580 (N_2580,N_1883,N_1770);
nand U2581 (N_2581,N_1305,N_1645);
xnor U2582 (N_2582,N_1016,N_1292);
nor U2583 (N_2583,N_1278,N_1006);
or U2584 (N_2584,N_1009,N_1864);
or U2585 (N_2585,N_1855,N_1743);
or U2586 (N_2586,N_1861,N_1618);
or U2587 (N_2587,N_1109,N_1315);
nand U2588 (N_2588,N_1984,N_1661);
or U2589 (N_2589,N_1364,N_1389);
or U2590 (N_2590,N_1055,N_1906);
nand U2591 (N_2591,N_1900,N_1784);
xor U2592 (N_2592,N_1772,N_1798);
nor U2593 (N_2593,N_1715,N_1814);
xor U2594 (N_2594,N_1995,N_1921);
nor U2595 (N_2595,N_1231,N_1305);
xor U2596 (N_2596,N_1189,N_1077);
nor U2597 (N_2597,N_1383,N_1170);
nand U2598 (N_2598,N_1267,N_1706);
nand U2599 (N_2599,N_1287,N_1456);
xor U2600 (N_2600,N_1053,N_1725);
nand U2601 (N_2601,N_1759,N_1130);
nor U2602 (N_2602,N_1201,N_1158);
xor U2603 (N_2603,N_1568,N_1575);
xnor U2604 (N_2604,N_1147,N_1320);
and U2605 (N_2605,N_1733,N_1686);
xor U2606 (N_2606,N_1403,N_1156);
xor U2607 (N_2607,N_1869,N_1397);
xor U2608 (N_2608,N_1329,N_1541);
nand U2609 (N_2609,N_1185,N_1041);
xor U2610 (N_2610,N_1769,N_1169);
xor U2611 (N_2611,N_1593,N_1444);
nor U2612 (N_2612,N_1347,N_1413);
and U2613 (N_2613,N_1469,N_1369);
nand U2614 (N_2614,N_1037,N_1230);
and U2615 (N_2615,N_1417,N_1960);
or U2616 (N_2616,N_1657,N_1754);
or U2617 (N_2617,N_1095,N_1380);
nand U2618 (N_2618,N_1353,N_1907);
or U2619 (N_2619,N_1297,N_1157);
nand U2620 (N_2620,N_1006,N_1726);
or U2621 (N_2621,N_1416,N_1444);
xnor U2622 (N_2622,N_1277,N_1024);
xor U2623 (N_2623,N_1455,N_1520);
nand U2624 (N_2624,N_1528,N_1112);
or U2625 (N_2625,N_1399,N_1024);
or U2626 (N_2626,N_1262,N_1828);
or U2627 (N_2627,N_1853,N_1813);
xor U2628 (N_2628,N_1584,N_1670);
xor U2629 (N_2629,N_1943,N_1301);
xor U2630 (N_2630,N_1263,N_1100);
and U2631 (N_2631,N_1207,N_1369);
nor U2632 (N_2632,N_1727,N_1708);
nor U2633 (N_2633,N_1363,N_1477);
or U2634 (N_2634,N_1647,N_1868);
xnor U2635 (N_2635,N_1814,N_1713);
nor U2636 (N_2636,N_1392,N_1088);
or U2637 (N_2637,N_1073,N_1210);
nand U2638 (N_2638,N_1695,N_1184);
and U2639 (N_2639,N_1783,N_1527);
xnor U2640 (N_2640,N_1345,N_1708);
nand U2641 (N_2641,N_1690,N_1276);
xnor U2642 (N_2642,N_1041,N_1087);
nor U2643 (N_2643,N_1541,N_1369);
nor U2644 (N_2644,N_1400,N_1895);
nand U2645 (N_2645,N_1000,N_1332);
nand U2646 (N_2646,N_1709,N_1061);
nand U2647 (N_2647,N_1978,N_1259);
xnor U2648 (N_2648,N_1270,N_1358);
xnor U2649 (N_2649,N_1915,N_1505);
xor U2650 (N_2650,N_1720,N_1287);
nor U2651 (N_2651,N_1664,N_1277);
or U2652 (N_2652,N_1981,N_1827);
nand U2653 (N_2653,N_1999,N_1867);
nand U2654 (N_2654,N_1487,N_1114);
xor U2655 (N_2655,N_1245,N_1972);
or U2656 (N_2656,N_1370,N_1495);
nand U2657 (N_2657,N_1640,N_1526);
nand U2658 (N_2658,N_1200,N_1103);
xor U2659 (N_2659,N_1085,N_1179);
and U2660 (N_2660,N_1836,N_1824);
nor U2661 (N_2661,N_1795,N_1083);
nor U2662 (N_2662,N_1658,N_1995);
and U2663 (N_2663,N_1472,N_1318);
nand U2664 (N_2664,N_1201,N_1527);
nor U2665 (N_2665,N_1987,N_1320);
and U2666 (N_2666,N_1879,N_1858);
xor U2667 (N_2667,N_1900,N_1660);
or U2668 (N_2668,N_1566,N_1773);
or U2669 (N_2669,N_1471,N_1424);
nand U2670 (N_2670,N_1113,N_1191);
xor U2671 (N_2671,N_1618,N_1187);
or U2672 (N_2672,N_1137,N_1788);
and U2673 (N_2673,N_1415,N_1108);
nand U2674 (N_2674,N_1075,N_1130);
nor U2675 (N_2675,N_1596,N_1735);
and U2676 (N_2676,N_1560,N_1909);
or U2677 (N_2677,N_1754,N_1704);
or U2678 (N_2678,N_1624,N_1784);
nor U2679 (N_2679,N_1514,N_1659);
nand U2680 (N_2680,N_1194,N_1846);
nor U2681 (N_2681,N_1840,N_1060);
and U2682 (N_2682,N_1437,N_1770);
and U2683 (N_2683,N_1658,N_1940);
or U2684 (N_2684,N_1053,N_1592);
xnor U2685 (N_2685,N_1667,N_1195);
xor U2686 (N_2686,N_1642,N_1853);
nand U2687 (N_2687,N_1371,N_1327);
xor U2688 (N_2688,N_1715,N_1899);
or U2689 (N_2689,N_1252,N_1780);
xor U2690 (N_2690,N_1567,N_1725);
and U2691 (N_2691,N_1699,N_1134);
nor U2692 (N_2692,N_1690,N_1543);
xor U2693 (N_2693,N_1487,N_1285);
nand U2694 (N_2694,N_1768,N_1067);
and U2695 (N_2695,N_1886,N_1510);
nor U2696 (N_2696,N_1003,N_1883);
xor U2697 (N_2697,N_1198,N_1881);
and U2698 (N_2698,N_1756,N_1187);
and U2699 (N_2699,N_1376,N_1417);
and U2700 (N_2700,N_1819,N_1342);
nand U2701 (N_2701,N_1925,N_1958);
or U2702 (N_2702,N_1640,N_1080);
nand U2703 (N_2703,N_1456,N_1633);
nor U2704 (N_2704,N_1153,N_1734);
xnor U2705 (N_2705,N_1475,N_1852);
nor U2706 (N_2706,N_1042,N_1852);
xor U2707 (N_2707,N_1478,N_1687);
or U2708 (N_2708,N_1397,N_1324);
and U2709 (N_2709,N_1948,N_1085);
xor U2710 (N_2710,N_1822,N_1089);
and U2711 (N_2711,N_1319,N_1506);
xor U2712 (N_2712,N_1506,N_1546);
xnor U2713 (N_2713,N_1797,N_1007);
nor U2714 (N_2714,N_1861,N_1479);
xnor U2715 (N_2715,N_1870,N_1320);
nor U2716 (N_2716,N_1442,N_1366);
xor U2717 (N_2717,N_1206,N_1146);
nand U2718 (N_2718,N_1697,N_1114);
xor U2719 (N_2719,N_1880,N_1998);
or U2720 (N_2720,N_1764,N_1773);
or U2721 (N_2721,N_1968,N_1349);
and U2722 (N_2722,N_1623,N_1964);
and U2723 (N_2723,N_1254,N_1378);
nor U2724 (N_2724,N_1780,N_1193);
xnor U2725 (N_2725,N_1469,N_1382);
xor U2726 (N_2726,N_1559,N_1332);
nor U2727 (N_2727,N_1277,N_1209);
xor U2728 (N_2728,N_1742,N_1335);
nor U2729 (N_2729,N_1556,N_1579);
and U2730 (N_2730,N_1862,N_1972);
nand U2731 (N_2731,N_1052,N_1202);
and U2732 (N_2732,N_1563,N_1539);
nor U2733 (N_2733,N_1974,N_1049);
or U2734 (N_2734,N_1273,N_1333);
nor U2735 (N_2735,N_1580,N_1276);
nand U2736 (N_2736,N_1231,N_1918);
xor U2737 (N_2737,N_1628,N_1225);
nand U2738 (N_2738,N_1320,N_1010);
and U2739 (N_2739,N_1335,N_1768);
or U2740 (N_2740,N_1632,N_1392);
or U2741 (N_2741,N_1283,N_1524);
nor U2742 (N_2742,N_1086,N_1412);
xor U2743 (N_2743,N_1829,N_1593);
and U2744 (N_2744,N_1559,N_1656);
xor U2745 (N_2745,N_1330,N_1566);
and U2746 (N_2746,N_1404,N_1358);
and U2747 (N_2747,N_1998,N_1467);
and U2748 (N_2748,N_1188,N_1754);
and U2749 (N_2749,N_1274,N_1913);
or U2750 (N_2750,N_1082,N_1159);
and U2751 (N_2751,N_1995,N_1100);
and U2752 (N_2752,N_1419,N_1988);
nor U2753 (N_2753,N_1669,N_1500);
or U2754 (N_2754,N_1710,N_1439);
xor U2755 (N_2755,N_1094,N_1654);
or U2756 (N_2756,N_1106,N_1712);
nand U2757 (N_2757,N_1672,N_1642);
xnor U2758 (N_2758,N_1604,N_1556);
or U2759 (N_2759,N_1131,N_1302);
or U2760 (N_2760,N_1931,N_1772);
nand U2761 (N_2761,N_1336,N_1960);
xor U2762 (N_2762,N_1824,N_1438);
nor U2763 (N_2763,N_1130,N_1503);
xnor U2764 (N_2764,N_1517,N_1280);
nand U2765 (N_2765,N_1064,N_1012);
nor U2766 (N_2766,N_1423,N_1653);
nor U2767 (N_2767,N_1663,N_1733);
nor U2768 (N_2768,N_1221,N_1765);
nand U2769 (N_2769,N_1484,N_1587);
or U2770 (N_2770,N_1793,N_1743);
and U2771 (N_2771,N_1718,N_1217);
nand U2772 (N_2772,N_1520,N_1131);
or U2773 (N_2773,N_1859,N_1289);
xnor U2774 (N_2774,N_1903,N_1825);
and U2775 (N_2775,N_1253,N_1638);
and U2776 (N_2776,N_1294,N_1074);
and U2777 (N_2777,N_1970,N_1094);
and U2778 (N_2778,N_1390,N_1423);
nand U2779 (N_2779,N_1143,N_1825);
and U2780 (N_2780,N_1551,N_1724);
xor U2781 (N_2781,N_1131,N_1455);
and U2782 (N_2782,N_1204,N_1918);
or U2783 (N_2783,N_1069,N_1833);
or U2784 (N_2784,N_1783,N_1041);
nor U2785 (N_2785,N_1614,N_1547);
xor U2786 (N_2786,N_1304,N_1537);
or U2787 (N_2787,N_1315,N_1748);
xor U2788 (N_2788,N_1495,N_1729);
nor U2789 (N_2789,N_1142,N_1937);
nand U2790 (N_2790,N_1879,N_1697);
nand U2791 (N_2791,N_1083,N_1653);
xor U2792 (N_2792,N_1729,N_1475);
and U2793 (N_2793,N_1833,N_1129);
and U2794 (N_2794,N_1859,N_1747);
and U2795 (N_2795,N_1442,N_1581);
and U2796 (N_2796,N_1574,N_1244);
and U2797 (N_2797,N_1428,N_1522);
and U2798 (N_2798,N_1953,N_1876);
nor U2799 (N_2799,N_1238,N_1982);
or U2800 (N_2800,N_1969,N_1052);
or U2801 (N_2801,N_1478,N_1966);
nor U2802 (N_2802,N_1094,N_1003);
xnor U2803 (N_2803,N_1796,N_1270);
nor U2804 (N_2804,N_1546,N_1428);
or U2805 (N_2805,N_1204,N_1269);
xnor U2806 (N_2806,N_1008,N_1953);
xnor U2807 (N_2807,N_1508,N_1622);
and U2808 (N_2808,N_1555,N_1373);
or U2809 (N_2809,N_1347,N_1820);
nand U2810 (N_2810,N_1784,N_1421);
nor U2811 (N_2811,N_1531,N_1591);
or U2812 (N_2812,N_1608,N_1473);
nand U2813 (N_2813,N_1713,N_1419);
and U2814 (N_2814,N_1683,N_1534);
or U2815 (N_2815,N_1305,N_1475);
or U2816 (N_2816,N_1931,N_1891);
nor U2817 (N_2817,N_1523,N_1199);
xor U2818 (N_2818,N_1391,N_1432);
nand U2819 (N_2819,N_1333,N_1260);
nand U2820 (N_2820,N_1980,N_1946);
or U2821 (N_2821,N_1593,N_1390);
nor U2822 (N_2822,N_1903,N_1215);
or U2823 (N_2823,N_1319,N_1085);
and U2824 (N_2824,N_1535,N_1741);
nor U2825 (N_2825,N_1411,N_1228);
or U2826 (N_2826,N_1851,N_1583);
nand U2827 (N_2827,N_1062,N_1233);
nor U2828 (N_2828,N_1456,N_1263);
nand U2829 (N_2829,N_1193,N_1532);
xnor U2830 (N_2830,N_1240,N_1908);
xor U2831 (N_2831,N_1913,N_1074);
nand U2832 (N_2832,N_1001,N_1663);
nand U2833 (N_2833,N_1578,N_1212);
nand U2834 (N_2834,N_1004,N_1418);
nor U2835 (N_2835,N_1169,N_1817);
nand U2836 (N_2836,N_1276,N_1795);
nor U2837 (N_2837,N_1321,N_1619);
xnor U2838 (N_2838,N_1129,N_1899);
or U2839 (N_2839,N_1328,N_1615);
or U2840 (N_2840,N_1841,N_1447);
and U2841 (N_2841,N_1897,N_1387);
or U2842 (N_2842,N_1863,N_1800);
or U2843 (N_2843,N_1447,N_1140);
nand U2844 (N_2844,N_1979,N_1448);
nand U2845 (N_2845,N_1442,N_1044);
and U2846 (N_2846,N_1776,N_1525);
nor U2847 (N_2847,N_1405,N_1353);
nand U2848 (N_2848,N_1841,N_1222);
xnor U2849 (N_2849,N_1864,N_1162);
and U2850 (N_2850,N_1588,N_1121);
or U2851 (N_2851,N_1018,N_1881);
or U2852 (N_2852,N_1684,N_1034);
and U2853 (N_2853,N_1821,N_1134);
or U2854 (N_2854,N_1139,N_1011);
or U2855 (N_2855,N_1581,N_1955);
xnor U2856 (N_2856,N_1350,N_1746);
and U2857 (N_2857,N_1644,N_1026);
nor U2858 (N_2858,N_1884,N_1255);
and U2859 (N_2859,N_1898,N_1799);
and U2860 (N_2860,N_1836,N_1026);
nor U2861 (N_2861,N_1574,N_1129);
nor U2862 (N_2862,N_1795,N_1698);
or U2863 (N_2863,N_1375,N_1013);
and U2864 (N_2864,N_1246,N_1688);
xnor U2865 (N_2865,N_1838,N_1903);
nor U2866 (N_2866,N_1973,N_1846);
nand U2867 (N_2867,N_1970,N_1668);
or U2868 (N_2868,N_1222,N_1697);
nor U2869 (N_2869,N_1983,N_1650);
xor U2870 (N_2870,N_1132,N_1029);
or U2871 (N_2871,N_1170,N_1473);
nand U2872 (N_2872,N_1477,N_1200);
and U2873 (N_2873,N_1832,N_1483);
xor U2874 (N_2874,N_1601,N_1519);
nand U2875 (N_2875,N_1997,N_1833);
xnor U2876 (N_2876,N_1692,N_1353);
xor U2877 (N_2877,N_1084,N_1722);
nor U2878 (N_2878,N_1710,N_1065);
and U2879 (N_2879,N_1138,N_1486);
nand U2880 (N_2880,N_1899,N_1524);
nand U2881 (N_2881,N_1045,N_1528);
or U2882 (N_2882,N_1432,N_1505);
nand U2883 (N_2883,N_1269,N_1202);
nor U2884 (N_2884,N_1089,N_1639);
and U2885 (N_2885,N_1764,N_1674);
and U2886 (N_2886,N_1637,N_1051);
nand U2887 (N_2887,N_1043,N_1080);
xor U2888 (N_2888,N_1614,N_1442);
nor U2889 (N_2889,N_1924,N_1316);
xor U2890 (N_2890,N_1258,N_1729);
nor U2891 (N_2891,N_1082,N_1999);
nand U2892 (N_2892,N_1124,N_1178);
and U2893 (N_2893,N_1050,N_1989);
and U2894 (N_2894,N_1766,N_1500);
nor U2895 (N_2895,N_1531,N_1698);
xnor U2896 (N_2896,N_1594,N_1707);
nand U2897 (N_2897,N_1448,N_1812);
nor U2898 (N_2898,N_1282,N_1320);
nor U2899 (N_2899,N_1079,N_1265);
xor U2900 (N_2900,N_1545,N_1692);
nor U2901 (N_2901,N_1447,N_1634);
or U2902 (N_2902,N_1509,N_1034);
nor U2903 (N_2903,N_1008,N_1534);
and U2904 (N_2904,N_1495,N_1170);
xor U2905 (N_2905,N_1120,N_1336);
or U2906 (N_2906,N_1472,N_1240);
and U2907 (N_2907,N_1854,N_1485);
xnor U2908 (N_2908,N_1471,N_1949);
or U2909 (N_2909,N_1760,N_1134);
nor U2910 (N_2910,N_1457,N_1175);
or U2911 (N_2911,N_1884,N_1464);
and U2912 (N_2912,N_1678,N_1416);
nor U2913 (N_2913,N_1317,N_1321);
nand U2914 (N_2914,N_1158,N_1281);
xor U2915 (N_2915,N_1985,N_1626);
or U2916 (N_2916,N_1307,N_1530);
nand U2917 (N_2917,N_1093,N_1359);
and U2918 (N_2918,N_1328,N_1422);
nand U2919 (N_2919,N_1423,N_1026);
nand U2920 (N_2920,N_1687,N_1767);
xnor U2921 (N_2921,N_1232,N_1589);
or U2922 (N_2922,N_1466,N_1773);
nand U2923 (N_2923,N_1924,N_1466);
xor U2924 (N_2924,N_1615,N_1162);
and U2925 (N_2925,N_1358,N_1963);
nor U2926 (N_2926,N_1888,N_1412);
or U2927 (N_2927,N_1992,N_1091);
and U2928 (N_2928,N_1473,N_1872);
nor U2929 (N_2929,N_1831,N_1247);
nand U2930 (N_2930,N_1835,N_1461);
xnor U2931 (N_2931,N_1216,N_1521);
and U2932 (N_2932,N_1588,N_1165);
or U2933 (N_2933,N_1063,N_1580);
or U2934 (N_2934,N_1881,N_1341);
and U2935 (N_2935,N_1899,N_1882);
nand U2936 (N_2936,N_1052,N_1483);
xnor U2937 (N_2937,N_1776,N_1586);
xnor U2938 (N_2938,N_1593,N_1402);
and U2939 (N_2939,N_1922,N_1166);
or U2940 (N_2940,N_1913,N_1997);
xnor U2941 (N_2941,N_1254,N_1363);
nand U2942 (N_2942,N_1661,N_1507);
xor U2943 (N_2943,N_1500,N_1103);
or U2944 (N_2944,N_1824,N_1359);
nand U2945 (N_2945,N_1865,N_1683);
xor U2946 (N_2946,N_1580,N_1298);
nand U2947 (N_2947,N_1279,N_1228);
or U2948 (N_2948,N_1308,N_1362);
nor U2949 (N_2949,N_1956,N_1054);
nor U2950 (N_2950,N_1299,N_1496);
nand U2951 (N_2951,N_1666,N_1530);
and U2952 (N_2952,N_1428,N_1794);
nor U2953 (N_2953,N_1801,N_1618);
nor U2954 (N_2954,N_1680,N_1026);
nor U2955 (N_2955,N_1410,N_1596);
nand U2956 (N_2956,N_1977,N_1367);
and U2957 (N_2957,N_1237,N_1355);
nand U2958 (N_2958,N_1822,N_1159);
xnor U2959 (N_2959,N_1876,N_1868);
and U2960 (N_2960,N_1406,N_1558);
and U2961 (N_2961,N_1211,N_1157);
nand U2962 (N_2962,N_1868,N_1889);
xnor U2963 (N_2963,N_1614,N_1645);
nand U2964 (N_2964,N_1281,N_1588);
nand U2965 (N_2965,N_1520,N_1278);
and U2966 (N_2966,N_1505,N_1734);
nand U2967 (N_2967,N_1157,N_1627);
or U2968 (N_2968,N_1644,N_1580);
or U2969 (N_2969,N_1535,N_1373);
nor U2970 (N_2970,N_1059,N_1795);
nor U2971 (N_2971,N_1892,N_1029);
or U2972 (N_2972,N_1640,N_1989);
nand U2973 (N_2973,N_1670,N_1866);
xor U2974 (N_2974,N_1306,N_1222);
or U2975 (N_2975,N_1290,N_1690);
or U2976 (N_2976,N_1953,N_1989);
or U2977 (N_2977,N_1065,N_1362);
or U2978 (N_2978,N_1284,N_1409);
xor U2979 (N_2979,N_1156,N_1883);
nand U2980 (N_2980,N_1373,N_1983);
nor U2981 (N_2981,N_1859,N_1663);
nor U2982 (N_2982,N_1705,N_1596);
nand U2983 (N_2983,N_1961,N_1358);
and U2984 (N_2984,N_1340,N_1848);
or U2985 (N_2985,N_1558,N_1785);
or U2986 (N_2986,N_1674,N_1431);
nand U2987 (N_2987,N_1420,N_1035);
nor U2988 (N_2988,N_1324,N_1323);
nor U2989 (N_2989,N_1546,N_1624);
and U2990 (N_2990,N_1141,N_1193);
nand U2991 (N_2991,N_1977,N_1162);
xnor U2992 (N_2992,N_1900,N_1681);
xor U2993 (N_2993,N_1742,N_1665);
or U2994 (N_2994,N_1441,N_1088);
nor U2995 (N_2995,N_1803,N_1655);
nand U2996 (N_2996,N_1622,N_1150);
or U2997 (N_2997,N_1595,N_1582);
and U2998 (N_2998,N_1938,N_1473);
or U2999 (N_2999,N_1901,N_1157);
xor U3000 (N_3000,N_2480,N_2517);
xnor U3001 (N_3001,N_2213,N_2221);
or U3002 (N_3002,N_2216,N_2981);
xor U3003 (N_3003,N_2312,N_2044);
xor U3004 (N_3004,N_2073,N_2561);
nand U3005 (N_3005,N_2944,N_2635);
nor U3006 (N_3006,N_2626,N_2406);
nand U3007 (N_3007,N_2449,N_2690);
xnor U3008 (N_3008,N_2060,N_2243);
or U3009 (N_3009,N_2979,N_2323);
and U3010 (N_3010,N_2651,N_2859);
and U3011 (N_3011,N_2028,N_2346);
or U3012 (N_3012,N_2585,N_2089);
xnor U3013 (N_3013,N_2744,N_2278);
or U3014 (N_3014,N_2362,N_2371);
or U3015 (N_3015,N_2775,N_2550);
xnor U3016 (N_3016,N_2311,N_2258);
nor U3017 (N_3017,N_2265,N_2074);
or U3018 (N_3018,N_2069,N_2732);
nor U3019 (N_3019,N_2932,N_2765);
xnor U3020 (N_3020,N_2888,N_2931);
and U3021 (N_3021,N_2023,N_2794);
nand U3022 (N_3022,N_2835,N_2576);
nor U3023 (N_3023,N_2219,N_2798);
nand U3024 (N_3024,N_2985,N_2112);
xor U3025 (N_3025,N_2827,N_2137);
or U3026 (N_3026,N_2793,N_2830);
nor U3027 (N_3027,N_2256,N_2053);
nand U3028 (N_3028,N_2152,N_2908);
and U3029 (N_3029,N_2810,N_2352);
and U3030 (N_3030,N_2735,N_2361);
and U3031 (N_3031,N_2686,N_2366);
and U3032 (N_3032,N_2970,N_2270);
and U3033 (N_3033,N_2994,N_2763);
xnor U3034 (N_3034,N_2729,N_2722);
or U3035 (N_3035,N_2092,N_2159);
nand U3036 (N_3036,N_2710,N_2544);
xor U3037 (N_3037,N_2506,N_2405);
nor U3038 (N_3038,N_2679,N_2495);
nand U3039 (N_3039,N_2855,N_2780);
nor U3040 (N_3040,N_2754,N_2695);
or U3041 (N_3041,N_2160,N_2937);
nand U3042 (N_3042,N_2683,N_2781);
or U3043 (N_3043,N_2663,N_2698);
xor U3044 (N_3044,N_2554,N_2719);
nor U3045 (N_3045,N_2815,N_2747);
nor U3046 (N_3046,N_2641,N_2012);
xnor U3047 (N_3047,N_2849,N_2422);
xor U3048 (N_3048,N_2887,N_2100);
or U3049 (N_3049,N_2058,N_2464);
and U3050 (N_3050,N_2388,N_2612);
and U3051 (N_3051,N_2475,N_2674);
and U3052 (N_3052,N_2106,N_2753);
or U3053 (N_3053,N_2501,N_2512);
nand U3054 (N_3054,N_2656,N_2942);
xor U3055 (N_3055,N_2518,N_2260);
xor U3056 (N_3056,N_2974,N_2108);
nor U3057 (N_3057,N_2597,N_2685);
and U3058 (N_3058,N_2766,N_2930);
or U3059 (N_3059,N_2086,N_2141);
nand U3060 (N_3060,N_2867,N_2292);
xnor U3061 (N_3061,N_2630,N_2463);
xnor U3062 (N_3062,N_2139,N_2914);
or U3063 (N_3063,N_2315,N_2750);
and U3064 (N_3064,N_2938,N_2555);
nor U3065 (N_3065,N_2749,N_2273);
nor U3066 (N_3066,N_2886,N_2821);
or U3067 (N_3067,N_2493,N_2148);
and U3068 (N_3068,N_2466,N_2569);
nand U3069 (N_3069,N_2600,N_2770);
nor U3070 (N_3070,N_2134,N_2474);
nand U3071 (N_3071,N_2647,N_2397);
xor U3072 (N_3072,N_2892,N_2689);
xor U3073 (N_3073,N_2521,N_2197);
and U3074 (N_3074,N_2844,N_2584);
nor U3075 (N_3075,N_2056,N_2824);
nor U3076 (N_3076,N_2812,N_2688);
xor U3077 (N_3077,N_2935,N_2170);
and U3078 (N_3078,N_2805,N_2856);
nand U3079 (N_3079,N_2013,N_2364);
and U3080 (N_3080,N_2715,N_2707);
xnor U3081 (N_3081,N_2603,N_2165);
nand U3082 (N_3082,N_2154,N_2210);
or U3083 (N_3083,N_2933,N_2175);
and U3084 (N_3084,N_2387,N_2649);
nor U3085 (N_3085,N_2087,N_2860);
and U3086 (N_3086,N_2136,N_2401);
nand U3087 (N_3087,N_2054,N_2229);
and U3088 (N_3088,N_2296,N_2540);
xnor U3089 (N_3089,N_2333,N_2613);
nor U3090 (N_3090,N_2426,N_2653);
xor U3091 (N_3091,N_2113,N_2486);
nand U3092 (N_3092,N_2669,N_2797);
xor U3093 (N_3093,N_2990,N_2709);
or U3094 (N_3094,N_2995,N_2923);
nor U3095 (N_3095,N_2564,N_2018);
xnor U3096 (N_3096,N_2907,N_2394);
and U3097 (N_3097,N_2169,N_2993);
nand U3098 (N_3098,N_2965,N_2926);
or U3099 (N_3099,N_2356,N_2648);
and U3100 (N_3100,N_2778,N_2402);
nor U3101 (N_3101,N_2180,N_2945);
nand U3102 (N_3102,N_2264,N_2309);
nor U3103 (N_3103,N_2999,N_2878);
or U3104 (N_3104,N_2488,N_2768);
and U3105 (N_3105,N_2740,N_2232);
xnor U3106 (N_3106,N_2654,N_2730);
nor U3107 (N_3107,N_2642,N_2290);
nand U3108 (N_3108,N_2204,N_2800);
and U3109 (N_3109,N_2407,N_2657);
and U3110 (N_3110,N_2948,N_2115);
xor U3111 (N_3111,N_2759,N_2183);
xnor U3112 (N_3112,N_2072,N_2530);
and U3113 (N_3113,N_2701,N_2850);
or U3114 (N_3114,N_2070,N_2173);
or U3115 (N_3115,N_2380,N_2306);
nand U3116 (N_3116,N_2791,N_2234);
and U3117 (N_3117,N_2271,N_2155);
and U3118 (N_3118,N_2419,N_2249);
nor U3119 (N_3119,N_2334,N_2218);
xnor U3120 (N_3120,N_2902,N_2116);
nand U3121 (N_3121,N_2446,N_2095);
nand U3122 (N_3122,N_2531,N_2904);
and U3123 (N_3123,N_2414,N_2840);
nand U3124 (N_3124,N_2400,N_2124);
nand U3125 (N_3125,N_2558,N_2454);
and U3126 (N_3126,N_2457,N_2529);
nor U3127 (N_3127,N_2969,N_2525);
or U3128 (N_3128,N_2967,N_2130);
xor U3129 (N_3129,N_2345,N_2910);
and U3130 (N_3130,N_2806,N_2037);
or U3131 (N_3131,N_2462,N_2043);
nand U3132 (N_3132,N_2602,N_2897);
and U3133 (N_3133,N_2538,N_2739);
nand U3134 (N_3134,N_2151,N_2682);
nand U3135 (N_3135,N_2348,N_2245);
and U3136 (N_3136,N_2332,N_2548);
xor U3137 (N_3137,N_2833,N_2848);
nand U3138 (N_3138,N_2138,N_2186);
and U3139 (N_3139,N_2237,N_2450);
or U3140 (N_3140,N_2675,N_2541);
nor U3141 (N_3141,N_2145,N_2403);
xor U3142 (N_3142,N_2829,N_2741);
nor U3143 (N_3143,N_2713,N_2971);
and U3144 (N_3144,N_2723,N_2898);
nor U3145 (N_3145,N_2852,N_2565);
nand U3146 (N_3146,N_2605,N_2157);
xor U3147 (N_3147,N_2034,N_2963);
xnor U3148 (N_3148,N_2560,N_2968);
or U3149 (N_3149,N_2890,N_2542);
or U3150 (N_3150,N_2357,N_2660);
and U3151 (N_3151,N_2527,N_2283);
and U3152 (N_3152,N_2076,N_2881);
xor U3153 (N_3153,N_2838,N_2000);
nand U3154 (N_3154,N_2021,N_2964);
xor U3155 (N_3155,N_2006,N_2767);
xnor U3156 (N_3156,N_2301,N_2962);
nand U3157 (N_3157,N_2697,N_2681);
and U3158 (N_3158,N_2310,N_2487);
nand U3159 (N_3159,N_2230,N_2862);
or U3160 (N_3160,N_2075,N_2212);
xor U3161 (N_3161,N_2639,N_2389);
xnor U3162 (N_3162,N_2953,N_2004);
xor U3163 (N_3163,N_2568,N_2293);
or U3164 (N_3164,N_2061,N_2619);
or U3165 (N_3165,N_2992,N_2955);
nor U3166 (N_3166,N_2019,N_2874);
and U3167 (N_3167,N_2007,N_2240);
nor U3168 (N_3168,N_2551,N_2431);
and U3169 (N_3169,N_2813,N_2279);
or U3170 (N_3170,N_2643,N_2658);
nor U3171 (N_3171,N_2442,N_2014);
and U3172 (N_3172,N_2254,N_2065);
or U3173 (N_3173,N_2746,N_2539);
nor U3174 (N_3174,N_2233,N_2420);
xnor U3175 (N_3175,N_2295,N_2826);
nand U3176 (N_3176,N_2338,N_2764);
and U3177 (N_3177,N_2928,N_2691);
nand U3178 (N_3178,N_2502,N_2771);
or U3179 (N_3179,N_2176,N_2001);
nor U3180 (N_3180,N_2973,N_2404);
nand U3181 (N_3181,N_2563,N_2864);
nor U3182 (N_3182,N_2132,N_2118);
nand U3183 (N_3183,N_2321,N_2150);
xor U3184 (N_3184,N_2328,N_2194);
nor U3185 (N_3185,N_2960,N_2496);
nand U3186 (N_3186,N_2049,N_2324);
nand U3187 (N_3187,N_2876,N_2756);
xor U3188 (N_3188,N_2162,N_2303);
nand U3189 (N_3189,N_2659,N_2248);
nor U3190 (N_3190,N_2574,N_2085);
nor U3191 (N_3191,N_2339,N_2869);
xnor U3192 (N_3192,N_2733,N_2179);
or U3193 (N_3193,N_2029,N_2453);
nand U3194 (N_3194,N_2040,N_2515);
nor U3195 (N_3195,N_2678,N_2492);
nor U3196 (N_3196,N_2809,N_2164);
nor U3197 (N_3197,N_2742,N_2490);
nand U3198 (N_3198,N_2077,N_2621);
and U3199 (N_3199,N_2680,N_2559);
or U3200 (N_3200,N_2351,N_2436);
or U3201 (N_3201,N_2451,N_2611);
nor U3202 (N_3202,N_2002,N_2636);
and U3203 (N_3203,N_2090,N_2415);
nor U3204 (N_3204,N_2631,N_2430);
and U3205 (N_3205,N_2267,N_2988);
nor U3206 (N_3206,N_2788,N_2819);
and U3207 (N_3207,N_2599,N_2836);
xnor U3208 (N_3208,N_2783,N_2491);
xor U3209 (N_3209,N_2877,N_2432);
xnor U3210 (N_3210,N_2208,N_2235);
and U3211 (N_3211,N_2593,N_2620);
or U3212 (N_3212,N_2711,N_2121);
nor U3213 (N_3213,N_2822,N_2662);
xor U3214 (N_3214,N_2182,N_2577);
and U3215 (N_3215,N_2314,N_2712);
nand U3216 (N_3216,N_2718,N_2231);
and U3217 (N_3217,N_2223,N_2755);
and U3218 (N_3218,N_2467,N_2322);
nor U3219 (N_3219,N_2858,N_2851);
and U3220 (N_3220,N_2027,N_2832);
nor U3221 (N_3221,N_2247,N_2181);
nand U3222 (N_3222,N_2059,N_2365);
and U3223 (N_3223,N_2342,N_2769);
nor U3224 (N_3224,N_2468,N_2667);
or U3225 (N_3225,N_2299,N_2983);
or U3226 (N_3226,N_2262,N_2284);
and U3227 (N_3227,N_2943,N_2408);
nand U3228 (N_3228,N_2634,N_2255);
nor U3229 (N_3229,N_2105,N_2784);
nand U3230 (N_3230,N_2716,N_2571);
nor U3231 (N_3231,N_2655,N_2596);
nand U3232 (N_3232,N_2785,N_2670);
or U3233 (N_3233,N_2929,N_2610);
nand U3234 (N_3234,N_2702,N_2135);
nand U3235 (N_3235,N_2880,N_2978);
nor U3236 (N_3236,N_2395,N_2045);
and U3237 (N_3237,N_2276,N_2016);
nor U3238 (N_3238,N_2714,N_2146);
nor U3239 (N_3239,N_2291,N_2423);
nand U3240 (N_3240,N_2140,N_2251);
nand U3241 (N_3241,N_2185,N_2174);
and U3242 (N_3242,N_2035,N_2206);
or U3243 (N_3243,N_2583,N_2048);
and U3244 (N_3244,N_2259,N_2355);
nand U3245 (N_3245,N_2298,N_2047);
xor U3246 (N_3246,N_2804,N_2640);
or U3247 (N_3247,N_2624,N_2760);
nand U3248 (N_3248,N_2782,N_2817);
nand U3249 (N_3249,N_2369,N_2752);
nor U3250 (N_3250,N_2687,N_2665);
nor U3251 (N_3251,N_2101,N_2834);
or U3252 (N_3252,N_2861,N_2927);
or U3253 (N_3253,N_2586,N_2854);
nand U3254 (N_3254,N_2917,N_2269);
and U3255 (N_3255,N_2511,N_2343);
nor U3256 (N_3256,N_2646,N_2863);
and U3257 (N_3257,N_2424,N_2104);
and U3258 (N_3258,N_2093,N_2313);
nor U3259 (N_3259,N_2190,N_2725);
or U3260 (N_3260,N_2872,N_2478);
nor U3261 (N_3261,N_2336,N_2396);
and U3262 (N_3262,N_2096,N_2133);
nor U3263 (N_3263,N_2811,N_2524);
and U3264 (N_3264,N_2383,N_2222);
nor U3265 (N_3265,N_2853,N_2025);
xor U3266 (N_3266,N_2772,N_2590);
and U3267 (N_3267,N_2814,N_2520);
and U3268 (N_3268,N_2470,N_2281);
nor U3269 (N_3269,N_2637,N_2316);
and U3270 (N_3270,N_2870,N_2084);
nand U3271 (N_3271,N_2894,N_2294);
nor U3272 (N_3272,N_2773,N_2057);
xnor U3273 (N_3273,N_2982,N_2010);
and U3274 (N_3274,N_2196,N_2706);
or U3275 (N_3275,N_2526,N_2425);
and U3276 (N_3276,N_2215,N_2111);
nor U3277 (N_3277,N_2980,N_2418);
and U3278 (N_3278,N_2708,N_2147);
nor U3279 (N_3279,N_2330,N_2916);
nand U3280 (N_3280,N_2445,N_2055);
or U3281 (N_3281,N_2846,N_2557);
and U3282 (N_3282,N_2042,N_2918);
nand U3283 (N_3283,N_2297,N_2427);
nor U3284 (N_3284,N_2158,N_2909);
nor U3285 (N_3285,N_2666,N_2919);
and U3286 (N_3286,N_2537,N_2319);
nor U3287 (N_3287,N_2376,N_2608);
xnor U3288 (N_3288,N_2738,N_2110);
nor U3289 (N_3289,N_2347,N_2692);
nand U3290 (N_3290,N_2941,N_2721);
xor U3291 (N_3291,N_2604,N_2149);
or U3292 (N_3292,N_2274,N_2694);
or U3293 (N_3293,N_2922,N_2318);
nand U3294 (N_3294,N_2308,N_2409);
nor U3295 (N_3295,N_2091,N_2616);
nor U3296 (N_3296,N_2789,N_2609);
and U3297 (N_3297,N_2252,N_2633);
nor U3298 (N_3298,N_2421,N_2949);
xnor U3299 (N_3299,N_2882,N_2167);
nand U3300 (N_3300,N_2924,N_2915);
nor U3301 (N_3301,N_2083,N_2220);
nor U3302 (N_3302,N_2504,N_2912);
and U3303 (N_3303,N_2331,N_2370);
and U3304 (N_3304,N_2349,N_2329);
xor U3305 (N_3305,N_2358,N_2300);
nand U3306 (N_3306,N_2381,N_2020);
nand U3307 (N_3307,N_2547,N_2239);
nor U3308 (N_3308,N_2022,N_2489);
or U3309 (N_3309,N_2051,N_2372);
nor U3310 (N_3310,N_2959,N_2579);
xor U3311 (N_3311,N_2940,N_2438);
and U3312 (N_3312,N_2071,N_2307);
and U3313 (N_3313,N_2614,N_2455);
nand U3314 (N_3314,N_2726,N_2039);
or U3315 (N_3315,N_2050,N_2479);
and U3316 (N_3316,N_2500,N_2211);
nor U3317 (N_3317,N_2808,N_2606);
or U3318 (N_3318,N_2866,N_2736);
and U3319 (N_3319,N_2956,N_2327);
and U3320 (N_3320,N_2360,N_2607);
xnor U3321 (N_3321,N_2905,N_2523);
nand U3322 (N_3322,N_2842,N_2828);
nand U3323 (N_3323,N_2818,N_2857);
nand U3324 (N_3324,N_2198,N_2337);
nand U3325 (N_3325,N_2661,N_2598);
nor U3326 (N_3326,N_2119,N_2217);
nand U3327 (N_3327,N_2494,N_2393);
or U3328 (N_3328,N_2505,N_2499);
and U3329 (N_3329,N_2673,N_2939);
and U3330 (N_3330,N_2335,N_2777);
and U3331 (N_3331,N_2030,N_2471);
xor U3332 (N_3332,N_2566,N_2519);
nor U3333 (N_3333,N_2015,N_2799);
or U3334 (N_3334,N_2459,N_2289);
nor U3335 (N_3335,N_2831,N_2129);
nor U3336 (N_3336,N_2473,N_2079);
or U3337 (N_3337,N_2437,N_2458);
nand U3338 (N_3338,N_2434,N_2758);
nor U3339 (N_3339,N_2201,N_2282);
and U3340 (N_3340,N_2224,N_2353);
and U3341 (N_3341,N_2776,N_2865);
xnor U3342 (N_3342,N_2997,N_2052);
xnor U3343 (N_3343,N_2200,N_2911);
nand U3344 (N_3344,N_2556,N_2128);
or U3345 (N_3345,N_2628,N_2192);
nor U3346 (N_3346,N_2417,N_2570);
xor U3347 (N_3347,N_2873,N_2677);
or U3348 (N_3348,N_2203,N_2627);
or U3349 (N_3349,N_2934,N_2761);
or U3350 (N_3350,N_2737,N_2026);
nor U3351 (N_3351,N_2325,N_2460);
or U3352 (N_3352,N_2594,N_2913);
nand U3353 (N_3353,N_2549,N_2632);
nor U3354 (N_3354,N_2341,N_2543);
xor U3355 (N_3355,N_2241,N_2131);
xnor U3356 (N_3356,N_2625,N_2433);
or U3357 (N_3357,N_2266,N_2246);
and U3358 (N_3358,N_2891,N_2484);
xor U3359 (N_3359,N_2003,N_2127);
and U3360 (N_3360,N_2705,N_2503);
or U3361 (N_3361,N_2081,N_2900);
nor U3362 (N_3362,N_2986,N_2591);
nor U3363 (N_3363,N_2317,N_2645);
or U3364 (N_3364,N_2906,N_2976);
xnor U3365 (N_3365,N_2845,N_2950);
nand U3366 (N_3366,N_2385,N_2429);
nand U3367 (N_3367,N_2534,N_2064);
and U3368 (N_3368,N_2440,N_2903);
xor U3369 (N_3369,N_2748,N_2589);
or U3370 (N_3370,N_2285,N_2801);
or U3371 (N_3371,N_2202,N_2277);
or U3372 (N_3372,N_2178,N_2373);
nand U3373 (N_3373,N_2552,N_2580);
or U3374 (N_3374,N_2510,N_2062);
and U3375 (N_3375,N_2899,N_2122);
and U3376 (N_3376,N_2172,N_2481);
and U3377 (N_3377,N_2103,N_2617);
or U3378 (N_3378,N_2823,N_2644);
and U3379 (N_3379,N_2416,N_2261);
xnor U3380 (N_3380,N_2263,N_2195);
nor U3381 (N_3381,N_2671,N_2731);
xor U3382 (N_3382,N_2946,N_2787);
and U3383 (N_3383,N_2024,N_2126);
or U3384 (N_3384,N_2441,N_2033);
nor U3385 (N_3385,N_2011,N_2790);
and U3386 (N_3386,N_2546,N_2413);
and U3387 (N_3387,N_2461,N_2144);
nor U3388 (N_3388,N_2412,N_2536);
xor U3389 (N_3389,N_2228,N_2895);
nor U3390 (N_3390,N_2984,N_2236);
xnor U3391 (N_3391,N_2280,N_2359);
nand U3392 (N_3392,N_2774,N_2036);
nor U3393 (N_3393,N_2989,N_2883);
and U3394 (N_3394,N_2483,N_2123);
nor U3395 (N_3395,N_2428,N_2304);
nand U3396 (N_3396,N_2120,N_2038);
nor U3397 (N_3397,N_2171,N_2996);
nand U3398 (N_3398,N_2094,N_2893);
xor U3399 (N_3399,N_2166,N_2302);
nor U3400 (N_3400,N_2498,N_2595);
nor U3401 (N_3401,N_2080,N_2226);
or U3402 (N_3402,N_2693,N_2622);
or U3403 (N_3403,N_2977,N_2199);
nand U3404 (N_3404,N_2391,N_2672);
nand U3405 (N_3405,N_2879,N_2320);
nor U3406 (N_3406,N_2063,N_2390);
and U3407 (N_3407,N_2456,N_2684);
nand U3408 (N_3408,N_2786,N_2191);
nand U3409 (N_3409,N_2485,N_2975);
nor U3410 (N_3410,N_2088,N_2469);
nor U3411 (N_3411,N_2507,N_2532);
xor U3412 (N_3412,N_2802,N_2444);
xnor U3413 (N_3413,N_2472,N_2399);
and U3414 (N_3414,N_2272,N_2363);
nand U3415 (N_3415,N_2209,N_2188);
nand U3416 (N_3416,N_2947,N_2901);
or U3417 (N_3417,N_2920,N_2623);
xor U3418 (N_3418,N_2588,N_2578);
xnor U3419 (N_3419,N_2008,N_2109);
or U3420 (N_3420,N_2587,N_2477);
or U3421 (N_3421,N_2189,N_2751);
xnor U3422 (N_3422,N_2921,N_2871);
or U3423 (N_3423,N_2275,N_2615);
nand U3424 (N_3424,N_2884,N_2326);
xnor U3425 (N_3425,N_2187,N_2286);
or U3426 (N_3426,N_2227,N_2168);
nand U3427 (N_3427,N_2447,N_2046);
nand U3428 (N_3428,N_2367,N_2066);
xor U3429 (N_3429,N_2107,N_2825);
and U3430 (N_3430,N_2225,N_2268);
or U3431 (N_3431,N_2936,N_2516);
xor U3432 (N_3432,N_2156,N_2508);
xnor U3433 (N_3433,N_2379,N_2257);
or U3434 (N_3434,N_2676,N_2005);
xnor U3435 (N_3435,N_2102,N_2184);
and U3436 (N_3436,N_2017,N_2448);
and U3437 (N_3437,N_2143,N_2954);
xnor U3438 (N_3438,N_2041,N_2885);
and U3439 (N_3439,N_2553,N_2031);
xor U3440 (N_3440,N_2757,N_2889);
nand U3441 (N_3441,N_2575,N_2803);
nor U3442 (N_3442,N_2497,N_2779);
and U3443 (N_3443,N_2410,N_2509);
and U3444 (N_3444,N_2344,N_2374);
or U3445 (N_3445,N_2652,N_2699);
and U3446 (N_3446,N_2386,N_2972);
nand U3447 (N_3447,N_2816,N_2392);
nor U3448 (N_3448,N_2350,N_2847);
xnor U3449 (N_3449,N_2650,N_2724);
nor U3450 (N_3450,N_2720,N_2998);
xor U3451 (N_3451,N_2238,N_2099);
or U3452 (N_3452,N_2078,N_2067);
or U3453 (N_3453,N_2837,N_2368);
xor U3454 (N_3454,N_2193,N_2377);
nand U3455 (N_3455,N_2664,N_2700);
xor U3456 (N_3456,N_2098,N_2573);
or U3457 (N_3457,N_2253,N_2841);
nor U3458 (N_3458,N_2250,N_2961);
xnor U3459 (N_3459,N_2522,N_2925);
nor U3460 (N_3460,N_2207,N_2465);
and U3461 (N_3461,N_2513,N_2242);
xnor U3462 (N_3462,N_2435,N_2629);
and U3463 (N_3463,N_2896,N_2638);
xnor U3464 (N_3464,N_2875,N_2009);
or U3465 (N_3465,N_2305,N_2734);
nand U3466 (N_3466,N_2567,N_2991);
and U3467 (N_3467,N_2727,N_2528);
nor U3468 (N_3468,N_2704,N_2745);
nand U3469 (N_3469,N_2082,N_2244);
and U3470 (N_3470,N_2601,N_2142);
nand U3471 (N_3471,N_2868,N_2951);
and U3472 (N_3472,N_2545,N_2533);
nand U3473 (N_3473,N_2382,N_2792);
or U3474 (N_3474,N_2514,N_2398);
nor U3475 (N_3475,N_2572,N_2668);
nand U3476 (N_3476,N_2163,N_2476);
nor U3477 (N_3477,N_2820,N_2582);
and U3478 (N_3478,N_2340,N_2728);
nand U3479 (N_3479,N_2288,N_2482);
nand U3480 (N_3480,N_2743,N_2843);
nor U3481 (N_3481,N_2032,N_2717);
xor U3482 (N_3482,N_2177,N_2592);
nor U3483 (N_3483,N_2439,N_2957);
or U3484 (N_3484,N_2535,N_2205);
or U3485 (N_3485,N_2703,N_2958);
nor U3486 (N_3486,N_2114,N_2214);
and U3487 (N_3487,N_2411,N_2762);
nand U3488 (N_3488,N_2966,N_2097);
xnor U3489 (N_3489,N_2562,N_2375);
nand U3490 (N_3490,N_2796,N_2696);
nand U3491 (N_3491,N_2161,N_2117);
nor U3492 (N_3492,N_2795,N_2839);
and U3493 (N_3493,N_2452,N_2384);
and U3494 (N_3494,N_2354,N_2987);
and U3495 (N_3495,N_2581,N_2125);
xnor U3496 (N_3496,N_2952,N_2618);
nor U3497 (N_3497,N_2068,N_2443);
nand U3498 (N_3498,N_2378,N_2153);
and U3499 (N_3499,N_2287,N_2807);
nor U3500 (N_3500,N_2318,N_2408);
and U3501 (N_3501,N_2490,N_2815);
or U3502 (N_3502,N_2745,N_2848);
xor U3503 (N_3503,N_2989,N_2640);
and U3504 (N_3504,N_2824,N_2706);
nor U3505 (N_3505,N_2969,N_2245);
xor U3506 (N_3506,N_2814,N_2767);
and U3507 (N_3507,N_2685,N_2675);
and U3508 (N_3508,N_2221,N_2142);
or U3509 (N_3509,N_2652,N_2315);
or U3510 (N_3510,N_2142,N_2880);
and U3511 (N_3511,N_2229,N_2225);
nor U3512 (N_3512,N_2931,N_2583);
nor U3513 (N_3513,N_2125,N_2531);
xnor U3514 (N_3514,N_2387,N_2956);
xor U3515 (N_3515,N_2834,N_2771);
xor U3516 (N_3516,N_2732,N_2353);
and U3517 (N_3517,N_2974,N_2918);
nand U3518 (N_3518,N_2245,N_2234);
nor U3519 (N_3519,N_2492,N_2559);
or U3520 (N_3520,N_2307,N_2922);
and U3521 (N_3521,N_2752,N_2940);
or U3522 (N_3522,N_2611,N_2130);
nand U3523 (N_3523,N_2460,N_2447);
or U3524 (N_3524,N_2008,N_2546);
xor U3525 (N_3525,N_2828,N_2405);
and U3526 (N_3526,N_2031,N_2491);
nor U3527 (N_3527,N_2347,N_2804);
or U3528 (N_3528,N_2738,N_2739);
nand U3529 (N_3529,N_2704,N_2791);
and U3530 (N_3530,N_2244,N_2386);
xnor U3531 (N_3531,N_2955,N_2691);
and U3532 (N_3532,N_2964,N_2360);
xor U3533 (N_3533,N_2116,N_2501);
or U3534 (N_3534,N_2191,N_2318);
and U3535 (N_3535,N_2099,N_2522);
nor U3536 (N_3536,N_2146,N_2578);
and U3537 (N_3537,N_2175,N_2294);
and U3538 (N_3538,N_2781,N_2430);
nor U3539 (N_3539,N_2872,N_2789);
nor U3540 (N_3540,N_2217,N_2932);
nand U3541 (N_3541,N_2729,N_2273);
and U3542 (N_3542,N_2618,N_2711);
and U3543 (N_3543,N_2909,N_2449);
and U3544 (N_3544,N_2220,N_2367);
or U3545 (N_3545,N_2080,N_2875);
or U3546 (N_3546,N_2309,N_2611);
and U3547 (N_3547,N_2381,N_2253);
or U3548 (N_3548,N_2383,N_2666);
xor U3549 (N_3549,N_2092,N_2002);
or U3550 (N_3550,N_2502,N_2345);
or U3551 (N_3551,N_2570,N_2539);
or U3552 (N_3552,N_2079,N_2814);
nand U3553 (N_3553,N_2189,N_2405);
nand U3554 (N_3554,N_2159,N_2981);
and U3555 (N_3555,N_2951,N_2581);
nand U3556 (N_3556,N_2995,N_2953);
and U3557 (N_3557,N_2625,N_2062);
and U3558 (N_3558,N_2303,N_2465);
nand U3559 (N_3559,N_2280,N_2530);
nor U3560 (N_3560,N_2282,N_2732);
xor U3561 (N_3561,N_2700,N_2120);
and U3562 (N_3562,N_2399,N_2712);
or U3563 (N_3563,N_2853,N_2703);
or U3564 (N_3564,N_2132,N_2956);
nor U3565 (N_3565,N_2965,N_2898);
nor U3566 (N_3566,N_2197,N_2874);
and U3567 (N_3567,N_2683,N_2911);
and U3568 (N_3568,N_2496,N_2554);
nor U3569 (N_3569,N_2625,N_2517);
nand U3570 (N_3570,N_2534,N_2181);
nand U3571 (N_3571,N_2222,N_2727);
and U3572 (N_3572,N_2264,N_2468);
and U3573 (N_3573,N_2757,N_2929);
nor U3574 (N_3574,N_2685,N_2937);
nor U3575 (N_3575,N_2942,N_2221);
xnor U3576 (N_3576,N_2529,N_2773);
xor U3577 (N_3577,N_2815,N_2322);
nand U3578 (N_3578,N_2801,N_2121);
or U3579 (N_3579,N_2628,N_2601);
and U3580 (N_3580,N_2722,N_2518);
nor U3581 (N_3581,N_2392,N_2820);
xor U3582 (N_3582,N_2367,N_2349);
nand U3583 (N_3583,N_2121,N_2838);
nand U3584 (N_3584,N_2832,N_2659);
and U3585 (N_3585,N_2780,N_2056);
xor U3586 (N_3586,N_2801,N_2167);
nor U3587 (N_3587,N_2703,N_2952);
nor U3588 (N_3588,N_2383,N_2420);
nand U3589 (N_3589,N_2511,N_2837);
xnor U3590 (N_3590,N_2137,N_2439);
nand U3591 (N_3591,N_2717,N_2639);
and U3592 (N_3592,N_2917,N_2658);
or U3593 (N_3593,N_2517,N_2919);
and U3594 (N_3594,N_2105,N_2454);
nor U3595 (N_3595,N_2206,N_2478);
xor U3596 (N_3596,N_2230,N_2305);
nor U3597 (N_3597,N_2579,N_2246);
or U3598 (N_3598,N_2413,N_2887);
nand U3599 (N_3599,N_2564,N_2668);
nand U3600 (N_3600,N_2407,N_2772);
nor U3601 (N_3601,N_2539,N_2552);
and U3602 (N_3602,N_2018,N_2842);
xor U3603 (N_3603,N_2872,N_2341);
xor U3604 (N_3604,N_2818,N_2456);
nor U3605 (N_3605,N_2557,N_2940);
and U3606 (N_3606,N_2374,N_2211);
and U3607 (N_3607,N_2708,N_2453);
nor U3608 (N_3608,N_2807,N_2132);
or U3609 (N_3609,N_2136,N_2538);
or U3610 (N_3610,N_2520,N_2023);
nor U3611 (N_3611,N_2852,N_2011);
nor U3612 (N_3612,N_2497,N_2071);
or U3613 (N_3613,N_2714,N_2088);
or U3614 (N_3614,N_2380,N_2669);
nand U3615 (N_3615,N_2253,N_2016);
nand U3616 (N_3616,N_2096,N_2146);
nand U3617 (N_3617,N_2530,N_2443);
nor U3618 (N_3618,N_2292,N_2325);
xnor U3619 (N_3619,N_2300,N_2290);
or U3620 (N_3620,N_2704,N_2435);
or U3621 (N_3621,N_2412,N_2778);
xnor U3622 (N_3622,N_2468,N_2093);
nand U3623 (N_3623,N_2637,N_2619);
and U3624 (N_3624,N_2069,N_2249);
xnor U3625 (N_3625,N_2593,N_2984);
and U3626 (N_3626,N_2643,N_2487);
and U3627 (N_3627,N_2621,N_2179);
nor U3628 (N_3628,N_2720,N_2444);
xor U3629 (N_3629,N_2685,N_2175);
xor U3630 (N_3630,N_2272,N_2301);
or U3631 (N_3631,N_2114,N_2433);
nor U3632 (N_3632,N_2079,N_2158);
and U3633 (N_3633,N_2279,N_2686);
and U3634 (N_3634,N_2265,N_2395);
nor U3635 (N_3635,N_2525,N_2806);
xnor U3636 (N_3636,N_2167,N_2105);
or U3637 (N_3637,N_2668,N_2657);
nor U3638 (N_3638,N_2481,N_2078);
or U3639 (N_3639,N_2130,N_2115);
xnor U3640 (N_3640,N_2073,N_2155);
nor U3641 (N_3641,N_2586,N_2613);
nand U3642 (N_3642,N_2511,N_2960);
or U3643 (N_3643,N_2662,N_2867);
or U3644 (N_3644,N_2170,N_2963);
and U3645 (N_3645,N_2340,N_2252);
nor U3646 (N_3646,N_2643,N_2128);
and U3647 (N_3647,N_2570,N_2180);
nor U3648 (N_3648,N_2510,N_2622);
nor U3649 (N_3649,N_2424,N_2705);
or U3650 (N_3650,N_2623,N_2788);
and U3651 (N_3651,N_2266,N_2025);
and U3652 (N_3652,N_2912,N_2480);
and U3653 (N_3653,N_2500,N_2142);
xor U3654 (N_3654,N_2741,N_2561);
nand U3655 (N_3655,N_2038,N_2477);
xor U3656 (N_3656,N_2466,N_2117);
nor U3657 (N_3657,N_2187,N_2592);
nand U3658 (N_3658,N_2237,N_2593);
nor U3659 (N_3659,N_2346,N_2399);
and U3660 (N_3660,N_2959,N_2858);
nand U3661 (N_3661,N_2019,N_2873);
nand U3662 (N_3662,N_2361,N_2356);
and U3663 (N_3663,N_2771,N_2021);
or U3664 (N_3664,N_2387,N_2846);
or U3665 (N_3665,N_2728,N_2601);
and U3666 (N_3666,N_2877,N_2589);
or U3667 (N_3667,N_2669,N_2130);
xnor U3668 (N_3668,N_2068,N_2027);
nor U3669 (N_3669,N_2111,N_2023);
xnor U3670 (N_3670,N_2067,N_2936);
nor U3671 (N_3671,N_2135,N_2444);
and U3672 (N_3672,N_2655,N_2869);
nand U3673 (N_3673,N_2694,N_2927);
nor U3674 (N_3674,N_2456,N_2736);
and U3675 (N_3675,N_2168,N_2187);
nor U3676 (N_3676,N_2315,N_2389);
xnor U3677 (N_3677,N_2764,N_2752);
and U3678 (N_3678,N_2269,N_2933);
and U3679 (N_3679,N_2337,N_2481);
and U3680 (N_3680,N_2141,N_2975);
nand U3681 (N_3681,N_2175,N_2546);
xor U3682 (N_3682,N_2692,N_2323);
nand U3683 (N_3683,N_2423,N_2182);
nor U3684 (N_3684,N_2952,N_2435);
and U3685 (N_3685,N_2727,N_2525);
and U3686 (N_3686,N_2763,N_2943);
or U3687 (N_3687,N_2302,N_2839);
nand U3688 (N_3688,N_2818,N_2770);
nor U3689 (N_3689,N_2919,N_2615);
nor U3690 (N_3690,N_2220,N_2928);
nand U3691 (N_3691,N_2885,N_2662);
xor U3692 (N_3692,N_2474,N_2016);
nand U3693 (N_3693,N_2695,N_2327);
nor U3694 (N_3694,N_2840,N_2596);
nand U3695 (N_3695,N_2985,N_2592);
or U3696 (N_3696,N_2194,N_2024);
nand U3697 (N_3697,N_2250,N_2886);
nand U3698 (N_3698,N_2193,N_2099);
xor U3699 (N_3699,N_2622,N_2046);
nand U3700 (N_3700,N_2773,N_2308);
nand U3701 (N_3701,N_2947,N_2140);
nand U3702 (N_3702,N_2319,N_2927);
or U3703 (N_3703,N_2896,N_2852);
nor U3704 (N_3704,N_2650,N_2452);
or U3705 (N_3705,N_2791,N_2664);
or U3706 (N_3706,N_2346,N_2508);
nor U3707 (N_3707,N_2223,N_2911);
and U3708 (N_3708,N_2426,N_2234);
or U3709 (N_3709,N_2086,N_2517);
nor U3710 (N_3710,N_2584,N_2732);
nor U3711 (N_3711,N_2465,N_2562);
or U3712 (N_3712,N_2686,N_2550);
or U3713 (N_3713,N_2314,N_2005);
xnor U3714 (N_3714,N_2025,N_2723);
or U3715 (N_3715,N_2535,N_2767);
nor U3716 (N_3716,N_2664,N_2306);
nor U3717 (N_3717,N_2194,N_2090);
and U3718 (N_3718,N_2938,N_2653);
or U3719 (N_3719,N_2210,N_2486);
or U3720 (N_3720,N_2943,N_2581);
xnor U3721 (N_3721,N_2041,N_2617);
xnor U3722 (N_3722,N_2731,N_2849);
and U3723 (N_3723,N_2444,N_2769);
nor U3724 (N_3724,N_2721,N_2811);
nor U3725 (N_3725,N_2907,N_2381);
xnor U3726 (N_3726,N_2723,N_2989);
and U3727 (N_3727,N_2650,N_2850);
and U3728 (N_3728,N_2545,N_2213);
or U3729 (N_3729,N_2735,N_2730);
and U3730 (N_3730,N_2873,N_2468);
or U3731 (N_3731,N_2249,N_2605);
and U3732 (N_3732,N_2239,N_2544);
xnor U3733 (N_3733,N_2910,N_2181);
or U3734 (N_3734,N_2364,N_2142);
nand U3735 (N_3735,N_2380,N_2874);
nand U3736 (N_3736,N_2957,N_2057);
nand U3737 (N_3737,N_2214,N_2569);
nor U3738 (N_3738,N_2449,N_2830);
nand U3739 (N_3739,N_2714,N_2708);
nor U3740 (N_3740,N_2763,N_2837);
nor U3741 (N_3741,N_2904,N_2820);
or U3742 (N_3742,N_2173,N_2994);
nor U3743 (N_3743,N_2259,N_2084);
or U3744 (N_3744,N_2402,N_2249);
or U3745 (N_3745,N_2725,N_2255);
xnor U3746 (N_3746,N_2699,N_2148);
or U3747 (N_3747,N_2193,N_2540);
xnor U3748 (N_3748,N_2483,N_2751);
and U3749 (N_3749,N_2175,N_2122);
xnor U3750 (N_3750,N_2112,N_2960);
xor U3751 (N_3751,N_2618,N_2722);
nand U3752 (N_3752,N_2844,N_2369);
nand U3753 (N_3753,N_2877,N_2234);
and U3754 (N_3754,N_2880,N_2910);
nor U3755 (N_3755,N_2745,N_2553);
nor U3756 (N_3756,N_2099,N_2479);
nand U3757 (N_3757,N_2789,N_2521);
or U3758 (N_3758,N_2173,N_2236);
and U3759 (N_3759,N_2895,N_2792);
nor U3760 (N_3760,N_2310,N_2065);
nand U3761 (N_3761,N_2886,N_2454);
or U3762 (N_3762,N_2922,N_2465);
xnor U3763 (N_3763,N_2430,N_2973);
nor U3764 (N_3764,N_2852,N_2933);
and U3765 (N_3765,N_2766,N_2486);
nor U3766 (N_3766,N_2351,N_2541);
xnor U3767 (N_3767,N_2181,N_2606);
nor U3768 (N_3768,N_2765,N_2891);
or U3769 (N_3769,N_2090,N_2700);
and U3770 (N_3770,N_2699,N_2260);
xnor U3771 (N_3771,N_2037,N_2936);
xnor U3772 (N_3772,N_2347,N_2113);
and U3773 (N_3773,N_2170,N_2825);
nand U3774 (N_3774,N_2102,N_2930);
nor U3775 (N_3775,N_2401,N_2469);
xnor U3776 (N_3776,N_2292,N_2528);
or U3777 (N_3777,N_2568,N_2982);
nor U3778 (N_3778,N_2660,N_2226);
nor U3779 (N_3779,N_2226,N_2200);
and U3780 (N_3780,N_2127,N_2926);
xnor U3781 (N_3781,N_2086,N_2768);
xnor U3782 (N_3782,N_2621,N_2197);
xnor U3783 (N_3783,N_2405,N_2216);
nand U3784 (N_3784,N_2766,N_2868);
or U3785 (N_3785,N_2058,N_2411);
and U3786 (N_3786,N_2365,N_2407);
nor U3787 (N_3787,N_2872,N_2014);
xor U3788 (N_3788,N_2458,N_2515);
nor U3789 (N_3789,N_2481,N_2676);
nor U3790 (N_3790,N_2395,N_2014);
and U3791 (N_3791,N_2935,N_2486);
nand U3792 (N_3792,N_2348,N_2873);
nand U3793 (N_3793,N_2878,N_2822);
or U3794 (N_3794,N_2328,N_2862);
nand U3795 (N_3795,N_2693,N_2635);
and U3796 (N_3796,N_2373,N_2530);
nor U3797 (N_3797,N_2273,N_2520);
nor U3798 (N_3798,N_2120,N_2846);
xnor U3799 (N_3799,N_2476,N_2060);
nor U3800 (N_3800,N_2728,N_2561);
xnor U3801 (N_3801,N_2943,N_2058);
nand U3802 (N_3802,N_2648,N_2610);
nor U3803 (N_3803,N_2574,N_2576);
and U3804 (N_3804,N_2187,N_2475);
nand U3805 (N_3805,N_2639,N_2691);
nor U3806 (N_3806,N_2457,N_2523);
or U3807 (N_3807,N_2169,N_2869);
xnor U3808 (N_3808,N_2505,N_2404);
and U3809 (N_3809,N_2432,N_2146);
nand U3810 (N_3810,N_2206,N_2387);
nor U3811 (N_3811,N_2097,N_2428);
nand U3812 (N_3812,N_2723,N_2287);
nand U3813 (N_3813,N_2873,N_2024);
nor U3814 (N_3814,N_2455,N_2412);
nand U3815 (N_3815,N_2716,N_2847);
and U3816 (N_3816,N_2319,N_2778);
or U3817 (N_3817,N_2634,N_2850);
and U3818 (N_3818,N_2547,N_2835);
or U3819 (N_3819,N_2692,N_2468);
or U3820 (N_3820,N_2106,N_2231);
xnor U3821 (N_3821,N_2394,N_2463);
and U3822 (N_3822,N_2645,N_2029);
nor U3823 (N_3823,N_2989,N_2956);
and U3824 (N_3824,N_2521,N_2849);
xnor U3825 (N_3825,N_2533,N_2379);
nor U3826 (N_3826,N_2375,N_2987);
or U3827 (N_3827,N_2611,N_2807);
nand U3828 (N_3828,N_2851,N_2662);
nand U3829 (N_3829,N_2767,N_2949);
nand U3830 (N_3830,N_2408,N_2571);
nor U3831 (N_3831,N_2942,N_2011);
or U3832 (N_3832,N_2572,N_2624);
nand U3833 (N_3833,N_2191,N_2597);
nand U3834 (N_3834,N_2726,N_2222);
or U3835 (N_3835,N_2916,N_2058);
and U3836 (N_3836,N_2117,N_2271);
nand U3837 (N_3837,N_2683,N_2885);
nand U3838 (N_3838,N_2237,N_2059);
and U3839 (N_3839,N_2811,N_2718);
nand U3840 (N_3840,N_2049,N_2977);
or U3841 (N_3841,N_2837,N_2708);
or U3842 (N_3842,N_2579,N_2164);
nand U3843 (N_3843,N_2828,N_2110);
xnor U3844 (N_3844,N_2505,N_2711);
or U3845 (N_3845,N_2879,N_2918);
or U3846 (N_3846,N_2468,N_2767);
or U3847 (N_3847,N_2295,N_2992);
or U3848 (N_3848,N_2335,N_2665);
xor U3849 (N_3849,N_2339,N_2643);
xor U3850 (N_3850,N_2838,N_2080);
nand U3851 (N_3851,N_2127,N_2729);
nor U3852 (N_3852,N_2215,N_2427);
xnor U3853 (N_3853,N_2936,N_2792);
or U3854 (N_3854,N_2441,N_2943);
nand U3855 (N_3855,N_2844,N_2848);
or U3856 (N_3856,N_2176,N_2577);
and U3857 (N_3857,N_2412,N_2452);
nand U3858 (N_3858,N_2132,N_2927);
nor U3859 (N_3859,N_2974,N_2726);
and U3860 (N_3860,N_2873,N_2591);
nor U3861 (N_3861,N_2926,N_2574);
or U3862 (N_3862,N_2861,N_2070);
nand U3863 (N_3863,N_2472,N_2910);
nor U3864 (N_3864,N_2580,N_2323);
nand U3865 (N_3865,N_2104,N_2123);
nor U3866 (N_3866,N_2278,N_2217);
xor U3867 (N_3867,N_2633,N_2243);
nand U3868 (N_3868,N_2095,N_2189);
xor U3869 (N_3869,N_2494,N_2007);
or U3870 (N_3870,N_2738,N_2211);
and U3871 (N_3871,N_2002,N_2364);
xnor U3872 (N_3872,N_2406,N_2651);
or U3873 (N_3873,N_2007,N_2232);
or U3874 (N_3874,N_2856,N_2173);
or U3875 (N_3875,N_2597,N_2645);
xor U3876 (N_3876,N_2633,N_2833);
and U3877 (N_3877,N_2878,N_2681);
nand U3878 (N_3878,N_2404,N_2892);
nor U3879 (N_3879,N_2751,N_2144);
nand U3880 (N_3880,N_2960,N_2947);
nand U3881 (N_3881,N_2347,N_2810);
or U3882 (N_3882,N_2177,N_2994);
and U3883 (N_3883,N_2935,N_2992);
nand U3884 (N_3884,N_2960,N_2577);
or U3885 (N_3885,N_2481,N_2170);
nand U3886 (N_3886,N_2145,N_2034);
and U3887 (N_3887,N_2976,N_2560);
or U3888 (N_3888,N_2869,N_2067);
nand U3889 (N_3889,N_2753,N_2681);
or U3890 (N_3890,N_2452,N_2577);
or U3891 (N_3891,N_2441,N_2029);
nand U3892 (N_3892,N_2447,N_2892);
nor U3893 (N_3893,N_2108,N_2972);
nand U3894 (N_3894,N_2584,N_2445);
nor U3895 (N_3895,N_2085,N_2976);
nor U3896 (N_3896,N_2350,N_2192);
or U3897 (N_3897,N_2968,N_2437);
and U3898 (N_3898,N_2320,N_2449);
xor U3899 (N_3899,N_2682,N_2245);
xor U3900 (N_3900,N_2195,N_2399);
xor U3901 (N_3901,N_2882,N_2533);
nand U3902 (N_3902,N_2013,N_2925);
nand U3903 (N_3903,N_2433,N_2141);
nor U3904 (N_3904,N_2245,N_2156);
nand U3905 (N_3905,N_2367,N_2819);
and U3906 (N_3906,N_2881,N_2243);
and U3907 (N_3907,N_2544,N_2256);
xnor U3908 (N_3908,N_2510,N_2565);
nand U3909 (N_3909,N_2789,N_2266);
and U3910 (N_3910,N_2936,N_2388);
nor U3911 (N_3911,N_2971,N_2169);
and U3912 (N_3912,N_2428,N_2928);
or U3913 (N_3913,N_2087,N_2747);
or U3914 (N_3914,N_2358,N_2208);
nor U3915 (N_3915,N_2392,N_2379);
nand U3916 (N_3916,N_2918,N_2865);
nor U3917 (N_3917,N_2843,N_2604);
and U3918 (N_3918,N_2510,N_2524);
nand U3919 (N_3919,N_2284,N_2684);
or U3920 (N_3920,N_2920,N_2028);
and U3921 (N_3921,N_2515,N_2375);
nor U3922 (N_3922,N_2751,N_2957);
nand U3923 (N_3923,N_2614,N_2786);
and U3924 (N_3924,N_2792,N_2409);
xor U3925 (N_3925,N_2912,N_2997);
and U3926 (N_3926,N_2404,N_2187);
and U3927 (N_3927,N_2483,N_2038);
and U3928 (N_3928,N_2225,N_2057);
xnor U3929 (N_3929,N_2672,N_2026);
nand U3930 (N_3930,N_2720,N_2866);
nor U3931 (N_3931,N_2284,N_2816);
xnor U3932 (N_3932,N_2913,N_2012);
and U3933 (N_3933,N_2627,N_2348);
xnor U3934 (N_3934,N_2205,N_2734);
nor U3935 (N_3935,N_2706,N_2084);
xor U3936 (N_3936,N_2346,N_2580);
or U3937 (N_3937,N_2150,N_2950);
xnor U3938 (N_3938,N_2053,N_2566);
nor U3939 (N_3939,N_2931,N_2896);
xnor U3940 (N_3940,N_2751,N_2933);
and U3941 (N_3941,N_2290,N_2192);
nor U3942 (N_3942,N_2073,N_2500);
and U3943 (N_3943,N_2585,N_2925);
and U3944 (N_3944,N_2865,N_2536);
or U3945 (N_3945,N_2189,N_2251);
or U3946 (N_3946,N_2820,N_2767);
or U3947 (N_3947,N_2133,N_2419);
nor U3948 (N_3948,N_2557,N_2595);
or U3949 (N_3949,N_2283,N_2628);
nand U3950 (N_3950,N_2558,N_2894);
xnor U3951 (N_3951,N_2295,N_2175);
nand U3952 (N_3952,N_2101,N_2357);
and U3953 (N_3953,N_2995,N_2806);
nand U3954 (N_3954,N_2794,N_2997);
or U3955 (N_3955,N_2910,N_2551);
or U3956 (N_3956,N_2287,N_2709);
xnor U3957 (N_3957,N_2150,N_2393);
and U3958 (N_3958,N_2698,N_2452);
nor U3959 (N_3959,N_2007,N_2500);
nor U3960 (N_3960,N_2538,N_2059);
and U3961 (N_3961,N_2798,N_2845);
nor U3962 (N_3962,N_2953,N_2780);
nor U3963 (N_3963,N_2191,N_2795);
nand U3964 (N_3964,N_2130,N_2330);
and U3965 (N_3965,N_2884,N_2382);
nand U3966 (N_3966,N_2522,N_2545);
nand U3967 (N_3967,N_2200,N_2023);
xnor U3968 (N_3968,N_2594,N_2625);
nand U3969 (N_3969,N_2570,N_2158);
xor U3970 (N_3970,N_2998,N_2909);
and U3971 (N_3971,N_2418,N_2370);
nand U3972 (N_3972,N_2905,N_2001);
and U3973 (N_3973,N_2728,N_2793);
and U3974 (N_3974,N_2144,N_2333);
xnor U3975 (N_3975,N_2659,N_2788);
and U3976 (N_3976,N_2001,N_2700);
or U3977 (N_3977,N_2093,N_2100);
or U3978 (N_3978,N_2630,N_2615);
nor U3979 (N_3979,N_2219,N_2206);
and U3980 (N_3980,N_2455,N_2330);
nand U3981 (N_3981,N_2130,N_2485);
xnor U3982 (N_3982,N_2657,N_2735);
and U3983 (N_3983,N_2223,N_2252);
nor U3984 (N_3984,N_2089,N_2870);
nor U3985 (N_3985,N_2917,N_2257);
nand U3986 (N_3986,N_2717,N_2595);
nor U3987 (N_3987,N_2411,N_2976);
and U3988 (N_3988,N_2114,N_2950);
and U3989 (N_3989,N_2747,N_2937);
xnor U3990 (N_3990,N_2664,N_2716);
or U3991 (N_3991,N_2884,N_2431);
and U3992 (N_3992,N_2394,N_2138);
nor U3993 (N_3993,N_2599,N_2412);
or U3994 (N_3994,N_2160,N_2438);
nand U3995 (N_3995,N_2220,N_2096);
or U3996 (N_3996,N_2085,N_2161);
xor U3997 (N_3997,N_2800,N_2556);
xnor U3998 (N_3998,N_2839,N_2384);
nor U3999 (N_3999,N_2007,N_2550);
or U4000 (N_4000,N_3077,N_3764);
and U4001 (N_4001,N_3407,N_3941);
and U4002 (N_4002,N_3674,N_3473);
nor U4003 (N_4003,N_3825,N_3837);
and U4004 (N_4004,N_3109,N_3740);
xor U4005 (N_4005,N_3430,N_3507);
or U4006 (N_4006,N_3349,N_3601);
xnor U4007 (N_4007,N_3503,N_3909);
and U4008 (N_4008,N_3558,N_3590);
nor U4009 (N_4009,N_3446,N_3708);
nand U4010 (N_4010,N_3947,N_3653);
nor U4011 (N_4011,N_3212,N_3681);
or U4012 (N_4012,N_3311,N_3834);
nor U4013 (N_4013,N_3651,N_3857);
nor U4014 (N_4014,N_3383,N_3898);
and U4015 (N_4015,N_3715,N_3358);
nand U4016 (N_4016,N_3922,N_3888);
or U4017 (N_4017,N_3238,N_3821);
xnor U4018 (N_4018,N_3805,N_3600);
nor U4019 (N_4019,N_3802,N_3999);
nand U4020 (N_4020,N_3610,N_3167);
nand U4021 (N_4021,N_3647,N_3052);
xnor U4022 (N_4022,N_3424,N_3344);
nand U4023 (N_4023,N_3916,N_3572);
nor U4024 (N_4024,N_3788,N_3047);
or U4025 (N_4025,N_3152,N_3139);
nand U4026 (N_4026,N_3867,N_3454);
xor U4027 (N_4027,N_3658,N_3900);
nand U4028 (N_4028,N_3712,N_3771);
or U4029 (N_4029,N_3186,N_3002);
xnor U4030 (N_4030,N_3725,N_3761);
and U4031 (N_4031,N_3975,N_3204);
nor U4032 (N_4032,N_3272,N_3846);
xnor U4033 (N_4033,N_3353,N_3505);
nor U4034 (N_4034,N_3923,N_3874);
or U4035 (N_4035,N_3736,N_3535);
and U4036 (N_4036,N_3908,N_3046);
and U4037 (N_4037,N_3244,N_3560);
xor U4038 (N_4038,N_3032,N_3648);
and U4039 (N_4039,N_3456,N_3483);
and U4040 (N_4040,N_3141,N_3745);
nor U4041 (N_4041,N_3132,N_3478);
xor U4042 (N_4042,N_3897,N_3369);
xnor U4043 (N_4043,N_3768,N_3758);
nand U4044 (N_4044,N_3532,N_3190);
nand U4045 (N_4045,N_3067,N_3952);
and U4046 (N_4046,N_3408,N_3950);
or U4047 (N_4047,N_3119,N_3113);
xnor U4048 (N_4048,N_3543,N_3733);
or U4049 (N_4049,N_3472,N_3022);
nor U4050 (N_4050,N_3288,N_3611);
nand U4051 (N_4051,N_3954,N_3638);
nand U4052 (N_4052,N_3176,N_3006);
nand U4053 (N_4053,N_3054,N_3692);
and U4054 (N_4054,N_3627,N_3631);
and U4055 (N_4055,N_3854,N_3342);
nor U4056 (N_4056,N_3877,N_3667);
nand U4057 (N_4057,N_3235,N_3123);
xor U4058 (N_4058,N_3596,N_3936);
nand U4059 (N_4059,N_3033,N_3556);
or U4060 (N_4060,N_3792,N_3071);
xnor U4061 (N_4061,N_3826,N_3907);
and U4062 (N_4062,N_3914,N_3830);
xor U4063 (N_4063,N_3892,N_3158);
xor U4064 (N_4064,N_3459,N_3973);
nand U4065 (N_4065,N_3078,N_3542);
nand U4066 (N_4066,N_3777,N_3436);
nor U4067 (N_4067,N_3106,N_3434);
nand U4068 (N_4068,N_3739,N_3561);
xnor U4069 (N_4069,N_3575,N_3347);
and U4070 (N_4070,N_3236,N_3426);
or U4071 (N_4071,N_3191,N_3637);
xor U4072 (N_4072,N_3544,N_3079);
xor U4073 (N_4073,N_3958,N_3640);
or U4074 (N_4074,N_3380,N_3980);
and U4075 (N_4075,N_3808,N_3809);
nor U4076 (N_4076,N_3604,N_3084);
and U4077 (N_4077,N_3428,N_3417);
or U4078 (N_4078,N_3420,N_3262);
and U4079 (N_4079,N_3850,N_3188);
nor U4080 (N_4080,N_3207,N_3378);
nor U4081 (N_4081,N_3030,N_3522);
and U4082 (N_4082,N_3260,N_3744);
xnor U4083 (N_4083,N_3121,N_3770);
or U4084 (N_4084,N_3474,N_3858);
nor U4085 (N_4085,N_3806,N_3061);
nor U4086 (N_4086,N_3324,N_3069);
or U4087 (N_4087,N_3114,N_3107);
xnor U4088 (N_4088,N_3406,N_3902);
nand U4089 (N_4089,N_3402,N_3865);
or U4090 (N_4090,N_3889,N_3643);
nand U4091 (N_4091,N_3416,N_3812);
nand U4092 (N_4092,N_3682,N_3634);
and U4093 (N_4093,N_3748,N_3290);
nand U4094 (N_4094,N_3133,N_3202);
nor U4095 (N_4095,N_3719,N_3623);
nor U4096 (N_4096,N_3977,N_3267);
xor U4097 (N_4097,N_3289,N_3278);
nand U4098 (N_4098,N_3512,N_3820);
and U4099 (N_4099,N_3211,N_3896);
xor U4100 (N_4100,N_3782,N_3237);
nor U4101 (N_4101,N_3752,N_3910);
nor U4102 (N_4102,N_3528,N_3751);
or U4103 (N_4103,N_3904,N_3774);
and U4104 (N_4104,N_3793,N_3527);
xor U4105 (N_4105,N_3060,N_3042);
or U4106 (N_4106,N_3285,N_3762);
xnor U4107 (N_4107,N_3799,N_3589);
nand U4108 (N_4108,N_3956,N_3763);
nor U4109 (N_4109,N_3495,N_3707);
nor U4110 (N_4110,N_3394,N_3189);
nand U4111 (N_4111,N_3964,N_3165);
xor U4112 (N_4112,N_3619,N_3673);
xor U4113 (N_4113,N_3435,N_3076);
or U4114 (N_4114,N_3146,N_3921);
and U4115 (N_4115,N_3192,N_3336);
or U4116 (N_4116,N_3912,N_3247);
or U4117 (N_4117,N_3471,N_3234);
xnor U4118 (N_4118,N_3592,N_3838);
nor U4119 (N_4119,N_3205,N_3476);
nand U4120 (N_4120,N_3804,N_3537);
and U4121 (N_4121,N_3924,N_3750);
and U4122 (N_4122,N_3790,N_3333);
and U4123 (N_4123,N_3754,N_3690);
xnor U4124 (N_4124,N_3635,N_3817);
and U4125 (N_4125,N_3957,N_3756);
nor U4126 (N_4126,N_3268,N_3074);
nand U4127 (N_4127,N_3531,N_3991);
nor U4128 (N_4128,N_3348,N_3683);
or U4129 (N_4129,N_3847,N_3431);
xor U4130 (N_4130,N_3618,N_3905);
xor U4131 (N_4131,N_3081,N_3961);
or U4132 (N_4132,N_3341,N_3546);
and U4133 (N_4133,N_3811,N_3582);
or U4134 (N_4134,N_3387,N_3917);
nand U4135 (N_4135,N_3376,N_3475);
or U4136 (N_4136,N_3704,N_3509);
nand U4137 (N_4137,N_3399,N_3019);
or U4138 (N_4138,N_3105,N_3853);
or U4139 (N_4139,N_3721,N_3816);
and U4140 (N_4140,N_3666,N_3553);
and U4141 (N_4141,N_3529,N_3020);
nand U4142 (N_4142,N_3965,N_3021);
and U4143 (N_4143,N_3685,N_3769);
nand U4144 (N_4144,N_3072,N_3603);
and U4145 (N_4145,N_3625,N_3617);
and U4146 (N_4146,N_3641,N_3229);
xor U4147 (N_4147,N_3354,N_3126);
nand U4148 (N_4148,N_3818,N_3959);
xnor U4149 (N_4149,N_3494,N_3421);
nand U4150 (N_4150,N_3286,N_3903);
nor U4151 (N_4151,N_3279,N_3918);
xor U4152 (N_4152,N_3265,N_3044);
or U4153 (N_4153,N_3058,N_3384);
nand U4154 (N_4154,N_3116,N_3514);
xnor U4155 (N_4155,N_3263,N_3028);
and U4156 (N_4156,N_3438,N_3845);
nor U4157 (N_4157,N_3566,N_3577);
and U4158 (N_4158,N_3179,N_3773);
xnor U4159 (N_4159,N_3995,N_3616);
and U4160 (N_4160,N_3962,N_3523);
nor U4161 (N_4161,N_3292,N_3082);
xnor U4162 (N_4162,N_3876,N_3287);
and U4163 (N_4163,N_3517,N_3310);
nor U4164 (N_4164,N_3415,N_3639);
and U4165 (N_4165,N_3729,N_3714);
or U4166 (N_4166,N_3864,N_3562);
and U4167 (N_4167,N_3781,N_3183);
nor U4168 (N_4168,N_3901,N_3632);
nor U4169 (N_4169,N_3148,N_3766);
or U4170 (N_4170,N_3662,N_3065);
nand U4171 (N_4171,N_3423,N_3484);
nand U4172 (N_4172,N_3025,N_3087);
nor U4173 (N_4173,N_3318,N_3791);
xnor U4174 (N_4174,N_3036,N_3095);
and U4175 (N_4175,N_3440,N_3598);
nand U4176 (N_4176,N_3366,N_3615);
nand U4177 (N_4177,N_3419,N_3501);
or U4178 (N_4178,N_3231,N_3429);
nor U4179 (N_4179,N_3579,N_3775);
or U4180 (N_4180,N_3026,N_3468);
nand U4181 (N_4181,N_3391,N_3645);
xnor U4182 (N_4182,N_3166,N_3242);
or U4183 (N_4183,N_3227,N_3689);
nor U4184 (N_4184,N_3023,N_3187);
and U4185 (N_4185,N_3097,N_3258);
and U4186 (N_4186,N_3252,N_3226);
xnor U4187 (N_4187,N_3539,N_3613);
nor U4188 (N_4188,N_3822,N_3986);
nand U4189 (N_4189,N_3088,N_3614);
or U4190 (N_4190,N_3913,N_3352);
nor U4191 (N_4191,N_3210,N_3937);
and U4192 (N_4192,N_3153,N_3570);
nand U4193 (N_4193,N_3480,N_3017);
and U4194 (N_4194,N_3269,N_3313);
nand U4195 (N_4195,N_3966,N_3098);
or U4196 (N_4196,N_3147,N_3624);
and U4197 (N_4197,N_3283,N_3228);
or U4198 (N_4198,N_3451,N_3270);
nand U4199 (N_4199,N_3320,N_3963);
nand U4200 (N_4200,N_3411,N_3515);
or U4201 (N_4201,N_3452,N_3711);
or U4202 (N_4202,N_3660,N_3599);
xor U4203 (N_4203,N_3266,N_3893);
and U4204 (N_4204,N_3005,N_3743);
or U4205 (N_4205,N_3698,N_3851);
xor U4206 (N_4206,N_3810,N_3524);
and U4207 (N_4207,N_3983,N_3457);
and U4208 (N_4208,N_3597,N_3979);
nor U4209 (N_4209,N_3776,N_3785);
nor U4210 (N_4210,N_3256,N_3856);
and U4211 (N_4211,N_3988,N_3671);
or U4212 (N_4212,N_3772,N_3753);
and U4213 (N_4213,N_3371,N_3306);
nor U4214 (N_4214,N_3724,N_3945);
nor U4215 (N_4215,N_3307,N_3414);
nor U4216 (N_4216,N_3465,N_3073);
nor U4217 (N_4217,N_3469,N_3209);
xnor U4218 (N_4218,N_3932,N_3159);
nor U4219 (N_4219,N_3949,N_3742);
and U4220 (N_4220,N_3053,N_3706);
or U4221 (N_4221,N_3377,N_3175);
or U4222 (N_4222,N_3703,N_3879);
nor U4223 (N_4223,N_3455,N_3299);
nor U4224 (N_4224,N_3008,N_3841);
xnor U4225 (N_4225,N_3241,N_3738);
xor U4226 (N_4226,N_3824,N_3254);
and U4227 (N_4227,N_3388,N_3112);
xor U4228 (N_4228,N_3092,N_3382);
nor U4229 (N_4229,N_3437,N_3564);
xnor U4230 (N_4230,N_3181,N_3894);
or U4231 (N_4231,N_3787,N_3933);
nor U4232 (N_4232,N_3878,N_3591);
and U4233 (N_4233,N_3545,N_3277);
and U4234 (N_4234,N_3346,N_3122);
nor U4235 (N_4235,N_3041,N_3246);
nand U4236 (N_4236,N_3654,N_3726);
xnor U4237 (N_4237,N_3606,N_3232);
nand U4238 (N_4238,N_3884,N_3068);
or U4239 (N_4239,N_3602,N_3140);
xnor U4240 (N_4240,N_3482,N_3233);
nor U4241 (N_4241,N_3677,N_3565);
or U4242 (N_4242,N_3548,N_3580);
xnor U4243 (N_4243,N_3872,N_3062);
nor U4244 (N_4244,N_3222,N_3134);
and U4245 (N_4245,N_3412,N_3303);
and U4246 (N_4246,N_3686,N_3281);
nor U4247 (N_4247,N_3997,N_3389);
nor U4248 (N_4248,N_3035,N_3086);
xnor U4249 (N_4249,N_3118,N_3011);
nand U4250 (N_4250,N_3938,N_3538);
nor U4251 (N_4251,N_3843,N_3305);
or U4252 (N_4252,N_3587,N_3361);
and U4253 (N_4253,N_3037,N_3275);
nand U4254 (N_4254,N_3261,N_3193);
or U4255 (N_4255,N_3803,N_3749);
and U4256 (N_4256,N_3883,N_3732);
or U4257 (N_4257,N_3955,N_3401);
or U4258 (N_4258,N_3518,N_3302);
nor U4259 (N_4259,N_3264,N_3144);
nor U4260 (N_4260,N_3747,N_3444);
xor U4261 (N_4261,N_3184,N_3869);
and U4262 (N_4262,N_3701,N_3636);
xnor U4263 (N_4263,N_3185,N_3737);
and U4264 (N_4264,N_3362,N_3511);
nand U4265 (N_4265,N_3767,N_3488);
and U4266 (N_4266,N_3013,N_3149);
or U4267 (N_4267,N_3547,N_3194);
nor U4268 (N_4268,N_3162,N_3576);
and U4269 (N_4269,N_3398,N_3293);
nor U4270 (N_4270,N_3108,N_3691);
nand U4271 (N_4271,N_3325,N_3064);
nand U4272 (N_4272,N_3374,N_3470);
and U4273 (N_4273,N_3493,N_3996);
nor U4274 (N_4274,N_3550,N_3009);
xor U4275 (N_4275,N_3447,N_3934);
and U4276 (N_4276,N_3206,N_3091);
or U4277 (N_4277,N_3218,N_3797);
nor U4278 (N_4278,N_3276,N_3439);
nor U4279 (N_4279,N_3508,N_3427);
and U4280 (N_4280,N_3038,N_3372);
and U4281 (N_4281,N_3066,N_3059);
or U4282 (N_4282,N_3160,N_3661);
nand U4283 (N_4283,N_3759,N_3578);
nand U4284 (N_4284,N_3432,N_3314);
nand U4285 (N_4285,N_3540,N_3899);
and U4286 (N_4286,N_3720,N_3819);
nand U4287 (N_4287,N_3607,N_3223);
or U4288 (N_4288,N_3855,N_3075);
and U4289 (N_4289,N_3882,N_3679);
or U4290 (N_4290,N_3669,N_3464);
nor U4291 (N_4291,N_3583,N_3168);
or U4292 (N_4292,N_3200,N_3367);
and U4293 (N_4293,N_3848,N_3827);
and U4294 (N_4294,N_3467,N_3029);
or U4295 (N_4295,N_3696,N_3807);
nand U4296 (N_4296,N_3612,N_3201);
nand U4297 (N_4297,N_3001,N_3784);
xor U4298 (N_4298,N_3693,N_3214);
nand U4299 (N_4299,N_3940,N_3502);
nor U4300 (N_4300,N_3115,N_3866);
or U4301 (N_4301,N_3757,N_3971);
xnor U4302 (N_4302,N_3151,N_3513);
and U4303 (N_4303,N_3368,N_3489);
nand U4304 (N_4304,N_3657,N_3911);
xnor U4305 (N_4305,N_3328,N_3626);
nor U4306 (N_4306,N_3094,N_3859);
nand U4307 (N_4307,N_3943,N_3968);
nand U4308 (N_4308,N_3213,N_3173);
nand U4309 (N_4309,N_3128,N_3220);
nand U4310 (N_4310,N_3702,N_3257);
nor U4311 (N_4311,N_3778,N_3828);
nor U4312 (N_4312,N_3500,N_3668);
and U4313 (N_4313,N_3208,N_3403);
nand U4314 (N_4314,N_3633,N_3230);
and U4315 (N_4315,N_3835,N_3350);
nand U4316 (N_4316,N_3057,N_3330);
and U4317 (N_4317,N_3195,N_3049);
xor U4318 (N_4318,N_3718,N_3137);
nor U4319 (N_4319,N_3196,N_3510);
nand U4320 (N_4320,N_3240,N_3274);
and U4321 (N_4321,N_3130,N_3760);
nor U4322 (N_4322,N_3381,N_3644);
xor U4323 (N_4323,N_3040,N_3881);
nor U4324 (N_4324,N_3433,N_3155);
and U4325 (N_4325,N_3014,N_3364);
nand U4326 (N_4326,N_3939,N_3331);
and U4327 (N_4327,N_3926,N_3870);
or U4328 (N_4328,N_3251,N_3944);
xor U4329 (N_4329,N_3171,N_3356);
or U4330 (N_4330,N_3814,N_3450);
and U4331 (N_4331,N_3534,N_3410);
xnor U4332 (N_4332,N_3441,N_3549);
or U4333 (N_4333,N_3765,N_3925);
and U4334 (N_4334,N_3297,N_3308);
or U4335 (N_4335,N_3294,N_3642);
xnor U4336 (N_4336,N_3375,N_3554);
or U4337 (N_4337,N_3316,N_3746);
or U4338 (N_4338,N_3629,N_3555);
nor U4339 (N_4339,N_3967,N_3031);
and U4340 (N_4340,N_3891,N_3728);
nor U4341 (N_4341,N_3124,N_3705);
xor U4342 (N_4342,N_3727,N_3630);
nand U4343 (N_4343,N_3111,N_3248);
nand U4344 (N_4344,N_3504,N_3687);
or U4345 (N_4345,N_3849,N_3448);
and U4346 (N_4346,N_3136,N_3050);
xor U4347 (N_4347,N_3920,N_3605);
nand U4348 (N_4348,N_3526,N_3861);
or U4349 (N_4349,N_3197,N_3255);
or U4350 (N_4350,N_3012,N_3863);
or U4351 (N_4351,N_3935,N_3823);
nor U4352 (N_4352,N_3571,N_3080);
and U4353 (N_4353,N_3163,N_3557);
nor U4354 (N_4354,N_3567,N_3741);
nor U4355 (N_4355,N_3497,N_3929);
xnor U4356 (N_4356,N_3034,N_3981);
nand U4357 (N_4357,N_3985,N_3177);
or U4358 (N_4358,N_3135,N_3243);
nor U4359 (N_4359,N_3043,N_3337);
nor U4360 (N_4360,N_3699,N_3982);
xor U4361 (N_4361,N_3085,N_3976);
xnor U4362 (N_4362,N_3652,N_3370);
nand U4363 (N_4363,N_3664,N_3974);
and U4364 (N_4364,N_3327,N_3852);
nand U4365 (N_4365,N_3443,N_3655);
xnor U4366 (N_4366,N_3326,N_3413);
nor U4367 (N_4367,N_3273,N_3551);
nor U4368 (N_4368,N_3154,N_3169);
or U4369 (N_4369,N_3335,N_3486);
nor U4370 (N_4370,N_3953,N_3688);
nand U4371 (N_4371,N_3461,N_3755);
nand U4372 (N_4372,N_3018,N_3730);
nand U4373 (N_4373,N_3397,N_3836);
nor U4374 (N_4374,N_3300,N_3678);
and U4375 (N_4375,N_3253,N_3045);
nand U4376 (N_4376,N_3386,N_3530);
or U4377 (N_4377,N_3385,N_3284);
xor U4378 (N_4378,N_3676,N_3731);
nor U4379 (N_4379,N_3024,N_3405);
xor U4380 (N_4380,N_3709,N_3735);
or U4381 (N_4381,N_3100,N_3466);
xnor U4382 (N_4382,N_3839,N_3479);
nand U4383 (N_4383,N_3585,N_3359);
or U4384 (N_4384,N_3533,N_3096);
xor U4385 (N_4385,N_3710,N_3586);
and U4386 (N_4386,N_3594,N_3919);
nor U4387 (N_4387,N_3315,N_3145);
xnor U4388 (N_4388,N_3271,N_3880);
and U4389 (N_4389,N_3915,N_3990);
or U4390 (N_4390,N_3506,N_3844);
nand U4391 (N_4391,N_3125,N_3083);
and U4392 (N_4392,N_3099,N_3317);
xnor U4393 (N_4393,N_3215,N_3117);
xor U4394 (N_4394,N_3831,N_3886);
xor U4395 (N_4395,N_3345,N_3161);
or U4396 (N_4396,N_3363,N_3110);
nor U4397 (N_4397,N_3395,N_3245);
xnor U4398 (N_4398,N_3104,N_3449);
and U4399 (N_4399,N_3373,N_3295);
or U4400 (N_4400,N_3951,N_3296);
or U4401 (N_4401,N_3588,N_3396);
nor U4402 (N_4402,N_3930,N_3339);
xnor U4403 (N_4403,N_3569,N_3906);
or U4404 (N_4404,N_3418,N_3960);
and U4405 (N_4405,N_3608,N_3801);
nor U4406 (N_4406,N_3595,N_3860);
and U4407 (N_4407,N_3978,N_3000);
or U4408 (N_4408,N_3453,N_3142);
or U4409 (N_4409,N_3536,N_3485);
xnor U4410 (N_4410,N_3568,N_3259);
nand U4411 (N_4411,N_3559,N_3563);
nor U4412 (N_4412,N_3697,N_3051);
or U4413 (N_4413,N_3055,N_3670);
or U4414 (N_4414,N_3521,N_3458);
xor U4415 (N_4415,N_3890,N_3129);
or U4416 (N_4416,N_3573,N_3593);
and U4417 (N_4417,N_3656,N_3895);
or U4418 (N_4418,N_3813,N_3649);
and U4419 (N_4419,N_3969,N_3390);
or U4420 (N_4420,N_3862,N_3016);
nor U4421 (N_4421,N_3887,N_3477);
and U4422 (N_4422,N_3481,N_3684);
or U4423 (N_4423,N_3621,N_3948);
nand U4424 (N_4424,N_3994,N_3552);
nor U4425 (N_4425,N_3794,N_3628);
nor U4426 (N_4426,N_3868,N_3717);
xnor U4427 (N_4427,N_3487,N_3993);
nor U4428 (N_4428,N_3650,N_3622);
nand U4429 (N_4429,N_3425,N_3779);
nand U4430 (N_4430,N_3581,N_3541);
xnor U4431 (N_4431,N_3620,N_3675);
nor U4432 (N_4432,N_3003,N_3379);
or U4433 (N_4433,N_3519,N_3716);
and U4434 (N_4434,N_3574,N_3680);
nand U4435 (N_4435,N_3298,N_3972);
nor U4436 (N_4436,N_3157,N_3492);
or U4437 (N_4437,N_3798,N_3217);
nand U4438 (N_4438,N_3056,N_3984);
nor U4439 (N_4439,N_3840,N_3156);
xor U4440 (N_4440,N_3089,N_3007);
nand U4441 (N_4441,N_3989,N_3795);
and U4442 (N_4442,N_3090,N_3663);
or U4443 (N_4443,N_3250,N_3291);
xor U4444 (N_4444,N_3409,N_3102);
xor U4445 (N_4445,N_3646,N_3357);
xnor U4446 (N_4446,N_3027,N_3239);
nor U4447 (N_4447,N_3249,N_3927);
or U4448 (N_4448,N_3282,N_3015);
and U4449 (N_4449,N_3103,N_3338);
xnor U4450 (N_4450,N_3659,N_3304);
xor U4451 (N_4451,N_3164,N_3343);
or U4452 (N_4452,N_3393,N_3039);
nand U4453 (N_4453,N_3225,N_3584);
nand U4454 (N_4454,N_3404,N_3832);
xor U4455 (N_4455,N_3010,N_3829);
xor U4456 (N_4456,N_3321,N_3694);
nand U4457 (N_4457,N_3334,N_3180);
xor U4458 (N_4458,N_3309,N_3198);
and U4459 (N_4459,N_3322,N_3462);
and U4460 (N_4460,N_3340,N_3445);
nand U4461 (N_4461,N_3131,N_3871);
and U4462 (N_4462,N_3004,N_3942);
xor U4463 (N_4463,N_3783,N_3172);
nor U4464 (N_4464,N_3873,N_3713);
xor U4465 (N_4465,N_3323,N_3360);
nor U4466 (N_4466,N_3789,N_3700);
nand U4467 (N_4467,N_3221,N_3665);
nand U4468 (N_4468,N_3301,N_3695);
and U4469 (N_4469,N_3224,N_3319);
nor U4470 (N_4470,N_3182,N_3442);
nand U4471 (N_4471,N_3460,N_3885);
nand U4472 (N_4472,N_3048,N_3723);
and U4473 (N_4473,N_3842,N_3786);
or U4474 (N_4474,N_3219,N_3174);
nor U4475 (N_4475,N_3520,N_3199);
or U4476 (N_4476,N_3987,N_3400);
nor U4477 (N_4477,N_3170,N_3875);
or U4478 (N_4478,N_3332,N_3998);
and U4479 (N_4479,N_3216,N_3203);
nand U4480 (N_4480,N_3992,N_3498);
or U4481 (N_4481,N_3499,N_3609);
xnor U4482 (N_4482,N_3312,N_3525);
and U4483 (N_4483,N_3722,N_3946);
nor U4484 (N_4484,N_3931,N_3422);
xor U4485 (N_4485,N_3355,N_3127);
nor U4486 (N_4486,N_3150,N_3392);
nor U4487 (N_4487,N_3463,N_3734);
and U4488 (N_4488,N_3833,N_3093);
or U4489 (N_4489,N_3101,N_3928);
and U4490 (N_4490,N_3970,N_3138);
nor U4491 (N_4491,N_3516,N_3491);
or U4492 (N_4492,N_3178,N_3365);
or U4493 (N_4493,N_3800,N_3815);
nor U4494 (N_4494,N_3143,N_3280);
xor U4495 (N_4495,N_3120,N_3351);
nand U4496 (N_4496,N_3796,N_3496);
nand U4497 (N_4497,N_3672,N_3070);
nor U4498 (N_4498,N_3063,N_3780);
or U4499 (N_4499,N_3490,N_3329);
nand U4500 (N_4500,N_3678,N_3091);
nand U4501 (N_4501,N_3585,N_3233);
nand U4502 (N_4502,N_3012,N_3177);
and U4503 (N_4503,N_3612,N_3573);
or U4504 (N_4504,N_3667,N_3571);
nand U4505 (N_4505,N_3464,N_3482);
xnor U4506 (N_4506,N_3760,N_3552);
and U4507 (N_4507,N_3610,N_3518);
xor U4508 (N_4508,N_3200,N_3269);
and U4509 (N_4509,N_3079,N_3621);
or U4510 (N_4510,N_3322,N_3851);
and U4511 (N_4511,N_3085,N_3780);
nor U4512 (N_4512,N_3849,N_3275);
nand U4513 (N_4513,N_3986,N_3241);
or U4514 (N_4514,N_3245,N_3493);
and U4515 (N_4515,N_3264,N_3999);
or U4516 (N_4516,N_3840,N_3886);
or U4517 (N_4517,N_3934,N_3037);
or U4518 (N_4518,N_3598,N_3356);
and U4519 (N_4519,N_3884,N_3752);
or U4520 (N_4520,N_3961,N_3701);
and U4521 (N_4521,N_3484,N_3218);
and U4522 (N_4522,N_3711,N_3092);
and U4523 (N_4523,N_3106,N_3671);
or U4524 (N_4524,N_3203,N_3418);
and U4525 (N_4525,N_3031,N_3182);
nor U4526 (N_4526,N_3350,N_3942);
and U4527 (N_4527,N_3179,N_3010);
xor U4528 (N_4528,N_3000,N_3020);
xnor U4529 (N_4529,N_3389,N_3869);
xor U4530 (N_4530,N_3827,N_3003);
xnor U4531 (N_4531,N_3102,N_3998);
xor U4532 (N_4532,N_3108,N_3378);
xnor U4533 (N_4533,N_3616,N_3790);
nor U4534 (N_4534,N_3499,N_3703);
nor U4535 (N_4535,N_3050,N_3889);
and U4536 (N_4536,N_3046,N_3293);
nor U4537 (N_4537,N_3765,N_3233);
nand U4538 (N_4538,N_3127,N_3881);
nand U4539 (N_4539,N_3206,N_3771);
nand U4540 (N_4540,N_3329,N_3966);
xnor U4541 (N_4541,N_3466,N_3030);
nor U4542 (N_4542,N_3689,N_3031);
xnor U4543 (N_4543,N_3451,N_3524);
nand U4544 (N_4544,N_3166,N_3836);
nand U4545 (N_4545,N_3972,N_3957);
nor U4546 (N_4546,N_3610,N_3463);
nand U4547 (N_4547,N_3052,N_3080);
nor U4548 (N_4548,N_3301,N_3256);
xor U4549 (N_4549,N_3514,N_3630);
xnor U4550 (N_4550,N_3937,N_3714);
and U4551 (N_4551,N_3695,N_3310);
and U4552 (N_4552,N_3856,N_3275);
or U4553 (N_4553,N_3661,N_3575);
and U4554 (N_4554,N_3067,N_3290);
nor U4555 (N_4555,N_3408,N_3925);
xor U4556 (N_4556,N_3487,N_3537);
xor U4557 (N_4557,N_3569,N_3498);
and U4558 (N_4558,N_3250,N_3986);
or U4559 (N_4559,N_3368,N_3178);
or U4560 (N_4560,N_3112,N_3282);
or U4561 (N_4561,N_3543,N_3625);
nor U4562 (N_4562,N_3967,N_3461);
xnor U4563 (N_4563,N_3344,N_3519);
nand U4564 (N_4564,N_3758,N_3219);
and U4565 (N_4565,N_3057,N_3118);
or U4566 (N_4566,N_3964,N_3160);
or U4567 (N_4567,N_3270,N_3282);
and U4568 (N_4568,N_3862,N_3522);
nor U4569 (N_4569,N_3709,N_3402);
nand U4570 (N_4570,N_3707,N_3630);
and U4571 (N_4571,N_3219,N_3292);
and U4572 (N_4572,N_3447,N_3245);
and U4573 (N_4573,N_3005,N_3062);
nor U4574 (N_4574,N_3114,N_3972);
and U4575 (N_4575,N_3114,N_3297);
nand U4576 (N_4576,N_3033,N_3298);
nor U4577 (N_4577,N_3463,N_3501);
xnor U4578 (N_4578,N_3740,N_3756);
xnor U4579 (N_4579,N_3273,N_3836);
nand U4580 (N_4580,N_3979,N_3354);
nand U4581 (N_4581,N_3524,N_3141);
or U4582 (N_4582,N_3419,N_3276);
nor U4583 (N_4583,N_3570,N_3863);
nor U4584 (N_4584,N_3047,N_3942);
nor U4585 (N_4585,N_3197,N_3228);
nand U4586 (N_4586,N_3156,N_3928);
nand U4587 (N_4587,N_3978,N_3275);
or U4588 (N_4588,N_3962,N_3782);
and U4589 (N_4589,N_3186,N_3633);
nand U4590 (N_4590,N_3123,N_3831);
and U4591 (N_4591,N_3725,N_3098);
and U4592 (N_4592,N_3571,N_3614);
and U4593 (N_4593,N_3574,N_3784);
nor U4594 (N_4594,N_3826,N_3300);
nand U4595 (N_4595,N_3854,N_3947);
or U4596 (N_4596,N_3723,N_3976);
and U4597 (N_4597,N_3260,N_3820);
and U4598 (N_4598,N_3392,N_3292);
nand U4599 (N_4599,N_3022,N_3863);
nor U4600 (N_4600,N_3432,N_3756);
and U4601 (N_4601,N_3991,N_3622);
nor U4602 (N_4602,N_3268,N_3267);
nor U4603 (N_4603,N_3627,N_3002);
or U4604 (N_4604,N_3927,N_3425);
xnor U4605 (N_4605,N_3045,N_3381);
nand U4606 (N_4606,N_3789,N_3833);
nand U4607 (N_4607,N_3524,N_3522);
or U4608 (N_4608,N_3228,N_3819);
nand U4609 (N_4609,N_3845,N_3001);
xnor U4610 (N_4610,N_3505,N_3057);
nand U4611 (N_4611,N_3043,N_3879);
xor U4612 (N_4612,N_3230,N_3828);
nand U4613 (N_4613,N_3384,N_3107);
xnor U4614 (N_4614,N_3396,N_3054);
or U4615 (N_4615,N_3049,N_3071);
or U4616 (N_4616,N_3515,N_3280);
and U4617 (N_4617,N_3833,N_3319);
or U4618 (N_4618,N_3081,N_3385);
nand U4619 (N_4619,N_3145,N_3640);
and U4620 (N_4620,N_3609,N_3870);
xnor U4621 (N_4621,N_3724,N_3869);
and U4622 (N_4622,N_3285,N_3158);
nand U4623 (N_4623,N_3406,N_3054);
nor U4624 (N_4624,N_3683,N_3330);
and U4625 (N_4625,N_3722,N_3312);
nand U4626 (N_4626,N_3107,N_3883);
nor U4627 (N_4627,N_3370,N_3718);
and U4628 (N_4628,N_3108,N_3298);
nor U4629 (N_4629,N_3108,N_3049);
or U4630 (N_4630,N_3491,N_3580);
xnor U4631 (N_4631,N_3596,N_3537);
nor U4632 (N_4632,N_3052,N_3099);
xor U4633 (N_4633,N_3774,N_3295);
or U4634 (N_4634,N_3003,N_3531);
xor U4635 (N_4635,N_3585,N_3966);
and U4636 (N_4636,N_3357,N_3305);
nand U4637 (N_4637,N_3931,N_3616);
nand U4638 (N_4638,N_3709,N_3475);
nand U4639 (N_4639,N_3585,N_3682);
or U4640 (N_4640,N_3394,N_3364);
or U4641 (N_4641,N_3129,N_3917);
and U4642 (N_4642,N_3058,N_3552);
nand U4643 (N_4643,N_3828,N_3531);
nand U4644 (N_4644,N_3735,N_3469);
nand U4645 (N_4645,N_3818,N_3666);
xor U4646 (N_4646,N_3950,N_3291);
and U4647 (N_4647,N_3561,N_3229);
nand U4648 (N_4648,N_3626,N_3563);
nand U4649 (N_4649,N_3004,N_3818);
nor U4650 (N_4650,N_3652,N_3931);
xnor U4651 (N_4651,N_3428,N_3745);
and U4652 (N_4652,N_3432,N_3021);
nor U4653 (N_4653,N_3978,N_3839);
xor U4654 (N_4654,N_3888,N_3745);
xor U4655 (N_4655,N_3194,N_3153);
or U4656 (N_4656,N_3042,N_3005);
or U4657 (N_4657,N_3389,N_3998);
xor U4658 (N_4658,N_3058,N_3419);
and U4659 (N_4659,N_3566,N_3859);
xor U4660 (N_4660,N_3023,N_3450);
or U4661 (N_4661,N_3224,N_3318);
and U4662 (N_4662,N_3231,N_3880);
or U4663 (N_4663,N_3689,N_3597);
nand U4664 (N_4664,N_3442,N_3350);
xnor U4665 (N_4665,N_3958,N_3441);
and U4666 (N_4666,N_3725,N_3216);
nand U4667 (N_4667,N_3656,N_3759);
nor U4668 (N_4668,N_3225,N_3474);
and U4669 (N_4669,N_3924,N_3878);
and U4670 (N_4670,N_3207,N_3405);
or U4671 (N_4671,N_3669,N_3776);
xor U4672 (N_4672,N_3367,N_3488);
and U4673 (N_4673,N_3371,N_3249);
xnor U4674 (N_4674,N_3596,N_3825);
nand U4675 (N_4675,N_3373,N_3389);
nor U4676 (N_4676,N_3053,N_3516);
xnor U4677 (N_4677,N_3891,N_3906);
nor U4678 (N_4678,N_3849,N_3369);
and U4679 (N_4679,N_3438,N_3115);
nand U4680 (N_4680,N_3706,N_3533);
nor U4681 (N_4681,N_3317,N_3389);
and U4682 (N_4682,N_3872,N_3120);
and U4683 (N_4683,N_3008,N_3859);
nand U4684 (N_4684,N_3814,N_3890);
or U4685 (N_4685,N_3753,N_3461);
xor U4686 (N_4686,N_3059,N_3112);
nand U4687 (N_4687,N_3878,N_3441);
nand U4688 (N_4688,N_3516,N_3587);
nor U4689 (N_4689,N_3485,N_3269);
nor U4690 (N_4690,N_3267,N_3126);
and U4691 (N_4691,N_3864,N_3220);
and U4692 (N_4692,N_3035,N_3334);
nor U4693 (N_4693,N_3197,N_3561);
or U4694 (N_4694,N_3029,N_3997);
and U4695 (N_4695,N_3605,N_3855);
xor U4696 (N_4696,N_3216,N_3764);
nand U4697 (N_4697,N_3595,N_3609);
xor U4698 (N_4698,N_3957,N_3034);
and U4699 (N_4699,N_3694,N_3897);
and U4700 (N_4700,N_3454,N_3209);
nand U4701 (N_4701,N_3485,N_3170);
nand U4702 (N_4702,N_3133,N_3983);
and U4703 (N_4703,N_3487,N_3841);
nand U4704 (N_4704,N_3326,N_3561);
or U4705 (N_4705,N_3099,N_3736);
xor U4706 (N_4706,N_3952,N_3827);
and U4707 (N_4707,N_3193,N_3266);
xor U4708 (N_4708,N_3096,N_3592);
or U4709 (N_4709,N_3499,N_3057);
nand U4710 (N_4710,N_3632,N_3975);
xnor U4711 (N_4711,N_3825,N_3758);
or U4712 (N_4712,N_3777,N_3263);
xor U4713 (N_4713,N_3664,N_3638);
and U4714 (N_4714,N_3648,N_3394);
xnor U4715 (N_4715,N_3126,N_3108);
and U4716 (N_4716,N_3682,N_3673);
and U4717 (N_4717,N_3237,N_3252);
and U4718 (N_4718,N_3861,N_3047);
and U4719 (N_4719,N_3003,N_3310);
xor U4720 (N_4720,N_3490,N_3916);
nor U4721 (N_4721,N_3329,N_3755);
or U4722 (N_4722,N_3242,N_3830);
and U4723 (N_4723,N_3831,N_3251);
and U4724 (N_4724,N_3307,N_3696);
and U4725 (N_4725,N_3360,N_3454);
or U4726 (N_4726,N_3669,N_3300);
nand U4727 (N_4727,N_3426,N_3682);
nand U4728 (N_4728,N_3549,N_3621);
nor U4729 (N_4729,N_3456,N_3975);
or U4730 (N_4730,N_3141,N_3931);
or U4731 (N_4731,N_3501,N_3564);
and U4732 (N_4732,N_3541,N_3009);
xor U4733 (N_4733,N_3490,N_3683);
or U4734 (N_4734,N_3247,N_3264);
nor U4735 (N_4735,N_3207,N_3112);
or U4736 (N_4736,N_3906,N_3849);
nor U4737 (N_4737,N_3271,N_3205);
xor U4738 (N_4738,N_3280,N_3409);
nor U4739 (N_4739,N_3393,N_3351);
nor U4740 (N_4740,N_3559,N_3526);
nand U4741 (N_4741,N_3698,N_3604);
xor U4742 (N_4742,N_3323,N_3785);
or U4743 (N_4743,N_3482,N_3833);
nand U4744 (N_4744,N_3928,N_3577);
nor U4745 (N_4745,N_3734,N_3529);
and U4746 (N_4746,N_3826,N_3123);
nor U4747 (N_4747,N_3434,N_3554);
xnor U4748 (N_4748,N_3227,N_3318);
nor U4749 (N_4749,N_3975,N_3689);
and U4750 (N_4750,N_3029,N_3247);
nand U4751 (N_4751,N_3654,N_3614);
nand U4752 (N_4752,N_3671,N_3504);
and U4753 (N_4753,N_3313,N_3814);
or U4754 (N_4754,N_3316,N_3138);
nand U4755 (N_4755,N_3046,N_3198);
or U4756 (N_4756,N_3433,N_3236);
or U4757 (N_4757,N_3520,N_3879);
xor U4758 (N_4758,N_3849,N_3821);
and U4759 (N_4759,N_3672,N_3778);
or U4760 (N_4760,N_3057,N_3667);
xor U4761 (N_4761,N_3534,N_3366);
or U4762 (N_4762,N_3603,N_3931);
or U4763 (N_4763,N_3157,N_3971);
nor U4764 (N_4764,N_3954,N_3545);
xor U4765 (N_4765,N_3485,N_3722);
or U4766 (N_4766,N_3812,N_3997);
nand U4767 (N_4767,N_3975,N_3588);
xor U4768 (N_4768,N_3557,N_3106);
nor U4769 (N_4769,N_3462,N_3417);
xor U4770 (N_4770,N_3522,N_3930);
xor U4771 (N_4771,N_3591,N_3436);
and U4772 (N_4772,N_3632,N_3311);
and U4773 (N_4773,N_3958,N_3218);
nand U4774 (N_4774,N_3568,N_3559);
and U4775 (N_4775,N_3916,N_3446);
nand U4776 (N_4776,N_3092,N_3088);
nand U4777 (N_4777,N_3535,N_3080);
xor U4778 (N_4778,N_3252,N_3054);
nor U4779 (N_4779,N_3570,N_3563);
and U4780 (N_4780,N_3206,N_3304);
or U4781 (N_4781,N_3127,N_3825);
nor U4782 (N_4782,N_3843,N_3203);
and U4783 (N_4783,N_3743,N_3480);
nand U4784 (N_4784,N_3528,N_3253);
and U4785 (N_4785,N_3005,N_3564);
or U4786 (N_4786,N_3347,N_3774);
and U4787 (N_4787,N_3032,N_3556);
nand U4788 (N_4788,N_3937,N_3415);
or U4789 (N_4789,N_3663,N_3940);
and U4790 (N_4790,N_3155,N_3418);
or U4791 (N_4791,N_3375,N_3639);
or U4792 (N_4792,N_3748,N_3049);
and U4793 (N_4793,N_3156,N_3020);
or U4794 (N_4794,N_3550,N_3596);
xnor U4795 (N_4795,N_3353,N_3832);
and U4796 (N_4796,N_3313,N_3377);
nor U4797 (N_4797,N_3771,N_3024);
xor U4798 (N_4798,N_3186,N_3998);
or U4799 (N_4799,N_3362,N_3244);
nor U4800 (N_4800,N_3934,N_3437);
and U4801 (N_4801,N_3613,N_3597);
and U4802 (N_4802,N_3860,N_3377);
nor U4803 (N_4803,N_3642,N_3146);
or U4804 (N_4804,N_3893,N_3143);
xor U4805 (N_4805,N_3442,N_3186);
xnor U4806 (N_4806,N_3260,N_3190);
or U4807 (N_4807,N_3775,N_3582);
xnor U4808 (N_4808,N_3524,N_3383);
or U4809 (N_4809,N_3147,N_3530);
xnor U4810 (N_4810,N_3744,N_3154);
nand U4811 (N_4811,N_3058,N_3959);
nand U4812 (N_4812,N_3358,N_3708);
nand U4813 (N_4813,N_3755,N_3688);
nor U4814 (N_4814,N_3581,N_3658);
xor U4815 (N_4815,N_3440,N_3901);
or U4816 (N_4816,N_3345,N_3961);
xor U4817 (N_4817,N_3298,N_3303);
xnor U4818 (N_4818,N_3965,N_3712);
nor U4819 (N_4819,N_3584,N_3382);
xnor U4820 (N_4820,N_3180,N_3795);
and U4821 (N_4821,N_3697,N_3589);
and U4822 (N_4822,N_3494,N_3650);
nand U4823 (N_4823,N_3153,N_3618);
or U4824 (N_4824,N_3460,N_3640);
nor U4825 (N_4825,N_3629,N_3403);
nand U4826 (N_4826,N_3212,N_3653);
and U4827 (N_4827,N_3870,N_3994);
or U4828 (N_4828,N_3109,N_3943);
or U4829 (N_4829,N_3538,N_3633);
nand U4830 (N_4830,N_3508,N_3134);
nor U4831 (N_4831,N_3785,N_3923);
nand U4832 (N_4832,N_3331,N_3739);
or U4833 (N_4833,N_3823,N_3896);
or U4834 (N_4834,N_3373,N_3892);
and U4835 (N_4835,N_3845,N_3579);
and U4836 (N_4836,N_3557,N_3034);
or U4837 (N_4837,N_3377,N_3063);
nand U4838 (N_4838,N_3194,N_3182);
nand U4839 (N_4839,N_3834,N_3049);
nor U4840 (N_4840,N_3875,N_3121);
nand U4841 (N_4841,N_3064,N_3721);
or U4842 (N_4842,N_3123,N_3745);
nand U4843 (N_4843,N_3219,N_3325);
or U4844 (N_4844,N_3029,N_3708);
nor U4845 (N_4845,N_3187,N_3168);
nand U4846 (N_4846,N_3166,N_3328);
or U4847 (N_4847,N_3591,N_3434);
xnor U4848 (N_4848,N_3079,N_3374);
or U4849 (N_4849,N_3300,N_3160);
xnor U4850 (N_4850,N_3194,N_3539);
or U4851 (N_4851,N_3898,N_3118);
nand U4852 (N_4852,N_3233,N_3535);
or U4853 (N_4853,N_3820,N_3188);
nand U4854 (N_4854,N_3767,N_3322);
xnor U4855 (N_4855,N_3516,N_3822);
or U4856 (N_4856,N_3807,N_3150);
or U4857 (N_4857,N_3191,N_3078);
or U4858 (N_4858,N_3623,N_3154);
and U4859 (N_4859,N_3074,N_3658);
nand U4860 (N_4860,N_3413,N_3795);
nor U4861 (N_4861,N_3807,N_3146);
and U4862 (N_4862,N_3356,N_3835);
and U4863 (N_4863,N_3437,N_3246);
and U4864 (N_4864,N_3627,N_3959);
nor U4865 (N_4865,N_3665,N_3705);
nand U4866 (N_4866,N_3748,N_3175);
xnor U4867 (N_4867,N_3905,N_3603);
or U4868 (N_4868,N_3014,N_3900);
or U4869 (N_4869,N_3303,N_3495);
and U4870 (N_4870,N_3861,N_3116);
nor U4871 (N_4871,N_3184,N_3913);
or U4872 (N_4872,N_3072,N_3477);
nor U4873 (N_4873,N_3770,N_3427);
xnor U4874 (N_4874,N_3288,N_3062);
and U4875 (N_4875,N_3184,N_3158);
and U4876 (N_4876,N_3830,N_3588);
nor U4877 (N_4877,N_3678,N_3724);
or U4878 (N_4878,N_3993,N_3703);
xnor U4879 (N_4879,N_3165,N_3238);
and U4880 (N_4880,N_3935,N_3383);
or U4881 (N_4881,N_3855,N_3554);
nor U4882 (N_4882,N_3470,N_3915);
nand U4883 (N_4883,N_3106,N_3080);
nand U4884 (N_4884,N_3871,N_3122);
or U4885 (N_4885,N_3271,N_3153);
or U4886 (N_4886,N_3146,N_3927);
and U4887 (N_4887,N_3888,N_3278);
and U4888 (N_4888,N_3462,N_3315);
xor U4889 (N_4889,N_3501,N_3269);
nand U4890 (N_4890,N_3994,N_3586);
and U4891 (N_4891,N_3029,N_3122);
and U4892 (N_4892,N_3801,N_3755);
xor U4893 (N_4893,N_3295,N_3930);
nor U4894 (N_4894,N_3166,N_3171);
and U4895 (N_4895,N_3622,N_3001);
or U4896 (N_4896,N_3958,N_3701);
nor U4897 (N_4897,N_3871,N_3920);
and U4898 (N_4898,N_3715,N_3542);
nand U4899 (N_4899,N_3891,N_3698);
nor U4900 (N_4900,N_3155,N_3781);
nor U4901 (N_4901,N_3996,N_3550);
nor U4902 (N_4902,N_3834,N_3638);
nand U4903 (N_4903,N_3712,N_3276);
nand U4904 (N_4904,N_3085,N_3662);
or U4905 (N_4905,N_3774,N_3013);
or U4906 (N_4906,N_3261,N_3905);
xnor U4907 (N_4907,N_3360,N_3253);
and U4908 (N_4908,N_3511,N_3589);
nor U4909 (N_4909,N_3635,N_3845);
xor U4910 (N_4910,N_3254,N_3043);
nand U4911 (N_4911,N_3237,N_3529);
nor U4912 (N_4912,N_3899,N_3291);
nor U4913 (N_4913,N_3319,N_3997);
nor U4914 (N_4914,N_3351,N_3489);
xor U4915 (N_4915,N_3602,N_3355);
and U4916 (N_4916,N_3340,N_3327);
nand U4917 (N_4917,N_3544,N_3957);
nor U4918 (N_4918,N_3162,N_3616);
nor U4919 (N_4919,N_3057,N_3343);
xor U4920 (N_4920,N_3260,N_3657);
nor U4921 (N_4921,N_3545,N_3671);
and U4922 (N_4922,N_3717,N_3095);
and U4923 (N_4923,N_3479,N_3475);
and U4924 (N_4924,N_3262,N_3278);
nor U4925 (N_4925,N_3542,N_3096);
and U4926 (N_4926,N_3263,N_3030);
nor U4927 (N_4927,N_3663,N_3450);
nor U4928 (N_4928,N_3876,N_3888);
xnor U4929 (N_4929,N_3932,N_3258);
nor U4930 (N_4930,N_3414,N_3534);
or U4931 (N_4931,N_3816,N_3125);
nand U4932 (N_4932,N_3168,N_3175);
nor U4933 (N_4933,N_3783,N_3484);
or U4934 (N_4934,N_3341,N_3467);
nor U4935 (N_4935,N_3528,N_3031);
nor U4936 (N_4936,N_3284,N_3914);
nand U4937 (N_4937,N_3291,N_3394);
or U4938 (N_4938,N_3293,N_3872);
or U4939 (N_4939,N_3464,N_3709);
nand U4940 (N_4940,N_3852,N_3924);
nand U4941 (N_4941,N_3018,N_3514);
nand U4942 (N_4942,N_3855,N_3353);
nand U4943 (N_4943,N_3164,N_3538);
and U4944 (N_4944,N_3608,N_3533);
xor U4945 (N_4945,N_3976,N_3973);
xnor U4946 (N_4946,N_3371,N_3922);
or U4947 (N_4947,N_3733,N_3133);
and U4948 (N_4948,N_3137,N_3203);
xor U4949 (N_4949,N_3474,N_3680);
xor U4950 (N_4950,N_3684,N_3350);
xnor U4951 (N_4951,N_3356,N_3510);
xnor U4952 (N_4952,N_3551,N_3473);
xor U4953 (N_4953,N_3099,N_3224);
and U4954 (N_4954,N_3330,N_3686);
or U4955 (N_4955,N_3548,N_3409);
nand U4956 (N_4956,N_3038,N_3059);
xnor U4957 (N_4957,N_3864,N_3884);
or U4958 (N_4958,N_3545,N_3558);
and U4959 (N_4959,N_3670,N_3559);
xnor U4960 (N_4960,N_3817,N_3122);
and U4961 (N_4961,N_3923,N_3714);
xor U4962 (N_4962,N_3261,N_3671);
nor U4963 (N_4963,N_3361,N_3148);
or U4964 (N_4964,N_3996,N_3564);
and U4965 (N_4965,N_3538,N_3061);
and U4966 (N_4966,N_3939,N_3070);
xnor U4967 (N_4967,N_3954,N_3246);
xnor U4968 (N_4968,N_3612,N_3428);
xor U4969 (N_4969,N_3715,N_3976);
xor U4970 (N_4970,N_3202,N_3918);
nand U4971 (N_4971,N_3918,N_3707);
and U4972 (N_4972,N_3931,N_3721);
xor U4973 (N_4973,N_3358,N_3056);
nor U4974 (N_4974,N_3700,N_3619);
nand U4975 (N_4975,N_3399,N_3511);
xnor U4976 (N_4976,N_3355,N_3409);
nand U4977 (N_4977,N_3467,N_3767);
or U4978 (N_4978,N_3152,N_3868);
or U4979 (N_4979,N_3779,N_3793);
nor U4980 (N_4980,N_3265,N_3773);
nor U4981 (N_4981,N_3483,N_3563);
and U4982 (N_4982,N_3760,N_3125);
nand U4983 (N_4983,N_3342,N_3430);
or U4984 (N_4984,N_3063,N_3349);
nand U4985 (N_4985,N_3873,N_3254);
or U4986 (N_4986,N_3066,N_3774);
or U4987 (N_4987,N_3363,N_3983);
nand U4988 (N_4988,N_3406,N_3152);
xnor U4989 (N_4989,N_3323,N_3345);
or U4990 (N_4990,N_3639,N_3134);
nand U4991 (N_4991,N_3232,N_3945);
and U4992 (N_4992,N_3686,N_3881);
or U4993 (N_4993,N_3099,N_3591);
or U4994 (N_4994,N_3572,N_3552);
xnor U4995 (N_4995,N_3106,N_3924);
nand U4996 (N_4996,N_3014,N_3318);
and U4997 (N_4997,N_3025,N_3035);
xor U4998 (N_4998,N_3001,N_3699);
nor U4999 (N_4999,N_3695,N_3977);
and U5000 (N_5000,N_4390,N_4075);
nor U5001 (N_5001,N_4443,N_4363);
xnor U5002 (N_5002,N_4810,N_4392);
nor U5003 (N_5003,N_4862,N_4701);
and U5004 (N_5004,N_4560,N_4345);
or U5005 (N_5005,N_4239,N_4680);
nand U5006 (N_5006,N_4347,N_4625);
xnor U5007 (N_5007,N_4951,N_4140);
nand U5008 (N_5008,N_4284,N_4935);
and U5009 (N_5009,N_4681,N_4070);
or U5010 (N_5010,N_4134,N_4520);
xor U5011 (N_5011,N_4992,N_4342);
nand U5012 (N_5012,N_4455,N_4203);
xnor U5013 (N_5013,N_4381,N_4469);
nor U5014 (N_5014,N_4216,N_4290);
and U5015 (N_5015,N_4404,N_4730);
or U5016 (N_5016,N_4936,N_4481);
or U5017 (N_5017,N_4424,N_4368);
or U5018 (N_5018,N_4108,N_4110);
nor U5019 (N_5019,N_4291,N_4830);
nand U5020 (N_5020,N_4444,N_4742);
or U5021 (N_5021,N_4942,N_4139);
and U5022 (N_5022,N_4036,N_4733);
or U5023 (N_5023,N_4842,N_4432);
and U5024 (N_5024,N_4006,N_4048);
nand U5025 (N_5025,N_4164,N_4557);
xnor U5026 (N_5026,N_4057,N_4780);
or U5027 (N_5027,N_4084,N_4453);
or U5028 (N_5028,N_4869,N_4043);
and U5029 (N_5029,N_4311,N_4802);
and U5030 (N_5030,N_4615,N_4235);
nand U5031 (N_5031,N_4587,N_4064);
nor U5032 (N_5032,N_4956,N_4030);
xor U5033 (N_5033,N_4369,N_4208);
xnor U5034 (N_5034,N_4083,N_4561);
or U5035 (N_5035,N_4524,N_4395);
xnor U5036 (N_5036,N_4737,N_4966);
or U5037 (N_5037,N_4771,N_4755);
nand U5038 (N_5038,N_4859,N_4867);
nand U5039 (N_5039,N_4195,N_4207);
and U5040 (N_5040,N_4371,N_4897);
and U5041 (N_5041,N_4967,N_4947);
or U5042 (N_5042,N_4971,N_4472);
xnor U5043 (N_5043,N_4653,N_4194);
or U5044 (N_5044,N_4225,N_4640);
and U5045 (N_5045,N_4712,N_4916);
or U5046 (N_5046,N_4550,N_4454);
xnor U5047 (N_5047,N_4761,N_4750);
or U5048 (N_5048,N_4421,N_4518);
nor U5049 (N_5049,N_4668,N_4637);
xor U5050 (N_5050,N_4766,N_4173);
and U5051 (N_5051,N_4768,N_4434);
nand U5052 (N_5052,N_4979,N_4344);
and U5053 (N_5053,N_4634,N_4298);
nand U5054 (N_5054,N_4868,N_4604);
nor U5055 (N_5055,N_4438,N_4969);
nor U5056 (N_5056,N_4078,N_4261);
xnor U5057 (N_5057,N_4309,N_4645);
and U5058 (N_5058,N_4873,N_4148);
nor U5059 (N_5059,N_4577,N_4321);
xor U5060 (N_5060,N_4101,N_4425);
nand U5061 (N_5061,N_4580,N_4360);
nand U5062 (N_5062,N_4820,N_4375);
nor U5063 (N_5063,N_4531,N_4315);
nor U5064 (N_5064,N_4643,N_4948);
xor U5065 (N_5065,N_4162,N_4044);
xnor U5066 (N_5066,N_4870,N_4046);
xor U5067 (N_5067,N_4541,N_4527);
nor U5068 (N_5068,N_4649,N_4813);
nor U5069 (N_5069,N_4756,N_4411);
and U5070 (N_5070,N_4970,N_4773);
xor U5071 (N_5071,N_4193,N_4609);
xnor U5072 (N_5072,N_4918,N_4274);
or U5073 (N_5073,N_4463,N_4985);
nor U5074 (N_5074,N_4686,N_4517);
and U5075 (N_5075,N_4510,N_4091);
nand U5076 (N_5076,N_4921,N_4415);
nor U5077 (N_5077,N_4166,N_4227);
or U5078 (N_5078,N_4275,N_4934);
or U5079 (N_5079,N_4707,N_4452);
or U5080 (N_5080,N_4687,N_4612);
nand U5081 (N_5081,N_4989,N_4512);
xor U5082 (N_5082,N_4703,N_4365);
xor U5083 (N_5083,N_4102,N_4198);
nor U5084 (N_5084,N_4223,N_4727);
or U5085 (N_5085,N_4350,N_4338);
or U5086 (N_5086,N_4589,N_4548);
nand U5087 (N_5087,N_4563,N_4474);
nor U5088 (N_5088,N_4984,N_4310);
or U5089 (N_5089,N_4839,N_4840);
nor U5090 (N_5090,N_4818,N_4708);
and U5091 (N_5091,N_4236,N_4807);
xnor U5092 (N_5092,N_4925,N_4117);
and U5093 (N_5093,N_4002,N_4475);
or U5094 (N_5094,N_4152,N_4220);
or U5095 (N_5095,N_4144,N_4297);
nand U5096 (N_5096,N_4762,N_4409);
or U5097 (N_5097,N_4206,N_4062);
nor U5098 (N_5098,N_4973,N_4628);
or U5099 (N_5099,N_4095,N_4549);
nor U5100 (N_5100,N_4608,N_4860);
and U5101 (N_5101,N_4927,N_4219);
nand U5102 (N_5102,N_4928,N_4808);
nand U5103 (N_5103,N_4978,N_4590);
and U5104 (N_5104,N_4187,N_4662);
xnor U5105 (N_5105,N_4564,N_4659);
or U5106 (N_5106,N_4211,N_4822);
nor U5107 (N_5107,N_4991,N_4729);
and U5108 (N_5108,N_4789,N_4702);
and U5109 (N_5109,N_4983,N_4841);
or U5110 (N_5110,N_4998,N_4210);
xnor U5111 (N_5111,N_4417,N_4156);
nand U5112 (N_5112,N_4241,N_4296);
xor U5113 (N_5113,N_4268,N_4749);
nand U5114 (N_5114,N_4535,N_4529);
nand U5115 (N_5115,N_4909,N_4570);
nor U5116 (N_5116,N_4538,N_4354);
and U5117 (N_5117,N_4081,N_4151);
xor U5118 (N_5118,N_4674,N_4184);
nand U5119 (N_5119,N_4440,N_4124);
nor U5120 (N_5120,N_4881,N_4500);
or U5121 (N_5121,N_4089,N_4059);
nor U5122 (N_5122,N_4552,N_4675);
nand U5123 (N_5123,N_4699,N_4537);
and U5124 (N_5124,N_4267,N_4571);
or U5125 (N_5125,N_4256,N_4781);
nor U5126 (N_5126,N_4805,N_4182);
and U5127 (N_5127,N_4855,N_4716);
nand U5128 (N_5128,N_4093,N_4528);
nor U5129 (N_5129,N_4126,N_4403);
and U5130 (N_5130,N_4303,N_4049);
or U5131 (N_5131,N_4846,N_4176);
nand U5132 (N_5132,N_4932,N_4950);
or U5133 (N_5133,N_4597,N_4019);
and U5134 (N_5134,N_4611,N_4283);
or U5135 (N_5135,N_4938,N_4994);
xnor U5136 (N_5136,N_4861,N_4694);
and U5137 (N_5137,N_4118,N_4719);
or U5138 (N_5138,N_4039,N_4798);
and U5139 (N_5139,N_4343,N_4300);
and U5140 (N_5140,N_4864,N_4437);
nand U5141 (N_5141,N_4278,N_4665);
xor U5142 (N_5142,N_4449,N_4063);
nor U5143 (N_5143,N_4871,N_4384);
nor U5144 (N_5144,N_4491,N_4149);
nand U5145 (N_5145,N_4367,N_4094);
nor U5146 (N_5146,N_4734,N_4397);
xor U5147 (N_5147,N_4362,N_4009);
xor U5148 (N_5148,N_4258,N_4495);
nor U5149 (N_5149,N_4904,N_4585);
nand U5150 (N_5150,N_4435,N_4451);
and U5151 (N_5151,N_4336,N_4565);
and U5152 (N_5152,N_4582,N_4460);
and U5153 (N_5153,N_4574,N_4960);
or U5154 (N_5154,N_4591,N_4185);
and U5155 (N_5155,N_4401,N_4486);
and U5156 (N_5156,N_4958,N_4010);
nor U5157 (N_5157,N_4067,N_4705);
nand U5158 (N_5158,N_4709,N_4175);
nand U5159 (N_5159,N_4885,N_4941);
and U5160 (N_5160,N_4504,N_4769);
nand U5161 (N_5161,N_4186,N_4850);
nor U5162 (N_5162,N_4112,N_4197);
or U5163 (N_5163,N_4431,N_4389);
or U5164 (N_5164,N_4098,N_4405);
nor U5165 (N_5165,N_4247,N_4279);
nand U5166 (N_5166,N_4005,N_4745);
or U5167 (N_5167,N_4014,N_4586);
nand U5168 (N_5168,N_4606,N_4123);
nand U5169 (N_5169,N_4572,N_4277);
or U5170 (N_5170,N_4376,N_4356);
and U5171 (N_5171,N_4483,N_4715);
or U5172 (N_5172,N_4974,N_4539);
nor U5173 (N_5173,N_4627,N_4631);
nand U5174 (N_5174,N_4217,N_4265);
and U5175 (N_5175,N_4426,N_4821);
and U5176 (N_5176,N_4205,N_4458);
nand U5177 (N_5177,N_4644,N_4304);
nor U5178 (N_5178,N_4450,N_4294);
or U5179 (N_5179,N_4340,N_4490);
xnor U5180 (N_5180,N_4379,N_4876);
nand U5181 (N_5181,N_4494,N_4683);
nand U5182 (N_5182,N_4191,N_4671);
nand U5183 (N_5183,N_4501,N_4929);
and U5184 (N_5184,N_4555,N_4327);
xnor U5185 (N_5185,N_4317,N_4339);
and U5186 (N_5186,N_4478,N_4556);
and U5187 (N_5187,N_4468,N_4908);
or U5188 (N_5188,N_4825,N_4677);
or U5189 (N_5189,N_4004,N_4353);
nand U5190 (N_5190,N_4981,N_4679);
nor U5191 (N_5191,N_4314,N_4359);
or U5192 (N_5192,N_4503,N_4045);
nor U5193 (N_5193,N_4926,N_4489);
and U5194 (N_5194,N_4540,N_4447);
nand U5195 (N_5195,N_4260,N_4388);
and U5196 (N_5196,N_4924,N_4779);
nor U5197 (N_5197,N_4467,N_4670);
and U5198 (N_5198,N_4115,N_4576);
nand U5199 (N_5199,N_4837,N_4446);
nor U5200 (N_5200,N_4324,N_4724);
or U5201 (N_5201,N_4913,N_4158);
nor U5202 (N_5202,N_4578,N_4109);
nand U5203 (N_5203,N_4498,N_4150);
and U5204 (N_5204,N_4079,N_4833);
xor U5205 (N_5205,N_4902,N_4133);
or U5206 (N_5206,N_4977,N_4757);
and U5207 (N_5207,N_4894,N_4812);
or U5208 (N_5208,N_4456,N_4252);
xnor U5209 (N_5209,N_4758,N_4439);
and U5210 (N_5210,N_4592,N_4135);
nor U5211 (N_5211,N_4700,N_4910);
xnor U5212 (N_5212,N_4121,N_4259);
xnor U5213 (N_5213,N_4382,N_4785);
nor U5214 (N_5214,N_4778,N_4726);
nor U5215 (N_5215,N_4299,N_4559);
xnor U5216 (N_5216,N_4251,N_4831);
or U5217 (N_5217,N_4116,N_4199);
xnor U5218 (N_5218,N_4652,N_4055);
and U5219 (N_5219,N_4465,N_4270);
or U5220 (N_5220,N_4028,N_4834);
or U5221 (N_5221,N_4142,N_4521);
nand U5222 (N_5222,N_4132,N_4848);
or U5223 (N_5223,N_4337,N_4420);
nand U5224 (N_5224,N_4533,N_4266);
nor U5225 (N_5225,N_4532,N_4972);
and U5226 (N_5226,N_4238,N_4325);
xnor U5227 (N_5227,N_4753,N_4018);
or U5228 (N_5228,N_4136,N_4982);
nand U5229 (N_5229,N_4836,N_4289);
nor U5230 (N_5230,N_4741,N_4900);
and U5231 (N_5231,N_4249,N_4738);
nor U5232 (N_5232,N_4598,N_4889);
xor U5233 (N_5233,N_4169,N_4511);
nor U5234 (N_5234,N_4740,N_4201);
or U5235 (N_5235,N_4603,N_4192);
xnor U5236 (N_5236,N_4607,N_4499);
nor U5237 (N_5237,N_4955,N_4349);
nor U5238 (N_5238,N_4962,N_4202);
and U5239 (N_5239,N_4377,N_4082);
or U5240 (N_5240,N_4050,N_4673);
or U5241 (N_5241,N_4413,N_4658);
nor U5242 (N_5242,N_4690,N_4313);
nand U5243 (N_5243,N_4547,N_4025);
nor U5244 (N_5244,N_4722,N_4269);
xnor U5245 (N_5245,N_4751,N_4806);
nand U5246 (N_5246,N_4281,N_4077);
nand U5247 (N_5247,N_4685,N_4562);
nand U5248 (N_5248,N_4965,N_4076);
nand U5249 (N_5249,N_4099,N_4573);
and U5250 (N_5250,N_4378,N_4937);
nand U5251 (N_5251,N_4215,N_4393);
xnor U5252 (N_5252,N_4060,N_4954);
xnor U5253 (N_5253,N_4880,N_4263);
or U5254 (N_5254,N_4273,N_4233);
or U5255 (N_5255,N_4240,N_4147);
and U5256 (N_5256,N_4968,N_4759);
xor U5257 (N_5257,N_4546,N_4179);
xor U5258 (N_5258,N_4835,N_4155);
nor U5259 (N_5259,N_4997,N_4554);
nand U5260 (N_5260,N_4448,N_4181);
and U5261 (N_5261,N_4416,N_4809);
nand U5262 (N_5262,N_4647,N_4221);
or U5263 (N_5263,N_4887,N_4792);
and U5264 (N_5264,N_4161,N_4817);
and U5265 (N_5265,N_4610,N_4513);
and U5266 (N_5266,N_4157,N_4348);
nand U5267 (N_5267,N_4657,N_4964);
xnor U5268 (N_5268,N_4328,N_4931);
and U5269 (N_5269,N_4307,N_4244);
or U5270 (N_5270,N_4605,N_4246);
xor U5271 (N_5271,N_4065,N_4224);
xnor U5272 (N_5272,N_4038,N_4302);
or U5273 (N_5273,N_4851,N_4655);
nand U5274 (N_5274,N_4961,N_4843);
and U5275 (N_5275,N_4096,N_4436);
or U5276 (N_5276,N_4706,N_4710);
nand U5277 (N_5277,N_4815,N_4790);
nand U5278 (N_5278,N_4856,N_4568);
xnor U5279 (N_5279,N_4787,N_4408);
or U5280 (N_5280,N_4714,N_4190);
or U5281 (N_5281,N_4536,N_4052);
or U5282 (N_5282,N_4824,N_4654);
nand U5283 (N_5283,N_4295,N_4558);
or U5284 (N_5284,N_4814,N_4949);
nand U5285 (N_5285,N_4613,N_4676);
nand U5286 (N_5286,N_4566,N_4250);
xnor U5287 (N_5287,N_4697,N_4844);
nor U5288 (N_5288,N_4986,N_4312);
or U5289 (N_5289,N_4308,N_4226);
and U5290 (N_5290,N_4786,N_4776);
and U5291 (N_5291,N_4784,N_4027);
xor U5292 (N_5292,N_4854,N_4646);
or U5293 (N_5293,N_4872,N_4693);
and U5294 (N_5294,N_4188,N_4515);
nand U5295 (N_5295,N_4051,N_4442);
or U5296 (N_5296,N_4530,N_4341);
nor U5297 (N_5297,N_4838,N_4796);
nand U5298 (N_5298,N_4332,N_4361);
or U5299 (N_5299,N_4963,N_4648);
nor U5300 (N_5300,N_4801,N_4433);
or U5301 (N_5301,N_4748,N_4462);
or U5302 (N_5302,N_4723,N_4286);
or U5303 (N_5303,N_4007,N_4485);
and U5304 (N_5304,N_4875,N_4721);
and U5305 (N_5305,N_4387,N_4008);
nor U5306 (N_5306,N_4072,N_4024);
nor U5307 (N_5307,N_4666,N_4656);
xnor U5308 (N_5308,N_4243,N_4905);
nor U5309 (N_5309,N_4143,N_4523);
nor U5310 (N_5310,N_4306,N_4428);
and U5311 (N_5311,N_4097,N_4103);
and U5312 (N_5312,N_4775,N_4899);
or U5313 (N_5313,N_4488,N_4765);
nor U5314 (N_5314,N_4248,N_4990);
and U5315 (N_5315,N_4791,N_4100);
or U5316 (N_5316,N_4725,N_4178);
nand U5317 (N_5317,N_4933,N_4579);
nand U5318 (N_5318,N_4023,N_4980);
or U5319 (N_5319,N_4476,N_4534);
nand U5320 (N_5320,N_4154,N_4920);
nor U5321 (N_5321,N_4667,N_4276);
nand U5322 (N_5322,N_4430,N_4545);
and U5323 (N_5323,N_4754,N_4542);
nand U5324 (N_5324,N_4782,N_4165);
and U5325 (N_5325,N_4105,N_4280);
xor U5326 (N_5326,N_4732,N_4911);
nand U5327 (N_5327,N_4543,N_4593);
and U5328 (N_5328,N_4713,N_4288);
xnor U5329 (N_5329,N_4020,N_4380);
nand U5330 (N_5330,N_4171,N_4583);
nor U5331 (N_5331,N_4896,N_4496);
nand U5332 (N_5332,N_4600,N_4879);
nand U5333 (N_5333,N_4914,N_4196);
nor U5334 (N_5334,N_4056,N_4509);
nor U5335 (N_5335,N_4282,N_4898);
nor U5336 (N_5336,N_4919,N_4923);
xor U5337 (N_5337,N_4874,N_4429);
nand U5338 (N_5338,N_4407,N_4594);
or U5339 (N_5339,N_4847,N_4764);
and U5340 (N_5340,N_4522,N_4272);
or U5341 (N_5341,N_4370,N_4826);
nand U5342 (N_5342,N_4318,N_4567);
and U5343 (N_5343,N_4943,N_4128);
and U5344 (N_5344,N_4040,N_4372);
nand U5345 (N_5345,N_4127,N_4718);
or U5346 (N_5346,N_4090,N_4596);
nor U5347 (N_5347,N_4222,N_4237);
nand U5348 (N_5348,N_4066,N_4080);
and U5349 (N_5349,N_4346,N_4641);
and U5350 (N_5350,N_4895,N_4678);
xnor U5351 (N_5351,N_4087,N_4253);
nand U5352 (N_5352,N_4691,N_4412);
and U5353 (N_5353,N_4003,N_4635);
and U5354 (N_5354,N_4254,N_4119);
and U5355 (N_5355,N_4493,N_4626);
nand U5356 (N_5356,N_4293,N_4398);
or U5357 (N_5357,N_4651,N_4364);
nor U5358 (N_5358,N_4170,N_4168);
and U5359 (N_5359,N_4695,N_4366);
and U5360 (N_5360,N_4125,N_4418);
nand U5361 (N_5361,N_4630,N_4042);
or U5362 (N_5362,N_4287,N_4772);
nand U5363 (N_5363,N_4642,N_4957);
nand U5364 (N_5364,N_4595,N_4209);
and U5365 (N_5365,N_4264,N_4915);
xor U5366 (N_5366,N_4614,N_4599);
xnor U5367 (N_5367,N_4514,N_4672);
and U5368 (N_5368,N_4746,N_4544);
or U5369 (N_5369,N_4660,N_4852);
or U5370 (N_5370,N_4172,N_4525);
nand U5371 (N_5371,N_4031,N_4022);
nand U5372 (N_5372,N_4901,N_4917);
nor U5373 (N_5373,N_4526,N_4086);
or U5374 (N_5374,N_4204,N_4035);
nor U5375 (N_5375,N_4912,N_4519);
nor U5376 (N_5376,N_4959,N_4698);
nor U5377 (N_5377,N_4414,N_4995);
nand U5378 (N_5378,N_4477,N_4423);
xor U5379 (N_5379,N_4183,N_4584);
nor U5380 (N_5380,N_4987,N_4242);
and U5381 (N_5381,N_4033,N_4996);
xor U5382 (N_5382,N_4731,N_4234);
and U5383 (N_5383,N_4026,N_4326);
nand U5384 (N_5384,N_4620,N_4484);
nor U5385 (N_5385,N_4457,N_4180);
nand U5386 (N_5386,N_4013,N_4399);
or U5387 (N_5387,N_4396,N_4351);
nor U5388 (N_5388,N_4029,N_4650);
or U5389 (N_5389,N_4827,N_4441);
nand U5390 (N_5390,N_4229,N_4141);
nor U5391 (N_5391,N_4034,N_4739);
nor U5392 (N_5392,N_4976,N_4107);
nand U5393 (N_5393,N_4882,N_4507);
and U5394 (N_5394,N_4629,N_4621);
nand U5395 (N_5395,N_4305,N_4129);
nor U5396 (N_5396,N_4069,N_4271);
and U5397 (N_5397,N_4823,N_4329);
nand U5398 (N_5398,N_4419,N_4114);
and U5399 (N_5399,N_4011,N_4760);
or U5400 (N_5400,N_4255,N_4068);
or U5401 (N_5401,N_4728,N_4878);
nand U5402 (N_5402,N_4120,N_4777);
nor U5403 (N_5403,N_4829,N_4669);
xor U5404 (N_5404,N_4053,N_4131);
or U5405 (N_5405,N_4487,N_4575);
and U5406 (N_5406,N_4232,N_4888);
nor U5407 (N_5407,N_4262,N_4624);
xnor U5408 (N_5408,N_4945,N_4553);
nand U5409 (N_5409,N_4111,N_4795);
or U5410 (N_5410,N_4720,N_4988);
nand U5411 (N_5411,N_4174,N_4301);
and U5412 (N_5412,N_4058,N_4865);
nor U5413 (N_5413,N_4793,N_4788);
nor U5414 (N_5414,N_4071,N_4632);
or U5415 (N_5415,N_4663,N_4717);
xor U5416 (N_5416,N_4482,N_4866);
xor U5417 (N_5417,N_4230,N_4892);
xnor U5418 (N_5418,N_4696,N_4245);
nand U5419 (N_5419,N_4054,N_4471);
or U5420 (N_5420,N_4884,N_4073);
and U5421 (N_5421,N_4975,N_4137);
and U5422 (N_5422,N_4400,N_4153);
and U5423 (N_5423,N_4569,N_4797);
nand U5424 (N_5424,N_4200,N_4104);
nor U5425 (N_5425,N_4330,N_4664);
nand U5426 (N_5426,N_4688,N_4092);
and U5427 (N_5427,N_4406,N_4177);
nand U5428 (N_5428,N_4214,N_4770);
xnor U5429 (N_5429,N_4228,N_4506);
xnor U5430 (N_5430,N_4189,N_4497);
nand U5431 (N_5431,N_4581,N_4993);
and U5432 (N_5432,N_4940,N_4159);
or U5433 (N_5433,N_4774,N_4858);
xnor U5434 (N_5434,N_4853,N_4374);
nor U5435 (N_5435,N_4383,N_4828);
nor U5436 (N_5436,N_4021,N_4684);
or U5437 (N_5437,N_4763,N_4502);
or U5438 (N_5438,N_4391,N_4138);
nor U5439 (N_5439,N_4106,N_4661);
xor U5440 (N_5440,N_4373,N_4047);
nand U5441 (N_5441,N_4953,N_4804);
nor U5442 (N_5442,N_4015,N_4886);
or U5443 (N_5443,N_4845,N_4952);
or U5444 (N_5444,N_4016,N_4877);
or U5445 (N_5445,N_4946,N_4508);
and U5446 (N_5446,N_4355,N_4001);
and U5447 (N_5447,N_4747,N_4334);
and U5448 (N_5448,N_4422,N_4883);
or U5449 (N_5449,N_4394,N_4212);
xnor U5450 (N_5450,N_4636,N_4999);
xnor U5451 (N_5451,N_4146,N_4682);
and U5452 (N_5452,N_4032,N_4800);
xnor U5453 (N_5453,N_4752,N_4466);
nor U5454 (N_5454,N_4333,N_4213);
nor U5455 (N_5455,N_4358,N_4459);
or U5456 (N_5456,N_4744,N_4167);
nor U5457 (N_5457,N_4319,N_4588);
nand U5458 (N_5458,N_4944,N_4017);
and U5459 (N_5459,N_4257,N_4819);
and U5460 (N_5460,N_4903,N_4402);
xnor U5461 (N_5461,N_4445,N_4891);
nor U5462 (N_5462,N_4505,N_4689);
nand U5463 (N_5463,N_4743,N_4331);
nand U5464 (N_5464,N_4619,N_4633);
or U5465 (N_5465,N_4711,N_4516);
or U5466 (N_5466,N_4906,N_4639);
or U5467 (N_5467,N_4618,N_4794);
xor U5468 (N_5468,N_4160,N_4783);
nor U5469 (N_5469,N_4163,N_4316);
xnor U5470 (N_5470,N_4085,N_4427);
or U5471 (N_5471,N_4479,N_4816);
and U5472 (N_5472,N_4736,N_4410);
nand U5473 (N_5473,N_4320,N_4735);
xnor U5474 (N_5474,N_4037,N_4692);
xnor U5475 (N_5475,N_4130,N_4601);
xor U5476 (N_5476,N_4470,N_4061);
xor U5477 (N_5477,N_4623,N_4464);
or U5478 (N_5478,N_4551,N_4323);
nor U5479 (N_5479,N_4832,N_4857);
nor U5480 (N_5480,N_4385,N_4803);
nor U5481 (N_5481,N_4811,N_4292);
nand U5482 (N_5482,N_4231,N_4218);
and U5483 (N_5483,N_4041,N_4145);
and U5484 (N_5484,N_4480,N_4930);
and U5485 (N_5485,N_4000,N_4122);
or U5486 (N_5486,N_4890,N_4849);
nor U5487 (N_5487,N_4473,N_4602);
nor U5488 (N_5488,N_4622,N_4863);
or U5489 (N_5489,N_4922,N_4799);
or U5490 (N_5490,N_4285,N_4767);
and U5491 (N_5491,N_4386,N_4335);
nor U5492 (N_5492,N_4322,N_4704);
nor U5493 (N_5493,N_4113,N_4616);
nand U5494 (N_5494,N_4893,N_4352);
nor U5495 (N_5495,N_4074,N_4638);
nor U5496 (N_5496,N_4461,N_4939);
xnor U5497 (N_5497,N_4492,N_4617);
or U5498 (N_5498,N_4012,N_4907);
and U5499 (N_5499,N_4357,N_4088);
and U5500 (N_5500,N_4162,N_4937);
xor U5501 (N_5501,N_4234,N_4303);
nor U5502 (N_5502,N_4334,N_4426);
and U5503 (N_5503,N_4435,N_4953);
nand U5504 (N_5504,N_4980,N_4187);
nand U5505 (N_5505,N_4775,N_4528);
or U5506 (N_5506,N_4009,N_4632);
or U5507 (N_5507,N_4814,N_4480);
and U5508 (N_5508,N_4466,N_4644);
nor U5509 (N_5509,N_4427,N_4651);
or U5510 (N_5510,N_4177,N_4034);
or U5511 (N_5511,N_4059,N_4376);
and U5512 (N_5512,N_4995,N_4698);
or U5513 (N_5513,N_4123,N_4432);
xnor U5514 (N_5514,N_4693,N_4225);
or U5515 (N_5515,N_4938,N_4847);
and U5516 (N_5516,N_4213,N_4643);
and U5517 (N_5517,N_4918,N_4599);
and U5518 (N_5518,N_4607,N_4661);
xor U5519 (N_5519,N_4609,N_4982);
or U5520 (N_5520,N_4669,N_4756);
and U5521 (N_5521,N_4406,N_4063);
and U5522 (N_5522,N_4650,N_4066);
xor U5523 (N_5523,N_4359,N_4532);
and U5524 (N_5524,N_4282,N_4351);
and U5525 (N_5525,N_4558,N_4427);
nand U5526 (N_5526,N_4001,N_4814);
or U5527 (N_5527,N_4045,N_4556);
xnor U5528 (N_5528,N_4050,N_4420);
nor U5529 (N_5529,N_4840,N_4763);
nand U5530 (N_5530,N_4277,N_4455);
or U5531 (N_5531,N_4048,N_4316);
and U5532 (N_5532,N_4075,N_4420);
or U5533 (N_5533,N_4741,N_4544);
and U5534 (N_5534,N_4850,N_4332);
xnor U5535 (N_5535,N_4549,N_4696);
or U5536 (N_5536,N_4614,N_4584);
xnor U5537 (N_5537,N_4847,N_4744);
nand U5538 (N_5538,N_4581,N_4822);
nand U5539 (N_5539,N_4767,N_4886);
or U5540 (N_5540,N_4701,N_4447);
nand U5541 (N_5541,N_4998,N_4619);
or U5542 (N_5542,N_4364,N_4866);
or U5543 (N_5543,N_4719,N_4619);
nor U5544 (N_5544,N_4490,N_4723);
nor U5545 (N_5545,N_4379,N_4683);
or U5546 (N_5546,N_4868,N_4042);
or U5547 (N_5547,N_4335,N_4870);
or U5548 (N_5548,N_4300,N_4201);
nor U5549 (N_5549,N_4919,N_4785);
nand U5550 (N_5550,N_4716,N_4433);
or U5551 (N_5551,N_4815,N_4720);
nor U5552 (N_5552,N_4888,N_4407);
xor U5553 (N_5553,N_4807,N_4566);
nand U5554 (N_5554,N_4948,N_4187);
nor U5555 (N_5555,N_4149,N_4560);
xnor U5556 (N_5556,N_4254,N_4460);
or U5557 (N_5557,N_4157,N_4134);
nand U5558 (N_5558,N_4518,N_4908);
nand U5559 (N_5559,N_4369,N_4934);
or U5560 (N_5560,N_4781,N_4951);
xnor U5561 (N_5561,N_4915,N_4695);
xnor U5562 (N_5562,N_4218,N_4704);
nand U5563 (N_5563,N_4130,N_4955);
nor U5564 (N_5564,N_4463,N_4958);
or U5565 (N_5565,N_4800,N_4313);
nand U5566 (N_5566,N_4457,N_4426);
xnor U5567 (N_5567,N_4847,N_4978);
or U5568 (N_5568,N_4230,N_4932);
or U5569 (N_5569,N_4377,N_4072);
and U5570 (N_5570,N_4771,N_4255);
nand U5571 (N_5571,N_4376,N_4222);
xnor U5572 (N_5572,N_4456,N_4781);
xnor U5573 (N_5573,N_4924,N_4974);
or U5574 (N_5574,N_4445,N_4709);
xnor U5575 (N_5575,N_4471,N_4122);
nand U5576 (N_5576,N_4416,N_4231);
and U5577 (N_5577,N_4222,N_4036);
xnor U5578 (N_5578,N_4339,N_4529);
nor U5579 (N_5579,N_4582,N_4147);
or U5580 (N_5580,N_4670,N_4380);
nand U5581 (N_5581,N_4909,N_4037);
nor U5582 (N_5582,N_4734,N_4062);
xnor U5583 (N_5583,N_4431,N_4201);
nand U5584 (N_5584,N_4372,N_4268);
and U5585 (N_5585,N_4783,N_4833);
and U5586 (N_5586,N_4953,N_4201);
xor U5587 (N_5587,N_4934,N_4983);
nand U5588 (N_5588,N_4743,N_4567);
xnor U5589 (N_5589,N_4181,N_4093);
nor U5590 (N_5590,N_4380,N_4658);
and U5591 (N_5591,N_4814,N_4065);
or U5592 (N_5592,N_4505,N_4971);
or U5593 (N_5593,N_4132,N_4801);
nor U5594 (N_5594,N_4724,N_4615);
nand U5595 (N_5595,N_4464,N_4201);
nand U5596 (N_5596,N_4645,N_4566);
xnor U5597 (N_5597,N_4357,N_4605);
and U5598 (N_5598,N_4157,N_4651);
nor U5599 (N_5599,N_4812,N_4944);
nand U5600 (N_5600,N_4934,N_4217);
or U5601 (N_5601,N_4696,N_4438);
and U5602 (N_5602,N_4799,N_4228);
xor U5603 (N_5603,N_4118,N_4270);
or U5604 (N_5604,N_4362,N_4602);
or U5605 (N_5605,N_4434,N_4950);
nor U5606 (N_5606,N_4849,N_4397);
xor U5607 (N_5607,N_4089,N_4531);
and U5608 (N_5608,N_4023,N_4321);
nand U5609 (N_5609,N_4971,N_4564);
nor U5610 (N_5610,N_4847,N_4420);
nand U5611 (N_5611,N_4626,N_4909);
nand U5612 (N_5612,N_4750,N_4275);
or U5613 (N_5613,N_4607,N_4131);
or U5614 (N_5614,N_4127,N_4051);
or U5615 (N_5615,N_4868,N_4608);
and U5616 (N_5616,N_4816,N_4099);
and U5617 (N_5617,N_4347,N_4986);
or U5618 (N_5618,N_4550,N_4555);
nand U5619 (N_5619,N_4165,N_4741);
xor U5620 (N_5620,N_4699,N_4965);
nor U5621 (N_5621,N_4158,N_4046);
and U5622 (N_5622,N_4091,N_4045);
and U5623 (N_5623,N_4581,N_4324);
nand U5624 (N_5624,N_4264,N_4664);
or U5625 (N_5625,N_4454,N_4286);
nor U5626 (N_5626,N_4906,N_4591);
and U5627 (N_5627,N_4910,N_4968);
or U5628 (N_5628,N_4070,N_4257);
nor U5629 (N_5629,N_4601,N_4578);
nand U5630 (N_5630,N_4354,N_4590);
nor U5631 (N_5631,N_4407,N_4691);
nor U5632 (N_5632,N_4098,N_4599);
nand U5633 (N_5633,N_4991,N_4308);
xnor U5634 (N_5634,N_4072,N_4144);
or U5635 (N_5635,N_4570,N_4059);
xor U5636 (N_5636,N_4887,N_4503);
nor U5637 (N_5637,N_4312,N_4705);
nor U5638 (N_5638,N_4038,N_4383);
xor U5639 (N_5639,N_4209,N_4109);
xnor U5640 (N_5640,N_4996,N_4963);
xnor U5641 (N_5641,N_4591,N_4969);
nor U5642 (N_5642,N_4198,N_4469);
nor U5643 (N_5643,N_4794,N_4946);
nor U5644 (N_5644,N_4678,N_4785);
nor U5645 (N_5645,N_4334,N_4413);
xnor U5646 (N_5646,N_4344,N_4392);
xnor U5647 (N_5647,N_4037,N_4571);
nand U5648 (N_5648,N_4788,N_4247);
xnor U5649 (N_5649,N_4219,N_4951);
or U5650 (N_5650,N_4063,N_4972);
or U5651 (N_5651,N_4756,N_4232);
or U5652 (N_5652,N_4096,N_4178);
nor U5653 (N_5653,N_4731,N_4870);
or U5654 (N_5654,N_4746,N_4390);
or U5655 (N_5655,N_4714,N_4078);
and U5656 (N_5656,N_4588,N_4939);
nor U5657 (N_5657,N_4110,N_4603);
nor U5658 (N_5658,N_4812,N_4174);
nand U5659 (N_5659,N_4058,N_4235);
xnor U5660 (N_5660,N_4090,N_4831);
nand U5661 (N_5661,N_4702,N_4439);
and U5662 (N_5662,N_4460,N_4244);
nand U5663 (N_5663,N_4542,N_4850);
or U5664 (N_5664,N_4998,N_4121);
xnor U5665 (N_5665,N_4957,N_4490);
and U5666 (N_5666,N_4008,N_4195);
and U5667 (N_5667,N_4242,N_4008);
or U5668 (N_5668,N_4047,N_4425);
and U5669 (N_5669,N_4515,N_4397);
or U5670 (N_5670,N_4602,N_4973);
nand U5671 (N_5671,N_4865,N_4699);
and U5672 (N_5672,N_4526,N_4572);
and U5673 (N_5673,N_4957,N_4130);
nor U5674 (N_5674,N_4427,N_4164);
and U5675 (N_5675,N_4191,N_4334);
and U5676 (N_5676,N_4147,N_4038);
xor U5677 (N_5677,N_4563,N_4772);
or U5678 (N_5678,N_4402,N_4831);
or U5679 (N_5679,N_4000,N_4567);
or U5680 (N_5680,N_4725,N_4586);
xor U5681 (N_5681,N_4962,N_4236);
xor U5682 (N_5682,N_4566,N_4720);
and U5683 (N_5683,N_4003,N_4294);
nor U5684 (N_5684,N_4073,N_4986);
and U5685 (N_5685,N_4593,N_4005);
xor U5686 (N_5686,N_4676,N_4773);
and U5687 (N_5687,N_4415,N_4235);
xor U5688 (N_5688,N_4471,N_4870);
xor U5689 (N_5689,N_4359,N_4537);
and U5690 (N_5690,N_4062,N_4690);
nand U5691 (N_5691,N_4568,N_4377);
xor U5692 (N_5692,N_4967,N_4048);
xnor U5693 (N_5693,N_4673,N_4406);
nor U5694 (N_5694,N_4508,N_4205);
nor U5695 (N_5695,N_4160,N_4712);
nand U5696 (N_5696,N_4657,N_4707);
and U5697 (N_5697,N_4253,N_4663);
and U5698 (N_5698,N_4173,N_4466);
nand U5699 (N_5699,N_4871,N_4389);
or U5700 (N_5700,N_4315,N_4945);
nand U5701 (N_5701,N_4907,N_4110);
nor U5702 (N_5702,N_4214,N_4246);
and U5703 (N_5703,N_4414,N_4745);
nor U5704 (N_5704,N_4825,N_4230);
xor U5705 (N_5705,N_4405,N_4948);
xor U5706 (N_5706,N_4434,N_4645);
nand U5707 (N_5707,N_4099,N_4668);
nand U5708 (N_5708,N_4413,N_4973);
or U5709 (N_5709,N_4521,N_4962);
and U5710 (N_5710,N_4163,N_4476);
xnor U5711 (N_5711,N_4495,N_4633);
xor U5712 (N_5712,N_4268,N_4393);
nor U5713 (N_5713,N_4523,N_4845);
nor U5714 (N_5714,N_4972,N_4924);
nand U5715 (N_5715,N_4660,N_4843);
or U5716 (N_5716,N_4764,N_4384);
and U5717 (N_5717,N_4180,N_4486);
or U5718 (N_5718,N_4548,N_4291);
xnor U5719 (N_5719,N_4107,N_4901);
nand U5720 (N_5720,N_4078,N_4867);
or U5721 (N_5721,N_4082,N_4952);
nor U5722 (N_5722,N_4853,N_4052);
xor U5723 (N_5723,N_4248,N_4015);
xor U5724 (N_5724,N_4750,N_4643);
and U5725 (N_5725,N_4277,N_4460);
and U5726 (N_5726,N_4312,N_4495);
nand U5727 (N_5727,N_4024,N_4684);
xor U5728 (N_5728,N_4019,N_4637);
xnor U5729 (N_5729,N_4473,N_4133);
or U5730 (N_5730,N_4853,N_4123);
or U5731 (N_5731,N_4431,N_4507);
or U5732 (N_5732,N_4356,N_4695);
or U5733 (N_5733,N_4216,N_4899);
and U5734 (N_5734,N_4740,N_4492);
nand U5735 (N_5735,N_4598,N_4198);
or U5736 (N_5736,N_4420,N_4614);
xor U5737 (N_5737,N_4087,N_4617);
or U5738 (N_5738,N_4087,N_4746);
or U5739 (N_5739,N_4227,N_4945);
or U5740 (N_5740,N_4119,N_4027);
and U5741 (N_5741,N_4569,N_4923);
and U5742 (N_5742,N_4831,N_4258);
and U5743 (N_5743,N_4886,N_4470);
nand U5744 (N_5744,N_4801,N_4327);
xor U5745 (N_5745,N_4719,N_4560);
and U5746 (N_5746,N_4588,N_4417);
or U5747 (N_5747,N_4542,N_4305);
and U5748 (N_5748,N_4388,N_4070);
nand U5749 (N_5749,N_4160,N_4952);
nand U5750 (N_5750,N_4353,N_4590);
xor U5751 (N_5751,N_4368,N_4608);
and U5752 (N_5752,N_4649,N_4569);
nor U5753 (N_5753,N_4597,N_4244);
xor U5754 (N_5754,N_4484,N_4793);
nand U5755 (N_5755,N_4276,N_4637);
nor U5756 (N_5756,N_4400,N_4965);
nor U5757 (N_5757,N_4801,N_4266);
and U5758 (N_5758,N_4321,N_4908);
nor U5759 (N_5759,N_4068,N_4856);
nor U5760 (N_5760,N_4081,N_4754);
xor U5761 (N_5761,N_4196,N_4699);
xnor U5762 (N_5762,N_4687,N_4992);
nand U5763 (N_5763,N_4637,N_4647);
xor U5764 (N_5764,N_4051,N_4765);
and U5765 (N_5765,N_4589,N_4030);
nand U5766 (N_5766,N_4189,N_4380);
xnor U5767 (N_5767,N_4621,N_4133);
or U5768 (N_5768,N_4906,N_4076);
xor U5769 (N_5769,N_4802,N_4115);
and U5770 (N_5770,N_4893,N_4596);
xor U5771 (N_5771,N_4499,N_4509);
or U5772 (N_5772,N_4982,N_4002);
or U5773 (N_5773,N_4376,N_4613);
nor U5774 (N_5774,N_4354,N_4848);
nand U5775 (N_5775,N_4095,N_4837);
xor U5776 (N_5776,N_4241,N_4594);
or U5777 (N_5777,N_4601,N_4288);
nand U5778 (N_5778,N_4934,N_4331);
and U5779 (N_5779,N_4006,N_4737);
nor U5780 (N_5780,N_4570,N_4259);
xnor U5781 (N_5781,N_4277,N_4293);
and U5782 (N_5782,N_4735,N_4750);
nand U5783 (N_5783,N_4761,N_4452);
nor U5784 (N_5784,N_4015,N_4410);
nor U5785 (N_5785,N_4047,N_4493);
or U5786 (N_5786,N_4542,N_4571);
and U5787 (N_5787,N_4368,N_4586);
nand U5788 (N_5788,N_4418,N_4927);
nor U5789 (N_5789,N_4352,N_4330);
or U5790 (N_5790,N_4067,N_4391);
nand U5791 (N_5791,N_4352,N_4839);
nand U5792 (N_5792,N_4586,N_4534);
and U5793 (N_5793,N_4841,N_4682);
xor U5794 (N_5794,N_4499,N_4836);
xor U5795 (N_5795,N_4357,N_4521);
and U5796 (N_5796,N_4087,N_4505);
or U5797 (N_5797,N_4237,N_4514);
nand U5798 (N_5798,N_4313,N_4873);
or U5799 (N_5799,N_4904,N_4650);
or U5800 (N_5800,N_4147,N_4185);
or U5801 (N_5801,N_4419,N_4534);
nand U5802 (N_5802,N_4947,N_4314);
nor U5803 (N_5803,N_4669,N_4596);
xor U5804 (N_5804,N_4978,N_4843);
and U5805 (N_5805,N_4271,N_4109);
xnor U5806 (N_5806,N_4790,N_4737);
or U5807 (N_5807,N_4095,N_4542);
and U5808 (N_5808,N_4664,N_4719);
or U5809 (N_5809,N_4677,N_4366);
or U5810 (N_5810,N_4487,N_4545);
xnor U5811 (N_5811,N_4297,N_4768);
or U5812 (N_5812,N_4713,N_4643);
nor U5813 (N_5813,N_4641,N_4538);
nor U5814 (N_5814,N_4923,N_4826);
xor U5815 (N_5815,N_4852,N_4482);
or U5816 (N_5816,N_4626,N_4311);
and U5817 (N_5817,N_4880,N_4301);
and U5818 (N_5818,N_4716,N_4101);
nand U5819 (N_5819,N_4193,N_4070);
nor U5820 (N_5820,N_4558,N_4172);
and U5821 (N_5821,N_4379,N_4707);
nor U5822 (N_5822,N_4230,N_4669);
nor U5823 (N_5823,N_4794,N_4152);
nor U5824 (N_5824,N_4907,N_4482);
or U5825 (N_5825,N_4001,N_4879);
nor U5826 (N_5826,N_4607,N_4682);
xor U5827 (N_5827,N_4406,N_4110);
xnor U5828 (N_5828,N_4229,N_4348);
nor U5829 (N_5829,N_4463,N_4590);
or U5830 (N_5830,N_4666,N_4522);
nor U5831 (N_5831,N_4405,N_4650);
nor U5832 (N_5832,N_4251,N_4988);
xor U5833 (N_5833,N_4351,N_4639);
xor U5834 (N_5834,N_4363,N_4226);
or U5835 (N_5835,N_4595,N_4193);
xnor U5836 (N_5836,N_4815,N_4569);
or U5837 (N_5837,N_4723,N_4951);
xnor U5838 (N_5838,N_4341,N_4955);
nand U5839 (N_5839,N_4512,N_4488);
xor U5840 (N_5840,N_4175,N_4050);
nor U5841 (N_5841,N_4147,N_4269);
and U5842 (N_5842,N_4862,N_4399);
or U5843 (N_5843,N_4111,N_4464);
and U5844 (N_5844,N_4261,N_4490);
xor U5845 (N_5845,N_4254,N_4927);
nand U5846 (N_5846,N_4699,N_4095);
or U5847 (N_5847,N_4486,N_4782);
nor U5848 (N_5848,N_4470,N_4435);
or U5849 (N_5849,N_4231,N_4467);
xnor U5850 (N_5850,N_4399,N_4214);
or U5851 (N_5851,N_4312,N_4172);
or U5852 (N_5852,N_4866,N_4844);
xor U5853 (N_5853,N_4853,N_4254);
nor U5854 (N_5854,N_4173,N_4135);
xor U5855 (N_5855,N_4848,N_4623);
or U5856 (N_5856,N_4963,N_4217);
nand U5857 (N_5857,N_4512,N_4775);
or U5858 (N_5858,N_4824,N_4735);
nand U5859 (N_5859,N_4224,N_4711);
or U5860 (N_5860,N_4264,N_4772);
or U5861 (N_5861,N_4323,N_4711);
nor U5862 (N_5862,N_4418,N_4582);
nand U5863 (N_5863,N_4036,N_4978);
nand U5864 (N_5864,N_4644,N_4053);
nor U5865 (N_5865,N_4904,N_4531);
and U5866 (N_5866,N_4592,N_4527);
nand U5867 (N_5867,N_4600,N_4264);
nor U5868 (N_5868,N_4746,N_4572);
and U5869 (N_5869,N_4841,N_4577);
xnor U5870 (N_5870,N_4117,N_4574);
nand U5871 (N_5871,N_4441,N_4886);
and U5872 (N_5872,N_4717,N_4833);
nor U5873 (N_5873,N_4771,N_4368);
xor U5874 (N_5874,N_4028,N_4574);
nand U5875 (N_5875,N_4311,N_4072);
and U5876 (N_5876,N_4956,N_4939);
xor U5877 (N_5877,N_4428,N_4081);
xor U5878 (N_5878,N_4658,N_4957);
xnor U5879 (N_5879,N_4324,N_4846);
nor U5880 (N_5880,N_4007,N_4637);
or U5881 (N_5881,N_4058,N_4982);
xnor U5882 (N_5882,N_4067,N_4028);
nor U5883 (N_5883,N_4712,N_4068);
and U5884 (N_5884,N_4331,N_4432);
and U5885 (N_5885,N_4130,N_4506);
nand U5886 (N_5886,N_4783,N_4703);
xnor U5887 (N_5887,N_4676,N_4918);
or U5888 (N_5888,N_4953,N_4695);
nor U5889 (N_5889,N_4334,N_4784);
and U5890 (N_5890,N_4402,N_4902);
xor U5891 (N_5891,N_4510,N_4561);
and U5892 (N_5892,N_4351,N_4959);
xor U5893 (N_5893,N_4537,N_4150);
and U5894 (N_5894,N_4448,N_4176);
nor U5895 (N_5895,N_4373,N_4671);
or U5896 (N_5896,N_4875,N_4330);
nor U5897 (N_5897,N_4698,N_4364);
or U5898 (N_5898,N_4762,N_4745);
nand U5899 (N_5899,N_4078,N_4139);
and U5900 (N_5900,N_4350,N_4253);
xnor U5901 (N_5901,N_4079,N_4089);
or U5902 (N_5902,N_4616,N_4922);
nor U5903 (N_5903,N_4313,N_4266);
nor U5904 (N_5904,N_4273,N_4852);
nand U5905 (N_5905,N_4380,N_4650);
nand U5906 (N_5906,N_4859,N_4944);
xnor U5907 (N_5907,N_4115,N_4756);
nand U5908 (N_5908,N_4941,N_4247);
xor U5909 (N_5909,N_4414,N_4656);
nand U5910 (N_5910,N_4616,N_4505);
nand U5911 (N_5911,N_4535,N_4021);
and U5912 (N_5912,N_4975,N_4810);
or U5913 (N_5913,N_4893,N_4505);
or U5914 (N_5914,N_4703,N_4918);
nor U5915 (N_5915,N_4932,N_4755);
and U5916 (N_5916,N_4741,N_4282);
xnor U5917 (N_5917,N_4268,N_4214);
xnor U5918 (N_5918,N_4229,N_4056);
or U5919 (N_5919,N_4980,N_4234);
nor U5920 (N_5920,N_4971,N_4886);
nand U5921 (N_5921,N_4349,N_4519);
xnor U5922 (N_5922,N_4656,N_4822);
and U5923 (N_5923,N_4667,N_4949);
or U5924 (N_5924,N_4335,N_4795);
xnor U5925 (N_5925,N_4042,N_4542);
nand U5926 (N_5926,N_4829,N_4908);
xnor U5927 (N_5927,N_4830,N_4466);
nand U5928 (N_5928,N_4246,N_4860);
and U5929 (N_5929,N_4710,N_4132);
or U5930 (N_5930,N_4756,N_4992);
xor U5931 (N_5931,N_4569,N_4244);
or U5932 (N_5932,N_4991,N_4947);
xor U5933 (N_5933,N_4037,N_4811);
xor U5934 (N_5934,N_4070,N_4278);
xnor U5935 (N_5935,N_4432,N_4251);
and U5936 (N_5936,N_4857,N_4264);
nand U5937 (N_5937,N_4660,N_4091);
xnor U5938 (N_5938,N_4386,N_4815);
nor U5939 (N_5939,N_4525,N_4536);
xor U5940 (N_5940,N_4640,N_4344);
xnor U5941 (N_5941,N_4954,N_4301);
or U5942 (N_5942,N_4477,N_4117);
xnor U5943 (N_5943,N_4190,N_4893);
or U5944 (N_5944,N_4908,N_4599);
or U5945 (N_5945,N_4216,N_4553);
nand U5946 (N_5946,N_4117,N_4610);
nor U5947 (N_5947,N_4219,N_4699);
nand U5948 (N_5948,N_4914,N_4078);
nand U5949 (N_5949,N_4737,N_4446);
or U5950 (N_5950,N_4005,N_4969);
and U5951 (N_5951,N_4368,N_4348);
and U5952 (N_5952,N_4956,N_4850);
nand U5953 (N_5953,N_4424,N_4372);
xnor U5954 (N_5954,N_4569,N_4950);
and U5955 (N_5955,N_4744,N_4444);
and U5956 (N_5956,N_4271,N_4650);
and U5957 (N_5957,N_4965,N_4939);
and U5958 (N_5958,N_4675,N_4571);
or U5959 (N_5959,N_4609,N_4844);
nor U5960 (N_5960,N_4711,N_4094);
xnor U5961 (N_5961,N_4339,N_4570);
and U5962 (N_5962,N_4337,N_4207);
nor U5963 (N_5963,N_4991,N_4887);
nand U5964 (N_5964,N_4306,N_4728);
nand U5965 (N_5965,N_4217,N_4173);
or U5966 (N_5966,N_4635,N_4840);
xor U5967 (N_5967,N_4508,N_4175);
nor U5968 (N_5968,N_4292,N_4086);
xor U5969 (N_5969,N_4036,N_4251);
nand U5970 (N_5970,N_4001,N_4893);
nor U5971 (N_5971,N_4416,N_4545);
nor U5972 (N_5972,N_4067,N_4920);
xor U5973 (N_5973,N_4736,N_4151);
xnor U5974 (N_5974,N_4660,N_4886);
nand U5975 (N_5975,N_4897,N_4275);
nor U5976 (N_5976,N_4074,N_4499);
nand U5977 (N_5977,N_4064,N_4147);
xor U5978 (N_5978,N_4053,N_4148);
xnor U5979 (N_5979,N_4694,N_4631);
xnor U5980 (N_5980,N_4056,N_4887);
nand U5981 (N_5981,N_4361,N_4267);
nor U5982 (N_5982,N_4943,N_4958);
and U5983 (N_5983,N_4544,N_4136);
nand U5984 (N_5984,N_4018,N_4883);
or U5985 (N_5985,N_4937,N_4399);
and U5986 (N_5986,N_4280,N_4812);
nand U5987 (N_5987,N_4015,N_4309);
xor U5988 (N_5988,N_4068,N_4617);
xor U5989 (N_5989,N_4500,N_4662);
or U5990 (N_5990,N_4245,N_4316);
xor U5991 (N_5991,N_4532,N_4710);
xnor U5992 (N_5992,N_4057,N_4525);
or U5993 (N_5993,N_4701,N_4773);
xor U5994 (N_5994,N_4394,N_4837);
nand U5995 (N_5995,N_4929,N_4708);
xor U5996 (N_5996,N_4412,N_4749);
nand U5997 (N_5997,N_4753,N_4403);
nand U5998 (N_5998,N_4916,N_4951);
or U5999 (N_5999,N_4560,N_4943);
and U6000 (N_6000,N_5054,N_5769);
xor U6001 (N_6001,N_5080,N_5431);
xor U6002 (N_6002,N_5762,N_5987);
and U6003 (N_6003,N_5001,N_5745);
and U6004 (N_6004,N_5962,N_5951);
or U6005 (N_6005,N_5771,N_5249);
nand U6006 (N_6006,N_5470,N_5624);
and U6007 (N_6007,N_5802,N_5486);
and U6008 (N_6008,N_5430,N_5239);
nand U6009 (N_6009,N_5741,N_5573);
xnor U6010 (N_6010,N_5899,N_5945);
or U6011 (N_6011,N_5213,N_5687);
nand U6012 (N_6012,N_5625,N_5627);
nor U6013 (N_6013,N_5197,N_5153);
nor U6014 (N_6014,N_5735,N_5123);
or U6015 (N_6015,N_5812,N_5324);
or U6016 (N_6016,N_5526,N_5079);
nand U6017 (N_6017,N_5510,N_5650);
and U6018 (N_6018,N_5699,N_5871);
and U6019 (N_6019,N_5633,N_5838);
xor U6020 (N_6020,N_5551,N_5960);
xnor U6021 (N_6021,N_5746,N_5384);
nor U6022 (N_6022,N_5293,N_5643);
and U6023 (N_6023,N_5007,N_5182);
and U6024 (N_6024,N_5955,N_5698);
nand U6025 (N_6025,N_5282,N_5559);
and U6026 (N_6026,N_5235,N_5364);
xnor U6027 (N_6027,N_5337,N_5408);
xor U6028 (N_6028,N_5676,N_5439);
and U6029 (N_6029,N_5133,N_5209);
or U6030 (N_6030,N_5928,N_5141);
or U6031 (N_6031,N_5243,N_5464);
nand U6032 (N_6032,N_5543,N_5936);
xnor U6033 (N_6033,N_5634,N_5806);
nor U6034 (N_6034,N_5664,N_5198);
xor U6035 (N_6035,N_5981,N_5948);
or U6036 (N_6036,N_5527,N_5314);
or U6037 (N_6037,N_5598,N_5031);
or U6038 (N_6038,N_5111,N_5246);
nand U6039 (N_6039,N_5301,N_5799);
nand U6040 (N_6040,N_5704,N_5791);
xor U6041 (N_6041,N_5017,N_5846);
xnor U6042 (N_6042,N_5742,N_5810);
and U6043 (N_6043,N_5331,N_5740);
or U6044 (N_6044,N_5567,N_5264);
or U6045 (N_6045,N_5095,N_5181);
and U6046 (N_6046,N_5018,N_5623);
nand U6047 (N_6047,N_5262,N_5353);
nor U6048 (N_6048,N_5541,N_5531);
nand U6049 (N_6049,N_5013,N_5338);
nor U6050 (N_6050,N_5026,N_5481);
xnor U6051 (N_6051,N_5577,N_5930);
and U6052 (N_6052,N_5117,N_5878);
nand U6053 (N_6053,N_5773,N_5009);
and U6054 (N_6054,N_5654,N_5042);
nand U6055 (N_6055,N_5880,N_5903);
and U6056 (N_6056,N_5874,N_5662);
xor U6057 (N_6057,N_5789,N_5589);
and U6058 (N_6058,N_5655,N_5750);
or U6059 (N_6059,N_5120,N_5852);
nor U6060 (N_6060,N_5516,N_5547);
or U6061 (N_6061,N_5944,N_5062);
nand U6062 (N_6062,N_5507,N_5569);
nand U6063 (N_6063,N_5142,N_5836);
xnor U6064 (N_6064,N_5394,N_5918);
or U6065 (N_6065,N_5058,N_5494);
nor U6066 (N_6066,N_5192,N_5232);
or U6067 (N_6067,N_5482,N_5942);
nor U6068 (N_6068,N_5994,N_5258);
or U6069 (N_6069,N_5612,N_5954);
or U6070 (N_6070,N_5252,N_5053);
or U6071 (N_6071,N_5440,N_5927);
xnor U6072 (N_6072,N_5362,N_5003);
nand U6073 (N_6073,N_5496,N_5963);
xnor U6074 (N_6074,N_5497,N_5719);
nand U6075 (N_6075,N_5418,N_5448);
xnor U6076 (N_6076,N_5420,N_5653);
nand U6077 (N_6077,N_5727,N_5863);
and U6078 (N_6078,N_5902,N_5862);
nand U6079 (N_6079,N_5522,N_5114);
nand U6080 (N_6080,N_5808,N_5816);
and U6081 (N_6081,N_5827,N_5593);
and U6082 (N_6082,N_5307,N_5467);
xnor U6083 (N_6083,N_5900,N_5309);
nor U6084 (N_6084,N_5753,N_5148);
nor U6085 (N_6085,N_5275,N_5012);
nor U6086 (N_6086,N_5377,N_5230);
and U6087 (N_6087,N_5629,N_5201);
and U6088 (N_6088,N_5221,N_5493);
or U6089 (N_6089,N_5390,N_5979);
or U6090 (N_6090,N_5595,N_5649);
nor U6091 (N_6091,N_5545,N_5885);
nor U6092 (N_6092,N_5733,N_5992);
and U6093 (N_6093,N_5028,N_5160);
nand U6094 (N_6094,N_5333,N_5202);
xor U6095 (N_6095,N_5501,N_5912);
and U6096 (N_6096,N_5705,N_5996);
or U6097 (N_6097,N_5894,N_5679);
or U6098 (N_6098,N_5147,N_5098);
and U6099 (N_6099,N_5882,N_5554);
nand U6100 (N_6100,N_5609,N_5100);
and U6101 (N_6101,N_5129,N_5724);
nor U6102 (N_6102,N_5535,N_5688);
xor U6103 (N_6103,N_5973,N_5958);
nand U6104 (N_6104,N_5970,N_5689);
or U6105 (N_6105,N_5596,N_5116);
or U6106 (N_6106,N_5835,N_5387);
nand U6107 (N_6107,N_5240,N_5093);
xnor U6108 (N_6108,N_5328,N_5382);
nor U6109 (N_6109,N_5847,N_5564);
nor U6110 (N_6110,N_5277,N_5823);
nand U6111 (N_6111,N_5159,N_5723);
nor U6112 (N_6112,N_5381,N_5082);
nor U6113 (N_6113,N_5236,N_5940);
nand U6114 (N_6114,N_5638,N_5509);
and U6115 (N_6115,N_5785,N_5647);
or U6116 (N_6116,N_5168,N_5030);
and U6117 (N_6117,N_5794,N_5599);
or U6118 (N_6118,N_5298,N_5580);
nor U6119 (N_6119,N_5626,N_5586);
nand U6120 (N_6120,N_5778,N_5392);
xnor U6121 (N_6121,N_5751,N_5020);
and U6122 (N_6122,N_5767,N_5225);
nor U6123 (N_6123,N_5619,N_5419);
xor U6124 (N_6124,N_5186,N_5367);
or U6125 (N_6125,N_5804,N_5045);
or U6126 (N_6126,N_5474,N_5779);
or U6127 (N_6127,N_5274,N_5081);
and U6128 (N_6128,N_5984,N_5811);
and U6129 (N_6129,N_5986,N_5477);
nand U6130 (N_6130,N_5563,N_5344);
nand U6131 (N_6131,N_5064,N_5303);
xor U6132 (N_6132,N_5658,N_5561);
nand U6133 (N_6133,N_5359,N_5965);
and U6134 (N_6134,N_5582,N_5226);
and U6135 (N_6135,N_5845,N_5245);
and U6136 (N_6136,N_5652,N_5269);
or U6137 (N_6137,N_5416,N_5669);
nor U6138 (N_6138,N_5834,N_5251);
and U6139 (N_6139,N_5991,N_5102);
and U6140 (N_6140,N_5155,N_5721);
nor U6141 (N_6141,N_5071,N_5128);
xnor U6142 (N_6142,N_5278,N_5161);
nand U6143 (N_6143,N_5857,N_5537);
or U6144 (N_6144,N_5046,N_5312);
or U6145 (N_6145,N_5280,N_5273);
nand U6146 (N_6146,N_5590,N_5043);
nor U6147 (N_6147,N_5261,N_5819);
nor U6148 (N_6148,N_5019,N_5397);
nor U6149 (N_6149,N_5241,N_5967);
nor U6150 (N_6150,N_5843,N_5920);
xnor U6151 (N_6151,N_5411,N_5438);
and U6152 (N_6152,N_5896,N_5460);
and U6153 (N_6153,N_5879,N_5413);
and U6154 (N_6154,N_5317,N_5714);
nor U6155 (N_6155,N_5718,N_5858);
xnor U6156 (N_6156,N_5790,N_5343);
or U6157 (N_6157,N_5105,N_5432);
or U6158 (N_6158,N_5259,N_5047);
xor U6159 (N_6159,N_5763,N_5572);
xnor U6160 (N_6160,N_5177,N_5780);
xnor U6161 (N_6161,N_5131,N_5622);
nand U6162 (N_6162,N_5883,N_5395);
nor U6163 (N_6163,N_5579,N_5491);
or U6164 (N_6164,N_5736,N_5844);
or U6165 (N_6165,N_5815,N_5352);
and U6166 (N_6166,N_5410,N_5950);
xnor U6167 (N_6167,N_5929,N_5399);
xnor U6168 (N_6168,N_5839,N_5985);
xnor U6169 (N_6169,N_5861,N_5453);
nor U6170 (N_6170,N_5611,N_5690);
and U6171 (N_6171,N_5566,N_5884);
nand U6172 (N_6172,N_5999,N_5330);
nand U6173 (N_6173,N_5754,N_5886);
or U6174 (N_6174,N_5150,N_5840);
xnor U6175 (N_6175,N_5592,N_5085);
nor U6176 (N_6176,N_5946,N_5010);
nor U6177 (N_6177,N_5975,N_5977);
nor U6178 (N_6178,N_5988,N_5311);
xor U6179 (N_6179,N_5925,N_5548);
or U6180 (N_6180,N_5171,N_5923);
or U6181 (N_6181,N_5210,N_5506);
and U6182 (N_6182,N_5725,N_5694);
or U6183 (N_6183,N_5693,N_5015);
nor U6184 (N_6184,N_5040,N_5403);
xor U6185 (N_6185,N_5898,N_5435);
nand U6186 (N_6186,N_5025,N_5480);
nand U6187 (N_6187,N_5208,N_5553);
or U6188 (N_6188,N_5520,N_5604);
and U6189 (N_6189,N_5833,N_5864);
nor U6190 (N_6190,N_5585,N_5254);
and U6191 (N_6191,N_5427,N_5890);
and U6192 (N_6192,N_5848,N_5222);
xor U6193 (N_6193,N_5409,N_5937);
or U6194 (N_6194,N_5373,N_5542);
nor U6195 (N_6195,N_5152,N_5692);
nand U6196 (N_6196,N_5630,N_5670);
and U6197 (N_6197,N_5326,N_5229);
or U6198 (N_6198,N_5027,N_5038);
nor U6199 (N_6199,N_5938,N_5821);
or U6200 (N_6200,N_5055,N_5966);
nor U6201 (N_6201,N_5747,N_5931);
xor U6202 (N_6202,N_5989,N_5351);
and U6203 (N_6203,N_5442,N_5648);
nand U6204 (N_6204,N_5014,N_5969);
and U6205 (N_6205,N_5299,N_5473);
and U6206 (N_6206,N_5617,N_5600);
nand U6207 (N_6207,N_5175,N_5683);
nor U6208 (N_6208,N_5214,N_5122);
nor U6209 (N_6209,N_5190,N_5228);
nand U6210 (N_6210,N_5841,N_5119);
or U6211 (N_6211,N_5907,N_5421);
nand U6212 (N_6212,N_5008,N_5517);
nor U6213 (N_6213,N_5734,N_5466);
nand U6214 (N_6214,N_5036,N_5876);
xor U6215 (N_6215,N_5540,N_5276);
nand U6216 (N_6216,N_5914,N_5107);
xnor U6217 (N_6217,N_5402,N_5901);
nand U6218 (N_6218,N_5078,N_5720);
or U6219 (N_6219,N_5178,N_5266);
or U6220 (N_6220,N_5933,N_5132);
nor U6221 (N_6221,N_5370,N_5795);
nand U6222 (N_6222,N_5345,N_5113);
nand U6223 (N_6223,N_5376,N_5726);
nor U6224 (N_6224,N_5378,N_5911);
and U6225 (N_6225,N_5656,N_5088);
and U6226 (N_6226,N_5452,N_5866);
nor U6227 (N_6227,N_5521,N_5552);
nor U6228 (N_6228,N_5730,N_5538);
and U6229 (N_6229,N_5528,N_5405);
xnor U6230 (N_6230,N_5905,N_5749);
and U6231 (N_6231,N_5711,N_5300);
or U6232 (N_6232,N_5350,N_5170);
nor U6233 (N_6233,N_5859,N_5060);
nand U6234 (N_6234,N_5587,N_5556);
or U6235 (N_6235,N_5072,N_5756);
or U6236 (N_6236,N_5760,N_5176);
or U6237 (N_6237,N_5490,N_5037);
nor U6238 (N_6238,N_5748,N_5233);
nor U6239 (N_6239,N_5358,N_5947);
xnor U6240 (N_6240,N_5185,N_5850);
or U6241 (N_6241,N_5529,N_5660);
xnor U6242 (N_6242,N_5605,N_5897);
and U6243 (N_6243,N_5423,N_5729);
nor U6244 (N_6244,N_5112,N_5283);
nor U6245 (N_6245,N_5562,N_5681);
and U6246 (N_6246,N_5052,N_5061);
nand U6247 (N_6247,N_5713,N_5519);
xor U6248 (N_6248,N_5515,N_5875);
nand U6249 (N_6249,N_5360,N_5825);
xnor U6250 (N_6250,N_5546,N_5908);
nor U6251 (N_6251,N_5101,N_5837);
and U6252 (N_6252,N_5069,N_5444);
and U6253 (N_6253,N_5635,N_5686);
or U6254 (N_6254,N_5982,N_5263);
xnor U6255 (N_6255,N_5104,N_5818);
and U6256 (N_6256,N_5505,N_5196);
xnor U6257 (N_6257,N_5602,N_5433);
nand U6258 (N_6258,N_5024,N_5504);
nand U6259 (N_6259,N_5379,N_5935);
and U6260 (N_6260,N_5469,N_5881);
or U6261 (N_6261,N_5797,N_5709);
xor U6262 (N_6262,N_5393,N_5077);
xor U6263 (N_6263,N_5800,N_5917);
and U6264 (N_6264,N_5220,N_5476);
xnor U6265 (N_6265,N_5135,N_5108);
or U6266 (N_6266,N_5479,N_5498);
nand U6267 (N_6267,N_5667,N_5887);
nand U6268 (N_6268,N_5584,N_5436);
xor U6269 (N_6269,N_5260,N_5005);
nand U6270 (N_6270,N_5755,N_5570);
nor U6271 (N_6271,N_5523,N_5006);
xnor U6272 (N_6272,N_5244,N_5456);
xnor U6273 (N_6273,N_5347,N_5073);
and U6274 (N_6274,N_5124,N_5086);
or U6275 (N_6275,N_5434,N_5842);
nor U6276 (N_6276,N_5739,N_5447);
xnor U6277 (N_6277,N_5820,N_5065);
and U6278 (N_6278,N_5211,N_5514);
nand U6279 (N_6279,N_5206,N_5136);
and U6280 (N_6280,N_5732,N_5500);
nor U6281 (N_6281,N_5856,N_5340);
xnor U6282 (N_6282,N_5461,N_5829);
and U6283 (N_6283,N_5285,N_5772);
xnor U6284 (N_6284,N_5286,N_5365);
xnor U6285 (N_6285,N_5004,N_5118);
or U6286 (N_6286,N_5889,N_5671);
nor U6287 (N_6287,N_5374,N_5029);
nor U6288 (N_6288,N_5388,N_5361);
xnor U6289 (N_6289,N_5675,N_5391);
or U6290 (N_6290,N_5781,N_5096);
or U6291 (N_6291,N_5615,N_5348);
nor U6292 (N_6292,N_5854,N_5227);
or U6293 (N_6293,N_5319,N_5865);
nand U6294 (N_6294,N_5425,N_5140);
or U6295 (N_6295,N_5488,N_5386);
and U6296 (N_6296,N_5616,N_5145);
and U6297 (N_6297,N_5059,N_5666);
or U6298 (N_6298,N_5591,N_5173);
nand U6299 (N_6299,N_5639,N_5400);
nand U6300 (N_6300,N_5092,N_5722);
and U6301 (N_6301,N_5256,N_5759);
and U6302 (N_6302,N_5308,N_5022);
and U6303 (N_6303,N_5315,N_5163);
nor U6304 (N_6304,N_5180,N_5558);
and U6305 (N_6305,N_5349,N_5939);
and U6306 (N_6306,N_5223,N_5659);
xnor U6307 (N_6307,N_5199,N_5606);
nand U6308 (N_6308,N_5106,N_5700);
and U6309 (N_6309,N_5696,N_5701);
xor U6310 (N_6310,N_5034,N_5137);
xnor U6311 (N_6311,N_5288,N_5809);
nand U6312 (N_6312,N_5305,N_5267);
and U6313 (N_6313,N_5422,N_5463);
and U6314 (N_6314,N_5524,N_5215);
nand U6315 (N_6315,N_5651,N_5188);
nand U6316 (N_6316,N_5325,N_5518);
xnor U6317 (N_6317,N_5039,N_5508);
xor U6318 (N_6318,N_5943,N_5455);
xnor U6319 (N_6319,N_5801,N_5503);
or U6320 (N_6320,N_5873,N_5250);
xor U6321 (N_6321,N_5000,N_5321);
xor U6322 (N_6322,N_5710,N_5478);
or U6323 (N_6323,N_5398,N_5238);
or U6324 (N_6324,N_5568,N_5224);
and U6325 (N_6325,N_5661,N_5091);
or U6326 (N_6326,N_5237,N_5891);
nand U6327 (N_6327,N_5777,N_5157);
nor U6328 (N_6328,N_5761,N_5798);
xnor U6329 (N_6329,N_5021,N_5849);
or U6330 (N_6330,N_5063,N_5297);
nor U6331 (N_6331,N_5860,N_5707);
and U6332 (N_6332,N_5796,N_5075);
nor U6333 (N_6333,N_5471,N_5407);
xnor U6334 (N_6334,N_5512,N_5764);
or U6335 (N_6335,N_5956,N_5271);
and U6336 (N_6336,N_5731,N_5995);
nand U6337 (N_6337,N_5533,N_5475);
or U6338 (N_6338,N_5787,N_5443);
nor U6339 (N_6339,N_5164,N_5070);
and U6340 (N_6340,N_5121,N_5357);
xor U6341 (N_6341,N_5680,N_5824);
nor U6342 (N_6342,N_5492,N_5212);
nand U6343 (N_6343,N_5255,N_5485);
or U6344 (N_6344,N_5099,N_5404);
or U6345 (N_6345,N_5597,N_5355);
xnor U6346 (N_6346,N_5621,N_5457);
and U6347 (N_6347,N_5576,N_5445);
nand U6348 (N_6348,N_5603,N_5002);
and U6349 (N_6349,N_5717,N_5926);
nor U6350 (N_6350,N_5231,N_5893);
nor U6351 (N_6351,N_5472,N_5765);
nand U6352 (N_6352,N_5032,N_5691);
nor U6353 (N_6353,N_5187,N_5204);
xnor U6354 (N_6354,N_5483,N_5921);
and U6355 (N_6355,N_5990,N_5162);
or U6356 (N_6356,N_5316,N_5334);
nor U6357 (N_6357,N_5284,N_5684);
or U6358 (N_6358,N_5998,N_5557);
xnor U6359 (N_6359,N_5703,N_5770);
and U6360 (N_6360,N_5744,N_5607);
xor U6361 (N_6361,N_5339,N_5203);
nor U6362 (N_6362,N_5620,N_5166);
nor U6363 (N_6363,N_5952,N_5143);
or U6364 (N_6364,N_5242,N_5855);
or U6365 (N_6365,N_5103,N_5877);
and U6366 (N_6366,N_5685,N_5363);
or U6367 (N_6367,N_5429,N_5127);
or U6368 (N_6368,N_5289,N_5830);
nand U6369 (N_6369,N_5997,N_5139);
nor U6370 (N_6370,N_5158,N_5601);
and U6371 (N_6371,N_5813,N_5169);
or U6372 (N_6372,N_5194,N_5156);
or U6373 (N_6373,N_5044,N_5291);
and U6374 (N_6374,N_5953,N_5428);
xor U6375 (N_6375,N_5869,N_5803);
or U6376 (N_6376,N_5910,N_5292);
or U6377 (N_6377,N_5502,N_5268);
nand U6378 (N_6378,N_5571,N_5657);
xnor U6379 (N_6379,N_5318,N_5642);
nor U6380 (N_6380,N_5641,N_5752);
or U6381 (N_6381,N_5578,N_5788);
or U6382 (N_6382,N_5867,N_5814);
xnor U6383 (N_6383,N_5087,N_5784);
xnor U6384 (N_6384,N_5290,N_5248);
xnor U6385 (N_6385,N_5441,N_5322);
nor U6386 (N_6386,N_5412,N_5468);
or U6387 (N_6387,N_5281,N_5459);
nand U6388 (N_6388,N_5805,N_5167);
or U6389 (N_6389,N_5396,N_5076);
and U6390 (N_6390,N_5851,N_5971);
nand U6391 (N_6391,N_5909,N_5919);
nor U6392 (N_6392,N_5183,N_5513);
and U6393 (N_6393,N_5668,N_5304);
and U6394 (N_6394,N_5594,N_5888);
nand U6395 (N_6395,N_5853,N_5383);
xor U6396 (N_6396,N_5941,N_5417);
or U6397 (N_6397,N_5449,N_5446);
nand U6398 (N_6398,N_5536,N_5870);
nor U6399 (N_6399,N_5544,N_5138);
or U6400 (N_6400,N_5993,N_5712);
and U6401 (N_6401,N_5310,N_5831);
nor U6402 (N_6402,N_5146,N_5041);
or U6403 (N_6403,N_5332,N_5151);
nor U6404 (N_6404,N_5892,N_5189);
nand U6405 (N_6405,N_5775,N_5766);
xor U6406 (N_6406,N_5066,N_5023);
nand U6407 (N_6407,N_5050,N_5961);
or U6408 (N_6408,N_5195,N_5640);
and U6409 (N_6409,N_5094,N_5172);
nand U6410 (N_6410,N_5932,N_5035);
nor U6411 (N_6411,N_5549,N_5499);
xnor U6412 (N_6412,N_5757,N_5375);
nand U6413 (N_6413,N_5828,N_5588);
nand U6414 (N_6414,N_5134,N_5327);
or U6415 (N_6415,N_5895,N_5495);
or U6416 (N_6416,N_5610,N_5636);
nand U6417 (N_6417,N_5306,N_5758);
xor U6418 (N_6418,N_5265,N_5356);
nor U6419 (N_6419,N_5462,N_5109);
and U6420 (N_6420,N_5272,N_5368);
or U6421 (N_6421,N_5978,N_5774);
or U6422 (N_6422,N_5279,N_5323);
nand U6423 (N_6423,N_5426,N_5628);
nand U6424 (N_6424,N_5980,N_5826);
xnor U6425 (N_6425,N_5964,N_5389);
xor U6426 (N_6426,N_5354,N_5335);
nand U6427 (N_6427,N_5565,N_5663);
xor U6428 (N_6428,N_5083,N_5807);
nand U6429 (N_6429,N_5179,N_5125);
and U6430 (N_6430,N_5346,N_5674);
nor U6431 (N_6431,N_5832,N_5530);
nor U6432 (N_6432,N_5184,N_5716);
xnor U6433 (N_6433,N_5057,N_5677);
nor U6434 (N_6434,N_5401,N_5257);
nor U6435 (N_6435,N_5632,N_5115);
nor U6436 (N_6436,N_5922,N_5695);
xor U6437 (N_6437,N_5555,N_5369);
xor U6438 (N_6438,N_5234,N_5016);
and U6439 (N_6439,N_5218,N_5974);
and U6440 (N_6440,N_5665,N_5165);
and U6441 (N_6441,N_5454,N_5253);
nor U6442 (N_6442,N_5702,N_5406);
and U6443 (N_6443,N_5424,N_5631);
or U6444 (N_6444,N_5645,N_5738);
xnor U6445 (N_6445,N_5782,N_5560);
or U6446 (N_6446,N_5637,N_5793);
or U6447 (N_6447,N_5051,N_5792);
nand U6448 (N_6448,N_5380,N_5916);
or U6449 (N_6449,N_5783,N_5247);
nor U6450 (N_6450,N_5097,N_5525);
and U6451 (N_6451,N_5972,N_5174);
nand U6452 (N_6452,N_5534,N_5465);
xor U6453 (N_6453,N_5341,N_5678);
nor U6454 (N_6454,N_5934,N_5608);
xor U6455 (N_6455,N_5074,N_5768);
nor U6456 (N_6456,N_5084,N_5450);
or U6457 (N_6457,N_5110,N_5414);
xor U6458 (N_6458,N_5049,N_5822);
nor U6459 (N_6459,N_5144,N_5320);
nor U6460 (N_6460,N_5776,N_5329);
xnor U6461 (N_6461,N_5968,N_5313);
and U6462 (N_6462,N_5484,N_5200);
or U6463 (N_6463,N_5371,N_5959);
xnor U6464 (N_6464,N_5715,N_5294);
and U6465 (N_6465,N_5614,N_5574);
and U6466 (N_6466,N_5270,N_5682);
nand U6467 (N_6467,N_5672,N_5868);
and U6468 (N_6468,N_5913,N_5906);
nor U6469 (N_6469,N_5539,N_5817);
or U6470 (N_6470,N_5743,N_5708);
nand U6471 (N_6471,N_5487,N_5983);
nand U6472 (N_6472,N_5737,N_5550);
xor U6473 (N_6473,N_5613,N_5089);
nor U6474 (N_6474,N_5451,N_5904);
or U6475 (N_6475,N_5644,N_5366);
nand U6476 (N_6476,N_5949,N_5385);
nor U6477 (N_6477,N_5924,N_5216);
xnor U6478 (N_6478,N_5915,N_5618);
xnor U6479 (N_6479,N_5193,N_5532);
and U6480 (N_6480,N_5296,N_5033);
nand U6481 (N_6481,N_5126,N_5646);
nand U6482 (N_6482,N_5207,N_5697);
nand U6483 (N_6483,N_5011,N_5130);
xnor U6484 (N_6484,N_5786,N_5458);
xnor U6485 (N_6485,N_5154,N_5336);
or U6486 (N_6486,N_5489,N_5706);
nand U6487 (N_6487,N_5205,N_5149);
and U6488 (N_6488,N_5581,N_5976);
or U6489 (N_6489,N_5342,N_5219);
xnor U6490 (N_6490,N_5575,N_5067);
or U6491 (N_6491,N_5287,N_5191);
or U6492 (N_6492,N_5415,N_5090);
nand U6493 (N_6493,N_5217,N_5068);
nor U6494 (N_6494,N_5511,N_5372);
and U6495 (N_6495,N_5048,N_5302);
nand U6496 (N_6496,N_5728,N_5437);
and U6497 (N_6497,N_5673,N_5872);
xor U6498 (N_6498,N_5583,N_5957);
nand U6499 (N_6499,N_5056,N_5295);
nand U6500 (N_6500,N_5093,N_5009);
nor U6501 (N_6501,N_5522,N_5334);
and U6502 (N_6502,N_5319,N_5982);
and U6503 (N_6503,N_5980,N_5067);
and U6504 (N_6504,N_5120,N_5723);
xnor U6505 (N_6505,N_5844,N_5325);
or U6506 (N_6506,N_5465,N_5665);
or U6507 (N_6507,N_5117,N_5744);
nand U6508 (N_6508,N_5184,N_5729);
and U6509 (N_6509,N_5441,N_5903);
and U6510 (N_6510,N_5208,N_5385);
xnor U6511 (N_6511,N_5277,N_5991);
or U6512 (N_6512,N_5244,N_5607);
or U6513 (N_6513,N_5519,N_5482);
nand U6514 (N_6514,N_5845,N_5624);
or U6515 (N_6515,N_5212,N_5092);
or U6516 (N_6516,N_5748,N_5436);
nand U6517 (N_6517,N_5605,N_5775);
or U6518 (N_6518,N_5308,N_5033);
and U6519 (N_6519,N_5012,N_5339);
nor U6520 (N_6520,N_5987,N_5021);
nor U6521 (N_6521,N_5871,N_5392);
and U6522 (N_6522,N_5737,N_5760);
nand U6523 (N_6523,N_5161,N_5203);
nor U6524 (N_6524,N_5583,N_5672);
and U6525 (N_6525,N_5129,N_5599);
or U6526 (N_6526,N_5906,N_5739);
or U6527 (N_6527,N_5610,N_5129);
nor U6528 (N_6528,N_5494,N_5022);
xnor U6529 (N_6529,N_5378,N_5365);
nor U6530 (N_6530,N_5943,N_5823);
xor U6531 (N_6531,N_5064,N_5439);
nor U6532 (N_6532,N_5274,N_5764);
or U6533 (N_6533,N_5531,N_5459);
or U6534 (N_6534,N_5603,N_5898);
nor U6535 (N_6535,N_5734,N_5913);
nand U6536 (N_6536,N_5158,N_5284);
or U6537 (N_6537,N_5526,N_5677);
and U6538 (N_6538,N_5943,N_5522);
xnor U6539 (N_6539,N_5490,N_5345);
nand U6540 (N_6540,N_5562,N_5927);
and U6541 (N_6541,N_5344,N_5763);
and U6542 (N_6542,N_5000,N_5763);
and U6543 (N_6543,N_5018,N_5523);
or U6544 (N_6544,N_5999,N_5257);
nand U6545 (N_6545,N_5276,N_5521);
nor U6546 (N_6546,N_5478,N_5746);
or U6547 (N_6547,N_5192,N_5146);
nor U6548 (N_6548,N_5959,N_5993);
or U6549 (N_6549,N_5626,N_5891);
or U6550 (N_6550,N_5131,N_5659);
and U6551 (N_6551,N_5046,N_5342);
nand U6552 (N_6552,N_5453,N_5549);
nand U6553 (N_6553,N_5646,N_5168);
nand U6554 (N_6554,N_5780,N_5662);
nor U6555 (N_6555,N_5760,N_5850);
or U6556 (N_6556,N_5270,N_5967);
or U6557 (N_6557,N_5719,N_5347);
nor U6558 (N_6558,N_5101,N_5789);
nand U6559 (N_6559,N_5999,N_5570);
nor U6560 (N_6560,N_5737,N_5954);
nand U6561 (N_6561,N_5143,N_5892);
nor U6562 (N_6562,N_5023,N_5075);
and U6563 (N_6563,N_5320,N_5701);
nand U6564 (N_6564,N_5973,N_5650);
xnor U6565 (N_6565,N_5218,N_5639);
nor U6566 (N_6566,N_5751,N_5911);
and U6567 (N_6567,N_5423,N_5371);
or U6568 (N_6568,N_5001,N_5112);
and U6569 (N_6569,N_5036,N_5402);
xnor U6570 (N_6570,N_5445,N_5231);
and U6571 (N_6571,N_5625,N_5471);
nor U6572 (N_6572,N_5851,N_5132);
nor U6573 (N_6573,N_5255,N_5101);
nor U6574 (N_6574,N_5242,N_5262);
and U6575 (N_6575,N_5907,N_5416);
or U6576 (N_6576,N_5903,N_5139);
or U6577 (N_6577,N_5429,N_5200);
xnor U6578 (N_6578,N_5362,N_5026);
nor U6579 (N_6579,N_5561,N_5575);
xnor U6580 (N_6580,N_5360,N_5773);
xor U6581 (N_6581,N_5887,N_5231);
nor U6582 (N_6582,N_5204,N_5112);
and U6583 (N_6583,N_5811,N_5238);
nand U6584 (N_6584,N_5843,N_5627);
nor U6585 (N_6585,N_5672,N_5621);
or U6586 (N_6586,N_5958,N_5299);
or U6587 (N_6587,N_5237,N_5598);
nand U6588 (N_6588,N_5192,N_5939);
xor U6589 (N_6589,N_5784,N_5099);
nor U6590 (N_6590,N_5446,N_5900);
xnor U6591 (N_6591,N_5560,N_5388);
nand U6592 (N_6592,N_5181,N_5417);
nor U6593 (N_6593,N_5129,N_5606);
xnor U6594 (N_6594,N_5658,N_5562);
and U6595 (N_6595,N_5627,N_5880);
xnor U6596 (N_6596,N_5702,N_5173);
nor U6597 (N_6597,N_5531,N_5814);
xnor U6598 (N_6598,N_5578,N_5168);
nor U6599 (N_6599,N_5572,N_5070);
nor U6600 (N_6600,N_5810,N_5897);
and U6601 (N_6601,N_5375,N_5869);
and U6602 (N_6602,N_5063,N_5142);
and U6603 (N_6603,N_5874,N_5235);
xor U6604 (N_6604,N_5216,N_5775);
or U6605 (N_6605,N_5460,N_5695);
or U6606 (N_6606,N_5372,N_5883);
xor U6607 (N_6607,N_5693,N_5346);
nor U6608 (N_6608,N_5950,N_5116);
nor U6609 (N_6609,N_5585,N_5442);
nor U6610 (N_6610,N_5636,N_5019);
xnor U6611 (N_6611,N_5791,N_5671);
or U6612 (N_6612,N_5331,N_5840);
nand U6613 (N_6613,N_5660,N_5349);
nand U6614 (N_6614,N_5231,N_5235);
or U6615 (N_6615,N_5026,N_5830);
and U6616 (N_6616,N_5980,N_5107);
nand U6617 (N_6617,N_5708,N_5940);
nor U6618 (N_6618,N_5363,N_5023);
nand U6619 (N_6619,N_5905,N_5158);
xnor U6620 (N_6620,N_5999,N_5993);
or U6621 (N_6621,N_5519,N_5251);
or U6622 (N_6622,N_5505,N_5873);
and U6623 (N_6623,N_5456,N_5276);
and U6624 (N_6624,N_5447,N_5436);
xnor U6625 (N_6625,N_5859,N_5307);
or U6626 (N_6626,N_5988,N_5659);
and U6627 (N_6627,N_5671,N_5284);
and U6628 (N_6628,N_5958,N_5275);
xnor U6629 (N_6629,N_5305,N_5095);
xor U6630 (N_6630,N_5284,N_5792);
and U6631 (N_6631,N_5209,N_5434);
and U6632 (N_6632,N_5321,N_5033);
nor U6633 (N_6633,N_5294,N_5527);
nor U6634 (N_6634,N_5871,N_5781);
and U6635 (N_6635,N_5552,N_5704);
xnor U6636 (N_6636,N_5800,N_5245);
and U6637 (N_6637,N_5501,N_5359);
nand U6638 (N_6638,N_5542,N_5341);
xor U6639 (N_6639,N_5850,N_5394);
nor U6640 (N_6640,N_5333,N_5398);
nand U6641 (N_6641,N_5237,N_5517);
xor U6642 (N_6642,N_5101,N_5449);
and U6643 (N_6643,N_5719,N_5039);
nor U6644 (N_6644,N_5204,N_5224);
nor U6645 (N_6645,N_5878,N_5722);
xor U6646 (N_6646,N_5253,N_5636);
nand U6647 (N_6647,N_5042,N_5311);
nand U6648 (N_6648,N_5079,N_5715);
nand U6649 (N_6649,N_5669,N_5509);
xor U6650 (N_6650,N_5290,N_5860);
nand U6651 (N_6651,N_5810,N_5738);
or U6652 (N_6652,N_5615,N_5572);
or U6653 (N_6653,N_5238,N_5643);
xor U6654 (N_6654,N_5930,N_5728);
and U6655 (N_6655,N_5594,N_5703);
xnor U6656 (N_6656,N_5726,N_5536);
or U6657 (N_6657,N_5219,N_5874);
nand U6658 (N_6658,N_5300,N_5613);
nor U6659 (N_6659,N_5398,N_5933);
nand U6660 (N_6660,N_5465,N_5681);
and U6661 (N_6661,N_5287,N_5799);
nor U6662 (N_6662,N_5362,N_5736);
nand U6663 (N_6663,N_5806,N_5276);
nor U6664 (N_6664,N_5890,N_5139);
nor U6665 (N_6665,N_5027,N_5405);
and U6666 (N_6666,N_5509,N_5714);
nor U6667 (N_6667,N_5183,N_5509);
and U6668 (N_6668,N_5858,N_5040);
or U6669 (N_6669,N_5936,N_5091);
or U6670 (N_6670,N_5171,N_5084);
or U6671 (N_6671,N_5511,N_5287);
xor U6672 (N_6672,N_5076,N_5407);
xor U6673 (N_6673,N_5065,N_5701);
and U6674 (N_6674,N_5644,N_5088);
nor U6675 (N_6675,N_5441,N_5912);
xor U6676 (N_6676,N_5948,N_5345);
xor U6677 (N_6677,N_5083,N_5619);
nand U6678 (N_6678,N_5492,N_5486);
xor U6679 (N_6679,N_5248,N_5830);
nand U6680 (N_6680,N_5769,N_5983);
nand U6681 (N_6681,N_5900,N_5919);
nand U6682 (N_6682,N_5692,N_5791);
xor U6683 (N_6683,N_5979,N_5348);
nor U6684 (N_6684,N_5698,N_5875);
xnor U6685 (N_6685,N_5253,N_5862);
xnor U6686 (N_6686,N_5439,N_5246);
nand U6687 (N_6687,N_5179,N_5478);
nand U6688 (N_6688,N_5731,N_5012);
nor U6689 (N_6689,N_5522,N_5271);
or U6690 (N_6690,N_5655,N_5566);
xnor U6691 (N_6691,N_5507,N_5900);
nor U6692 (N_6692,N_5619,N_5247);
and U6693 (N_6693,N_5679,N_5198);
xnor U6694 (N_6694,N_5867,N_5130);
and U6695 (N_6695,N_5501,N_5217);
nor U6696 (N_6696,N_5106,N_5670);
and U6697 (N_6697,N_5693,N_5734);
xor U6698 (N_6698,N_5512,N_5869);
and U6699 (N_6699,N_5115,N_5786);
and U6700 (N_6700,N_5756,N_5796);
and U6701 (N_6701,N_5939,N_5722);
xor U6702 (N_6702,N_5919,N_5128);
and U6703 (N_6703,N_5757,N_5033);
nand U6704 (N_6704,N_5153,N_5402);
or U6705 (N_6705,N_5500,N_5224);
xor U6706 (N_6706,N_5103,N_5595);
and U6707 (N_6707,N_5339,N_5041);
nand U6708 (N_6708,N_5018,N_5063);
nand U6709 (N_6709,N_5712,N_5314);
and U6710 (N_6710,N_5290,N_5958);
and U6711 (N_6711,N_5165,N_5612);
or U6712 (N_6712,N_5697,N_5429);
nand U6713 (N_6713,N_5703,N_5520);
or U6714 (N_6714,N_5954,N_5185);
xor U6715 (N_6715,N_5513,N_5816);
and U6716 (N_6716,N_5019,N_5950);
and U6717 (N_6717,N_5954,N_5462);
and U6718 (N_6718,N_5675,N_5253);
or U6719 (N_6719,N_5519,N_5010);
or U6720 (N_6720,N_5072,N_5669);
nor U6721 (N_6721,N_5113,N_5480);
nand U6722 (N_6722,N_5965,N_5493);
nand U6723 (N_6723,N_5164,N_5567);
and U6724 (N_6724,N_5506,N_5391);
or U6725 (N_6725,N_5418,N_5850);
nand U6726 (N_6726,N_5809,N_5085);
nor U6727 (N_6727,N_5288,N_5140);
and U6728 (N_6728,N_5717,N_5164);
nand U6729 (N_6729,N_5652,N_5277);
or U6730 (N_6730,N_5156,N_5351);
xor U6731 (N_6731,N_5417,N_5759);
xor U6732 (N_6732,N_5704,N_5974);
nand U6733 (N_6733,N_5512,N_5484);
nor U6734 (N_6734,N_5201,N_5866);
and U6735 (N_6735,N_5280,N_5523);
nor U6736 (N_6736,N_5603,N_5894);
or U6737 (N_6737,N_5009,N_5081);
nor U6738 (N_6738,N_5196,N_5127);
and U6739 (N_6739,N_5689,N_5773);
or U6740 (N_6740,N_5580,N_5592);
xor U6741 (N_6741,N_5364,N_5994);
xnor U6742 (N_6742,N_5788,N_5718);
and U6743 (N_6743,N_5399,N_5888);
xnor U6744 (N_6744,N_5778,N_5827);
nor U6745 (N_6745,N_5451,N_5375);
nand U6746 (N_6746,N_5411,N_5884);
nand U6747 (N_6747,N_5087,N_5556);
and U6748 (N_6748,N_5929,N_5310);
nand U6749 (N_6749,N_5196,N_5359);
nor U6750 (N_6750,N_5068,N_5514);
nand U6751 (N_6751,N_5262,N_5295);
and U6752 (N_6752,N_5194,N_5070);
nand U6753 (N_6753,N_5169,N_5323);
xnor U6754 (N_6754,N_5928,N_5946);
xor U6755 (N_6755,N_5421,N_5625);
xor U6756 (N_6756,N_5285,N_5489);
and U6757 (N_6757,N_5677,N_5414);
nand U6758 (N_6758,N_5144,N_5858);
nor U6759 (N_6759,N_5282,N_5782);
nor U6760 (N_6760,N_5006,N_5984);
nand U6761 (N_6761,N_5383,N_5872);
nand U6762 (N_6762,N_5532,N_5068);
nor U6763 (N_6763,N_5796,N_5689);
xor U6764 (N_6764,N_5471,N_5447);
nand U6765 (N_6765,N_5949,N_5628);
xnor U6766 (N_6766,N_5638,N_5763);
or U6767 (N_6767,N_5177,N_5223);
xnor U6768 (N_6768,N_5339,N_5180);
nor U6769 (N_6769,N_5978,N_5301);
nand U6770 (N_6770,N_5175,N_5852);
xnor U6771 (N_6771,N_5221,N_5627);
xnor U6772 (N_6772,N_5220,N_5761);
nand U6773 (N_6773,N_5503,N_5796);
xor U6774 (N_6774,N_5816,N_5335);
nor U6775 (N_6775,N_5318,N_5286);
and U6776 (N_6776,N_5253,N_5176);
nand U6777 (N_6777,N_5445,N_5456);
nor U6778 (N_6778,N_5350,N_5367);
nand U6779 (N_6779,N_5679,N_5962);
xnor U6780 (N_6780,N_5327,N_5045);
nor U6781 (N_6781,N_5035,N_5461);
and U6782 (N_6782,N_5462,N_5584);
and U6783 (N_6783,N_5961,N_5253);
or U6784 (N_6784,N_5573,N_5224);
xnor U6785 (N_6785,N_5401,N_5089);
and U6786 (N_6786,N_5742,N_5887);
nand U6787 (N_6787,N_5001,N_5752);
xor U6788 (N_6788,N_5403,N_5882);
nor U6789 (N_6789,N_5948,N_5935);
and U6790 (N_6790,N_5498,N_5998);
xor U6791 (N_6791,N_5902,N_5882);
nand U6792 (N_6792,N_5965,N_5766);
or U6793 (N_6793,N_5384,N_5000);
nor U6794 (N_6794,N_5733,N_5388);
and U6795 (N_6795,N_5906,N_5501);
nand U6796 (N_6796,N_5919,N_5035);
or U6797 (N_6797,N_5206,N_5513);
and U6798 (N_6798,N_5297,N_5773);
or U6799 (N_6799,N_5955,N_5904);
nand U6800 (N_6800,N_5675,N_5081);
or U6801 (N_6801,N_5917,N_5073);
nand U6802 (N_6802,N_5764,N_5054);
or U6803 (N_6803,N_5892,N_5961);
nor U6804 (N_6804,N_5367,N_5858);
nand U6805 (N_6805,N_5264,N_5500);
nor U6806 (N_6806,N_5739,N_5337);
nand U6807 (N_6807,N_5775,N_5162);
and U6808 (N_6808,N_5561,N_5847);
or U6809 (N_6809,N_5649,N_5076);
and U6810 (N_6810,N_5425,N_5266);
and U6811 (N_6811,N_5596,N_5509);
nor U6812 (N_6812,N_5031,N_5479);
or U6813 (N_6813,N_5776,N_5655);
nand U6814 (N_6814,N_5390,N_5506);
and U6815 (N_6815,N_5842,N_5718);
or U6816 (N_6816,N_5865,N_5523);
nand U6817 (N_6817,N_5140,N_5176);
xnor U6818 (N_6818,N_5414,N_5383);
nor U6819 (N_6819,N_5915,N_5146);
xor U6820 (N_6820,N_5473,N_5719);
nor U6821 (N_6821,N_5208,N_5896);
and U6822 (N_6822,N_5206,N_5808);
or U6823 (N_6823,N_5192,N_5621);
nor U6824 (N_6824,N_5831,N_5086);
and U6825 (N_6825,N_5769,N_5071);
nand U6826 (N_6826,N_5502,N_5253);
nand U6827 (N_6827,N_5848,N_5036);
or U6828 (N_6828,N_5386,N_5876);
or U6829 (N_6829,N_5461,N_5673);
nand U6830 (N_6830,N_5142,N_5361);
nor U6831 (N_6831,N_5133,N_5432);
or U6832 (N_6832,N_5065,N_5832);
and U6833 (N_6833,N_5526,N_5976);
or U6834 (N_6834,N_5618,N_5643);
xor U6835 (N_6835,N_5679,N_5839);
nor U6836 (N_6836,N_5656,N_5704);
or U6837 (N_6837,N_5759,N_5646);
and U6838 (N_6838,N_5839,N_5432);
xor U6839 (N_6839,N_5754,N_5436);
and U6840 (N_6840,N_5435,N_5831);
nor U6841 (N_6841,N_5784,N_5532);
nand U6842 (N_6842,N_5394,N_5979);
nor U6843 (N_6843,N_5347,N_5105);
xnor U6844 (N_6844,N_5791,N_5529);
and U6845 (N_6845,N_5955,N_5164);
and U6846 (N_6846,N_5231,N_5592);
and U6847 (N_6847,N_5428,N_5391);
nor U6848 (N_6848,N_5005,N_5903);
or U6849 (N_6849,N_5871,N_5424);
nor U6850 (N_6850,N_5945,N_5627);
nor U6851 (N_6851,N_5684,N_5052);
or U6852 (N_6852,N_5250,N_5391);
or U6853 (N_6853,N_5948,N_5169);
xnor U6854 (N_6854,N_5545,N_5615);
and U6855 (N_6855,N_5157,N_5285);
xor U6856 (N_6856,N_5553,N_5574);
nand U6857 (N_6857,N_5145,N_5740);
and U6858 (N_6858,N_5104,N_5037);
nor U6859 (N_6859,N_5851,N_5058);
and U6860 (N_6860,N_5194,N_5137);
nor U6861 (N_6861,N_5910,N_5733);
xor U6862 (N_6862,N_5009,N_5211);
nor U6863 (N_6863,N_5364,N_5283);
and U6864 (N_6864,N_5149,N_5144);
nor U6865 (N_6865,N_5365,N_5778);
nor U6866 (N_6866,N_5882,N_5641);
nand U6867 (N_6867,N_5766,N_5504);
and U6868 (N_6868,N_5886,N_5930);
nand U6869 (N_6869,N_5907,N_5785);
nand U6870 (N_6870,N_5700,N_5052);
xnor U6871 (N_6871,N_5028,N_5697);
or U6872 (N_6872,N_5617,N_5511);
and U6873 (N_6873,N_5280,N_5328);
nor U6874 (N_6874,N_5539,N_5150);
and U6875 (N_6875,N_5335,N_5989);
nand U6876 (N_6876,N_5635,N_5127);
or U6877 (N_6877,N_5734,N_5529);
nand U6878 (N_6878,N_5343,N_5920);
nand U6879 (N_6879,N_5587,N_5583);
and U6880 (N_6880,N_5839,N_5214);
or U6881 (N_6881,N_5859,N_5340);
and U6882 (N_6882,N_5199,N_5138);
or U6883 (N_6883,N_5835,N_5017);
xnor U6884 (N_6884,N_5397,N_5979);
or U6885 (N_6885,N_5211,N_5580);
xnor U6886 (N_6886,N_5735,N_5523);
xor U6887 (N_6887,N_5096,N_5321);
and U6888 (N_6888,N_5757,N_5997);
nand U6889 (N_6889,N_5162,N_5154);
nand U6890 (N_6890,N_5593,N_5672);
and U6891 (N_6891,N_5057,N_5776);
xnor U6892 (N_6892,N_5026,N_5736);
or U6893 (N_6893,N_5115,N_5140);
nor U6894 (N_6894,N_5313,N_5979);
and U6895 (N_6895,N_5104,N_5654);
nor U6896 (N_6896,N_5404,N_5861);
xnor U6897 (N_6897,N_5004,N_5482);
or U6898 (N_6898,N_5511,N_5098);
nand U6899 (N_6899,N_5016,N_5535);
xor U6900 (N_6900,N_5856,N_5137);
nand U6901 (N_6901,N_5630,N_5929);
xor U6902 (N_6902,N_5348,N_5567);
nor U6903 (N_6903,N_5962,N_5837);
xnor U6904 (N_6904,N_5010,N_5501);
or U6905 (N_6905,N_5459,N_5284);
and U6906 (N_6906,N_5155,N_5643);
nand U6907 (N_6907,N_5909,N_5491);
and U6908 (N_6908,N_5486,N_5517);
and U6909 (N_6909,N_5314,N_5373);
and U6910 (N_6910,N_5153,N_5759);
or U6911 (N_6911,N_5939,N_5049);
nand U6912 (N_6912,N_5860,N_5174);
and U6913 (N_6913,N_5918,N_5973);
xor U6914 (N_6914,N_5678,N_5267);
and U6915 (N_6915,N_5943,N_5026);
nand U6916 (N_6916,N_5519,N_5202);
xnor U6917 (N_6917,N_5110,N_5717);
nand U6918 (N_6918,N_5852,N_5170);
xor U6919 (N_6919,N_5336,N_5270);
xor U6920 (N_6920,N_5902,N_5926);
nand U6921 (N_6921,N_5961,N_5043);
and U6922 (N_6922,N_5491,N_5291);
xnor U6923 (N_6923,N_5146,N_5287);
nor U6924 (N_6924,N_5028,N_5759);
and U6925 (N_6925,N_5494,N_5318);
and U6926 (N_6926,N_5227,N_5475);
nand U6927 (N_6927,N_5419,N_5380);
and U6928 (N_6928,N_5461,N_5890);
and U6929 (N_6929,N_5070,N_5648);
xnor U6930 (N_6930,N_5169,N_5121);
xnor U6931 (N_6931,N_5857,N_5509);
xnor U6932 (N_6932,N_5474,N_5233);
nand U6933 (N_6933,N_5684,N_5531);
xor U6934 (N_6934,N_5026,N_5676);
nand U6935 (N_6935,N_5101,N_5889);
nand U6936 (N_6936,N_5090,N_5770);
nand U6937 (N_6937,N_5483,N_5256);
nand U6938 (N_6938,N_5586,N_5116);
nor U6939 (N_6939,N_5390,N_5470);
and U6940 (N_6940,N_5265,N_5848);
and U6941 (N_6941,N_5362,N_5903);
xor U6942 (N_6942,N_5859,N_5800);
and U6943 (N_6943,N_5359,N_5895);
xnor U6944 (N_6944,N_5036,N_5029);
xnor U6945 (N_6945,N_5701,N_5208);
xor U6946 (N_6946,N_5336,N_5078);
nor U6947 (N_6947,N_5464,N_5939);
nor U6948 (N_6948,N_5407,N_5403);
nor U6949 (N_6949,N_5195,N_5473);
nand U6950 (N_6950,N_5471,N_5643);
nand U6951 (N_6951,N_5033,N_5556);
xor U6952 (N_6952,N_5578,N_5857);
and U6953 (N_6953,N_5670,N_5952);
or U6954 (N_6954,N_5829,N_5151);
nand U6955 (N_6955,N_5909,N_5793);
and U6956 (N_6956,N_5909,N_5925);
nor U6957 (N_6957,N_5771,N_5992);
or U6958 (N_6958,N_5826,N_5925);
and U6959 (N_6959,N_5564,N_5214);
or U6960 (N_6960,N_5849,N_5127);
and U6961 (N_6961,N_5252,N_5958);
nor U6962 (N_6962,N_5892,N_5057);
nor U6963 (N_6963,N_5704,N_5054);
or U6964 (N_6964,N_5675,N_5019);
xor U6965 (N_6965,N_5774,N_5042);
nand U6966 (N_6966,N_5658,N_5321);
and U6967 (N_6967,N_5676,N_5644);
nand U6968 (N_6968,N_5346,N_5353);
nand U6969 (N_6969,N_5552,N_5215);
nor U6970 (N_6970,N_5188,N_5829);
nor U6971 (N_6971,N_5757,N_5061);
nor U6972 (N_6972,N_5334,N_5731);
and U6973 (N_6973,N_5120,N_5572);
xor U6974 (N_6974,N_5068,N_5454);
nor U6975 (N_6975,N_5664,N_5870);
and U6976 (N_6976,N_5836,N_5940);
and U6977 (N_6977,N_5767,N_5390);
xor U6978 (N_6978,N_5773,N_5495);
and U6979 (N_6979,N_5817,N_5069);
xnor U6980 (N_6980,N_5357,N_5341);
nor U6981 (N_6981,N_5802,N_5267);
nor U6982 (N_6982,N_5818,N_5765);
xnor U6983 (N_6983,N_5420,N_5780);
xor U6984 (N_6984,N_5909,N_5388);
or U6985 (N_6985,N_5579,N_5052);
xor U6986 (N_6986,N_5134,N_5883);
xor U6987 (N_6987,N_5318,N_5677);
xor U6988 (N_6988,N_5511,N_5653);
or U6989 (N_6989,N_5339,N_5294);
or U6990 (N_6990,N_5207,N_5128);
nor U6991 (N_6991,N_5020,N_5448);
nor U6992 (N_6992,N_5422,N_5265);
nor U6993 (N_6993,N_5990,N_5277);
nand U6994 (N_6994,N_5447,N_5983);
or U6995 (N_6995,N_5205,N_5965);
nand U6996 (N_6996,N_5808,N_5863);
or U6997 (N_6997,N_5836,N_5179);
xor U6998 (N_6998,N_5738,N_5606);
nand U6999 (N_6999,N_5034,N_5773);
or U7000 (N_7000,N_6923,N_6315);
xor U7001 (N_7001,N_6463,N_6859);
nor U7002 (N_7002,N_6055,N_6603);
or U7003 (N_7003,N_6319,N_6595);
xnor U7004 (N_7004,N_6614,N_6140);
nor U7005 (N_7005,N_6577,N_6156);
or U7006 (N_7006,N_6978,N_6877);
nand U7007 (N_7007,N_6266,N_6599);
xor U7008 (N_7008,N_6081,N_6321);
xor U7009 (N_7009,N_6890,N_6540);
and U7010 (N_7010,N_6930,N_6450);
nand U7011 (N_7011,N_6063,N_6001);
nand U7012 (N_7012,N_6416,N_6099);
and U7013 (N_7013,N_6491,N_6992);
or U7014 (N_7014,N_6823,N_6171);
nand U7015 (N_7015,N_6670,N_6863);
and U7016 (N_7016,N_6498,N_6429);
nand U7017 (N_7017,N_6672,N_6418);
or U7018 (N_7018,N_6914,N_6068);
or U7019 (N_7019,N_6257,N_6015);
or U7020 (N_7020,N_6348,N_6986);
nor U7021 (N_7021,N_6184,N_6387);
nor U7022 (N_7022,N_6717,N_6868);
nand U7023 (N_7023,N_6052,N_6518);
nor U7024 (N_7024,N_6311,N_6270);
nor U7025 (N_7025,N_6486,N_6940);
nor U7026 (N_7026,N_6697,N_6324);
xnor U7027 (N_7027,N_6118,N_6427);
nor U7028 (N_7028,N_6051,N_6803);
and U7029 (N_7029,N_6981,N_6901);
and U7030 (N_7030,N_6556,N_6912);
or U7031 (N_7031,N_6925,N_6080);
or U7032 (N_7032,N_6719,N_6283);
nor U7033 (N_7033,N_6759,N_6881);
and U7034 (N_7034,N_6846,N_6316);
or U7035 (N_7035,N_6012,N_6292);
nor U7036 (N_7036,N_6249,N_6618);
and U7037 (N_7037,N_6422,N_6627);
nor U7038 (N_7038,N_6400,N_6189);
nor U7039 (N_7039,N_6641,N_6751);
nand U7040 (N_7040,N_6048,N_6535);
or U7041 (N_7041,N_6737,N_6936);
and U7042 (N_7042,N_6245,N_6836);
nor U7043 (N_7043,N_6182,N_6820);
or U7044 (N_7044,N_6109,N_6061);
nand U7045 (N_7045,N_6433,N_6659);
xnor U7046 (N_7046,N_6769,N_6529);
xor U7047 (N_7047,N_6917,N_6044);
nor U7048 (N_7048,N_6758,N_6456);
nor U7049 (N_7049,N_6875,N_6882);
nor U7050 (N_7050,N_6223,N_6632);
nor U7051 (N_7051,N_6970,N_6442);
nand U7052 (N_7052,N_6306,N_6447);
or U7053 (N_7053,N_6354,N_6723);
and U7054 (N_7054,N_6232,N_6927);
nand U7055 (N_7055,N_6384,N_6642);
nor U7056 (N_7056,N_6459,N_6715);
nand U7057 (N_7057,N_6713,N_6916);
and U7058 (N_7058,N_6607,N_6476);
xnor U7059 (N_7059,N_6772,N_6106);
nand U7060 (N_7060,N_6299,N_6691);
or U7061 (N_7061,N_6902,N_6307);
nor U7062 (N_7062,N_6405,N_6924);
xnor U7063 (N_7063,N_6764,N_6669);
or U7064 (N_7064,N_6471,N_6839);
nand U7065 (N_7065,N_6013,N_6372);
nand U7066 (N_7066,N_6496,N_6796);
or U7067 (N_7067,N_6129,N_6609);
xnor U7068 (N_7068,N_6520,N_6141);
xnor U7069 (N_7069,N_6009,N_6120);
or U7070 (N_7070,N_6660,N_6236);
or U7071 (N_7071,N_6760,N_6615);
and U7072 (N_7072,N_6147,N_6745);
xor U7073 (N_7073,N_6512,N_6532);
nand U7074 (N_7074,N_6302,N_6473);
nor U7075 (N_7075,N_6227,N_6122);
nor U7076 (N_7076,N_6775,N_6159);
nand U7077 (N_7077,N_6948,N_6583);
xor U7078 (N_7078,N_6822,N_6551);
or U7079 (N_7079,N_6967,N_6298);
and U7080 (N_7080,N_6467,N_6439);
xnor U7081 (N_7081,N_6907,N_6766);
or U7082 (N_7082,N_6199,N_6169);
or U7083 (N_7083,N_6550,N_6167);
and U7084 (N_7084,N_6074,N_6272);
nor U7085 (N_7085,N_6706,N_6938);
nor U7086 (N_7086,N_6260,N_6087);
and U7087 (N_7087,N_6395,N_6630);
nand U7088 (N_7088,N_6698,N_6945);
or U7089 (N_7089,N_6606,N_6460);
nand U7090 (N_7090,N_6489,N_6869);
xnor U7091 (N_7091,N_6284,N_6452);
nand U7092 (N_7092,N_6033,N_6380);
or U7093 (N_7093,N_6552,N_6214);
or U7094 (N_7094,N_6020,N_6179);
nor U7095 (N_7095,N_6424,N_6941);
xor U7096 (N_7096,N_6225,N_6993);
xnor U7097 (N_7097,N_6317,N_6515);
nand U7098 (N_7098,N_6041,N_6493);
or U7099 (N_7099,N_6743,N_6218);
and U7100 (N_7100,N_6586,N_6206);
nor U7101 (N_7101,N_6144,N_6036);
xnor U7102 (N_7102,N_6497,N_6326);
nor U7103 (N_7103,N_6776,N_6542);
or U7104 (N_7104,N_6029,N_6633);
or U7105 (N_7105,N_6246,N_6406);
and U7106 (N_7106,N_6662,N_6997);
xnor U7107 (N_7107,N_6782,N_6534);
and U7108 (N_7108,N_6414,N_6440);
xnor U7109 (N_7109,N_6749,N_6193);
and U7110 (N_7110,N_6024,N_6340);
nor U7111 (N_7111,N_6777,N_6248);
and U7112 (N_7112,N_6409,N_6856);
xnor U7113 (N_7113,N_6721,N_6522);
xnor U7114 (N_7114,N_6408,N_6794);
or U7115 (N_7115,N_6007,N_6346);
xor U7116 (N_7116,N_6038,N_6666);
or U7117 (N_7117,N_6059,N_6176);
and U7118 (N_7118,N_6990,N_6752);
nor U7119 (N_7119,N_6658,N_6593);
or U7120 (N_7120,N_6037,N_6181);
and U7121 (N_7121,N_6438,N_6343);
nand U7122 (N_7122,N_6410,N_6965);
nor U7123 (N_7123,N_6386,N_6533);
nand U7124 (N_7124,N_6928,N_6098);
nand U7125 (N_7125,N_6728,N_6964);
nor U7126 (N_7126,N_6237,N_6815);
nor U7127 (N_7127,N_6664,N_6499);
or U7128 (N_7128,N_6116,N_6350);
xnor U7129 (N_7129,N_6904,N_6108);
and U7130 (N_7130,N_6332,N_6274);
and U7131 (N_7131,N_6300,N_6119);
nand U7132 (N_7132,N_6867,N_6774);
or U7133 (N_7133,N_6799,N_6834);
xor U7134 (N_7134,N_6661,N_6800);
nor U7135 (N_7135,N_6314,N_6401);
nand U7136 (N_7136,N_6251,N_6514);
nor U7137 (N_7137,N_6710,N_6268);
nand U7138 (N_7138,N_6151,N_6654);
xnor U7139 (N_7139,N_6053,N_6216);
xor U7140 (N_7140,N_6154,N_6297);
or U7141 (N_7141,N_6714,N_6622);
nor U7142 (N_7142,N_6561,N_6973);
xor U7143 (N_7143,N_6788,N_6860);
xnor U7144 (N_7144,N_6072,N_6444);
and U7145 (N_7145,N_6265,N_6420);
xnor U7146 (N_7146,N_6356,N_6634);
xor U7147 (N_7147,N_6239,N_6908);
xor U7148 (N_7148,N_6761,N_6589);
or U7149 (N_7149,N_6682,N_6631);
xor U7150 (N_7150,N_6798,N_6918);
nand U7151 (N_7151,N_6293,N_6353);
nand U7152 (N_7152,N_6187,N_6352);
xor U7153 (N_7153,N_6909,N_6730);
or U7154 (N_7154,N_6177,N_6736);
and U7155 (N_7155,N_6318,N_6261);
xnor U7156 (N_7156,N_6046,N_6235);
xor U7157 (N_7157,N_6503,N_6831);
or U7158 (N_7158,N_6695,N_6271);
and U7159 (N_7159,N_6853,N_6139);
or U7160 (N_7160,N_6005,N_6011);
nor U7161 (N_7161,N_6826,N_6162);
nor U7162 (N_7162,N_6365,N_6191);
nor U7163 (N_7163,N_6485,N_6519);
xnor U7164 (N_7164,N_6146,N_6819);
nand U7165 (N_7165,N_6309,N_6379);
nand U7166 (N_7166,N_6840,N_6767);
nor U7167 (N_7167,N_6732,N_6864);
nor U7168 (N_7168,N_6557,N_6871);
xnor U7169 (N_7169,N_6349,N_6537);
or U7170 (N_7170,N_6359,N_6602);
xor U7171 (N_7171,N_6821,N_6295);
xnor U7172 (N_7172,N_6887,N_6802);
nor U7173 (N_7173,N_6903,N_6524);
or U7174 (N_7174,N_6555,N_6455);
or U7175 (N_7175,N_6791,N_6880);
and U7176 (N_7176,N_6441,N_6402);
or U7177 (N_7177,N_6288,N_6885);
nand U7178 (N_7178,N_6852,N_6818);
xnor U7179 (N_7179,N_6208,N_6035);
and U7180 (N_7180,N_6166,N_6412);
xor U7181 (N_7181,N_6170,N_6138);
and U7182 (N_7182,N_6959,N_6010);
xnor U7183 (N_7183,N_6377,N_6152);
or U7184 (N_7184,N_6221,N_6827);
nor U7185 (N_7185,N_6204,N_6130);
nor U7186 (N_7186,N_6947,N_6958);
nor U7187 (N_7187,N_6996,N_6762);
nor U7188 (N_7188,N_6089,N_6194);
nand U7189 (N_7189,N_6809,N_6619);
nand U7190 (N_7190,N_6644,N_6338);
and U7191 (N_7191,N_6647,N_6203);
or U7192 (N_7192,N_6581,N_6107);
xor U7193 (N_7193,N_6164,N_6829);
and U7194 (N_7194,N_6105,N_6848);
and U7195 (N_7195,N_6378,N_6462);
or U7196 (N_7196,N_6962,N_6124);
and U7197 (N_7197,N_6276,N_6689);
xor U7198 (N_7198,N_6886,N_6753);
nor U7199 (N_7199,N_6653,N_6510);
and U7200 (N_7200,N_6768,N_6388);
or U7201 (N_7201,N_6244,N_6587);
nor U7202 (N_7202,N_6501,N_6961);
xnor U7203 (N_7203,N_6126,N_6031);
or U7204 (N_7204,N_6370,N_6070);
nor U7205 (N_7205,N_6580,N_6573);
or U7206 (N_7206,N_6845,N_6163);
nand U7207 (N_7207,N_6757,N_6718);
and U7208 (N_7208,N_6373,N_6937);
nor U7209 (N_7209,N_6974,N_6481);
nand U7210 (N_7210,N_6312,N_6115);
xnor U7211 (N_7211,N_6657,N_6252);
nand U7212 (N_7212,N_6103,N_6466);
and U7213 (N_7213,N_6617,N_6243);
and U7214 (N_7214,N_6242,N_6582);
nor U7215 (N_7215,N_6620,N_6113);
xnor U7216 (N_7216,N_6854,N_6469);
or U7217 (N_7217,N_6468,N_6180);
or U7218 (N_7218,N_6549,N_6135);
nand U7219 (N_7219,N_6683,N_6559);
nand U7220 (N_7220,N_6256,N_6003);
or U7221 (N_7221,N_6536,N_6376);
nand U7222 (N_7222,N_6982,N_6382);
nand U7223 (N_7223,N_6746,N_6999);
or U7224 (N_7224,N_6547,N_6004);
nor U7225 (N_7225,N_6470,N_6207);
nor U7226 (N_7226,N_6240,N_6765);
nor U7227 (N_7227,N_6727,N_6475);
nor U7228 (N_7228,N_6693,N_6733);
nand U7229 (N_7229,N_6842,N_6213);
xor U7230 (N_7230,N_6711,N_6502);
or U7231 (N_7231,N_6874,N_6304);
or U7232 (N_7232,N_6097,N_6161);
or U7233 (N_7233,N_6335,N_6696);
and U7234 (N_7234,N_6562,N_6892);
xor U7235 (N_7235,N_6626,N_6770);
nand U7236 (N_7236,N_6687,N_6042);
nor U7237 (N_7237,N_6328,N_6136);
or U7238 (N_7238,N_6342,N_6432);
nor U7239 (N_7239,N_6064,N_6021);
and U7240 (N_7240,N_6043,N_6153);
or U7241 (N_7241,N_6708,N_6910);
xnor U7242 (N_7242,N_6419,N_6527);
nand U7243 (N_7243,N_6876,N_6201);
or U7244 (N_7244,N_6453,N_6495);
nor U7245 (N_7245,N_6411,N_6079);
nor U7246 (N_7246,N_6568,N_6525);
or U7247 (N_7247,N_6979,N_6748);
and U7248 (N_7248,N_6464,N_6506);
or U7249 (N_7249,N_6571,N_6933);
and U7250 (N_7250,N_6804,N_6394);
or U7251 (N_7251,N_6262,N_6102);
nor U7252 (N_7252,N_6991,N_6258);
or U7253 (N_7253,N_6747,N_6709);
nor U7254 (N_7254,N_6543,N_6508);
or U7255 (N_7255,N_6722,N_6734);
and U7256 (N_7256,N_6778,N_6362);
and U7257 (N_7257,N_6544,N_6197);
xor U7258 (N_7258,N_6391,N_6645);
nor U7259 (N_7259,N_6448,N_6703);
xor U7260 (N_7260,N_6374,N_6896);
nor U7261 (N_7261,N_6128,N_6112);
xor U7262 (N_7262,N_6357,N_6133);
or U7263 (N_7263,N_6132,N_6094);
and U7264 (N_7264,N_6539,N_6333);
nor U7265 (N_7265,N_6480,N_6364);
nor U7266 (N_7266,N_6920,N_6117);
nand U7267 (N_7267,N_6946,N_6142);
or U7268 (N_7268,N_6049,N_6200);
and U7269 (N_7269,N_6145,N_6814);
or U7270 (N_7270,N_6039,N_6785);
or U7271 (N_7271,N_6289,N_6360);
nor U7272 (N_7272,N_6810,N_6667);
nand U7273 (N_7273,N_6741,N_6492);
nand U7274 (N_7274,N_6030,N_6792);
nand U7275 (N_7275,N_6255,N_6415);
or U7276 (N_7276,N_6638,N_6546);
nand U7277 (N_7277,N_6841,N_6801);
xnor U7278 (N_7278,N_6584,N_6596);
xnor U7279 (N_7279,N_6604,N_6123);
or U7280 (N_7280,N_6889,N_6598);
or U7281 (N_7281,N_6553,N_6608);
and U7282 (N_7282,N_6294,N_6673);
xor U7283 (N_7283,N_6729,N_6057);
nand U7284 (N_7284,N_6174,N_6229);
or U7285 (N_7285,N_6677,N_6578);
nand U7286 (N_7286,N_6269,N_6396);
nor U7287 (N_7287,N_6833,N_6088);
nand U7288 (N_7288,N_6849,N_6873);
or U7289 (N_7289,N_6942,N_6790);
and U7290 (N_7290,N_6375,N_6674);
or U7291 (N_7291,N_6157,N_6891);
nand U7292 (N_7292,N_6613,N_6230);
or U7293 (N_7293,N_6541,N_6389);
xnor U7294 (N_7294,N_6594,N_6784);
nor U7295 (N_7295,N_6056,N_6327);
nand U7296 (N_7296,N_6034,N_6217);
or U7297 (N_7297,N_6972,N_6472);
or U7298 (N_7298,N_6110,N_6040);
xor U7299 (N_7299,N_6955,N_6078);
nand U7300 (N_7300,N_6341,N_6296);
nand U7301 (N_7301,N_6234,N_6062);
xor U7302 (N_7302,N_6511,N_6090);
and U7303 (N_7303,N_6323,N_6228);
or U7304 (N_7304,N_6220,N_6313);
nand U7305 (N_7305,N_6983,N_6944);
and U7306 (N_7306,N_6701,N_6019);
nand U7307 (N_7307,N_6461,N_6465);
nor U7308 (N_7308,N_6330,N_6643);
nor U7309 (N_7309,N_6665,N_6308);
nor U7310 (N_7310,N_6787,N_6183);
and U7311 (N_7311,N_6096,N_6148);
nor U7312 (N_7312,N_6032,N_6755);
xor U7313 (N_7313,N_6828,N_6344);
nor U7314 (N_7314,N_6943,N_6303);
nor U7315 (N_7315,N_6368,N_6700);
and U7316 (N_7316,N_6279,N_6807);
nor U7317 (N_7317,N_6155,N_6224);
nor U7318 (N_7318,N_6731,N_6780);
and U7319 (N_7319,N_6984,N_6280);
xnor U7320 (N_7320,N_6509,N_6725);
nand U7321 (N_7321,N_6702,N_6825);
xnor U7322 (N_7322,N_6425,N_6726);
nand U7323 (N_7323,N_6505,N_6143);
and U7324 (N_7324,N_6149,N_6781);
and U7325 (N_7325,N_6951,N_6686);
and U7326 (N_7326,N_6478,N_6866);
and U7327 (N_7327,N_6554,N_6334);
or U7328 (N_7328,N_6275,N_6173);
xor U7329 (N_7329,N_6091,N_6668);
nor U7330 (N_7330,N_6084,N_6685);
or U7331 (N_7331,N_6487,N_6957);
or U7332 (N_7332,N_6835,N_6205);
nand U7333 (N_7333,N_6320,N_6381);
and U7334 (N_7334,N_6186,N_6385);
nand U7335 (N_7335,N_6712,N_6635);
or U7336 (N_7336,N_6851,N_6190);
nor U7337 (N_7337,N_6361,N_6222);
nor U7338 (N_7338,N_6651,N_6652);
nor U7339 (N_7339,N_6282,N_6329);
nand U7340 (N_7340,N_6339,N_6565);
xnor U7341 (N_7341,N_6656,N_6254);
nor U7342 (N_7342,N_6008,N_6650);
and U7343 (N_7343,N_6210,N_6857);
or U7344 (N_7344,N_6572,N_6872);
xor U7345 (N_7345,N_6884,N_6071);
xnor U7346 (N_7346,N_6490,N_6637);
nand U7347 (N_7347,N_6325,N_6369);
nor U7348 (N_7348,N_6987,N_6134);
nand U7349 (N_7349,N_6484,N_6915);
or U7350 (N_7350,N_6567,N_6345);
xor U7351 (N_7351,N_6060,N_6158);
or U7352 (N_7352,N_6366,N_6738);
nor U7353 (N_7353,N_6621,N_6678);
and U7354 (N_7354,N_6301,N_6893);
nand U7355 (N_7355,N_6844,N_6998);
nand U7356 (N_7356,N_6956,N_6754);
nand U7357 (N_7357,N_6436,N_6172);
nand U7358 (N_7358,N_6824,N_6531);
or U7359 (N_7359,N_6932,N_6054);
or U7360 (N_7360,N_6430,N_6290);
nor U7361 (N_7361,N_6952,N_6862);
and U7362 (N_7362,N_6023,N_6457);
or U7363 (N_7363,N_6574,N_6897);
nand U7364 (N_7364,N_6310,N_6198);
nand U7365 (N_7365,N_6264,N_6047);
nand U7366 (N_7366,N_6988,N_6101);
nor U7367 (N_7367,N_6837,N_6560);
nor U7368 (N_7368,N_6434,N_6779);
and U7369 (N_7369,N_6083,N_6805);
nand U7370 (N_7370,N_6684,N_6994);
nor U7371 (N_7371,N_6291,N_6027);
and U7372 (N_7372,N_6954,N_6215);
or U7373 (N_7373,N_6563,N_6209);
xor U7374 (N_7374,N_6050,N_6287);
nor U7375 (N_7375,N_6403,N_6281);
or U7376 (N_7376,N_6797,N_6899);
xnor U7377 (N_7377,N_6663,N_6392);
and U7378 (N_7378,N_6421,N_6795);
nor U7379 (N_7379,N_6014,N_6742);
nor U7380 (N_7380,N_6002,N_6950);
xnor U7381 (N_7381,N_6934,N_6211);
or U7382 (N_7382,N_6393,N_6263);
and U7383 (N_7383,N_6783,N_6570);
nand U7384 (N_7384,N_6086,N_6789);
xor U7385 (N_7385,N_6649,N_6267);
and U7386 (N_7386,N_6259,N_6763);
and U7387 (N_7387,N_6114,N_6771);
xnor U7388 (N_7388,N_6305,N_6488);
nor U7389 (N_7389,N_6989,N_6233);
nand U7390 (N_7390,N_6681,N_6073);
xor U7391 (N_7391,N_6398,N_6812);
nor U7392 (N_7392,N_6579,N_6076);
or U7393 (N_7393,N_6131,N_6277);
nand U7394 (N_7394,N_6625,N_6740);
nand U7395 (N_7395,N_6953,N_6680);
nor U7396 (N_7396,N_6628,N_6196);
nor U7397 (N_7397,N_6646,N_6929);
or U7398 (N_7398,N_6610,N_6597);
xnor U7399 (N_7399,N_6692,N_6337);
nand U7400 (N_7400,N_6600,N_6588);
or U7401 (N_7401,N_6006,N_6690);
nand U7402 (N_7402,N_6045,N_6085);
and U7403 (N_7403,N_6616,N_6065);
nor U7404 (N_7404,N_6640,N_6092);
and U7405 (N_7405,N_6975,N_6175);
nand U7406 (N_7406,N_6513,N_6523);
and U7407 (N_7407,N_6808,N_6482);
xor U7408 (N_7408,N_6966,N_6336);
xor U7409 (N_7409,N_6939,N_6995);
nor U7410 (N_7410,N_6516,N_6739);
xnor U7411 (N_7411,N_6705,N_6921);
nand U7412 (N_7412,N_6926,N_6351);
nor U7413 (N_7413,N_6458,N_6075);
and U7414 (N_7414,N_6435,N_6431);
or U7415 (N_7415,N_6253,N_6121);
nand U7416 (N_7416,N_6906,N_6397);
xnor U7417 (N_7417,N_6811,N_6592);
nor U7418 (N_7418,N_6545,N_6095);
or U7419 (N_7419,N_6022,N_6793);
xor U7420 (N_7420,N_6949,N_6445);
and U7421 (N_7421,N_6724,N_6331);
nand U7422 (N_7422,N_6454,N_6226);
nor U7423 (N_7423,N_6756,N_6504);
or U7424 (N_7424,N_6564,N_6241);
nor U7425 (N_7425,N_6575,N_6894);
nand U7426 (N_7426,N_6025,N_6150);
nand U7427 (N_7427,N_6750,N_6679);
nor U7428 (N_7428,N_6016,N_6911);
nand U7429 (N_7429,N_6426,N_6250);
nand U7430 (N_7430,N_6905,N_6437);
xor U7431 (N_7431,N_6566,N_6067);
nor U7432 (N_7432,N_6816,N_6878);
nand U7433 (N_7433,N_6069,N_6585);
or U7434 (N_7434,N_6188,N_6185);
and U7435 (N_7435,N_6879,N_6985);
nand U7436 (N_7436,N_6813,N_6913);
nand U7437 (N_7437,N_6898,N_6363);
and U7438 (N_7438,N_6390,N_6699);
nand U7439 (N_7439,N_6530,N_6526);
xor U7440 (N_7440,N_6371,N_6832);
xnor U7441 (N_7441,N_6569,N_6969);
xor U7442 (N_7442,N_6500,N_6238);
nor U7443 (N_7443,N_6017,N_6963);
nand U7444 (N_7444,N_6000,N_6285);
and U7445 (N_7445,N_6195,N_6538);
xor U7446 (N_7446,N_6922,N_6694);
or U7447 (N_7447,N_6786,N_6624);
nand U7448 (N_7448,N_6026,N_6675);
xnor U7449 (N_7449,N_6483,N_6521);
or U7450 (N_7450,N_6900,N_6980);
and U7451 (N_7451,N_6125,N_6160);
nor U7452 (N_7452,N_6648,N_6399);
or U7453 (N_7453,N_6704,N_6605);
nor U7454 (N_7454,N_6028,N_6931);
nand U7455 (N_7455,N_6817,N_6707);
or U7456 (N_7456,N_6127,N_6383);
nor U7457 (N_7457,N_6623,N_6413);
or U7458 (N_7458,N_6066,N_6960);
and U7459 (N_7459,N_6601,N_6137);
nor U7460 (N_7460,N_6018,N_6202);
and U7461 (N_7461,N_6716,N_6865);
xor U7462 (N_7462,N_6192,N_6735);
nand U7463 (N_7463,N_6494,N_6858);
nor U7464 (N_7464,N_6919,N_6671);
nor U7465 (N_7465,N_6847,N_6367);
xnor U7466 (N_7466,N_6548,N_6111);
nand U7467 (N_7467,N_6231,N_6636);
or U7468 (N_7468,N_6611,N_6895);
or U7469 (N_7469,N_6077,N_6446);
or U7470 (N_7470,N_6888,N_6474);
or U7471 (N_7471,N_6417,N_6806);
nand U7472 (N_7472,N_6507,N_6273);
or U7473 (N_7473,N_6322,N_6178);
xnor U7474 (N_7474,N_6861,N_6479);
nand U7475 (N_7475,N_6870,N_6720);
and U7476 (N_7476,N_6528,N_6247);
nor U7477 (N_7477,N_6093,N_6165);
xor U7478 (N_7478,N_6168,N_6629);
xor U7479 (N_7479,N_6855,N_6212);
xnor U7480 (N_7480,N_6935,N_6104);
or U7481 (N_7481,N_6100,N_6576);
nand U7482 (N_7482,N_6676,N_6968);
xor U7483 (N_7483,N_6058,N_6612);
and U7484 (N_7484,N_6451,N_6404);
nand U7485 (N_7485,N_6843,N_6347);
nor U7486 (N_7486,N_6977,N_6358);
xnor U7487 (N_7487,N_6883,N_6850);
and U7488 (N_7488,N_6423,N_6773);
and U7489 (N_7489,N_6443,N_6655);
nor U7490 (N_7490,N_6278,N_6286);
or U7491 (N_7491,N_6971,N_6407);
nand U7492 (N_7492,N_6219,N_6744);
nor U7493 (N_7493,N_6830,N_6477);
or U7494 (N_7494,N_6355,N_6976);
and U7495 (N_7495,N_6591,N_6428);
nor U7496 (N_7496,N_6449,N_6517);
nand U7497 (N_7497,N_6082,N_6688);
nand U7498 (N_7498,N_6639,N_6558);
nor U7499 (N_7499,N_6590,N_6838);
nand U7500 (N_7500,N_6348,N_6235);
or U7501 (N_7501,N_6522,N_6946);
xnor U7502 (N_7502,N_6333,N_6552);
nor U7503 (N_7503,N_6323,N_6098);
xor U7504 (N_7504,N_6724,N_6646);
nor U7505 (N_7505,N_6469,N_6417);
or U7506 (N_7506,N_6674,N_6034);
and U7507 (N_7507,N_6318,N_6970);
nor U7508 (N_7508,N_6545,N_6357);
xnor U7509 (N_7509,N_6385,N_6822);
nand U7510 (N_7510,N_6061,N_6582);
or U7511 (N_7511,N_6070,N_6431);
and U7512 (N_7512,N_6361,N_6736);
nor U7513 (N_7513,N_6800,N_6612);
nand U7514 (N_7514,N_6926,N_6617);
nand U7515 (N_7515,N_6933,N_6293);
xnor U7516 (N_7516,N_6714,N_6234);
and U7517 (N_7517,N_6110,N_6939);
or U7518 (N_7518,N_6856,N_6715);
xnor U7519 (N_7519,N_6950,N_6496);
nor U7520 (N_7520,N_6115,N_6628);
nand U7521 (N_7521,N_6064,N_6203);
xor U7522 (N_7522,N_6626,N_6231);
nor U7523 (N_7523,N_6491,N_6433);
nor U7524 (N_7524,N_6623,N_6801);
or U7525 (N_7525,N_6941,N_6755);
xor U7526 (N_7526,N_6865,N_6114);
and U7527 (N_7527,N_6488,N_6742);
nand U7528 (N_7528,N_6966,N_6555);
nand U7529 (N_7529,N_6757,N_6537);
nor U7530 (N_7530,N_6246,N_6838);
or U7531 (N_7531,N_6326,N_6615);
or U7532 (N_7532,N_6100,N_6099);
and U7533 (N_7533,N_6227,N_6854);
nor U7534 (N_7534,N_6873,N_6507);
nor U7535 (N_7535,N_6918,N_6024);
and U7536 (N_7536,N_6061,N_6471);
nand U7537 (N_7537,N_6031,N_6678);
xor U7538 (N_7538,N_6912,N_6536);
nand U7539 (N_7539,N_6639,N_6865);
nand U7540 (N_7540,N_6196,N_6262);
or U7541 (N_7541,N_6509,N_6478);
nor U7542 (N_7542,N_6318,N_6538);
nand U7543 (N_7543,N_6430,N_6979);
xor U7544 (N_7544,N_6954,N_6288);
and U7545 (N_7545,N_6526,N_6228);
nand U7546 (N_7546,N_6855,N_6293);
or U7547 (N_7547,N_6702,N_6352);
and U7548 (N_7548,N_6097,N_6577);
nor U7549 (N_7549,N_6487,N_6513);
nand U7550 (N_7550,N_6864,N_6380);
xnor U7551 (N_7551,N_6642,N_6697);
nor U7552 (N_7552,N_6227,N_6667);
nand U7553 (N_7553,N_6399,N_6157);
xnor U7554 (N_7554,N_6677,N_6787);
nand U7555 (N_7555,N_6647,N_6115);
nand U7556 (N_7556,N_6621,N_6438);
or U7557 (N_7557,N_6598,N_6934);
nand U7558 (N_7558,N_6419,N_6605);
or U7559 (N_7559,N_6836,N_6181);
xor U7560 (N_7560,N_6278,N_6583);
or U7561 (N_7561,N_6753,N_6653);
nand U7562 (N_7562,N_6710,N_6485);
nor U7563 (N_7563,N_6735,N_6181);
nand U7564 (N_7564,N_6427,N_6213);
and U7565 (N_7565,N_6500,N_6941);
and U7566 (N_7566,N_6055,N_6601);
nand U7567 (N_7567,N_6729,N_6843);
or U7568 (N_7568,N_6256,N_6460);
nand U7569 (N_7569,N_6689,N_6583);
nor U7570 (N_7570,N_6991,N_6748);
nor U7571 (N_7571,N_6339,N_6889);
nor U7572 (N_7572,N_6662,N_6486);
or U7573 (N_7573,N_6748,N_6970);
or U7574 (N_7574,N_6256,N_6449);
nor U7575 (N_7575,N_6113,N_6739);
nand U7576 (N_7576,N_6649,N_6638);
and U7577 (N_7577,N_6517,N_6484);
xor U7578 (N_7578,N_6421,N_6191);
nand U7579 (N_7579,N_6596,N_6899);
xnor U7580 (N_7580,N_6754,N_6964);
or U7581 (N_7581,N_6894,N_6968);
nand U7582 (N_7582,N_6562,N_6001);
nand U7583 (N_7583,N_6646,N_6180);
or U7584 (N_7584,N_6163,N_6513);
or U7585 (N_7585,N_6209,N_6504);
and U7586 (N_7586,N_6982,N_6251);
nor U7587 (N_7587,N_6217,N_6009);
nand U7588 (N_7588,N_6111,N_6194);
nor U7589 (N_7589,N_6322,N_6259);
and U7590 (N_7590,N_6408,N_6198);
nor U7591 (N_7591,N_6489,N_6499);
nor U7592 (N_7592,N_6085,N_6783);
or U7593 (N_7593,N_6836,N_6113);
and U7594 (N_7594,N_6193,N_6667);
and U7595 (N_7595,N_6062,N_6538);
or U7596 (N_7596,N_6643,N_6288);
nor U7597 (N_7597,N_6592,N_6371);
nand U7598 (N_7598,N_6699,N_6571);
and U7599 (N_7599,N_6889,N_6860);
or U7600 (N_7600,N_6092,N_6404);
xnor U7601 (N_7601,N_6030,N_6851);
and U7602 (N_7602,N_6240,N_6846);
nor U7603 (N_7603,N_6201,N_6939);
xnor U7604 (N_7604,N_6405,N_6202);
nand U7605 (N_7605,N_6762,N_6624);
and U7606 (N_7606,N_6985,N_6750);
or U7607 (N_7607,N_6551,N_6750);
nor U7608 (N_7608,N_6091,N_6855);
and U7609 (N_7609,N_6363,N_6413);
nand U7610 (N_7610,N_6177,N_6759);
xor U7611 (N_7611,N_6578,N_6010);
and U7612 (N_7612,N_6482,N_6723);
nand U7613 (N_7613,N_6601,N_6798);
nor U7614 (N_7614,N_6729,N_6594);
xnor U7615 (N_7615,N_6998,N_6399);
or U7616 (N_7616,N_6250,N_6016);
or U7617 (N_7617,N_6341,N_6325);
and U7618 (N_7618,N_6032,N_6581);
or U7619 (N_7619,N_6442,N_6318);
or U7620 (N_7620,N_6131,N_6436);
nor U7621 (N_7621,N_6701,N_6533);
nand U7622 (N_7622,N_6051,N_6520);
or U7623 (N_7623,N_6650,N_6330);
nand U7624 (N_7624,N_6066,N_6910);
xnor U7625 (N_7625,N_6729,N_6983);
nor U7626 (N_7626,N_6958,N_6354);
nand U7627 (N_7627,N_6323,N_6010);
nor U7628 (N_7628,N_6075,N_6926);
nand U7629 (N_7629,N_6942,N_6072);
and U7630 (N_7630,N_6040,N_6946);
xor U7631 (N_7631,N_6814,N_6694);
xnor U7632 (N_7632,N_6525,N_6764);
and U7633 (N_7633,N_6982,N_6936);
nor U7634 (N_7634,N_6823,N_6856);
or U7635 (N_7635,N_6502,N_6364);
nand U7636 (N_7636,N_6446,N_6709);
xor U7637 (N_7637,N_6935,N_6570);
and U7638 (N_7638,N_6872,N_6731);
and U7639 (N_7639,N_6288,N_6961);
nor U7640 (N_7640,N_6397,N_6517);
nand U7641 (N_7641,N_6369,N_6196);
or U7642 (N_7642,N_6629,N_6997);
nand U7643 (N_7643,N_6632,N_6834);
nand U7644 (N_7644,N_6632,N_6010);
nor U7645 (N_7645,N_6602,N_6601);
or U7646 (N_7646,N_6672,N_6934);
xnor U7647 (N_7647,N_6799,N_6097);
nand U7648 (N_7648,N_6757,N_6684);
nand U7649 (N_7649,N_6215,N_6728);
xor U7650 (N_7650,N_6706,N_6980);
xor U7651 (N_7651,N_6737,N_6515);
or U7652 (N_7652,N_6246,N_6573);
xor U7653 (N_7653,N_6228,N_6658);
and U7654 (N_7654,N_6828,N_6746);
nor U7655 (N_7655,N_6423,N_6145);
nand U7656 (N_7656,N_6479,N_6239);
or U7657 (N_7657,N_6782,N_6370);
xor U7658 (N_7658,N_6490,N_6557);
and U7659 (N_7659,N_6087,N_6955);
or U7660 (N_7660,N_6546,N_6841);
and U7661 (N_7661,N_6360,N_6781);
and U7662 (N_7662,N_6761,N_6025);
or U7663 (N_7663,N_6207,N_6959);
nand U7664 (N_7664,N_6791,N_6064);
or U7665 (N_7665,N_6708,N_6902);
or U7666 (N_7666,N_6054,N_6110);
nor U7667 (N_7667,N_6130,N_6636);
nor U7668 (N_7668,N_6726,N_6064);
and U7669 (N_7669,N_6529,N_6384);
or U7670 (N_7670,N_6123,N_6900);
nand U7671 (N_7671,N_6573,N_6293);
nand U7672 (N_7672,N_6485,N_6222);
or U7673 (N_7673,N_6888,N_6032);
and U7674 (N_7674,N_6703,N_6142);
xnor U7675 (N_7675,N_6120,N_6858);
nor U7676 (N_7676,N_6223,N_6506);
or U7677 (N_7677,N_6281,N_6769);
or U7678 (N_7678,N_6534,N_6162);
xor U7679 (N_7679,N_6877,N_6549);
xor U7680 (N_7680,N_6640,N_6458);
nor U7681 (N_7681,N_6013,N_6010);
or U7682 (N_7682,N_6186,N_6031);
and U7683 (N_7683,N_6313,N_6818);
nor U7684 (N_7684,N_6296,N_6635);
and U7685 (N_7685,N_6185,N_6637);
nand U7686 (N_7686,N_6169,N_6539);
and U7687 (N_7687,N_6452,N_6765);
nor U7688 (N_7688,N_6341,N_6044);
and U7689 (N_7689,N_6961,N_6598);
nand U7690 (N_7690,N_6097,N_6686);
or U7691 (N_7691,N_6819,N_6149);
or U7692 (N_7692,N_6034,N_6315);
nand U7693 (N_7693,N_6977,N_6505);
and U7694 (N_7694,N_6107,N_6279);
nand U7695 (N_7695,N_6847,N_6315);
nor U7696 (N_7696,N_6323,N_6994);
nand U7697 (N_7697,N_6117,N_6901);
and U7698 (N_7698,N_6100,N_6487);
or U7699 (N_7699,N_6443,N_6116);
nand U7700 (N_7700,N_6699,N_6973);
nand U7701 (N_7701,N_6662,N_6898);
xor U7702 (N_7702,N_6468,N_6930);
nand U7703 (N_7703,N_6699,N_6244);
and U7704 (N_7704,N_6350,N_6446);
nand U7705 (N_7705,N_6318,N_6515);
nor U7706 (N_7706,N_6240,N_6353);
xor U7707 (N_7707,N_6136,N_6046);
nor U7708 (N_7708,N_6535,N_6018);
or U7709 (N_7709,N_6001,N_6744);
xor U7710 (N_7710,N_6046,N_6208);
nand U7711 (N_7711,N_6726,N_6680);
nor U7712 (N_7712,N_6147,N_6391);
or U7713 (N_7713,N_6124,N_6547);
nor U7714 (N_7714,N_6421,N_6582);
nor U7715 (N_7715,N_6373,N_6089);
and U7716 (N_7716,N_6745,N_6514);
nand U7717 (N_7717,N_6166,N_6538);
nand U7718 (N_7718,N_6192,N_6708);
or U7719 (N_7719,N_6601,N_6019);
or U7720 (N_7720,N_6700,N_6238);
nand U7721 (N_7721,N_6398,N_6755);
nand U7722 (N_7722,N_6937,N_6621);
xnor U7723 (N_7723,N_6823,N_6097);
xnor U7724 (N_7724,N_6070,N_6288);
nor U7725 (N_7725,N_6714,N_6200);
xnor U7726 (N_7726,N_6819,N_6742);
and U7727 (N_7727,N_6640,N_6995);
and U7728 (N_7728,N_6414,N_6734);
nand U7729 (N_7729,N_6958,N_6774);
xnor U7730 (N_7730,N_6717,N_6881);
or U7731 (N_7731,N_6660,N_6675);
nand U7732 (N_7732,N_6361,N_6280);
xnor U7733 (N_7733,N_6494,N_6830);
or U7734 (N_7734,N_6317,N_6044);
or U7735 (N_7735,N_6536,N_6015);
or U7736 (N_7736,N_6730,N_6106);
or U7737 (N_7737,N_6573,N_6701);
or U7738 (N_7738,N_6867,N_6677);
and U7739 (N_7739,N_6181,N_6693);
and U7740 (N_7740,N_6152,N_6942);
xor U7741 (N_7741,N_6940,N_6742);
nand U7742 (N_7742,N_6588,N_6060);
nand U7743 (N_7743,N_6077,N_6187);
nor U7744 (N_7744,N_6235,N_6916);
nor U7745 (N_7745,N_6969,N_6231);
or U7746 (N_7746,N_6895,N_6261);
nor U7747 (N_7747,N_6300,N_6781);
xnor U7748 (N_7748,N_6133,N_6534);
nand U7749 (N_7749,N_6238,N_6980);
and U7750 (N_7750,N_6326,N_6565);
xnor U7751 (N_7751,N_6574,N_6726);
and U7752 (N_7752,N_6384,N_6639);
and U7753 (N_7753,N_6089,N_6256);
xor U7754 (N_7754,N_6137,N_6682);
and U7755 (N_7755,N_6718,N_6904);
or U7756 (N_7756,N_6353,N_6389);
nor U7757 (N_7757,N_6444,N_6188);
and U7758 (N_7758,N_6432,N_6020);
and U7759 (N_7759,N_6964,N_6752);
nand U7760 (N_7760,N_6138,N_6388);
or U7761 (N_7761,N_6527,N_6454);
nor U7762 (N_7762,N_6100,N_6333);
nand U7763 (N_7763,N_6793,N_6755);
nand U7764 (N_7764,N_6212,N_6025);
or U7765 (N_7765,N_6436,N_6486);
and U7766 (N_7766,N_6658,N_6185);
xnor U7767 (N_7767,N_6903,N_6324);
xnor U7768 (N_7768,N_6737,N_6141);
nand U7769 (N_7769,N_6809,N_6450);
xor U7770 (N_7770,N_6809,N_6001);
or U7771 (N_7771,N_6987,N_6126);
and U7772 (N_7772,N_6245,N_6944);
xor U7773 (N_7773,N_6725,N_6476);
and U7774 (N_7774,N_6518,N_6275);
nor U7775 (N_7775,N_6058,N_6708);
and U7776 (N_7776,N_6792,N_6384);
nor U7777 (N_7777,N_6824,N_6845);
xor U7778 (N_7778,N_6686,N_6687);
nand U7779 (N_7779,N_6122,N_6397);
nor U7780 (N_7780,N_6575,N_6825);
or U7781 (N_7781,N_6083,N_6516);
and U7782 (N_7782,N_6290,N_6163);
or U7783 (N_7783,N_6994,N_6266);
and U7784 (N_7784,N_6990,N_6160);
nor U7785 (N_7785,N_6467,N_6640);
xor U7786 (N_7786,N_6526,N_6943);
or U7787 (N_7787,N_6853,N_6542);
xnor U7788 (N_7788,N_6589,N_6968);
and U7789 (N_7789,N_6355,N_6520);
nand U7790 (N_7790,N_6403,N_6852);
xnor U7791 (N_7791,N_6415,N_6923);
nand U7792 (N_7792,N_6693,N_6183);
nand U7793 (N_7793,N_6275,N_6075);
and U7794 (N_7794,N_6377,N_6925);
nand U7795 (N_7795,N_6194,N_6977);
nor U7796 (N_7796,N_6595,N_6885);
nand U7797 (N_7797,N_6833,N_6025);
xor U7798 (N_7798,N_6278,N_6909);
nor U7799 (N_7799,N_6093,N_6798);
or U7800 (N_7800,N_6202,N_6861);
nor U7801 (N_7801,N_6187,N_6371);
or U7802 (N_7802,N_6854,N_6947);
nand U7803 (N_7803,N_6988,N_6997);
and U7804 (N_7804,N_6760,N_6172);
nor U7805 (N_7805,N_6566,N_6227);
xor U7806 (N_7806,N_6043,N_6755);
xor U7807 (N_7807,N_6554,N_6183);
and U7808 (N_7808,N_6642,N_6006);
and U7809 (N_7809,N_6578,N_6744);
nand U7810 (N_7810,N_6435,N_6798);
nor U7811 (N_7811,N_6817,N_6057);
or U7812 (N_7812,N_6741,N_6758);
or U7813 (N_7813,N_6007,N_6128);
and U7814 (N_7814,N_6381,N_6183);
nor U7815 (N_7815,N_6904,N_6627);
nand U7816 (N_7816,N_6063,N_6720);
nor U7817 (N_7817,N_6664,N_6863);
xor U7818 (N_7818,N_6494,N_6197);
nand U7819 (N_7819,N_6252,N_6199);
nand U7820 (N_7820,N_6708,N_6142);
or U7821 (N_7821,N_6377,N_6806);
nor U7822 (N_7822,N_6922,N_6966);
or U7823 (N_7823,N_6104,N_6199);
xor U7824 (N_7824,N_6045,N_6185);
or U7825 (N_7825,N_6805,N_6893);
and U7826 (N_7826,N_6516,N_6388);
nor U7827 (N_7827,N_6263,N_6165);
or U7828 (N_7828,N_6785,N_6489);
nor U7829 (N_7829,N_6598,N_6574);
xor U7830 (N_7830,N_6417,N_6816);
nand U7831 (N_7831,N_6402,N_6767);
xnor U7832 (N_7832,N_6885,N_6984);
nor U7833 (N_7833,N_6508,N_6440);
nand U7834 (N_7834,N_6570,N_6276);
or U7835 (N_7835,N_6480,N_6232);
xor U7836 (N_7836,N_6851,N_6551);
nand U7837 (N_7837,N_6015,N_6269);
or U7838 (N_7838,N_6588,N_6105);
and U7839 (N_7839,N_6824,N_6571);
xor U7840 (N_7840,N_6597,N_6839);
or U7841 (N_7841,N_6604,N_6354);
nand U7842 (N_7842,N_6347,N_6906);
and U7843 (N_7843,N_6825,N_6164);
nand U7844 (N_7844,N_6028,N_6982);
xor U7845 (N_7845,N_6274,N_6125);
xnor U7846 (N_7846,N_6076,N_6306);
nor U7847 (N_7847,N_6382,N_6462);
nand U7848 (N_7848,N_6273,N_6421);
nand U7849 (N_7849,N_6756,N_6031);
xnor U7850 (N_7850,N_6678,N_6471);
and U7851 (N_7851,N_6141,N_6212);
nor U7852 (N_7852,N_6644,N_6953);
or U7853 (N_7853,N_6390,N_6696);
nand U7854 (N_7854,N_6500,N_6769);
nand U7855 (N_7855,N_6841,N_6315);
xnor U7856 (N_7856,N_6953,N_6309);
nand U7857 (N_7857,N_6970,N_6179);
xnor U7858 (N_7858,N_6651,N_6981);
nor U7859 (N_7859,N_6765,N_6850);
nor U7860 (N_7860,N_6633,N_6058);
nand U7861 (N_7861,N_6163,N_6400);
nand U7862 (N_7862,N_6637,N_6840);
and U7863 (N_7863,N_6682,N_6029);
xor U7864 (N_7864,N_6695,N_6422);
nand U7865 (N_7865,N_6479,N_6791);
xnor U7866 (N_7866,N_6691,N_6379);
nor U7867 (N_7867,N_6842,N_6279);
xnor U7868 (N_7868,N_6942,N_6136);
nor U7869 (N_7869,N_6799,N_6548);
and U7870 (N_7870,N_6787,N_6779);
xnor U7871 (N_7871,N_6098,N_6033);
and U7872 (N_7872,N_6936,N_6250);
and U7873 (N_7873,N_6331,N_6623);
and U7874 (N_7874,N_6726,N_6795);
or U7875 (N_7875,N_6274,N_6490);
nor U7876 (N_7876,N_6498,N_6382);
nand U7877 (N_7877,N_6399,N_6126);
nand U7878 (N_7878,N_6960,N_6063);
nand U7879 (N_7879,N_6216,N_6201);
and U7880 (N_7880,N_6002,N_6925);
and U7881 (N_7881,N_6432,N_6030);
or U7882 (N_7882,N_6263,N_6124);
xor U7883 (N_7883,N_6342,N_6231);
xnor U7884 (N_7884,N_6935,N_6096);
xor U7885 (N_7885,N_6260,N_6478);
xor U7886 (N_7886,N_6551,N_6041);
or U7887 (N_7887,N_6726,N_6922);
nand U7888 (N_7888,N_6948,N_6719);
nand U7889 (N_7889,N_6051,N_6759);
nand U7890 (N_7890,N_6667,N_6511);
nor U7891 (N_7891,N_6019,N_6418);
xor U7892 (N_7892,N_6059,N_6757);
and U7893 (N_7893,N_6096,N_6853);
or U7894 (N_7894,N_6479,N_6988);
nor U7895 (N_7895,N_6239,N_6028);
or U7896 (N_7896,N_6705,N_6309);
nor U7897 (N_7897,N_6237,N_6778);
or U7898 (N_7898,N_6294,N_6221);
nor U7899 (N_7899,N_6806,N_6199);
nor U7900 (N_7900,N_6115,N_6812);
nor U7901 (N_7901,N_6251,N_6508);
or U7902 (N_7902,N_6092,N_6435);
and U7903 (N_7903,N_6404,N_6128);
xnor U7904 (N_7904,N_6344,N_6598);
and U7905 (N_7905,N_6252,N_6117);
nand U7906 (N_7906,N_6563,N_6371);
nor U7907 (N_7907,N_6434,N_6135);
xnor U7908 (N_7908,N_6659,N_6217);
and U7909 (N_7909,N_6052,N_6648);
xor U7910 (N_7910,N_6162,N_6252);
nand U7911 (N_7911,N_6009,N_6050);
nand U7912 (N_7912,N_6755,N_6442);
or U7913 (N_7913,N_6796,N_6055);
or U7914 (N_7914,N_6638,N_6496);
xnor U7915 (N_7915,N_6418,N_6666);
nand U7916 (N_7916,N_6150,N_6966);
and U7917 (N_7917,N_6100,N_6256);
nor U7918 (N_7918,N_6534,N_6721);
nand U7919 (N_7919,N_6582,N_6977);
nor U7920 (N_7920,N_6675,N_6539);
or U7921 (N_7921,N_6022,N_6884);
and U7922 (N_7922,N_6214,N_6806);
and U7923 (N_7923,N_6121,N_6228);
or U7924 (N_7924,N_6032,N_6162);
or U7925 (N_7925,N_6701,N_6519);
nand U7926 (N_7926,N_6816,N_6038);
nand U7927 (N_7927,N_6271,N_6631);
xnor U7928 (N_7928,N_6080,N_6999);
or U7929 (N_7929,N_6789,N_6409);
nor U7930 (N_7930,N_6273,N_6704);
or U7931 (N_7931,N_6473,N_6871);
and U7932 (N_7932,N_6356,N_6576);
and U7933 (N_7933,N_6079,N_6905);
nor U7934 (N_7934,N_6433,N_6056);
nor U7935 (N_7935,N_6500,N_6671);
or U7936 (N_7936,N_6208,N_6031);
or U7937 (N_7937,N_6613,N_6662);
and U7938 (N_7938,N_6359,N_6639);
nand U7939 (N_7939,N_6435,N_6445);
and U7940 (N_7940,N_6279,N_6934);
xor U7941 (N_7941,N_6793,N_6939);
nand U7942 (N_7942,N_6573,N_6191);
or U7943 (N_7943,N_6527,N_6015);
xnor U7944 (N_7944,N_6673,N_6442);
nand U7945 (N_7945,N_6920,N_6456);
nand U7946 (N_7946,N_6762,N_6887);
or U7947 (N_7947,N_6841,N_6523);
or U7948 (N_7948,N_6719,N_6219);
and U7949 (N_7949,N_6827,N_6599);
nor U7950 (N_7950,N_6320,N_6165);
nand U7951 (N_7951,N_6010,N_6574);
xnor U7952 (N_7952,N_6828,N_6260);
or U7953 (N_7953,N_6450,N_6830);
xnor U7954 (N_7954,N_6702,N_6687);
nor U7955 (N_7955,N_6603,N_6927);
nand U7956 (N_7956,N_6355,N_6714);
xor U7957 (N_7957,N_6244,N_6503);
or U7958 (N_7958,N_6700,N_6247);
or U7959 (N_7959,N_6586,N_6250);
or U7960 (N_7960,N_6920,N_6843);
or U7961 (N_7961,N_6009,N_6902);
xor U7962 (N_7962,N_6306,N_6913);
nand U7963 (N_7963,N_6291,N_6759);
and U7964 (N_7964,N_6462,N_6984);
nand U7965 (N_7965,N_6472,N_6879);
or U7966 (N_7966,N_6496,N_6492);
xnor U7967 (N_7967,N_6921,N_6484);
xnor U7968 (N_7968,N_6761,N_6296);
nand U7969 (N_7969,N_6560,N_6818);
nor U7970 (N_7970,N_6479,N_6554);
or U7971 (N_7971,N_6718,N_6232);
nor U7972 (N_7972,N_6103,N_6855);
or U7973 (N_7973,N_6579,N_6687);
xor U7974 (N_7974,N_6664,N_6086);
nor U7975 (N_7975,N_6724,N_6215);
and U7976 (N_7976,N_6107,N_6008);
xnor U7977 (N_7977,N_6694,N_6628);
nand U7978 (N_7978,N_6728,N_6075);
nor U7979 (N_7979,N_6156,N_6494);
or U7980 (N_7980,N_6611,N_6932);
xnor U7981 (N_7981,N_6187,N_6255);
nor U7982 (N_7982,N_6956,N_6276);
or U7983 (N_7983,N_6679,N_6452);
or U7984 (N_7984,N_6749,N_6294);
and U7985 (N_7985,N_6124,N_6893);
xor U7986 (N_7986,N_6164,N_6690);
nor U7987 (N_7987,N_6466,N_6680);
nor U7988 (N_7988,N_6407,N_6893);
or U7989 (N_7989,N_6075,N_6552);
xor U7990 (N_7990,N_6356,N_6771);
nor U7991 (N_7991,N_6485,N_6928);
nor U7992 (N_7992,N_6098,N_6253);
nor U7993 (N_7993,N_6565,N_6873);
nor U7994 (N_7994,N_6909,N_6041);
or U7995 (N_7995,N_6642,N_6878);
nor U7996 (N_7996,N_6051,N_6529);
or U7997 (N_7997,N_6564,N_6576);
nand U7998 (N_7998,N_6649,N_6864);
or U7999 (N_7999,N_6734,N_6516);
nor U8000 (N_8000,N_7162,N_7744);
xor U8001 (N_8001,N_7010,N_7759);
nor U8002 (N_8002,N_7555,N_7218);
xnor U8003 (N_8003,N_7772,N_7845);
xor U8004 (N_8004,N_7444,N_7850);
nor U8005 (N_8005,N_7078,N_7748);
or U8006 (N_8006,N_7344,N_7229);
xnor U8007 (N_8007,N_7724,N_7276);
nor U8008 (N_8008,N_7102,N_7662);
nor U8009 (N_8009,N_7129,N_7397);
nand U8010 (N_8010,N_7996,N_7970);
nor U8011 (N_8011,N_7709,N_7428);
nor U8012 (N_8012,N_7161,N_7495);
or U8013 (N_8013,N_7360,N_7095);
or U8014 (N_8014,N_7238,N_7223);
xnor U8015 (N_8015,N_7215,N_7658);
or U8016 (N_8016,N_7034,N_7666);
and U8017 (N_8017,N_7565,N_7804);
xnor U8018 (N_8018,N_7227,N_7522);
and U8019 (N_8019,N_7037,N_7336);
or U8020 (N_8020,N_7571,N_7028);
xnor U8021 (N_8021,N_7601,N_7096);
nand U8022 (N_8022,N_7306,N_7511);
xnor U8023 (N_8023,N_7520,N_7889);
or U8024 (N_8024,N_7137,N_7974);
nor U8025 (N_8025,N_7813,N_7041);
nand U8026 (N_8026,N_7901,N_7530);
and U8027 (N_8027,N_7870,N_7302);
and U8028 (N_8028,N_7543,N_7998);
nor U8029 (N_8029,N_7320,N_7125);
nand U8030 (N_8030,N_7688,N_7613);
and U8031 (N_8031,N_7127,N_7819);
nand U8032 (N_8032,N_7443,N_7358);
xor U8033 (N_8033,N_7698,N_7062);
and U8034 (N_8034,N_7986,N_7001);
and U8035 (N_8035,N_7859,N_7132);
xnor U8036 (N_8036,N_7179,N_7875);
xor U8037 (N_8037,N_7529,N_7664);
nor U8038 (N_8038,N_7092,N_7867);
and U8039 (N_8039,N_7059,N_7591);
or U8040 (N_8040,N_7676,N_7356);
or U8041 (N_8041,N_7071,N_7145);
or U8042 (N_8042,N_7108,N_7960);
nor U8043 (N_8043,N_7536,N_7372);
or U8044 (N_8044,N_7888,N_7142);
nor U8045 (N_8045,N_7131,N_7368);
nor U8046 (N_8046,N_7708,N_7098);
and U8047 (N_8047,N_7439,N_7113);
and U8048 (N_8048,N_7089,N_7749);
nor U8049 (N_8049,N_7138,N_7479);
or U8050 (N_8050,N_7921,N_7279);
nor U8051 (N_8051,N_7902,N_7349);
nor U8052 (N_8052,N_7296,N_7419);
and U8053 (N_8053,N_7564,N_7180);
or U8054 (N_8054,N_7115,N_7105);
and U8055 (N_8055,N_7795,N_7788);
or U8056 (N_8056,N_7898,N_7166);
and U8057 (N_8057,N_7422,N_7021);
nand U8058 (N_8058,N_7140,N_7608);
or U8059 (N_8059,N_7736,N_7348);
and U8060 (N_8060,N_7371,N_7618);
or U8061 (N_8061,N_7810,N_7820);
xnor U8062 (N_8062,N_7539,N_7080);
xnor U8063 (N_8063,N_7169,N_7338);
or U8064 (N_8064,N_7391,N_7032);
xor U8065 (N_8065,N_7009,N_7049);
nor U8066 (N_8066,N_7833,N_7713);
or U8067 (N_8067,N_7677,N_7993);
xnor U8068 (N_8068,N_7815,N_7366);
xnor U8069 (N_8069,N_7044,N_7357);
xnor U8070 (N_8070,N_7074,N_7103);
or U8071 (N_8071,N_7375,N_7863);
or U8072 (N_8072,N_7082,N_7448);
or U8073 (N_8073,N_7752,N_7560);
xor U8074 (N_8074,N_7421,N_7058);
nor U8075 (N_8075,N_7959,N_7350);
nor U8076 (N_8076,N_7864,N_7346);
or U8077 (N_8077,N_7650,N_7274);
nor U8078 (N_8078,N_7455,N_7353);
and U8079 (N_8079,N_7226,N_7172);
or U8080 (N_8080,N_7470,N_7068);
xnor U8081 (N_8081,N_7013,N_7139);
or U8082 (N_8082,N_7471,N_7619);
or U8083 (N_8083,N_7042,N_7386);
or U8084 (N_8084,N_7466,N_7681);
xor U8085 (N_8085,N_7485,N_7484);
xor U8086 (N_8086,N_7237,N_7355);
xnor U8087 (N_8087,N_7019,N_7198);
xnor U8088 (N_8088,N_7966,N_7651);
or U8089 (N_8089,N_7119,N_7763);
and U8090 (N_8090,N_7908,N_7678);
and U8091 (N_8091,N_7114,N_7278);
and U8092 (N_8092,N_7794,N_7155);
nand U8093 (N_8093,N_7652,N_7186);
or U8094 (N_8094,N_7896,N_7519);
or U8095 (N_8095,N_7580,N_7527);
xnor U8096 (N_8096,N_7880,N_7022);
and U8097 (N_8097,N_7656,N_7200);
and U8098 (N_8098,N_7906,N_7853);
and U8099 (N_8099,N_7997,N_7628);
and U8100 (N_8100,N_7508,N_7644);
or U8101 (N_8101,N_7924,N_7909);
nand U8102 (N_8102,N_7240,N_7154);
and U8103 (N_8103,N_7940,N_7351);
xnor U8104 (N_8104,N_7712,N_7693);
nand U8105 (N_8105,N_7282,N_7367);
and U8106 (N_8106,N_7012,N_7039);
and U8107 (N_8107,N_7680,N_7827);
nand U8108 (N_8108,N_7634,N_7980);
and U8109 (N_8109,N_7562,N_7181);
nand U8110 (N_8110,N_7463,N_7595);
nand U8111 (N_8111,N_7531,N_7257);
xnor U8112 (N_8112,N_7232,N_7177);
nor U8113 (N_8113,N_7070,N_7394);
or U8114 (N_8114,N_7510,N_7047);
and U8115 (N_8115,N_7755,N_7625);
or U8116 (N_8116,N_7493,N_7590);
nor U8117 (N_8117,N_7064,N_7729);
nand U8118 (N_8118,N_7566,N_7382);
or U8119 (N_8119,N_7572,N_7739);
nor U8120 (N_8120,N_7874,N_7799);
or U8121 (N_8121,N_7483,N_7597);
nor U8122 (N_8122,N_7961,N_7361);
xor U8123 (N_8123,N_7574,N_7459);
and U8124 (N_8124,N_7319,N_7660);
or U8125 (N_8125,N_7018,N_7971);
nand U8126 (N_8126,N_7433,N_7876);
nor U8127 (N_8127,N_7609,N_7538);
or U8128 (N_8128,N_7554,N_7899);
xnor U8129 (N_8129,N_7411,N_7723);
or U8130 (N_8130,N_7937,N_7745);
nor U8131 (N_8131,N_7976,N_7923);
nand U8132 (N_8132,N_7434,N_7480);
and U8133 (N_8133,N_7501,N_7380);
xor U8134 (N_8134,N_7280,N_7751);
nand U8135 (N_8135,N_7482,N_7486);
xnor U8136 (N_8136,N_7373,N_7249);
nand U8137 (N_8137,N_7189,N_7738);
or U8138 (N_8138,N_7151,N_7488);
and U8139 (N_8139,N_7667,N_7825);
nor U8140 (N_8140,N_7582,N_7904);
or U8141 (N_8141,N_7461,N_7570);
xor U8142 (N_8142,N_7984,N_7231);
or U8143 (N_8143,N_7728,N_7526);
and U8144 (N_8144,N_7568,N_7150);
nor U8145 (N_8145,N_7523,N_7852);
nor U8146 (N_8146,N_7040,N_7143);
nand U8147 (N_8147,N_7184,N_7316);
nor U8148 (N_8148,N_7477,N_7604);
nor U8149 (N_8149,N_7561,N_7051);
or U8150 (N_8150,N_7083,N_7174);
and U8151 (N_8151,N_7112,N_7610);
or U8152 (N_8152,N_7968,N_7197);
nand U8153 (N_8153,N_7903,N_7178);
nand U8154 (N_8154,N_7286,N_7206);
and U8155 (N_8155,N_7163,N_7091);
xor U8156 (N_8156,N_7823,N_7235);
and U8157 (N_8157,N_7292,N_7830);
nand U8158 (N_8158,N_7101,N_7977);
nand U8159 (N_8159,N_7800,N_7866);
nor U8160 (N_8160,N_7699,N_7265);
nand U8161 (N_8161,N_7654,N_7701);
or U8162 (N_8162,N_7547,N_7762);
nand U8163 (N_8163,N_7170,N_7243);
nor U8164 (N_8164,N_7173,N_7690);
and U8165 (N_8165,N_7141,N_7244);
or U8166 (N_8166,N_7248,N_7737);
or U8167 (N_8167,N_7719,N_7259);
nor U8168 (N_8168,N_7873,N_7931);
xor U8169 (N_8169,N_7939,N_7110);
or U8170 (N_8170,N_7423,N_7318);
and U8171 (N_8171,N_7757,N_7623);
nor U8172 (N_8172,N_7106,N_7994);
or U8173 (N_8173,N_7216,N_7457);
xnor U8174 (N_8174,N_7385,N_7297);
xor U8175 (N_8175,N_7207,N_7337);
or U8176 (N_8176,N_7503,N_7441);
and U8177 (N_8177,N_7395,N_7705);
nand U8178 (N_8178,N_7147,N_7435);
or U8179 (N_8179,N_7792,N_7111);
nor U8180 (N_8180,N_7187,N_7928);
nor U8181 (N_8181,N_7291,N_7857);
nor U8182 (N_8182,N_7774,N_7587);
nor U8183 (N_8183,N_7777,N_7253);
and U8184 (N_8184,N_7204,N_7258);
nor U8185 (N_8185,N_7416,N_7836);
nor U8186 (N_8186,N_7657,N_7584);
or U8187 (N_8187,N_7490,N_7842);
nand U8188 (N_8188,N_7449,N_7330);
and U8189 (N_8189,N_7636,N_7951);
nand U8190 (N_8190,N_7393,N_7431);
and U8191 (N_8191,N_7878,N_7388);
and U8192 (N_8192,N_7315,N_7084);
and U8193 (N_8193,N_7639,N_7946);
and U8194 (N_8194,N_7811,N_7914);
nor U8195 (N_8195,N_7061,N_7266);
xnor U8196 (N_8196,N_7653,N_7152);
nand U8197 (N_8197,N_7586,N_7962);
nand U8198 (N_8198,N_7967,N_7404);
xor U8199 (N_8199,N_7665,N_7381);
or U8200 (N_8200,N_7935,N_7990);
xnor U8201 (N_8201,N_7505,N_7066);
and U8202 (N_8202,N_7094,N_7474);
xnor U8203 (N_8203,N_7387,N_7934);
xor U8204 (N_8204,N_7014,N_7185);
and U8205 (N_8205,N_7254,N_7784);
xor U8206 (N_8206,N_7721,N_7376);
xor U8207 (N_8207,N_7473,N_7640);
nor U8208 (N_8208,N_7104,N_7400);
nand U8209 (N_8209,N_7979,N_7011);
xnor U8210 (N_8210,N_7965,N_7541);
nand U8211 (N_8211,N_7689,N_7392);
nor U8212 (N_8212,N_7427,N_7500);
nor U8213 (N_8213,N_7824,N_7600);
xnor U8214 (N_8214,N_7453,N_7563);
nor U8215 (N_8215,N_7950,N_7947);
and U8216 (N_8216,N_7789,N_7556);
or U8217 (N_8217,N_7507,N_7126);
nand U8218 (N_8218,N_7630,N_7841);
and U8219 (N_8219,N_7516,N_7420);
nand U8220 (N_8220,N_7537,N_7304);
or U8221 (N_8221,N_7532,N_7317);
nand U8222 (N_8222,N_7287,N_7323);
nand U8223 (N_8223,N_7548,N_7374);
and U8224 (N_8224,N_7578,N_7342);
nand U8225 (N_8225,N_7299,N_7284);
and U8226 (N_8226,N_7559,N_7002);
and U8227 (N_8227,N_7504,N_7881);
nor U8228 (N_8228,N_7334,N_7305);
nor U8229 (N_8229,N_7321,N_7213);
nand U8230 (N_8230,N_7897,N_7991);
xor U8231 (N_8231,N_7109,N_7188);
or U8232 (N_8232,N_7707,N_7158);
nand U8233 (N_8233,N_7851,N_7932);
and U8234 (N_8234,N_7551,N_7929);
and U8235 (N_8235,N_7585,N_7005);
nor U8236 (N_8236,N_7731,N_7691);
and U8237 (N_8237,N_7770,N_7133);
xor U8238 (N_8238,N_7217,N_7004);
and U8239 (N_8239,N_7879,N_7714);
xor U8240 (N_8240,N_7497,N_7612);
nand U8241 (N_8241,N_7849,N_7922);
and U8242 (N_8242,N_7620,N_7785);
or U8243 (N_8243,N_7535,N_7195);
and U8244 (N_8244,N_7569,N_7343);
or U8245 (N_8245,N_7558,N_7854);
and U8246 (N_8246,N_7632,N_7430);
nand U8247 (N_8247,N_7130,N_7176);
nor U8248 (N_8248,N_7773,N_7452);
or U8249 (N_8249,N_7606,N_7872);
nand U8250 (N_8250,N_7865,N_7646);
xnor U8251 (N_8251,N_7577,N_7264);
nor U8252 (N_8252,N_7858,N_7648);
and U8253 (N_8253,N_7467,N_7413);
nor U8254 (N_8254,N_7964,N_7643);
nand U8255 (N_8255,N_7927,N_7629);
xnor U8256 (N_8256,N_7885,N_7308);
nand U8257 (N_8257,N_7027,N_7534);
xnor U8258 (N_8258,N_7743,N_7877);
or U8259 (N_8259,N_7917,N_7182);
xnor U8260 (N_8260,N_7469,N_7786);
xnor U8261 (N_8261,N_7135,N_7941);
nand U8262 (N_8262,N_7201,N_7809);
or U8263 (N_8263,N_7999,N_7515);
xnor U8264 (N_8264,N_7703,N_7332);
or U8265 (N_8265,N_7686,N_7153);
and U8266 (N_8266,N_7675,N_7412);
nor U8267 (N_8267,N_7912,N_7687);
nand U8268 (N_8268,N_7202,N_7672);
or U8269 (N_8269,N_7390,N_7491);
nor U8270 (N_8270,N_7075,N_7289);
nand U8271 (N_8271,N_7742,N_7642);
or U8272 (N_8272,N_7512,N_7425);
nand U8273 (N_8273,N_7583,N_7871);
and U8274 (N_8274,N_7900,N_7099);
nand U8275 (N_8275,N_7383,N_7806);
xnor U8276 (N_8276,N_7989,N_7635);
and U8277 (N_8277,N_7615,N_7359);
and U8278 (N_8278,N_7476,N_7079);
and U8279 (N_8279,N_7300,N_7722);
nor U8280 (N_8280,N_7415,N_7295);
xor U8281 (N_8281,N_7916,N_7599);
nor U8282 (N_8282,N_7190,N_7930);
nor U8283 (N_8283,N_7760,N_7481);
nor U8284 (N_8284,N_7684,N_7862);
xnor U8285 (N_8285,N_7589,N_7692);
nand U8286 (N_8286,N_7124,N_7553);
or U8287 (N_8287,N_7171,N_7052);
xnor U8288 (N_8288,N_7886,N_7364);
xor U8289 (N_8289,N_7808,N_7593);
and U8290 (N_8290,N_7409,N_7882);
or U8291 (N_8291,N_7250,N_7456);
or U8292 (N_8292,N_7312,N_7611);
nor U8293 (N_8293,N_7509,N_7093);
nor U8294 (N_8294,N_7592,N_7436);
nor U8295 (N_8295,N_7156,N_7805);
nand U8296 (N_8296,N_7165,N_7987);
nor U8297 (N_8297,N_7498,N_7269);
and U8298 (N_8298,N_7290,N_7236);
and U8299 (N_8299,N_7831,N_7146);
nor U8300 (N_8300,N_7442,N_7087);
nand U8301 (N_8301,N_7241,N_7525);
and U8302 (N_8302,N_7725,N_7884);
and U8303 (N_8303,N_7550,N_7633);
xor U8304 (N_8304,N_7938,N_7097);
xnor U8305 (N_8305,N_7776,N_7239);
nand U8306 (N_8306,N_7370,N_7622);
nor U8307 (N_8307,N_7616,N_7552);
nor U8308 (N_8308,N_7398,N_7796);
and U8309 (N_8309,N_7983,N_7328);
xnor U8310 (N_8310,N_7234,N_7379);
or U8311 (N_8311,N_7918,N_7262);
nor U8312 (N_8312,N_7659,N_7298);
xnor U8313 (N_8313,N_7203,N_7679);
nor U8314 (N_8314,N_7761,N_7454);
and U8315 (N_8315,N_7985,N_7579);
nand U8316 (N_8316,N_7271,N_7003);
and U8317 (N_8317,N_7502,N_7050);
or U8318 (N_8318,N_7822,N_7267);
nand U8319 (N_8319,N_7191,N_7157);
and U8320 (N_8320,N_7437,N_7747);
nor U8321 (N_8321,N_7085,N_7352);
nand U8322 (N_8322,N_7647,N_7432);
nand U8323 (N_8323,N_7575,N_7017);
and U8324 (N_8324,N_7056,N_7440);
nand U8325 (N_8325,N_7160,N_7627);
or U8326 (N_8326,N_7309,N_7159);
nand U8327 (N_8327,N_7655,N_7086);
and U8328 (N_8328,N_7779,N_7026);
and U8329 (N_8329,N_7925,N_7088);
xnor U8330 (N_8330,N_7782,N_7006);
xor U8331 (N_8331,N_7369,N_7429);
nand U8332 (N_8332,N_7706,N_7702);
nand U8333 (N_8333,N_7015,N_7401);
nor U8334 (N_8334,N_7521,N_7478);
xnor U8335 (N_8335,N_7362,N_7817);
nor U8336 (N_8336,N_7716,N_7958);
xor U8337 (N_8337,N_7220,N_7033);
nor U8338 (N_8338,N_7720,N_7069);
nor U8339 (N_8339,N_7288,N_7624);
nand U8340 (N_8340,N_7952,N_7233);
nand U8341 (N_8341,N_7780,N_7314);
and U8342 (N_8342,N_7840,N_7710);
nor U8343 (N_8343,N_7843,N_7683);
nor U8344 (N_8344,N_7975,N_7329);
xor U8345 (N_8345,N_7389,N_7767);
nand U8346 (N_8346,N_7008,N_7384);
nand U8347 (N_8347,N_7260,N_7447);
and U8348 (N_8348,N_7230,N_7043);
and U8349 (N_8349,N_7740,N_7617);
xnor U8350 (N_8350,N_7926,N_7090);
nor U8351 (N_8351,N_7696,N_7268);
nand U8352 (N_8352,N_7038,N_7816);
nand U8353 (N_8353,N_7396,N_7905);
and U8354 (N_8354,N_7301,N_7222);
and U8355 (N_8355,N_7860,N_7000);
and U8356 (N_8356,N_7758,N_7164);
xor U8357 (N_8357,N_7861,N_7046);
xor U8358 (N_8358,N_7894,N_7828);
and U8359 (N_8359,N_7120,N_7915);
xor U8360 (N_8360,N_7517,N_7790);
xnor U8361 (N_8361,N_7718,N_7557);
nor U8362 (N_8362,N_7148,N_7489);
nor U8363 (N_8363,N_7293,N_7199);
nand U8364 (N_8364,N_7594,N_7492);
and U8365 (N_8365,N_7307,N_7913);
nor U8366 (N_8366,N_7765,N_7327);
and U8367 (N_8367,N_7494,N_7311);
xnor U8368 (N_8368,N_7783,N_7848);
and U8369 (N_8369,N_7107,N_7771);
nor U8370 (N_8370,N_7117,N_7669);
and U8371 (N_8371,N_7313,N_7715);
or U8372 (N_8372,N_7183,N_7285);
nand U8373 (N_8373,N_7054,N_7637);
or U8374 (N_8374,N_7460,N_7414);
nor U8375 (N_8375,N_7700,N_7208);
nor U8376 (N_8376,N_7528,N_7263);
nand U8377 (N_8377,N_7573,N_7402);
and U8378 (N_8378,N_7540,N_7766);
and U8379 (N_8379,N_7546,N_7281);
nand U8380 (N_8380,N_7196,N_7814);
or U8381 (N_8381,N_7123,N_7242);
nor U8382 (N_8382,N_7408,N_7741);
and U8383 (N_8383,N_7116,N_7793);
nand U8384 (N_8384,N_7487,N_7036);
or U8385 (N_8385,N_7403,N_7077);
and U8386 (N_8386,N_7803,N_7545);
nor U8387 (N_8387,N_7953,N_7121);
and U8388 (N_8388,N_7945,N_7065);
and U8389 (N_8389,N_7462,N_7007);
nor U8390 (N_8390,N_7868,N_7598);
and U8391 (N_8391,N_7936,N_7340);
or U8392 (N_8392,N_7542,N_7753);
or U8393 (N_8393,N_7544,N_7685);
or U8394 (N_8394,N_7246,N_7219);
or U8395 (N_8395,N_7856,N_7072);
and U8396 (N_8396,N_7883,N_7067);
nand U8397 (N_8397,N_7410,N_7969);
nand U8398 (N_8398,N_7798,N_7303);
and U8399 (N_8399,N_7671,N_7855);
or U8400 (N_8400,N_7446,N_7057);
xnor U8401 (N_8401,N_7209,N_7895);
nand U8402 (N_8402,N_7136,N_7645);
nor U8403 (N_8403,N_7055,N_7347);
and U8404 (N_8404,N_7499,N_7294);
or U8405 (N_8405,N_7122,N_7081);
nand U8406 (N_8406,N_7801,N_7907);
nor U8407 (N_8407,N_7826,N_7048);
nor U8408 (N_8408,N_7310,N_7735);
or U8409 (N_8409,N_7732,N_7649);
nor U8410 (N_8410,N_7277,N_7674);
nand U8411 (N_8411,N_7641,N_7025);
nand U8412 (N_8412,N_7272,N_7832);
nand U8413 (N_8413,N_7275,N_7030);
or U8414 (N_8414,N_7445,N_7944);
and U8415 (N_8415,N_7345,N_7354);
nor U8416 (N_8416,N_7465,N_7424);
and U8417 (N_8417,N_7175,N_7661);
nor U8418 (N_8418,N_7768,N_7167);
and U8419 (N_8419,N_7603,N_7211);
or U8420 (N_8420,N_7957,N_7333);
nand U8421 (N_8421,N_7475,N_7128);
nor U8422 (N_8422,N_7118,N_7533);
nand U8423 (N_8423,N_7638,N_7192);
or U8424 (N_8424,N_7829,N_7992);
and U8425 (N_8425,N_7458,N_7844);
and U8426 (N_8426,N_7363,N_7273);
or U8427 (N_8427,N_7549,N_7956);
nand U8428 (N_8428,N_7031,N_7910);
nor U8429 (N_8429,N_7697,N_7734);
xor U8430 (N_8430,N_7035,N_7775);
xnor U8431 (N_8431,N_7134,N_7668);
xor U8432 (N_8432,N_7261,N_7221);
or U8433 (N_8433,N_7518,N_7324);
and U8434 (N_8434,N_7045,N_7614);
and U8435 (N_8435,N_7787,N_7228);
nand U8436 (N_8436,N_7331,N_7891);
nand U8437 (N_8437,N_7911,N_7663);
nor U8438 (N_8438,N_7890,N_7496);
nor U8439 (N_8439,N_7954,N_7727);
nand U8440 (N_8440,N_7995,N_7626);
or U8441 (N_8441,N_7377,N_7682);
xor U8442 (N_8442,N_7839,N_7695);
and U8443 (N_8443,N_7506,N_7023);
xnor U8444 (N_8444,N_7988,N_7212);
or U8445 (N_8445,N_7405,N_7978);
xnor U8446 (N_8446,N_7588,N_7869);
xnor U8447 (N_8447,N_7812,N_7972);
xor U8448 (N_8448,N_7837,N_7438);
and U8449 (N_8449,N_7746,N_7673);
nand U8450 (N_8450,N_7892,N_7621);
or U8451 (N_8451,N_7513,N_7607);
and U8452 (N_8452,N_7717,N_7955);
nand U8453 (N_8453,N_7807,N_7893);
xor U8454 (N_8454,N_7322,N_7847);
and U8455 (N_8455,N_7631,N_7245);
nor U8456 (N_8456,N_7399,N_7224);
nand U8457 (N_8457,N_7943,N_7754);
and U8458 (N_8458,N_7670,N_7205);
nor U8459 (N_8459,N_7270,N_7016);
xor U8460 (N_8460,N_7524,N_7973);
xor U8461 (N_8461,N_7335,N_7778);
and U8462 (N_8462,N_7576,N_7769);
nor U8463 (N_8463,N_7919,N_7602);
and U8464 (N_8464,N_7596,N_7764);
and U8465 (N_8465,N_7063,N_7251);
xor U8466 (N_8466,N_7949,N_7834);
nand U8467 (N_8467,N_7450,N_7407);
xnor U8468 (N_8468,N_7073,N_7963);
nor U8469 (N_8469,N_7255,N_7451);
and U8470 (N_8470,N_7791,N_7468);
xnor U8471 (N_8471,N_7567,N_7417);
and U8472 (N_8472,N_7076,N_7933);
or U8473 (N_8473,N_7193,N_7326);
or U8474 (N_8474,N_7711,N_7756);
and U8475 (N_8475,N_7835,N_7406);
nor U8476 (N_8476,N_7514,N_7060);
nand U8477 (N_8477,N_7464,N_7887);
or U8478 (N_8478,N_7942,N_7283);
or U8479 (N_8479,N_7818,N_7472);
nor U8480 (N_8480,N_7020,N_7225);
nand U8481 (N_8481,N_7733,N_7426);
xnor U8482 (N_8482,N_7100,N_7821);
or U8483 (N_8483,N_7214,N_7982);
nand U8484 (N_8484,N_7252,N_7694);
and U8485 (N_8485,N_7920,N_7247);
or U8486 (N_8486,N_7256,N_7168);
or U8487 (N_8487,N_7194,N_7149);
or U8488 (N_8488,N_7797,N_7750);
xnor U8489 (N_8489,N_7378,N_7605);
xnor U8490 (N_8490,N_7029,N_7726);
xor U8491 (N_8491,N_7210,N_7341);
and U8492 (N_8492,N_7838,N_7339);
nand U8493 (N_8493,N_7581,N_7024);
nor U8494 (N_8494,N_7325,N_7948);
xor U8495 (N_8495,N_7418,N_7846);
nand U8496 (N_8496,N_7730,N_7781);
nor U8497 (N_8497,N_7365,N_7144);
or U8498 (N_8498,N_7053,N_7802);
nor U8499 (N_8499,N_7981,N_7704);
xnor U8500 (N_8500,N_7208,N_7827);
and U8501 (N_8501,N_7529,N_7149);
and U8502 (N_8502,N_7423,N_7352);
and U8503 (N_8503,N_7245,N_7096);
nand U8504 (N_8504,N_7072,N_7854);
and U8505 (N_8505,N_7330,N_7135);
nand U8506 (N_8506,N_7303,N_7999);
xor U8507 (N_8507,N_7588,N_7339);
or U8508 (N_8508,N_7347,N_7417);
or U8509 (N_8509,N_7471,N_7719);
nand U8510 (N_8510,N_7740,N_7215);
xor U8511 (N_8511,N_7557,N_7055);
or U8512 (N_8512,N_7337,N_7997);
nand U8513 (N_8513,N_7400,N_7995);
nor U8514 (N_8514,N_7417,N_7104);
nor U8515 (N_8515,N_7935,N_7937);
nand U8516 (N_8516,N_7982,N_7386);
xor U8517 (N_8517,N_7586,N_7377);
nor U8518 (N_8518,N_7363,N_7848);
nor U8519 (N_8519,N_7172,N_7143);
xor U8520 (N_8520,N_7513,N_7961);
xor U8521 (N_8521,N_7230,N_7638);
and U8522 (N_8522,N_7960,N_7962);
nor U8523 (N_8523,N_7326,N_7956);
nand U8524 (N_8524,N_7341,N_7441);
and U8525 (N_8525,N_7551,N_7698);
or U8526 (N_8526,N_7607,N_7234);
and U8527 (N_8527,N_7410,N_7098);
nor U8528 (N_8528,N_7722,N_7588);
and U8529 (N_8529,N_7416,N_7755);
and U8530 (N_8530,N_7302,N_7567);
nor U8531 (N_8531,N_7530,N_7356);
and U8532 (N_8532,N_7962,N_7774);
xor U8533 (N_8533,N_7567,N_7705);
xnor U8534 (N_8534,N_7763,N_7757);
nand U8535 (N_8535,N_7243,N_7357);
nand U8536 (N_8536,N_7983,N_7424);
and U8537 (N_8537,N_7608,N_7492);
xor U8538 (N_8538,N_7541,N_7752);
or U8539 (N_8539,N_7908,N_7961);
xor U8540 (N_8540,N_7426,N_7994);
nor U8541 (N_8541,N_7214,N_7656);
nand U8542 (N_8542,N_7618,N_7172);
xnor U8543 (N_8543,N_7358,N_7314);
or U8544 (N_8544,N_7243,N_7231);
and U8545 (N_8545,N_7537,N_7734);
or U8546 (N_8546,N_7032,N_7508);
nor U8547 (N_8547,N_7392,N_7653);
nor U8548 (N_8548,N_7903,N_7689);
or U8549 (N_8549,N_7172,N_7757);
and U8550 (N_8550,N_7066,N_7941);
nand U8551 (N_8551,N_7821,N_7700);
or U8552 (N_8552,N_7977,N_7261);
nor U8553 (N_8553,N_7542,N_7360);
nor U8554 (N_8554,N_7532,N_7841);
nor U8555 (N_8555,N_7151,N_7344);
or U8556 (N_8556,N_7809,N_7247);
xnor U8557 (N_8557,N_7975,N_7797);
and U8558 (N_8558,N_7970,N_7975);
xnor U8559 (N_8559,N_7939,N_7283);
nor U8560 (N_8560,N_7792,N_7121);
xnor U8561 (N_8561,N_7196,N_7976);
or U8562 (N_8562,N_7818,N_7066);
or U8563 (N_8563,N_7814,N_7838);
nand U8564 (N_8564,N_7067,N_7635);
nand U8565 (N_8565,N_7176,N_7521);
or U8566 (N_8566,N_7423,N_7381);
nand U8567 (N_8567,N_7712,N_7063);
xnor U8568 (N_8568,N_7157,N_7753);
xor U8569 (N_8569,N_7329,N_7134);
and U8570 (N_8570,N_7386,N_7199);
xor U8571 (N_8571,N_7422,N_7713);
xnor U8572 (N_8572,N_7603,N_7074);
xnor U8573 (N_8573,N_7888,N_7855);
nand U8574 (N_8574,N_7737,N_7813);
nor U8575 (N_8575,N_7193,N_7013);
or U8576 (N_8576,N_7938,N_7597);
xnor U8577 (N_8577,N_7421,N_7613);
and U8578 (N_8578,N_7689,N_7137);
and U8579 (N_8579,N_7843,N_7923);
or U8580 (N_8580,N_7893,N_7353);
xnor U8581 (N_8581,N_7722,N_7826);
nor U8582 (N_8582,N_7522,N_7414);
xor U8583 (N_8583,N_7456,N_7772);
or U8584 (N_8584,N_7676,N_7261);
xor U8585 (N_8585,N_7188,N_7683);
nand U8586 (N_8586,N_7477,N_7407);
or U8587 (N_8587,N_7378,N_7676);
or U8588 (N_8588,N_7897,N_7884);
xor U8589 (N_8589,N_7241,N_7966);
and U8590 (N_8590,N_7721,N_7237);
nor U8591 (N_8591,N_7421,N_7172);
nor U8592 (N_8592,N_7344,N_7895);
nor U8593 (N_8593,N_7271,N_7043);
and U8594 (N_8594,N_7334,N_7486);
xnor U8595 (N_8595,N_7716,N_7812);
or U8596 (N_8596,N_7819,N_7071);
or U8597 (N_8597,N_7575,N_7547);
nor U8598 (N_8598,N_7363,N_7764);
nor U8599 (N_8599,N_7032,N_7453);
xnor U8600 (N_8600,N_7212,N_7267);
xnor U8601 (N_8601,N_7804,N_7298);
xnor U8602 (N_8602,N_7631,N_7715);
nand U8603 (N_8603,N_7164,N_7937);
or U8604 (N_8604,N_7276,N_7880);
nand U8605 (N_8605,N_7821,N_7880);
nand U8606 (N_8606,N_7926,N_7011);
and U8607 (N_8607,N_7008,N_7064);
xnor U8608 (N_8608,N_7507,N_7566);
nand U8609 (N_8609,N_7034,N_7934);
nand U8610 (N_8610,N_7943,N_7532);
or U8611 (N_8611,N_7737,N_7905);
xnor U8612 (N_8612,N_7600,N_7861);
or U8613 (N_8613,N_7112,N_7503);
nand U8614 (N_8614,N_7742,N_7567);
and U8615 (N_8615,N_7170,N_7388);
nand U8616 (N_8616,N_7641,N_7818);
xnor U8617 (N_8617,N_7027,N_7226);
nand U8618 (N_8618,N_7783,N_7882);
nand U8619 (N_8619,N_7154,N_7671);
nor U8620 (N_8620,N_7580,N_7346);
nand U8621 (N_8621,N_7325,N_7612);
nor U8622 (N_8622,N_7333,N_7171);
nand U8623 (N_8623,N_7681,N_7998);
xnor U8624 (N_8624,N_7750,N_7393);
nand U8625 (N_8625,N_7571,N_7274);
nor U8626 (N_8626,N_7884,N_7774);
or U8627 (N_8627,N_7809,N_7994);
xnor U8628 (N_8628,N_7382,N_7774);
nor U8629 (N_8629,N_7879,N_7554);
or U8630 (N_8630,N_7410,N_7971);
nand U8631 (N_8631,N_7595,N_7541);
and U8632 (N_8632,N_7998,N_7478);
xnor U8633 (N_8633,N_7533,N_7177);
nor U8634 (N_8634,N_7021,N_7941);
nor U8635 (N_8635,N_7756,N_7020);
nor U8636 (N_8636,N_7601,N_7789);
xor U8637 (N_8637,N_7705,N_7324);
nor U8638 (N_8638,N_7023,N_7275);
nor U8639 (N_8639,N_7773,N_7682);
and U8640 (N_8640,N_7378,N_7285);
nor U8641 (N_8641,N_7636,N_7480);
and U8642 (N_8642,N_7959,N_7535);
nor U8643 (N_8643,N_7566,N_7883);
nand U8644 (N_8644,N_7609,N_7700);
or U8645 (N_8645,N_7073,N_7236);
nand U8646 (N_8646,N_7076,N_7485);
or U8647 (N_8647,N_7074,N_7194);
and U8648 (N_8648,N_7589,N_7388);
or U8649 (N_8649,N_7598,N_7846);
and U8650 (N_8650,N_7679,N_7396);
and U8651 (N_8651,N_7428,N_7153);
nand U8652 (N_8652,N_7299,N_7328);
xor U8653 (N_8653,N_7572,N_7374);
nor U8654 (N_8654,N_7487,N_7829);
xor U8655 (N_8655,N_7191,N_7844);
nand U8656 (N_8656,N_7230,N_7010);
or U8657 (N_8657,N_7177,N_7481);
nor U8658 (N_8658,N_7688,N_7880);
or U8659 (N_8659,N_7106,N_7224);
or U8660 (N_8660,N_7399,N_7392);
and U8661 (N_8661,N_7417,N_7915);
and U8662 (N_8662,N_7241,N_7612);
and U8663 (N_8663,N_7145,N_7004);
and U8664 (N_8664,N_7678,N_7855);
nor U8665 (N_8665,N_7072,N_7488);
xnor U8666 (N_8666,N_7543,N_7299);
nand U8667 (N_8667,N_7612,N_7979);
nand U8668 (N_8668,N_7224,N_7114);
or U8669 (N_8669,N_7387,N_7502);
nor U8670 (N_8670,N_7140,N_7432);
or U8671 (N_8671,N_7644,N_7873);
xor U8672 (N_8672,N_7406,N_7341);
nor U8673 (N_8673,N_7760,N_7004);
and U8674 (N_8674,N_7296,N_7066);
nand U8675 (N_8675,N_7510,N_7569);
xnor U8676 (N_8676,N_7417,N_7366);
nand U8677 (N_8677,N_7177,N_7100);
nor U8678 (N_8678,N_7864,N_7582);
or U8679 (N_8679,N_7755,N_7222);
xor U8680 (N_8680,N_7437,N_7027);
or U8681 (N_8681,N_7598,N_7363);
nor U8682 (N_8682,N_7214,N_7811);
or U8683 (N_8683,N_7815,N_7755);
nor U8684 (N_8684,N_7136,N_7186);
or U8685 (N_8685,N_7503,N_7460);
and U8686 (N_8686,N_7677,N_7765);
xnor U8687 (N_8687,N_7957,N_7058);
xnor U8688 (N_8688,N_7811,N_7036);
xnor U8689 (N_8689,N_7535,N_7997);
nand U8690 (N_8690,N_7670,N_7667);
nand U8691 (N_8691,N_7654,N_7035);
or U8692 (N_8692,N_7830,N_7305);
nand U8693 (N_8693,N_7256,N_7128);
and U8694 (N_8694,N_7689,N_7348);
and U8695 (N_8695,N_7665,N_7243);
or U8696 (N_8696,N_7654,N_7512);
nand U8697 (N_8697,N_7277,N_7271);
xnor U8698 (N_8698,N_7189,N_7546);
xor U8699 (N_8699,N_7025,N_7463);
nand U8700 (N_8700,N_7932,N_7198);
nand U8701 (N_8701,N_7511,N_7784);
or U8702 (N_8702,N_7646,N_7690);
xor U8703 (N_8703,N_7644,N_7754);
or U8704 (N_8704,N_7591,N_7347);
xor U8705 (N_8705,N_7272,N_7122);
or U8706 (N_8706,N_7561,N_7240);
xor U8707 (N_8707,N_7235,N_7629);
nand U8708 (N_8708,N_7347,N_7032);
nor U8709 (N_8709,N_7372,N_7926);
and U8710 (N_8710,N_7719,N_7409);
or U8711 (N_8711,N_7280,N_7945);
and U8712 (N_8712,N_7612,N_7305);
or U8713 (N_8713,N_7694,N_7666);
or U8714 (N_8714,N_7737,N_7706);
nand U8715 (N_8715,N_7224,N_7107);
xor U8716 (N_8716,N_7098,N_7187);
and U8717 (N_8717,N_7062,N_7075);
xnor U8718 (N_8718,N_7491,N_7534);
nand U8719 (N_8719,N_7690,N_7760);
and U8720 (N_8720,N_7488,N_7663);
or U8721 (N_8721,N_7704,N_7025);
nor U8722 (N_8722,N_7481,N_7635);
or U8723 (N_8723,N_7962,N_7204);
or U8724 (N_8724,N_7922,N_7712);
or U8725 (N_8725,N_7123,N_7545);
xnor U8726 (N_8726,N_7753,N_7287);
nor U8727 (N_8727,N_7722,N_7889);
xnor U8728 (N_8728,N_7787,N_7519);
and U8729 (N_8729,N_7307,N_7316);
or U8730 (N_8730,N_7558,N_7453);
or U8731 (N_8731,N_7014,N_7424);
and U8732 (N_8732,N_7158,N_7019);
or U8733 (N_8733,N_7480,N_7616);
nand U8734 (N_8734,N_7727,N_7689);
xor U8735 (N_8735,N_7779,N_7500);
xnor U8736 (N_8736,N_7847,N_7116);
nand U8737 (N_8737,N_7142,N_7196);
or U8738 (N_8738,N_7337,N_7846);
nand U8739 (N_8739,N_7050,N_7474);
xor U8740 (N_8740,N_7990,N_7925);
and U8741 (N_8741,N_7989,N_7055);
xnor U8742 (N_8742,N_7792,N_7604);
nor U8743 (N_8743,N_7903,N_7931);
xnor U8744 (N_8744,N_7277,N_7712);
nor U8745 (N_8745,N_7752,N_7679);
and U8746 (N_8746,N_7998,N_7830);
nand U8747 (N_8747,N_7293,N_7224);
nor U8748 (N_8748,N_7929,N_7417);
nand U8749 (N_8749,N_7352,N_7459);
and U8750 (N_8750,N_7632,N_7459);
and U8751 (N_8751,N_7167,N_7220);
xor U8752 (N_8752,N_7944,N_7898);
xor U8753 (N_8753,N_7966,N_7792);
or U8754 (N_8754,N_7706,N_7061);
nor U8755 (N_8755,N_7115,N_7410);
nor U8756 (N_8756,N_7627,N_7537);
and U8757 (N_8757,N_7654,N_7170);
xnor U8758 (N_8758,N_7321,N_7682);
xor U8759 (N_8759,N_7741,N_7183);
and U8760 (N_8760,N_7235,N_7067);
nand U8761 (N_8761,N_7968,N_7650);
or U8762 (N_8762,N_7401,N_7379);
and U8763 (N_8763,N_7690,N_7424);
nand U8764 (N_8764,N_7028,N_7116);
or U8765 (N_8765,N_7642,N_7752);
xnor U8766 (N_8766,N_7405,N_7326);
nand U8767 (N_8767,N_7667,N_7335);
nor U8768 (N_8768,N_7011,N_7895);
and U8769 (N_8769,N_7930,N_7455);
nor U8770 (N_8770,N_7045,N_7864);
xnor U8771 (N_8771,N_7923,N_7816);
xor U8772 (N_8772,N_7984,N_7917);
nand U8773 (N_8773,N_7296,N_7054);
and U8774 (N_8774,N_7958,N_7049);
and U8775 (N_8775,N_7351,N_7483);
nand U8776 (N_8776,N_7242,N_7010);
or U8777 (N_8777,N_7790,N_7959);
nor U8778 (N_8778,N_7532,N_7879);
nor U8779 (N_8779,N_7101,N_7765);
and U8780 (N_8780,N_7628,N_7187);
and U8781 (N_8781,N_7594,N_7165);
and U8782 (N_8782,N_7473,N_7297);
or U8783 (N_8783,N_7264,N_7211);
nand U8784 (N_8784,N_7985,N_7695);
and U8785 (N_8785,N_7230,N_7020);
nor U8786 (N_8786,N_7947,N_7119);
nor U8787 (N_8787,N_7019,N_7696);
nand U8788 (N_8788,N_7647,N_7756);
nor U8789 (N_8789,N_7581,N_7492);
nor U8790 (N_8790,N_7317,N_7717);
and U8791 (N_8791,N_7097,N_7664);
or U8792 (N_8792,N_7892,N_7218);
nor U8793 (N_8793,N_7896,N_7791);
or U8794 (N_8794,N_7753,N_7875);
nand U8795 (N_8795,N_7047,N_7737);
nand U8796 (N_8796,N_7365,N_7989);
nand U8797 (N_8797,N_7895,N_7833);
or U8798 (N_8798,N_7497,N_7043);
nor U8799 (N_8799,N_7165,N_7844);
nand U8800 (N_8800,N_7384,N_7338);
nand U8801 (N_8801,N_7849,N_7845);
nand U8802 (N_8802,N_7349,N_7076);
nand U8803 (N_8803,N_7022,N_7004);
and U8804 (N_8804,N_7414,N_7060);
nand U8805 (N_8805,N_7111,N_7541);
and U8806 (N_8806,N_7965,N_7868);
nor U8807 (N_8807,N_7806,N_7504);
nor U8808 (N_8808,N_7837,N_7282);
or U8809 (N_8809,N_7343,N_7495);
and U8810 (N_8810,N_7410,N_7647);
or U8811 (N_8811,N_7023,N_7723);
nor U8812 (N_8812,N_7369,N_7941);
nor U8813 (N_8813,N_7473,N_7116);
or U8814 (N_8814,N_7793,N_7662);
nand U8815 (N_8815,N_7588,N_7656);
and U8816 (N_8816,N_7315,N_7956);
or U8817 (N_8817,N_7226,N_7511);
nand U8818 (N_8818,N_7418,N_7023);
or U8819 (N_8819,N_7130,N_7110);
or U8820 (N_8820,N_7820,N_7327);
xor U8821 (N_8821,N_7714,N_7648);
xnor U8822 (N_8822,N_7143,N_7983);
nor U8823 (N_8823,N_7935,N_7773);
xor U8824 (N_8824,N_7503,N_7752);
xor U8825 (N_8825,N_7282,N_7071);
xnor U8826 (N_8826,N_7053,N_7508);
or U8827 (N_8827,N_7139,N_7291);
nor U8828 (N_8828,N_7861,N_7386);
and U8829 (N_8829,N_7344,N_7101);
and U8830 (N_8830,N_7968,N_7640);
nor U8831 (N_8831,N_7380,N_7159);
xor U8832 (N_8832,N_7974,N_7288);
nand U8833 (N_8833,N_7411,N_7850);
or U8834 (N_8834,N_7590,N_7509);
nand U8835 (N_8835,N_7018,N_7488);
xnor U8836 (N_8836,N_7530,N_7967);
nand U8837 (N_8837,N_7231,N_7816);
nand U8838 (N_8838,N_7478,N_7968);
and U8839 (N_8839,N_7716,N_7756);
nor U8840 (N_8840,N_7355,N_7676);
and U8841 (N_8841,N_7493,N_7017);
xor U8842 (N_8842,N_7768,N_7635);
or U8843 (N_8843,N_7482,N_7009);
xor U8844 (N_8844,N_7031,N_7628);
and U8845 (N_8845,N_7794,N_7503);
xor U8846 (N_8846,N_7563,N_7628);
and U8847 (N_8847,N_7695,N_7047);
and U8848 (N_8848,N_7929,N_7384);
or U8849 (N_8849,N_7026,N_7069);
xnor U8850 (N_8850,N_7599,N_7095);
nand U8851 (N_8851,N_7582,N_7877);
nor U8852 (N_8852,N_7372,N_7124);
xor U8853 (N_8853,N_7150,N_7043);
and U8854 (N_8854,N_7775,N_7428);
xnor U8855 (N_8855,N_7638,N_7145);
xor U8856 (N_8856,N_7969,N_7452);
or U8857 (N_8857,N_7933,N_7728);
nor U8858 (N_8858,N_7658,N_7800);
or U8859 (N_8859,N_7450,N_7060);
nor U8860 (N_8860,N_7319,N_7731);
xnor U8861 (N_8861,N_7136,N_7540);
xnor U8862 (N_8862,N_7696,N_7417);
or U8863 (N_8863,N_7764,N_7849);
and U8864 (N_8864,N_7529,N_7924);
nor U8865 (N_8865,N_7238,N_7878);
and U8866 (N_8866,N_7347,N_7577);
nor U8867 (N_8867,N_7148,N_7433);
and U8868 (N_8868,N_7305,N_7762);
or U8869 (N_8869,N_7720,N_7561);
or U8870 (N_8870,N_7532,N_7422);
nor U8871 (N_8871,N_7298,N_7028);
nor U8872 (N_8872,N_7979,N_7351);
and U8873 (N_8873,N_7439,N_7568);
xor U8874 (N_8874,N_7279,N_7032);
nand U8875 (N_8875,N_7283,N_7093);
xnor U8876 (N_8876,N_7762,N_7137);
and U8877 (N_8877,N_7446,N_7080);
xor U8878 (N_8878,N_7545,N_7070);
nand U8879 (N_8879,N_7092,N_7422);
nor U8880 (N_8880,N_7684,N_7763);
xor U8881 (N_8881,N_7776,N_7398);
nor U8882 (N_8882,N_7555,N_7953);
and U8883 (N_8883,N_7636,N_7497);
xnor U8884 (N_8884,N_7168,N_7274);
xnor U8885 (N_8885,N_7743,N_7031);
or U8886 (N_8886,N_7273,N_7629);
and U8887 (N_8887,N_7322,N_7200);
nand U8888 (N_8888,N_7199,N_7758);
or U8889 (N_8889,N_7700,N_7603);
or U8890 (N_8890,N_7358,N_7260);
and U8891 (N_8891,N_7797,N_7399);
xor U8892 (N_8892,N_7825,N_7649);
xor U8893 (N_8893,N_7104,N_7529);
nor U8894 (N_8894,N_7350,N_7980);
nor U8895 (N_8895,N_7348,N_7603);
and U8896 (N_8896,N_7579,N_7871);
and U8897 (N_8897,N_7132,N_7351);
or U8898 (N_8898,N_7094,N_7329);
xnor U8899 (N_8899,N_7056,N_7817);
nand U8900 (N_8900,N_7363,N_7916);
xor U8901 (N_8901,N_7244,N_7025);
and U8902 (N_8902,N_7030,N_7053);
xnor U8903 (N_8903,N_7890,N_7187);
nand U8904 (N_8904,N_7792,N_7545);
or U8905 (N_8905,N_7573,N_7609);
xnor U8906 (N_8906,N_7918,N_7555);
nand U8907 (N_8907,N_7953,N_7557);
xor U8908 (N_8908,N_7384,N_7480);
xnor U8909 (N_8909,N_7444,N_7252);
or U8910 (N_8910,N_7525,N_7700);
xnor U8911 (N_8911,N_7200,N_7744);
nand U8912 (N_8912,N_7951,N_7884);
and U8913 (N_8913,N_7701,N_7712);
xnor U8914 (N_8914,N_7223,N_7885);
xor U8915 (N_8915,N_7140,N_7254);
and U8916 (N_8916,N_7406,N_7876);
nand U8917 (N_8917,N_7118,N_7321);
or U8918 (N_8918,N_7957,N_7195);
and U8919 (N_8919,N_7438,N_7843);
xor U8920 (N_8920,N_7242,N_7760);
or U8921 (N_8921,N_7141,N_7763);
nand U8922 (N_8922,N_7241,N_7214);
xor U8923 (N_8923,N_7151,N_7188);
nor U8924 (N_8924,N_7093,N_7775);
nor U8925 (N_8925,N_7299,N_7811);
and U8926 (N_8926,N_7153,N_7168);
or U8927 (N_8927,N_7820,N_7719);
and U8928 (N_8928,N_7696,N_7735);
nand U8929 (N_8929,N_7231,N_7762);
nor U8930 (N_8930,N_7218,N_7491);
nor U8931 (N_8931,N_7612,N_7834);
nor U8932 (N_8932,N_7035,N_7350);
nand U8933 (N_8933,N_7250,N_7817);
and U8934 (N_8934,N_7915,N_7849);
nand U8935 (N_8935,N_7727,N_7893);
nor U8936 (N_8936,N_7762,N_7785);
nand U8937 (N_8937,N_7009,N_7152);
and U8938 (N_8938,N_7897,N_7043);
xor U8939 (N_8939,N_7346,N_7225);
xor U8940 (N_8940,N_7473,N_7639);
xnor U8941 (N_8941,N_7996,N_7608);
or U8942 (N_8942,N_7039,N_7855);
or U8943 (N_8943,N_7937,N_7529);
and U8944 (N_8944,N_7490,N_7721);
nor U8945 (N_8945,N_7424,N_7488);
and U8946 (N_8946,N_7152,N_7357);
nor U8947 (N_8947,N_7007,N_7169);
or U8948 (N_8948,N_7545,N_7798);
xnor U8949 (N_8949,N_7216,N_7065);
nor U8950 (N_8950,N_7800,N_7055);
xnor U8951 (N_8951,N_7343,N_7137);
nand U8952 (N_8952,N_7781,N_7387);
or U8953 (N_8953,N_7493,N_7114);
nor U8954 (N_8954,N_7301,N_7556);
nor U8955 (N_8955,N_7073,N_7522);
and U8956 (N_8956,N_7732,N_7583);
nor U8957 (N_8957,N_7599,N_7834);
xnor U8958 (N_8958,N_7031,N_7625);
nor U8959 (N_8959,N_7348,N_7043);
nor U8960 (N_8960,N_7451,N_7693);
xor U8961 (N_8961,N_7074,N_7079);
nor U8962 (N_8962,N_7541,N_7579);
or U8963 (N_8963,N_7742,N_7578);
or U8964 (N_8964,N_7396,N_7074);
nor U8965 (N_8965,N_7961,N_7116);
and U8966 (N_8966,N_7826,N_7755);
nor U8967 (N_8967,N_7796,N_7652);
nand U8968 (N_8968,N_7389,N_7124);
or U8969 (N_8969,N_7385,N_7674);
nand U8970 (N_8970,N_7963,N_7326);
and U8971 (N_8971,N_7959,N_7834);
and U8972 (N_8972,N_7508,N_7921);
and U8973 (N_8973,N_7912,N_7351);
and U8974 (N_8974,N_7099,N_7472);
or U8975 (N_8975,N_7775,N_7132);
xnor U8976 (N_8976,N_7853,N_7028);
nor U8977 (N_8977,N_7840,N_7846);
nand U8978 (N_8978,N_7642,N_7071);
and U8979 (N_8979,N_7387,N_7909);
and U8980 (N_8980,N_7004,N_7675);
xor U8981 (N_8981,N_7474,N_7802);
and U8982 (N_8982,N_7185,N_7702);
and U8983 (N_8983,N_7740,N_7521);
or U8984 (N_8984,N_7399,N_7488);
xor U8985 (N_8985,N_7716,N_7455);
xnor U8986 (N_8986,N_7951,N_7245);
or U8987 (N_8987,N_7274,N_7984);
and U8988 (N_8988,N_7601,N_7101);
or U8989 (N_8989,N_7410,N_7640);
nor U8990 (N_8990,N_7943,N_7121);
nand U8991 (N_8991,N_7646,N_7479);
nand U8992 (N_8992,N_7291,N_7030);
and U8993 (N_8993,N_7557,N_7176);
nor U8994 (N_8994,N_7708,N_7374);
and U8995 (N_8995,N_7901,N_7020);
xor U8996 (N_8996,N_7875,N_7533);
and U8997 (N_8997,N_7001,N_7375);
nor U8998 (N_8998,N_7236,N_7043);
and U8999 (N_8999,N_7229,N_7795);
nand U9000 (N_9000,N_8800,N_8756);
nor U9001 (N_9001,N_8382,N_8921);
and U9002 (N_9002,N_8551,N_8373);
or U9003 (N_9003,N_8839,N_8063);
xnor U9004 (N_9004,N_8436,N_8245);
and U9005 (N_9005,N_8579,N_8202);
nor U9006 (N_9006,N_8682,N_8770);
or U9007 (N_9007,N_8392,N_8652);
nand U9008 (N_9008,N_8901,N_8528);
and U9009 (N_9009,N_8697,N_8851);
nor U9010 (N_9010,N_8386,N_8473);
and U9011 (N_9011,N_8044,N_8902);
or U9012 (N_9012,N_8308,N_8025);
and U9013 (N_9013,N_8254,N_8206);
xnor U9014 (N_9014,N_8628,N_8763);
xnor U9015 (N_9015,N_8422,N_8434);
nand U9016 (N_9016,N_8844,N_8925);
nand U9017 (N_9017,N_8592,N_8097);
nor U9018 (N_9018,N_8356,N_8663);
nand U9019 (N_9019,N_8446,N_8014);
xnor U9020 (N_9020,N_8140,N_8156);
nor U9021 (N_9021,N_8300,N_8781);
or U9022 (N_9022,N_8240,N_8562);
xnor U9023 (N_9023,N_8113,N_8067);
nor U9024 (N_9024,N_8909,N_8270);
xor U9025 (N_9025,N_8758,N_8132);
or U9026 (N_9026,N_8601,N_8124);
and U9027 (N_9027,N_8748,N_8737);
and U9028 (N_9028,N_8584,N_8893);
and U9029 (N_9029,N_8280,N_8725);
nor U9030 (N_9030,N_8217,N_8913);
nor U9031 (N_9031,N_8058,N_8732);
nor U9032 (N_9032,N_8459,N_8670);
nor U9033 (N_9033,N_8543,N_8537);
nand U9034 (N_9034,N_8546,N_8509);
nand U9035 (N_9035,N_8218,N_8702);
or U9036 (N_9036,N_8004,N_8147);
nand U9037 (N_9037,N_8785,N_8742);
or U9038 (N_9038,N_8615,N_8089);
nand U9039 (N_9039,N_8503,N_8019);
nand U9040 (N_9040,N_8419,N_8167);
and U9041 (N_9041,N_8624,N_8250);
or U9042 (N_9042,N_8786,N_8148);
or U9043 (N_9043,N_8618,N_8507);
xor U9044 (N_9044,N_8887,N_8407);
nor U9045 (N_9045,N_8357,N_8984);
or U9046 (N_9046,N_8056,N_8621);
or U9047 (N_9047,N_8006,N_8052);
xor U9048 (N_9048,N_8332,N_8049);
nor U9049 (N_9049,N_8677,N_8573);
nand U9050 (N_9050,N_8387,N_8418);
nor U9051 (N_9051,N_8325,N_8606);
xor U9052 (N_9052,N_8944,N_8164);
xnor U9053 (N_9053,N_8121,N_8403);
or U9054 (N_9054,N_8144,N_8223);
nand U9055 (N_9055,N_8169,N_8687);
nand U9056 (N_9056,N_8723,N_8029);
nand U9057 (N_9057,N_8972,N_8066);
nand U9058 (N_9058,N_8421,N_8349);
xor U9059 (N_9059,N_8484,N_8559);
nor U9060 (N_9060,N_8865,N_8142);
nor U9061 (N_9061,N_8681,N_8203);
xor U9062 (N_9062,N_8690,N_8461);
and U9063 (N_9063,N_8774,N_8924);
xnor U9064 (N_9064,N_8940,N_8072);
nand U9065 (N_9065,N_8453,N_8700);
nor U9066 (N_9066,N_8005,N_8840);
nand U9067 (N_9067,N_8733,N_8252);
and U9068 (N_9068,N_8717,N_8751);
xor U9069 (N_9069,N_8975,N_8731);
or U9070 (N_9070,N_8087,N_8661);
or U9071 (N_9071,N_8582,N_8249);
xor U9072 (N_9072,N_8784,N_8013);
or U9073 (N_9073,N_8627,N_8266);
nand U9074 (N_9074,N_8205,N_8879);
nand U9075 (N_9075,N_8374,N_8655);
and U9076 (N_9076,N_8305,N_8965);
nor U9077 (N_9077,N_8511,N_8799);
or U9078 (N_9078,N_8368,N_8157);
nand U9079 (N_9079,N_8499,N_8881);
and U9080 (N_9080,N_8900,N_8173);
nand U9081 (N_9081,N_8111,N_8302);
and U9082 (N_9082,N_8523,N_8318);
nor U9083 (N_9083,N_8754,N_8316);
or U9084 (N_9084,N_8378,N_8815);
nor U9085 (N_9085,N_8420,N_8221);
xor U9086 (N_9086,N_8172,N_8787);
and U9087 (N_9087,N_8504,N_8480);
and U9088 (N_9088,N_8607,N_8662);
nand U9089 (N_9089,N_8194,N_8365);
or U9090 (N_9090,N_8567,N_8450);
nor U9091 (N_9091,N_8323,N_8908);
xor U9092 (N_9092,N_8428,N_8439);
and U9093 (N_9093,N_8744,N_8103);
or U9094 (N_9094,N_8435,N_8855);
xnor U9095 (N_9095,N_8059,N_8791);
and U9096 (N_9096,N_8296,N_8307);
or U9097 (N_9097,N_8824,N_8856);
and U9098 (N_9098,N_8634,N_8050);
nand U9099 (N_9099,N_8686,N_8916);
or U9100 (N_9100,N_8466,N_8168);
and U9101 (N_9101,N_8035,N_8017);
nor U9102 (N_9102,N_8427,N_8312);
xnor U9103 (N_9103,N_8967,N_8570);
xor U9104 (N_9104,N_8135,N_8971);
nand U9105 (N_9105,N_8355,N_8021);
nand U9106 (N_9106,N_8952,N_8083);
nand U9107 (N_9107,N_8423,N_8798);
nand U9108 (N_9108,N_8888,N_8572);
nor U9109 (N_9109,N_8076,N_8379);
and U9110 (N_9110,N_8062,N_8350);
xor U9111 (N_9111,N_8348,N_8891);
or U9112 (N_9112,N_8271,N_8342);
nor U9113 (N_9113,N_8729,N_8396);
or U9114 (N_9114,N_8992,N_8811);
xor U9115 (N_9115,N_8789,N_8264);
or U9116 (N_9116,N_8657,N_8228);
and U9117 (N_9117,N_8796,N_8255);
nand U9118 (N_9118,N_8073,N_8701);
and U9119 (N_9119,N_8912,N_8694);
nor U9120 (N_9120,N_8776,N_8287);
nor U9121 (N_9121,N_8110,N_8558);
nand U9122 (N_9122,N_8877,N_8120);
or U9123 (N_9123,N_8740,N_8492);
xor U9124 (N_9124,N_8755,N_8177);
nor U9125 (N_9125,N_8531,N_8874);
nor U9126 (N_9126,N_8125,N_8198);
nand U9127 (N_9127,N_8917,N_8163);
or U9128 (N_9128,N_8415,N_8096);
or U9129 (N_9129,N_8208,N_8922);
xor U9130 (N_9130,N_8061,N_8759);
or U9131 (N_9131,N_8892,N_8850);
xnor U9132 (N_9132,N_8611,N_8640);
and U9133 (N_9133,N_8158,N_8105);
nand U9134 (N_9134,N_8878,N_8767);
nand U9135 (N_9135,N_8768,N_8806);
and U9136 (N_9136,N_8919,N_8589);
and U9137 (N_9137,N_8054,N_8793);
or U9138 (N_9138,N_8540,N_8956);
nand U9139 (N_9139,N_8460,N_8950);
nand U9140 (N_9140,N_8630,N_8539);
nand U9141 (N_9141,N_8053,N_8290);
and U9142 (N_9142,N_8042,N_8506);
nand U9143 (N_9143,N_8283,N_8684);
or U9144 (N_9144,N_8286,N_8894);
or U9145 (N_9145,N_8711,N_8243);
nand U9146 (N_9146,N_8846,N_8020);
or U9147 (N_9147,N_8384,N_8358);
and U9148 (N_9148,N_8612,N_8366);
nand U9149 (N_9149,N_8788,N_8849);
xor U9150 (N_9150,N_8822,N_8672);
or U9151 (N_9151,N_8968,N_8735);
nand U9152 (N_9152,N_8211,N_8385);
or U9153 (N_9153,N_8244,N_8039);
xor U9154 (N_9154,N_8556,N_8333);
or U9155 (N_9155,N_8997,N_8225);
nand U9156 (N_9156,N_8406,N_8669);
nand U9157 (N_9157,N_8159,N_8993);
nor U9158 (N_9158,N_8576,N_8795);
or U9159 (N_9159,N_8638,N_8226);
nand U9160 (N_9160,N_8186,N_8613);
xor U9161 (N_9161,N_8081,N_8995);
nor U9162 (N_9162,N_8519,N_8693);
and U9163 (N_9163,N_8635,N_8279);
nand U9164 (N_9164,N_8691,N_8027);
nand U9165 (N_9165,N_8478,N_8360);
nor U9166 (N_9166,N_8721,N_8747);
nor U9167 (N_9167,N_8571,N_8903);
xnor U9168 (N_9168,N_8516,N_8870);
nand U9169 (N_9169,N_8602,N_8381);
and U9170 (N_9170,N_8297,N_8346);
nand U9171 (N_9171,N_8497,N_8857);
nor U9172 (N_9172,N_8549,N_8141);
and U9173 (N_9173,N_8835,N_8698);
nand U9174 (N_9174,N_8896,N_8311);
nand U9175 (N_9175,N_8015,N_8914);
nand U9176 (N_9176,N_8003,N_8170);
nor U9177 (N_9177,N_8032,N_8685);
or U9178 (N_9178,N_8468,N_8915);
and U9179 (N_9179,N_8676,N_8253);
xor U9180 (N_9180,N_8837,N_8843);
nand U9181 (N_9181,N_8077,N_8367);
and U9182 (N_9182,N_8750,N_8265);
nor U9183 (N_9183,N_8958,N_8749);
or U9184 (N_9184,N_8500,N_8114);
xnor U9185 (N_9185,N_8372,N_8183);
and U9186 (N_9186,N_8472,N_8433);
nand U9187 (N_9187,N_8778,N_8364);
nand U9188 (N_9188,N_8370,N_8109);
or U9189 (N_9189,N_8819,N_8889);
nand U9190 (N_9190,N_8040,N_8345);
and U9191 (N_9191,N_8552,N_8561);
xor U9192 (N_9192,N_8301,N_8743);
nand U9193 (N_9193,N_8859,N_8978);
nand U9194 (N_9194,N_8309,N_8091);
xnor U9195 (N_9195,N_8152,N_8505);
xor U9196 (N_9196,N_8398,N_8961);
nor U9197 (N_9197,N_8586,N_8236);
xor U9198 (N_9198,N_8939,N_8585);
nor U9199 (N_9199,N_8610,N_8619);
or U9200 (N_9200,N_8658,N_8022);
or U9201 (N_9201,N_8028,N_8327);
nor U9202 (N_9202,N_8873,N_8391);
xnor U9203 (N_9203,N_8649,N_8547);
nor U9204 (N_9204,N_8119,N_8990);
nand U9205 (N_9205,N_8578,N_8727);
nand U9206 (N_9206,N_8529,N_8193);
nand U9207 (N_9207,N_8431,N_8128);
nand U9208 (N_9208,N_8769,N_8777);
xor U9209 (N_9209,N_8942,N_8339);
nor U9210 (N_9210,N_8425,N_8895);
xor U9211 (N_9211,N_8192,N_8093);
and U9212 (N_9212,N_8477,N_8046);
or U9213 (N_9213,N_8078,N_8175);
xnor U9214 (N_9214,N_8234,N_8617);
nand U9215 (N_9215,N_8149,N_8263);
nor U9216 (N_9216,N_8320,N_8598);
nand U9217 (N_9217,N_8051,N_8179);
or U9218 (N_9218,N_8771,N_8359);
nor U9219 (N_9219,N_8581,N_8550);
and U9220 (N_9220,N_8825,N_8591);
and U9221 (N_9221,N_8739,N_8836);
and U9222 (N_9222,N_8007,N_8935);
nor U9223 (N_9223,N_8294,N_8008);
nor U9224 (N_9224,N_8165,N_8444);
or U9225 (N_9225,N_8470,N_8475);
or U9226 (N_9226,N_8564,N_8184);
nor U9227 (N_9227,N_8577,N_8931);
xnor U9228 (N_9228,N_8282,N_8488);
nor U9229 (N_9229,N_8970,N_8981);
xnor U9230 (N_9230,N_8929,N_8651);
nand U9231 (N_9231,N_8195,N_8298);
nand U9232 (N_9232,N_8980,N_8115);
xor U9233 (N_9233,N_8947,N_8112);
and U9234 (N_9234,N_8928,N_8314);
or U9235 (N_9235,N_8988,N_8371);
nor U9236 (N_9236,N_8313,N_8196);
nand U9237 (N_9237,N_8842,N_8490);
nand U9238 (N_9238,N_8375,N_8092);
or U9239 (N_9239,N_8389,N_8829);
nand U9240 (N_9240,N_8304,N_8764);
and U9241 (N_9241,N_8369,N_8853);
nor U9242 (N_9242,N_8449,N_8716);
nor U9243 (N_9243,N_8963,N_8641);
nor U9244 (N_9244,N_8522,N_8817);
and U9245 (N_9245,N_8395,N_8945);
xor U9246 (N_9246,N_8934,N_8251);
xor U9247 (N_9247,N_8229,N_8991);
nand U9248 (N_9248,N_8455,N_8650);
nand U9249 (N_9249,N_8321,N_8803);
xnor U9250 (N_9250,N_8692,N_8329);
nor U9251 (N_9251,N_8084,N_8966);
or U9252 (N_9252,N_8773,N_8487);
nand U9253 (N_9253,N_8154,N_8224);
nand U9254 (N_9254,N_8603,N_8680);
nand U9255 (N_9255,N_8043,N_8653);
xor U9256 (N_9256,N_8994,N_8190);
nor U9257 (N_9257,N_8214,N_8599);
and U9258 (N_9258,N_8639,N_8979);
or U9259 (N_9259,N_8131,N_8590);
nand U9260 (N_9260,N_8261,N_8838);
xnor U9261 (N_9261,N_8937,N_8098);
nor U9262 (N_9262,N_8536,N_8476);
nand U9263 (N_9263,N_8237,N_8133);
nand U9264 (N_9264,N_8269,N_8210);
and U9265 (N_9265,N_8812,N_8608);
and U9266 (N_9266,N_8334,N_8841);
nor U9267 (N_9267,N_8495,N_8456);
nand U9268 (N_9268,N_8647,N_8510);
and U9269 (N_9269,N_8719,N_8447);
and U9270 (N_9270,N_8104,N_8792);
or U9271 (N_9271,N_8703,N_8180);
nand U9272 (N_9272,N_8143,N_8426);
nand U9273 (N_9273,N_8411,N_8090);
xor U9274 (N_9274,N_8974,N_8408);
or U9275 (N_9275,N_8996,N_8730);
nand U9276 (N_9276,N_8918,N_8959);
xor U9277 (N_9277,N_8710,N_8766);
nand U9278 (N_9278,N_8910,N_8593);
nand U9279 (N_9279,N_8830,N_8762);
nand U9280 (N_9280,N_8099,N_8782);
or U9281 (N_9281,N_8757,N_8438);
and U9282 (N_9282,N_8813,N_8233);
xnor U9283 (N_9283,N_8187,N_8609);
or U9284 (N_9284,N_8055,N_8752);
and U9285 (N_9285,N_8064,N_8033);
nor U9286 (N_9286,N_8377,N_8380);
nand U9287 (N_9287,N_8828,N_8361);
or U9288 (N_9288,N_8779,N_8563);
and U9289 (N_9289,N_8905,N_8048);
nor U9290 (N_9290,N_8134,N_8343);
nor U9291 (N_9291,N_8341,N_8845);
xor U9292 (N_9292,N_8741,N_8262);
nand U9293 (N_9293,N_8363,N_8906);
xnor U9294 (N_9294,N_8648,N_8679);
nand U9295 (N_9295,N_8864,N_8498);
xnor U9296 (N_9296,N_8715,N_8285);
nor U9297 (N_9297,N_8069,N_8409);
and U9298 (N_9298,N_8106,N_8854);
nand U9299 (N_9299,N_8102,N_8258);
or U9300 (N_9300,N_8277,N_8580);
nand U9301 (N_9301,N_8868,N_8821);
and U9302 (N_9302,N_8432,N_8955);
or U9303 (N_9303,N_8883,N_8319);
nand U9304 (N_9304,N_8116,N_8000);
xnor U9305 (N_9305,N_8181,N_8726);
or U9306 (N_9306,N_8414,N_8976);
xor U9307 (N_9307,N_8724,N_8930);
xor U9308 (N_9308,N_8852,N_8867);
xnor U9309 (N_9309,N_8594,N_8161);
or U9310 (N_9310,N_8448,N_8036);
or U9311 (N_9311,N_8220,N_8969);
nor U9312 (N_9312,N_8568,N_8616);
nor U9313 (N_9313,N_8885,N_8954);
and U9314 (N_9314,N_8001,N_8412);
xor U9315 (N_9315,N_8441,N_8464);
nor U9316 (N_9316,N_8227,N_8898);
nor U9317 (N_9317,N_8642,N_8532);
xnor U9318 (N_9318,N_8646,N_8151);
xnor U9319 (N_9319,N_8794,N_8026);
and U9320 (N_9320,N_8704,N_8807);
xor U9321 (N_9321,N_8554,N_8278);
nand U9322 (N_9322,N_8065,N_8204);
nor U9323 (N_9323,N_8437,N_8016);
xor U9324 (N_9324,N_8080,N_8197);
and U9325 (N_9325,N_8595,N_8268);
and U9326 (N_9326,N_8805,N_8376);
and U9327 (N_9327,N_8513,N_8284);
nor U9328 (N_9328,N_8946,N_8943);
and U9329 (N_9329,N_8247,N_8215);
nor U9330 (N_9330,N_8317,N_8699);
nor U9331 (N_9331,N_8508,N_8353);
or U9332 (N_9332,N_8442,N_8212);
xor U9333 (N_9333,N_8239,N_8689);
and U9334 (N_9334,N_8485,N_8031);
nor U9335 (N_9335,N_8521,N_8289);
or U9336 (N_9336,N_8189,N_8660);
nand U9337 (N_9337,N_8587,N_8705);
and U9338 (N_9338,N_8722,N_8765);
xnor U9339 (N_9339,N_8797,N_8292);
or U9340 (N_9340,N_8230,N_8760);
xnor U9341 (N_9341,N_8075,N_8718);
nand U9342 (N_9342,N_8858,N_8604);
nor U9343 (N_9343,N_8520,N_8808);
nand U9344 (N_9344,N_8823,N_8273);
or U9345 (N_9345,N_8315,N_8517);
xor U9346 (N_9346,N_8625,N_8614);
nor U9347 (N_9347,N_8695,N_8259);
nor U9348 (N_9348,N_8977,N_8986);
nand U9349 (N_9349,N_8827,N_8533);
nand U9350 (N_9350,N_8107,N_8274);
or U9351 (N_9351,N_8162,N_8150);
nand U9352 (N_9352,N_8869,N_8941);
nor U9353 (N_9353,N_8527,N_8293);
nor U9354 (N_9354,N_8569,N_8201);
and U9355 (N_9355,N_8555,N_8038);
and U9356 (N_9356,N_8736,N_8809);
nand U9357 (N_9357,N_8082,N_8136);
xnor U9358 (N_9358,N_8011,N_8213);
nand U9359 (N_9359,N_8002,N_8079);
nand U9360 (N_9360,N_8753,N_8458);
and U9361 (N_9361,N_8451,N_8182);
nor U9362 (N_9362,N_8667,N_8330);
and U9363 (N_9363,N_8688,N_8071);
nor U9364 (N_9364,N_8037,N_8160);
nand U9365 (N_9365,N_8863,N_8574);
nor U9366 (N_9366,N_8964,N_8362);
or U9367 (N_9367,N_8153,N_8445);
nor U9368 (N_9368,N_8872,N_8880);
nor U9369 (N_9369,N_8085,N_8626);
xor U9370 (N_9370,N_8932,N_8605);
or U9371 (N_9371,N_8122,N_8340);
and U9372 (N_9372,N_8397,N_8600);
or U9373 (N_9373,N_8938,N_8074);
xor U9374 (N_9374,N_8034,N_8538);
or U9375 (N_9375,N_8665,N_8518);
or U9376 (N_9376,N_8416,N_8772);
nand U9377 (N_9377,N_8454,N_8525);
or U9378 (N_9378,N_8814,N_8714);
nand U9379 (N_9379,N_8745,N_8405);
and U9380 (N_9380,N_8095,N_8720);
and U9381 (N_9381,N_8544,N_8636);
or U9382 (N_9382,N_8404,N_8326);
and U9383 (N_9383,N_8012,N_8394);
nand U9384 (N_9384,N_8139,N_8178);
or U9385 (N_9385,N_8656,N_8545);
or U9386 (N_9386,N_8862,N_8481);
xnor U9387 (N_9387,N_8024,N_8272);
xnor U9388 (N_9388,N_8117,N_8440);
or U9389 (N_9389,N_8088,N_8583);
nand U9390 (N_9390,N_8138,N_8267);
nor U9391 (N_9391,N_8907,N_8548);
nand U9392 (N_9392,N_8644,N_8260);
or U9393 (N_9393,N_8542,N_8496);
nor U9394 (N_9394,N_8565,N_8171);
xnor U9395 (N_9395,N_8347,N_8402);
nand U9396 (N_9396,N_8351,N_8041);
xnor U9397 (N_9397,N_8288,N_8462);
nand U9398 (N_9398,N_8235,N_8535);
xor U9399 (N_9399,N_8336,N_8401);
and U9400 (N_9400,N_8775,N_8328);
nand U9401 (N_9401,N_8962,N_8783);
xnor U9402 (N_9402,N_8191,N_8474);
nand U9403 (N_9403,N_8761,N_8541);
and U9404 (N_9404,N_8712,N_8246);
or U9405 (N_9405,N_8155,N_8030);
nor U9406 (N_9406,N_8494,N_8471);
nor U9407 (N_9407,N_8337,N_8489);
nor U9408 (N_9408,N_8130,N_8018);
xnor U9409 (N_9409,N_8904,N_8256);
nand U9410 (N_9410,N_8390,N_8486);
nor U9411 (N_9411,N_8622,N_8557);
nand U9412 (N_9412,N_8248,N_8746);
or U9413 (N_9413,N_8185,N_8118);
nand U9414 (N_9414,N_8623,N_8452);
xnor U9415 (N_9415,N_8281,N_8231);
nor U9416 (N_9416,N_8933,N_8832);
xor U9417 (N_9417,N_8324,N_8831);
and U9418 (N_9418,N_8674,N_8866);
or U9419 (N_9419,N_8491,N_8524);
nand U9420 (N_9420,N_8514,N_8983);
or U9421 (N_9421,N_8515,N_8199);
nand U9422 (N_9422,N_8876,N_8553);
nor U9423 (N_9423,N_8344,N_8291);
nand U9424 (N_9424,N_8512,N_8070);
and U9425 (N_9425,N_8383,N_8457);
or U9426 (N_9426,N_8826,N_8429);
nand U9427 (N_9427,N_8241,N_8707);
nor U9428 (N_9428,N_8790,N_8479);
xnor U9429 (N_9429,N_8999,N_8804);
nor U9430 (N_9430,N_8534,N_8242);
xor U9431 (N_9431,N_8126,N_8659);
xor U9432 (N_9432,N_8633,N_8989);
or U9433 (N_9433,N_8886,N_8645);
xor U9434 (N_9434,N_8501,N_8666);
nor U9435 (N_9435,N_8848,N_8295);
or U9436 (N_9436,N_8232,N_8413);
xnor U9437 (N_9437,N_8166,N_8108);
and U9438 (N_9438,N_8207,N_8129);
nor U9439 (N_9439,N_8575,N_8238);
or U9440 (N_9440,N_8306,N_8219);
xor U9441 (N_9441,N_8675,N_8145);
nor U9442 (N_9442,N_8884,N_8820);
xor U9443 (N_9443,N_8123,N_8009);
nand U9444 (N_9444,N_8936,N_8631);
xor U9445 (N_9445,N_8664,N_8926);
and U9446 (N_9446,N_8276,N_8222);
and U9447 (N_9447,N_8818,N_8728);
nor U9448 (N_9448,N_8973,N_8951);
and U9449 (N_9449,N_8871,N_8637);
and U9450 (N_9450,N_8709,N_8816);
and U9451 (N_9451,N_8188,N_8257);
nand U9452 (N_9452,N_8899,N_8927);
nor U9453 (N_9453,N_8696,N_8467);
xnor U9454 (N_9454,N_8530,N_8060);
or U9455 (N_9455,N_8985,N_8566);
nand U9456 (N_9456,N_8393,N_8209);
nor U9457 (N_9457,N_8708,N_8673);
nor U9458 (N_9458,N_8174,N_8982);
nor U9459 (N_9459,N_8632,N_8668);
xnor U9460 (N_9460,N_8352,N_8890);
or U9461 (N_9461,N_8465,N_8200);
and U9462 (N_9462,N_8463,N_8482);
or U9463 (N_9463,N_8957,N_8713);
xnor U9464 (N_9464,N_8010,N_8216);
nand U9465 (N_9465,N_8526,N_8810);
nor U9466 (N_9466,N_8310,N_8875);
xnor U9467 (N_9467,N_8780,N_8920);
nor U9468 (N_9468,N_8706,N_8596);
or U9469 (N_9469,N_8045,N_8094);
xor U9470 (N_9470,N_8620,N_8923);
xor U9471 (N_9471,N_8802,N_8861);
xor U9472 (N_9472,N_8303,N_8100);
xnor U9473 (N_9473,N_8417,N_8299);
and U9474 (N_9474,N_8654,N_8678);
nor U9475 (N_9475,N_8502,N_8911);
nor U9476 (N_9476,N_8834,N_8897);
nand U9477 (N_9477,N_8424,N_8047);
and U9478 (N_9478,N_8671,N_8629);
xnor U9479 (N_9479,N_8948,N_8400);
and U9480 (N_9480,N_8560,N_8987);
xnor U9481 (N_9481,N_8137,N_8086);
nor U9482 (N_9482,N_8493,N_8469);
nand U9483 (N_9483,N_8176,N_8597);
xor U9484 (N_9484,N_8023,N_8331);
or U9485 (N_9485,N_8322,N_8683);
xnor U9486 (N_9486,N_8410,N_8275);
nor U9487 (N_9487,N_8960,N_8949);
xnor U9488 (N_9488,N_8738,N_8860);
nor U9489 (N_9489,N_8588,N_8833);
and U9490 (N_9490,N_8882,N_8399);
nor U9491 (N_9491,N_8068,N_8354);
or U9492 (N_9492,N_8127,N_8388);
and U9493 (N_9493,N_8146,N_8953);
xor U9494 (N_9494,N_8335,N_8801);
nor U9495 (N_9495,N_8101,N_8443);
and U9496 (N_9496,N_8847,N_8643);
nand U9497 (N_9497,N_8734,N_8998);
nor U9498 (N_9498,N_8057,N_8430);
xor U9499 (N_9499,N_8338,N_8483);
nor U9500 (N_9500,N_8451,N_8421);
and U9501 (N_9501,N_8967,N_8471);
or U9502 (N_9502,N_8416,N_8664);
and U9503 (N_9503,N_8162,N_8055);
and U9504 (N_9504,N_8116,N_8944);
and U9505 (N_9505,N_8347,N_8602);
nand U9506 (N_9506,N_8281,N_8423);
or U9507 (N_9507,N_8904,N_8779);
nor U9508 (N_9508,N_8001,N_8908);
nand U9509 (N_9509,N_8524,N_8028);
xnor U9510 (N_9510,N_8758,N_8179);
or U9511 (N_9511,N_8047,N_8123);
nor U9512 (N_9512,N_8431,N_8992);
xnor U9513 (N_9513,N_8926,N_8916);
nor U9514 (N_9514,N_8229,N_8673);
nand U9515 (N_9515,N_8364,N_8727);
or U9516 (N_9516,N_8210,N_8117);
nand U9517 (N_9517,N_8758,N_8304);
nor U9518 (N_9518,N_8339,N_8868);
or U9519 (N_9519,N_8503,N_8074);
nor U9520 (N_9520,N_8641,N_8623);
nor U9521 (N_9521,N_8192,N_8320);
or U9522 (N_9522,N_8925,N_8922);
xor U9523 (N_9523,N_8480,N_8479);
nor U9524 (N_9524,N_8434,N_8617);
and U9525 (N_9525,N_8297,N_8483);
xor U9526 (N_9526,N_8494,N_8835);
and U9527 (N_9527,N_8584,N_8726);
xnor U9528 (N_9528,N_8126,N_8855);
nand U9529 (N_9529,N_8414,N_8956);
or U9530 (N_9530,N_8272,N_8436);
or U9531 (N_9531,N_8736,N_8285);
nand U9532 (N_9532,N_8289,N_8931);
or U9533 (N_9533,N_8002,N_8054);
xnor U9534 (N_9534,N_8012,N_8683);
xnor U9535 (N_9535,N_8125,N_8861);
or U9536 (N_9536,N_8718,N_8728);
and U9537 (N_9537,N_8188,N_8308);
xor U9538 (N_9538,N_8425,N_8137);
nand U9539 (N_9539,N_8676,N_8624);
nor U9540 (N_9540,N_8742,N_8278);
nand U9541 (N_9541,N_8650,N_8522);
nor U9542 (N_9542,N_8910,N_8745);
or U9543 (N_9543,N_8594,N_8964);
xnor U9544 (N_9544,N_8021,N_8538);
xnor U9545 (N_9545,N_8207,N_8440);
and U9546 (N_9546,N_8956,N_8481);
nor U9547 (N_9547,N_8312,N_8774);
nor U9548 (N_9548,N_8896,N_8291);
or U9549 (N_9549,N_8114,N_8344);
or U9550 (N_9550,N_8238,N_8943);
xnor U9551 (N_9551,N_8018,N_8174);
nand U9552 (N_9552,N_8537,N_8795);
xor U9553 (N_9553,N_8997,N_8123);
xor U9554 (N_9554,N_8212,N_8959);
nand U9555 (N_9555,N_8872,N_8853);
xor U9556 (N_9556,N_8894,N_8300);
or U9557 (N_9557,N_8634,N_8415);
xnor U9558 (N_9558,N_8283,N_8237);
or U9559 (N_9559,N_8831,N_8587);
nand U9560 (N_9560,N_8527,N_8509);
and U9561 (N_9561,N_8960,N_8435);
nor U9562 (N_9562,N_8888,N_8713);
nor U9563 (N_9563,N_8406,N_8604);
or U9564 (N_9564,N_8993,N_8233);
or U9565 (N_9565,N_8714,N_8966);
nor U9566 (N_9566,N_8838,N_8977);
and U9567 (N_9567,N_8102,N_8790);
xor U9568 (N_9568,N_8457,N_8370);
xor U9569 (N_9569,N_8832,N_8158);
xnor U9570 (N_9570,N_8612,N_8042);
or U9571 (N_9571,N_8017,N_8109);
and U9572 (N_9572,N_8153,N_8261);
or U9573 (N_9573,N_8394,N_8798);
or U9574 (N_9574,N_8553,N_8294);
and U9575 (N_9575,N_8371,N_8860);
xnor U9576 (N_9576,N_8888,N_8413);
and U9577 (N_9577,N_8718,N_8865);
and U9578 (N_9578,N_8712,N_8399);
and U9579 (N_9579,N_8144,N_8227);
nor U9580 (N_9580,N_8764,N_8483);
nand U9581 (N_9581,N_8828,N_8271);
nor U9582 (N_9582,N_8127,N_8261);
or U9583 (N_9583,N_8449,N_8675);
xnor U9584 (N_9584,N_8283,N_8343);
or U9585 (N_9585,N_8705,N_8777);
nand U9586 (N_9586,N_8129,N_8005);
nand U9587 (N_9587,N_8964,N_8949);
or U9588 (N_9588,N_8757,N_8823);
or U9589 (N_9589,N_8819,N_8445);
and U9590 (N_9590,N_8047,N_8379);
xnor U9591 (N_9591,N_8751,N_8412);
xnor U9592 (N_9592,N_8444,N_8889);
nor U9593 (N_9593,N_8913,N_8375);
nand U9594 (N_9594,N_8525,N_8911);
and U9595 (N_9595,N_8940,N_8910);
and U9596 (N_9596,N_8627,N_8649);
or U9597 (N_9597,N_8470,N_8495);
nor U9598 (N_9598,N_8949,N_8568);
nor U9599 (N_9599,N_8264,N_8988);
nor U9600 (N_9600,N_8219,N_8842);
nand U9601 (N_9601,N_8535,N_8857);
and U9602 (N_9602,N_8365,N_8524);
and U9603 (N_9603,N_8789,N_8320);
nor U9604 (N_9604,N_8484,N_8439);
or U9605 (N_9605,N_8981,N_8183);
nand U9606 (N_9606,N_8484,N_8882);
nand U9607 (N_9607,N_8911,N_8825);
and U9608 (N_9608,N_8659,N_8651);
xor U9609 (N_9609,N_8044,N_8978);
xor U9610 (N_9610,N_8898,N_8909);
and U9611 (N_9611,N_8446,N_8032);
nand U9612 (N_9612,N_8546,N_8278);
and U9613 (N_9613,N_8858,N_8606);
nand U9614 (N_9614,N_8116,N_8083);
or U9615 (N_9615,N_8753,N_8771);
and U9616 (N_9616,N_8665,N_8929);
and U9617 (N_9617,N_8869,N_8561);
nand U9618 (N_9618,N_8214,N_8931);
or U9619 (N_9619,N_8847,N_8096);
and U9620 (N_9620,N_8367,N_8132);
and U9621 (N_9621,N_8412,N_8445);
nor U9622 (N_9622,N_8970,N_8408);
xor U9623 (N_9623,N_8877,N_8376);
nor U9624 (N_9624,N_8739,N_8250);
xor U9625 (N_9625,N_8878,N_8923);
or U9626 (N_9626,N_8413,N_8338);
and U9627 (N_9627,N_8869,N_8564);
nor U9628 (N_9628,N_8041,N_8131);
nand U9629 (N_9629,N_8569,N_8052);
nor U9630 (N_9630,N_8095,N_8918);
or U9631 (N_9631,N_8153,N_8297);
or U9632 (N_9632,N_8675,N_8415);
nand U9633 (N_9633,N_8057,N_8224);
nor U9634 (N_9634,N_8879,N_8277);
or U9635 (N_9635,N_8166,N_8144);
and U9636 (N_9636,N_8604,N_8070);
nor U9637 (N_9637,N_8701,N_8305);
nand U9638 (N_9638,N_8289,N_8044);
nand U9639 (N_9639,N_8813,N_8730);
xor U9640 (N_9640,N_8349,N_8861);
or U9641 (N_9641,N_8483,N_8093);
nand U9642 (N_9642,N_8201,N_8142);
nand U9643 (N_9643,N_8260,N_8054);
nor U9644 (N_9644,N_8345,N_8404);
xnor U9645 (N_9645,N_8553,N_8617);
nand U9646 (N_9646,N_8017,N_8892);
xor U9647 (N_9647,N_8124,N_8810);
xnor U9648 (N_9648,N_8641,N_8525);
nor U9649 (N_9649,N_8090,N_8072);
and U9650 (N_9650,N_8453,N_8526);
and U9651 (N_9651,N_8554,N_8117);
nand U9652 (N_9652,N_8729,N_8181);
and U9653 (N_9653,N_8394,N_8997);
xnor U9654 (N_9654,N_8340,N_8575);
nand U9655 (N_9655,N_8338,N_8831);
nand U9656 (N_9656,N_8934,N_8474);
nor U9657 (N_9657,N_8133,N_8730);
or U9658 (N_9658,N_8226,N_8511);
nor U9659 (N_9659,N_8505,N_8000);
xnor U9660 (N_9660,N_8410,N_8346);
nor U9661 (N_9661,N_8799,N_8161);
nor U9662 (N_9662,N_8476,N_8150);
or U9663 (N_9663,N_8322,N_8111);
xnor U9664 (N_9664,N_8068,N_8773);
nand U9665 (N_9665,N_8548,N_8833);
xor U9666 (N_9666,N_8741,N_8245);
nand U9667 (N_9667,N_8084,N_8137);
nand U9668 (N_9668,N_8577,N_8845);
or U9669 (N_9669,N_8722,N_8742);
nor U9670 (N_9670,N_8432,N_8842);
and U9671 (N_9671,N_8006,N_8812);
nand U9672 (N_9672,N_8318,N_8533);
and U9673 (N_9673,N_8637,N_8338);
xor U9674 (N_9674,N_8414,N_8661);
nand U9675 (N_9675,N_8965,N_8445);
and U9676 (N_9676,N_8959,N_8569);
nand U9677 (N_9677,N_8848,N_8915);
or U9678 (N_9678,N_8698,N_8724);
nand U9679 (N_9679,N_8913,N_8393);
nor U9680 (N_9680,N_8672,N_8099);
nor U9681 (N_9681,N_8087,N_8441);
xor U9682 (N_9682,N_8156,N_8521);
xnor U9683 (N_9683,N_8413,N_8276);
or U9684 (N_9684,N_8912,N_8158);
xnor U9685 (N_9685,N_8826,N_8401);
and U9686 (N_9686,N_8429,N_8831);
or U9687 (N_9687,N_8746,N_8934);
nand U9688 (N_9688,N_8858,N_8288);
xor U9689 (N_9689,N_8591,N_8123);
nor U9690 (N_9690,N_8294,N_8310);
or U9691 (N_9691,N_8100,N_8266);
nand U9692 (N_9692,N_8237,N_8569);
and U9693 (N_9693,N_8637,N_8989);
and U9694 (N_9694,N_8481,N_8302);
nor U9695 (N_9695,N_8916,N_8691);
xnor U9696 (N_9696,N_8572,N_8334);
and U9697 (N_9697,N_8388,N_8021);
and U9698 (N_9698,N_8490,N_8922);
or U9699 (N_9699,N_8667,N_8985);
xor U9700 (N_9700,N_8474,N_8704);
or U9701 (N_9701,N_8359,N_8302);
or U9702 (N_9702,N_8255,N_8208);
nand U9703 (N_9703,N_8518,N_8434);
xor U9704 (N_9704,N_8811,N_8988);
and U9705 (N_9705,N_8837,N_8075);
nor U9706 (N_9706,N_8224,N_8060);
xnor U9707 (N_9707,N_8925,N_8619);
xor U9708 (N_9708,N_8519,N_8321);
and U9709 (N_9709,N_8593,N_8297);
and U9710 (N_9710,N_8352,N_8648);
nand U9711 (N_9711,N_8294,N_8442);
nor U9712 (N_9712,N_8429,N_8236);
and U9713 (N_9713,N_8703,N_8785);
nand U9714 (N_9714,N_8708,N_8713);
xor U9715 (N_9715,N_8080,N_8184);
nand U9716 (N_9716,N_8455,N_8861);
nand U9717 (N_9717,N_8048,N_8670);
nand U9718 (N_9718,N_8823,N_8070);
and U9719 (N_9719,N_8411,N_8577);
nor U9720 (N_9720,N_8387,N_8628);
or U9721 (N_9721,N_8290,N_8304);
or U9722 (N_9722,N_8514,N_8371);
and U9723 (N_9723,N_8366,N_8883);
nor U9724 (N_9724,N_8554,N_8414);
or U9725 (N_9725,N_8413,N_8403);
nand U9726 (N_9726,N_8497,N_8783);
and U9727 (N_9727,N_8932,N_8634);
or U9728 (N_9728,N_8275,N_8456);
xnor U9729 (N_9729,N_8312,N_8391);
or U9730 (N_9730,N_8446,N_8207);
and U9731 (N_9731,N_8469,N_8103);
nor U9732 (N_9732,N_8009,N_8799);
xor U9733 (N_9733,N_8891,N_8973);
or U9734 (N_9734,N_8117,N_8957);
and U9735 (N_9735,N_8355,N_8963);
nor U9736 (N_9736,N_8615,N_8779);
nor U9737 (N_9737,N_8562,N_8212);
or U9738 (N_9738,N_8041,N_8570);
xor U9739 (N_9739,N_8398,N_8096);
nor U9740 (N_9740,N_8101,N_8427);
nor U9741 (N_9741,N_8466,N_8719);
or U9742 (N_9742,N_8708,N_8956);
nand U9743 (N_9743,N_8650,N_8156);
xnor U9744 (N_9744,N_8193,N_8034);
xor U9745 (N_9745,N_8651,N_8860);
and U9746 (N_9746,N_8219,N_8670);
or U9747 (N_9747,N_8790,N_8465);
nor U9748 (N_9748,N_8076,N_8482);
nor U9749 (N_9749,N_8594,N_8134);
and U9750 (N_9750,N_8285,N_8317);
xnor U9751 (N_9751,N_8107,N_8918);
xnor U9752 (N_9752,N_8651,N_8068);
xnor U9753 (N_9753,N_8496,N_8899);
nand U9754 (N_9754,N_8005,N_8907);
or U9755 (N_9755,N_8264,N_8036);
nand U9756 (N_9756,N_8904,N_8553);
or U9757 (N_9757,N_8914,N_8641);
or U9758 (N_9758,N_8327,N_8708);
or U9759 (N_9759,N_8742,N_8135);
or U9760 (N_9760,N_8548,N_8005);
xor U9761 (N_9761,N_8111,N_8128);
or U9762 (N_9762,N_8893,N_8563);
nand U9763 (N_9763,N_8043,N_8654);
xor U9764 (N_9764,N_8870,N_8634);
xnor U9765 (N_9765,N_8510,N_8102);
nor U9766 (N_9766,N_8038,N_8147);
nor U9767 (N_9767,N_8419,N_8496);
xor U9768 (N_9768,N_8318,N_8201);
xor U9769 (N_9769,N_8801,N_8872);
nor U9770 (N_9770,N_8012,N_8439);
and U9771 (N_9771,N_8091,N_8167);
nor U9772 (N_9772,N_8972,N_8944);
nand U9773 (N_9773,N_8311,N_8996);
xnor U9774 (N_9774,N_8657,N_8604);
xor U9775 (N_9775,N_8901,N_8182);
and U9776 (N_9776,N_8762,N_8247);
or U9777 (N_9777,N_8287,N_8790);
and U9778 (N_9778,N_8336,N_8669);
nand U9779 (N_9779,N_8884,N_8039);
and U9780 (N_9780,N_8845,N_8052);
and U9781 (N_9781,N_8832,N_8378);
nand U9782 (N_9782,N_8366,N_8637);
and U9783 (N_9783,N_8243,N_8867);
or U9784 (N_9784,N_8143,N_8632);
nand U9785 (N_9785,N_8310,N_8528);
and U9786 (N_9786,N_8055,N_8465);
nor U9787 (N_9787,N_8739,N_8826);
or U9788 (N_9788,N_8886,N_8901);
nor U9789 (N_9789,N_8206,N_8490);
or U9790 (N_9790,N_8674,N_8806);
or U9791 (N_9791,N_8676,N_8841);
xnor U9792 (N_9792,N_8480,N_8662);
nor U9793 (N_9793,N_8468,N_8154);
nand U9794 (N_9794,N_8384,N_8154);
xnor U9795 (N_9795,N_8055,N_8090);
and U9796 (N_9796,N_8844,N_8230);
nor U9797 (N_9797,N_8450,N_8537);
xnor U9798 (N_9798,N_8583,N_8484);
or U9799 (N_9799,N_8787,N_8471);
and U9800 (N_9800,N_8445,N_8454);
xor U9801 (N_9801,N_8766,N_8370);
xor U9802 (N_9802,N_8991,N_8935);
and U9803 (N_9803,N_8287,N_8818);
and U9804 (N_9804,N_8754,N_8881);
or U9805 (N_9805,N_8001,N_8794);
or U9806 (N_9806,N_8058,N_8309);
or U9807 (N_9807,N_8291,N_8084);
nand U9808 (N_9808,N_8742,N_8011);
nor U9809 (N_9809,N_8761,N_8528);
and U9810 (N_9810,N_8495,N_8925);
xnor U9811 (N_9811,N_8837,N_8239);
xor U9812 (N_9812,N_8157,N_8958);
nor U9813 (N_9813,N_8056,N_8559);
or U9814 (N_9814,N_8349,N_8581);
xnor U9815 (N_9815,N_8747,N_8376);
or U9816 (N_9816,N_8303,N_8055);
nor U9817 (N_9817,N_8502,N_8559);
or U9818 (N_9818,N_8163,N_8720);
xnor U9819 (N_9819,N_8320,N_8352);
nand U9820 (N_9820,N_8327,N_8602);
and U9821 (N_9821,N_8534,N_8217);
and U9822 (N_9822,N_8148,N_8682);
nor U9823 (N_9823,N_8137,N_8824);
or U9824 (N_9824,N_8837,N_8973);
and U9825 (N_9825,N_8140,N_8248);
and U9826 (N_9826,N_8420,N_8387);
and U9827 (N_9827,N_8563,N_8686);
nand U9828 (N_9828,N_8238,N_8057);
and U9829 (N_9829,N_8618,N_8821);
nor U9830 (N_9830,N_8764,N_8336);
and U9831 (N_9831,N_8474,N_8417);
nor U9832 (N_9832,N_8209,N_8755);
and U9833 (N_9833,N_8586,N_8401);
and U9834 (N_9834,N_8594,N_8869);
nand U9835 (N_9835,N_8861,N_8115);
and U9836 (N_9836,N_8417,N_8612);
and U9837 (N_9837,N_8068,N_8367);
or U9838 (N_9838,N_8192,N_8325);
nor U9839 (N_9839,N_8990,N_8862);
xor U9840 (N_9840,N_8713,N_8473);
nand U9841 (N_9841,N_8386,N_8761);
xnor U9842 (N_9842,N_8360,N_8191);
or U9843 (N_9843,N_8538,N_8226);
xor U9844 (N_9844,N_8727,N_8446);
xnor U9845 (N_9845,N_8652,N_8071);
nand U9846 (N_9846,N_8024,N_8780);
or U9847 (N_9847,N_8267,N_8650);
nand U9848 (N_9848,N_8089,N_8214);
xor U9849 (N_9849,N_8400,N_8541);
or U9850 (N_9850,N_8340,N_8445);
xor U9851 (N_9851,N_8893,N_8064);
and U9852 (N_9852,N_8729,N_8030);
nand U9853 (N_9853,N_8964,N_8838);
xor U9854 (N_9854,N_8316,N_8321);
nand U9855 (N_9855,N_8776,N_8362);
or U9856 (N_9856,N_8265,N_8063);
nand U9857 (N_9857,N_8937,N_8465);
xnor U9858 (N_9858,N_8136,N_8484);
xor U9859 (N_9859,N_8177,N_8060);
xnor U9860 (N_9860,N_8121,N_8434);
or U9861 (N_9861,N_8719,N_8527);
or U9862 (N_9862,N_8731,N_8480);
or U9863 (N_9863,N_8491,N_8315);
xnor U9864 (N_9864,N_8659,N_8116);
nor U9865 (N_9865,N_8898,N_8352);
and U9866 (N_9866,N_8785,N_8064);
nand U9867 (N_9867,N_8564,N_8309);
nor U9868 (N_9868,N_8131,N_8487);
or U9869 (N_9869,N_8757,N_8143);
xnor U9870 (N_9870,N_8016,N_8130);
and U9871 (N_9871,N_8890,N_8076);
nand U9872 (N_9872,N_8928,N_8656);
or U9873 (N_9873,N_8784,N_8797);
or U9874 (N_9874,N_8925,N_8001);
nor U9875 (N_9875,N_8817,N_8311);
nand U9876 (N_9876,N_8475,N_8677);
nor U9877 (N_9877,N_8593,N_8148);
and U9878 (N_9878,N_8459,N_8633);
xnor U9879 (N_9879,N_8751,N_8041);
xnor U9880 (N_9880,N_8251,N_8074);
xnor U9881 (N_9881,N_8237,N_8138);
nor U9882 (N_9882,N_8032,N_8604);
xor U9883 (N_9883,N_8087,N_8690);
xnor U9884 (N_9884,N_8544,N_8490);
or U9885 (N_9885,N_8565,N_8292);
nand U9886 (N_9886,N_8104,N_8381);
nor U9887 (N_9887,N_8252,N_8048);
nand U9888 (N_9888,N_8654,N_8203);
nand U9889 (N_9889,N_8277,N_8856);
nand U9890 (N_9890,N_8012,N_8300);
or U9891 (N_9891,N_8303,N_8631);
or U9892 (N_9892,N_8379,N_8560);
nand U9893 (N_9893,N_8342,N_8671);
nand U9894 (N_9894,N_8840,N_8825);
nor U9895 (N_9895,N_8528,N_8718);
nand U9896 (N_9896,N_8348,N_8644);
nor U9897 (N_9897,N_8580,N_8135);
or U9898 (N_9898,N_8489,N_8321);
nand U9899 (N_9899,N_8713,N_8448);
nand U9900 (N_9900,N_8570,N_8644);
xor U9901 (N_9901,N_8667,N_8104);
nor U9902 (N_9902,N_8589,N_8101);
nor U9903 (N_9903,N_8400,N_8715);
nor U9904 (N_9904,N_8087,N_8259);
nor U9905 (N_9905,N_8317,N_8329);
nand U9906 (N_9906,N_8346,N_8429);
or U9907 (N_9907,N_8316,N_8798);
xor U9908 (N_9908,N_8627,N_8793);
nor U9909 (N_9909,N_8401,N_8870);
xnor U9910 (N_9910,N_8875,N_8559);
and U9911 (N_9911,N_8573,N_8237);
xor U9912 (N_9912,N_8052,N_8341);
xor U9913 (N_9913,N_8364,N_8467);
nand U9914 (N_9914,N_8815,N_8658);
or U9915 (N_9915,N_8127,N_8396);
or U9916 (N_9916,N_8309,N_8376);
nor U9917 (N_9917,N_8368,N_8622);
xor U9918 (N_9918,N_8400,N_8987);
nand U9919 (N_9919,N_8210,N_8364);
xor U9920 (N_9920,N_8525,N_8819);
xor U9921 (N_9921,N_8218,N_8363);
or U9922 (N_9922,N_8200,N_8211);
or U9923 (N_9923,N_8066,N_8028);
or U9924 (N_9924,N_8791,N_8111);
and U9925 (N_9925,N_8203,N_8266);
nand U9926 (N_9926,N_8581,N_8044);
or U9927 (N_9927,N_8426,N_8360);
nand U9928 (N_9928,N_8070,N_8356);
xnor U9929 (N_9929,N_8983,N_8509);
or U9930 (N_9930,N_8338,N_8233);
and U9931 (N_9931,N_8579,N_8296);
and U9932 (N_9932,N_8988,N_8885);
xor U9933 (N_9933,N_8538,N_8058);
or U9934 (N_9934,N_8954,N_8333);
xor U9935 (N_9935,N_8075,N_8359);
and U9936 (N_9936,N_8890,N_8977);
nand U9937 (N_9937,N_8641,N_8187);
or U9938 (N_9938,N_8853,N_8006);
nor U9939 (N_9939,N_8891,N_8193);
nand U9940 (N_9940,N_8674,N_8663);
xor U9941 (N_9941,N_8730,N_8070);
or U9942 (N_9942,N_8772,N_8508);
nand U9943 (N_9943,N_8331,N_8972);
or U9944 (N_9944,N_8293,N_8406);
nand U9945 (N_9945,N_8666,N_8476);
or U9946 (N_9946,N_8654,N_8598);
and U9947 (N_9947,N_8376,N_8976);
or U9948 (N_9948,N_8530,N_8568);
or U9949 (N_9949,N_8166,N_8457);
and U9950 (N_9950,N_8012,N_8686);
and U9951 (N_9951,N_8776,N_8573);
or U9952 (N_9952,N_8988,N_8468);
or U9953 (N_9953,N_8381,N_8035);
nor U9954 (N_9954,N_8221,N_8829);
nand U9955 (N_9955,N_8407,N_8575);
nor U9956 (N_9956,N_8815,N_8558);
and U9957 (N_9957,N_8025,N_8285);
xnor U9958 (N_9958,N_8784,N_8255);
or U9959 (N_9959,N_8873,N_8505);
or U9960 (N_9960,N_8571,N_8979);
nor U9961 (N_9961,N_8606,N_8466);
or U9962 (N_9962,N_8981,N_8654);
and U9963 (N_9963,N_8672,N_8581);
xor U9964 (N_9964,N_8004,N_8876);
and U9965 (N_9965,N_8590,N_8363);
nor U9966 (N_9966,N_8363,N_8892);
nand U9967 (N_9967,N_8694,N_8834);
xnor U9968 (N_9968,N_8308,N_8118);
or U9969 (N_9969,N_8988,N_8217);
or U9970 (N_9970,N_8266,N_8420);
nand U9971 (N_9971,N_8581,N_8836);
nand U9972 (N_9972,N_8669,N_8593);
nand U9973 (N_9973,N_8935,N_8514);
xor U9974 (N_9974,N_8311,N_8027);
nand U9975 (N_9975,N_8216,N_8484);
xor U9976 (N_9976,N_8969,N_8346);
or U9977 (N_9977,N_8112,N_8201);
nor U9978 (N_9978,N_8901,N_8796);
and U9979 (N_9979,N_8207,N_8101);
xnor U9980 (N_9980,N_8487,N_8950);
nor U9981 (N_9981,N_8018,N_8214);
nand U9982 (N_9982,N_8817,N_8714);
and U9983 (N_9983,N_8114,N_8959);
nor U9984 (N_9984,N_8310,N_8230);
nor U9985 (N_9985,N_8307,N_8048);
and U9986 (N_9986,N_8531,N_8088);
nand U9987 (N_9987,N_8781,N_8973);
nor U9988 (N_9988,N_8945,N_8871);
and U9989 (N_9989,N_8965,N_8094);
and U9990 (N_9990,N_8322,N_8782);
nand U9991 (N_9991,N_8764,N_8644);
or U9992 (N_9992,N_8186,N_8004);
and U9993 (N_9993,N_8169,N_8759);
and U9994 (N_9994,N_8019,N_8035);
or U9995 (N_9995,N_8360,N_8852);
and U9996 (N_9996,N_8387,N_8319);
or U9997 (N_9997,N_8038,N_8251);
and U9998 (N_9998,N_8442,N_8618);
nor U9999 (N_9999,N_8407,N_8162);
nor U10000 (N_10000,N_9737,N_9070);
xor U10001 (N_10001,N_9058,N_9712);
or U10002 (N_10002,N_9738,N_9096);
nand U10003 (N_10003,N_9476,N_9972);
xnor U10004 (N_10004,N_9925,N_9966);
and U10005 (N_10005,N_9048,N_9587);
nor U10006 (N_10006,N_9185,N_9748);
or U10007 (N_10007,N_9574,N_9824);
xnor U10008 (N_10008,N_9817,N_9341);
nor U10009 (N_10009,N_9197,N_9195);
xor U10010 (N_10010,N_9324,N_9657);
and U10011 (N_10011,N_9434,N_9672);
or U10012 (N_10012,N_9991,N_9759);
nor U10013 (N_10013,N_9377,N_9273);
nor U10014 (N_10014,N_9219,N_9035);
nand U10015 (N_10015,N_9913,N_9045);
xor U10016 (N_10016,N_9911,N_9469);
and U10017 (N_10017,N_9092,N_9255);
nor U10018 (N_10018,N_9477,N_9954);
xor U10019 (N_10019,N_9366,N_9566);
nor U10020 (N_10020,N_9177,N_9963);
or U10021 (N_10021,N_9472,N_9387);
xnor U10022 (N_10022,N_9621,N_9208);
nor U10023 (N_10023,N_9025,N_9021);
or U10024 (N_10024,N_9711,N_9808);
or U10025 (N_10025,N_9589,N_9804);
or U10026 (N_10026,N_9551,N_9953);
nor U10027 (N_10027,N_9501,N_9344);
nor U10028 (N_10028,N_9281,N_9732);
and U10029 (N_10029,N_9989,N_9140);
xor U10030 (N_10030,N_9371,N_9723);
nand U10031 (N_10031,N_9073,N_9649);
xor U10032 (N_10032,N_9119,N_9405);
and U10033 (N_10033,N_9543,N_9661);
xnor U10034 (N_10034,N_9135,N_9293);
or U10035 (N_10035,N_9253,N_9625);
or U10036 (N_10036,N_9685,N_9796);
or U10037 (N_10037,N_9705,N_9463);
xnor U10038 (N_10038,N_9353,N_9651);
nand U10039 (N_10039,N_9006,N_9000);
and U10040 (N_10040,N_9342,N_9052);
nor U10041 (N_10041,N_9396,N_9165);
or U10042 (N_10042,N_9029,N_9181);
nand U10043 (N_10043,N_9532,N_9461);
xnor U10044 (N_10044,N_9013,N_9761);
and U10045 (N_10045,N_9794,N_9232);
and U10046 (N_10046,N_9334,N_9921);
or U10047 (N_10047,N_9065,N_9557);
xnor U10048 (N_10048,N_9294,N_9339);
nand U10049 (N_10049,N_9230,N_9388);
and U10050 (N_10050,N_9613,N_9784);
xnor U10051 (N_10051,N_9274,N_9949);
nand U10052 (N_10052,N_9320,N_9576);
nand U10053 (N_10053,N_9741,N_9162);
nand U10054 (N_10054,N_9571,N_9164);
xnor U10055 (N_10055,N_9414,N_9102);
xor U10056 (N_10056,N_9883,N_9053);
nor U10057 (N_10057,N_9871,N_9080);
nor U10058 (N_10058,N_9365,N_9179);
nand U10059 (N_10059,N_9533,N_9321);
or U10060 (N_10060,N_9504,N_9735);
and U10061 (N_10061,N_9585,N_9187);
xor U10062 (N_10062,N_9158,N_9731);
xor U10063 (N_10063,N_9858,N_9412);
and U10064 (N_10064,N_9724,N_9771);
nor U10065 (N_10065,N_9299,N_9718);
and U10066 (N_10066,N_9199,N_9999);
and U10067 (N_10067,N_9675,N_9357);
or U10068 (N_10068,N_9237,N_9751);
nor U10069 (N_10069,N_9774,N_9990);
nand U10070 (N_10070,N_9312,N_9516);
nand U10071 (N_10071,N_9236,N_9530);
or U10072 (N_10072,N_9482,N_9263);
or U10073 (N_10073,N_9245,N_9003);
nor U10074 (N_10074,N_9077,N_9929);
xor U10075 (N_10075,N_9581,N_9280);
nand U10076 (N_10076,N_9155,N_9359);
xor U10077 (N_10077,N_9257,N_9345);
nand U10078 (N_10078,N_9679,N_9934);
nor U10079 (N_10079,N_9389,N_9994);
or U10080 (N_10080,N_9746,N_9494);
nor U10081 (N_10081,N_9413,N_9818);
and U10082 (N_10082,N_9311,N_9959);
nand U10083 (N_10083,N_9578,N_9607);
nor U10084 (N_10084,N_9699,N_9307);
or U10085 (N_10085,N_9676,N_9089);
nor U10086 (N_10086,N_9580,N_9060);
nand U10087 (N_10087,N_9868,N_9957);
or U10088 (N_10088,N_9433,N_9876);
nor U10089 (N_10089,N_9196,N_9335);
nand U10090 (N_10090,N_9183,N_9665);
xnor U10091 (N_10091,N_9099,N_9787);
or U10092 (N_10092,N_9605,N_9684);
xnor U10093 (N_10093,N_9979,N_9776);
nand U10094 (N_10094,N_9832,N_9860);
nand U10095 (N_10095,N_9385,N_9854);
nand U10096 (N_10096,N_9023,N_9228);
xnor U10097 (N_10097,N_9127,N_9030);
nor U10098 (N_10098,N_9271,N_9662);
and U10099 (N_10099,N_9464,N_9659);
nor U10100 (N_10100,N_9419,N_9332);
xnor U10101 (N_10101,N_9515,N_9791);
or U10102 (N_10102,N_9424,N_9885);
or U10103 (N_10103,N_9430,N_9535);
or U10104 (N_10104,N_9638,N_9241);
xor U10105 (N_10105,N_9108,N_9295);
or U10106 (N_10106,N_9250,N_9351);
nand U10107 (N_10107,N_9628,N_9779);
nand U10108 (N_10108,N_9626,N_9895);
xor U10109 (N_10109,N_9548,N_9667);
nor U10110 (N_10110,N_9734,N_9286);
and U10111 (N_10111,N_9243,N_9756);
nor U10112 (N_10112,N_9207,N_9952);
xor U10113 (N_10113,N_9223,N_9213);
nor U10114 (N_10114,N_9570,N_9736);
nor U10115 (N_10115,N_9360,N_9141);
or U10116 (N_10116,N_9943,N_9766);
or U10117 (N_10117,N_9151,N_9123);
nand U10118 (N_10118,N_9289,N_9588);
and U10119 (N_10119,N_9471,N_9234);
xor U10120 (N_10120,N_9411,N_9869);
and U10121 (N_10121,N_9362,N_9846);
xor U10122 (N_10122,N_9752,N_9282);
and U10123 (N_10123,N_9121,N_9950);
and U10124 (N_10124,N_9034,N_9435);
nand U10125 (N_10125,N_9190,N_9802);
and U10126 (N_10126,N_9502,N_9850);
or U10127 (N_10127,N_9475,N_9393);
or U10128 (N_10128,N_9429,N_9483);
nor U10129 (N_10129,N_9009,N_9064);
nand U10130 (N_10130,N_9272,N_9349);
or U10131 (N_10131,N_9133,N_9401);
or U10132 (N_10132,N_9278,N_9720);
xor U10133 (N_10133,N_9800,N_9507);
xnor U10134 (N_10134,N_9379,N_9864);
nor U10135 (N_10135,N_9783,N_9998);
nor U10136 (N_10136,N_9806,N_9163);
nor U10137 (N_10137,N_9329,N_9128);
nand U10138 (N_10138,N_9773,N_9593);
and U10139 (N_10139,N_9923,N_9031);
nand U10140 (N_10140,N_9455,N_9848);
and U10141 (N_10141,N_9967,N_9384);
nand U10142 (N_10142,N_9325,N_9402);
xor U10143 (N_10143,N_9799,N_9235);
and U10144 (N_10144,N_9322,N_9193);
or U10145 (N_10145,N_9706,N_9634);
nand U10146 (N_10146,N_9085,N_9612);
xnor U10147 (N_10147,N_9652,N_9291);
or U10148 (N_10148,N_9452,N_9894);
nor U10149 (N_10149,N_9466,N_9105);
and U10150 (N_10150,N_9555,N_9372);
nor U10151 (N_10151,N_9202,N_9837);
nor U10152 (N_10152,N_9317,N_9100);
xor U10153 (N_10153,N_9691,N_9528);
nor U10154 (N_10154,N_9617,N_9572);
nand U10155 (N_10155,N_9873,N_9627);
xor U10156 (N_10156,N_9001,N_9015);
nor U10157 (N_10157,N_9238,N_9907);
nor U10158 (N_10158,N_9240,N_9258);
xnor U10159 (N_10159,N_9422,N_9326);
nand U10160 (N_10160,N_9906,N_9930);
xnor U10161 (N_10161,N_9426,N_9044);
nand U10162 (N_10162,N_9525,N_9057);
xor U10163 (N_10163,N_9936,N_9346);
and U10164 (N_10164,N_9304,N_9742);
nand U10165 (N_10165,N_9584,N_9231);
or U10166 (N_10166,N_9352,N_9109);
nand U10167 (N_10167,N_9714,N_9184);
nor U10168 (N_10168,N_9910,N_9693);
nand U10169 (N_10169,N_9664,N_9498);
xnor U10170 (N_10170,N_9117,N_9916);
and U10171 (N_10171,N_9855,N_9478);
and U10172 (N_10172,N_9319,N_9618);
nand U10173 (N_10173,N_9636,N_9409);
nand U10174 (N_10174,N_9188,N_9903);
xnor U10175 (N_10175,N_9562,N_9816);
nor U10176 (N_10176,N_9026,N_9768);
and U10177 (N_10177,N_9552,N_9150);
or U10178 (N_10178,N_9391,N_9394);
nor U10179 (N_10179,N_9630,N_9890);
or U10180 (N_10180,N_9054,N_9524);
nor U10181 (N_10181,N_9211,N_9702);
nor U10182 (N_10182,N_9609,N_9316);
nand U10183 (N_10183,N_9838,N_9086);
nor U10184 (N_10184,N_9602,N_9055);
and U10185 (N_10185,N_9194,N_9945);
nor U10186 (N_10186,N_9460,N_9840);
and U10187 (N_10187,N_9867,N_9596);
and U10188 (N_10188,N_9897,N_9915);
xnor U10189 (N_10189,N_9614,N_9018);
nor U10190 (N_10190,N_9892,N_9283);
nor U10191 (N_10191,N_9300,N_9306);
nor U10192 (N_10192,N_9347,N_9971);
or U10193 (N_10193,N_9601,N_9264);
or U10194 (N_10194,N_9423,N_9186);
and U10195 (N_10195,N_9172,N_9467);
xor U10196 (N_10196,N_9019,N_9169);
and U10197 (N_10197,N_9113,N_9110);
nand U10198 (N_10198,N_9813,N_9677);
xnor U10199 (N_10199,N_9616,N_9069);
and U10200 (N_10200,N_9719,N_9681);
or U10201 (N_10201,N_9451,N_9459);
xnor U10202 (N_10202,N_9523,N_9658);
xnor U10203 (N_10203,N_9275,N_9062);
xor U10204 (N_10204,N_9399,N_9743);
nand U10205 (N_10205,N_9042,N_9554);
or U10206 (N_10206,N_9767,N_9279);
or U10207 (N_10207,N_9835,N_9680);
nand U10208 (N_10208,N_9157,N_9314);
nor U10209 (N_10209,N_9066,N_9760);
nor U10210 (N_10210,N_9932,N_9153);
and U10211 (N_10211,N_9448,N_9305);
nor U10212 (N_10212,N_9595,N_9938);
nand U10213 (N_10213,N_9889,N_9191);
and U10214 (N_10214,N_9287,N_9933);
nor U10215 (N_10215,N_9330,N_9338);
or U10216 (N_10216,N_9978,N_9182);
and U10217 (N_10217,N_9529,N_9037);
and U10218 (N_10218,N_9754,N_9750);
nor U10219 (N_10219,N_9829,N_9450);
nand U10220 (N_10220,N_9792,N_9820);
and U10221 (N_10221,N_9438,N_9297);
nand U10222 (N_10222,N_9538,N_9487);
nand U10223 (N_10223,N_9481,N_9201);
xor U10224 (N_10224,N_9834,N_9418);
nand U10225 (N_10225,N_9221,N_9358);
and U10226 (N_10226,N_9505,N_9653);
and U10227 (N_10227,N_9553,N_9036);
and U10228 (N_10228,N_9795,N_9982);
xnor U10229 (N_10229,N_9249,N_9381);
and U10230 (N_10230,N_9740,N_9407);
xnor U10231 (N_10231,N_9369,N_9917);
and U10232 (N_10232,N_9541,N_9666);
xnor U10233 (N_10233,N_9129,N_9038);
xor U10234 (N_10234,N_9027,N_9775);
xor U10235 (N_10235,N_9645,N_9142);
and U10236 (N_10236,N_9880,N_9171);
nand U10237 (N_10237,N_9458,N_9156);
xor U10238 (N_10238,N_9701,N_9200);
xnor U10239 (N_10239,N_9508,N_9856);
xor U10240 (N_10240,N_9076,N_9893);
xnor U10241 (N_10241,N_9040,N_9484);
and U10242 (N_10242,N_9205,N_9383);
nor U10243 (N_10243,N_9660,N_9814);
xnor U10244 (N_10244,N_9298,N_9154);
nor U10245 (N_10245,N_9721,N_9447);
xor U10246 (N_10246,N_9843,N_9203);
xnor U10247 (N_10247,N_9390,N_9703);
and U10248 (N_10248,N_9313,N_9285);
and U10249 (N_10249,N_9598,N_9340);
nor U10250 (N_10250,N_9083,N_9709);
xnor U10251 (N_10251,N_9518,N_9446);
xor U10252 (N_10252,N_9431,N_9710);
nand U10253 (N_10253,N_9261,N_9836);
xnor U10254 (N_10254,N_9098,N_9097);
nand U10255 (N_10255,N_9788,N_9683);
nor U10256 (N_10256,N_9397,N_9361);
or U10257 (N_10257,N_9198,N_9514);
and U10258 (N_10258,N_9270,N_9115);
nand U10259 (N_10259,N_9328,N_9539);
or U10260 (N_10260,N_9220,N_9561);
nor U10261 (N_10261,N_9454,N_9877);
nand U10262 (N_10262,N_9682,N_9739);
or U10263 (N_10263,N_9975,N_9993);
nor U10264 (N_10264,N_9863,N_9985);
or U10265 (N_10265,N_9827,N_9688);
or U10266 (N_10266,N_9124,N_9668);
or U10267 (N_10267,N_9729,N_9988);
xor U10268 (N_10268,N_9908,N_9226);
xnor U10269 (N_10269,N_9216,N_9542);
nand U10270 (N_10270,N_9266,N_9537);
or U10271 (N_10271,N_9655,N_9002);
or U10272 (N_10272,N_9011,N_9276);
or U10273 (N_10273,N_9331,N_9567);
and U10274 (N_10274,N_9056,N_9974);
and U10275 (N_10275,N_9079,N_9640);
and U10276 (N_10276,N_9209,N_9445);
nor U10277 (N_10277,N_9318,N_9425);
xor U10278 (N_10278,N_9671,N_9984);
and U10279 (N_10279,N_9695,N_9862);
xor U10280 (N_10280,N_9088,N_9786);
nor U10281 (N_10281,N_9506,N_9995);
xnor U10282 (N_10282,N_9465,N_9147);
nand U10283 (N_10283,N_9944,N_9798);
nor U10284 (N_10284,N_9696,N_9067);
xor U10285 (N_10285,N_9336,N_9503);
nor U10286 (N_10286,N_9842,N_9087);
nand U10287 (N_10287,N_9830,N_9939);
and U10288 (N_10288,N_9259,N_9632);
xnor U10289 (N_10289,N_9747,N_9152);
nand U10290 (N_10290,N_9262,N_9606);
nand U10291 (N_10291,N_9292,N_9497);
nor U10292 (N_10292,N_9189,N_9049);
xnor U10293 (N_10293,N_9386,N_9777);
nand U10294 (N_10294,N_9192,N_9343);
xor U10295 (N_10295,N_9964,N_9546);
or U10296 (N_10296,N_9215,N_9020);
nand U10297 (N_10297,N_9753,N_9246);
nor U10298 (N_10298,N_9509,N_9690);
or U10299 (N_10299,N_9380,N_9790);
and U10300 (N_10300,N_9356,N_9355);
and U10301 (N_10301,N_9486,N_9865);
or U10302 (N_10302,N_9206,N_9265);
and U10303 (N_10303,N_9849,N_9488);
or U10304 (N_10304,N_9233,N_9886);
nor U10305 (N_10305,N_9948,N_9081);
or U10306 (N_10306,N_9902,N_9178);
and U10307 (N_10307,N_9499,N_9046);
nor U10308 (N_10308,N_9161,N_9449);
and U10309 (N_10309,N_9725,N_9656);
xnor U10310 (N_10310,N_9758,N_9084);
nand U10311 (N_10311,N_9122,N_9765);
or U10312 (N_10312,N_9940,N_9935);
and U10313 (N_10313,N_9986,N_9284);
xor U10314 (N_10314,N_9222,N_9809);
nor U10315 (N_10315,N_9091,N_9007);
nor U10316 (N_10316,N_9973,N_9698);
xor U10317 (N_10317,N_9093,N_9582);
and U10318 (N_10318,N_9296,N_9914);
and U10319 (N_10319,N_9797,N_9457);
or U10320 (N_10320,N_9014,N_9125);
nand U10321 (N_10321,N_9323,N_9823);
xnor U10322 (N_10322,N_9955,N_9583);
or U10323 (N_10323,N_9891,N_9764);
or U10324 (N_10324,N_9600,N_9131);
and U10325 (N_10325,N_9565,N_9337);
xor U10326 (N_10326,N_9149,N_9267);
nor U10327 (N_10327,N_9364,N_9540);
or U10328 (N_10328,N_9114,N_9641);
or U10329 (N_10329,N_9210,N_9781);
nand U10330 (N_10330,N_9861,N_9111);
xor U10331 (N_10331,N_9410,N_9715);
nor U10332 (N_10332,N_9051,N_9851);
nor U10333 (N_10333,N_9981,N_9225);
xor U10334 (N_10334,N_9408,N_9793);
or U10335 (N_10335,N_9575,N_9490);
xor U10336 (N_10336,N_9648,N_9428);
nor U10337 (N_10337,N_9227,N_9647);
xnor U10338 (N_10338,N_9819,N_9983);
nand U10339 (N_10339,N_9931,N_9350);
and U10340 (N_10340,N_9733,N_9022);
nand U10341 (N_10341,N_9363,N_9116);
nand U10342 (N_10342,N_9654,N_9145);
nor U10343 (N_10343,N_9047,N_9315);
nand U10344 (N_10344,N_9252,N_9919);
nand U10345 (N_10345,N_9260,N_9839);
nor U10346 (N_10346,N_9961,N_9874);
nor U10347 (N_10347,N_9900,N_9167);
or U10348 (N_10348,N_9496,N_9610);
nor U10349 (N_10349,N_9597,N_9103);
nand U10350 (N_10350,N_9962,N_9008);
nand U10351 (N_10351,N_9400,N_9559);
nor U10352 (N_10352,N_9132,N_9674);
xnor U10353 (N_10353,N_9859,N_9631);
and U10354 (N_10354,N_9374,N_9126);
nor U10355 (N_10355,N_9847,N_9663);
or U10356 (N_10356,N_9462,N_9888);
nor U10357 (N_10357,N_9174,N_9556);
nand U10358 (N_10358,N_9395,N_9248);
nor U10359 (N_10359,N_9547,N_9780);
and U10360 (N_10360,N_9442,N_9642);
xnor U10361 (N_10361,N_9722,N_9420);
or U10362 (N_10362,N_9005,N_9905);
and U10363 (N_10363,N_9212,N_9043);
and U10364 (N_10364,N_9039,N_9526);
nor U10365 (N_10365,N_9619,N_9977);
or U10366 (N_10366,N_9176,N_9782);
or U10367 (N_10367,N_9090,N_9904);
xor U10368 (N_10368,N_9370,N_9882);
nand U10369 (N_10369,N_9708,N_9239);
nand U10370 (N_10370,N_9309,N_9879);
and U10371 (N_10371,N_9144,N_9244);
nand U10372 (N_10372,N_9624,N_9996);
nor U10373 (N_10373,N_9204,N_9500);
nor U10374 (N_10374,N_9120,N_9956);
and U10375 (N_10375,N_9398,N_9694);
xnor U10376 (N_10376,N_9063,N_9730);
and U10377 (N_10377,N_9432,N_9909);
nor U10378 (N_10378,N_9012,N_9927);
and U10379 (N_10379,N_9762,N_9558);
xnor U10380 (N_10380,N_9218,N_9082);
and U10381 (N_10381,N_9517,N_9492);
and U10382 (N_10382,N_9826,N_9303);
xor U10383 (N_10383,N_9522,N_9010);
or U10384 (N_10384,N_9277,N_9687);
xnor U10385 (N_10385,N_9810,N_9884);
nand U10386 (N_10386,N_9717,N_9247);
and U10387 (N_10387,N_9180,N_9853);
or U10388 (N_10388,N_9118,N_9563);
and U10389 (N_10389,N_9622,N_9633);
nand U10390 (N_10390,N_9644,N_9175);
or U10391 (N_10391,N_9106,N_9134);
nor U10392 (N_10392,N_9924,N_9749);
xor U10393 (N_10393,N_9444,N_9544);
nor U10394 (N_10394,N_9269,N_9637);
nand U10395 (N_10395,N_9406,N_9623);
xnor U10396 (N_10396,N_9521,N_9421);
nor U10397 (N_10397,N_9852,N_9173);
and U10398 (N_10398,N_9473,N_9815);
and U10399 (N_10399,N_9639,N_9635);
xnor U10400 (N_10400,N_9327,N_9901);
xor U10401 (N_10401,N_9130,N_9592);
nand U10402 (N_10402,N_9772,N_9104);
nor U10403 (N_10403,N_9569,N_9579);
and U10404 (N_10404,N_9976,N_9997);
or U10405 (N_10405,N_9493,N_9168);
nand U10406 (N_10406,N_9143,N_9301);
nor U10407 (N_10407,N_9573,N_9456);
xnor U10408 (N_10408,N_9136,N_9947);
or U10409 (N_10409,N_9094,N_9302);
xnor U10410 (N_10410,N_9669,N_9778);
nor U10411 (N_10411,N_9594,N_9785);
or U10412 (N_10412,N_9958,N_9604);
or U10413 (N_10413,N_9857,N_9375);
nor U10414 (N_10414,N_9560,N_9479);
nand U10415 (N_10415,N_9716,N_9896);
and U10416 (N_10416,N_9755,N_9440);
and U10417 (N_10417,N_9480,N_9288);
or U10418 (N_10418,N_9531,N_9878);
or U10419 (N_10419,N_9159,N_9348);
xnor U10420 (N_10420,N_9214,N_9650);
nand U10421 (N_10421,N_9382,N_9912);
and U10422 (N_10422,N_9436,N_9536);
nand U10423 (N_10423,N_9068,N_9427);
xnor U10424 (N_10424,N_9095,N_9415);
nor U10425 (N_10425,N_9378,N_9920);
and U10426 (N_10426,N_9881,N_9112);
and U10427 (N_10427,N_9992,N_9519);
nand U10428 (N_10428,N_9591,N_9367);
nor U10429 (N_10429,N_9937,N_9887);
and U10430 (N_10430,N_9564,N_9139);
xor U10431 (N_10431,N_9268,N_9333);
nand U10432 (N_10432,N_9831,N_9803);
nor U10433 (N_10433,N_9160,N_9254);
nor U10434 (N_10434,N_9437,N_9075);
and U10435 (N_10435,N_9727,N_9670);
xor U10436 (N_10436,N_9615,N_9510);
and U10437 (N_10437,N_9485,N_9704);
and U10438 (N_10438,N_9726,N_9373);
nand U10439 (N_10439,N_9707,N_9577);
or U10440 (N_10440,N_9611,N_9028);
nand U10441 (N_10441,N_9805,N_9700);
and U10442 (N_10442,N_9608,N_9033);
xor U10443 (N_10443,N_9697,N_9922);
xnor U10444 (N_10444,N_9825,N_9368);
and U10445 (N_10445,N_9078,N_9769);
nor U10446 (N_10446,N_9678,N_9017);
or U10447 (N_10447,N_9692,N_9811);
or U10448 (N_10448,N_9527,N_9549);
xor U10449 (N_10449,N_9403,N_9545);
and U10450 (N_10450,N_9416,N_9256);
or U10451 (N_10451,N_9629,N_9757);
and U10452 (N_10452,N_9599,N_9016);
xnor U10453 (N_10453,N_9474,N_9468);
nor U10454 (N_10454,N_9673,N_9686);
or U10455 (N_10455,N_9217,N_9745);
nand U10456 (N_10456,N_9980,N_9872);
or U10457 (N_10457,N_9453,N_9032);
nand U10458 (N_10458,N_9101,N_9137);
nand U10459 (N_10459,N_9968,N_9946);
or U10460 (N_10460,N_9004,N_9960);
nor U10461 (N_10461,N_9443,N_9620);
nor U10462 (N_10462,N_9550,N_9024);
or U10463 (N_10463,N_9308,N_9534);
or U10464 (N_10464,N_9812,N_9050);
or U10465 (N_10465,N_9590,N_9470);
or U10466 (N_10466,N_9170,N_9568);
nor U10467 (N_10467,N_9822,N_9290);
or U10468 (N_10468,N_9251,N_9491);
or U10469 (N_10469,N_9138,N_9146);
xor U10470 (N_10470,N_9586,N_9821);
xnor U10471 (N_10471,N_9513,N_9310);
nor U10472 (N_10472,N_9242,N_9392);
nand U10473 (N_10473,N_9845,N_9646);
nor U10474 (N_10474,N_9439,N_9928);
xnor U10475 (N_10475,N_9951,N_9744);
nor U10476 (N_10476,N_9166,N_9833);
xor U10477 (N_10477,N_9376,N_9074);
and U10478 (N_10478,N_9941,N_9071);
nor U10479 (N_10479,N_9713,N_9969);
nand U10480 (N_10480,N_9489,N_9987);
xor U10481 (N_10481,N_9441,N_9041);
nor U10482 (N_10482,N_9148,N_9643);
or U10483 (N_10483,N_9763,N_9520);
nand U10484 (N_10484,N_9107,N_9061);
xor U10485 (N_10485,N_9728,N_9970);
and U10486 (N_10486,N_9965,N_9603);
or U10487 (N_10487,N_9354,N_9807);
nor U10488 (N_10488,N_9770,N_9841);
xnor U10489 (N_10489,N_9789,N_9942);
or U10490 (N_10490,N_9404,N_9866);
nor U10491 (N_10491,N_9229,N_9059);
nor U10492 (N_10492,N_9801,N_9072);
and U10493 (N_10493,N_9875,N_9918);
or U10494 (N_10494,N_9828,N_9926);
xnor U10495 (N_10495,N_9495,N_9417);
nor U10496 (N_10496,N_9898,N_9899);
nor U10497 (N_10497,N_9512,N_9870);
or U10498 (N_10498,N_9224,N_9844);
nand U10499 (N_10499,N_9511,N_9689);
or U10500 (N_10500,N_9286,N_9502);
and U10501 (N_10501,N_9919,N_9992);
nand U10502 (N_10502,N_9383,N_9744);
and U10503 (N_10503,N_9700,N_9755);
xor U10504 (N_10504,N_9917,N_9227);
nand U10505 (N_10505,N_9111,N_9586);
or U10506 (N_10506,N_9740,N_9052);
nor U10507 (N_10507,N_9353,N_9315);
and U10508 (N_10508,N_9235,N_9924);
xor U10509 (N_10509,N_9538,N_9650);
xor U10510 (N_10510,N_9702,N_9934);
or U10511 (N_10511,N_9614,N_9039);
and U10512 (N_10512,N_9012,N_9633);
nand U10513 (N_10513,N_9661,N_9364);
nand U10514 (N_10514,N_9957,N_9427);
or U10515 (N_10515,N_9554,N_9157);
xor U10516 (N_10516,N_9384,N_9647);
nor U10517 (N_10517,N_9479,N_9504);
or U10518 (N_10518,N_9876,N_9094);
xor U10519 (N_10519,N_9686,N_9456);
or U10520 (N_10520,N_9132,N_9078);
and U10521 (N_10521,N_9995,N_9284);
xor U10522 (N_10522,N_9312,N_9819);
or U10523 (N_10523,N_9762,N_9014);
or U10524 (N_10524,N_9939,N_9086);
or U10525 (N_10525,N_9799,N_9033);
nand U10526 (N_10526,N_9059,N_9941);
nor U10527 (N_10527,N_9937,N_9311);
xnor U10528 (N_10528,N_9043,N_9053);
and U10529 (N_10529,N_9870,N_9531);
and U10530 (N_10530,N_9372,N_9395);
nor U10531 (N_10531,N_9358,N_9604);
or U10532 (N_10532,N_9326,N_9504);
nor U10533 (N_10533,N_9453,N_9495);
and U10534 (N_10534,N_9034,N_9429);
xor U10535 (N_10535,N_9721,N_9860);
nor U10536 (N_10536,N_9651,N_9926);
or U10537 (N_10537,N_9491,N_9242);
xor U10538 (N_10538,N_9842,N_9155);
xor U10539 (N_10539,N_9196,N_9849);
or U10540 (N_10540,N_9134,N_9787);
nand U10541 (N_10541,N_9969,N_9493);
xnor U10542 (N_10542,N_9760,N_9206);
or U10543 (N_10543,N_9456,N_9589);
nor U10544 (N_10544,N_9161,N_9483);
nor U10545 (N_10545,N_9432,N_9266);
nor U10546 (N_10546,N_9621,N_9142);
nand U10547 (N_10547,N_9826,N_9976);
nor U10548 (N_10548,N_9236,N_9128);
nor U10549 (N_10549,N_9895,N_9333);
nand U10550 (N_10550,N_9436,N_9440);
nor U10551 (N_10551,N_9297,N_9704);
and U10552 (N_10552,N_9552,N_9788);
nor U10553 (N_10553,N_9432,N_9466);
and U10554 (N_10554,N_9870,N_9213);
nand U10555 (N_10555,N_9491,N_9714);
and U10556 (N_10556,N_9960,N_9117);
nor U10557 (N_10557,N_9671,N_9699);
xor U10558 (N_10558,N_9899,N_9877);
and U10559 (N_10559,N_9554,N_9655);
xnor U10560 (N_10560,N_9618,N_9620);
and U10561 (N_10561,N_9082,N_9949);
or U10562 (N_10562,N_9180,N_9515);
and U10563 (N_10563,N_9089,N_9539);
nor U10564 (N_10564,N_9007,N_9343);
nand U10565 (N_10565,N_9554,N_9134);
xor U10566 (N_10566,N_9970,N_9832);
xnor U10567 (N_10567,N_9621,N_9555);
nand U10568 (N_10568,N_9158,N_9390);
and U10569 (N_10569,N_9455,N_9601);
nor U10570 (N_10570,N_9096,N_9753);
or U10571 (N_10571,N_9835,N_9927);
nand U10572 (N_10572,N_9709,N_9680);
nor U10573 (N_10573,N_9845,N_9634);
nor U10574 (N_10574,N_9862,N_9774);
xor U10575 (N_10575,N_9920,N_9861);
xor U10576 (N_10576,N_9891,N_9138);
nor U10577 (N_10577,N_9274,N_9984);
nand U10578 (N_10578,N_9607,N_9969);
nor U10579 (N_10579,N_9718,N_9852);
or U10580 (N_10580,N_9714,N_9664);
and U10581 (N_10581,N_9499,N_9395);
nor U10582 (N_10582,N_9413,N_9191);
xor U10583 (N_10583,N_9513,N_9899);
nand U10584 (N_10584,N_9334,N_9451);
nor U10585 (N_10585,N_9951,N_9406);
or U10586 (N_10586,N_9466,N_9827);
or U10587 (N_10587,N_9807,N_9114);
xnor U10588 (N_10588,N_9413,N_9458);
xnor U10589 (N_10589,N_9530,N_9065);
xnor U10590 (N_10590,N_9188,N_9087);
or U10591 (N_10591,N_9612,N_9636);
nor U10592 (N_10592,N_9288,N_9462);
or U10593 (N_10593,N_9758,N_9439);
xor U10594 (N_10594,N_9813,N_9432);
or U10595 (N_10595,N_9545,N_9443);
xnor U10596 (N_10596,N_9231,N_9509);
xor U10597 (N_10597,N_9148,N_9446);
nand U10598 (N_10598,N_9122,N_9693);
nand U10599 (N_10599,N_9616,N_9615);
or U10600 (N_10600,N_9789,N_9001);
nor U10601 (N_10601,N_9221,N_9092);
and U10602 (N_10602,N_9927,N_9431);
nand U10603 (N_10603,N_9114,N_9332);
or U10604 (N_10604,N_9081,N_9825);
and U10605 (N_10605,N_9341,N_9623);
nor U10606 (N_10606,N_9697,N_9190);
or U10607 (N_10607,N_9029,N_9935);
nand U10608 (N_10608,N_9502,N_9084);
xnor U10609 (N_10609,N_9500,N_9269);
or U10610 (N_10610,N_9543,N_9133);
nor U10611 (N_10611,N_9870,N_9346);
and U10612 (N_10612,N_9120,N_9564);
xnor U10613 (N_10613,N_9600,N_9146);
and U10614 (N_10614,N_9350,N_9247);
nor U10615 (N_10615,N_9059,N_9232);
xor U10616 (N_10616,N_9762,N_9097);
or U10617 (N_10617,N_9815,N_9017);
or U10618 (N_10618,N_9655,N_9596);
xnor U10619 (N_10619,N_9908,N_9629);
nor U10620 (N_10620,N_9919,N_9679);
and U10621 (N_10621,N_9633,N_9232);
or U10622 (N_10622,N_9773,N_9905);
nor U10623 (N_10623,N_9428,N_9069);
nand U10624 (N_10624,N_9961,N_9211);
and U10625 (N_10625,N_9123,N_9317);
nand U10626 (N_10626,N_9831,N_9421);
and U10627 (N_10627,N_9495,N_9484);
nor U10628 (N_10628,N_9299,N_9325);
and U10629 (N_10629,N_9106,N_9836);
xnor U10630 (N_10630,N_9993,N_9845);
nand U10631 (N_10631,N_9710,N_9536);
nand U10632 (N_10632,N_9291,N_9683);
nand U10633 (N_10633,N_9009,N_9668);
and U10634 (N_10634,N_9381,N_9995);
or U10635 (N_10635,N_9014,N_9791);
nand U10636 (N_10636,N_9448,N_9650);
and U10637 (N_10637,N_9011,N_9895);
nor U10638 (N_10638,N_9925,N_9814);
or U10639 (N_10639,N_9832,N_9256);
nand U10640 (N_10640,N_9115,N_9523);
nand U10641 (N_10641,N_9552,N_9111);
and U10642 (N_10642,N_9590,N_9529);
or U10643 (N_10643,N_9751,N_9123);
xnor U10644 (N_10644,N_9328,N_9527);
nand U10645 (N_10645,N_9505,N_9957);
nor U10646 (N_10646,N_9573,N_9590);
nor U10647 (N_10647,N_9922,N_9160);
and U10648 (N_10648,N_9486,N_9991);
and U10649 (N_10649,N_9163,N_9802);
nand U10650 (N_10650,N_9357,N_9725);
xnor U10651 (N_10651,N_9568,N_9043);
or U10652 (N_10652,N_9231,N_9552);
or U10653 (N_10653,N_9351,N_9556);
or U10654 (N_10654,N_9121,N_9375);
nor U10655 (N_10655,N_9811,N_9317);
and U10656 (N_10656,N_9514,N_9315);
or U10657 (N_10657,N_9313,N_9098);
nand U10658 (N_10658,N_9800,N_9907);
nor U10659 (N_10659,N_9504,N_9149);
nand U10660 (N_10660,N_9331,N_9055);
or U10661 (N_10661,N_9425,N_9874);
and U10662 (N_10662,N_9507,N_9301);
nand U10663 (N_10663,N_9020,N_9336);
and U10664 (N_10664,N_9995,N_9749);
nand U10665 (N_10665,N_9517,N_9190);
nand U10666 (N_10666,N_9226,N_9336);
and U10667 (N_10667,N_9186,N_9817);
or U10668 (N_10668,N_9238,N_9347);
and U10669 (N_10669,N_9605,N_9401);
nor U10670 (N_10670,N_9519,N_9605);
nor U10671 (N_10671,N_9288,N_9964);
nor U10672 (N_10672,N_9310,N_9623);
or U10673 (N_10673,N_9638,N_9342);
xnor U10674 (N_10674,N_9658,N_9164);
xnor U10675 (N_10675,N_9765,N_9902);
and U10676 (N_10676,N_9534,N_9959);
or U10677 (N_10677,N_9539,N_9514);
nand U10678 (N_10678,N_9685,N_9452);
nand U10679 (N_10679,N_9909,N_9030);
xor U10680 (N_10680,N_9958,N_9693);
or U10681 (N_10681,N_9177,N_9676);
nand U10682 (N_10682,N_9227,N_9188);
or U10683 (N_10683,N_9215,N_9927);
and U10684 (N_10684,N_9530,N_9471);
and U10685 (N_10685,N_9757,N_9438);
nand U10686 (N_10686,N_9420,N_9559);
xnor U10687 (N_10687,N_9428,N_9597);
xor U10688 (N_10688,N_9018,N_9783);
nand U10689 (N_10689,N_9978,N_9823);
xor U10690 (N_10690,N_9337,N_9953);
nand U10691 (N_10691,N_9517,N_9113);
or U10692 (N_10692,N_9762,N_9094);
nor U10693 (N_10693,N_9781,N_9835);
nand U10694 (N_10694,N_9790,N_9296);
xor U10695 (N_10695,N_9925,N_9471);
and U10696 (N_10696,N_9018,N_9522);
nand U10697 (N_10697,N_9725,N_9543);
nand U10698 (N_10698,N_9773,N_9545);
xor U10699 (N_10699,N_9743,N_9533);
nor U10700 (N_10700,N_9871,N_9085);
nand U10701 (N_10701,N_9230,N_9668);
nand U10702 (N_10702,N_9798,N_9834);
and U10703 (N_10703,N_9758,N_9405);
nor U10704 (N_10704,N_9525,N_9558);
nand U10705 (N_10705,N_9914,N_9927);
xnor U10706 (N_10706,N_9338,N_9561);
nor U10707 (N_10707,N_9378,N_9352);
or U10708 (N_10708,N_9835,N_9789);
and U10709 (N_10709,N_9244,N_9185);
nand U10710 (N_10710,N_9173,N_9232);
nor U10711 (N_10711,N_9435,N_9313);
xor U10712 (N_10712,N_9272,N_9386);
or U10713 (N_10713,N_9213,N_9847);
and U10714 (N_10714,N_9258,N_9968);
xor U10715 (N_10715,N_9884,N_9659);
and U10716 (N_10716,N_9697,N_9756);
xnor U10717 (N_10717,N_9851,N_9143);
or U10718 (N_10718,N_9474,N_9769);
nand U10719 (N_10719,N_9765,N_9476);
xor U10720 (N_10720,N_9023,N_9224);
nand U10721 (N_10721,N_9180,N_9203);
nand U10722 (N_10722,N_9914,N_9688);
nor U10723 (N_10723,N_9328,N_9012);
nor U10724 (N_10724,N_9257,N_9978);
xor U10725 (N_10725,N_9247,N_9609);
xor U10726 (N_10726,N_9962,N_9168);
nor U10727 (N_10727,N_9434,N_9695);
or U10728 (N_10728,N_9910,N_9511);
or U10729 (N_10729,N_9505,N_9794);
nor U10730 (N_10730,N_9544,N_9758);
nor U10731 (N_10731,N_9144,N_9155);
or U10732 (N_10732,N_9077,N_9127);
nand U10733 (N_10733,N_9458,N_9153);
nand U10734 (N_10734,N_9284,N_9338);
and U10735 (N_10735,N_9503,N_9580);
and U10736 (N_10736,N_9384,N_9142);
or U10737 (N_10737,N_9125,N_9141);
or U10738 (N_10738,N_9829,N_9906);
or U10739 (N_10739,N_9517,N_9144);
or U10740 (N_10740,N_9929,N_9036);
and U10741 (N_10741,N_9664,N_9472);
nand U10742 (N_10742,N_9460,N_9098);
and U10743 (N_10743,N_9925,N_9678);
or U10744 (N_10744,N_9142,N_9241);
or U10745 (N_10745,N_9725,N_9413);
nand U10746 (N_10746,N_9066,N_9047);
or U10747 (N_10747,N_9467,N_9772);
xnor U10748 (N_10748,N_9884,N_9452);
nand U10749 (N_10749,N_9939,N_9746);
xnor U10750 (N_10750,N_9656,N_9361);
or U10751 (N_10751,N_9091,N_9372);
nand U10752 (N_10752,N_9036,N_9025);
nor U10753 (N_10753,N_9710,N_9482);
or U10754 (N_10754,N_9405,N_9320);
xor U10755 (N_10755,N_9730,N_9639);
and U10756 (N_10756,N_9090,N_9624);
and U10757 (N_10757,N_9971,N_9384);
nand U10758 (N_10758,N_9229,N_9672);
nand U10759 (N_10759,N_9561,N_9209);
or U10760 (N_10760,N_9059,N_9227);
and U10761 (N_10761,N_9780,N_9424);
nor U10762 (N_10762,N_9209,N_9088);
xnor U10763 (N_10763,N_9021,N_9756);
nor U10764 (N_10764,N_9599,N_9120);
and U10765 (N_10765,N_9572,N_9886);
xor U10766 (N_10766,N_9450,N_9070);
and U10767 (N_10767,N_9714,N_9030);
nor U10768 (N_10768,N_9490,N_9764);
or U10769 (N_10769,N_9227,N_9782);
nor U10770 (N_10770,N_9493,N_9609);
or U10771 (N_10771,N_9081,N_9468);
nor U10772 (N_10772,N_9373,N_9387);
and U10773 (N_10773,N_9457,N_9180);
nor U10774 (N_10774,N_9920,N_9421);
nor U10775 (N_10775,N_9818,N_9781);
and U10776 (N_10776,N_9562,N_9465);
xor U10777 (N_10777,N_9931,N_9668);
nand U10778 (N_10778,N_9329,N_9668);
xnor U10779 (N_10779,N_9284,N_9324);
and U10780 (N_10780,N_9277,N_9187);
and U10781 (N_10781,N_9591,N_9455);
nor U10782 (N_10782,N_9569,N_9564);
nand U10783 (N_10783,N_9350,N_9869);
or U10784 (N_10784,N_9198,N_9819);
nand U10785 (N_10785,N_9804,N_9826);
nand U10786 (N_10786,N_9953,N_9986);
nor U10787 (N_10787,N_9725,N_9174);
xnor U10788 (N_10788,N_9467,N_9108);
nand U10789 (N_10789,N_9698,N_9107);
nand U10790 (N_10790,N_9326,N_9207);
and U10791 (N_10791,N_9100,N_9697);
nor U10792 (N_10792,N_9663,N_9493);
or U10793 (N_10793,N_9984,N_9929);
and U10794 (N_10794,N_9940,N_9071);
xnor U10795 (N_10795,N_9852,N_9621);
or U10796 (N_10796,N_9110,N_9199);
and U10797 (N_10797,N_9638,N_9837);
nand U10798 (N_10798,N_9956,N_9579);
or U10799 (N_10799,N_9780,N_9787);
xnor U10800 (N_10800,N_9435,N_9286);
and U10801 (N_10801,N_9201,N_9290);
nor U10802 (N_10802,N_9254,N_9123);
and U10803 (N_10803,N_9931,N_9448);
or U10804 (N_10804,N_9964,N_9576);
or U10805 (N_10805,N_9416,N_9388);
and U10806 (N_10806,N_9176,N_9876);
and U10807 (N_10807,N_9297,N_9504);
nand U10808 (N_10808,N_9892,N_9777);
or U10809 (N_10809,N_9013,N_9041);
and U10810 (N_10810,N_9192,N_9338);
and U10811 (N_10811,N_9690,N_9137);
and U10812 (N_10812,N_9141,N_9972);
nor U10813 (N_10813,N_9029,N_9220);
or U10814 (N_10814,N_9451,N_9262);
or U10815 (N_10815,N_9606,N_9862);
nand U10816 (N_10816,N_9138,N_9078);
or U10817 (N_10817,N_9540,N_9635);
or U10818 (N_10818,N_9154,N_9771);
and U10819 (N_10819,N_9934,N_9402);
nor U10820 (N_10820,N_9688,N_9292);
xnor U10821 (N_10821,N_9025,N_9848);
xnor U10822 (N_10822,N_9727,N_9712);
xnor U10823 (N_10823,N_9511,N_9063);
or U10824 (N_10824,N_9137,N_9493);
nor U10825 (N_10825,N_9402,N_9799);
nand U10826 (N_10826,N_9663,N_9553);
nor U10827 (N_10827,N_9701,N_9634);
and U10828 (N_10828,N_9300,N_9540);
xor U10829 (N_10829,N_9946,N_9260);
nor U10830 (N_10830,N_9154,N_9260);
and U10831 (N_10831,N_9034,N_9137);
nand U10832 (N_10832,N_9540,N_9189);
or U10833 (N_10833,N_9125,N_9458);
nand U10834 (N_10834,N_9807,N_9563);
nor U10835 (N_10835,N_9545,N_9549);
or U10836 (N_10836,N_9194,N_9771);
and U10837 (N_10837,N_9288,N_9229);
or U10838 (N_10838,N_9885,N_9193);
or U10839 (N_10839,N_9830,N_9115);
or U10840 (N_10840,N_9300,N_9326);
nand U10841 (N_10841,N_9830,N_9196);
or U10842 (N_10842,N_9549,N_9060);
xor U10843 (N_10843,N_9072,N_9531);
nand U10844 (N_10844,N_9550,N_9770);
and U10845 (N_10845,N_9342,N_9663);
nor U10846 (N_10846,N_9524,N_9541);
or U10847 (N_10847,N_9910,N_9537);
nor U10848 (N_10848,N_9108,N_9640);
or U10849 (N_10849,N_9033,N_9040);
nand U10850 (N_10850,N_9348,N_9884);
and U10851 (N_10851,N_9837,N_9391);
or U10852 (N_10852,N_9909,N_9203);
xor U10853 (N_10853,N_9701,N_9962);
or U10854 (N_10854,N_9921,N_9122);
xnor U10855 (N_10855,N_9508,N_9940);
xor U10856 (N_10856,N_9648,N_9449);
nor U10857 (N_10857,N_9607,N_9310);
and U10858 (N_10858,N_9441,N_9377);
xnor U10859 (N_10859,N_9920,N_9910);
and U10860 (N_10860,N_9424,N_9790);
xor U10861 (N_10861,N_9952,N_9923);
nand U10862 (N_10862,N_9116,N_9876);
nor U10863 (N_10863,N_9258,N_9528);
and U10864 (N_10864,N_9119,N_9510);
or U10865 (N_10865,N_9037,N_9036);
nor U10866 (N_10866,N_9255,N_9392);
nor U10867 (N_10867,N_9058,N_9580);
and U10868 (N_10868,N_9580,N_9007);
nand U10869 (N_10869,N_9773,N_9494);
or U10870 (N_10870,N_9971,N_9707);
nand U10871 (N_10871,N_9959,N_9899);
or U10872 (N_10872,N_9579,N_9214);
nand U10873 (N_10873,N_9710,N_9091);
nor U10874 (N_10874,N_9222,N_9868);
and U10875 (N_10875,N_9363,N_9142);
or U10876 (N_10876,N_9172,N_9645);
and U10877 (N_10877,N_9548,N_9298);
nand U10878 (N_10878,N_9447,N_9133);
and U10879 (N_10879,N_9228,N_9413);
or U10880 (N_10880,N_9386,N_9514);
or U10881 (N_10881,N_9074,N_9747);
nor U10882 (N_10882,N_9256,N_9730);
or U10883 (N_10883,N_9774,N_9259);
nor U10884 (N_10884,N_9193,N_9849);
or U10885 (N_10885,N_9837,N_9644);
nand U10886 (N_10886,N_9550,N_9913);
and U10887 (N_10887,N_9418,N_9875);
and U10888 (N_10888,N_9960,N_9439);
nor U10889 (N_10889,N_9628,N_9362);
xnor U10890 (N_10890,N_9367,N_9295);
nor U10891 (N_10891,N_9711,N_9528);
or U10892 (N_10892,N_9860,N_9178);
and U10893 (N_10893,N_9767,N_9087);
nor U10894 (N_10894,N_9914,N_9032);
or U10895 (N_10895,N_9839,N_9476);
and U10896 (N_10896,N_9438,N_9322);
xnor U10897 (N_10897,N_9710,N_9309);
and U10898 (N_10898,N_9740,N_9567);
nor U10899 (N_10899,N_9622,N_9812);
or U10900 (N_10900,N_9830,N_9357);
nor U10901 (N_10901,N_9514,N_9732);
and U10902 (N_10902,N_9110,N_9796);
nor U10903 (N_10903,N_9132,N_9852);
or U10904 (N_10904,N_9080,N_9767);
nand U10905 (N_10905,N_9438,N_9992);
xor U10906 (N_10906,N_9979,N_9440);
nor U10907 (N_10907,N_9676,N_9699);
and U10908 (N_10908,N_9445,N_9561);
xor U10909 (N_10909,N_9984,N_9256);
and U10910 (N_10910,N_9925,N_9545);
and U10911 (N_10911,N_9255,N_9162);
or U10912 (N_10912,N_9477,N_9482);
xnor U10913 (N_10913,N_9722,N_9541);
and U10914 (N_10914,N_9537,N_9650);
or U10915 (N_10915,N_9556,N_9704);
or U10916 (N_10916,N_9016,N_9197);
xnor U10917 (N_10917,N_9149,N_9320);
or U10918 (N_10918,N_9840,N_9084);
and U10919 (N_10919,N_9221,N_9308);
and U10920 (N_10920,N_9801,N_9721);
or U10921 (N_10921,N_9229,N_9853);
nand U10922 (N_10922,N_9450,N_9897);
nand U10923 (N_10923,N_9928,N_9374);
and U10924 (N_10924,N_9581,N_9112);
or U10925 (N_10925,N_9889,N_9003);
and U10926 (N_10926,N_9976,N_9269);
xor U10927 (N_10927,N_9087,N_9262);
xnor U10928 (N_10928,N_9930,N_9421);
or U10929 (N_10929,N_9635,N_9909);
or U10930 (N_10930,N_9201,N_9581);
and U10931 (N_10931,N_9472,N_9212);
nand U10932 (N_10932,N_9220,N_9843);
or U10933 (N_10933,N_9754,N_9663);
nor U10934 (N_10934,N_9047,N_9853);
or U10935 (N_10935,N_9164,N_9280);
nor U10936 (N_10936,N_9822,N_9089);
or U10937 (N_10937,N_9169,N_9932);
or U10938 (N_10938,N_9651,N_9894);
nand U10939 (N_10939,N_9877,N_9448);
nand U10940 (N_10940,N_9671,N_9376);
nor U10941 (N_10941,N_9441,N_9821);
or U10942 (N_10942,N_9522,N_9189);
and U10943 (N_10943,N_9663,N_9929);
and U10944 (N_10944,N_9260,N_9623);
or U10945 (N_10945,N_9527,N_9092);
or U10946 (N_10946,N_9632,N_9857);
xnor U10947 (N_10947,N_9789,N_9273);
and U10948 (N_10948,N_9795,N_9673);
xnor U10949 (N_10949,N_9362,N_9632);
nand U10950 (N_10950,N_9095,N_9234);
nand U10951 (N_10951,N_9744,N_9646);
or U10952 (N_10952,N_9790,N_9398);
nor U10953 (N_10953,N_9422,N_9146);
xnor U10954 (N_10954,N_9944,N_9377);
nor U10955 (N_10955,N_9619,N_9167);
nor U10956 (N_10956,N_9669,N_9950);
or U10957 (N_10957,N_9804,N_9415);
nor U10958 (N_10958,N_9486,N_9799);
nand U10959 (N_10959,N_9755,N_9919);
nor U10960 (N_10960,N_9443,N_9031);
and U10961 (N_10961,N_9838,N_9143);
nand U10962 (N_10962,N_9696,N_9076);
or U10963 (N_10963,N_9671,N_9747);
nand U10964 (N_10964,N_9704,N_9262);
nor U10965 (N_10965,N_9762,N_9602);
nor U10966 (N_10966,N_9895,N_9476);
and U10967 (N_10967,N_9391,N_9701);
and U10968 (N_10968,N_9624,N_9021);
nor U10969 (N_10969,N_9984,N_9169);
nand U10970 (N_10970,N_9380,N_9752);
or U10971 (N_10971,N_9155,N_9112);
nand U10972 (N_10972,N_9233,N_9456);
nand U10973 (N_10973,N_9516,N_9254);
xor U10974 (N_10974,N_9614,N_9843);
and U10975 (N_10975,N_9167,N_9946);
xnor U10976 (N_10976,N_9369,N_9746);
xor U10977 (N_10977,N_9383,N_9614);
nand U10978 (N_10978,N_9235,N_9154);
nor U10979 (N_10979,N_9837,N_9370);
nand U10980 (N_10980,N_9115,N_9639);
xor U10981 (N_10981,N_9449,N_9928);
or U10982 (N_10982,N_9676,N_9925);
nor U10983 (N_10983,N_9338,N_9018);
nand U10984 (N_10984,N_9172,N_9399);
nor U10985 (N_10985,N_9938,N_9721);
nor U10986 (N_10986,N_9745,N_9454);
and U10987 (N_10987,N_9166,N_9570);
or U10988 (N_10988,N_9920,N_9962);
xnor U10989 (N_10989,N_9140,N_9341);
or U10990 (N_10990,N_9004,N_9583);
nand U10991 (N_10991,N_9285,N_9907);
nor U10992 (N_10992,N_9736,N_9339);
and U10993 (N_10993,N_9898,N_9045);
nor U10994 (N_10994,N_9211,N_9883);
xor U10995 (N_10995,N_9610,N_9976);
and U10996 (N_10996,N_9007,N_9256);
nand U10997 (N_10997,N_9134,N_9835);
or U10998 (N_10998,N_9970,N_9039);
and U10999 (N_10999,N_9196,N_9627);
and U11000 (N_11000,N_10716,N_10649);
and U11001 (N_11001,N_10040,N_10950);
xnor U11002 (N_11002,N_10968,N_10852);
xor U11003 (N_11003,N_10883,N_10887);
nand U11004 (N_11004,N_10110,N_10564);
xnor U11005 (N_11005,N_10194,N_10869);
nand U11006 (N_11006,N_10168,N_10212);
or U11007 (N_11007,N_10135,N_10123);
and U11008 (N_11008,N_10332,N_10926);
nor U11009 (N_11009,N_10327,N_10560);
nand U11010 (N_11010,N_10092,N_10153);
xor U11011 (N_11011,N_10938,N_10744);
nor U11012 (N_11012,N_10970,N_10606);
nand U11013 (N_11013,N_10301,N_10009);
nand U11014 (N_11014,N_10389,N_10801);
xor U11015 (N_11015,N_10767,N_10066);
and U11016 (N_11016,N_10895,N_10988);
nor U11017 (N_11017,N_10300,N_10315);
and U11018 (N_11018,N_10520,N_10489);
or U11019 (N_11019,N_10287,N_10912);
nand U11020 (N_11020,N_10414,N_10838);
nor U11021 (N_11021,N_10139,N_10855);
and U11022 (N_11022,N_10458,N_10675);
xor U11023 (N_11023,N_10086,N_10863);
nand U11024 (N_11024,N_10395,N_10367);
nand U11025 (N_11025,N_10507,N_10992);
nor U11026 (N_11026,N_10751,N_10383);
nand U11027 (N_11027,N_10178,N_10755);
nand U11028 (N_11028,N_10486,N_10515);
nand U11029 (N_11029,N_10387,N_10888);
xnor U11030 (N_11030,N_10693,N_10686);
nor U11031 (N_11031,N_10371,N_10457);
xor U11032 (N_11032,N_10103,N_10236);
or U11033 (N_11033,N_10118,N_10575);
xor U11034 (N_11034,N_10243,N_10469);
or U11035 (N_11035,N_10430,N_10821);
nand U11036 (N_11036,N_10813,N_10282);
xnor U11037 (N_11037,N_10014,N_10891);
xor U11038 (N_11038,N_10095,N_10131);
nand U11039 (N_11039,N_10476,N_10002);
and U11040 (N_11040,N_10679,N_10845);
and U11041 (N_11041,N_10922,N_10714);
xnor U11042 (N_11042,N_10233,N_10292);
nand U11043 (N_11043,N_10244,N_10800);
and U11044 (N_11044,N_10842,N_10848);
or U11045 (N_11045,N_10406,N_10256);
nor U11046 (N_11046,N_10657,N_10816);
nor U11047 (N_11047,N_10288,N_10510);
nand U11048 (N_11048,N_10196,N_10592);
nand U11049 (N_11049,N_10474,N_10420);
and U11050 (N_11050,N_10382,N_10322);
nor U11051 (N_11051,N_10127,N_10843);
nand U11052 (N_11052,N_10145,N_10392);
xor U11053 (N_11053,N_10370,N_10728);
nand U11054 (N_11054,N_10147,N_10343);
xor U11055 (N_11055,N_10351,N_10302);
xnor U11056 (N_11056,N_10633,N_10769);
nor U11057 (N_11057,N_10772,N_10729);
and U11058 (N_11058,N_10811,N_10546);
or U11059 (N_11059,N_10273,N_10715);
and U11060 (N_11060,N_10830,N_10875);
and U11061 (N_11061,N_10849,N_10384);
or U11062 (N_11062,N_10834,N_10949);
xor U11063 (N_11063,N_10963,N_10815);
or U11064 (N_11064,N_10381,N_10920);
xor U11065 (N_11065,N_10219,N_10410);
nor U11066 (N_11066,N_10688,N_10033);
nor U11067 (N_11067,N_10019,N_10481);
xor U11068 (N_11068,N_10543,N_10905);
nor U11069 (N_11069,N_10077,N_10105);
xor U11070 (N_11070,N_10783,N_10579);
and U11071 (N_11071,N_10334,N_10513);
nand U11072 (N_11072,N_10622,N_10470);
or U11073 (N_11073,N_10156,N_10656);
or U11074 (N_11074,N_10578,N_10016);
nor U11075 (N_11075,N_10403,N_10449);
and U11076 (N_11076,N_10438,N_10943);
nand U11077 (N_11077,N_10150,N_10107);
xnor U11078 (N_11078,N_10043,N_10473);
xnor U11079 (N_11079,N_10494,N_10999);
or U11080 (N_11080,N_10415,N_10396);
nor U11081 (N_11081,N_10029,N_10166);
and U11082 (N_11082,N_10133,N_10789);
and U11083 (N_11083,N_10208,N_10443);
xnor U11084 (N_11084,N_10587,N_10251);
and U11085 (N_11085,N_10614,N_10278);
nand U11086 (N_11086,N_10659,N_10709);
or U11087 (N_11087,N_10246,N_10159);
and U11088 (N_11088,N_10788,N_10862);
xnor U11089 (N_11089,N_10076,N_10207);
or U11090 (N_11090,N_10252,N_10423);
or U11091 (N_11091,N_10625,N_10213);
nor U11092 (N_11092,N_10027,N_10448);
nor U11093 (N_11093,N_10065,N_10792);
nand U11094 (N_11094,N_10739,N_10655);
nor U11095 (N_11095,N_10761,N_10588);
nand U11096 (N_11096,N_10984,N_10765);
nor U11097 (N_11097,N_10202,N_10893);
nor U11098 (N_11098,N_10930,N_10031);
nand U11099 (N_11099,N_10941,N_10652);
and U11100 (N_11100,N_10480,N_10525);
xnor U11101 (N_11101,N_10336,N_10923);
xnor U11102 (N_11102,N_10931,N_10240);
nor U11103 (N_11103,N_10154,N_10768);
nor U11104 (N_11104,N_10230,N_10115);
nand U11105 (N_11105,N_10902,N_10871);
nand U11106 (N_11106,N_10827,N_10928);
xor U11107 (N_11107,N_10356,N_10824);
nand U11108 (N_11108,N_10733,N_10405);
xor U11109 (N_11109,N_10493,N_10121);
nand U11110 (N_11110,N_10089,N_10143);
and U11111 (N_11111,N_10508,N_10399);
xor U11112 (N_11112,N_10929,N_10964);
and U11113 (N_11113,N_10781,N_10333);
or U11114 (N_11114,N_10453,N_10619);
xnor U11115 (N_11115,N_10311,N_10994);
nor U11116 (N_11116,N_10646,N_10954);
or U11117 (N_11117,N_10390,N_10743);
or U11118 (N_11118,N_10264,N_10638);
and U11119 (N_11119,N_10960,N_10439);
nand U11120 (N_11120,N_10787,N_10726);
nand U11121 (N_11121,N_10348,N_10042);
and U11122 (N_11122,N_10102,N_10011);
or U11123 (N_11123,N_10257,N_10364);
xor U11124 (N_11124,N_10025,N_10354);
xnor U11125 (N_11125,N_10705,N_10548);
nor U11126 (N_11126,N_10155,N_10967);
nor U11127 (N_11127,N_10516,N_10184);
and U11128 (N_11128,N_10071,N_10250);
nand U11129 (N_11129,N_10283,N_10804);
or U11130 (N_11130,N_10959,N_10130);
or U11131 (N_11131,N_10010,N_10004);
nand U11132 (N_11132,N_10710,N_10023);
nor U11133 (N_11133,N_10366,N_10140);
nor U11134 (N_11134,N_10148,N_10098);
nand U11135 (N_11135,N_10122,N_10746);
xor U11136 (N_11136,N_10001,N_10707);
nand U11137 (N_11137,N_10083,N_10975);
nor U11138 (N_11138,N_10088,N_10426);
or U11139 (N_11139,N_10660,N_10175);
and U11140 (N_11140,N_10321,N_10731);
and U11141 (N_11141,N_10341,N_10756);
xnor U11142 (N_11142,N_10053,N_10497);
xor U11143 (N_11143,N_10262,N_10450);
nor U11144 (N_11144,N_10151,N_10590);
nand U11145 (N_11145,N_10719,N_10868);
nand U11146 (N_11146,N_10152,N_10277);
nand U11147 (N_11147,N_10199,N_10401);
xor U11148 (N_11148,N_10223,N_10683);
nor U11149 (N_11149,N_10198,N_10720);
and U11150 (N_11150,N_10472,N_10220);
nand U11151 (N_11151,N_10687,N_10078);
xor U11152 (N_11152,N_10442,N_10276);
or U11153 (N_11153,N_10445,N_10030);
or U11154 (N_11154,N_10512,N_10365);
and U11155 (N_11155,N_10253,N_10214);
and U11156 (N_11156,N_10907,N_10038);
and U11157 (N_11157,N_10499,N_10350);
xor U11158 (N_11158,N_10291,N_10627);
xnor U11159 (N_11159,N_10459,N_10226);
and U11160 (N_11160,N_10149,N_10850);
nand U11161 (N_11161,N_10722,N_10629);
nand U11162 (N_11162,N_10620,N_10081);
or U11163 (N_11163,N_10248,N_10164);
nor U11164 (N_11164,N_10643,N_10528);
or U11165 (N_11165,N_10460,N_10778);
xnor U11166 (N_11166,N_10313,N_10180);
nand U11167 (N_11167,N_10612,N_10829);
and U11168 (N_11168,N_10237,N_10752);
and U11169 (N_11169,N_10502,N_10073);
xor U11170 (N_11170,N_10036,N_10962);
nor U11171 (N_11171,N_10290,N_10980);
xnor U11172 (N_11172,N_10613,N_10634);
and U11173 (N_11173,N_10055,N_10573);
nand U11174 (N_11174,N_10070,N_10437);
and U11175 (N_11175,N_10805,N_10644);
nand U11176 (N_11176,N_10866,N_10757);
nor U11177 (N_11177,N_10203,N_10583);
xnor U11178 (N_11178,N_10097,N_10444);
nand U11179 (N_11179,N_10521,N_10044);
or U11180 (N_11180,N_10851,N_10295);
nor U11181 (N_11181,N_10305,N_10680);
or U11182 (N_11182,N_10340,N_10584);
and U11183 (N_11183,N_10440,N_10666);
or U11184 (N_11184,N_10385,N_10889);
xor U11185 (N_11185,N_10375,N_10872);
nor U11186 (N_11186,N_10903,N_10927);
and U11187 (N_11187,N_10839,N_10758);
nand U11188 (N_11188,N_10617,N_10279);
xor U11189 (N_11189,N_10640,N_10774);
nor U11190 (N_11190,N_10704,N_10242);
nor U11191 (N_11191,N_10455,N_10897);
nor U11192 (N_11192,N_10116,N_10581);
nand U11193 (N_11193,N_10338,N_10732);
and U11194 (N_11194,N_10873,N_10079);
nor U11195 (N_11195,N_10298,N_10369);
nand U11196 (N_11196,N_10221,N_10607);
or U11197 (N_11197,N_10478,N_10012);
nor U11198 (N_11198,N_10550,N_10120);
or U11199 (N_11199,N_10809,N_10518);
and U11200 (N_11200,N_10008,N_10361);
nand U11201 (N_11201,N_10645,N_10067);
nand U11202 (N_11202,N_10328,N_10621);
and U11203 (N_11203,N_10776,N_10063);
or U11204 (N_11204,N_10536,N_10712);
xnor U11205 (N_11205,N_10421,N_10393);
and U11206 (N_11206,N_10183,N_10847);
xnor U11207 (N_11207,N_10346,N_10270);
nor U11208 (N_11208,N_10635,N_10671);
nand U11209 (N_11209,N_10072,N_10228);
nand U11210 (N_11210,N_10754,N_10225);
and U11211 (N_11211,N_10378,N_10037);
and U11212 (N_11212,N_10413,N_10054);
and U11213 (N_11213,N_10400,N_10491);
nor U11214 (N_11214,N_10691,N_10335);
xnor U11215 (N_11215,N_10174,N_10886);
xnor U11216 (N_11216,N_10818,N_10484);
and U11217 (N_11217,N_10900,N_10201);
or U11218 (N_11218,N_10206,N_10837);
and U11219 (N_11219,N_10094,N_10087);
or U11220 (N_11220,N_10993,N_10377);
or U11221 (N_11221,N_10812,N_10464);
or U11222 (N_11222,N_10314,N_10132);
nand U11223 (N_11223,N_10211,N_10698);
nor U11224 (N_11224,N_10961,N_10238);
or U11225 (N_11225,N_10391,N_10522);
and U11226 (N_11226,N_10547,N_10940);
nand U11227 (N_11227,N_10763,N_10216);
or U11228 (N_11228,N_10885,N_10566);
xor U11229 (N_11229,N_10747,N_10397);
xnor U11230 (N_11230,N_10750,N_10320);
or U11231 (N_11231,N_10925,N_10604);
nand U11232 (N_11232,N_10945,N_10146);
and U11233 (N_11233,N_10259,N_10119);
nand U11234 (N_11234,N_10535,N_10870);
and U11235 (N_11235,N_10694,N_10972);
or U11236 (N_11236,N_10736,N_10234);
xnor U11237 (N_11237,N_10689,N_10062);
xnor U11238 (N_11238,N_10749,N_10021);
or U11239 (N_11239,N_10374,N_10468);
or U11240 (N_11240,N_10597,N_10137);
nand U11241 (N_11241,N_10013,N_10339);
nand U11242 (N_11242,N_10695,N_10610);
or U11243 (N_11243,N_10163,N_10568);
nor U11244 (N_11244,N_10068,N_10682);
and U11245 (N_11245,N_10601,N_10661);
nor U11246 (N_11246,N_10128,N_10005);
nor U11247 (N_11247,N_10965,N_10594);
xor U11248 (N_11248,N_10700,N_10734);
nand U11249 (N_11249,N_10359,N_10254);
and U11250 (N_11250,N_10762,N_10669);
or U11251 (N_11251,N_10235,N_10505);
nor U11252 (N_11252,N_10901,N_10544);
and U11253 (N_11253,N_10007,N_10495);
xor U11254 (N_11254,N_10859,N_10745);
nand U11255 (N_11255,N_10263,N_10018);
and U11256 (N_11256,N_10618,N_10775);
xor U11257 (N_11257,N_10409,N_10488);
xor U11258 (N_11258,N_10773,N_10541);
and U11259 (N_11259,N_10134,N_10260);
or U11260 (N_11260,N_10176,N_10160);
or U11261 (N_11261,N_10814,N_10632);
nor U11262 (N_11262,N_10057,N_10501);
nand U11263 (N_11263,N_10910,N_10692);
xor U11264 (N_11264,N_10991,N_10108);
xor U11265 (N_11265,N_10737,N_10304);
and U11266 (N_11266,N_10890,N_10049);
or U11267 (N_11267,N_10408,N_10585);
nor U11268 (N_11268,N_10721,N_10557);
or U11269 (N_11269,N_10785,N_10349);
nand U11270 (N_11270,N_10347,N_10471);
and U11271 (N_11271,N_10161,N_10858);
xor U11272 (N_11272,N_10609,N_10239);
nand U11273 (N_11273,N_10485,N_10530);
and U11274 (N_11274,N_10976,N_10820);
nor U11275 (N_11275,N_10266,N_10099);
xnor U11276 (N_11276,N_10642,N_10701);
xnor U11277 (N_11277,N_10402,N_10524);
or U11278 (N_11278,N_10917,N_10831);
or U11279 (N_11279,N_10690,N_10939);
and U11280 (N_11280,N_10538,N_10452);
nand U11281 (N_11281,N_10357,N_10952);
nor U11282 (N_11282,N_10551,N_10265);
nor U11283 (N_11283,N_10275,N_10117);
xor U11284 (N_11284,N_10881,N_10173);
and U11285 (N_11285,N_10268,N_10157);
nand U11286 (N_11286,N_10217,N_10565);
nor U11287 (N_11287,N_10312,N_10188);
nand U11288 (N_11288,N_10527,N_10879);
and U11289 (N_11289,N_10914,N_10836);
and U11290 (N_11290,N_10685,N_10075);
xor U11291 (N_11291,N_10059,N_10977);
and U11292 (N_11292,N_10353,N_10559);
nand U11293 (N_11293,N_10599,N_10696);
xor U11294 (N_11294,N_10571,N_10906);
xnor U11295 (N_11295,N_10857,N_10844);
nand U11296 (N_11296,N_10446,N_10267);
or U11297 (N_11297,N_10670,N_10718);
or U11298 (N_11298,N_10771,N_10373);
nor U11299 (N_11299,N_10504,N_10981);
and U11300 (N_11300,N_10653,N_10258);
nor U11301 (N_11301,N_10344,N_10319);
nand U11302 (N_11302,N_10487,N_10624);
nor U11303 (N_11303,N_10285,N_10828);
nand U11304 (N_11304,N_10286,N_10894);
or U11305 (N_11305,N_10598,N_10424);
and U11306 (N_11306,N_10593,N_10003);
nor U11307 (N_11307,N_10492,N_10989);
and U11308 (N_11308,N_10318,N_10218);
nand U11309 (N_11309,N_10269,N_10362);
nor U11310 (N_11310,N_10650,N_10281);
xor U11311 (N_11311,N_10125,N_10562);
or U11312 (N_11312,N_10880,N_10162);
xor U11313 (N_11313,N_10434,N_10222);
xor U11314 (N_11314,N_10558,N_10953);
nand U11315 (N_11315,N_10165,N_10129);
xnor U11316 (N_11316,N_10416,N_10490);
xnor U11317 (N_11317,N_10840,N_10172);
and U11318 (N_11318,N_10136,N_10748);
or U11319 (N_11319,N_10983,N_10948);
and U11320 (N_11320,N_10529,N_10937);
xor U11321 (N_11321,N_10456,N_10046);
xor U11322 (N_11322,N_10600,N_10064);
xnor U11323 (N_11323,N_10864,N_10231);
nor U11324 (N_11324,N_10703,N_10289);
nor U11325 (N_11325,N_10574,N_10570);
or U11326 (N_11326,N_10956,N_10832);
nor U11327 (N_11327,N_10227,N_10919);
nand U11328 (N_11328,N_10197,N_10532);
or U11329 (N_11329,N_10215,N_10819);
nor U11330 (N_11330,N_10461,N_10668);
nor U11331 (N_11331,N_10825,N_10060);
and U11332 (N_11332,N_10177,N_10786);
nand U11333 (N_11333,N_10272,N_10794);
and U11334 (N_11334,N_10182,N_10144);
and U11335 (N_11335,N_10308,N_10951);
nand U11336 (N_11336,N_10780,N_10051);
xnor U11337 (N_11337,N_10569,N_10229);
xor U11338 (N_11338,N_10802,N_10896);
nand U11339 (N_11339,N_10331,N_10483);
nand U11340 (N_11340,N_10477,N_10435);
or U11341 (N_11341,N_10190,N_10908);
or U11342 (N_11342,N_10966,N_10418);
nor U11343 (N_11343,N_10232,N_10104);
nand U11344 (N_11344,N_10542,N_10052);
nand U11345 (N_11345,N_10770,N_10717);
nor U11346 (N_11346,N_10623,N_10799);
and U11347 (N_11347,N_10608,N_10368);
xnor U11348 (N_11348,N_10386,N_10611);
xor U11349 (N_11349,N_10628,N_10957);
nand U11350 (N_11350,N_10061,N_10360);
nor U11351 (N_11351,N_10662,N_10779);
and U11352 (N_11352,N_10380,N_10947);
nor U11353 (N_11353,N_10921,N_10572);
nand U11354 (N_11354,N_10605,N_10639);
or U11355 (N_11355,N_10944,N_10101);
xor U11356 (N_11356,N_10808,N_10998);
nor U11357 (N_11357,N_10158,N_10109);
and U11358 (N_11358,N_10823,N_10526);
xor U11359 (N_11359,N_10942,N_10026);
and U11360 (N_11360,N_10496,N_10325);
and U11361 (N_11361,N_10667,N_10441);
nand U11362 (N_11362,N_10727,N_10978);
and U11363 (N_11363,N_10436,N_10241);
or U11364 (N_11364,N_10296,N_10138);
and U11365 (N_11365,N_10846,N_10856);
nand U11366 (N_11366,N_10303,N_10898);
nor U11367 (N_11367,N_10540,N_10017);
xnor U11368 (N_11368,N_10093,N_10294);
xor U11369 (N_11369,N_10782,N_10506);
xor U11370 (N_11370,N_10187,N_10210);
nand U11371 (N_11371,N_10337,N_10323);
nand U11372 (N_11372,N_10982,N_10990);
nor U11373 (N_11373,N_10000,N_10822);
xor U11374 (N_11374,N_10681,N_10358);
nor U11375 (N_11375,N_10647,N_10245);
xnor U11376 (N_11376,N_10412,N_10056);
nor U11377 (N_11377,N_10539,N_10082);
xor U11378 (N_11378,N_10482,N_10985);
nor U11379 (N_11379,N_10022,N_10058);
nand U11380 (N_11380,N_10911,N_10035);
nand U11381 (N_11381,N_10616,N_10549);
xnor U11382 (N_11382,N_10723,N_10651);
nand U11383 (N_11383,N_10995,N_10854);
xnor U11384 (N_11384,N_10462,N_10224);
and U11385 (N_11385,N_10648,N_10015);
or U11386 (N_11386,N_10195,N_10577);
xnor U11387 (N_11387,N_10725,N_10833);
or U11388 (N_11388,N_10636,N_10793);
xor U11389 (N_11389,N_10509,N_10591);
nor U11390 (N_11390,N_10106,N_10803);
and U11391 (N_11391,N_10432,N_10554);
nor U11392 (N_11392,N_10425,N_10741);
or U11393 (N_11393,N_10179,N_10958);
and U11394 (N_11394,N_10817,N_10113);
nand U11395 (N_11395,N_10631,N_10428);
nand U11396 (N_11396,N_10463,N_10735);
xor U11397 (N_11397,N_10186,N_10324);
and U11398 (N_11398,N_10969,N_10615);
nor U11399 (N_11399,N_10533,N_10935);
xor U11400 (N_11400,N_10523,N_10996);
and U11401 (N_11401,N_10602,N_10209);
or U11402 (N_11402,N_10979,N_10519);
xor U11403 (N_11403,N_10091,N_10674);
and U11404 (N_11404,N_10561,N_10084);
nor U11405 (N_11405,N_10876,N_10247);
or U11406 (N_11406,N_10419,N_10169);
and U11407 (N_11407,N_10200,N_10658);
and U11408 (N_11408,N_10111,N_10345);
nor U11409 (N_11409,N_10913,N_10924);
and U11410 (N_11410,N_10699,N_10552);
xor U11411 (N_11411,N_10537,N_10626);
or U11412 (N_11412,N_10841,N_10379);
and U11413 (N_11413,N_10797,N_10730);
xnor U11414 (N_11414,N_10475,N_10498);
nor U11415 (N_11415,N_10563,N_10205);
nor U11416 (N_11416,N_10742,N_10170);
nor U11417 (N_11417,N_10708,N_10664);
or U11418 (N_11418,N_10467,N_10024);
nand U11419 (N_11419,N_10777,N_10047);
nand U11420 (N_11420,N_10904,N_10677);
xor U11421 (N_11421,N_10665,N_10433);
or U11422 (N_11422,N_10284,N_10918);
and U11423 (N_11423,N_10050,N_10916);
or U11424 (N_11424,N_10861,N_10429);
xnor U11425 (N_11425,N_10454,N_10466);
nor U11426 (N_11426,N_10032,N_10791);
and U11427 (N_11427,N_10447,N_10427);
nor U11428 (N_11428,N_10330,N_10545);
or U11429 (N_11429,N_10738,N_10317);
nand U11430 (N_11430,N_10882,N_10204);
and U11431 (N_11431,N_10372,N_10580);
or U11432 (N_11432,N_10192,N_10892);
or U11433 (N_11433,N_10293,N_10933);
or U11434 (N_11434,N_10316,N_10997);
and U11435 (N_11435,N_10637,N_10932);
nor U11436 (N_11436,N_10048,N_10431);
nand U11437 (N_11437,N_10376,N_10028);
nor U11438 (N_11438,N_10865,N_10867);
or U11439 (N_11439,N_10596,N_10045);
xnor U11440 (N_11440,N_10090,N_10309);
nor U11441 (N_11441,N_10678,N_10553);
and U11442 (N_11442,N_10124,N_10189);
and U11443 (N_11443,N_10307,N_10641);
and U11444 (N_11444,N_10555,N_10884);
or U11445 (N_11445,N_10112,N_10630);
nor U11446 (N_11446,N_10096,N_10702);
nand U11447 (N_11447,N_10352,N_10039);
nand U11448 (N_11448,N_10500,N_10407);
nor U11449 (N_11449,N_10193,N_10041);
or U11450 (N_11450,N_10974,N_10790);
xnor U11451 (N_11451,N_10759,N_10724);
nand U11452 (N_11452,N_10271,N_10987);
or U11453 (N_11453,N_10946,N_10280);
xor U11454 (N_11454,N_10713,N_10255);
xor U11455 (N_11455,N_10654,N_10404);
nor U11456 (N_11456,N_10973,N_10874);
xor U11457 (N_11457,N_10853,N_10576);
xor U11458 (N_11458,N_10310,N_10514);
nor U11459 (N_11459,N_10422,N_10249);
and U11460 (N_11460,N_10807,N_10142);
nor U11461 (N_11461,N_10363,N_10595);
and U11462 (N_11462,N_10810,N_10020);
xor U11463 (N_11463,N_10141,N_10971);
nand U11464 (N_11464,N_10355,N_10706);
xor U11465 (N_11465,N_10126,N_10479);
nor U11466 (N_11466,N_10329,N_10511);
nor U11467 (N_11467,N_10411,N_10582);
xnor U11468 (N_11468,N_10074,N_10185);
nor U11469 (N_11469,N_10697,N_10784);
and U11470 (N_11470,N_10191,N_10080);
nand U11471 (N_11471,N_10878,N_10417);
or U11472 (N_11472,N_10326,N_10398);
nand U11473 (N_11473,N_10503,N_10909);
and U11474 (N_11474,N_10167,N_10006);
and U11475 (N_11475,N_10274,N_10753);
and U11476 (N_11476,N_10603,N_10531);
or U11477 (N_11477,N_10069,N_10297);
xor U11478 (N_11478,N_10100,N_10299);
nand U11479 (N_11479,N_10936,N_10261);
nand U11480 (N_11480,N_10955,N_10589);
and U11481 (N_11481,N_10806,N_10860);
xor U11482 (N_11482,N_10877,N_10394);
xor U11483 (N_11483,N_10711,N_10306);
xor U11484 (N_11484,N_10663,N_10798);
nand U11485 (N_11485,N_10672,N_10534);
or U11486 (N_11486,N_10760,N_10517);
xnor U11487 (N_11487,N_10766,N_10171);
or U11488 (N_11488,N_10586,N_10796);
and U11489 (N_11489,N_10556,N_10567);
nor U11490 (N_11490,N_10465,N_10899);
nand U11491 (N_11491,N_10673,N_10034);
xor U11492 (N_11492,N_10986,N_10684);
nand U11493 (N_11493,N_10740,N_10676);
or U11494 (N_11494,N_10114,N_10934);
or U11495 (N_11495,N_10085,N_10915);
or U11496 (N_11496,N_10342,N_10181);
nand U11497 (N_11497,N_10451,N_10835);
and U11498 (N_11498,N_10795,N_10388);
nor U11499 (N_11499,N_10826,N_10764);
xor U11500 (N_11500,N_10365,N_10545);
or U11501 (N_11501,N_10278,N_10161);
nand U11502 (N_11502,N_10560,N_10062);
xnor U11503 (N_11503,N_10987,N_10076);
xnor U11504 (N_11504,N_10103,N_10118);
nor U11505 (N_11505,N_10184,N_10503);
xor U11506 (N_11506,N_10935,N_10079);
and U11507 (N_11507,N_10775,N_10194);
or U11508 (N_11508,N_10064,N_10774);
or U11509 (N_11509,N_10276,N_10838);
nor U11510 (N_11510,N_10301,N_10021);
or U11511 (N_11511,N_10140,N_10348);
nor U11512 (N_11512,N_10697,N_10554);
and U11513 (N_11513,N_10816,N_10549);
and U11514 (N_11514,N_10326,N_10986);
or U11515 (N_11515,N_10413,N_10614);
and U11516 (N_11516,N_10416,N_10106);
and U11517 (N_11517,N_10141,N_10324);
nor U11518 (N_11518,N_10501,N_10631);
nand U11519 (N_11519,N_10265,N_10843);
or U11520 (N_11520,N_10645,N_10571);
nand U11521 (N_11521,N_10938,N_10730);
or U11522 (N_11522,N_10546,N_10065);
xnor U11523 (N_11523,N_10927,N_10677);
or U11524 (N_11524,N_10571,N_10598);
or U11525 (N_11525,N_10396,N_10782);
and U11526 (N_11526,N_10554,N_10400);
nand U11527 (N_11527,N_10931,N_10314);
xnor U11528 (N_11528,N_10524,N_10670);
and U11529 (N_11529,N_10148,N_10526);
xor U11530 (N_11530,N_10440,N_10089);
xor U11531 (N_11531,N_10001,N_10958);
nand U11532 (N_11532,N_10629,N_10315);
and U11533 (N_11533,N_10439,N_10382);
and U11534 (N_11534,N_10456,N_10496);
nor U11535 (N_11535,N_10665,N_10349);
xnor U11536 (N_11536,N_10034,N_10402);
nor U11537 (N_11537,N_10374,N_10875);
xnor U11538 (N_11538,N_10636,N_10164);
and U11539 (N_11539,N_10199,N_10112);
xor U11540 (N_11540,N_10640,N_10162);
nor U11541 (N_11541,N_10932,N_10152);
and U11542 (N_11542,N_10527,N_10091);
nor U11543 (N_11543,N_10948,N_10263);
xor U11544 (N_11544,N_10443,N_10917);
or U11545 (N_11545,N_10866,N_10218);
xor U11546 (N_11546,N_10768,N_10709);
xnor U11547 (N_11547,N_10374,N_10637);
xor U11548 (N_11548,N_10161,N_10467);
nor U11549 (N_11549,N_10159,N_10766);
xor U11550 (N_11550,N_10007,N_10912);
or U11551 (N_11551,N_10839,N_10977);
and U11552 (N_11552,N_10191,N_10724);
or U11553 (N_11553,N_10487,N_10703);
or U11554 (N_11554,N_10361,N_10842);
and U11555 (N_11555,N_10663,N_10988);
nor U11556 (N_11556,N_10738,N_10493);
and U11557 (N_11557,N_10926,N_10302);
nand U11558 (N_11558,N_10381,N_10437);
and U11559 (N_11559,N_10476,N_10603);
nor U11560 (N_11560,N_10682,N_10255);
nand U11561 (N_11561,N_10316,N_10189);
xor U11562 (N_11562,N_10506,N_10775);
and U11563 (N_11563,N_10367,N_10794);
or U11564 (N_11564,N_10953,N_10300);
nor U11565 (N_11565,N_10963,N_10744);
and U11566 (N_11566,N_10970,N_10027);
xnor U11567 (N_11567,N_10876,N_10880);
nand U11568 (N_11568,N_10040,N_10705);
nor U11569 (N_11569,N_10586,N_10731);
and U11570 (N_11570,N_10143,N_10739);
nor U11571 (N_11571,N_10270,N_10788);
nand U11572 (N_11572,N_10213,N_10632);
and U11573 (N_11573,N_10277,N_10661);
and U11574 (N_11574,N_10588,N_10657);
and U11575 (N_11575,N_10382,N_10346);
or U11576 (N_11576,N_10088,N_10169);
nand U11577 (N_11577,N_10152,N_10964);
xor U11578 (N_11578,N_10685,N_10490);
nand U11579 (N_11579,N_10373,N_10498);
xor U11580 (N_11580,N_10571,N_10587);
and U11581 (N_11581,N_10292,N_10236);
and U11582 (N_11582,N_10649,N_10336);
and U11583 (N_11583,N_10282,N_10052);
nand U11584 (N_11584,N_10079,N_10748);
nor U11585 (N_11585,N_10309,N_10712);
nand U11586 (N_11586,N_10137,N_10697);
xor U11587 (N_11587,N_10674,N_10071);
xor U11588 (N_11588,N_10563,N_10743);
xor U11589 (N_11589,N_10826,N_10639);
xnor U11590 (N_11590,N_10085,N_10150);
or U11591 (N_11591,N_10908,N_10164);
and U11592 (N_11592,N_10724,N_10953);
or U11593 (N_11593,N_10390,N_10558);
nand U11594 (N_11594,N_10254,N_10991);
or U11595 (N_11595,N_10674,N_10339);
or U11596 (N_11596,N_10488,N_10822);
nand U11597 (N_11597,N_10375,N_10346);
and U11598 (N_11598,N_10858,N_10968);
nand U11599 (N_11599,N_10340,N_10135);
xnor U11600 (N_11600,N_10275,N_10574);
and U11601 (N_11601,N_10974,N_10468);
and U11602 (N_11602,N_10260,N_10223);
nand U11603 (N_11603,N_10583,N_10898);
xnor U11604 (N_11604,N_10784,N_10853);
and U11605 (N_11605,N_10881,N_10217);
nor U11606 (N_11606,N_10663,N_10090);
nor U11607 (N_11607,N_10347,N_10348);
and U11608 (N_11608,N_10949,N_10199);
nand U11609 (N_11609,N_10936,N_10362);
nor U11610 (N_11610,N_10141,N_10442);
and U11611 (N_11611,N_10479,N_10005);
xnor U11612 (N_11612,N_10490,N_10449);
nor U11613 (N_11613,N_10139,N_10325);
and U11614 (N_11614,N_10291,N_10153);
nor U11615 (N_11615,N_10397,N_10224);
nand U11616 (N_11616,N_10956,N_10542);
nor U11617 (N_11617,N_10457,N_10607);
nor U11618 (N_11618,N_10866,N_10031);
nand U11619 (N_11619,N_10186,N_10593);
nand U11620 (N_11620,N_10087,N_10519);
nor U11621 (N_11621,N_10898,N_10726);
and U11622 (N_11622,N_10563,N_10032);
nand U11623 (N_11623,N_10287,N_10335);
and U11624 (N_11624,N_10199,N_10044);
xnor U11625 (N_11625,N_10577,N_10253);
xnor U11626 (N_11626,N_10877,N_10812);
and U11627 (N_11627,N_10451,N_10119);
nand U11628 (N_11628,N_10774,N_10399);
and U11629 (N_11629,N_10971,N_10389);
and U11630 (N_11630,N_10249,N_10595);
and U11631 (N_11631,N_10854,N_10445);
nor U11632 (N_11632,N_10708,N_10460);
xnor U11633 (N_11633,N_10268,N_10028);
or U11634 (N_11634,N_10042,N_10926);
and U11635 (N_11635,N_10492,N_10690);
xor U11636 (N_11636,N_10463,N_10787);
nor U11637 (N_11637,N_10353,N_10250);
nor U11638 (N_11638,N_10813,N_10193);
nand U11639 (N_11639,N_10943,N_10212);
nor U11640 (N_11640,N_10014,N_10276);
and U11641 (N_11641,N_10324,N_10968);
nor U11642 (N_11642,N_10124,N_10465);
nor U11643 (N_11643,N_10012,N_10986);
and U11644 (N_11644,N_10239,N_10774);
nor U11645 (N_11645,N_10444,N_10577);
nand U11646 (N_11646,N_10317,N_10203);
and U11647 (N_11647,N_10407,N_10993);
or U11648 (N_11648,N_10495,N_10059);
and U11649 (N_11649,N_10388,N_10030);
xnor U11650 (N_11650,N_10252,N_10460);
xor U11651 (N_11651,N_10599,N_10335);
nor U11652 (N_11652,N_10252,N_10893);
or U11653 (N_11653,N_10356,N_10159);
xnor U11654 (N_11654,N_10934,N_10239);
or U11655 (N_11655,N_10030,N_10875);
nor U11656 (N_11656,N_10442,N_10592);
nor U11657 (N_11657,N_10609,N_10828);
or U11658 (N_11658,N_10022,N_10296);
nand U11659 (N_11659,N_10568,N_10179);
and U11660 (N_11660,N_10219,N_10852);
nand U11661 (N_11661,N_10291,N_10076);
nor U11662 (N_11662,N_10845,N_10387);
nor U11663 (N_11663,N_10086,N_10589);
or U11664 (N_11664,N_10954,N_10982);
xor U11665 (N_11665,N_10891,N_10098);
and U11666 (N_11666,N_10415,N_10489);
or U11667 (N_11667,N_10429,N_10511);
xnor U11668 (N_11668,N_10892,N_10406);
nor U11669 (N_11669,N_10603,N_10292);
and U11670 (N_11670,N_10665,N_10628);
xor U11671 (N_11671,N_10746,N_10203);
nor U11672 (N_11672,N_10411,N_10748);
nor U11673 (N_11673,N_10393,N_10483);
xor U11674 (N_11674,N_10635,N_10384);
or U11675 (N_11675,N_10783,N_10722);
and U11676 (N_11676,N_10740,N_10759);
or U11677 (N_11677,N_10946,N_10080);
and U11678 (N_11678,N_10592,N_10091);
nor U11679 (N_11679,N_10648,N_10714);
or U11680 (N_11680,N_10600,N_10360);
and U11681 (N_11681,N_10511,N_10649);
nand U11682 (N_11682,N_10867,N_10561);
and U11683 (N_11683,N_10110,N_10424);
or U11684 (N_11684,N_10701,N_10908);
and U11685 (N_11685,N_10638,N_10036);
nand U11686 (N_11686,N_10006,N_10518);
nor U11687 (N_11687,N_10203,N_10345);
and U11688 (N_11688,N_10514,N_10093);
xor U11689 (N_11689,N_10182,N_10460);
or U11690 (N_11690,N_10894,N_10826);
xor U11691 (N_11691,N_10287,N_10898);
and U11692 (N_11692,N_10534,N_10434);
or U11693 (N_11693,N_10767,N_10250);
xor U11694 (N_11694,N_10217,N_10030);
and U11695 (N_11695,N_10884,N_10226);
xnor U11696 (N_11696,N_10464,N_10043);
or U11697 (N_11697,N_10395,N_10464);
xnor U11698 (N_11698,N_10462,N_10999);
nor U11699 (N_11699,N_10449,N_10842);
xnor U11700 (N_11700,N_10762,N_10231);
and U11701 (N_11701,N_10872,N_10009);
or U11702 (N_11702,N_10111,N_10890);
and U11703 (N_11703,N_10685,N_10648);
and U11704 (N_11704,N_10812,N_10011);
nor U11705 (N_11705,N_10793,N_10340);
and U11706 (N_11706,N_10494,N_10560);
xnor U11707 (N_11707,N_10377,N_10336);
and U11708 (N_11708,N_10261,N_10581);
or U11709 (N_11709,N_10214,N_10245);
or U11710 (N_11710,N_10713,N_10554);
xnor U11711 (N_11711,N_10008,N_10801);
nand U11712 (N_11712,N_10125,N_10435);
xnor U11713 (N_11713,N_10621,N_10561);
or U11714 (N_11714,N_10428,N_10637);
nand U11715 (N_11715,N_10353,N_10747);
xor U11716 (N_11716,N_10568,N_10269);
and U11717 (N_11717,N_10083,N_10811);
and U11718 (N_11718,N_10187,N_10241);
nor U11719 (N_11719,N_10704,N_10948);
nand U11720 (N_11720,N_10036,N_10289);
nor U11721 (N_11721,N_10701,N_10100);
xnor U11722 (N_11722,N_10550,N_10270);
xnor U11723 (N_11723,N_10234,N_10935);
nand U11724 (N_11724,N_10416,N_10936);
and U11725 (N_11725,N_10055,N_10687);
xor U11726 (N_11726,N_10033,N_10598);
xor U11727 (N_11727,N_10807,N_10735);
nand U11728 (N_11728,N_10421,N_10086);
nor U11729 (N_11729,N_10698,N_10440);
xor U11730 (N_11730,N_10692,N_10979);
xnor U11731 (N_11731,N_10259,N_10210);
nor U11732 (N_11732,N_10237,N_10303);
nor U11733 (N_11733,N_10730,N_10315);
xor U11734 (N_11734,N_10953,N_10363);
and U11735 (N_11735,N_10791,N_10063);
xnor U11736 (N_11736,N_10350,N_10527);
nor U11737 (N_11737,N_10218,N_10650);
nor U11738 (N_11738,N_10395,N_10119);
nor U11739 (N_11739,N_10845,N_10789);
or U11740 (N_11740,N_10254,N_10112);
and U11741 (N_11741,N_10033,N_10151);
xnor U11742 (N_11742,N_10888,N_10507);
nor U11743 (N_11743,N_10962,N_10055);
nor U11744 (N_11744,N_10997,N_10389);
xor U11745 (N_11745,N_10822,N_10850);
nand U11746 (N_11746,N_10114,N_10738);
and U11747 (N_11747,N_10108,N_10751);
xor U11748 (N_11748,N_10536,N_10717);
or U11749 (N_11749,N_10145,N_10121);
and U11750 (N_11750,N_10398,N_10831);
and U11751 (N_11751,N_10674,N_10680);
and U11752 (N_11752,N_10954,N_10043);
xor U11753 (N_11753,N_10462,N_10478);
nor U11754 (N_11754,N_10244,N_10487);
nor U11755 (N_11755,N_10233,N_10894);
nand U11756 (N_11756,N_10379,N_10906);
or U11757 (N_11757,N_10618,N_10097);
nor U11758 (N_11758,N_10485,N_10931);
nand U11759 (N_11759,N_10581,N_10313);
nor U11760 (N_11760,N_10044,N_10501);
and U11761 (N_11761,N_10151,N_10188);
xor U11762 (N_11762,N_10504,N_10681);
nand U11763 (N_11763,N_10247,N_10535);
nor U11764 (N_11764,N_10662,N_10335);
xnor U11765 (N_11765,N_10047,N_10179);
nand U11766 (N_11766,N_10266,N_10722);
nand U11767 (N_11767,N_10851,N_10321);
or U11768 (N_11768,N_10535,N_10541);
xor U11769 (N_11769,N_10966,N_10301);
nand U11770 (N_11770,N_10572,N_10951);
nand U11771 (N_11771,N_10656,N_10382);
nand U11772 (N_11772,N_10593,N_10753);
nand U11773 (N_11773,N_10419,N_10569);
xnor U11774 (N_11774,N_10852,N_10714);
or U11775 (N_11775,N_10221,N_10928);
or U11776 (N_11776,N_10499,N_10676);
nor U11777 (N_11777,N_10903,N_10364);
and U11778 (N_11778,N_10720,N_10596);
nor U11779 (N_11779,N_10807,N_10885);
nor U11780 (N_11780,N_10603,N_10390);
xnor U11781 (N_11781,N_10955,N_10794);
and U11782 (N_11782,N_10516,N_10811);
nor U11783 (N_11783,N_10854,N_10062);
nor U11784 (N_11784,N_10442,N_10950);
nand U11785 (N_11785,N_10403,N_10557);
xor U11786 (N_11786,N_10784,N_10277);
or U11787 (N_11787,N_10929,N_10251);
and U11788 (N_11788,N_10243,N_10744);
and U11789 (N_11789,N_10498,N_10927);
nor U11790 (N_11790,N_10241,N_10668);
and U11791 (N_11791,N_10610,N_10894);
or U11792 (N_11792,N_10563,N_10109);
or U11793 (N_11793,N_10746,N_10405);
nor U11794 (N_11794,N_10769,N_10437);
or U11795 (N_11795,N_10723,N_10313);
nor U11796 (N_11796,N_10736,N_10130);
xor U11797 (N_11797,N_10866,N_10252);
nor U11798 (N_11798,N_10263,N_10873);
or U11799 (N_11799,N_10637,N_10246);
xnor U11800 (N_11800,N_10352,N_10972);
xor U11801 (N_11801,N_10624,N_10613);
and U11802 (N_11802,N_10397,N_10688);
or U11803 (N_11803,N_10892,N_10753);
nor U11804 (N_11804,N_10717,N_10454);
nand U11805 (N_11805,N_10822,N_10540);
and U11806 (N_11806,N_10536,N_10086);
nor U11807 (N_11807,N_10275,N_10253);
nand U11808 (N_11808,N_10562,N_10131);
nand U11809 (N_11809,N_10102,N_10147);
xor U11810 (N_11810,N_10564,N_10890);
xnor U11811 (N_11811,N_10005,N_10726);
and U11812 (N_11812,N_10247,N_10296);
and U11813 (N_11813,N_10434,N_10218);
xor U11814 (N_11814,N_10106,N_10609);
nand U11815 (N_11815,N_10817,N_10953);
nand U11816 (N_11816,N_10147,N_10067);
or U11817 (N_11817,N_10103,N_10889);
xor U11818 (N_11818,N_10115,N_10593);
xor U11819 (N_11819,N_10316,N_10685);
nand U11820 (N_11820,N_10140,N_10135);
nor U11821 (N_11821,N_10077,N_10208);
and U11822 (N_11822,N_10238,N_10668);
or U11823 (N_11823,N_10716,N_10285);
xnor U11824 (N_11824,N_10314,N_10243);
or U11825 (N_11825,N_10910,N_10817);
and U11826 (N_11826,N_10885,N_10242);
nand U11827 (N_11827,N_10452,N_10394);
nor U11828 (N_11828,N_10068,N_10234);
nor U11829 (N_11829,N_10153,N_10517);
or U11830 (N_11830,N_10712,N_10159);
nor U11831 (N_11831,N_10732,N_10339);
nand U11832 (N_11832,N_10725,N_10929);
or U11833 (N_11833,N_10703,N_10319);
xnor U11834 (N_11834,N_10331,N_10101);
xor U11835 (N_11835,N_10752,N_10202);
nor U11836 (N_11836,N_10219,N_10964);
nand U11837 (N_11837,N_10429,N_10560);
nand U11838 (N_11838,N_10815,N_10274);
nor U11839 (N_11839,N_10375,N_10291);
or U11840 (N_11840,N_10240,N_10611);
nand U11841 (N_11841,N_10784,N_10097);
nand U11842 (N_11842,N_10881,N_10682);
nor U11843 (N_11843,N_10070,N_10800);
xnor U11844 (N_11844,N_10392,N_10774);
xor U11845 (N_11845,N_10532,N_10975);
nor U11846 (N_11846,N_10834,N_10074);
xnor U11847 (N_11847,N_10893,N_10543);
xor U11848 (N_11848,N_10272,N_10921);
xnor U11849 (N_11849,N_10048,N_10542);
and U11850 (N_11850,N_10463,N_10018);
xor U11851 (N_11851,N_10500,N_10256);
nand U11852 (N_11852,N_10376,N_10481);
nor U11853 (N_11853,N_10111,N_10786);
or U11854 (N_11854,N_10101,N_10292);
xnor U11855 (N_11855,N_10269,N_10064);
and U11856 (N_11856,N_10190,N_10827);
and U11857 (N_11857,N_10261,N_10414);
and U11858 (N_11858,N_10092,N_10190);
nand U11859 (N_11859,N_10849,N_10646);
nor U11860 (N_11860,N_10897,N_10866);
xor U11861 (N_11861,N_10096,N_10021);
and U11862 (N_11862,N_10194,N_10325);
xor U11863 (N_11863,N_10738,N_10912);
xnor U11864 (N_11864,N_10704,N_10697);
and U11865 (N_11865,N_10328,N_10364);
nand U11866 (N_11866,N_10334,N_10331);
or U11867 (N_11867,N_10870,N_10685);
and U11868 (N_11868,N_10848,N_10028);
or U11869 (N_11869,N_10124,N_10475);
nor U11870 (N_11870,N_10169,N_10774);
xor U11871 (N_11871,N_10751,N_10278);
or U11872 (N_11872,N_10874,N_10409);
xnor U11873 (N_11873,N_10032,N_10255);
nand U11874 (N_11874,N_10109,N_10266);
xnor U11875 (N_11875,N_10143,N_10259);
nor U11876 (N_11876,N_10456,N_10895);
nand U11877 (N_11877,N_10284,N_10489);
nor U11878 (N_11878,N_10689,N_10450);
or U11879 (N_11879,N_10312,N_10539);
xnor U11880 (N_11880,N_10259,N_10736);
or U11881 (N_11881,N_10076,N_10400);
or U11882 (N_11882,N_10911,N_10798);
nor U11883 (N_11883,N_10058,N_10666);
xor U11884 (N_11884,N_10638,N_10311);
xnor U11885 (N_11885,N_10704,N_10188);
and U11886 (N_11886,N_10860,N_10269);
xnor U11887 (N_11887,N_10108,N_10467);
nand U11888 (N_11888,N_10526,N_10271);
nor U11889 (N_11889,N_10443,N_10842);
nor U11890 (N_11890,N_10191,N_10687);
nand U11891 (N_11891,N_10311,N_10925);
nor U11892 (N_11892,N_10938,N_10617);
and U11893 (N_11893,N_10762,N_10278);
and U11894 (N_11894,N_10237,N_10761);
nor U11895 (N_11895,N_10278,N_10910);
nand U11896 (N_11896,N_10952,N_10887);
nor U11897 (N_11897,N_10471,N_10969);
nor U11898 (N_11898,N_10536,N_10586);
nand U11899 (N_11899,N_10065,N_10940);
xnor U11900 (N_11900,N_10430,N_10411);
nor U11901 (N_11901,N_10966,N_10809);
or U11902 (N_11902,N_10772,N_10093);
or U11903 (N_11903,N_10166,N_10324);
and U11904 (N_11904,N_10285,N_10164);
and U11905 (N_11905,N_10662,N_10077);
xnor U11906 (N_11906,N_10211,N_10477);
xor U11907 (N_11907,N_10395,N_10060);
and U11908 (N_11908,N_10184,N_10968);
or U11909 (N_11909,N_10459,N_10551);
nand U11910 (N_11910,N_10915,N_10157);
xor U11911 (N_11911,N_10337,N_10633);
or U11912 (N_11912,N_10638,N_10068);
nand U11913 (N_11913,N_10542,N_10849);
nor U11914 (N_11914,N_10028,N_10139);
or U11915 (N_11915,N_10211,N_10710);
xnor U11916 (N_11916,N_10088,N_10562);
nand U11917 (N_11917,N_10588,N_10120);
or U11918 (N_11918,N_10538,N_10864);
or U11919 (N_11919,N_10153,N_10389);
nor U11920 (N_11920,N_10368,N_10816);
or U11921 (N_11921,N_10205,N_10530);
or U11922 (N_11922,N_10370,N_10719);
and U11923 (N_11923,N_10648,N_10090);
nand U11924 (N_11924,N_10718,N_10476);
nand U11925 (N_11925,N_10485,N_10412);
nand U11926 (N_11926,N_10024,N_10910);
or U11927 (N_11927,N_10402,N_10860);
nor U11928 (N_11928,N_10634,N_10494);
or U11929 (N_11929,N_10337,N_10244);
nand U11930 (N_11930,N_10364,N_10634);
nor U11931 (N_11931,N_10391,N_10031);
nor U11932 (N_11932,N_10827,N_10791);
and U11933 (N_11933,N_10579,N_10359);
or U11934 (N_11934,N_10018,N_10627);
nand U11935 (N_11935,N_10070,N_10394);
nor U11936 (N_11936,N_10772,N_10958);
xnor U11937 (N_11937,N_10465,N_10980);
and U11938 (N_11938,N_10479,N_10737);
and U11939 (N_11939,N_10007,N_10667);
or U11940 (N_11940,N_10249,N_10239);
nand U11941 (N_11941,N_10800,N_10686);
xor U11942 (N_11942,N_10717,N_10734);
nand U11943 (N_11943,N_10805,N_10991);
nand U11944 (N_11944,N_10083,N_10794);
nor U11945 (N_11945,N_10361,N_10970);
and U11946 (N_11946,N_10805,N_10531);
xnor U11947 (N_11947,N_10727,N_10471);
nor U11948 (N_11948,N_10469,N_10587);
or U11949 (N_11949,N_10929,N_10729);
nand U11950 (N_11950,N_10019,N_10074);
nand U11951 (N_11951,N_10158,N_10862);
and U11952 (N_11952,N_10512,N_10990);
xor U11953 (N_11953,N_10921,N_10036);
or U11954 (N_11954,N_10268,N_10804);
or U11955 (N_11955,N_10372,N_10390);
nor U11956 (N_11956,N_10480,N_10163);
or U11957 (N_11957,N_10009,N_10275);
nand U11958 (N_11958,N_10633,N_10306);
or U11959 (N_11959,N_10750,N_10725);
nand U11960 (N_11960,N_10398,N_10905);
nor U11961 (N_11961,N_10360,N_10702);
nor U11962 (N_11962,N_10115,N_10454);
nand U11963 (N_11963,N_10000,N_10839);
nand U11964 (N_11964,N_10123,N_10471);
or U11965 (N_11965,N_10361,N_10586);
xnor U11966 (N_11966,N_10471,N_10894);
nor U11967 (N_11967,N_10597,N_10936);
and U11968 (N_11968,N_10085,N_10725);
nand U11969 (N_11969,N_10544,N_10711);
nor U11970 (N_11970,N_10959,N_10062);
or U11971 (N_11971,N_10337,N_10470);
or U11972 (N_11972,N_10666,N_10012);
nand U11973 (N_11973,N_10372,N_10114);
and U11974 (N_11974,N_10161,N_10896);
and U11975 (N_11975,N_10544,N_10954);
xnor U11976 (N_11976,N_10503,N_10374);
or U11977 (N_11977,N_10924,N_10049);
nor U11978 (N_11978,N_10491,N_10587);
or U11979 (N_11979,N_10519,N_10898);
nor U11980 (N_11980,N_10005,N_10507);
nand U11981 (N_11981,N_10470,N_10370);
nor U11982 (N_11982,N_10490,N_10256);
and U11983 (N_11983,N_10868,N_10268);
or U11984 (N_11984,N_10398,N_10209);
nor U11985 (N_11985,N_10733,N_10797);
or U11986 (N_11986,N_10157,N_10334);
or U11987 (N_11987,N_10396,N_10831);
xnor U11988 (N_11988,N_10786,N_10873);
nand U11989 (N_11989,N_10932,N_10614);
and U11990 (N_11990,N_10935,N_10733);
nand U11991 (N_11991,N_10913,N_10876);
and U11992 (N_11992,N_10899,N_10343);
nand U11993 (N_11993,N_10880,N_10551);
or U11994 (N_11994,N_10428,N_10183);
or U11995 (N_11995,N_10259,N_10804);
and U11996 (N_11996,N_10475,N_10172);
and U11997 (N_11997,N_10044,N_10192);
nor U11998 (N_11998,N_10582,N_10090);
or U11999 (N_11999,N_10995,N_10562);
and U12000 (N_12000,N_11515,N_11697);
or U12001 (N_12001,N_11488,N_11689);
and U12002 (N_12002,N_11586,N_11838);
or U12003 (N_12003,N_11897,N_11217);
and U12004 (N_12004,N_11195,N_11019);
and U12005 (N_12005,N_11245,N_11623);
nand U12006 (N_12006,N_11320,N_11328);
or U12007 (N_12007,N_11249,N_11125);
and U12008 (N_12008,N_11531,N_11762);
nor U12009 (N_12009,N_11828,N_11085);
or U12010 (N_12010,N_11244,N_11717);
or U12011 (N_12011,N_11778,N_11734);
nor U12012 (N_12012,N_11648,N_11731);
and U12013 (N_12013,N_11312,N_11463);
nand U12014 (N_12014,N_11390,N_11363);
nand U12015 (N_12015,N_11696,N_11012);
and U12016 (N_12016,N_11445,N_11402);
or U12017 (N_12017,N_11609,N_11637);
xor U12018 (N_12018,N_11846,N_11517);
and U12019 (N_12019,N_11995,N_11391);
nor U12020 (N_12020,N_11510,N_11535);
or U12021 (N_12021,N_11679,N_11880);
nand U12022 (N_12022,N_11822,N_11694);
nand U12023 (N_12023,N_11285,N_11074);
nor U12024 (N_12024,N_11016,N_11505);
nand U12025 (N_12025,N_11111,N_11824);
xnor U12026 (N_12026,N_11765,N_11157);
and U12027 (N_12027,N_11304,N_11108);
nand U12028 (N_12028,N_11053,N_11169);
nor U12029 (N_12029,N_11769,N_11842);
or U12030 (N_12030,N_11819,N_11025);
nor U12031 (N_12031,N_11232,N_11314);
or U12032 (N_12032,N_11130,N_11932);
nand U12033 (N_12033,N_11851,N_11375);
nand U12034 (N_12034,N_11110,N_11829);
xor U12035 (N_12035,N_11761,N_11103);
nor U12036 (N_12036,N_11844,N_11072);
or U12037 (N_12037,N_11212,N_11567);
nor U12038 (N_12038,N_11136,N_11707);
nor U12039 (N_12039,N_11092,N_11729);
nor U12040 (N_12040,N_11224,N_11268);
xnor U12041 (N_12041,N_11216,N_11049);
xor U12042 (N_12042,N_11321,N_11643);
or U12043 (N_12043,N_11754,N_11413);
or U12044 (N_12044,N_11953,N_11023);
or U12045 (N_12045,N_11832,N_11070);
and U12046 (N_12046,N_11907,N_11471);
or U12047 (N_12047,N_11068,N_11554);
nand U12048 (N_12048,N_11067,N_11758);
or U12049 (N_12049,N_11161,N_11766);
or U12050 (N_12050,N_11459,N_11789);
or U12051 (N_12051,N_11594,N_11972);
nor U12052 (N_12052,N_11360,N_11090);
nand U12053 (N_12053,N_11214,N_11941);
xnor U12054 (N_12054,N_11931,N_11954);
xor U12055 (N_12055,N_11200,N_11845);
or U12056 (N_12056,N_11010,N_11276);
nor U12057 (N_12057,N_11102,N_11760);
and U12058 (N_12058,N_11836,N_11676);
nor U12059 (N_12059,N_11383,N_11509);
nor U12060 (N_12060,N_11142,N_11007);
nand U12061 (N_12061,N_11477,N_11563);
or U12062 (N_12062,N_11750,N_11981);
nor U12063 (N_12063,N_11475,N_11978);
nor U12064 (N_12064,N_11324,N_11065);
nor U12065 (N_12065,N_11417,N_11179);
nor U12066 (N_12066,N_11456,N_11184);
xnor U12067 (N_12067,N_11549,N_11300);
or U12068 (N_12068,N_11211,N_11529);
or U12069 (N_12069,N_11129,N_11794);
nor U12070 (N_12070,N_11776,N_11120);
nor U12071 (N_12071,N_11665,N_11308);
nand U12072 (N_12072,N_11343,N_11044);
xnor U12073 (N_12073,N_11578,N_11809);
nor U12074 (N_12074,N_11124,N_11787);
nand U12075 (N_12075,N_11935,N_11154);
and U12076 (N_12076,N_11668,N_11749);
xor U12077 (N_12077,N_11831,N_11796);
nor U12078 (N_12078,N_11958,N_11163);
nor U12079 (N_12079,N_11550,N_11864);
nand U12080 (N_12080,N_11334,N_11654);
nor U12081 (N_12081,N_11234,N_11647);
and U12082 (N_12082,N_11774,N_11674);
nand U12083 (N_12083,N_11626,N_11024);
or U12084 (N_12084,N_11925,N_11979);
and U12085 (N_12085,N_11620,N_11266);
nor U12086 (N_12086,N_11411,N_11716);
or U12087 (N_12087,N_11345,N_11660);
and U12088 (N_12088,N_11943,N_11407);
nor U12089 (N_12089,N_11060,N_11558);
xnor U12090 (N_12090,N_11847,N_11933);
xnor U12091 (N_12091,N_11858,N_11562);
xnor U12092 (N_12092,N_11143,N_11898);
xor U12093 (N_12093,N_11265,N_11811);
xor U12094 (N_12094,N_11015,N_11171);
and U12095 (N_12095,N_11893,N_11923);
nor U12096 (N_12096,N_11569,N_11570);
nand U12097 (N_12097,N_11737,N_11657);
xnor U12098 (N_12098,N_11152,N_11231);
nand U12099 (N_12099,N_11104,N_11084);
xnor U12100 (N_12100,N_11975,N_11087);
nor U12101 (N_12101,N_11455,N_11856);
nor U12102 (N_12102,N_11722,N_11326);
nor U12103 (N_12103,N_11080,N_11681);
xnor U12104 (N_12104,N_11307,N_11180);
nor U12105 (N_12105,N_11297,N_11850);
nor U12106 (N_12106,N_11219,N_11046);
nor U12107 (N_12107,N_11501,N_11703);
xor U12108 (N_12108,N_11122,N_11038);
and U12109 (N_12109,N_11521,N_11624);
and U12110 (N_12110,N_11977,N_11823);
and U12111 (N_12111,N_11281,N_11377);
nor U12112 (N_12112,N_11194,N_11058);
and U12113 (N_12113,N_11480,N_11610);
and U12114 (N_12114,N_11011,N_11983);
nand U12115 (N_12115,N_11651,N_11453);
nor U12116 (N_12116,N_11430,N_11653);
xnor U12117 (N_12117,N_11645,N_11951);
or U12118 (N_12118,N_11803,N_11534);
nand U12119 (N_12119,N_11584,N_11193);
and U12120 (N_12120,N_11565,N_11223);
or U12121 (N_12121,N_11040,N_11793);
or U12122 (N_12122,N_11711,N_11618);
nand U12123 (N_12123,N_11773,N_11047);
nand U12124 (N_12124,N_11001,N_11539);
nor U12125 (N_12125,N_11944,N_11885);
and U12126 (N_12126,N_11246,N_11474);
nand U12127 (N_12127,N_11272,N_11018);
and U12128 (N_12128,N_11573,N_11118);
nand U12129 (N_12129,N_11270,N_11917);
nor U12130 (N_12130,N_11107,N_11863);
nor U12131 (N_12131,N_11661,N_11890);
xnor U12132 (N_12132,N_11870,N_11968);
or U12133 (N_12133,N_11177,N_11814);
nor U12134 (N_12134,N_11976,N_11128);
nand U12135 (N_12135,N_11601,N_11699);
nand U12136 (N_12136,N_11017,N_11994);
nand U12137 (N_12137,N_11640,N_11867);
or U12138 (N_12138,N_11834,N_11387);
and U12139 (N_12139,N_11054,N_11079);
or U12140 (N_12140,N_11915,N_11380);
or U12141 (N_12141,N_11155,N_11914);
or U12142 (N_12142,N_11993,N_11205);
or U12143 (N_12143,N_11006,N_11848);
nand U12144 (N_12144,N_11020,N_11512);
and U12145 (N_12145,N_11405,N_11013);
or U12146 (N_12146,N_11322,N_11239);
xnor U12147 (N_12147,N_11371,N_11685);
and U12148 (N_12148,N_11868,N_11790);
xnor U12149 (N_12149,N_11949,N_11162);
or U12150 (N_12150,N_11482,N_11538);
nor U12151 (N_12151,N_11327,N_11394);
nand U12152 (N_12152,N_11422,N_11818);
nand U12153 (N_12153,N_11255,N_11302);
xnor U12154 (N_12154,N_11997,N_11805);
or U12155 (N_12155,N_11613,N_11004);
xnor U12156 (N_12156,N_11593,N_11396);
xnor U12157 (N_12157,N_11595,N_11784);
nor U12158 (N_12158,N_11582,N_11088);
and U12159 (N_12159,N_11305,N_11221);
xor U12160 (N_12160,N_11421,N_11415);
xor U12161 (N_12161,N_11034,N_11202);
nand U12162 (N_12162,N_11469,N_11615);
and U12163 (N_12163,N_11775,N_11050);
and U12164 (N_12164,N_11262,N_11678);
and U12165 (N_12165,N_11030,N_11437);
nor U12166 (N_12166,N_11936,N_11833);
nor U12167 (N_12167,N_11132,N_11319);
and U12168 (N_12168,N_11695,N_11081);
and U12169 (N_12169,N_11075,N_11166);
xor U12170 (N_12170,N_11197,N_11311);
nor U12171 (N_12171,N_11635,N_11918);
nand U12172 (N_12172,N_11806,N_11884);
nor U12173 (N_12173,N_11188,N_11490);
or U12174 (N_12174,N_11743,N_11514);
and U12175 (N_12175,N_11920,N_11346);
and U12176 (N_12176,N_11447,N_11701);
nor U12177 (N_12177,N_11106,N_11959);
nor U12178 (N_12178,N_11622,N_11359);
nand U12179 (N_12179,N_11964,N_11274);
nand U12180 (N_12180,N_11423,N_11191);
and U12181 (N_12181,N_11029,N_11499);
xnor U12182 (N_12182,N_11506,N_11516);
xor U12183 (N_12183,N_11662,N_11659);
and U12184 (N_12184,N_11031,N_11057);
nand U12185 (N_12185,N_11233,N_11768);
or U12186 (N_12186,N_11650,N_11256);
xor U12187 (N_12187,N_11435,N_11332);
and U12188 (N_12188,N_11633,N_11099);
nor U12189 (N_12189,N_11061,N_11289);
nand U12190 (N_12190,N_11418,N_11753);
or U12191 (N_12191,N_11980,N_11349);
and U12192 (N_12192,N_11795,N_11508);
or U12193 (N_12193,N_11644,N_11439);
nand U12194 (N_12194,N_11082,N_11782);
or U12195 (N_12195,N_11882,N_11204);
xor U12196 (N_12196,N_11687,N_11638);
nor U12197 (N_12197,N_11684,N_11062);
nand U12198 (N_12198,N_11617,N_11614);
or U12199 (N_12199,N_11780,N_11114);
xor U12200 (N_12200,N_11339,N_11649);
xor U12201 (N_12201,N_11298,N_11741);
and U12202 (N_12202,N_11816,N_11258);
nor U12203 (N_12203,N_11370,N_11952);
and U12204 (N_12204,N_11399,N_11874);
and U12205 (N_12205,N_11817,N_11379);
and U12206 (N_12206,N_11263,N_11472);
nor U12207 (N_12207,N_11369,N_11059);
or U12208 (N_12208,N_11666,N_11454);
nand U12209 (N_12209,N_11800,N_11872);
or U12210 (N_12210,N_11519,N_11781);
or U12211 (N_12211,N_11408,N_11928);
or U12212 (N_12212,N_11916,N_11014);
nand U12213 (N_12213,N_11912,N_11998);
and U12214 (N_12214,N_11160,N_11756);
nor U12215 (N_12215,N_11619,N_11492);
nand U12216 (N_12216,N_11990,N_11295);
or U12217 (N_12217,N_11966,N_11576);
nand U12218 (N_12218,N_11876,N_11350);
nand U12219 (N_12219,N_11574,N_11937);
or U12220 (N_12220,N_11473,N_11725);
nand U12221 (N_12221,N_11902,N_11543);
and U12222 (N_12222,N_11172,N_11428);
nand U12223 (N_12223,N_11094,N_11198);
nand U12224 (N_12224,N_11807,N_11755);
xor U12225 (N_12225,N_11486,N_11260);
and U12226 (N_12226,N_11672,N_11548);
or U12227 (N_12227,N_11680,N_11939);
or U12228 (N_12228,N_11227,N_11409);
and U12229 (N_12229,N_11218,N_11176);
nand U12230 (N_12230,N_11804,N_11942);
and U12231 (N_12231,N_11207,N_11904);
xor U12232 (N_12232,N_11201,N_11236);
and U12233 (N_12233,N_11967,N_11628);
nand U12234 (N_12234,N_11228,N_11746);
or U12235 (N_12235,N_11283,N_11905);
nand U12236 (N_12236,N_11173,N_11727);
nor U12237 (N_12237,N_11287,N_11692);
nand U12238 (N_12238,N_11945,N_11724);
nand U12239 (N_12239,N_11602,N_11098);
nor U12240 (N_12240,N_11403,N_11271);
xnor U12241 (N_12241,N_11785,N_11895);
nand U12242 (N_12242,N_11852,N_11210);
nand U12243 (N_12243,N_11779,N_11636);
xnor U12244 (N_12244,N_11608,N_11841);
xor U12245 (N_12245,N_11987,N_11675);
and U12246 (N_12246,N_11446,N_11306);
nor U12247 (N_12247,N_11443,N_11713);
or U12248 (N_12248,N_11877,N_11797);
xnor U12249 (N_12249,N_11606,N_11362);
and U12250 (N_12250,N_11751,N_11721);
nor U12251 (N_12251,N_11434,N_11185);
nand U12252 (N_12252,N_11384,N_11052);
and U12253 (N_12253,N_11386,N_11865);
xor U12254 (N_12254,N_11892,N_11487);
xnor U12255 (N_12255,N_11996,N_11181);
nor U12256 (N_12256,N_11929,N_11461);
or U12257 (N_12257,N_11551,N_11131);
or U12258 (N_12258,N_11891,N_11427);
or U12259 (N_12259,N_11000,N_11752);
nor U12260 (N_12260,N_11373,N_11559);
and U12261 (N_12261,N_11083,N_11267);
nand U12262 (N_12262,N_11432,N_11237);
or U12263 (N_12263,N_11688,N_11259);
nand U12264 (N_12264,N_11464,N_11045);
nor U12265 (N_12265,N_11078,N_11280);
and U12266 (N_12266,N_11424,N_11495);
and U12267 (N_12267,N_11553,N_11433);
nor U12268 (N_12268,N_11385,N_11389);
nor U12269 (N_12269,N_11127,N_11008);
or U12270 (N_12270,N_11686,N_11333);
or U12271 (N_12271,N_11329,N_11632);
xnor U12272 (N_12272,N_11147,N_11801);
nand U12273 (N_12273,N_11726,N_11148);
xor U12274 (N_12274,N_11604,N_11041);
and U12275 (N_12275,N_11159,N_11957);
nand U12276 (N_12276,N_11862,N_11973);
nor U12277 (N_12277,N_11658,N_11372);
and U12278 (N_12278,N_11922,N_11572);
nor U12279 (N_12279,N_11340,N_11507);
nor U12280 (N_12280,N_11664,N_11027);
xor U12281 (N_12281,N_11174,N_11264);
nor U12282 (N_12282,N_11698,N_11069);
or U12283 (N_12283,N_11144,N_11589);
and U12284 (N_12284,N_11886,N_11183);
nand U12285 (N_12285,N_11431,N_11926);
nor U12286 (N_12286,N_11605,N_11927);
or U12287 (N_12287,N_11225,N_11991);
nor U12288 (N_12288,N_11580,N_11100);
nand U12289 (N_12289,N_11542,N_11291);
nor U12290 (N_12290,N_11603,N_11557);
xnor U12291 (N_12291,N_11896,N_11444);
and U12292 (N_12292,N_11873,N_11241);
nand U12293 (N_12293,N_11468,N_11420);
xnor U12294 (N_12294,N_11064,N_11470);
and U12295 (N_12295,N_11467,N_11894);
nor U12296 (N_12296,N_11733,N_11235);
nand U12297 (N_12297,N_11460,N_11073);
nor U12298 (N_12298,N_11700,N_11331);
nand U12299 (N_12299,N_11043,N_11416);
and U12300 (N_12300,N_11119,N_11577);
nor U12301 (N_12301,N_11076,N_11401);
and U12302 (N_12302,N_11536,N_11693);
or U12303 (N_12303,N_11527,N_11251);
nor U12304 (N_12304,N_11187,N_11513);
nand U12305 (N_12305,N_11117,N_11330);
nand U12306 (N_12306,N_11440,N_11310);
nand U12307 (N_12307,N_11960,N_11382);
nand U12308 (N_12308,N_11048,N_11625);
and U12309 (N_12309,N_11764,N_11419);
or U12310 (N_12310,N_11849,N_11367);
nor U12311 (N_12311,N_11887,N_11066);
xor U12312 (N_12312,N_11631,N_11560);
nor U12313 (N_12313,N_11156,N_11376);
nor U12314 (N_12314,N_11909,N_11277);
or U12315 (N_12315,N_11133,N_11579);
and U12316 (N_12316,N_11655,N_11571);
and U12317 (N_12317,N_11598,N_11101);
or U12318 (N_12318,N_11134,N_11581);
nand U12319 (N_12319,N_11229,N_11940);
or U12320 (N_12320,N_11400,N_11338);
and U12321 (N_12321,N_11575,N_11466);
nor U12322 (N_12322,N_11555,N_11528);
and U12323 (N_12323,N_11532,N_11190);
nand U12324 (N_12324,N_11511,N_11410);
and U12325 (N_12325,N_11253,N_11121);
or U12326 (N_12326,N_11189,N_11151);
nand U12327 (N_12327,N_11425,N_11113);
or U12328 (N_12328,N_11999,N_11491);
nand U12329 (N_12329,N_11351,N_11381);
xnor U12330 (N_12330,N_11854,N_11203);
nor U12331 (N_12331,N_11730,N_11323);
or U12332 (N_12332,N_11222,N_11629);
xnor U12333 (N_12333,N_11641,N_11961);
and U12334 (N_12334,N_11767,N_11723);
nand U12335 (N_12335,N_11465,N_11748);
or U12336 (N_12336,N_11525,N_11533);
or U12337 (N_12337,N_11436,N_11597);
nand U12338 (N_12338,N_11522,N_11962);
nor U12339 (N_12339,N_11518,N_11950);
nand U12340 (N_12340,N_11093,N_11970);
nand U12341 (N_12341,N_11705,N_11158);
and U12342 (N_12342,N_11071,N_11690);
and U12343 (N_12343,N_11670,N_11969);
nand U12344 (N_12344,N_11502,N_11826);
nand U12345 (N_12345,N_11252,N_11042);
nor U12346 (N_12346,N_11164,N_11663);
xor U12347 (N_12347,N_11039,N_11985);
or U12348 (N_12348,N_11357,N_11303);
nor U12349 (N_12349,N_11313,N_11520);
and U12350 (N_12350,N_11881,N_11496);
nor U12351 (N_12351,N_11747,N_11347);
nand U12352 (N_12352,N_11537,N_11992);
nor U12353 (N_12353,N_11546,N_11984);
nand U12354 (N_12354,N_11206,N_11908);
and U12355 (N_12355,N_11911,N_11588);
and U12356 (N_12356,N_11612,N_11630);
xor U12357 (N_12357,N_11783,N_11002);
nor U12358 (N_12358,N_11667,N_11165);
nor U12359 (N_12359,N_11116,N_11745);
xnor U12360 (N_12360,N_11462,N_11974);
nand U12361 (N_12361,N_11378,N_11392);
xnor U12362 (N_12362,N_11859,N_11627);
nand U12363 (N_12363,N_11820,N_11438);
or U12364 (N_12364,N_11564,N_11352);
nor U12365 (N_12365,N_11247,N_11028);
nor U12366 (N_12366,N_11250,N_11368);
or U12367 (N_12367,N_11450,N_11607);
nor U12368 (N_12368,N_11494,N_11033);
xnor U12369 (N_12369,N_11899,N_11592);
xor U12370 (N_12370,N_11137,N_11036);
xnor U12371 (N_12371,N_11903,N_11683);
nand U12372 (N_12372,N_11178,N_11839);
nand U12373 (N_12373,N_11947,N_11547);
and U12374 (N_12374,N_11294,N_11341);
nand U12375 (N_12375,N_11853,N_11772);
or U12376 (N_12376,N_11135,N_11566);
and U12377 (N_12377,N_11192,N_11673);
nor U12378 (N_12378,N_11710,N_11055);
or U12379 (N_12379,N_11540,N_11971);
xnor U12380 (N_12380,N_11485,N_11037);
nand U12381 (N_12381,N_11286,N_11702);
nor U12382 (N_12382,N_11921,N_11337);
nor U12383 (N_12383,N_11830,N_11213);
nand U12384 (N_12384,N_11889,N_11366);
or U12385 (N_12385,N_11167,N_11742);
or U12386 (N_12386,N_11835,N_11149);
or U12387 (N_12387,N_11261,N_11869);
nand U12388 (N_12388,N_11720,N_11704);
or U12389 (N_12389,N_11353,N_11348);
and U12390 (N_12390,N_11652,N_11316);
or U12391 (N_12391,N_11530,N_11948);
nand U12392 (N_12392,N_11956,N_11883);
or U12393 (N_12393,N_11738,N_11095);
xor U12394 (N_12394,N_11503,N_11709);
xnor U12395 (N_12395,N_11599,N_11600);
and U12396 (N_12396,N_11355,N_11861);
and U12397 (N_12397,N_11634,N_11282);
or U12398 (N_12398,N_11096,N_11646);
or U12399 (N_12399,N_11315,N_11523);
and U12400 (N_12400,N_11452,N_11344);
or U12401 (N_12401,N_11669,N_11293);
xnor U12402 (N_12402,N_11759,N_11799);
nand U12403 (N_12403,N_11682,N_11757);
nor U12404 (N_12404,N_11526,N_11815);
nand U12405 (N_12405,N_11788,N_11919);
nor U12406 (N_12406,N_11810,N_11051);
nor U12407 (N_12407,N_11354,N_11857);
or U12408 (N_12408,N_11364,N_11561);
or U12409 (N_12409,N_11484,N_11358);
or U12410 (N_12410,N_11196,N_11254);
nand U12411 (N_12411,N_11708,N_11552);
and U12412 (N_12412,N_11924,N_11802);
or U12413 (N_12413,N_11404,N_11005);
and U12414 (N_12414,N_11930,N_11269);
nand U12415 (N_12415,N_11112,N_11056);
xnor U12416 (N_12416,N_11226,N_11483);
nor U12417 (N_12417,N_11706,N_11813);
nor U12418 (N_12418,N_11086,N_11812);
nand U12419 (N_12419,N_11763,N_11989);
or U12420 (N_12420,N_11168,N_11825);
and U12421 (N_12421,N_11591,N_11365);
xnor U12422 (N_12422,N_11871,N_11458);
nor U12423 (N_12423,N_11003,N_11336);
or U12424 (N_12424,N_11097,N_11986);
or U12425 (N_12425,N_11022,N_11275);
or U12426 (N_12426,N_11792,N_11827);
and U12427 (N_12427,N_11318,N_11642);
nand U12428 (N_12428,N_11035,N_11317);
nand U12429 (N_12429,N_11238,N_11616);
nand U12430 (N_12430,N_11109,N_11677);
or U12431 (N_12431,N_11963,N_11639);
xnor U12432 (N_12432,N_11808,N_11442);
and U12433 (N_12433,N_11497,N_11441);
nand U12434 (N_12434,N_11278,N_11077);
nand U12435 (N_12435,N_11309,N_11296);
and U12436 (N_12436,N_11715,N_11123);
nor U12437 (N_12437,N_11821,N_11913);
or U12438 (N_12438,N_11299,N_11139);
and U12439 (N_12439,N_11938,N_11524);
or U12440 (N_12440,N_11493,N_11860);
nor U12441 (N_12441,N_11955,N_11965);
xnor U12442 (N_12442,N_11021,N_11479);
xor U12443 (N_12443,N_11843,N_11744);
or U12444 (N_12444,N_11220,N_11412);
and U12445 (N_12445,N_11791,N_11091);
nand U12446 (N_12446,N_11063,N_11449);
and U12447 (N_12447,N_11583,N_11208);
nor U12448 (N_12448,N_11946,N_11489);
and U12449 (N_12449,N_11771,N_11879);
nand U12450 (N_12450,N_11032,N_11718);
nor U12451 (N_12451,N_11585,N_11910);
nor U12452 (N_12452,N_11855,N_11182);
nor U12453 (N_12453,N_11500,N_11568);
xor U12454 (N_12454,N_11292,N_11740);
xnor U12455 (N_12455,N_11590,N_11875);
xnor U12456 (N_12456,N_11476,N_11900);
xnor U12457 (N_12457,N_11215,N_11279);
xnor U12458 (N_12458,N_11393,N_11089);
or U12459 (N_12459,N_11356,N_11199);
and U12460 (N_12460,N_11798,N_11478);
and U12461 (N_12461,N_11451,N_11395);
nor U12462 (N_12462,N_11712,N_11209);
and U12463 (N_12463,N_11342,N_11170);
and U12464 (N_12464,N_11325,N_11374);
or U12465 (N_12465,N_11026,N_11284);
or U12466 (N_12466,N_11240,N_11736);
nor U12467 (N_12467,N_11248,N_11429);
or U12468 (N_12468,N_11115,N_11388);
or U12469 (N_12469,N_11126,N_11786);
or U12470 (N_12470,N_11732,N_11719);
nor U12471 (N_12471,N_11596,N_11288);
nor U12472 (N_12472,N_11691,N_11426);
nand U12473 (N_12473,N_11397,N_11878);
xor U12474 (N_12474,N_11541,N_11301);
or U12475 (N_12475,N_11545,N_11105);
nor U12476 (N_12476,N_11257,N_11739);
nor U12477 (N_12477,N_11587,N_11145);
xor U12478 (N_12478,N_11406,N_11906);
nor U12479 (N_12479,N_11138,N_11398);
nor U12480 (N_12480,N_11457,N_11009);
xor U12481 (N_12481,N_11728,N_11621);
nor U12482 (N_12482,N_11735,N_11611);
xor U12483 (N_12483,N_11481,N_11498);
xnor U12484 (N_12484,N_11141,N_11671);
or U12485 (N_12485,N_11175,N_11242);
xor U12486 (N_12486,N_11290,N_11777);
or U12487 (N_12487,N_11335,N_11150);
or U12488 (N_12488,N_11770,N_11243);
nand U12489 (N_12489,N_11544,N_11888);
xor U12490 (N_12490,N_11866,N_11186);
or U12491 (N_12491,N_11934,N_11556);
nor U12492 (N_12492,N_11153,N_11448);
nor U12493 (N_12493,N_11837,N_11146);
nor U12494 (N_12494,N_11656,N_11714);
nor U12495 (N_12495,N_11901,N_11840);
nor U12496 (N_12496,N_11361,N_11414);
and U12497 (N_12497,N_11504,N_11988);
and U12498 (N_12498,N_11230,N_11140);
nand U12499 (N_12499,N_11982,N_11273);
nor U12500 (N_12500,N_11568,N_11304);
nor U12501 (N_12501,N_11381,N_11991);
and U12502 (N_12502,N_11055,N_11241);
nor U12503 (N_12503,N_11649,N_11514);
xor U12504 (N_12504,N_11368,N_11739);
nand U12505 (N_12505,N_11283,N_11287);
xor U12506 (N_12506,N_11470,N_11327);
nor U12507 (N_12507,N_11169,N_11982);
xor U12508 (N_12508,N_11679,N_11773);
nand U12509 (N_12509,N_11310,N_11824);
or U12510 (N_12510,N_11331,N_11929);
nand U12511 (N_12511,N_11374,N_11762);
nor U12512 (N_12512,N_11221,N_11563);
or U12513 (N_12513,N_11516,N_11052);
xnor U12514 (N_12514,N_11759,N_11592);
nor U12515 (N_12515,N_11627,N_11995);
nand U12516 (N_12516,N_11138,N_11179);
nand U12517 (N_12517,N_11686,N_11171);
xnor U12518 (N_12518,N_11316,N_11493);
nor U12519 (N_12519,N_11896,N_11750);
and U12520 (N_12520,N_11173,N_11806);
or U12521 (N_12521,N_11529,N_11466);
or U12522 (N_12522,N_11770,N_11876);
or U12523 (N_12523,N_11861,N_11525);
or U12524 (N_12524,N_11606,N_11818);
nand U12525 (N_12525,N_11582,N_11776);
nor U12526 (N_12526,N_11151,N_11508);
xor U12527 (N_12527,N_11622,N_11831);
nor U12528 (N_12528,N_11819,N_11253);
and U12529 (N_12529,N_11853,N_11584);
and U12530 (N_12530,N_11555,N_11855);
nor U12531 (N_12531,N_11254,N_11690);
or U12532 (N_12532,N_11133,N_11115);
nor U12533 (N_12533,N_11481,N_11467);
and U12534 (N_12534,N_11495,N_11779);
xor U12535 (N_12535,N_11231,N_11692);
and U12536 (N_12536,N_11219,N_11201);
or U12537 (N_12537,N_11057,N_11998);
nor U12538 (N_12538,N_11994,N_11982);
and U12539 (N_12539,N_11161,N_11866);
xor U12540 (N_12540,N_11918,N_11312);
nor U12541 (N_12541,N_11538,N_11792);
xor U12542 (N_12542,N_11498,N_11786);
nand U12543 (N_12543,N_11069,N_11874);
nand U12544 (N_12544,N_11996,N_11174);
nand U12545 (N_12545,N_11446,N_11410);
nand U12546 (N_12546,N_11829,N_11407);
or U12547 (N_12547,N_11225,N_11818);
or U12548 (N_12548,N_11219,N_11424);
xnor U12549 (N_12549,N_11682,N_11905);
or U12550 (N_12550,N_11665,N_11890);
xor U12551 (N_12551,N_11076,N_11590);
xnor U12552 (N_12552,N_11060,N_11914);
xor U12553 (N_12553,N_11612,N_11678);
and U12554 (N_12554,N_11977,N_11633);
or U12555 (N_12555,N_11468,N_11252);
nand U12556 (N_12556,N_11792,N_11181);
xnor U12557 (N_12557,N_11612,N_11910);
nor U12558 (N_12558,N_11932,N_11552);
xnor U12559 (N_12559,N_11797,N_11970);
or U12560 (N_12560,N_11131,N_11614);
nand U12561 (N_12561,N_11411,N_11114);
nor U12562 (N_12562,N_11396,N_11727);
nand U12563 (N_12563,N_11775,N_11310);
xor U12564 (N_12564,N_11737,N_11644);
nand U12565 (N_12565,N_11543,N_11576);
and U12566 (N_12566,N_11150,N_11434);
nor U12567 (N_12567,N_11703,N_11527);
nand U12568 (N_12568,N_11206,N_11894);
or U12569 (N_12569,N_11926,N_11738);
nor U12570 (N_12570,N_11639,N_11818);
or U12571 (N_12571,N_11283,N_11223);
xnor U12572 (N_12572,N_11440,N_11535);
xnor U12573 (N_12573,N_11119,N_11591);
or U12574 (N_12574,N_11827,N_11629);
nor U12575 (N_12575,N_11356,N_11505);
or U12576 (N_12576,N_11027,N_11610);
or U12577 (N_12577,N_11639,N_11438);
or U12578 (N_12578,N_11246,N_11665);
xnor U12579 (N_12579,N_11130,N_11935);
nand U12580 (N_12580,N_11831,N_11259);
or U12581 (N_12581,N_11301,N_11083);
nor U12582 (N_12582,N_11512,N_11361);
nor U12583 (N_12583,N_11782,N_11109);
nor U12584 (N_12584,N_11098,N_11464);
or U12585 (N_12585,N_11778,N_11615);
nor U12586 (N_12586,N_11939,N_11398);
or U12587 (N_12587,N_11958,N_11847);
xnor U12588 (N_12588,N_11049,N_11522);
nand U12589 (N_12589,N_11083,N_11130);
or U12590 (N_12590,N_11251,N_11379);
and U12591 (N_12591,N_11341,N_11028);
nand U12592 (N_12592,N_11546,N_11723);
and U12593 (N_12593,N_11285,N_11208);
or U12594 (N_12594,N_11490,N_11081);
nor U12595 (N_12595,N_11499,N_11406);
and U12596 (N_12596,N_11126,N_11485);
and U12597 (N_12597,N_11770,N_11554);
or U12598 (N_12598,N_11514,N_11741);
xor U12599 (N_12599,N_11425,N_11458);
nand U12600 (N_12600,N_11415,N_11943);
xnor U12601 (N_12601,N_11230,N_11570);
nor U12602 (N_12602,N_11029,N_11846);
nand U12603 (N_12603,N_11503,N_11980);
nand U12604 (N_12604,N_11095,N_11473);
and U12605 (N_12605,N_11586,N_11376);
xor U12606 (N_12606,N_11871,N_11546);
nor U12607 (N_12607,N_11580,N_11829);
nand U12608 (N_12608,N_11503,N_11322);
nor U12609 (N_12609,N_11667,N_11118);
nand U12610 (N_12610,N_11269,N_11015);
nand U12611 (N_12611,N_11008,N_11548);
nand U12612 (N_12612,N_11822,N_11437);
and U12613 (N_12613,N_11510,N_11560);
or U12614 (N_12614,N_11122,N_11332);
nor U12615 (N_12615,N_11047,N_11573);
and U12616 (N_12616,N_11793,N_11765);
xor U12617 (N_12617,N_11378,N_11190);
or U12618 (N_12618,N_11251,N_11684);
or U12619 (N_12619,N_11232,N_11372);
and U12620 (N_12620,N_11322,N_11738);
nand U12621 (N_12621,N_11526,N_11497);
and U12622 (N_12622,N_11889,N_11435);
nand U12623 (N_12623,N_11035,N_11750);
nand U12624 (N_12624,N_11822,N_11014);
xor U12625 (N_12625,N_11229,N_11117);
and U12626 (N_12626,N_11291,N_11937);
nand U12627 (N_12627,N_11781,N_11054);
nor U12628 (N_12628,N_11971,N_11313);
xnor U12629 (N_12629,N_11797,N_11680);
and U12630 (N_12630,N_11046,N_11277);
nand U12631 (N_12631,N_11916,N_11544);
nand U12632 (N_12632,N_11396,N_11253);
or U12633 (N_12633,N_11574,N_11228);
xor U12634 (N_12634,N_11868,N_11343);
xnor U12635 (N_12635,N_11418,N_11118);
nand U12636 (N_12636,N_11668,N_11123);
xor U12637 (N_12637,N_11653,N_11381);
and U12638 (N_12638,N_11938,N_11074);
nand U12639 (N_12639,N_11808,N_11190);
nand U12640 (N_12640,N_11703,N_11451);
nor U12641 (N_12641,N_11365,N_11636);
nand U12642 (N_12642,N_11595,N_11941);
nor U12643 (N_12643,N_11815,N_11613);
nor U12644 (N_12644,N_11636,N_11866);
xnor U12645 (N_12645,N_11309,N_11083);
and U12646 (N_12646,N_11794,N_11195);
xnor U12647 (N_12647,N_11339,N_11096);
xnor U12648 (N_12648,N_11868,N_11779);
or U12649 (N_12649,N_11758,N_11999);
or U12650 (N_12650,N_11939,N_11735);
and U12651 (N_12651,N_11421,N_11521);
nor U12652 (N_12652,N_11506,N_11852);
xnor U12653 (N_12653,N_11972,N_11937);
nand U12654 (N_12654,N_11696,N_11667);
nand U12655 (N_12655,N_11394,N_11107);
nor U12656 (N_12656,N_11807,N_11736);
and U12657 (N_12657,N_11805,N_11613);
or U12658 (N_12658,N_11082,N_11030);
and U12659 (N_12659,N_11990,N_11742);
or U12660 (N_12660,N_11046,N_11711);
xor U12661 (N_12661,N_11549,N_11251);
xor U12662 (N_12662,N_11666,N_11171);
and U12663 (N_12663,N_11168,N_11229);
and U12664 (N_12664,N_11300,N_11781);
and U12665 (N_12665,N_11555,N_11306);
nand U12666 (N_12666,N_11663,N_11500);
nand U12667 (N_12667,N_11586,N_11661);
nand U12668 (N_12668,N_11869,N_11583);
or U12669 (N_12669,N_11641,N_11647);
nand U12670 (N_12670,N_11624,N_11484);
or U12671 (N_12671,N_11213,N_11336);
nor U12672 (N_12672,N_11089,N_11991);
xnor U12673 (N_12673,N_11145,N_11578);
or U12674 (N_12674,N_11689,N_11998);
and U12675 (N_12675,N_11391,N_11465);
nor U12676 (N_12676,N_11665,N_11723);
or U12677 (N_12677,N_11445,N_11890);
or U12678 (N_12678,N_11963,N_11888);
or U12679 (N_12679,N_11477,N_11038);
nand U12680 (N_12680,N_11812,N_11036);
nand U12681 (N_12681,N_11009,N_11639);
or U12682 (N_12682,N_11294,N_11691);
nand U12683 (N_12683,N_11291,N_11633);
nor U12684 (N_12684,N_11310,N_11402);
and U12685 (N_12685,N_11649,N_11460);
or U12686 (N_12686,N_11257,N_11194);
nor U12687 (N_12687,N_11773,N_11950);
nor U12688 (N_12688,N_11112,N_11365);
nand U12689 (N_12689,N_11717,N_11680);
or U12690 (N_12690,N_11876,N_11990);
nand U12691 (N_12691,N_11968,N_11853);
nand U12692 (N_12692,N_11013,N_11091);
xnor U12693 (N_12693,N_11349,N_11375);
or U12694 (N_12694,N_11296,N_11256);
nand U12695 (N_12695,N_11203,N_11938);
or U12696 (N_12696,N_11239,N_11183);
or U12697 (N_12697,N_11689,N_11383);
xnor U12698 (N_12698,N_11742,N_11563);
nand U12699 (N_12699,N_11655,N_11401);
or U12700 (N_12700,N_11652,N_11767);
xor U12701 (N_12701,N_11184,N_11987);
nand U12702 (N_12702,N_11063,N_11219);
nor U12703 (N_12703,N_11311,N_11383);
nand U12704 (N_12704,N_11096,N_11658);
xor U12705 (N_12705,N_11315,N_11567);
nand U12706 (N_12706,N_11146,N_11830);
xor U12707 (N_12707,N_11947,N_11010);
nor U12708 (N_12708,N_11406,N_11486);
nor U12709 (N_12709,N_11540,N_11360);
nor U12710 (N_12710,N_11753,N_11790);
nand U12711 (N_12711,N_11632,N_11073);
nand U12712 (N_12712,N_11218,N_11987);
and U12713 (N_12713,N_11868,N_11757);
nand U12714 (N_12714,N_11974,N_11803);
nand U12715 (N_12715,N_11797,N_11532);
and U12716 (N_12716,N_11205,N_11445);
nor U12717 (N_12717,N_11037,N_11683);
xor U12718 (N_12718,N_11016,N_11282);
and U12719 (N_12719,N_11521,N_11155);
or U12720 (N_12720,N_11451,N_11366);
nand U12721 (N_12721,N_11550,N_11809);
and U12722 (N_12722,N_11541,N_11863);
and U12723 (N_12723,N_11541,N_11166);
or U12724 (N_12724,N_11085,N_11131);
nor U12725 (N_12725,N_11718,N_11005);
or U12726 (N_12726,N_11819,N_11223);
or U12727 (N_12727,N_11392,N_11767);
xor U12728 (N_12728,N_11599,N_11787);
nor U12729 (N_12729,N_11081,N_11383);
and U12730 (N_12730,N_11026,N_11692);
nand U12731 (N_12731,N_11092,N_11071);
or U12732 (N_12732,N_11755,N_11173);
nor U12733 (N_12733,N_11992,N_11530);
nor U12734 (N_12734,N_11921,N_11031);
or U12735 (N_12735,N_11124,N_11088);
nand U12736 (N_12736,N_11195,N_11212);
and U12737 (N_12737,N_11410,N_11083);
nand U12738 (N_12738,N_11353,N_11250);
xor U12739 (N_12739,N_11842,N_11191);
nor U12740 (N_12740,N_11466,N_11812);
xor U12741 (N_12741,N_11627,N_11804);
nor U12742 (N_12742,N_11246,N_11927);
nand U12743 (N_12743,N_11252,N_11969);
nor U12744 (N_12744,N_11400,N_11875);
and U12745 (N_12745,N_11459,N_11465);
or U12746 (N_12746,N_11172,N_11472);
nor U12747 (N_12747,N_11186,N_11996);
nor U12748 (N_12748,N_11977,N_11488);
xnor U12749 (N_12749,N_11810,N_11533);
nor U12750 (N_12750,N_11717,N_11768);
or U12751 (N_12751,N_11088,N_11995);
xnor U12752 (N_12752,N_11102,N_11522);
nand U12753 (N_12753,N_11766,N_11877);
and U12754 (N_12754,N_11831,N_11846);
nor U12755 (N_12755,N_11895,N_11603);
nor U12756 (N_12756,N_11939,N_11674);
and U12757 (N_12757,N_11198,N_11060);
and U12758 (N_12758,N_11836,N_11644);
or U12759 (N_12759,N_11120,N_11476);
nand U12760 (N_12760,N_11184,N_11597);
nor U12761 (N_12761,N_11948,N_11779);
and U12762 (N_12762,N_11061,N_11604);
and U12763 (N_12763,N_11649,N_11810);
xor U12764 (N_12764,N_11547,N_11229);
or U12765 (N_12765,N_11551,N_11001);
xnor U12766 (N_12766,N_11061,N_11292);
nor U12767 (N_12767,N_11259,N_11949);
or U12768 (N_12768,N_11810,N_11732);
nor U12769 (N_12769,N_11439,N_11309);
xnor U12770 (N_12770,N_11945,N_11258);
and U12771 (N_12771,N_11758,N_11092);
and U12772 (N_12772,N_11962,N_11476);
nor U12773 (N_12773,N_11577,N_11023);
or U12774 (N_12774,N_11960,N_11203);
or U12775 (N_12775,N_11955,N_11610);
nor U12776 (N_12776,N_11496,N_11198);
and U12777 (N_12777,N_11959,N_11147);
and U12778 (N_12778,N_11860,N_11586);
nor U12779 (N_12779,N_11514,N_11241);
and U12780 (N_12780,N_11852,N_11902);
xor U12781 (N_12781,N_11798,N_11979);
and U12782 (N_12782,N_11260,N_11118);
and U12783 (N_12783,N_11374,N_11329);
nor U12784 (N_12784,N_11107,N_11688);
nand U12785 (N_12785,N_11274,N_11421);
nor U12786 (N_12786,N_11642,N_11536);
xnor U12787 (N_12787,N_11751,N_11449);
nand U12788 (N_12788,N_11502,N_11468);
nand U12789 (N_12789,N_11263,N_11452);
nor U12790 (N_12790,N_11803,N_11039);
or U12791 (N_12791,N_11971,N_11488);
nor U12792 (N_12792,N_11552,N_11301);
nand U12793 (N_12793,N_11482,N_11319);
nand U12794 (N_12794,N_11082,N_11632);
nor U12795 (N_12795,N_11391,N_11785);
nand U12796 (N_12796,N_11536,N_11537);
or U12797 (N_12797,N_11767,N_11084);
nor U12798 (N_12798,N_11232,N_11689);
nor U12799 (N_12799,N_11742,N_11352);
nor U12800 (N_12800,N_11101,N_11748);
xor U12801 (N_12801,N_11090,N_11781);
nand U12802 (N_12802,N_11283,N_11956);
nor U12803 (N_12803,N_11836,N_11624);
nand U12804 (N_12804,N_11319,N_11272);
xnor U12805 (N_12805,N_11920,N_11288);
nor U12806 (N_12806,N_11616,N_11864);
nor U12807 (N_12807,N_11114,N_11137);
nand U12808 (N_12808,N_11026,N_11290);
or U12809 (N_12809,N_11850,N_11351);
and U12810 (N_12810,N_11108,N_11055);
xor U12811 (N_12811,N_11865,N_11943);
nor U12812 (N_12812,N_11044,N_11496);
and U12813 (N_12813,N_11142,N_11120);
xnor U12814 (N_12814,N_11232,N_11498);
and U12815 (N_12815,N_11722,N_11247);
nor U12816 (N_12816,N_11678,N_11267);
and U12817 (N_12817,N_11891,N_11093);
xor U12818 (N_12818,N_11552,N_11539);
xnor U12819 (N_12819,N_11329,N_11852);
or U12820 (N_12820,N_11008,N_11092);
or U12821 (N_12821,N_11299,N_11179);
and U12822 (N_12822,N_11516,N_11150);
nand U12823 (N_12823,N_11254,N_11180);
xnor U12824 (N_12824,N_11883,N_11192);
and U12825 (N_12825,N_11979,N_11609);
nor U12826 (N_12826,N_11124,N_11061);
xnor U12827 (N_12827,N_11400,N_11132);
and U12828 (N_12828,N_11506,N_11216);
or U12829 (N_12829,N_11339,N_11322);
and U12830 (N_12830,N_11127,N_11173);
nor U12831 (N_12831,N_11132,N_11296);
and U12832 (N_12832,N_11073,N_11219);
nand U12833 (N_12833,N_11336,N_11856);
or U12834 (N_12834,N_11133,N_11215);
xnor U12835 (N_12835,N_11546,N_11875);
xor U12836 (N_12836,N_11495,N_11016);
and U12837 (N_12837,N_11446,N_11267);
nand U12838 (N_12838,N_11271,N_11618);
xor U12839 (N_12839,N_11070,N_11324);
nand U12840 (N_12840,N_11091,N_11688);
nand U12841 (N_12841,N_11793,N_11945);
nor U12842 (N_12842,N_11925,N_11882);
or U12843 (N_12843,N_11467,N_11221);
and U12844 (N_12844,N_11068,N_11569);
or U12845 (N_12845,N_11741,N_11307);
or U12846 (N_12846,N_11630,N_11799);
and U12847 (N_12847,N_11330,N_11160);
xor U12848 (N_12848,N_11057,N_11249);
xnor U12849 (N_12849,N_11949,N_11013);
xnor U12850 (N_12850,N_11345,N_11720);
xor U12851 (N_12851,N_11584,N_11907);
and U12852 (N_12852,N_11308,N_11877);
nand U12853 (N_12853,N_11187,N_11002);
or U12854 (N_12854,N_11075,N_11752);
or U12855 (N_12855,N_11981,N_11653);
nor U12856 (N_12856,N_11625,N_11996);
or U12857 (N_12857,N_11918,N_11364);
nor U12858 (N_12858,N_11303,N_11448);
or U12859 (N_12859,N_11038,N_11390);
or U12860 (N_12860,N_11917,N_11601);
and U12861 (N_12861,N_11067,N_11699);
xor U12862 (N_12862,N_11755,N_11863);
xor U12863 (N_12863,N_11764,N_11825);
nor U12864 (N_12864,N_11904,N_11052);
xor U12865 (N_12865,N_11913,N_11904);
nand U12866 (N_12866,N_11589,N_11350);
xor U12867 (N_12867,N_11173,N_11193);
or U12868 (N_12868,N_11700,N_11200);
and U12869 (N_12869,N_11044,N_11269);
nor U12870 (N_12870,N_11655,N_11635);
xor U12871 (N_12871,N_11358,N_11766);
or U12872 (N_12872,N_11128,N_11873);
nand U12873 (N_12873,N_11093,N_11977);
nand U12874 (N_12874,N_11123,N_11730);
xnor U12875 (N_12875,N_11170,N_11812);
nand U12876 (N_12876,N_11704,N_11683);
and U12877 (N_12877,N_11869,N_11846);
or U12878 (N_12878,N_11655,N_11432);
xor U12879 (N_12879,N_11435,N_11427);
nor U12880 (N_12880,N_11713,N_11309);
and U12881 (N_12881,N_11968,N_11434);
xor U12882 (N_12882,N_11781,N_11130);
xor U12883 (N_12883,N_11767,N_11436);
nor U12884 (N_12884,N_11849,N_11276);
or U12885 (N_12885,N_11278,N_11389);
xor U12886 (N_12886,N_11601,N_11887);
or U12887 (N_12887,N_11234,N_11591);
nand U12888 (N_12888,N_11976,N_11214);
or U12889 (N_12889,N_11161,N_11437);
or U12890 (N_12890,N_11367,N_11737);
or U12891 (N_12891,N_11622,N_11552);
nor U12892 (N_12892,N_11113,N_11914);
or U12893 (N_12893,N_11767,N_11530);
nand U12894 (N_12894,N_11902,N_11307);
nor U12895 (N_12895,N_11450,N_11687);
nand U12896 (N_12896,N_11094,N_11592);
xor U12897 (N_12897,N_11020,N_11519);
and U12898 (N_12898,N_11728,N_11841);
nand U12899 (N_12899,N_11112,N_11308);
or U12900 (N_12900,N_11884,N_11056);
nor U12901 (N_12901,N_11757,N_11909);
or U12902 (N_12902,N_11146,N_11159);
xnor U12903 (N_12903,N_11799,N_11943);
and U12904 (N_12904,N_11392,N_11004);
xor U12905 (N_12905,N_11282,N_11656);
and U12906 (N_12906,N_11371,N_11739);
nand U12907 (N_12907,N_11196,N_11139);
and U12908 (N_12908,N_11980,N_11754);
and U12909 (N_12909,N_11228,N_11737);
nor U12910 (N_12910,N_11239,N_11156);
nor U12911 (N_12911,N_11447,N_11875);
or U12912 (N_12912,N_11452,N_11365);
and U12913 (N_12913,N_11561,N_11439);
or U12914 (N_12914,N_11619,N_11956);
and U12915 (N_12915,N_11425,N_11872);
and U12916 (N_12916,N_11411,N_11020);
or U12917 (N_12917,N_11967,N_11378);
xor U12918 (N_12918,N_11996,N_11664);
or U12919 (N_12919,N_11907,N_11345);
nor U12920 (N_12920,N_11538,N_11149);
xor U12921 (N_12921,N_11333,N_11162);
xor U12922 (N_12922,N_11903,N_11016);
or U12923 (N_12923,N_11615,N_11249);
xnor U12924 (N_12924,N_11638,N_11111);
and U12925 (N_12925,N_11541,N_11615);
xor U12926 (N_12926,N_11625,N_11560);
or U12927 (N_12927,N_11966,N_11746);
nor U12928 (N_12928,N_11761,N_11651);
nor U12929 (N_12929,N_11734,N_11613);
nand U12930 (N_12930,N_11715,N_11053);
nand U12931 (N_12931,N_11601,N_11069);
or U12932 (N_12932,N_11568,N_11758);
or U12933 (N_12933,N_11857,N_11429);
and U12934 (N_12934,N_11364,N_11474);
or U12935 (N_12935,N_11674,N_11348);
and U12936 (N_12936,N_11912,N_11609);
nand U12937 (N_12937,N_11724,N_11026);
xnor U12938 (N_12938,N_11386,N_11299);
nor U12939 (N_12939,N_11048,N_11375);
nor U12940 (N_12940,N_11013,N_11615);
nor U12941 (N_12941,N_11439,N_11633);
nand U12942 (N_12942,N_11332,N_11061);
or U12943 (N_12943,N_11526,N_11697);
nor U12944 (N_12944,N_11272,N_11557);
nor U12945 (N_12945,N_11694,N_11034);
and U12946 (N_12946,N_11689,N_11167);
or U12947 (N_12947,N_11081,N_11718);
and U12948 (N_12948,N_11276,N_11744);
nor U12949 (N_12949,N_11045,N_11291);
nand U12950 (N_12950,N_11222,N_11550);
nor U12951 (N_12951,N_11411,N_11518);
and U12952 (N_12952,N_11450,N_11956);
nor U12953 (N_12953,N_11168,N_11428);
nor U12954 (N_12954,N_11529,N_11340);
nor U12955 (N_12955,N_11729,N_11118);
nand U12956 (N_12956,N_11032,N_11603);
nor U12957 (N_12957,N_11685,N_11425);
nor U12958 (N_12958,N_11308,N_11380);
xor U12959 (N_12959,N_11519,N_11385);
xor U12960 (N_12960,N_11989,N_11942);
nand U12961 (N_12961,N_11549,N_11304);
xnor U12962 (N_12962,N_11505,N_11239);
or U12963 (N_12963,N_11053,N_11402);
or U12964 (N_12964,N_11330,N_11738);
nand U12965 (N_12965,N_11542,N_11216);
xor U12966 (N_12966,N_11864,N_11156);
or U12967 (N_12967,N_11947,N_11401);
and U12968 (N_12968,N_11444,N_11543);
xor U12969 (N_12969,N_11431,N_11897);
or U12970 (N_12970,N_11866,N_11410);
nor U12971 (N_12971,N_11613,N_11769);
or U12972 (N_12972,N_11846,N_11749);
and U12973 (N_12973,N_11180,N_11012);
nor U12974 (N_12974,N_11994,N_11212);
or U12975 (N_12975,N_11852,N_11285);
and U12976 (N_12976,N_11419,N_11649);
or U12977 (N_12977,N_11839,N_11572);
nor U12978 (N_12978,N_11217,N_11791);
xor U12979 (N_12979,N_11760,N_11790);
xor U12980 (N_12980,N_11009,N_11825);
nand U12981 (N_12981,N_11921,N_11912);
or U12982 (N_12982,N_11340,N_11648);
nand U12983 (N_12983,N_11402,N_11521);
or U12984 (N_12984,N_11665,N_11979);
nor U12985 (N_12985,N_11753,N_11484);
or U12986 (N_12986,N_11210,N_11636);
nor U12987 (N_12987,N_11613,N_11214);
xor U12988 (N_12988,N_11296,N_11598);
nand U12989 (N_12989,N_11455,N_11680);
nor U12990 (N_12990,N_11742,N_11091);
nor U12991 (N_12991,N_11979,N_11421);
and U12992 (N_12992,N_11981,N_11587);
and U12993 (N_12993,N_11323,N_11225);
xor U12994 (N_12994,N_11328,N_11100);
xor U12995 (N_12995,N_11554,N_11224);
or U12996 (N_12996,N_11214,N_11912);
xor U12997 (N_12997,N_11258,N_11229);
or U12998 (N_12998,N_11191,N_11363);
or U12999 (N_12999,N_11557,N_11115);
and U13000 (N_13000,N_12485,N_12594);
nand U13001 (N_13001,N_12365,N_12360);
xor U13002 (N_13002,N_12284,N_12916);
and U13003 (N_13003,N_12888,N_12155);
nand U13004 (N_13004,N_12641,N_12024);
nor U13005 (N_13005,N_12402,N_12100);
or U13006 (N_13006,N_12309,N_12023);
and U13007 (N_13007,N_12630,N_12156);
nand U13008 (N_13008,N_12821,N_12112);
and U13009 (N_13009,N_12478,N_12054);
or U13010 (N_13010,N_12083,N_12537);
nand U13011 (N_13011,N_12885,N_12801);
nor U13012 (N_13012,N_12538,N_12279);
xor U13013 (N_13013,N_12524,N_12527);
and U13014 (N_13014,N_12443,N_12231);
nor U13015 (N_13015,N_12976,N_12462);
and U13016 (N_13016,N_12132,N_12130);
nand U13017 (N_13017,N_12922,N_12242);
nand U13018 (N_13018,N_12094,N_12610);
and U13019 (N_13019,N_12590,N_12535);
nor U13020 (N_13020,N_12341,N_12247);
nor U13021 (N_13021,N_12985,N_12109);
nand U13022 (N_13022,N_12545,N_12404);
xor U13023 (N_13023,N_12992,N_12064);
nor U13024 (N_13024,N_12855,N_12308);
xor U13025 (N_13025,N_12771,N_12474);
xor U13026 (N_13026,N_12297,N_12603);
nor U13027 (N_13027,N_12748,N_12999);
nor U13028 (N_13028,N_12160,N_12219);
xnor U13029 (N_13029,N_12166,N_12546);
nand U13030 (N_13030,N_12446,N_12549);
nor U13031 (N_13031,N_12361,N_12298);
and U13032 (N_13032,N_12306,N_12802);
xnor U13033 (N_13033,N_12528,N_12456);
and U13034 (N_13034,N_12548,N_12810);
or U13035 (N_13035,N_12710,N_12269);
nor U13036 (N_13036,N_12792,N_12719);
and U13037 (N_13037,N_12529,N_12206);
or U13038 (N_13038,N_12048,N_12775);
and U13039 (N_13039,N_12099,N_12292);
or U13040 (N_13040,N_12941,N_12628);
nor U13041 (N_13041,N_12723,N_12749);
xor U13042 (N_13042,N_12962,N_12965);
xnor U13043 (N_13043,N_12479,N_12335);
or U13044 (N_13044,N_12761,N_12173);
xnor U13045 (N_13045,N_12424,N_12319);
or U13046 (N_13046,N_12518,N_12271);
nand U13047 (N_13047,N_12035,N_12949);
nand U13048 (N_13048,N_12872,N_12191);
and U13049 (N_13049,N_12832,N_12891);
xor U13050 (N_13050,N_12374,N_12724);
and U13051 (N_13051,N_12451,N_12412);
and U13052 (N_13052,N_12522,N_12889);
xor U13053 (N_13053,N_12551,N_12531);
xnor U13054 (N_13054,N_12447,N_12364);
nand U13055 (N_13055,N_12260,N_12880);
or U13056 (N_13056,N_12349,N_12919);
or U13057 (N_13057,N_12979,N_12849);
or U13058 (N_13058,N_12777,N_12744);
and U13059 (N_13059,N_12815,N_12542);
nand U13060 (N_13060,N_12585,N_12042);
nor U13061 (N_13061,N_12974,N_12987);
xnor U13062 (N_13062,N_12826,N_12726);
xor U13063 (N_13063,N_12986,N_12669);
xor U13064 (N_13064,N_12058,N_12684);
nand U13065 (N_13065,N_12452,N_12805);
and U13066 (N_13066,N_12977,N_12138);
nand U13067 (N_13067,N_12275,N_12214);
nand U13068 (N_13068,N_12003,N_12601);
or U13069 (N_13069,N_12510,N_12147);
and U13070 (N_13070,N_12140,N_12526);
xor U13071 (N_13071,N_12783,N_12468);
nor U13072 (N_13072,N_12914,N_12934);
xor U13073 (N_13073,N_12505,N_12569);
xnor U13074 (N_13074,N_12366,N_12073);
xor U13075 (N_13075,N_12770,N_12253);
and U13076 (N_13076,N_12653,N_12691);
nand U13077 (N_13077,N_12852,N_12091);
or U13078 (N_13078,N_12090,N_12146);
and U13079 (N_13079,N_12069,N_12346);
nand U13080 (N_13080,N_12718,N_12932);
and U13081 (N_13081,N_12781,N_12520);
nor U13082 (N_13082,N_12325,N_12912);
xor U13083 (N_13083,N_12359,N_12400);
nor U13084 (N_13084,N_12337,N_12107);
or U13085 (N_13085,N_12800,N_12789);
and U13086 (N_13086,N_12621,N_12564);
xnor U13087 (N_13087,N_12642,N_12989);
nor U13088 (N_13088,N_12387,N_12172);
nand U13089 (N_13089,N_12116,N_12455);
nand U13090 (N_13090,N_12980,N_12931);
and U13091 (N_13091,N_12790,N_12115);
and U13092 (N_13092,N_12706,N_12611);
nand U13093 (N_13093,N_12288,N_12908);
nand U13094 (N_13094,N_12961,N_12806);
and U13095 (N_13095,N_12694,N_12082);
nor U13096 (N_13096,N_12756,N_12878);
and U13097 (N_13097,N_12933,N_12597);
nand U13098 (N_13098,N_12263,N_12238);
xnor U13099 (N_13099,N_12157,N_12791);
nor U13100 (N_13100,N_12016,N_12123);
nand U13101 (N_13101,N_12311,N_12390);
or U13102 (N_13102,N_12993,N_12001);
or U13103 (N_13103,N_12521,N_12689);
xnor U13104 (N_13104,N_12576,N_12406);
and U13105 (N_13105,N_12525,N_12385);
xnor U13106 (N_13106,N_12063,N_12409);
nor U13107 (N_13107,N_12228,N_12798);
or U13108 (N_13108,N_12093,N_12799);
and U13109 (N_13109,N_12418,N_12469);
or U13110 (N_13110,N_12760,N_12489);
xnor U13111 (N_13111,N_12465,N_12725);
nor U13112 (N_13112,N_12286,N_12301);
nor U13113 (N_13113,N_12786,N_12274);
or U13114 (N_13114,N_12907,N_12321);
nor U13115 (N_13115,N_12210,N_12644);
xnor U13116 (N_13116,N_12680,N_12667);
nand U13117 (N_13117,N_12072,N_12473);
nand U13118 (N_13118,N_12794,N_12948);
nand U13119 (N_13119,N_12512,N_12595);
and U13120 (N_13120,N_12212,N_12126);
and U13121 (N_13121,N_12764,N_12327);
nor U13122 (N_13122,N_12445,N_12394);
nand U13123 (N_13123,N_12250,N_12399);
xnor U13124 (N_13124,N_12646,N_12753);
or U13125 (N_13125,N_12436,N_12398);
xnor U13126 (N_13126,N_12196,N_12830);
or U13127 (N_13127,N_12532,N_12060);
and U13128 (N_13128,N_12937,N_12076);
and U13129 (N_13129,N_12788,N_12056);
xnor U13130 (N_13130,N_12197,N_12005);
or U13131 (N_13131,N_12833,N_12230);
and U13132 (N_13132,N_12763,N_12491);
xnor U13133 (N_13133,N_12281,N_12362);
nor U13134 (N_13134,N_12876,N_12998);
nor U13135 (N_13135,N_12894,N_12618);
or U13136 (N_13136,N_12735,N_12939);
xnor U13137 (N_13137,N_12515,N_12258);
xor U13138 (N_13138,N_12517,N_12293);
xor U13139 (N_13139,N_12136,N_12671);
xor U13140 (N_13140,N_12434,N_12395);
xor U13141 (N_13141,N_12114,N_12245);
or U13142 (N_13142,N_12108,N_12079);
xnor U13143 (N_13143,N_12829,N_12075);
nor U13144 (N_13144,N_12938,N_12541);
or U13145 (N_13145,N_12127,N_12354);
nand U13146 (N_13146,N_12303,N_12012);
or U13147 (N_13147,N_12313,N_12622);
nand U13148 (N_13148,N_12088,N_12851);
or U13149 (N_13149,N_12645,N_12233);
or U13150 (N_13150,N_12928,N_12574);
xor U13151 (N_13151,N_12222,N_12033);
nor U13152 (N_13152,N_12808,N_12831);
or U13153 (N_13153,N_12209,N_12811);
xor U13154 (N_13154,N_12995,N_12699);
and U13155 (N_13155,N_12251,N_12007);
nor U13156 (N_13156,N_12070,N_12417);
xnor U13157 (N_13157,N_12199,N_12432);
or U13158 (N_13158,N_12128,N_12778);
nand U13159 (N_13159,N_12170,N_12825);
nor U13160 (N_13160,N_12623,N_12580);
xor U13161 (N_13161,N_12501,N_12591);
or U13162 (N_13162,N_12759,N_12617);
and U13163 (N_13163,N_12187,N_12375);
nor U13164 (N_13164,N_12442,N_12865);
nand U13165 (N_13165,N_12037,N_12913);
or U13166 (N_13166,N_12860,N_12910);
xor U13167 (N_13167,N_12869,N_12282);
xor U13168 (N_13168,N_12670,N_12936);
nor U13169 (N_13169,N_12660,N_12807);
nand U13170 (N_13170,N_12066,N_12661);
and U13171 (N_13171,N_12722,N_12785);
and U13172 (N_13172,N_12539,N_12158);
nor U13173 (N_13173,N_12514,N_12113);
and U13174 (N_13174,N_12729,N_12483);
or U13175 (N_13175,N_12071,N_12034);
nand U13176 (N_13176,N_12502,N_12596);
or U13177 (N_13177,N_12384,N_12973);
xnor U13178 (N_13178,N_12150,N_12148);
xor U13179 (N_13179,N_12612,N_12078);
xor U13180 (N_13180,N_12896,N_12427);
xnor U13181 (N_13181,N_12015,N_12420);
or U13182 (N_13182,N_12813,N_12847);
nand U13183 (N_13183,N_12262,N_12178);
xor U13184 (N_13184,N_12708,N_12019);
xnor U13185 (N_13185,N_12240,N_12946);
and U13186 (N_13186,N_12296,N_12453);
xor U13187 (N_13187,N_12353,N_12081);
nand U13188 (N_13188,N_12804,N_12217);
or U13189 (N_13189,N_12853,N_12487);
nand U13190 (N_13190,N_12448,N_12200);
nand U13191 (N_13191,N_12905,N_12457);
xnor U13192 (N_13192,N_12709,N_12086);
or U13193 (N_13193,N_12589,N_12803);
or U13194 (N_13194,N_12039,N_12310);
xor U13195 (N_13195,N_12599,N_12105);
nand U13196 (N_13196,N_12678,N_12643);
nor U13197 (N_13197,N_12864,N_12440);
nor U13198 (N_13198,N_12267,N_12782);
or U13199 (N_13199,N_12774,N_12673);
and U13200 (N_13200,N_12499,N_12571);
nor U13201 (N_13201,N_12085,N_12425);
and U13202 (N_13202,N_12903,N_12547);
nand U13203 (N_13203,N_12882,N_12111);
xor U13204 (N_13204,N_12714,N_12958);
nand U13205 (N_13205,N_12002,N_12413);
or U13206 (N_13206,N_12924,N_12117);
and U13207 (N_13207,N_12615,N_12221);
nor U13208 (N_13208,N_12106,N_12318);
nor U13209 (N_13209,N_12236,N_12963);
and U13210 (N_13210,N_12376,N_12859);
and U13211 (N_13211,N_12686,N_12655);
or U13212 (N_13212,N_12017,N_12020);
nor U13213 (N_13213,N_12061,N_12488);
nand U13214 (N_13214,N_12225,N_12969);
nor U13215 (N_13215,N_12193,N_12736);
nor U13216 (N_13216,N_12386,N_12049);
and U13217 (N_13217,N_12142,N_12681);
and U13218 (N_13218,N_12895,N_12254);
and U13219 (N_13219,N_12947,N_12863);
or U13220 (N_13220,N_12837,N_12243);
nor U13221 (N_13221,N_12649,N_12836);
xnor U13222 (N_13222,N_12294,N_12171);
or U13223 (N_13223,N_12339,N_12110);
nor U13224 (N_13224,N_12183,N_12163);
or U13225 (N_13225,N_12819,N_12139);
and U13226 (N_13226,N_12059,N_12356);
nor U13227 (N_13227,N_12982,N_12264);
and U13228 (N_13228,N_12496,N_12768);
nand U13229 (N_13229,N_12135,N_12368);
or U13230 (N_13230,N_12161,N_12227);
and U13231 (N_13231,N_12181,N_12165);
or U13232 (N_13232,N_12118,N_12342);
or U13233 (N_13233,N_12614,N_12504);
nand U13234 (N_13234,N_12031,N_12248);
xnor U13235 (N_13235,N_12272,N_12122);
and U13236 (N_13236,N_12021,N_12654);
and U13237 (N_13237,N_12244,N_12917);
or U13238 (N_13238,N_12096,N_12182);
xor U13239 (N_13239,N_12040,N_12822);
or U13240 (N_13240,N_12103,N_12897);
and U13241 (N_13241,N_12834,N_12340);
nand U13242 (N_13242,N_12416,N_12755);
xor U13243 (N_13243,N_12757,N_12769);
xnor U13244 (N_13244,N_12553,N_12698);
xnor U13245 (N_13245,N_12246,N_12902);
xnor U13246 (N_13246,N_12584,N_12273);
or U13247 (N_13247,N_12509,N_12014);
nor U13248 (N_13248,N_12960,N_12942);
xor U13249 (N_13249,N_12751,N_12666);
and U13250 (N_13250,N_12018,N_12046);
and U13251 (N_13251,N_12787,N_12711);
or U13252 (N_13252,N_12923,N_12036);
nor U13253 (N_13253,N_12044,N_12577);
or U13254 (N_13254,N_12195,N_12415);
and U13255 (N_13255,N_12350,N_12629);
nand U13256 (N_13256,N_12846,N_12475);
xor U13257 (N_13257,N_12506,N_12077);
xnor U13258 (N_13258,N_12372,N_12433);
or U13259 (N_13259,N_12378,N_12430);
and U13260 (N_13260,N_12188,N_12557);
nand U13261 (N_13261,N_12270,N_12743);
or U13262 (N_13262,N_12682,N_12991);
or U13263 (N_13263,N_12935,N_12609);
or U13264 (N_13264,N_12676,N_12164);
and U13265 (N_13265,N_12028,N_12940);
or U13266 (N_13266,N_12280,N_12561);
or U13267 (N_13267,N_12032,N_12022);
xor U13268 (N_13268,N_12693,N_12008);
and U13269 (N_13269,N_12728,N_12844);
and U13270 (N_13270,N_12556,N_12582);
nor U13271 (N_13271,N_12784,N_12981);
xor U13272 (N_13272,N_12702,N_12766);
xnor U13273 (N_13273,N_12652,N_12009);
nand U13274 (N_13274,N_12396,N_12747);
and U13275 (N_13275,N_12431,N_12593);
xnor U13276 (N_13276,N_12915,N_12382);
or U13277 (N_13277,N_12131,N_12441);
and U13278 (N_13278,N_12369,N_12712);
nand U13279 (N_13279,N_12348,N_12381);
and U13280 (N_13280,N_12237,N_12920);
nand U13281 (N_13281,N_12814,N_12823);
nand U13282 (N_13282,N_12167,N_12675);
or U13283 (N_13283,N_12256,N_12632);
nor U13284 (N_13284,N_12773,N_12926);
nor U13285 (N_13285,N_12363,N_12624);
and U13286 (N_13286,N_12705,N_12930);
or U13287 (N_13287,N_12845,N_12011);
nor U13288 (N_13288,N_12423,N_12168);
or U13289 (N_13289,N_12216,N_12704);
xor U13290 (N_13290,N_12765,N_12638);
nand U13291 (N_13291,N_12635,N_12334);
xnor U13292 (N_13292,N_12276,N_12658);
xor U13293 (N_13293,N_12358,N_12426);
nor U13294 (N_13294,N_12038,N_12964);
or U13295 (N_13295,N_12707,N_12184);
and U13296 (N_13296,N_12174,N_12687);
nand U13297 (N_13297,N_12041,N_12450);
and U13298 (N_13298,N_12600,N_12731);
and U13299 (N_13299,N_12534,N_12218);
nand U13300 (N_13300,N_12563,N_12169);
xnor U13301 (N_13301,N_12486,N_12383);
and U13302 (N_13302,N_12133,N_12640);
or U13303 (N_13303,N_12898,N_12498);
nand U13304 (N_13304,N_12300,N_12631);
and U13305 (N_13305,N_12223,N_12467);
or U13306 (N_13306,N_12662,N_12740);
xor U13307 (N_13307,N_12820,N_12320);
or U13308 (N_13308,N_12151,N_12047);
xnor U13309 (N_13309,N_12175,N_12824);
and U13310 (N_13310,N_12067,N_12929);
nor U13311 (N_13311,N_12862,N_12754);
nand U13312 (N_13312,N_12809,N_12454);
or U13313 (N_13313,N_12881,N_12438);
nand U13314 (N_13314,N_12145,N_12429);
xnor U13315 (N_13315,N_12351,N_12516);
nor U13316 (N_13316,N_12154,N_12659);
xor U13317 (N_13317,N_12816,N_12153);
nand U13318 (N_13318,N_12536,N_12886);
and U13319 (N_13319,N_12951,N_12758);
nand U13320 (N_13320,N_12180,N_12010);
nand U13321 (N_13321,N_12051,N_12968);
xor U13322 (N_13322,N_12605,N_12877);
and U13323 (N_13323,N_12975,N_12795);
and U13324 (N_13324,N_12205,N_12772);
xor U13325 (N_13325,N_12344,N_12411);
or U13326 (N_13326,N_12634,N_12767);
and U13327 (N_13327,N_12879,N_12393);
nand U13328 (N_13328,N_12857,N_12084);
nor U13329 (N_13329,N_12890,N_12224);
nor U13330 (N_13330,N_12204,N_12668);
nor U13331 (N_13331,N_12651,N_12636);
xor U13332 (N_13332,N_12746,N_12573);
nand U13333 (N_13333,N_12970,N_12866);
nand U13334 (N_13334,N_12586,N_12388);
or U13335 (N_13335,N_12291,N_12098);
and U13336 (N_13336,N_12149,N_12484);
and U13337 (N_13337,N_12997,N_12435);
and U13338 (N_13338,N_12285,N_12322);
nor U13339 (N_13339,N_12555,N_12259);
and U13340 (N_13340,N_12332,N_12732);
and U13341 (N_13341,N_12373,N_12377);
or U13342 (N_13342,N_12690,N_12883);
nand U13343 (N_13343,N_12215,N_12730);
xnor U13344 (N_13344,N_12656,N_12232);
and U13345 (N_13345,N_12087,N_12608);
and U13346 (N_13346,N_12871,N_12190);
nor U13347 (N_13347,N_12013,N_12550);
or U13348 (N_13348,N_12302,N_12950);
xnor U13349 (N_13349,N_12352,N_12533);
nand U13350 (N_13350,N_12620,N_12065);
nor U13351 (N_13351,N_12925,N_12328);
and U13352 (N_13352,N_12570,N_12868);
nor U13353 (N_13353,N_12848,N_12026);
nand U13354 (N_13354,N_12884,N_12208);
or U13355 (N_13355,N_12124,N_12952);
nand U13356 (N_13356,N_12125,N_12818);
and U13357 (N_13357,N_12639,N_12305);
or U13358 (N_13358,N_12422,N_12598);
or U13359 (N_13359,N_12141,N_12207);
xor U13360 (N_13360,N_12477,N_12439);
or U13361 (N_13361,N_12480,N_12226);
or U13362 (N_13362,N_12906,N_12476);
or U13363 (N_13363,N_12336,N_12578);
or U13364 (N_13364,N_12494,N_12089);
nand U13365 (N_13365,N_12458,N_12472);
or U13366 (N_13366,N_12616,N_12873);
nand U13367 (N_13367,N_12921,N_12397);
nor U13368 (N_13368,N_12568,N_12481);
nand U13369 (N_13369,N_12410,N_12945);
nand U13370 (N_13370,N_12095,N_12025);
xnor U13371 (N_13371,N_12552,N_12892);
nand U13372 (N_13372,N_12482,N_12750);
or U13373 (N_13373,N_12911,N_12606);
xor U13374 (N_13374,N_12211,N_12490);
nor U13375 (N_13375,N_12198,N_12459);
or U13376 (N_13376,N_12203,N_12062);
or U13377 (N_13377,N_12742,N_12967);
nand U13378 (N_13378,N_12403,N_12843);
nor U13379 (N_13379,N_12613,N_12672);
or U13380 (N_13380,N_12572,N_12000);
nand U13381 (N_13381,N_12371,N_12194);
nand U13382 (N_13382,N_12978,N_12045);
nor U13383 (N_13383,N_12213,N_12647);
and U13384 (N_13384,N_12796,N_12343);
xnor U13385 (N_13385,N_12324,N_12329);
and U13386 (N_13386,N_12717,N_12817);
and U13387 (N_13387,N_12893,N_12887);
and U13388 (N_13388,N_12650,N_12289);
and U13389 (N_13389,N_12752,N_12055);
xor U13390 (N_13390,N_12626,N_12850);
and U13391 (N_13391,N_12900,N_12414);
nand U13392 (N_13392,N_12657,N_12720);
or U13393 (N_13393,N_12307,N_12239);
nand U13394 (N_13394,N_12953,N_12513);
xor U13395 (N_13395,N_12575,N_12841);
xor U13396 (N_13396,N_12421,N_12287);
nand U13397 (N_13397,N_12201,N_12129);
nor U13398 (N_13398,N_12856,N_12314);
or U13399 (N_13399,N_12665,N_12053);
xnor U13400 (N_13400,N_12102,N_12990);
or U13401 (N_13401,N_12004,N_12176);
nor U13402 (N_13402,N_12252,N_12779);
nor U13403 (N_13403,N_12104,N_12700);
xnor U13404 (N_13404,N_12966,N_12317);
nor U13405 (N_13405,N_12470,N_12762);
or U13406 (N_13406,N_12554,N_12234);
nand U13407 (N_13407,N_12345,N_12428);
xor U13408 (N_13408,N_12583,N_12793);
nor U13409 (N_13409,N_12648,N_12544);
and U13410 (N_13410,N_12523,N_12492);
or U13411 (N_13411,N_12664,N_12179);
xor U13412 (N_13412,N_12738,N_12679);
nand U13413 (N_13413,N_12683,N_12592);
and U13414 (N_13414,N_12315,N_12955);
nor U13415 (N_13415,N_12074,N_12331);
xnor U13416 (N_13416,N_12299,N_12715);
xor U13417 (N_13417,N_12565,N_12838);
or U13418 (N_13418,N_12134,N_12677);
and U13419 (N_13419,N_12347,N_12092);
xnor U13420 (N_13420,N_12627,N_12685);
or U13421 (N_13421,N_12407,N_12701);
or U13422 (N_13422,N_12994,N_12290);
nor U13423 (N_13423,N_12943,N_12192);
or U13424 (N_13424,N_12737,N_12029);
or U13425 (N_13425,N_12828,N_12721);
or U13426 (N_13426,N_12278,N_12562);
or U13427 (N_13427,N_12466,N_12121);
xnor U13428 (N_13428,N_12152,N_12137);
nor U13429 (N_13429,N_12101,N_12493);
nor U13430 (N_13430,N_12006,N_12739);
nand U13431 (N_13431,N_12380,N_12229);
nor U13432 (N_13432,N_12904,N_12674);
nand U13433 (N_13433,N_12326,N_12027);
nor U13434 (N_13434,N_12954,N_12776);
nor U13435 (N_13435,N_12835,N_12697);
nor U13436 (N_13436,N_12268,N_12560);
and U13437 (N_13437,N_12875,N_12080);
nand U13438 (N_13438,N_12870,N_12604);
nand U13439 (N_13439,N_12909,N_12255);
nand U13440 (N_13440,N_12405,N_12588);
nand U13441 (N_13441,N_12177,N_12696);
nand U13442 (N_13442,N_12367,N_12607);
xnor U13443 (N_13443,N_12097,N_12745);
xor U13444 (N_13444,N_12330,N_12444);
xnor U13445 (N_13445,N_12530,N_12392);
and U13446 (N_13446,N_12780,N_12688);
nor U13447 (N_13447,N_12304,N_12261);
xor U13448 (N_13448,N_12323,N_12988);
or U13449 (N_13449,N_12495,N_12497);
nand U13450 (N_13450,N_12463,N_12068);
and U13451 (N_13451,N_12333,N_12241);
nor U13452 (N_13452,N_12389,N_12692);
xor U13453 (N_13453,N_12663,N_12316);
nand U13454 (N_13454,N_12713,N_12867);
nand U13455 (N_13455,N_12186,N_12419);
nand U13456 (N_13456,N_12312,N_12842);
and U13457 (N_13457,N_12401,N_12119);
and U13458 (N_13458,N_12500,N_12727);
or U13459 (N_13459,N_12567,N_12460);
and U13460 (N_13460,N_12357,N_12901);
nor U13461 (N_13461,N_12143,N_12741);
xnor U13462 (N_13462,N_12840,N_12858);
nand U13463 (N_13463,N_12959,N_12052);
xor U13464 (N_13464,N_12983,N_12559);
and U13465 (N_13465,N_12503,N_12159);
nor U13466 (N_13466,N_12519,N_12277);
or U13467 (N_13467,N_12266,N_12695);
xnor U13468 (N_13468,N_12972,N_12566);
nor U13469 (N_13469,N_12543,N_12633);
nand U13470 (N_13470,N_12120,N_12637);
and U13471 (N_13471,N_12581,N_12057);
xor U13472 (N_13472,N_12619,N_12189);
and U13473 (N_13473,N_12144,N_12956);
or U13474 (N_13474,N_12162,N_12507);
xor U13475 (N_13475,N_12235,N_12957);
nand U13476 (N_13476,N_12471,N_12971);
nand U13477 (N_13477,N_12703,N_12257);
xnor U13478 (N_13478,N_12602,N_12812);
or U13479 (N_13479,N_12391,N_12511);
nand U13480 (N_13480,N_12734,N_12827);
xor U13481 (N_13481,N_12355,N_12370);
nor U13482 (N_13482,N_12338,N_12220);
and U13483 (N_13483,N_12944,N_12899);
nand U13484 (N_13484,N_12797,N_12050);
or U13485 (N_13485,N_12625,N_12249);
nand U13486 (N_13486,N_12854,N_12861);
nor U13487 (N_13487,N_12379,N_12508);
and U13488 (N_13488,N_12874,N_12927);
xor U13489 (N_13489,N_12283,N_12839);
and U13490 (N_13490,N_12464,N_12408);
xnor U13491 (N_13491,N_12265,N_12461);
nand U13492 (N_13492,N_12540,N_12185);
nor U13493 (N_13493,N_12558,N_12295);
and U13494 (N_13494,N_12202,N_12449);
nor U13495 (N_13495,N_12579,N_12043);
xor U13496 (N_13496,N_12733,N_12587);
xnor U13497 (N_13497,N_12716,N_12030);
and U13498 (N_13498,N_12984,N_12996);
and U13499 (N_13499,N_12918,N_12437);
and U13500 (N_13500,N_12512,N_12857);
nor U13501 (N_13501,N_12245,N_12465);
nand U13502 (N_13502,N_12559,N_12187);
xor U13503 (N_13503,N_12488,N_12080);
and U13504 (N_13504,N_12104,N_12631);
nor U13505 (N_13505,N_12611,N_12467);
and U13506 (N_13506,N_12839,N_12355);
xnor U13507 (N_13507,N_12759,N_12028);
nor U13508 (N_13508,N_12901,N_12174);
and U13509 (N_13509,N_12664,N_12098);
nand U13510 (N_13510,N_12448,N_12996);
and U13511 (N_13511,N_12628,N_12720);
nand U13512 (N_13512,N_12986,N_12899);
nor U13513 (N_13513,N_12301,N_12995);
nor U13514 (N_13514,N_12865,N_12949);
xnor U13515 (N_13515,N_12679,N_12695);
nor U13516 (N_13516,N_12868,N_12656);
xor U13517 (N_13517,N_12452,N_12530);
xnor U13518 (N_13518,N_12480,N_12547);
xnor U13519 (N_13519,N_12474,N_12340);
nor U13520 (N_13520,N_12541,N_12957);
xor U13521 (N_13521,N_12530,N_12154);
or U13522 (N_13522,N_12530,N_12433);
xnor U13523 (N_13523,N_12123,N_12277);
and U13524 (N_13524,N_12792,N_12661);
and U13525 (N_13525,N_12869,N_12359);
nor U13526 (N_13526,N_12534,N_12372);
and U13527 (N_13527,N_12997,N_12053);
or U13528 (N_13528,N_12708,N_12006);
nor U13529 (N_13529,N_12569,N_12688);
or U13530 (N_13530,N_12428,N_12622);
or U13531 (N_13531,N_12767,N_12814);
and U13532 (N_13532,N_12405,N_12894);
and U13533 (N_13533,N_12542,N_12579);
xnor U13534 (N_13534,N_12714,N_12117);
nor U13535 (N_13535,N_12340,N_12448);
and U13536 (N_13536,N_12374,N_12765);
and U13537 (N_13537,N_12180,N_12739);
and U13538 (N_13538,N_12306,N_12699);
nand U13539 (N_13539,N_12996,N_12771);
and U13540 (N_13540,N_12481,N_12664);
or U13541 (N_13541,N_12768,N_12100);
or U13542 (N_13542,N_12064,N_12365);
or U13543 (N_13543,N_12686,N_12205);
and U13544 (N_13544,N_12098,N_12750);
and U13545 (N_13545,N_12454,N_12887);
nor U13546 (N_13546,N_12466,N_12911);
nand U13547 (N_13547,N_12740,N_12311);
nor U13548 (N_13548,N_12589,N_12785);
and U13549 (N_13549,N_12798,N_12358);
xnor U13550 (N_13550,N_12362,N_12602);
nand U13551 (N_13551,N_12743,N_12828);
nor U13552 (N_13552,N_12793,N_12148);
or U13553 (N_13553,N_12529,N_12922);
nor U13554 (N_13554,N_12989,N_12860);
or U13555 (N_13555,N_12463,N_12553);
xnor U13556 (N_13556,N_12899,N_12052);
or U13557 (N_13557,N_12856,N_12279);
or U13558 (N_13558,N_12896,N_12244);
xnor U13559 (N_13559,N_12254,N_12982);
or U13560 (N_13560,N_12611,N_12297);
and U13561 (N_13561,N_12811,N_12292);
nor U13562 (N_13562,N_12957,N_12310);
nor U13563 (N_13563,N_12425,N_12068);
nand U13564 (N_13564,N_12468,N_12218);
or U13565 (N_13565,N_12528,N_12725);
and U13566 (N_13566,N_12774,N_12650);
xnor U13567 (N_13567,N_12455,N_12060);
nand U13568 (N_13568,N_12789,N_12238);
nor U13569 (N_13569,N_12046,N_12567);
nand U13570 (N_13570,N_12928,N_12072);
or U13571 (N_13571,N_12428,N_12868);
and U13572 (N_13572,N_12279,N_12313);
and U13573 (N_13573,N_12829,N_12303);
xor U13574 (N_13574,N_12830,N_12278);
nor U13575 (N_13575,N_12275,N_12047);
xnor U13576 (N_13576,N_12644,N_12533);
xor U13577 (N_13577,N_12185,N_12228);
xnor U13578 (N_13578,N_12783,N_12256);
xor U13579 (N_13579,N_12117,N_12725);
nor U13580 (N_13580,N_12501,N_12007);
or U13581 (N_13581,N_12915,N_12752);
nor U13582 (N_13582,N_12238,N_12875);
or U13583 (N_13583,N_12528,N_12640);
nor U13584 (N_13584,N_12080,N_12881);
or U13585 (N_13585,N_12736,N_12908);
nor U13586 (N_13586,N_12104,N_12043);
nor U13587 (N_13587,N_12309,N_12552);
or U13588 (N_13588,N_12711,N_12065);
and U13589 (N_13589,N_12189,N_12845);
or U13590 (N_13590,N_12195,N_12901);
nor U13591 (N_13591,N_12091,N_12512);
nor U13592 (N_13592,N_12247,N_12178);
or U13593 (N_13593,N_12187,N_12994);
nand U13594 (N_13594,N_12025,N_12405);
nor U13595 (N_13595,N_12819,N_12959);
xor U13596 (N_13596,N_12643,N_12906);
xor U13597 (N_13597,N_12493,N_12040);
xnor U13598 (N_13598,N_12067,N_12410);
nor U13599 (N_13599,N_12725,N_12255);
and U13600 (N_13600,N_12991,N_12426);
and U13601 (N_13601,N_12541,N_12976);
or U13602 (N_13602,N_12283,N_12678);
nor U13603 (N_13603,N_12793,N_12819);
or U13604 (N_13604,N_12137,N_12531);
or U13605 (N_13605,N_12621,N_12766);
or U13606 (N_13606,N_12320,N_12227);
or U13607 (N_13607,N_12094,N_12900);
or U13608 (N_13608,N_12021,N_12720);
nor U13609 (N_13609,N_12433,N_12716);
nand U13610 (N_13610,N_12145,N_12658);
or U13611 (N_13611,N_12943,N_12655);
xor U13612 (N_13612,N_12178,N_12361);
or U13613 (N_13613,N_12486,N_12556);
xnor U13614 (N_13614,N_12879,N_12402);
nand U13615 (N_13615,N_12079,N_12761);
nand U13616 (N_13616,N_12025,N_12603);
and U13617 (N_13617,N_12764,N_12504);
nand U13618 (N_13618,N_12526,N_12222);
xnor U13619 (N_13619,N_12865,N_12692);
nand U13620 (N_13620,N_12761,N_12206);
xor U13621 (N_13621,N_12243,N_12656);
xor U13622 (N_13622,N_12942,N_12415);
and U13623 (N_13623,N_12941,N_12313);
xnor U13624 (N_13624,N_12501,N_12195);
or U13625 (N_13625,N_12881,N_12072);
xor U13626 (N_13626,N_12664,N_12596);
or U13627 (N_13627,N_12729,N_12260);
nand U13628 (N_13628,N_12994,N_12283);
nor U13629 (N_13629,N_12905,N_12569);
or U13630 (N_13630,N_12766,N_12511);
xor U13631 (N_13631,N_12280,N_12344);
and U13632 (N_13632,N_12720,N_12669);
nand U13633 (N_13633,N_12319,N_12000);
nand U13634 (N_13634,N_12993,N_12005);
xor U13635 (N_13635,N_12105,N_12997);
xor U13636 (N_13636,N_12734,N_12581);
nor U13637 (N_13637,N_12376,N_12100);
and U13638 (N_13638,N_12791,N_12036);
or U13639 (N_13639,N_12361,N_12548);
or U13640 (N_13640,N_12832,N_12872);
or U13641 (N_13641,N_12666,N_12347);
and U13642 (N_13642,N_12696,N_12384);
nor U13643 (N_13643,N_12036,N_12554);
nor U13644 (N_13644,N_12487,N_12876);
xnor U13645 (N_13645,N_12726,N_12498);
nor U13646 (N_13646,N_12431,N_12223);
nor U13647 (N_13647,N_12137,N_12134);
nor U13648 (N_13648,N_12920,N_12844);
nor U13649 (N_13649,N_12093,N_12223);
and U13650 (N_13650,N_12921,N_12538);
or U13651 (N_13651,N_12327,N_12793);
or U13652 (N_13652,N_12975,N_12726);
xnor U13653 (N_13653,N_12196,N_12674);
nand U13654 (N_13654,N_12830,N_12208);
and U13655 (N_13655,N_12693,N_12682);
or U13656 (N_13656,N_12945,N_12353);
nor U13657 (N_13657,N_12034,N_12363);
nand U13658 (N_13658,N_12814,N_12827);
nor U13659 (N_13659,N_12587,N_12263);
or U13660 (N_13660,N_12864,N_12834);
nand U13661 (N_13661,N_12706,N_12600);
and U13662 (N_13662,N_12719,N_12831);
nand U13663 (N_13663,N_12111,N_12119);
nand U13664 (N_13664,N_12676,N_12501);
xnor U13665 (N_13665,N_12135,N_12892);
nand U13666 (N_13666,N_12584,N_12540);
and U13667 (N_13667,N_12926,N_12664);
xor U13668 (N_13668,N_12069,N_12290);
nand U13669 (N_13669,N_12947,N_12490);
nor U13670 (N_13670,N_12715,N_12477);
and U13671 (N_13671,N_12221,N_12780);
nand U13672 (N_13672,N_12974,N_12606);
or U13673 (N_13673,N_12893,N_12117);
xnor U13674 (N_13674,N_12092,N_12383);
nand U13675 (N_13675,N_12272,N_12815);
nor U13676 (N_13676,N_12369,N_12600);
nor U13677 (N_13677,N_12336,N_12611);
xor U13678 (N_13678,N_12331,N_12351);
or U13679 (N_13679,N_12972,N_12876);
or U13680 (N_13680,N_12647,N_12100);
and U13681 (N_13681,N_12308,N_12093);
and U13682 (N_13682,N_12492,N_12858);
xor U13683 (N_13683,N_12450,N_12769);
or U13684 (N_13684,N_12246,N_12767);
xor U13685 (N_13685,N_12892,N_12595);
nor U13686 (N_13686,N_12394,N_12529);
xor U13687 (N_13687,N_12115,N_12401);
or U13688 (N_13688,N_12776,N_12318);
xor U13689 (N_13689,N_12792,N_12958);
xnor U13690 (N_13690,N_12954,N_12785);
xnor U13691 (N_13691,N_12284,N_12178);
xor U13692 (N_13692,N_12611,N_12627);
and U13693 (N_13693,N_12312,N_12334);
or U13694 (N_13694,N_12346,N_12088);
or U13695 (N_13695,N_12946,N_12291);
nand U13696 (N_13696,N_12280,N_12569);
or U13697 (N_13697,N_12785,N_12444);
and U13698 (N_13698,N_12691,N_12827);
and U13699 (N_13699,N_12932,N_12507);
or U13700 (N_13700,N_12085,N_12605);
nand U13701 (N_13701,N_12379,N_12844);
and U13702 (N_13702,N_12671,N_12515);
nand U13703 (N_13703,N_12539,N_12417);
xnor U13704 (N_13704,N_12182,N_12353);
xnor U13705 (N_13705,N_12495,N_12230);
or U13706 (N_13706,N_12310,N_12241);
or U13707 (N_13707,N_12108,N_12655);
and U13708 (N_13708,N_12647,N_12604);
and U13709 (N_13709,N_12736,N_12698);
xnor U13710 (N_13710,N_12868,N_12971);
and U13711 (N_13711,N_12897,N_12491);
nor U13712 (N_13712,N_12976,N_12238);
nand U13713 (N_13713,N_12009,N_12276);
nand U13714 (N_13714,N_12415,N_12465);
or U13715 (N_13715,N_12981,N_12645);
nand U13716 (N_13716,N_12831,N_12254);
nand U13717 (N_13717,N_12643,N_12602);
nand U13718 (N_13718,N_12054,N_12651);
xor U13719 (N_13719,N_12704,N_12050);
and U13720 (N_13720,N_12361,N_12521);
nor U13721 (N_13721,N_12044,N_12892);
nor U13722 (N_13722,N_12491,N_12062);
and U13723 (N_13723,N_12209,N_12835);
xnor U13724 (N_13724,N_12855,N_12686);
and U13725 (N_13725,N_12635,N_12849);
xnor U13726 (N_13726,N_12715,N_12736);
nand U13727 (N_13727,N_12773,N_12574);
and U13728 (N_13728,N_12871,N_12526);
xnor U13729 (N_13729,N_12606,N_12745);
and U13730 (N_13730,N_12795,N_12451);
nor U13731 (N_13731,N_12982,N_12535);
nand U13732 (N_13732,N_12620,N_12882);
or U13733 (N_13733,N_12605,N_12257);
xor U13734 (N_13734,N_12993,N_12623);
nor U13735 (N_13735,N_12013,N_12755);
xnor U13736 (N_13736,N_12136,N_12759);
nor U13737 (N_13737,N_12969,N_12452);
nand U13738 (N_13738,N_12912,N_12622);
xnor U13739 (N_13739,N_12526,N_12476);
or U13740 (N_13740,N_12940,N_12141);
or U13741 (N_13741,N_12485,N_12951);
or U13742 (N_13742,N_12029,N_12617);
nor U13743 (N_13743,N_12672,N_12577);
nand U13744 (N_13744,N_12875,N_12662);
nor U13745 (N_13745,N_12672,N_12738);
nand U13746 (N_13746,N_12961,N_12968);
nand U13747 (N_13747,N_12134,N_12397);
nor U13748 (N_13748,N_12181,N_12336);
nand U13749 (N_13749,N_12058,N_12481);
and U13750 (N_13750,N_12130,N_12552);
nand U13751 (N_13751,N_12729,N_12690);
or U13752 (N_13752,N_12279,N_12770);
xor U13753 (N_13753,N_12555,N_12118);
and U13754 (N_13754,N_12712,N_12117);
xor U13755 (N_13755,N_12560,N_12761);
or U13756 (N_13756,N_12766,N_12523);
xor U13757 (N_13757,N_12867,N_12664);
or U13758 (N_13758,N_12109,N_12798);
and U13759 (N_13759,N_12454,N_12955);
nand U13760 (N_13760,N_12785,N_12277);
nor U13761 (N_13761,N_12019,N_12146);
and U13762 (N_13762,N_12622,N_12672);
nand U13763 (N_13763,N_12311,N_12440);
xnor U13764 (N_13764,N_12283,N_12848);
nor U13765 (N_13765,N_12455,N_12587);
xnor U13766 (N_13766,N_12422,N_12884);
or U13767 (N_13767,N_12375,N_12113);
nor U13768 (N_13768,N_12147,N_12643);
and U13769 (N_13769,N_12970,N_12628);
nand U13770 (N_13770,N_12164,N_12379);
or U13771 (N_13771,N_12348,N_12161);
xor U13772 (N_13772,N_12903,N_12413);
nand U13773 (N_13773,N_12388,N_12491);
xor U13774 (N_13774,N_12857,N_12434);
nand U13775 (N_13775,N_12470,N_12792);
xor U13776 (N_13776,N_12912,N_12839);
nand U13777 (N_13777,N_12690,N_12989);
nor U13778 (N_13778,N_12644,N_12837);
nand U13779 (N_13779,N_12514,N_12384);
nand U13780 (N_13780,N_12819,N_12842);
nand U13781 (N_13781,N_12712,N_12622);
or U13782 (N_13782,N_12025,N_12790);
and U13783 (N_13783,N_12105,N_12653);
nand U13784 (N_13784,N_12521,N_12559);
nor U13785 (N_13785,N_12583,N_12225);
nor U13786 (N_13786,N_12966,N_12115);
and U13787 (N_13787,N_12658,N_12354);
xnor U13788 (N_13788,N_12651,N_12712);
or U13789 (N_13789,N_12447,N_12234);
or U13790 (N_13790,N_12118,N_12340);
nor U13791 (N_13791,N_12090,N_12019);
and U13792 (N_13792,N_12603,N_12878);
and U13793 (N_13793,N_12535,N_12960);
and U13794 (N_13794,N_12708,N_12201);
and U13795 (N_13795,N_12794,N_12886);
and U13796 (N_13796,N_12899,N_12204);
xnor U13797 (N_13797,N_12717,N_12698);
and U13798 (N_13798,N_12578,N_12494);
or U13799 (N_13799,N_12430,N_12664);
xnor U13800 (N_13800,N_12111,N_12992);
xnor U13801 (N_13801,N_12479,N_12258);
or U13802 (N_13802,N_12187,N_12645);
and U13803 (N_13803,N_12144,N_12698);
or U13804 (N_13804,N_12688,N_12009);
xor U13805 (N_13805,N_12994,N_12496);
nand U13806 (N_13806,N_12277,N_12337);
or U13807 (N_13807,N_12558,N_12334);
or U13808 (N_13808,N_12953,N_12570);
xnor U13809 (N_13809,N_12632,N_12084);
xnor U13810 (N_13810,N_12110,N_12625);
xor U13811 (N_13811,N_12932,N_12619);
nand U13812 (N_13812,N_12598,N_12658);
and U13813 (N_13813,N_12482,N_12467);
or U13814 (N_13814,N_12215,N_12917);
xor U13815 (N_13815,N_12982,N_12666);
or U13816 (N_13816,N_12817,N_12943);
or U13817 (N_13817,N_12014,N_12465);
xor U13818 (N_13818,N_12074,N_12152);
or U13819 (N_13819,N_12552,N_12821);
nand U13820 (N_13820,N_12857,N_12032);
and U13821 (N_13821,N_12192,N_12132);
xnor U13822 (N_13822,N_12174,N_12039);
nand U13823 (N_13823,N_12926,N_12662);
nor U13824 (N_13824,N_12576,N_12403);
nor U13825 (N_13825,N_12370,N_12943);
xor U13826 (N_13826,N_12764,N_12705);
nand U13827 (N_13827,N_12797,N_12451);
nor U13828 (N_13828,N_12821,N_12115);
and U13829 (N_13829,N_12927,N_12911);
xor U13830 (N_13830,N_12152,N_12312);
and U13831 (N_13831,N_12438,N_12313);
nand U13832 (N_13832,N_12039,N_12414);
nor U13833 (N_13833,N_12805,N_12222);
nand U13834 (N_13834,N_12061,N_12877);
nand U13835 (N_13835,N_12279,N_12944);
or U13836 (N_13836,N_12547,N_12114);
nand U13837 (N_13837,N_12565,N_12651);
and U13838 (N_13838,N_12070,N_12407);
xor U13839 (N_13839,N_12078,N_12004);
and U13840 (N_13840,N_12417,N_12382);
nor U13841 (N_13841,N_12984,N_12689);
or U13842 (N_13842,N_12899,N_12651);
nand U13843 (N_13843,N_12186,N_12786);
nand U13844 (N_13844,N_12241,N_12923);
xnor U13845 (N_13845,N_12895,N_12817);
or U13846 (N_13846,N_12214,N_12946);
nor U13847 (N_13847,N_12908,N_12428);
nand U13848 (N_13848,N_12014,N_12989);
nand U13849 (N_13849,N_12602,N_12673);
nand U13850 (N_13850,N_12283,N_12228);
or U13851 (N_13851,N_12233,N_12787);
and U13852 (N_13852,N_12066,N_12736);
nor U13853 (N_13853,N_12873,N_12016);
nor U13854 (N_13854,N_12656,N_12379);
nor U13855 (N_13855,N_12874,N_12751);
or U13856 (N_13856,N_12169,N_12599);
or U13857 (N_13857,N_12996,N_12797);
xnor U13858 (N_13858,N_12008,N_12301);
nand U13859 (N_13859,N_12370,N_12199);
nor U13860 (N_13860,N_12181,N_12426);
and U13861 (N_13861,N_12398,N_12012);
xnor U13862 (N_13862,N_12676,N_12673);
xor U13863 (N_13863,N_12137,N_12077);
and U13864 (N_13864,N_12734,N_12688);
nand U13865 (N_13865,N_12645,N_12883);
xor U13866 (N_13866,N_12893,N_12927);
nor U13867 (N_13867,N_12010,N_12922);
and U13868 (N_13868,N_12241,N_12149);
and U13869 (N_13869,N_12001,N_12411);
nand U13870 (N_13870,N_12410,N_12031);
or U13871 (N_13871,N_12763,N_12401);
nor U13872 (N_13872,N_12121,N_12631);
xnor U13873 (N_13873,N_12416,N_12101);
nor U13874 (N_13874,N_12818,N_12747);
and U13875 (N_13875,N_12690,N_12037);
nand U13876 (N_13876,N_12529,N_12792);
and U13877 (N_13877,N_12138,N_12360);
and U13878 (N_13878,N_12874,N_12577);
xor U13879 (N_13879,N_12394,N_12685);
nand U13880 (N_13880,N_12024,N_12255);
nand U13881 (N_13881,N_12678,N_12384);
xor U13882 (N_13882,N_12024,N_12111);
nand U13883 (N_13883,N_12031,N_12373);
or U13884 (N_13884,N_12468,N_12374);
and U13885 (N_13885,N_12860,N_12391);
nor U13886 (N_13886,N_12319,N_12204);
nand U13887 (N_13887,N_12080,N_12165);
nor U13888 (N_13888,N_12827,N_12631);
or U13889 (N_13889,N_12753,N_12588);
or U13890 (N_13890,N_12584,N_12883);
xor U13891 (N_13891,N_12221,N_12812);
nor U13892 (N_13892,N_12096,N_12170);
or U13893 (N_13893,N_12713,N_12021);
nor U13894 (N_13894,N_12220,N_12192);
and U13895 (N_13895,N_12468,N_12239);
and U13896 (N_13896,N_12622,N_12732);
or U13897 (N_13897,N_12385,N_12333);
nor U13898 (N_13898,N_12733,N_12990);
nor U13899 (N_13899,N_12778,N_12348);
xor U13900 (N_13900,N_12390,N_12429);
nand U13901 (N_13901,N_12159,N_12510);
nand U13902 (N_13902,N_12784,N_12595);
and U13903 (N_13903,N_12551,N_12767);
xnor U13904 (N_13904,N_12511,N_12172);
xor U13905 (N_13905,N_12265,N_12837);
nand U13906 (N_13906,N_12387,N_12987);
nor U13907 (N_13907,N_12620,N_12990);
nand U13908 (N_13908,N_12189,N_12573);
nor U13909 (N_13909,N_12724,N_12155);
nand U13910 (N_13910,N_12018,N_12264);
nand U13911 (N_13911,N_12646,N_12639);
and U13912 (N_13912,N_12929,N_12352);
nor U13913 (N_13913,N_12914,N_12495);
nor U13914 (N_13914,N_12110,N_12694);
or U13915 (N_13915,N_12927,N_12140);
and U13916 (N_13916,N_12656,N_12244);
nand U13917 (N_13917,N_12627,N_12645);
or U13918 (N_13918,N_12926,N_12858);
or U13919 (N_13919,N_12376,N_12020);
nor U13920 (N_13920,N_12983,N_12231);
xor U13921 (N_13921,N_12886,N_12795);
xnor U13922 (N_13922,N_12232,N_12790);
nor U13923 (N_13923,N_12446,N_12524);
xor U13924 (N_13924,N_12497,N_12414);
nand U13925 (N_13925,N_12722,N_12719);
or U13926 (N_13926,N_12537,N_12663);
and U13927 (N_13927,N_12502,N_12745);
nand U13928 (N_13928,N_12687,N_12341);
and U13929 (N_13929,N_12397,N_12697);
nor U13930 (N_13930,N_12713,N_12420);
or U13931 (N_13931,N_12167,N_12516);
nand U13932 (N_13932,N_12551,N_12592);
nor U13933 (N_13933,N_12501,N_12814);
or U13934 (N_13934,N_12716,N_12983);
or U13935 (N_13935,N_12233,N_12379);
or U13936 (N_13936,N_12948,N_12674);
nor U13937 (N_13937,N_12975,N_12625);
xnor U13938 (N_13938,N_12771,N_12859);
nor U13939 (N_13939,N_12565,N_12151);
nor U13940 (N_13940,N_12001,N_12655);
xor U13941 (N_13941,N_12241,N_12054);
or U13942 (N_13942,N_12134,N_12115);
nor U13943 (N_13943,N_12350,N_12523);
nor U13944 (N_13944,N_12011,N_12572);
or U13945 (N_13945,N_12099,N_12494);
and U13946 (N_13946,N_12615,N_12262);
and U13947 (N_13947,N_12855,N_12667);
and U13948 (N_13948,N_12720,N_12269);
xnor U13949 (N_13949,N_12093,N_12698);
xnor U13950 (N_13950,N_12522,N_12826);
nor U13951 (N_13951,N_12535,N_12879);
and U13952 (N_13952,N_12903,N_12811);
and U13953 (N_13953,N_12296,N_12580);
nand U13954 (N_13954,N_12453,N_12924);
xor U13955 (N_13955,N_12396,N_12335);
nand U13956 (N_13956,N_12181,N_12974);
nand U13957 (N_13957,N_12538,N_12199);
or U13958 (N_13958,N_12250,N_12322);
nor U13959 (N_13959,N_12055,N_12392);
xor U13960 (N_13960,N_12240,N_12024);
nand U13961 (N_13961,N_12598,N_12052);
or U13962 (N_13962,N_12903,N_12180);
nor U13963 (N_13963,N_12922,N_12638);
and U13964 (N_13964,N_12356,N_12898);
xnor U13965 (N_13965,N_12706,N_12220);
or U13966 (N_13966,N_12489,N_12602);
xor U13967 (N_13967,N_12535,N_12543);
xnor U13968 (N_13968,N_12335,N_12887);
xor U13969 (N_13969,N_12763,N_12672);
or U13970 (N_13970,N_12989,N_12102);
nand U13971 (N_13971,N_12601,N_12327);
nor U13972 (N_13972,N_12867,N_12610);
or U13973 (N_13973,N_12566,N_12412);
xnor U13974 (N_13974,N_12881,N_12621);
or U13975 (N_13975,N_12521,N_12173);
xor U13976 (N_13976,N_12823,N_12323);
and U13977 (N_13977,N_12104,N_12417);
or U13978 (N_13978,N_12032,N_12023);
nor U13979 (N_13979,N_12338,N_12834);
nand U13980 (N_13980,N_12567,N_12391);
nand U13981 (N_13981,N_12797,N_12722);
nor U13982 (N_13982,N_12712,N_12291);
xnor U13983 (N_13983,N_12627,N_12029);
or U13984 (N_13984,N_12289,N_12240);
xor U13985 (N_13985,N_12469,N_12299);
nand U13986 (N_13986,N_12246,N_12606);
or U13987 (N_13987,N_12672,N_12863);
nand U13988 (N_13988,N_12391,N_12951);
and U13989 (N_13989,N_12316,N_12689);
nor U13990 (N_13990,N_12970,N_12055);
xnor U13991 (N_13991,N_12995,N_12189);
nand U13992 (N_13992,N_12958,N_12225);
nand U13993 (N_13993,N_12119,N_12522);
or U13994 (N_13994,N_12277,N_12062);
and U13995 (N_13995,N_12522,N_12748);
or U13996 (N_13996,N_12802,N_12715);
nand U13997 (N_13997,N_12145,N_12587);
or U13998 (N_13998,N_12471,N_12262);
or U13999 (N_13999,N_12254,N_12237);
or U14000 (N_14000,N_13277,N_13433);
or U14001 (N_14001,N_13973,N_13995);
nand U14002 (N_14002,N_13547,N_13473);
and U14003 (N_14003,N_13145,N_13043);
nor U14004 (N_14004,N_13363,N_13111);
nand U14005 (N_14005,N_13828,N_13093);
nor U14006 (N_14006,N_13164,N_13534);
nand U14007 (N_14007,N_13570,N_13532);
nor U14008 (N_14008,N_13034,N_13374);
and U14009 (N_14009,N_13727,N_13630);
nor U14010 (N_14010,N_13046,N_13495);
nor U14011 (N_14011,N_13471,N_13724);
xor U14012 (N_14012,N_13704,N_13010);
and U14013 (N_14013,N_13530,N_13194);
nor U14014 (N_14014,N_13737,N_13291);
nand U14015 (N_14015,N_13982,N_13065);
nand U14016 (N_14016,N_13347,N_13193);
nor U14017 (N_14017,N_13875,N_13036);
xnor U14018 (N_14018,N_13684,N_13083);
xor U14019 (N_14019,N_13538,N_13814);
nor U14020 (N_14020,N_13930,N_13897);
nand U14021 (N_14021,N_13966,N_13574);
nor U14022 (N_14022,N_13493,N_13186);
nor U14023 (N_14023,N_13149,N_13414);
xor U14024 (N_14024,N_13185,N_13019);
nand U14025 (N_14025,N_13263,N_13925);
or U14026 (N_14026,N_13183,N_13654);
xnor U14027 (N_14027,N_13406,N_13513);
or U14028 (N_14028,N_13954,N_13343);
nand U14029 (N_14029,N_13572,N_13494);
nor U14030 (N_14030,N_13150,N_13861);
or U14031 (N_14031,N_13795,N_13319);
xor U14032 (N_14032,N_13753,N_13822);
and U14033 (N_14033,N_13154,N_13956);
nor U14034 (N_14034,N_13090,N_13222);
or U14035 (N_14035,N_13799,N_13415);
xnor U14036 (N_14036,N_13215,N_13793);
nor U14037 (N_14037,N_13801,N_13927);
and U14038 (N_14038,N_13445,N_13352);
and U14039 (N_14039,N_13564,N_13477);
or U14040 (N_14040,N_13688,N_13628);
and U14041 (N_14041,N_13082,N_13266);
and U14042 (N_14042,N_13329,N_13852);
nand U14043 (N_14043,N_13562,N_13696);
xnor U14044 (N_14044,N_13555,N_13812);
xor U14045 (N_14045,N_13606,N_13807);
or U14046 (N_14046,N_13219,N_13836);
nor U14047 (N_14047,N_13057,N_13529);
and U14048 (N_14048,N_13965,N_13718);
or U14049 (N_14049,N_13693,N_13617);
and U14050 (N_14050,N_13285,N_13980);
and U14051 (N_14051,N_13928,N_13269);
or U14052 (N_14052,N_13134,N_13012);
xnor U14053 (N_14053,N_13069,N_13674);
nor U14054 (N_14054,N_13869,N_13197);
and U14055 (N_14055,N_13054,N_13881);
or U14056 (N_14056,N_13413,N_13049);
or U14057 (N_14057,N_13993,N_13920);
and U14058 (N_14058,N_13857,N_13620);
or U14059 (N_14059,N_13220,N_13158);
nor U14060 (N_14060,N_13166,N_13138);
and U14061 (N_14061,N_13450,N_13479);
nand U14062 (N_14062,N_13227,N_13207);
and U14063 (N_14063,N_13748,N_13039);
or U14064 (N_14064,N_13451,N_13307);
xnor U14065 (N_14065,N_13863,N_13217);
nand U14066 (N_14066,N_13761,N_13751);
or U14067 (N_14067,N_13366,N_13918);
nand U14068 (N_14068,N_13978,N_13786);
xnor U14069 (N_14069,N_13058,N_13976);
nor U14070 (N_14070,N_13528,N_13026);
xor U14071 (N_14071,N_13951,N_13489);
xnor U14072 (N_14072,N_13360,N_13434);
or U14073 (N_14073,N_13330,N_13949);
xnor U14074 (N_14074,N_13962,N_13270);
or U14075 (N_14075,N_13084,N_13959);
nor U14076 (N_14076,N_13755,N_13905);
xnor U14077 (N_14077,N_13264,N_13350);
or U14078 (N_14078,N_13757,N_13779);
xnor U14079 (N_14079,N_13236,N_13539);
and U14080 (N_14080,N_13323,N_13018);
nor U14081 (N_14081,N_13913,N_13576);
xor U14082 (N_14082,N_13017,N_13624);
nand U14083 (N_14083,N_13732,N_13651);
nor U14084 (N_14084,N_13212,N_13712);
and U14085 (N_14085,N_13563,N_13253);
and U14086 (N_14086,N_13963,N_13256);
nand U14087 (N_14087,N_13311,N_13989);
nor U14088 (N_14088,N_13697,N_13108);
and U14089 (N_14089,N_13646,N_13802);
or U14090 (N_14090,N_13225,N_13671);
or U14091 (N_14091,N_13496,N_13669);
or U14092 (N_14092,N_13664,N_13475);
nand U14093 (N_14093,N_13364,N_13052);
and U14094 (N_14094,N_13623,N_13890);
or U14095 (N_14095,N_13171,N_13005);
xor U14096 (N_14096,N_13419,N_13556);
xnor U14097 (N_14097,N_13522,N_13680);
nor U14098 (N_14098,N_13250,N_13791);
and U14099 (N_14099,N_13463,N_13432);
and U14100 (N_14100,N_13768,N_13118);
nand U14101 (N_14101,N_13206,N_13817);
xor U14102 (N_14102,N_13068,N_13862);
xnor U14103 (N_14103,N_13866,N_13089);
or U14104 (N_14104,N_13251,N_13660);
xnor U14105 (N_14105,N_13454,N_13957);
nand U14106 (N_14106,N_13540,N_13213);
xnor U14107 (N_14107,N_13709,N_13914);
nand U14108 (N_14108,N_13749,N_13009);
and U14109 (N_14109,N_13731,N_13879);
and U14110 (N_14110,N_13701,N_13594);
or U14111 (N_14111,N_13125,N_13591);
nor U14112 (N_14112,N_13355,N_13716);
nor U14113 (N_14113,N_13932,N_13910);
nor U14114 (N_14114,N_13868,N_13754);
nor U14115 (N_14115,N_13232,N_13103);
xnor U14116 (N_14116,N_13784,N_13760);
and U14117 (N_14117,N_13279,N_13580);
xor U14118 (N_14118,N_13602,N_13066);
nand U14119 (N_14119,N_13014,N_13242);
xnor U14120 (N_14120,N_13015,N_13675);
and U14121 (N_14121,N_13805,N_13705);
xor U14122 (N_14122,N_13518,N_13265);
and U14123 (N_14123,N_13127,N_13393);
and U14124 (N_14124,N_13211,N_13707);
nor U14125 (N_14125,N_13990,N_13521);
xnor U14126 (N_14126,N_13899,N_13315);
and U14127 (N_14127,N_13934,N_13258);
and U14128 (N_14128,N_13045,N_13417);
and U14129 (N_14129,N_13173,N_13523);
xor U14130 (N_14130,N_13723,N_13614);
or U14131 (N_14131,N_13783,N_13105);
nor U14132 (N_14132,N_13611,N_13072);
nor U14133 (N_14133,N_13887,N_13581);
nor U14134 (N_14134,N_13179,N_13498);
xnor U14135 (N_14135,N_13923,N_13334);
xor U14136 (N_14136,N_13616,N_13703);
nor U14137 (N_14137,N_13509,N_13850);
and U14138 (N_14138,N_13508,N_13059);
xor U14139 (N_14139,N_13661,N_13855);
nor U14140 (N_14140,N_13273,N_13953);
and U14141 (N_14141,N_13441,N_13283);
or U14142 (N_14142,N_13968,N_13667);
xor U14143 (N_14143,N_13060,N_13790);
or U14144 (N_14144,N_13140,N_13048);
nand U14145 (N_14145,N_13035,N_13235);
nand U14146 (N_14146,N_13621,N_13744);
nand U14147 (N_14147,N_13935,N_13029);
xor U14148 (N_14148,N_13176,N_13759);
and U14149 (N_14149,N_13734,N_13300);
nor U14150 (N_14150,N_13603,N_13367);
and U14151 (N_14151,N_13794,N_13497);
xor U14152 (N_14152,N_13991,N_13998);
xor U14153 (N_14153,N_13711,N_13804);
or U14154 (N_14154,N_13798,N_13040);
nor U14155 (N_14155,N_13136,N_13823);
or U14156 (N_14156,N_13764,N_13296);
and U14157 (N_14157,N_13245,N_13524);
xnor U14158 (N_14158,N_13372,N_13486);
or U14159 (N_14159,N_13061,N_13595);
or U14160 (N_14160,N_13738,N_13337);
xor U14161 (N_14161,N_13815,N_13342);
nand U14162 (N_14162,N_13357,N_13032);
xor U14163 (N_14163,N_13573,N_13199);
or U14164 (N_14164,N_13947,N_13946);
nor U14165 (N_14165,N_13282,N_13637);
nand U14166 (N_14166,N_13420,N_13062);
nor U14167 (N_14167,N_13233,N_13668);
or U14168 (N_14168,N_13682,N_13865);
or U14169 (N_14169,N_13690,N_13933);
and U14170 (N_14170,N_13608,N_13520);
nand U14171 (N_14171,N_13402,N_13379);
xnor U14172 (N_14172,N_13666,N_13728);
nor U14173 (N_14173,N_13588,N_13501);
nor U14174 (N_14174,N_13948,N_13557);
nand U14175 (N_14175,N_13305,N_13871);
or U14176 (N_14176,N_13437,N_13986);
nand U14177 (N_14177,N_13468,N_13161);
nand U14178 (N_14178,N_13605,N_13338);
nor U14179 (N_14179,N_13829,N_13351);
nor U14180 (N_14180,N_13182,N_13849);
xor U14181 (N_14181,N_13299,N_13346);
and U14182 (N_14182,N_13792,N_13845);
nand U14183 (N_14183,N_13888,N_13558);
nor U14184 (N_14184,N_13657,N_13101);
xor U14185 (N_14185,N_13915,N_13770);
nand U14186 (N_14186,N_13559,N_13882);
xor U14187 (N_14187,N_13370,N_13885);
xor U14188 (N_14188,N_13536,N_13649);
or U14189 (N_14189,N_13774,N_13141);
nand U14190 (N_14190,N_13604,N_13729);
or U14191 (N_14191,N_13846,N_13816);
nand U14192 (N_14192,N_13478,N_13387);
nor U14193 (N_14193,N_13984,N_13365);
nand U14194 (N_14194,N_13788,N_13597);
or U14195 (N_14195,N_13272,N_13892);
xnor U14196 (N_14196,N_13924,N_13544);
nand U14197 (N_14197,N_13230,N_13808);
and U14198 (N_14198,N_13598,N_13492);
nor U14199 (N_14199,N_13169,N_13552);
or U14200 (N_14200,N_13455,N_13067);
nand U14201 (N_14201,N_13025,N_13535);
and U14202 (N_14202,N_13440,N_13821);
or U14203 (N_14203,N_13135,N_13405);
and U14204 (N_14204,N_13702,N_13255);
or U14205 (N_14205,N_13908,N_13571);
nand U14206 (N_14206,N_13516,N_13710);
xor U14207 (N_14207,N_13326,N_13988);
and U14208 (N_14208,N_13316,N_13038);
or U14209 (N_14209,N_13271,N_13904);
or U14210 (N_14210,N_13099,N_13943);
nor U14211 (N_14211,N_13607,N_13113);
nor U14212 (N_14212,N_13047,N_13244);
or U14213 (N_14213,N_13175,N_13708);
nor U14214 (N_14214,N_13359,N_13683);
nor U14215 (N_14215,N_13027,N_13579);
or U14216 (N_14216,N_13126,N_13781);
nor U14217 (N_14217,N_13332,N_13361);
nand U14218 (N_14218,N_13331,N_13385);
and U14219 (N_14219,N_13304,N_13488);
nor U14220 (N_14220,N_13819,N_13502);
nand U14221 (N_14221,N_13964,N_13527);
and U14222 (N_14222,N_13349,N_13985);
nor U14223 (N_14223,N_13378,N_13028);
or U14224 (N_14224,N_13411,N_13726);
nand U14225 (N_14225,N_13587,N_13839);
and U14226 (N_14226,N_13741,N_13511);
nand U14227 (N_14227,N_13458,N_13833);
and U14228 (N_14228,N_13599,N_13268);
nand U14229 (N_14229,N_13635,N_13132);
nand U14230 (N_14230,N_13131,N_13053);
xor U14231 (N_14231,N_13686,N_13813);
nand U14232 (N_14232,N_13714,N_13916);
xor U14233 (N_14233,N_13421,N_13425);
nor U14234 (N_14234,N_13457,N_13842);
and U14235 (N_14235,N_13358,N_13292);
xor U14236 (N_14236,N_13546,N_13577);
xnor U14237 (N_14237,N_13678,N_13961);
nor U14238 (N_14238,N_13583,N_13006);
and U14239 (N_14239,N_13446,N_13567);
nor U14240 (N_14240,N_13835,N_13214);
nand U14241 (N_14241,N_13341,N_13950);
nor U14242 (N_14242,N_13389,N_13643);
or U14243 (N_14243,N_13837,N_13593);
xor U14244 (N_14244,N_13545,N_13549);
or U14245 (N_14245,N_13187,N_13626);
xor U14246 (N_14246,N_13080,N_13767);
xnor U14247 (N_14247,N_13160,N_13143);
nand U14248 (N_14248,N_13022,N_13515);
nor U14249 (N_14249,N_13384,N_13582);
and U14250 (N_14250,N_13130,N_13771);
and U14251 (N_14251,N_13841,N_13864);
and U14252 (N_14252,N_13172,N_13876);
nor U14253 (N_14253,N_13644,N_13936);
xnor U14254 (N_14254,N_13344,N_13736);
and U14255 (N_14255,N_13706,N_13640);
nor U14256 (N_14256,N_13809,N_13151);
and U14257 (N_14257,N_13123,N_13720);
nor U14258 (N_14258,N_13191,N_13873);
nor U14259 (N_14259,N_13368,N_13306);
nor U14260 (N_14260,N_13153,N_13645);
and U14261 (N_14261,N_13972,N_13878);
nand U14262 (N_14262,N_13408,N_13431);
or U14263 (N_14263,N_13838,N_13237);
nor U14264 (N_14264,N_13952,N_13653);
xnor U14265 (N_14265,N_13743,N_13147);
or U14266 (N_14266,N_13403,N_13204);
nand U14267 (N_14267,N_13003,N_13224);
or U14268 (N_14268,N_13137,N_13551);
or U14269 (N_14269,N_13485,N_13938);
nand U14270 (N_14270,N_13554,N_13261);
nor U14271 (N_14271,N_13994,N_13210);
and U14272 (N_14272,N_13426,N_13503);
xnor U14273 (N_14273,N_13853,N_13100);
nand U14274 (N_14274,N_13380,N_13159);
nand U14275 (N_14275,N_13505,N_13373);
nor U14276 (N_14276,N_13321,N_13397);
xnor U14277 (N_14277,N_13618,N_13248);
nand U14278 (N_14278,N_13023,N_13129);
xor U14279 (N_14279,N_13676,N_13955);
xor U14280 (N_14280,N_13202,N_13730);
or U14281 (N_14281,N_13880,N_13257);
or U14282 (N_14282,N_13267,N_13252);
or U14283 (N_14283,N_13911,N_13464);
nor U14284 (N_14284,N_13088,N_13531);
nand U14285 (N_14285,N_13806,N_13785);
xnor U14286 (N_14286,N_13107,N_13362);
nand U14287 (N_14287,N_13410,N_13917);
and U14288 (N_14288,N_13525,N_13238);
nor U14289 (N_14289,N_13655,N_13262);
nor U14290 (N_14290,N_13778,N_13625);
and U14291 (N_14291,N_13124,N_13700);
or U14292 (N_14292,N_13165,N_13746);
and U14293 (N_14293,N_13466,N_13647);
nand U14294 (N_14294,N_13001,N_13996);
nand U14295 (N_14295,N_13412,N_13076);
or U14296 (N_14296,N_13750,N_13601);
nand U14297 (N_14297,N_13184,N_13490);
and U14298 (N_14298,N_13320,N_13416);
nor U14299 (N_14299,N_13223,N_13286);
and U14300 (N_14300,N_13939,N_13484);
and U14301 (N_14301,N_13290,N_13717);
and U14302 (N_14302,N_13423,N_13428);
nor U14303 (N_14303,N_13476,N_13922);
nand U14304 (N_14304,N_13699,N_13803);
nand U14305 (N_14305,N_13997,N_13831);
xnor U14306 (N_14306,N_13243,N_13152);
or U14307 (N_14307,N_13340,N_13533);
nor U14308 (N_14308,N_13071,N_13691);
and U14309 (N_14309,N_13177,N_13287);
and U14310 (N_14310,N_13826,N_13309);
xnor U14311 (N_14311,N_13526,N_13575);
and U14312 (N_14312,N_13339,N_13336);
and U14313 (N_14313,N_13568,N_13399);
or U14314 (N_14314,N_13335,N_13418);
nand U14315 (N_14315,N_13438,N_13470);
or U14316 (N_14316,N_13313,N_13375);
nor U14317 (N_14317,N_13896,N_13979);
xnor U14318 (N_14318,N_13274,N_13942);
and U14319 (N_14319,N_13190,N_13247);
nor U14320 (N_14320,N_13293,N_13900);
or U14321 (N_14321,N_13391,N_13453);
nor U14322 (N_14322,N_13241,N_13436);
nand U14323 (N_14323,N_13877,N_13325);
nor U14324 (N_14324,N_13740,N_13481);
xnor U14325 (N_14325,N_13456,N_13912);
and U14326 (N_14326,N_13376,N_13442);
xnor U14327 (N_14327,N_13514,N_13480);
nor U14328 (N_14328,N_13085,N_13613);
or U14329 (N_14329,N_13112,N_13318);
and U14330 (N_14330,N_13081,N_13208);
nand U14331 (N_14331,N_13079,N_13281);
and U14332 (N_14332,N_13312,N_13443);
xnor U14333 (N_14333,N_13584,N_13181);
and U14334 (N_14334,N_13310,N_13847);
or U14335 (N_14335,N_13078,N_13926);
or U14336 (N_14336,N_13596,N_13196);
or U14337 (N_14337,N_13317,N_13919);
or U14338 (N_14338,N_13507,N_13400);
xnor U14339 (N_14339,N_13632,N_13077);
and U14340 (N_14340,N_13109,N_13627);
nor U14341 (N_14341,N_13940,N_13610);
and U14342 (N_14342,N_13681,N_13745);
xnor U14343 (N_14343,N_13569,N_13992);
or U14344 (N_14344,N_13094,N_13452);
nand U14345 (N_14345,N_13328,N_13280);
nand U14346 (N_14346,N_13371,N_13119);
and U14347 (N_14347,N_13465,N_13860);
xor U14348 (N_14348,N_13429,N_13142);
xnor U14349 (N_14349,N_13658,N_13000);
or U14350 (N_14350,N_13685,N_13752);
or U14351 (N_14351,N_13561,N_13776);
and U14352 (N_14352,N_13369,N_13636);
nor U14353 (N_14353,N_13687,N_13504);
nand U14354 (N_14354,N_13506,N_13472);
nand U14355 (N_14355,N_13578,N_13157);
or U14356 (N_14356,N_13091,N_13007);
xnor U14357 (N_14357,N_13016,N_13780);
and U14358 (N_14358,N_13301,N_13381);
nand U14359 (N_14359,N_13324,N_13333);
nand U14360 (N_14360,N_13162,N_13097);
or U14361 (N_14361,N_13641,N_13075);
nor U14362 (N_14362,N_13677,N_13874);
nor U14363 (N_14363,N_13216,N_13500);
or U14364 (N_14364,N_13543,N_13859);
or U14365 (N_14365,N_13469,N_13218);
or U14366 (N_14366,N_13353,N_13987);
or U14367 (N_14367,N_13308,N_13548);
or U14368 (N_14368,N_13840,N_13585);
nand U14369 (N_14369,N_13763,N_13971);
xor U14370 (N_14370,N_13758,N_13030);
xor U14371 (N_14371,N_13246,N_13168);
or U14372 (N_14372,N_13715,N_13021);
or U14373 (N_14373,N_13474,N_13024);
nor U14374 (N_14374,N_13354,N_13037);
nor U14375 (N_14375,N_13872,N_13095);
and U14376 (N_14376,N_13944,N_13612);
xnor U14377 (N_14377,N_13074,N_13903);
xor U14378 (N_14378,N_13102,N_13189);
or U14379 (N_14379,N_13725,N_13844);
nor U14380 (N_14380,N_13114,N_13435);
or U14381 (N_14381,N_13600,N_13827);
or U14382 (N_14382,N_13388,N_13008);
nor U14383 (N_14383,N_13377,N_13180);
and U14384 (N_14384,N_13541,N_13073);
and U14385 (N_14385,N_13797,N_13044);
xnor U14386 (N_14386,N_13200,N_13519);
nand U14387 (N_14387,N_13483,N_13459);
and U14388 (N_14388,N_13769,N_13395);
nand U14389 (N_14389,N_13834,N_13884);
nor U14390 (N_14390,N_13619,N_13974);
or U14391 (N_14391,N_13448,N_13106);
nand U14392 (N_14392,N_13692,N_13295);
xor U14393 (N_14393,N_13775,N_13228);
and U14394 (N_14394,N_13122,N_13401);
nor U14395 (N_14395,N_13345,N_13120);
nor U14396 (N_14396,N_13139,N_13195);
or U14397 (N_14397,N_13422,N_13133);
and U14398 (N_14398,N_13394,N_13777);
and U14399 (N_14399,N_13670,N_13772);
and U14400 (N_14400,N_13178,N_13733);
xnor U14401 (N_14401,N_13883,N_13055);
nand U14402 (N_14402,N_13977,N_13735);
or U14403 (N_14403,N_13820,N_13694);
nor U14404 (N_14404,N_13205,N_13742);
nand U14405 (N_14405,N_13303,N_13542);
xor U14406 (N_14406,N_13648,N_13889);
or U14407 (N_14407,N_13960,N_13921);
and U14408 (N_14408,N_13652,N_13398);
nor U14409 (N_14409,N_13893,N_13537);
xor U14410 (N_14410,N_13895,N_13294);
and U14411 (N_14411,N_13592,N_13560);
and U14412 (N_14412,N_13396,N_13510);
nor U14413 (N_14413,N_13392,N_13020);
xor U14414 (N_14414,N_13382,N_13383);
and U14415 (N_14415,N_13656,N_13999);
xnor U14416 (N_14416,N_13444,N_13086);
xor U14417 (N_14417,N_13221,N_13589);
nand U14418 (N_14418,N_13449,N_13121);
xor U14419 (N_14419,N_13631,N_13969);
or U14420 (N_14420,N_13689,N_13615);
nor U14421 (N_14421,N_13260,N_13096);
and U14422 (N_14422,N_13240,N_13234);
and U14423 (N_14423,N_13945,N_13843);
nand U14424 (N_14424,N_13239,N_13155);
or U14425 (N_14425,N_13832,N_13586);
and U14426 (N_14426,N_13856,N_13051);
nand U14427 (N_14427,N_13789,N_13642);
or U14428 (N_14428,N_13170,N_13314);
nor U14429 (N_14429,N_13116,N_13174);
nand U14430 (N_14430,N_13629,N_13226);
or U14431 (N_14431,N_13633,N_13275);
xor U14432 (N_14432,N_13787,N_13407);
nand U14433 (N_14433,N_13144,N_13854);
nand U14434 (N_14434,N_13163,N_13722);
nand U14435 (N_14435,N_13851,N_13092);
and U14436 (N_14436,N_13858,N_13115);
or U14437 (N_14437,N_13302,N_13739);
xnor U14438 (N_14438,N_13609,N_13013);
or U14439 (N_14439,N_13698,N_13713);
nand U14440 (N_14440,N_13482,N_13983);
nor U14441 (N_14441,N_13663,N_13461);
and U14442 (N_14442,N_13259,N_13278);
nor U14443 (N_14443,N_13886,N_13356);
xnor U14444 (N_14444,N_13229,N_13941);
nor U14445 (N_14445,N_13042,N_13662);
xor U14446 (N_14446,N_13937,N_13870);
nor U14447 (N_14447,N_13297,N_13254);
and U14448 (N_14448,N_13284,N_13128);
nand U14449 (N_14449,N_13198,N_13901);
or U14450 (N_14450,N_13907,N_13231);
nand U14451 (N_14451,N_13929,N_13192);
nor U14452 (N_14452,N_13659,N_13117);
and U14453 (N_14453,N_13638,N_13011);
nor U14454 (N_14454,N_13424,N_13004);
nor U14455 (N_14455,N_13800,N_13512);
and U14456 (N_14456,N_13167,N_13188);
nand U14457 (N_14457,N_13811,N_13818);
or U14458 (N_14458,N_13766,N_13070);
and U14459 (N_14459,N_13467,N_13002);
xor U14460 (N_14460,N_13056,N_13679);
and U14461 (N_14461,N_13902,N_13050);
nor U14462 (N_14462,N_13719,N_13782);
nand U14463 (N_14463,N_13796,N_13146);
xor U14464 (N_14464,N_13386,N_13634);
and U14465 (N_14465,N_13898,N_13430);
and U14466 (N_14466,N_13550,N_13031);
xor U14467 (N_14467,N_13033,N_13439);
or U14468 (N_14468,N_13460,N_13981);
xnor U14469 (N_14469,N_13672,N_13327);
or U14470 (N_14470,N_13462,N_13041);
or U14471 (N_14471,N_13087,N_13098);
xnor U14472 (N_14472,N_13404,N_13156);
nand U14473 (N_14473,N_13665,N_13148);
or U14474 (N_14474,N_13487,N_13298);
nor U14475 (N_14475,N_13830,N_13348);
and U14476 (N_14476,N_13390,N_13931);
nor U14477 (N_14477,N_13427,N_13499);
xnor U14478 (N_14478,N_13566,N_13249);
nand U14479 (N_14479,N_13894,N_13447);
or U14480 (N_14480,N_13756,N_13064);
and U14481 (N_14481,N_13765,N_13975);
or U14482 (N_14482,N_13409,N_13289);
or U14483 (N_14483,N_13891,N_13622);
or U14484 (N_14484,N_13590,N_13773);
nor U14485 (N_14485,N_13650,N_13276);
nand U14486 (N_14486,N_13288,N_13825);
nor U14487 (N_14487,N_13322,N_13810);
or U14488 (N_14488,N_13673,N_13565);
and U14489 (N_14489,N_13203,N_13209);
xnor U14490 (N_14490,N_13491,N_13639);
and U14491 (N_14491,N_13970,N_13958);
nor U14492 (N_14492,N_13553,N_13967);
and U14493 (N_14493,N_13110,N_13517);
and U14494 (N_14494,N_13747,N_13824);
and U14495 (N_14495,N_13721,N_13762);
nor U14496 (N_14496,N_13909,N_13695);
nor U14497 (N_14497,N_13201,N_13906);
nand U14498 (N_14498,N_13867,N_13848);
and U14499 (N_14499,N_13063,N_13104);
nand U14500 (N_14500,N_13768,N_13459);
nand U14501 (N_14501,N_13311,N_13132);
nand U14502 (N_14502,N_13110,N_13689);
and U14503 (N_14503,N_13396,N_13819);
xor U14504 (N_14504,N_13217,N_13519);
xnor U14505 (N_14505,N_13553,N_13408);
nor U14506 (N_14506,N_13474,N_13919);
or U14507 (N_14507,N_13514,N_13518);
xor U14508 (N_14508,N_13607,N_13579);
nor U14509 (N_14509,N_13748,N_13254);
nand U14510 (N_14510,N_13132,N_13175);
nor U14511 (N_14511,N_13428,N_13347);
xnor U14512 (N_14512,N_13964,N_13663);
nand U14513 (N_14513,N_13649,N_13503);
nor U14514 (N_14514,N_13746,N_13161);
xor U14515 (N_14515,N_13508,N_13348);
nor U14516 (N_14516,N_13974,N_13402);
nor U14517 (N_14517,N_13575,N_13321);
xnor U14518 (N_14518,N_13134,N_13464);
xnor U14519 (N_14519,N_13560,N_13358);
nor U14520 (N_14520,N_13231,N_13450);
or U14521 (N_14521,N_13761,N_13182);
and U14522 (N_14522,N_13342,N_13201);
xor U14523 (N_14523,N_13635,N_13452);
nand U14524 (N_14524,N_13731,N_13365);
xnor U14525 (N_14525,N_13540,N_13851);
or U14526 (N_14526,N_13725,N_13769);
nor U14527 (N_14527,N_13566,N_13614);
or U14528 (N_14528,N_13687,N_13820);
and U14529 (N_14529,N_13063,N_13905);
nor U14530 (N_14530,N_13328,N_13723);
xnor U14531 (N_14531,N_13762,N_13083);
and U14532 (N_14532,N_13376,N_13078);
or U14533 (N_14533,N_13031,N_13934);
or U14534 (N_14534,N_13355,N_13207);
and U14535 (N_14535,N_13307,N_13306);
xnor U14536 (N_14536,N_13687,N_13788);
or U14537 (N_14537,N_13152,N_13351);
and U14538 (N_14538,N_13774,N_13278);
or U14539 (N_14539,N_13745,N_13960);
nand U14540 (N_14540,N_13408,N_13468);
nor U14541 (N_14541,N_13784,N_13456);
nor U14542 (N_14542,N_13187,N_13520);
nor U14543 (N_14543,N_13284,N_13867);
and U14544 (N_14544,N_13970,N_13369);
nand U14545 (N_14545,N_13698,N_13353);
xnor U14546 (N_14546,N_13742,N_13258);
xor U14547 (N_14547,N_13302,N_13545);
and U14548 (N_14548,N_13983,N_13365);
xor U14549 (N_14549,N_13594,N_13957);
nand U14550 (N_14550,N_13151,N_13935);
and U14551 (N_14551,N_13578,N_13298);
or U14552 (N_14552,N_13147,N_13040);
or U14553 (N_14553,N_13154,N_13629);
xor U14554 (N_14554,N_13065,N_13383);
and U14555 (N_14555,N_13300,N_13878);
or U14556 (N_14556,N_13424,N_13419);
or U14557 (N_14557,N_13948,N_13799);
or U14558 (N_14558,N_13078,N_13036);
and U14559 (N_14559,N_13699,N_13416);
and U14560 (N_14560,N_13301,N_13805);
nand U14561 (N_14561,N_13507,N_13688);
and U14562 (N_14562,N_13661,N_13408);
nor U14563 (N_14563,N_13040,N_13046);
nand U14564 (N_14564,N_13564,N_13191);
xor U14565 (N_14565,N_13834,N_13778);
xnor U14566 (N_14566,N_13563,N_13449);
and U14567 (N_14567,N_13246,N_13369);
or U14568 (N_14568,N_13597,N_13816);
nor U14569 (N_14569,N_13261,N_13256);
nor U14570 (N_14570,N_13321,N_13805);
and U14571 (N_14571,N_13230,N_13618);
and U14572 (N_14572,N_13335,N_13792);
xnor U14573 (N_14573,N_13434,N_13194);
nand U14574 (N_14574,N_13375,N_13248);
xor U14575 (N_14575,N_13415,N_13932);
or U14576 (N_14576,N_13543,N_13637);
nand U14577 (N_14577,N_13915,N_13361);
nand U14578 (N_14578,N_13147,N_13008);
nor U14579 (N_14579,N_13091,N_13742);
nand U14580 (N_14580,N_13582,N_13202);
nand U14581 (N_14581,N_13475,N_13181);
xor U14582 (N_14582,N_13887,N_13335);
nor U14583 (N_14583,N_13133,N_13323);
or U14584 (N_14584,N_13913,N_13795);
xnor U14585 (N_14585,N_13072,N_13434);
and U14586 (N_14586,N_13326,N_13095);
nand U14587 (N_14587,N_13765,N_13618);
and U14588 (N_14588,N_13866,N_13631);
nor U14589 (N_14589,N_13624,N_13795);
and U14590 (N_14590,N_13271,N_13200);
nor U14591 (N_14591,N_13484,N_13874);
and U14592 (N_14592,N_13312,N_13203);
nor U14593 (N_14593,N_13644,N_13278);
or U14594 (N_14594,N_13176,N_13000);
nor U14595 (N_14595,N_13734,N_13104);
or U14596 (N_14596,N_13646,N_13949);
or U14597 (N_14597,N_13238,N_13922);
nor U14598 (N_14598,N_13835,N_13979);
or U14599 (N_14599,N_13315,N_13296);
and U14600 (N_14600,N_13849,N_13506);
xor U14601 (N_14601,N_13613,N_13069);
or U14602 (N_14602,N_13010,N_13373);
and U14603 (N_14603,N_13402,N_13191);
nand U14604 (N_14604,N_13297,N_13174);
nor U14605 (N_14605,N_13814,N_13195);
nand U14606 (N_14606,N_13803,N_13343);
nand U14607 (N_14607,N_13175,N_13551);
or U14608 (N_14608,N_13527,N_13500);
and U14609 (N_14609,N_13148,N_13305);
and U14610 (N_14610,N_13906,N_13765);
xnor U14611 (N_14611,N_13162,N_13475);
xnor U14612 (N_14612,N_13184,N_13866);
and U14613 (N_14613,N_13384,N_13461);
or U14614 (N_14614,N_13651,N_13675);
xor U14615 (N_14615,N_13061,N_13487);
nor U14616 (N_14616,N_13181,N_13721);
nand U14617 (N_14617,N_13772,N_13972);
nor U14618 (N_14618,N_13355,N_13775);
and U14619 (N_14619,N_13212,N_13802);
nand U14620 (N_14620,N_13716,N_13054);
nor U14621 (N_14621,N_13339,N_13441);
or U14622 (N_14622,N_13667,N_13716);
nor U14623 (N_14623,N_13319,N_13624);
nor U14624 (N_14624,N_13109,N_13856);
xor U14625 (N_14625,N_13841,N_13392);
and U14626 (N_14626,N_13183,N_13139);
nor U14627 (N_14627,N_13730,N_13559);
nor U14628 (N_14628,N_13431,N_13740);
nand U14629 (N_14629,N_13356,N_13266);
nand U14630 (N_14630,N_13696,N_13033);
nor U14631 (N_14631,N_13840,N_13823);
or U14632 (N_14632,N_13058,N_13752);
xnor U14633 (N_14633,N_13506,N_13858);
nand U14634 (N_14634,N_13626,N_13900);
nor U14635 (N_14635,N_13139,N_13755);
or U14636 (N_14636,N_13741,N_13474);
nor U14637 (N_14637,N_13976,N_13090);
nand U14638 (N_14638,N_13033,N_13994);
nor U14639 (N_14639,N_13338,N_13996);
xor U14640 (N_14640,N_13340,N_13734);
xor U14641 (N_14641,N_13274,N_13794);
and U14642 (N_14642,N_13659,N_13838);
nor U14643 (N_14643,N_13662,N_13751);
xnor U14644 (N_14644,N_13123,N_13060);
nor U14645 (N_14645,N_13148,N_13559);
and U14646 (N_14646,N_13720,N_13858);
xor U14647 (N_14647,N_13702,N_13886);
and U14648 (N_14648,N_13979,N_13999);
nand U14649 (N_14649,N_13849,N_13592);
xor U14650 (N_14650,N_13822,N_13752);
xor U14651 (N_14651,N_13197,N_13580);
xnor U14652 (N_14652,N_13098,N_13867);
nor U14653 (N_14653,N_13754,N_13215);
and U14654 (N_14654,N_13246,N_13486);
and U14655 (N_14655,N_13635,N_13847);
xnor U14656 (N_14656,N_13096,N_13744);
xnor U14657 (N_14657,N_13260,N_13398);
and U14658 (N_14658,N_13493,N_13145);
xnor U14659 (N_14659,N_13279,N_13989);
nand U14660 (N_14660,N_13313,N_13132);
nor U14661 (N_14661,N_13925,N_13188);
nor U14662 (N_14662,N_13405,N_13384);
nand U14663 (N_14663,N_13552,N_13037);
nor U14664 (N_14664,N_13034,N_13206);
and U14665 (N_14665,N_13751,N_13277);
nand U14666 (N_14666,N_13692,N_13342);
xor U14667 (N_14667,N_13898,N_13998);
or U14668 (N_14668,N_13300,N_13847);
and U14669 (N_14669,N_13040,N_13375);
xor U14670 (N_14670,N_13537,N_13643);
nor U14671 (N_14671,N_13291,N_13490);
nor U14672 (N_14672,N_13473,N_13099);
and U14673 (N_14673,N_13415,N_13219);
and U14674 (N_14674,N_13907,N_13028);
xor U14675 (N_14675,N_13146,N_13415);
nor U14676 (N_14676,N_13976,N_13514);
nor U14677 (N_14677,N_13573,N_13718);
and U14678 (N_14678,N_13585,N_13240);
and U14679 (N_14679,N_13535,N_13459);
and U14680 (N_14680,N_13021,N_13929);
or U14681 (N_14681,N_13147,N_13944);
xnor U14682 (N_14682,N_13402,N_13923);
xor U14683 (N_14683,N_13648,N_13843);
nor U14684 (N_14684,N_13926,N_13246);
and U14685 (N_14685,N_13224,N_13907);
nor U14686 (N_14686,N_13875,N_13530);
xor U14687 (N_14687,N_13743,N_13722);
xnor U14688 (N_14688,N_13310,N_13889);
nand U14689 (N_14689,N_13541,N_13792);
and U14690 (N_14690,N_13210,N_13085);
nor U14691 (N_14691,N_13657,N_13210);
nor U14692 (N_14692,N_13836,N_13386);
and U14693 (N_14693,N_13131,N_13517);
or U14694 (N_14694,N_13913,N_13145);
xnor U14695 (N_14695,N_13889,N_13155);
and U14696 (N_14696,N_13016,N_13601);
nor U14697 (N_14697,N_13372,N_13555);
and U14698 (N_14698,N_13927,N_13702);
and U14699 (N_14699,N_13032,N_13024);
xor U14700 (N_14700,N_13306,N_13741);
nand U14701 (N_14701,N_13343,N_13133);
nand U14702 (N_14702,N_13098,N_13948);
nand U14703 (N_14703,N_13327,N_13401);
nand U14704 (N_14704,N_13584,N_13786);
and U14705 (N_14705,N_13574,N_13225);
nor U14706 (N_14706,N_13227,N_13707);
nand U14707 (N_14707,N_13272,N_13856);
nand U14708 (N_14708,N_13197,N_13909);
and U14709 (N_14709,N_13476,N_13534);
and U14710 (N_14710,N_13186,N_13263);
nor U14711 (N_14711,N_13913,N_13527);
xor U14712 (N_14712,N_13852,N_13197);
and U14713 (N_14713,N_13850,N_13307);
and U14714 (N_14714,N_13302,N_13962);
nor U14715 (N_14715,N_13418,N_13397);
nand U14716 (N_14716,N_13982,N_13268);
nor U14717 (N_14717,N_13888,N_13593);
nor U14718 (N_14718,N_13601,N_13617);
xnor U14719 (N_14719,N_13144,N_13636);
xnor U14720 (N_14720,N_13233,N_13694);
or U14721 (N_14721,N_13484,N_13074);
nand U14722 (N_14722,N_13879,N_13108);
and U14723 (N_14723,N_13272,N_13196);
nand U14724 (N_14724,N_13059,N_13261);
or U14725 (N_14725,N_13922,N_13913);
nand U14726 (N_14726,N_13800,N_13749);
nand U14727 (N_14727,N_13215,N_13718);
or U14728 (N_14728,N_13872,N_13170);
nand U14729 (N_14729,N_13500,N_13604);
or U14730 (N_14730,N_13832,N_13377);
nand U14731 (N_14731,N_13039,N_13616);
xor U14732 (N_14732,N_13988,N_13359);
nor U14733 (N_14733,N_13233,N_13753);
or U14734 (N_14734,N_13154,N_13858);
nand U14735 (N_14735,N_13689,N_13385);
xnor U14736 (N_14736,N_13401,N_13794);
and U14737 (N_14737,N_13051,N_13467);
xor U14738 (N_14738,N_13105,N_13438);
nor U14739 (N_14739,N_13706,N_13648);
xnor U14740 (N_14740,N_13104,N_13045);
xnor U14741 (N_14741,N_13158,N_13095);
or U14742 (N_14742,N_13265,N_13701);
nand U14743 (N_14743,N_13620,N_13227);
and U14744 (N_14744,N_13960,N_13016);
xor U14745 (N_14745,N_13854,N_13730);
nor U14746 (N_14746,N_13040,N_13699);
and U14747 (N_14747,N_13249,N_13151);
and U14748 (N_14748,N_13285,N_13595);
nor U14749 (N_14749,N_13878,N_13567);
xor U14750 (N_14750,N_13407,N_13262);
nor U14751 (N_14751,N_13646,N_13307);
and U14752 (N_14752,N_13416,N_13792);
or U14753 (N_14753,N_13440,N_13323);
xnor U14754 (N_14754,N_13093,N_13634);
and U14755 (N_14755,N_13399,N_13740);
xnor U14756 (N_14756,N_13430,N_13807);
nor U14757 (N_14757,N_13895,N_13339);
or U14758 (N_14758,N_13929,N_13575);
or U14759 (N_14759,N_13590,N_13223);
nor U14760 (N_14760,N_13007,N_13099);
and U14761 (N_14761,N_13955,N_13660);
nand U14762 (N_14762,N_13593,N_13598);
or U14763 (N_14763,N_13285,N_13704);
or U14764 (N_14764,N_13140,N_13784);
nor U14765 (N_14765,N_13968,N_13427);
xor U14766 (N_14766,N_13666,N_13635);
and U14767 (N_14767,N_13982,N_13129);
nor U14768 (N_14768,N_13608,N_13410);
nand U14769 (N_14769,N_13092,N_13968);
nand U14770 (N_14770,N_13980,N_13258);
or U14771 (N_14771,N_13642,N_13514);
and U14772 (N_14772,N_13086,N_13995);
or U14773 (N_14773,N_13602,N_13528);
nor U14774 (N_14774,N_13720,N_13271);
nor U14775 (N_14775,N_13695,N_13387);
nor U14776 (N_14776,N_13444,N_13281);
xnor U14777 (N_14777,N_13410,N_13060);
and U14778 (N_14778,N_13902,N_13980);
xnor U14779 (N_14779,N_13585,N_13809);
and U14780 (N_14780,N_13547,N_13437);
nor U14781 (N_14781,N_13307,N_13658);
or U14782 (N_14782,N_13822,N_13717);
nor U14783 (N_14783,N_13922,N_13545);
nor U14784 (N_14784,N_13370,N_13113);
and U14785 (N_14785,N_13844,N_13657);
nor U14786 (N_14786,N_13357,N_13592);
nor U14787 (N_14787,N_13774,N_13103);
nand U14788 (N_14788,N_13089,N_13822);
nor U14789 (N_14789,N_13130,N_13404);
xnor U14790 (N_14790,N_13705,N_13437);
or U14791 (N_14791,N_13724,N_13431);
xor U14792 (N_14792,N_13649,N_13174);
or U14793 (N_14793,N_13939,N_13925);
nand U14794 (N_14794,N_13867,N_13493);
xnor U14795 (N_14795,N_13082,N_13941);
xnor U14796 (N_14796,N_13514,N_13024);
nor U14797 (N_14797,N_13439,N_13301);
and U14798 (N_14798,N_13066,N_13734);
and U14799 (N_14799,N_13297,N_13855);
and U14800 (N_14800,N_13430,N_13078);
and U14801 (N_14801,N_13733,N_13021);
nand U14802 (N_14802,N_13316,N_13260);
and U14803 (N_14803,N_13853,N_13408);
nand U14804 (N_14804,N_13235,N_13172);
and U14805 (N_14805,N_13568,N_13417);
and U14806 (N_14806,N_13129,N_13910);
nand U14807 (N_14807,N_13274,N_13272);
or U14808 (N_14808,N_13794,N_13212);
nand U14809 (N_14809,N_13723,N_13427);
and U14810 (N_14810,N_13890,N_13446);
or U14811 (N_14811,N_13747,N_13233);
and U14812 (N_14812,N_13699,N_13214);
and U14813 (N_14813,N_13462,N_13605);
nor U14814 (N_14814,N_13295,N_13788);
xnor U14815 (N_14815,N_13362,N_13461);
xor U14816 (N_14816,N_13541,N_13192);
nor U14817 (N_14817,N_13032,N_13464);
nand U14818 (N_14818,N_13254,N_13955);
and U14819 (N_14819,N_13139,N_13941);
or U14820 (N_14820,N_13366,N_13590);
and U14821 (N_14821,N_13791,N_13038);
nor U14822 (N_14822,N_13965,N_13512);
nor U14823 (N_14823,N_13314,N_13316);
nand U14824 (N_14824,N_13800,N_13763);
or U14825 (N_14825,N_13079,N_13797);
nand U14826 (N_14826,N_13820,N_13073);
nand U14827 (N_14827,N_13841,N_13931);
and U14828 (N_14828,N_13072,N_13762);
xnor U14829 (N_14829,N_13514,N_13280);
nor U14830 (N_14830,N_13310,N_13015);
nor U14831 (N_14831,N_13637,N_13408);
or U14832 (N_14832,N_13152,N_13299);
nand U14833 (N_14833,N_13646,N_13789);
and U14834 (N_14834,N_13202,N_13570);
or U14835 (N_14835,N_13608,N_13997);
xnor U14836 (N_14836,N_13021,N_13623);
xor U14837 (N_14837,N_13100,N_13017);
xnor U14838 (N_14838,N_13921,N_13938);
or U14839 (N_14839,N_13644,N_13070);
or U14840 (N_14840,N_13945,N_13483);
and U14841 (N_14841,N_13020,N_13045);
xnor U14842 (N_14842,N_13994,N_13083);
xor U14843 (N_14843,N_13219,N_13158);
and U14844 (N_14844,N_13767,N_13580);
and U14845 (N_14845,N_13636,N_13374);
nand U14846 (N_14846,N_13781,N_13731);
and U14847 (N_14847,N_13663,N_13040);
nor U14848 (N_14848,N_13962,N_13937);
nand U14849 (N_14849,N_13627,N_13509);
nor U14850 (N_14850,N_13838,N_13260);
or U14851 (N_14851,N_13036,N_13391);
and U14852 (N_14852,N_13912,N_13055);
and U14853 (N_14853,N_13848,N_13297);
xor U14854 (N_14854,N_13103,N_13473);
nor U14855 (N_14855,N_13658,N_13551);
xor U14856 (N_14856,N_13534,N_13184);
nand U14857 (N_14857,N_13285,N_13637);
xor U14858 (N_14858,N_13706,N_13649);
or U14859 (N_14859,N_13103,N_13111);
nand U14860 (N_14860,N_13734,N_13082);
xor U14861 (N_14861,N_13394,N_13248);
and U14862 (N_14862,N_13133,N_13813);
nand U14863 (N_14863,N_13228,N_13370);
and U14864 (N_14864,N_13345,N_13775);
nor U14865 (N_14865,N_13360,N_13249);
nand U14866 (N_14866,N_13183,N_13889);
and U14867 (N_14867,N_13154,N_13408);
xnor U14868 (N_14868,N_13291,N_13032);
nor U14869 (N_14869,N_13410,N_13888);
nor U14870 (N_14870,N_13070,N_13832);
nor U14871 (N_14871,N_13327,N_13790);
nand U14872 (N_14872,N_13903,N_13080);
and U14873 (N_14873,N_13189,N_13239);
nand U14874 (N_14874,N_13603,N_13690);
nand U14875 (N_14875,N_13754,N_13082);
xnor U14876 (N_14876,N_13860,N_13101);
nand U14877 (N_14877,N_13883,N_13819);
and U14878 (N_14878,N_13339,N_13803);
nand U14879 (N_14879,N_13728,N_13676);
nor U14880 (N_14880,N_13876,N_13024);
nand U14881 (N_14881,N_13432,N_13588);
and U14882 (N_14882,N_13104,N_13445);
or U14883 (N_14883,N_13190,N_13849);
nand U14884 (N_14884,N_13498,N_13138);
nor U14885 (N_14885,N_13059,N_13214);
and U14886 (N_14886,N_13356,N_13200);
xnor U14887 (N_14887,N_13789,N_13476);
nand U14888 (N_14888,N_13714,N_13703);
or U14889 (N_14889,N_13830,N_13027);
nand U14890 (N_14890,N_13066,N_13942);
xnor U14891 (N_14891,N_13640,N_13604);
nor U14892 (N_14892,N_13440,N_13478);
nand U14893 (N_14893,N_13615,N_13352);
nor U14894 (N_14894,N_13712,N_13740);
or U14895 (N_14895,N_13691,N_13000);
nand U14896 (N_14896,N_13650,N_13666);
xnor U14897 (N_14897,N_13744,N_13450);
xor U14898 (N_14898,N_13345,N_13172);
or U14899 (N_14899,N_13149,N_13265);
xnor U14900 (N_14900,N_13640,N_13808);
nand U14901 (N_14901,N_13947,N_13198);
and U14902 (N_14902,N_13675,N_13783);
nand U14903 (N_14903,N_13871,N_13523);
nand U14904 (N_14904,N_13804,N_13726);
nand U14905 (N_14905,N_13122,N_13073);
nor U14906 (N_14906,N_13203,N_13014);
or U14907 (N_14907,N_13766,N_13570);
nor U14908 (N_14908,N_13502,N_13433);
xnor U14909 (N_14909,N_13703,N_13355);
and U14910 (N_14910,N_13640,N_13174);
or U14911 (N_14911,N_13854,N_13189);
and U14912 (N_14912,N_13093,N_13987);
nor U14913 (N_14913,N_13657,N_13522);
xor U14914 (N_14914,N_13354,N_13312);
and U14915 (N_14915,N_13212,N_13862);
nor U14916 (N_14916,N_13139,N_13391);
xnor U14917 (N_14917,N_13274,N_13112);
or U14918 (N_14918,N_13098,N_13355);
and U14919 (N_14919,N_13190,N_13932);
nand U14920 (N_14920,N_13366,N_13034);
and U14921 (N_14921,N_13750,N_13969);
or U14922 (N_14922,N_13904,N_13091);
nand U14923 (N_14923,N_13182,N_13926);
xor U14924 (N_14924,N_13189,N_13172);
and U14925 (N_14925,N_13647,N_13239);
or U14926 (N_14926,N_13529,N_13382);
or U14927 (N_14927,N_13831,N_13704);
nand U14928 (N_14928,N_13539,N_13161);
and U14929 (N_14929,N_13766,N_13073);
and U14930 (N_14930,N_13530,N_13860);
and U14931 (N_14931,N_13561,N_13116);
xor U14932 (N_14932,N_13102,N_13302);
nor U14933 (N_14933,N_13212,N_13366);
nor U14934 (N_14934,N_13609,N_13453);
xor U14935 (N_14935,N_13240,N_13932);
xnor U14936 (N_14936,N_13426,N_13274);
and U14937 (N_14937,N_13277,N_13472);
nand U14938 (N_14938,N_13105,N_13209);
or U14939 (N_14939,N_13693,N_13431);
xnor U14940 (N_14940,N_13595,N_13158);
nor U14941 (N_14941,N_13952,N_13333);
or U14942 (N_14942,N_13490,N_13296);
and U14943 (N_14943,N_13220,N_13989);
and U14944 (N_14944,N_13543,N_13315);
nand U14945 (N_14945,N_13768,N_13871);
xor U14946 (N_14946,N_13210,N_13270);
xor U14947 (N_14947,N_13776,N_13630);
xor U14948 (N_14948,N_13005,N_13519);
nand U14949 (N_14949,N_13296,N_13883);
or U14950 (N_14950,N_13261,N_13778);
or U14951 (N_14951,N_13043,N_13921);
or U14952 (N_14952,N_13114,N_13014);
nor U14953 (N_14953,N_13413,N_13082);
and U14954 (N_14954,N_13042,N_13985);
and U14955 (N_14955,N_13309,N_13246);
or U14956 (N_14956,N_13112,N_13901);
xor U14957 (N_14957,N_13075,N_13462);
and U14958 (N_14958,N_13874,N_13204);
xnor U14959 (N_14959,N_13110,N_13024);
nor U14960 (N_14960,N_13874,N_13088);
or U14961 (N_14961,N_13782,N_13904);
nand U14962 (N_14962,N_13601,N_13773);
nand U14963 (N_14963,N_13862,N_13363);
nor U14964 (N_14964,N_13368,N_13371);
and U14965 (N_14965,N_13452,N_13967);
and U14966 (N_14966,N_13048,N_13464);
and U14967 (N_14967,N_13414,N_13932);
nor U14968 (N_14968,N_13841,N_13313);
or U14969 (N_14969,N_13696,N_13856);
nand U14970 (N_14970,N_13612,N_13321);
and U14971 (N_14971,N_13811,N_13631);
nand U14972 (N_14972,N_13001,N_13265);
xor U14973 (N_14973,N_13130,N_13069);
nor U14974 (N_14974,N_13896,N_13956);
and U14975 (N_14975,N_13066,N_13551);
and U14976 (N_14976,N_13516,N_13476);
nand U14977 (N_14977,N_13662,N_13821);
nand U14978 (N_14978,N_13235,N_13505);
or U14979 (N_14979,N_13827,N_13209);
and U14980 (N_14980,N_13008,N_13000);
xnor U14981 (N_14981,N_13782,N_13309);
and U14982 (N_14982,N_13825,N_13578);
or U14983 (N_14983,N_13912,N_13040);
nand U14984 (N_14984,N_13349,N_13944);
nand U14985 (N_14985,N_13825,N_13172);
nor U14986 (N_14986,N_13929,N_13097);
or U14987 (N_14987,N_13587,N_13043);
or U14988 (N_14988,N_13527,N_13715);
xnor U14989 (N_14989,N_13905,N_13005);
nor U14990 (N_14990,N_13687,N_13239);
or U14991 (N_14991,N_13064,N_13239);
xor U14992 (N_14992,N_13236,N_13489);
and U14993 (N_14993,N_13123,N_13376);
xnor U14994 (N_14994,N_13400,N_13202);
and U14995 (N_14995,N_13312,N_13235);
nand U14996 (N_14996,N_13959,N_13269);
or U14997 (N_14997,N_13457,N_13514);
or U14998 (N_14998,N_13237,N_13708);
or U14999 (N_14999,N_13319,N_13625);
xor U15000 (N_15000,N_14085,N_14176);
xnor U15001 (N_15001,N_14999,N_14296);
and U15002 (N_15002,N_14791,N_14720);
or U15003 (N_15003,N_14067,N_14520);
nor U15004 (N_15004,N_14024,N_14097);
and U15005 (N_15005,N_14310,N_14727);
nor U15006 (N_15006,N_14729,N_14361);
nor U15007 (N_15007,N_14429,N_14351);
nand U15008 (N_15008,N_14061,N_14594);
nand U15009 (N_15009,N_14106,N_14491);
xnor U15010 (N_15010,N_14398,N_14741);
nand U15011 (N_15011,N_14707,N_14991);
nand U15012 (N_15012,N_14845,N_14743);
nor U15013 (N_15013,N_14937,N_14156);
and U15014 (N_15014,N_14619,N_14411);
and U15015 (N_15015,N_14812,N_14205);
and U15016 (N_15016,N_14759,N_14464);
and U15017 (N_15017,N_14614,N_14158);
or U15018 (N_15018,N_14955,N_14944);
or U15019 (N_15019,N_14823,N_14073);
or U15020 (N_15020,N_14961,N_14988);
nand U15021 (N_15021,N_14503,N_14080);
nor U15022 (N_15022,N_14826,N_14144);
xnor U15023 (N_15023,N_14328,N_14905);
nand U15024 (N_15024,N_14348,N_14596);
nand U15025 (N_15025,N_14324,N_14957);
and U15026 (N_15026,N_14409,N_14533);
or U15027 (N_15027,N_14781,N_14337);
or U15028 (N_15028,N_14603,N_14753);
or U15029 (N_15029,N_14629,N_14269);
nand U15030 (N_15030,N_14693,N_14213);
xnor U15031 (N_15031,N_14069,N_14399);
xnor U15032 (N_15032,N_14167,N_14347);
and U15033 (N_15033,N_14066,N_14048);
nand U15034 (N_15034,N_14865,N_14873);
and U15035 (N_15035,N_14912,N_14016);
xnor U15036 (N_15036,N_14728,N_14185);
or U15037 (N_15037,N_14768,N_14239);
nand U15038 (N_15038,N_14022,N_14565);
or U15039 (N_15039,N_14881,N_14631);
xnor U15040 (N_15040,N_14730,N_14461);
and U15041 (N_15041,N_14434,N_14457);
and U15042 (N_15042,N_14956,N_14656);
nand U15043 (N_15043,N_14088,N_14612);
xnor U15044 (N_15044,N_14868,N_14815);
nor U15045 (N_15045,N_14018,N_14257);
nand U15046 (N_15046,N_14688,N_14841);
or U15047 (N_15047,N_14618,N_14780);
nor U15048 (N_15048,N_14960,N_14786);
or U15049 (N_15049,N_14009,N_14722);
and U15050 (N_15050,N_14017,N_14810);
nand U15051 (N_15051,N_14314,N_14380);
xor U15052 (N_15052,N_14953,N_14182);
and U15053 (N_15053,N_14668,N_14684);
nor U15054 (N_15054,N_14276,N_14431);
and U15055 (N_15055,N_14173,N_14896);
nand U15056 (N_15056,N_14542,N_14078);
nand U15057 (N_15057,N_14419,N_14968);
or U15058 (N_15058,N_14571,N_14095);
and U15059 (N_15059,N_14280,N_14566);
and U15060 (N_15060,N_14998,N_14825);
xor U15061 (N_15061,N_14330,N_14975);
nor U15062 (N_15062,N_14447,N_14417);
xor U15063 (N_15063,N_14402,N_14083);
nand U15064 (N_15064,N_14426,N_14180);
nand U15065 (N_15065,N_14237,N_14884);
or U15066 (N_15066,N_14654,N_14904);
xor U15067 (N_15067,N_14110,N_14748);
nor U15068 (N_15068,N_14104,N_14371);
nand U15069 (N_15069,N_14861,N_14026);
or U15070 (N_15070,N_14375,N_14844);
nor U15071 (N_15071,N_14444,N_14495);
xor U15072 (N_15072,N_14818,N_14258);
xor U15073 (N_15073,N_14797,N_14293);
and U15074 (N_15074,N_14806,N_14362);
or U15075 (N_15075,N_14057,N_14517);
and U15076 (N_15076,N_14479,N_14400);
and U15077 (N_15077,N_14680,N_14763);
xnor U15078 (N_15078,N_14068,N_14789);
xnor U15079 (N_15079,N_14472,N_14767);
nor U15080 (N_15080,N_14734,N_14385);
nor U15081 (N_15081,N_14485,N_14278);
xnor U15082 (N_15082,N_14949,N_14309);
nor U15083 (N_15083,N_14135,N_14509);
nor U15084 (N_15084,N_14321,N_14271);
or U15085 (N_15085,N_14422,N_14799);
nor U15086 (N_15086,N_14887,N_14672);
nor U15087 (N_15087,N_14383,N_14969);
xnor U15088 (N_15088,N_14289,N_14811);
and U15089 (N_15089,N_14802,N_14248);
or U15090 (N_15090,N_14487,N_14268);
nor U15091 (N_15091,N_14441,N_14723);
nand U15092 (N_15092,N_14139,N_14138);
xor U15093 (N_15093,N_14386,N_14287);
nand U15094 (N_15094,N_14907,N_14519);
and U15095 (N_15095,N_14587,N_14382);
or U15096 (N_15096,N_14948,N_14628);
xnor U15097 (N_15097,N_14794,N_14658);
nand U15098 (N_15098,N_14754,N_14942);
xor U15099 (N_15099,N_14554,N_14625);
xnor U15100 (N_15100,N_14545,N_14240);
nand U15101 (N_15101,N_14558,N_14539);
nand U15102 (N_15102,N_14316,N_14987);
or U15103 (N_15103,N_14186,N_14021);
xnor U15104 (N_15104,N_14506,N_14977);
or U15105 (N_15105,N_14002,N_14690);
nand U15106 (N_15106,N_14200,N_14702);
nand U15107 (N_15107,N_14651,N_14005);
nand U15108 (N_15108,N_14013,N_14535);
xor U15109 (N_15109,N_14890,N_14254);
nand U15110 (N_15110,N_14114,N_14195);
nor U15111 (N_15111,N_14105,N_14401);
xnor U15112 (N_15112,N_14323,N_14164);
nor U15113 (N_15113,N_14776,N_14965);
and U15114 (N_15114,N_14389,N_14032);
nor U15115 (N_15115,N_14169,N_14559);
and U15116 (N_15116,N_14649,N_14994);
or U15117 (N_15117,N_14538,N_14475);
and U15118 (N_15118,N_14130,N_14885);
nand U15119 (N_15119,N_14986,N_14855);
xor U15120 (N_15120,N_14827,N_14121);
nor U15121 (N_15121,N_14007,N_14537);
and U15122 (N_15122,N_14008,N_14893);
nand U15123 (N_15123,N_14196,N_14358);
and U15124 (N_15124,N_14415,N_14548);
and U15125 (N_15125,N_14959,N_14151);
nand U15126 (N_15126,N_14163,N_14642);
nand U15127 (N_15127,N_14427,N_14939);
or U15128 (N_15128,N_14320,N_14072);
or U15129 (N_15129,N_14983,N_14867);
xor U15130 (N_15130,N_14049,N_14604);
nand U15131 (N_15131,N_14172,N_14835);
nor U15132 (N_15132,N_14266,N_14421);
or U15133 (N_15133,N_14911,N_14241);
or U15134 (N_15134,N_14750,N_14997);
xor U15135 (N_15135,N_14458,N_14148);
xor U15136 (N_15136,N_14063,N_14544);
or U15137 (N_15137,N_14100,N_14039);
nor U15138 (N_15138,N_14259,N_14735);
and U15139 (N_15139,N_14368,N_14075);
or U15140 (N_15140,N_14712,N_14635);
or U15141 (N_15141,N_14197,N_14641);
nand U15142 (N_15142,N_14346,N_14384);
xor U15143 (N_15143,N_14663,N_14655);
xnor U15144 (N_15144,N_14489,N_14837);
nor U15145 (N_15145,N_14507,N_14198);
xnor U15146 (N_15146,N_14985,N_14137);
and U15147 (N_15147,N_14101,N_14143);
and U15148 (N_15148,N_14476,N_14504);
xor U15149 (N_15149,N_14123,N_14115);
nand U15150 (N_15150,N_14903,N_14010);
and U15151 (N_15151,N_14037,N_14880);
and U15152 (N_15152,N_14500,N_14602);
xnor U15153 (N_15153,N_14512,N_14046);
nor U15154 (N_15154,N_14670,N_14652);
xor U15155 (N_15155,N_14263,N_14099);
nand U15156 (N_15156,N_14090,N_14440);
and U15157 (N_15157,N_14626,N_14343);
nand U15158 (N_15158,N_14557,N_14521);
xnor U15159 (N_15159,N_14820,N_14952);
nand U15160 (N_15160,N_14660,N_14891);
nand U15161 (N_15161,N_14929,N_14028);
or U15162 (N_15162,N_14225,N_14443);
nand U15163 (N_15163,N_14179,N_14305);
nand U15164 (N_15164,N_14265,N_14665);
xor U15165 (N_15165,N_14681,N_14214);
or U15166 (N_15166,N_14103,N_14919);
or U15167 (N_15167,N_14901,N_14292);
or U15168 (N_15168,N_14313,N_14738);
and U15169 (N_15169,N_14423,N_14875);
and U15170 (N_15170,N_14474,N_14951);
nor U15171 (N_15171,N_14524,N_14562);
xor U15172 (N_15172,N_14395,N_14486);
and U15173 (N_15173,N_14212,N_14771);
nand U15174 (N_15174,N_14803,N_14160);
nor U15175 (N_15175,N_14913,N_14129);
or U15176 (N_15176,N_14247,N_14726);
nand U15177 (N_15177,N_14255,N_14468);
or U15178 (N_15178,N_14192,N_14623);
nand U15179 (N_15179,N_14785,N_14581);
nand U15180 (N_15180,N_14992,N_14019);
nor U15181 (N_15181,N_14677,N_14526);
nand U15182 (N_15182,N_14001,N_14798);
nand U15183 (N_15183,N_14757,N_14071);
and U15184 (N_15184,N_14394,N_14555);
nand U15185 (N_15185,N_14250,N_14459);
nand U15186 (N_15186,N_14393,N_14126);
nand U15187 (N_15187,N_14349,N_14971);
or U15188 (N_15188,N_14369,N_14284);
nor U15189 (N_15189,N_14228,N_14640);
nor U15190 (N_15190,N_14011,N_14601);
nand U15191 (N_15191,N_14168,N_14674);
nor U15192 (N_15192,N_14373,N_14606);
nor U15193 (N_15193,N_14232,N_14588);
or U15194 (N_15194,N_14513,N_14737);
or U15195 (N_15195,N_14838,N_14416);
and U15196 (N_15196,N_14678,N_14854);
and U15197 (N_15197,N_14713,N_14546);
and U15198 (N_15198,N_14570,N_14249);
or U15199 (N_15199,N_14418,N_14940);
or U15200 (N_15200,N_14454,N_14439);
or U15201 (N_15201,N_14575,N_14523);
and U15202 (N_15202,N_14692,N_14062);
or U15203 (N_15203,N_14162,N_14847);
xor U15204 (N_15204,N_14446,N_14208);
xor U15205 (N_15205,N_14270,N_14091);
xor U15206 (N_15206,N_14834,N_14607);
nor U15207 (N_15207,N_14092,N_14831);
nand U15208 (N_15208,N_14215,N_14157);
and U15209 (N_15209,N_14245,N_14227);
nor U15210 (N_15210,N_14033,N_14632);
xnor U15211 (N_15211,N_14332,N_14928);
xor U15212 (N_15212,N_14014,N_14000);
nor U15213 (N_15213,N_14034,N_14877);
nand U15214 (N_15214,N_14125,N_14136);
xnor U15215 (N_15215,N_14897,N_14611);
and U15216 (N_15216,N_14627,N_14600);
or U15217 (N_15217,N_14716,N_14231);
nand U15218 (N_15218,N_14435,N_14808);
nor U15219 (N_15219,N_14433,N_14751);
nand U15220 (N_15220,N_14756,N_14857);
or U15221 (N_15221,N_14989,N_14609);
and U15222 (N_15222,N_14675,N_14696);
nor U15223 (N_15223,N_14664,N_14578);
or U15224 (N_15224,N_14483,N_14059);
or U15225 (N_15225,N_14536,N_14350);
and U15226 (N_15226,N_14899,N_14190);
xor U15227 (N_15227,N_14406,N_14087);
xnor U15228 (N_15228,N_14451,N_14391);
or U15229 (N_15229,N_14849,N_14943);
xnor U15230 (N_15230,N_14954,N_14964);
or U15231 (N_15231,N_14341,N_14866);
and U15232 (N_15232,N_14584,N_14045);
or U15233 (N_15233,N_14982,N_14335);
nor U15234 (N_15234,N_14970,N_14622);
and U15235 (N_15235,N_14437,N_14822);
nor U15236 (N_15236,N_14745,N_14608);
and U15237 (N_15237,N_14731,N_14181);
and U15238 (N_15238,N_14282,N_14807);
xnor U15239 (N_15239,N_14900,N_14084);
or U15240 (N_15240,N_14359,N_14553);
or U15241 (N_15241,N_14824,N_14438);
and U15242 (N_15242,N_14645,N_14442);
nand U15243 (N_15243,N_14921,N_14082);
nand U15244 (N_15244,N_14322,N_14843);
xor U15245 (N_15245,N_14736,N_14089);
nor U15246 (N_15246,N_14445,N_14770);
xor U15247 (N_15247,N_14779,N_14027);
nand U15248 (N_15248,N_14342,N_14315);
nand U15249 (N_15249,N_14869,N_14706);
and U15250 (N_15250,N_14079,N_14209);
nor U15251 (N_15251,N_14428,N_14990);
nor U15252 (N_15252,N_14760,N_14145);
xnor U15253 (N_15253,N_14256,N_14141);
nand U15254 (N_15254,N_14146,N_14211);
nand U15255 (N_15255,N_14119,N_14846);
xnor U15256 (N_15256,N_14593,N_14586);
or U15257 (N_15257,N_14591,N_14221);
nand U15258 (N_15258,N_14892,N_14829);
nor U15259 (N_15259,N_14518,N_14840);
nor U15260 (N_15260,N_14777,N_14908);
xnor U15261 (N_15261,N_14605,N_14993);
nor U15262 (N_15262,N_14804,N_14070);
xor U15263 (N_15263,N_14460,N_14590);
and U15264 (N_15264,N_14345,N_14117);
xor U15265 (N_15265,N_14933,N_14568);
xor U15266 (N_15266,N_14355,N_14783);
xor U15267 (N_15267,N_14790,N_14718);
or U15268 (N_15268,N_14876,N_14326);
or U15269 (N_15269,N_14889,N_14065);
or U15270 (N_15270,N_14294,N_14938);
or U15271 (N_15271,N_14683,N_14187);
xor U15272 (N_15272,N_14772,N_14633);
nor U15273 (N_15273,N_14170,N_14700);
or U15274 (N_15274,N_14295,N_14035);
nand U15275 (N_15275,N_14924,N_14682);
nor U15276 (N_15276,N_14710,N_14872);
nor U15277 (N_15277,N_14381,N_14274);
nand U15278 (N_15278,N_14234,N_14246);
nand U15279 (N_15279,N_14550,N_14004);
nand U15280 (N_15280,N_14450,N_14592);
or U15281 (N_15281,N_14492,N_14410);
nor U15282 (N_15282,N_14895,N_14556);
nor U15283 (N_15283,N_14661,N_14188);
and U15284 (N_15284,N_14177,N_14473);
and U15285 (N_15285,N_14074,N_14025);
nor U15286 (N_15286,N_14639,N_14354);
nand U15287 (N_15287,N_14816,N_14356);
nor U15288 (N_15288,N_14530,N_14981);
nor U15289 (N_15289,N_14449,N_14746);
xnor U15290 (N_15290,N_14366,N_14508);
xor U15291 (N_15291,N_14836,N_14910);
nand U15292 (N_15292,N_14687,N_14733);
nor U15293 (N_15293,N_14229,N_14425);
nand U15294 (N_15294,N_14576,N_14226);
xor U15295 (N_15295,N_14814,N_14930);
and U15296 (N_15296,N_14334,N_14396);
nand U15297 (N_15297,N_14708,N_14813);
or U15298 (N_15298,N_14936,N_14327);
and U15299 (N_15299,N_14093,N_14076);
or U15300 (N_15300,N_14036,N_14471);
xor U15301 (N_15301,N_14784,N_14666);
nand U15302 (N_15302,N_14020,N_14950);
and U15303 (N_15303,N_14113,N_14273);
and U15304 (N_15304,N_14318,N_14297);
or U15305 (N_15305,N_14765,N_14914);
and U15306 (N_15306,N_14392,N_14947);
nor U15307 (N_15307,N_14671,N_14253);
nor U15308 (N_15308,N_14223,N_14528);
nor U15309 (N_15309,N_14980,N_14560);
and U15310 (N_15310,N_14886,N_14448);
nor U15311 (N_15311,N_14299,N_14819);
nor U15312 (N_15312,N_14552,N_14599);
or U15313 (N_15313,N_14298,N_14744);
nand U15314 (N_15314,N_14224,N_14527);
nand U15315 (N_15315,N_14572,N_14621);
nand U15316 (N_15316,N_14963,N_14041);
or U15317 (N_15317,N_14055,N_14470);
and U15318 (N_15318,N_14404,N_14860);
nor U15319 (N_15319,N_14617,N_14243);
nor U15320 (N_15320,N_14598,N_14699);
nor U15321 (N_15321,N_14363,N_14329);
xor U15322 (N_15322,N_14060,N_14709);
or U15323 (N_15323,N_14755,N_14108);
and U15324 (N_15324,N_14301,N_14149);
nand U15325 (N_15325,N_14585,N_14918);
nand U15326 (N_15326,N_14372,N_14615);
xor U15327 (N_15327,N_14766,N_14976);
or U15328 (N_15328,N_14452,N_14325);
nand U15329 (N_15329,N_14264,N_14279);
and U15330 (N_15330,N_14833,N_14597);
xor U15331 (N_15331,N_14408,N_14481);
or U15332 (N_15332,N_14272,N_14233);
xor U15333 (N_15333,N_14543,N_14882);
nor U15334 (N_15334,N_14573,N_14252);
or U15335 (N_15335,N_14667,N_14374);
and U15336 (N_15336,N_14051,N_14966);
or U15337 (N_15337,N_14870,N_14219);
xnor U15338 (N_15338,N_14782,N_14477);
xnor U15339 (N_15339,N_14133,N_14926);
nor U15340 (N_15340,N_14420,N_14319);
xor U15341 (N_15341,N_14493,N_14569);
nand U15342 (N_15342,N_14673,N_14365);
nand U15343 (N_15343,N_14222,N_14580);
or U15344 (N_15344,N_14171,N_14691);
xnor U15345 (N_15345,N_14430,N_14958);
or U15346 (N_15346,N_14775,N_14344);
or U15347 (N_15347,N_14769,N_14236);
nor U15348 (N_15348,N_14453,N_14788);
nor U15349 (N_15349,N_14613,N_14577);
xnor U15350 (N_15350,N_14800,N_14502);
nand U15351 (N_15351,N_14561,N_14705);
xnor U15352 (N_15352,N_14102,N_14006);
xor U15353 (N_15353,N_14370,N_14174);
or U15354 (N_15354,N_14131,N_14303);
or U15355 (N_15355,N_14510,N_14064);
nand U15356 (N_15356,N_14793,N_14821);
and U15357 (N_15357,N_14859,N_14862);
nand U15358 (N_15358,N_14497,N_14367);
and U15359 (N_15359,N_14740,N_14281);
and U15360 (N_15360,N_14467,N_14676);
and U15361 (N_15361,N_14407,N_14762);
or U15362 (N_15362,N_14262,N_14719);
or U15363 (N_15363,N_14054,N_14828);
nor U15364 (N_15364,N_14044,N_14946);
and U15365 (N_15365,N_14053,N_14086);
nand U15366 (N_15366,N_14047,N_14317);
xnor U15367 (N_15367,N_14056,N_14302);
xnor U15368 (N_15368,N_14582,N_14934);
or U15369 (N_15369,N_14387,N_14331);
and U15370 (N_15370,N_14184,N_14686);
xor U15371 (N_15371,N_14403,N_14077);
and U15372 (N_15372,N_14111,N_14094);
or U15373 (N_15373,N_14352,N_14307);
xnor U15374 (N_15374,N_14275,N_14193);
or U15375 (N_15375,N_14050,N_14379);
and U15376 (N_15376,N_14166,N_14340);
or U15377 (N_15377,N_14484,N_14194);
nand U15378 (N_15378,N_14290,N_14796);
xnor U15379 (N_15379,N_14494,N_14721);
xor U15380 (N_15380,N_14888,N_14817);
xnor U15381 (N_15381,N_14984,N_14636);
nor U15382 (N_15382,N_14267,N_14758);
xor U15383 (N_15383,N_14805,N_14979);
or U15384 (N_15384,N_14583,N_14206);
nor U15385 (N_15385,N_14511,N_14207);
xnor U15386 (N_15386,N_14878,N_14199);
and U15387 (N_15387,N_14175,N_14698);
xnor U15388 (N_15388,N_14701,N_14043);
nor U15389 (N_15389,N_14336,N_14288);
nor U15390 (N_15390,N_14496,N_14178);
or U15391 (N_15391,N_14285,N_14853);
and U15392 (N_15392,N_14353,N_14927);
xor U15393 (N_15393,N_14286,N_14124);
nand U15394 (N_15394,N_14541,N_14851);
and U15395 (N_15395,N_14109,N_14778);
nand U15396 (N_15396,N_14773,N_14659);
nor U15397 (N_15397,N_14291,N_14724);
and U15398 (N_15398,N_14414,N_14832);
nor U15399 (N_15399,N_14132,N_14397);
nor U15400 (N_15400,N_14023,N_14218);
nand U15401 (N_15401,N_14916,N_14216);
and U15402 (N_15402,N_14030,N_14159);
nand U15403 (N_15403,N_14116,N_14098);
nand U15404 (N_15404,N_14120,N_14972);
or U15405 (N_15405,N_14516,N_14669);
or U15406 (N_15406,N_14747,N_14540);
nand U15407 (N_15407,N_14142,N_14277);
nor U15408 (N_15408,N_14685,N_14456);
xnor U15409 (N_15409,N_14941,N_14711);
and U15410 (N_15410,N_14898,N_14140);
xor U15411 (N_15411,N_14436,N_14842);
xor U15412 (N_15412,N_14695,N_14210);
nand U15413 (N_15413,N_14052,N_14220);
nand U15414 (N_15414,N_14150,N_14152);
nor U15415 (N_15415,N_14795,N_14463);
nand U15416 (N_15416,N_14412,N_14764);
and U15417 (N_15417,N_14742,N_14505);
xor U15418 (N_15418,N_14931,N_14749);
nand U15419 (N_15419,N_14694,N_14155);
xor U15420 (N_15420,N_14529,N_14189);
xnor U15421 (N_15421,N_14902,N_14920);
xor U15422 (N_15422,N_14809,N_14871);
nand U15423 (N_15423,N_14333,N_14300);
or U15424 (N_15424,N_14634,N_14850);
and U15425 (N_15425,N_14306,N_14015);
nor U15426 (N_15426,N_14567,N_14653);
xor U15427 (N_15427,N_14251,N_14935);
and U15428 (N_15428,N_14490,N_14127);
nand U15429 (N_15429,N_14703,N_14128);
nand U15430 (N_15430,N_14499,N_14338);
or U15431 (N_15431,N_14858,N_14643);
nand U15432 (N_15432,N_14413,N_14357);
xor U15433 (N_15433,N_14201,N_14040);
and U15434 (N_15434,N_14432,N_14107);
nand U15435 (N_15435,N_14549,N_14308);
xnor U15436 (N_15436,N_14388,N_14217);
nor U15437 (N_15437,N_14112,N_14364);
nand U15438 (N_15438,N_14311,N_14647);
xnor U15439 (N_15439,N_14147,N_14122);
nand U15440 (N_15440,N_14906,N_14894);
nand U15441 (N_15441,N_14165,N_14376);
xor U15442 (N_15442,N_14183,N_14534);
and U15443 (N_15443,N_14515,N_14244);
nor U15444 (N_15444,N_14962,N_14405);
nand U15445 (N_15445,N_14465,N_14390);
xnor U15446 (N_15446,N_14646,N_14774);
xnor U15447 (N_15447,N_14915,N_14191);
xnor U15448 (N_15448,N_14909,N_14974);
or U15449 (N_15449,N_14637,N_14482);
or U15450 (N_15450,N_14455,N_14466);
xnor U15451 (N_15451,N_14469,N_14488);
and U15452 (N_15452,N_14378,N_14579);
nor U15453 (N_15453,N_14801,N_14996);
or U15454 (N_15454,N_14787,N_14624);
xor U15455 (N_15455,N_14312,N_14864);
nand U15456 (N_15456,N_14973,N_14242);
or U15457 (N_15457,N_14616,N_14725);
xnor U15458 (N_15458,N_14657,N_14551);
and U15459 (N_15459,N_14704,N_14715);
nor U15460 (N_15460,N_14514,N_14638);
nor U15461 (N_15461,N_14739,N_14839);
xor U15462 (N_15462,N_14563,N_14863);
and U15463 (N_15463,N_14081,N_14230);
nand U15464 (N_15464,N_14153,N_14792);
xnor U15465 (N_15465,N_14925,N_14031);
nor U15466 (N_15466,N_14154,N_14478);
nor U15467 (N_15467,N_14874,N_14945);
nor U15468 (N_15468,N_14203,N_14501);
xnor U15469 (N_15469,N_14204,N_14531);
xnor U15470 (N_15470,N_14697,N_14610);
xnor U15471 (N_15471,N_14620,N_14134);
or U15472 (N_15472,N_14498,N_14012);
or U15473 (N_15473,N_14830,N_14732);
and U15474 (N_15474,N_14304,N_14283);
nor U15475 (N_15475,N_14360,N_14260);
and U15476 (N_15476,N_14852,N_14922);
or U15477 (N_15477,N_14532,N_14644);
nand U15478 (N_15478,N_14630,N_14879);
nor U15479 (N_15479,N_14714,N_14564);
xor U15480 (N_15480,N_14978,N_14235);
nor U15481 (N_15481,N_14339,N_14161);
and U15482 (N_15482,N_14967,N_14589);
or U15483 (N_15483,N_14424,N_14480);
xnor U15484 (N_15484,N_14038,N_14029);
nand U15485 (N_15485,N_14096,N_14202);
or U15486 (N_15486,N_14761,N_14883);
xnor U15487 (N_15487,N_14923,N_14547);
or U15488 (N_15488,N_14058,N_14525);
xor U15489 (N_15489,N_14377,N_14648);
xnor U15490 (N_15490,N_14042,N_14238);
or U15491 (N_15491,N_14261,N_14932);
xor U15492 (N_15492,N_14679,N_14752);
and U15493 (N_15493,N_14848,N_14856);
or U15494 (N_15494,N_14462,N_14003);
nor U15495 (N_15495,N_14917,N_14650);
nand U15496 (N_15496,N_14995,N_14662);
and U15497 (N_15497,N_14574,N_14689);
or U15498 (N_15498,N_14118,N_14522);
or U15499 (N_15499,N_14595,N_14717);
nor U15500 (N_15500,N_14504,N_14578);
xor U15501 (N_15501,N_14265,N_14212);
nand U15502 (N_15502,N_14409,N_14341);
xnor U15503 (N_15503,N_14982,N_14373);
or U15504 (N_15504,N_14418,N_14054);
nor U15505 (N_15505,N_14476,N_14738);
and U15506 (N_15506,N_14615,N_14972);
and U15507 (N_15507,N_14856,N_14656);
and U15508 (N_15508,N_14975,N_14994);
nor U15509 (N_15509,N_14122,N_14658);
or U15510 (N_15510,N_14472,N_14745);
xnor U15511 (N_15511,N_14143,N_14391);
and U15512 (N_15512,N_14510,N_14981);
xor U15513 (N_15513,N_14999,N_14391);
nand U15514 (N_15514,N_14848,N_14042);
nand U15515 (N_15515,N_14304,N_14831);
or U15516 (N_15516,N_14285,N_14716);
nor U15517 (N_15517,N_14123,N_14872);
or U15518 (N_15518,N_14344,N_14747);
and U15519 (N_15519,N_14551,N_14987);
nand U15520 (N_15520,N_14747,N_14212);
and U15521 (N_15521,N_14825,N_14154);
nand U15522 (N_15522,N_14758,N_14874);
xor U15523 (N_15523,N_14060,N_14929);
or U15524 (N_15524,N_14631,N_14237);
or U15525 (N_15525,N_14892,N_14840);
nor U15526 (N_15526,N_14861,N_14825);
and U15527 (N_15527,N_14466,N_14938);
xnor U15528 (N_15528,N_14119,N_14190);
or U15529 (N_15529,N_14329,N_14620);
and U15530 (N_15530,N_14048,N_14620);
and U15531 (N_15531,N_14271,N_14785);
nor U15532 (N_15532,N_14658,N_14368);
xnor U15533 (N_15533,N_14644,N_14413);
xor U15534 (N_15534,N_14793,N_14076);
xnor U15535 (N_15535,N_14251,N_14173);
or U15536 (N_15536,N_14024,N_14165);
xor U15537 (N_15537,N_14094,N_14785);
xor U15538 (N_15538,N_14562,N_14031);
xnor U15539 (N_15539,N_14224,N_14538);
or U15540 (N_15540,N_14333,N_14729);
or U15541 (N_15541,N_14852,N_14101);
and U15542 (N_15542,N_14652,N_14860);
xor U15543 (N_15543,N_14145,N_14942);
nand U15544 (N_15544,N_14592,N_14430);
nand U15545 (N_15545,N_14274,N_14886);
nor U15546 (N_15546,N_14394,N_14048);
nor U15547 (N_15547,N_14109,N_14118);
or U15548 (N_15548,N_14909,N_14146);
nand U15549 (N_15549,N_14928,N_14010);
nand U15550 (N_15550,N_14479,N_14781);
nand U15551 (N_15551,N_14077,N_14935);
nor U15552 (N_15552,N_14539,N_14062);
or U15553 (N_15553,N_14016,N_14816);
nand U15554 (N_15554,N_14548,N_14407);
nand U15555 (N_15555,N_14997,N_14732);
nor U15556 (N_15556,N_14049,N_14975);
and U15557 (N_15557,N_14516,N_14230);
and U15558 (N_15558,N_14276,N_14361);
and U15559 (N_15559,N_14769,N_14623);
xnor U15560 (N_15560,N_14415,N_14242);
or U15561 (N_15561,N_14352,N_14090);
and U15562 (N_15562,N_14507,N_14801);
and U15563 (N_15563,N_14317,N_14123);
nand U15564 (N_15564,N_14036,N_14055);
nand U15565 (N_15565,N_14744,N_14313);
and U15566 (N_15566,N_14097,N_14312);
nand U15567 (N_15567,N_14902,N_14425);
nand U15568 (N_15568,N_14159,N_14593);
or U15569 (N_15569,N_14901,N_14705);
or U15570 (N_15570,N_14515,N_14806);
and U15571 (N_15571,N_14049,N_14796);
nor U15572 (N_15572,N_14194,N_14660);
or U15573 (N_15573,N_14263,N_14773);
or U15574 (N_15574,N_14634,N_14651);
or U15575 (N_15575,N_14628,N_14242);
and U15576 (N_15576,N_14239,N_14773);
and U15577 (N_15577,N_14984,N_14388);
or U15578 (N_15578,N_14774,N_14819);
nand U15579 (N_15579,N_14555,N_14061);
nor U15580 (N_15580,N_14726,N_14233);
nor U15581 (N_15581,N_14171,N_14093);
and U15582 (N_15582,N_14890,N_14895);
nor U15583 (N_15583,N_14252,N_14468);
and U15584 (N_15584,N_14807,N_14008);
and U15585 (N_15585,N_14709,N_14176);
or U15586 (N_15586,N_14490,N_14010);
and U15587 (N_15587,N_14916,N_14814);
nand U15588 (N_15588,N_14532,N_14270);
nand U15589 (N_15589,N_14239,N_14420);
or U15590 (N_15590,N_14741,N_14883);
xnor U15591 (N_15591,N_14751,N_14796);
nor U15592 (N_15592,N_14054,N_14253);
and U15593 (N_15593,N_14547,N_14991);
xnor U15594 (N_15594,N_14259,N_14580);
nand U15595 (N_15595,N_14050,N_14553);
and U15596 (N_15596,N_14888,N_14362);
or U15597 (N_15597,N_14768,N_14014);
nand U15598 (N_15598,N_14232,N_14206);
or U15599 (N_15599,N_14287,N_14566);
nor U15600 (N_15600,N_14169,N_14488);
or U15601 (N_15601,N_14002,N_14114);
nand U15602 (N_15602,N_14141,N_14089);
or U15603 (N_15603,N_14196,N_14353);
nand U15604 (N_15604,N_14255,N_14402);
and U15605 (N_15605,N_14833,N_14116);
xnor U15606 (N_15606,N_14720,N_14648);
xnor U15607 (N_15607,N_14030,N_14967);
nor U15608 (N_15608,N_14953,N_14947);
or U15609 (N_15609,N_14801,N_14024);
nand U15610 (N_15610,N_14613,N_14678);
or U15611 (N_15611,N_14517,N_14160);
and U15612 (N_15612,N_14619,N_14287);
and U15613 (N_15613,N_14494,N_14700);
and U15614 (N_15614,N_14149,N_14117);
nor U15615 (N_15615,N_14964,N_14956);
and U15616 (N_15616,N_14124,N_14251);
and U15617 (N_15617,N_14719,N_14318);
nor U15618 (N_15618,N_14757,N_14460);
or U15619 (N_15619,N_14934,N_14512);
or U15620 (N_15620,N_14660,N_14502);
and U15621 (N_15621,N_14307,N_14904);
nor U15622 (N_15622,N_14599,N_14355);
nor U15623 (N_15623,N_14757,N_14777);
xor U15624 (N_15624,N_14165,N_14866);
or U15625 (N_15625,N_14544,N_14919);
xnor U15626 (N_15626,N_14266,N_14111);
nor U15627 (N_15627,N_14085,N_14756);
or U15628 (N_15628,N_14015,N_14706);
nor U15629 (N_15629,N_14948,N_14966);
or U15630 (N_15630,N_14446,N_14469);
nor U15631 (N_15631,N_14014,N_14884);
and U15632 (N_15632,N_14547,N_14043);
and U15633 (N_15633,N_14592,N_14694);
and U15634 (N_15634,N_14588,N_14878);
or U15635 (N_15635,N_14757,N_14373);
or U15636 (N_15636,N_14414,N_14165);
nand U15637 (N_15637,N_14097,N_14292);
or U15638 (N_15638,N_14158,N_14993);
nor U15639 (N_15639,N_14837,N_14273);
nor U15640 (N_15640,N_14421,N_14055);
or U15641 (N_15641,N_14919,N_14178);
and U15642 (N_15642,N_14235,N_14901);
xnor U15643 (N_15643,N_14414,N_14707);
nand U15644 (N_15644,N_14599,N_14394);
and U15645 (N_15645,N_14230,N_14335);
nor U15646 (N_15646,N_14993,N_14848);
or U15647 (N_15647,N_14442,N_14854);
or U15648 (N_15648,N_14421,N_14401);
or U15649 (N_15649,N_14367,N_14574);
nor U15650 (N_15650,N_14147,N_14697);
nor U15651 (N_15651,N_14422,N_14968);
xor U15652 (N_15652,N_14259,N_14710);
nor U15653 (N_15653,N_14853,N_14938);
nor U15654 (N_15654,N_14277,N_14689);
xor U15655 (N_15655,N_14281,N_14312);
and U15656 (N_15656,N_14790,N_14219);
nor U15657 (N_15657,N_14277,N_14788);
xor U15658 (N_15658,N_14124,N_14927);
xor U15659 (N_15659,N_14654,N_14081);
nor U15660 (N_15660,N_14588,N_14164);
or U15661 (N_15661,N_14521,N_14431);
or U15662 (N_15662,N_14425,N_14938);
or U15663 (N_15663,N_14173,N_14364);
nand U15664 (N_15664,N_14366,N_14858);
and U15665 (N_15665,N_14760,N_14749);
xnor U15666 (N_15666,N_14968,N_14251);
or U15667 (N_15667,N_14774,N_14270);
nand U15668 (N_15668,N_14509,N_14400);
and U15669 (N_15669,N_14402,N_14820);
or U15670 (N_15670,N_14537,N_14395);
and U15671 (N_15671,N_14562,N_14245);
or U15672 (N_15672,N_14219,N_14233);
or U15673 (N_15673,N_14402,N_14824);
and U15674 (N_15674,N_14387,N_14763);
xnor U15675 (N_15675,N_14717,N_14358);
nand U15676 (N_15676,N_14199,N_14909);
or U15677 (N_15677,N_14640,N_14454);
nor U15678 (N_15678,N_14236,N_14921);
nand U15679 (N_15679,N_14195,N_14465);
or U15680 (N_15680,N_14045,N_14653);
xor U15681 (N_15681,N_14623,N_14181);
or U15682 (N_15682,N_14427,N_14559);
nor U15683 (N_15683,N_14839,N_14644);
nand U15684 (N_15684,N_14698,N_14412);
or U15685 (N_15685,N_14668,N_14864);
nand U15686 (N_15686,N_14951,N_14775);
nor U15687 (N_15687,N_14142,N_14426);
nand U15688 (N_15688,N_14108,N_14611);
and U15689 (N_15689,N_14887,N_14893);
nor U15690 (N_15690,N_14750,N_14985);
xor U15691 (N_15691,N_14588,N_14209);
nor U15692 (N_15692,N_14017,N_14599);
nor U15693 (N_15693,N_14075,N_14891);
and U15694 (N_15694,N_14720,N_14853);
or U15695 (N_15695,N_14716,N_14300);
nor U15696 (N_15696,N_14891,N_14342);
nand U15697 (N_15697,N_14161,N_14599);
nor U15698 (N_15698,N_14056,N_14524);
or U15699 (N_15699,N_14714,N_14427);
or U15700 (N_15700,N_14844,N_14172);
xor U15701 (N_15701,N_14376,N_14194);
nand U15702 (N_15702,N_14508,N_14477);
xor U15703 (N_15703,N_14053,N_14885);
or U15704 (N_15704,N_14991,N_14246);
xor U15705 (N_15705,N_14695,N_14601);
nor U15706 (N_15706,N_14804,N_14157);
and U15707 (N_15707,N_14535,N_14144);
and U15708 (N_15708,N_14096,N_14616);
and U15709 (N_15709,N_14581,N_14556);
xnor U15710 (N_15710,N_14177,N_14951);
nand U15711 (N_15711,N_14052,N_14145);
or U15712 (N_15712,N_14757,N_14826);
nor U15713 (N_15713,N_14035,N_14538);
xnor U15714 (N_15714,N_14699,N_14357);
and U15715 (N_15715,N_14645,N_14253);
xor U15716 (N_15716,N_14618,N_14627);
or U15717 (N_15717,N_14815,N_14540);
xor U15718 (N_15718,N_14766,N_14686);
or U15719 (N_15719,N_14479,N_14256);
nand U15720 (N_15720,N_14866,N_14947);
nand U15721 (N_15721,N_14433,N_14931);
and U15722 (N_15722,N_14305,N_14616);
or U15723 (N_15723,N_14625,N_14600);
nor U15724 (N_15724,N_14109,N_14978);
nor U15725 (N_15725,N_14132,N_14430);
and U15726 (N_15726,N_14837,N_14864);
nand U15727 (N_15727,N_14383,N_14437);
nand U15728 (N_15728,N_14896,N_14219);
or U15729 (N_15729,N_14571,N_14130);
nor U15730 (N_15730,N_14525,N_14562);
or U15731 (N_15731,N_14621,N_14699);
and U15732 (N_15732,N_14297,N_14432);
xor U15733 (N_15733,N_14791,N_14437);
xnor U15734 (N_15734,N_14123,N_14353);
or U15735 (N_15735,N_14054,N_14674);
or U15736 (N_15736,N_14600,N_14475);
nand U15737 (N_15737,N_14215,N_14541);
xnor U15738 (N_15738,N_14529,N_14080);
nand U15739 (N_15739,N_14490,N_14399);
xnor U15740 (N_15740,N_14948,N_14439);
xnor U15741 (N_15741,N_14508,N_14700);
or U15742 (N_15742,N_14848,N_14509);
and U15743 (N_15743,N_14471,N_14799);
nand U15744 (N_15744,N_14802,N_14950);
and U15745 (N_15745,N_14799,N_14440);
nor U15746 (N_15746,N_14211,N_14632);
nor U15747 (N_15747,N_14235,N_14890);
nand U15748 (N_15748,N_14537,N_14785);
and U15749 (N_15749,N_14561,N_14173);
nand U15750 (N_15750,N_14094,N_14387);
and U15751 (N_15751,N_14369,N_14689);
and U15752 (N_15752,N_14182,N_14834);
or U15753 (N_15753,N_14045,N_14774);
or U15754 (N_15754,N_14382,N_14308);
and U15755 (N_15755,N_14486,N_14785);
xnor U15756 (N_15756,N_14487,N_14534);
or U15757 (N_15757,N_14835,N_14631);
nor U15758 (N_15758,N_14638,N_14843);
nor U15759 (N_15759,N_14158,N_14710);
xnor U15760 (N_15760,N_14445,N_14948);
nand U15761 (N_15761,N_14999,N_14990);
xnor U15762 (N_15762,N_14891,N_14271);
or U15763 (N_15763,N_14333,N_14179);
xnor U15764 (N_15764,N_14492,N_14011);
and U15765 (N_15765,N_14775,N_14592);
xnor U15766 (N_15766,N_14795,N_14207);
xnor U15767 (N_15767,N_14421,N_14381);
nand U15768 (N_15768,N_14495,N_14273);
and U15769 (N_15769,N_14614,N_14630);
or U15770 (N_15770,N_14966,N_14064);
or U15771 (N_15771,N_14173,N_14292);
or U15772 (N_15772,N_14891,N_14886);
nand U15773 (N_15773,N_14824,N_14949);
and U15774 (N_15774,N_14166,N_14514);
nor U15775 (N_15775,N_14689,N_14937);
xnor U15776 (N_15776,N_14228,N_14856);
and U15777 (N_15777,N_14925,N_14012);
nor U15778 (N_15778,N_14145,N_14629);
and U15779 (N_15779,N_14380,N_14267);
and U15780 (N_15780,N_14710,N_14910);
nor U15781 (N_15781,N_14435,N_14502);
or U15782 (N_15782,N_14945,N_14178);
nand U15783 (N_15783,N_14016,N_14199);
nand U15784 (N_15784,N_14135,N_14604);
or U15785 (N_15785,N_14315,N_14046);
xnor U15786 (N_15786,N_14178,N_14938);
nand U15787 (N_15787,N_14681,N_14998);
nor U15788 (N_15788,N_14540,N_14499);
xor U15789 (N_15789,N_14086,N_14585);
nand U15790 (N_15790,N_14914,N_14971);
or U15791 (N_15791,N_14243,N_14931);
nand U15792 (N_15792,N_14130,N_14119);
nor U15793 (N_15793,N_14140,N_14715);
xnor U15794 (N_15794,N_14741,N_14406);
and U15795 (N_15795,N_14864,N_14392);
and U15796 (N_15796,N_14371,N_14612);
nand U15797 (N_15797,N_14204,N_14896);
xor U15798 (N_15798,N_14177,N_14741);
nand U15799 (N_15799,N_14958,N_14280);
nand U15800 (N_15800,N_14222,N_14971);
nor U15801 (N_15801,N_14660,N_14128);
nor U15802 (N_15802,N_14413,N_14640);
or U15803 (N_15803,N_14108,N_14515);
nand U15804 (N_15804,N_14179,N_14089);
xnor U15805 (N_15805,N_14300,N_14048);
nand U15806 (N_15806,N_14173,N_14368);
nand U15807 (N_15807,N_14612,N_14361);
nor U15808 (N_15808,N_14675,N_14746);
nand U15809 (N_15809,N_14168,N_14707);
nand U15810 (N_15810,N_14855,N_14048);
nor U15811 (N_15811,N_14984,N_14924);
nand U15812 (N_15812,N_14974,N_14153);
nand U15813 (N_15813,N_14873,N_14980);
xor U15814 (N_15814,N_14435,N_14560);
nand U15815 (N_15815,N_14596,N_14224);
xor U15816 (N_15816,N_14848,N_14777);
or U15817 (N_15817,N_14516,N_14585);
and U15818 (N_15818,N_14734,N_14879);
nand U15819 (N_15819,N_14808,N_14012);
xor U15820 (N_15820,N_14275,N_14406);
nand U15821 (N_15821,N_14397,N_14079);
xor U15822 (N_15822,N_14735,N_14242);
nand U15823 (N_15823,N_14238,N_14310);
nand U15824 (N_15824,N_14075,N_14445);
or U15825 (N_15825,N_14799,N_14666);
nand U15826 (N_15826,N_14499,N_14447);
xor U15827 (N_15827,N_14206,N_14099);
and U15828 (N_15828,N_14757,N_14634);
nor U15829 (N_15829,N_14000,N_14824);
or U15830 (N_15830,N_14753,N_14344);
xor U15831 (N_15831,N_14726,N_14701);
and U15832 (N_15832,N_14521,N_14790);
xnor U15833 (N_15833,N_14806,N_14398);
and U15834 (N_15834,N_14334,N_14131);
xnor U15835 (N_15835,N_14575,N_14869);
nor U15836 (N_15836,N_14998,N_14567);
nand U15837 (N_15837,N_14093,N_14152);
nor U15838 (N_15838,N_14249,N_14854);
or U15839 (N_15839,N_14352,N_14033);
nor U15840 (N_15840,N_14645,N_14671);
and U15841 (N_15841,N_14130,N_14672);
nand U15842 (N_15842,N_14421,N_14914);
or U15843 (N_15843,N_14806,N_14130);
nor U15844 (N_15844,N_14083,N_14594);
or U15845 (N_15845,N_14341,N_14820);
nand U15846 (N_15846,N_14645,N_14797);
nor U15847 (N_15847,N_14796,N_14346);
xnor U15848 (N_15848,N_14311,N_14256);
or U15849 (N_15849,N_14173,N_14921);
or U15850 (N_15850,N_14068,N_14806);
nand U15851 (N_15851,N_14828,N_14508);
or U15852 (N_15852,N_14101,N_14287);
nor U15853 (N_15853,N_14000,N_14639);
nor U15854 (N_15854,N_14131,N_14415);
xnor U15855 (N_15855,N_14583,N_14859);
xor U15856 (N_15856,N_14636,N_14966);
or U15857 (N_15857,N_14326,N_14401);
xor U15858 (N_15858,N_14455,N_14023);
nand U15859 (N_15859,N_14023,N_14247);
or U15860 (N_15860,N_14509,N_14654);
xnor U15861 (N_15861,N_14463,N_14876);
and U15862 (N_15862,N_14006,N_14899);
nor U15863 (N_15863,N_14906,N_14408);
nand U15864 (N_15864,N_14978,N_14690);
nor U15865 (N_15865,N_14329,N_14755);
xnor U15866 (N_15866,N_14919,N_14800);
xor U15867 (N_15867,N_14212,N_14757);
nor U15868 (N_15868,N_14038,N_14310);
nand U15869 (N_15869,N_14097,N_14095);
or U15870 (N_15870,N_14747,N_14314);
and U15871 (N_15871,N_14450,N_14777);
and U15872 (N_15872,N_14982,N_14444);
and U15873 (N_15873,N_14456,N_14380);
or U15874 (N_15874,N_14346,N_14839);
and U15875 (N_15875,N_14511,N_14332);
or U15876 (N_15876,N_14580,N_14696);
and U15877 (N_15877,N_14622,N_14753);
or U15878 (N_15878,N_14125,N_14902);
xnor U15879 (N_15879,N_14829,N_14695);
nand U15880 (N_15880,N_14176,N_14880);
xor U15881 (N_15881,N_14528,N_14472);
nand U15882 (N_15882,N_14235,N_14467);
nand U15883 (N_15883,N_14794,N_14149);
xnor U15884 (N_15884,N_14335,N_14977);
xnor U15885 (N_15885,N_14214,N_14545);
xnor U15886 (N_15886,N_14633,N_14310);
nor U15887 (N_15887,N_14109,N_14061);
and U15888 (N_15888,N_14872,N_14779);
xnor U15889 (N_15889,N_14690,N_14694);
and U15890 (N_15890,N_14868,N_14414);
xnor U15891 (N_15891,N_14167,N_14021);
xor U15892 (N_15892,N_14780,N_14158);
xor U15893 (N_15893,N_14981,N_14163);
nand U15894 (N_15894,N_14934,N_14094);
and U15895 (N_15895,N_14392,N_14067);
or U15896 (N_15896,N_14168,N_14009);
nor U15897 (N_15897,N_14392,N_14910);
nand U15898 (N_15898,N_14891,N_14802);
or U15899 (N_15899,N_14345,N_14772);
xor U15900 (N_15900,N_14559,N_14346);
and U15901 (N_15901,N_14256,N_14769);
and U15902 (N_15902,N_14972,N_14436);
nor U15903 (N_15903,N_14911,N_14004);
xor U15904 (N_15904,N_14939,N_14742);
nand U15905 (N_15905,N_14461,N_14303);
nor U15906 (N_15906,N_14835,N_14672);
nand U15907 (N_15907,N_14218,N_14028);
nand U15908 (N_15908,N_14489,N_14634);
nand U15909 (N_15909,N_14477,N_14146);
xnor U15910 (N_15910,N_14886,N_14440);
nand U15911 (N_15911,N_14427,N_14020);
and U15912 (N_15912,N_14678,N_14267);
nand U15913 (N_15913,N_14321,N_14956);
and U15914 (N_15914,N_14445,N_14363);
nor U15915 (N_15915,N_14123,N_14431);
and U15916 (N_15916,N_14818,N_14977);
and U15917 (N_15917,N_14171,N_14970);
xor U15918 (N_15918,N_14142,N_14369);
and U15919 (N_15919,N_14705,N_14174);
nor U15920 (N_15920,N_14776,N_14752);
nand U15921 (N_15921,N_14146,N_14516);
nor U15922 (N_15922,N_14708,N_14375);
or U15923 (N_15923,N_14277,N_14136);
nor U15924 (N_15924,N_14090,N_14980);
nand U15925 (N_15925,N_14660,N_14066);
nand U15926 (N_15926,N_14537,N_14207);
nand U15927 (N_15927,N_14490,N_14864);
nor U15928 (N_15928,N_14945,N_14270);
xor U15929 (N_15929,N_14208,N_14093);
xnor U15930 (N_15930,N_14249,N_14168);
xnor U15931 (N_15931,N_14381,N_14542);
and U15932 (N_15932,N_14070,N_14395);
nor U15933 (N_15933,N_14024,N_14180);
and U15934 (N_15934,N_14952,N_14296);
nand U15935 (N_15935,N_14280,N_14638);
and U15936 (N_15936,N_14421,N_14311);
and U15937 (N_15937,N_14595,N_14648);
or U15938 (N_15938,N_14936,N_14415);
nor U15939 (N_15939,N_14091,N_14194);
xnor U15940 (N_15940,N_14500,N_14616);
xor U15941 (N_15941,N_14852,N_14988);
xnor U15942 (N_15942,N_14760,N_14214);
nor U15943 (N_15943,N_14086,N_14295);
nand U15944 (N_15944,N_14586,N_14326);
nand U15945 (N_15945,N_14425,N_14043);
xor U15946 (N_15946,N_14837,N_14959);
xnor U15947 (N_15947,N_14874,N_14746);
or U15948 (N_15948,N_14622,N_14233);
or U15949 (N_15949,N_14446,N_14300);
xor U15950 (N_15950,N_14689,N_14732);
or U15951 (N_15951,N_14115,N_14812);
nand U15952 (N_15952,N_14270,N_14915);
nand U15953 (N_15953,N_14203,N_14580);
nor U15954 (N_15954,N_14190,N_14854);
and U15955 (N_15955,N_14850,N_14937);
nand U15956 (N_15956,N_14392,N_14080);
nand U15957 (N_15957,N_14551,N_14704);
and U15958 (N_15958,N_14835,N_14374);
nor U15959 (N_15959,N_14301,N_14483);
xnor U15960 (N_15960,N_14610,N_14480);
and U15961 (N_15961,N_14654,N_14314);
nand U15962 (N_15962,N_14162,N_14654);
nor U15963 (N_15963,N_14640,N_14324);
nor U15964 (N_15964,N_14489,N_14274);
and U15965 (N_15965,N_14038,N_14457);
xnor U15966 (N_15966,N_14793,N_14653);
nor U15967 (N_15967,N_14064,N_14814);
nor U15968 (N_15968,N_14480,N_14165);
xnor U15969 (N_15969,N_14709,N_14724);
and U15970 (N_15970,N_14378,N_14112);
and U15971 (N_15971,N_14290,N_14538);
nand U15972 (N_15972,N_14037,N_14676);
and U15973 (N_15973,N_14735,N_14649);
xnor U15974 (N_15974,N_14173,N_14129);
xnor U15975 (N_15975,N_14998,N_14565);
or U15976 (N_15976,N_14494,N_14532);
nor U15977 (N_15977,N_14776,N_14791);
xor U15978 (N_15978,N_14048,N_14612);
or U15979 (N_15979,N_14778,N_14636);
xor U15980 (N_15980,N_14475,N_14495);
or U15981 (N_15981,N_14192,N_14026);
or U15982 (N_15982,N_14134,N_14817);
nor U15983 (N_15983,N_14140,N_14369);
xor U15984 (N_15984,N_14412,N_14771);
nor U15985 (N_15985,N_14427,N_14845);
nor U15986 (N_15986,N_14307,N_14552);
xor U15987 (N_15987,N_14804,N_14578);
or U15988 (N_15988,N_14163,N_14648);
and U15989 (N_15989,N_14063,N_14873);
nand U15990 (N_15990,N_14540,N_14704);
nor U15991 (N_15991,N_14876,N_14340);
or U15992 (N_15992,N_14792,N_14958);
xnor U15993 (N_15993,N_14583,N_14861);
nor U15994 (N_15994,N_14036,N_14790);
xor U15995 (N_15995,N_14861,N_14127);
or U15996 (N_15996,N_14936,N_14701);
nand U15997 (N_15997,N_14308,N_14032);
nand U15998 (N_15998,N_14528,N_14265);
nor U15999 (N_15999,N_14679,N_14120);
and U16000 (N_16000,N_15136,N_15693);
and U16001 (N_16001,N_15086,N_15676);
and U16002 (N_16002,N_15093,N_15096);
xnor U16003 (N_16003,N_15555,N_15483);
and U16004 (N_16004,N_15443,N_15370);
and U16005 (N_16005,N_15017,N_15120);
nor U16006 (N_16006,N_15384,N_15235);
and U16007 (N_16007,N_15129,N_15655);
nand U16008 (N_16008,N_15089,N_15471);
and U16009 (N_16009,N_15790,N_15466);
or U16010 (N_16010,N_15157,N_15703);
and U16011 (N_16011,N_15989,N_15691);
xnor U16012 (N_16012,N_15648,N_15361);
or U16013 (N_16013,N_15953,N_15885);
nor U16014 (N_16014,N_15763,N_15316);
or U16015 (N_16015,N_15686,N_15201);
nor U16016 (N_16016,N_15991,N_15331);
nand U16017 (N_16017,N_15163,N_15253);
or U16018 (N_16018,N_15199,N_15931);
or U16019 (N_16019,N_15977,N_15627);
nor U16020 (N_16020,N_15533,N_15787);
nor U16021 (N_16021,N_15146,N_15553);
and U16022 (N_16022,N_15234,N_15155);
nand U16023 (N_16023,N_15218,N_15418);
or U16024 (N_16024,N_15314,N_15293);
xor U16025 (N_16025,N_15079,N_15150);
nand U16026 (N_16026,N_15734,N_15057);
or U16027 (N_16027,N_15566,N_15924);
and U16028 (N_16028,N_15156,N_15240);
or U16029 (N_16029,N_15855,N_15695);
or U16030 (N_16030,N_15732,N_15356);
and U16031 (N_16031,N_15792,N_15375);
nor U16032 (N_16032,N_15069,N_15274);
and U16033 (N_16033,N_15256,N_15144);
or U16034 (N_16034,N_15397,N_15108);
xor U16035 (N_16035,N_15581,N_15700);
or U16036 (N_16036,N_15490,N_15765);
or U16037 (N_16037,N_15629,N_15460);
nand U16038 (N_16038,N_15962,N_15118);
nor U16039 (N_16039,N_15717,N_15399);
nand U16040 (N_16040,N_15639,N_15051);
nand U16041 (N_16041,N_15796,N_15066);
xnor U16042 (N_16042,N_15360,N_15635);
nand U16043 (N_16043,N_15744,N_15641);
xnor U16044 (N_16044,N_15650,N_15245);
and U16045 (N_16045,N_15509,N_15799);
or U16046 (N_16046,N_15898,N_15585);
nor U16047 (N_16047,N_15087,N_15236);
nand U16048 (N_16048,N_15781,N_15432);
and U16049 (N_16049,N_15248,N_15575);
nor U16050 (N_16050,N_15423,N_15965);
xor U16051 (N_16051,N_15659,N_15651);
or U16052 (N_16052,N_15012,N_15020);
nor U16053 (N_16053,N_15182,N_15172);
nor U16054 (N_16054,N_15847,N_15049);
or U16055 (N_16055,N_15554,N_15882);
nor U16056 (N_16056,N_15968,N_15672);
nand U16057 (N_16057,N_15865,N_15297);
and U16058 (N_16058,N_15834,N_15334);
nor U16059 (N_16059,N_15205,N_15436);
and U16060 (N_16060,N_15203,N_15495);
nand U16061 (N_16061,N_15442,N_15395);
nor U16062 (N_16062,N_15282,N_15197);
nand U16063 (N_16063,N_15178,N_15420);
nor U16064 (N_16064,N_15663,N_15671);
nand U16065 (N_16065,N_15474,N_15897);
xnor U16066 (N_16066,N_15188,N_15771);
and U16067 (N_16067,N_15391,N_15213);
xor U16068 (N_16068,N_15081,N_15615);
nor U16069 (N_16069,N_15307,N_15347);
or U16070 (N_16070,N_15278,N_15273);
nor U16071 (N_16071,N_15811,N_15603);
xnor U16072 (N_16072,N_15194,N_15401);
nor U16073 (N_16073,N_15883,N_15404);
and U16074 (N_16074,N_15364,N_15216);
and U16075 (N_16075,N_15955,N_15091);
nor U16076 (N_16076,N_15861,N_15382);
nor U16077 (N_16077,N_15767,N_15579);
nand U16078 (N_16078,N_15985,N_15995);
or U16079 (N_16079,N_15330,N_15284);
or U16080 (N_16080,N_15764,N_15301);
and U16081 (N_16081,N_15043,N_15348);
nand U16082 (N_16082,N_15183,N_15335);
and U16083 (N_16083,N_15266,N_15230);
nand U16084 (N_16084,N_15594,N_15611);
or U16085 (N_16085,N_15160,N_15685);
xor U16086 (N_16086,N_15353,N_15943);
or U16087 (N_16087,N_15488,N_15457);
and U16088 (N_16088,N_15626,N_15392);
or U16089 (N_16089,N_15130,N_15251);
or U16090 (N_16090,N_15678,N_15794);
nand U16091 (N_16091,N_15327,N_15545);
nor U16092 (N_16092,N_15954,N_15904);
or U16093 (N_16093,N_15591,N_15212);
xnor U16094 (N_16094,N_15867,N_15903);
or U16095 (N_16095,N_15009,N_15547);
or U16096 (N_16096,N_15682,N_15637);
nand U16097 (N_16097,N_15520,N_15596);
nand U16098 (N_16098,N_15192,N_15803);
or U16099 (N_16099,N_15106,N_15048);
xor U16100 (N_16100,N_15414,N_15708);
nor U16101 (N_16101,N_15735,N_15856);
nor U16102 (N_16102,N_15805,N_15938);
nor U16103 (N_16103,N_15500,N_15345);
and U16104 (N_16104,N_15149,N_15974);
nand U16105 (N_16105,N_15383,N_15768);
or U16106 (N_16106,N_15715,N_15281);
nor U16107 (N_16107,N_15934,N_15123);
or U16108 (N_16108,N_15970,N_15696);
xnor U16109 (N_16109,N_15342,N_15850);
nand U16110 (N_16110,N_15411,N_15412);
xor U16111 (N_16111,N_15625,N_15694);
xor U16112 (N_16112,N_15909,N_15452);
nand U16113 (N_16113,N_15426,N_15489);
nor U16114 (N_16114,N_15373,N_15941);
or U16115 (N_16115,N_15486,N_15134);
nor U16116 (N_16116,N_15802,N_15047);
or U16117 (N_16117,N_15170,N_15518);
or U16118 (N_16118,N_15262,N_15588);
xnor U16119 (N_16119,N_15413,N_15076);
nor U16120 (N_16120,N_15709,N_15932);
and U16121 (N_16121,N_15761,N_15719);
nand U16122 (N_16122,N_15535,N_15926);
nor U16123 (N_16123,N_15422,N_15832);
or U16124 (N_16124,N_15877,N_15595);
and U16125 (N_16125,N_15394,N_15675);
xnor U16126 (N_16126,N_15945,N_15598);
and U16127 (N_16127,N_15326,N_15058);
or U16128 (N_16128,N_15631,N_15731);
xnor U16129 (N_16129,N_15558,N_15055);
xnor U16130 (N_16130,N_15584,N_15922);
or U16131 (N_16131,N_15942,N_15793);
nand U16132 (N_16132,N_15578,N_15239);
nand U16133 (N_16133,N_15910,N_15433);
xnor U16134 (N_16134,N_15396,N_15747);
and U16135 (N_16135,N_15807,N_15369);
nand U16136 (N_16136,N_15393,N_15762);
or U16137 (N_16137,N_15892,N_15035);
nand U16138 (N_16138,N_15828,N_15366);
xnor U16139 (N_16139,N_15797,N_15153);
nand U16140 (N_16140,N_15127,N_15465);
and U16141 (N_16141,N_15435,N_15313);
or U16142 (N_16142,N_15439,N_15109);
or U16143 (N_16143,N_15121,N_15410);
and U16144 (N_16144,N_15008,N_15010);
xnor U16145 (N_16145,N_15280,N_15513);
and U16146 (N_16146,N_15895,N_15021);
and U16147 (N_16147,N_15998,N_15718);
xor U16148 (N_16148,N_15602,N_15871);
or U16149 (N_16149,N_15633,N_15227);
or U16150 (N_16150,N_15548,N_15788);
or U16151 (N_16151,N_15528,N_15774);
nor U16152 (N_16152,N_15561,N_15056);
or U16153 (N_16153,N_15687,N_15317);
xnor U16154 (N_16154,N_15532,N_15033);
or U16155 (N_16155,N_15878,N_15609);
or U16156 (N_16156,N_15791,N_15067);
nor U16157 (N_16157,N_15920,N_15223);
or U16158 (N_16158,N_15211,N_15884);
and U16159 (N_16159,N_15463,N_15484);
nand U16160 (N_16160,N_15947,N_15960);
nor U16161 (N_16161,N_15823,N_15138);
and U16162 (N_16162,N_15721,N_15472);
xnor U16163 (N_16163,N_15097,N_15501);
or U16164 (N_16164,N_15408,N_15099);
xnor U16165 (N_16165,N_15538,N_15844);
nand U16166 (N_16166,N_15210,N_15225);
nand U16167 (N_16167,N_15859,N_15980);
nor U16168 (N_16168,N_15377,N_15034);
xor U16169 (N_16169,N_15333,N_15986);
xor U16170 (N_16170,N_15740,N_15101);
or U16171 (N_16171,N_15214,N_15961);
nor U16172 (N_16172,N_15175,N_15996);
or U16173 (N_16173,N_15565,N_15652);
xor U16174 (N_16174,N_15956,N_15402);
xnor U16175 (N_16175,N_15729,N_15562);
nand U16176 (N_16176,N_15219,N_15543);
xor U16177 (N_16177,N_15690,N_15406);
and U16178 (N_16178,N_15125,N_15876);
xnor U16179 (N_16179,N_15372,N_15933);
nor U16180 (N_16180,N_15024,N_15312);
xnor U16181 (N_16181,N_15869,N_15870);
or U16182 (N_16182,N_15743,N_15654);
or U16183 (N_16183,N_15405,N_15050);
or U16184 (N_16184,N_15858,N_15344);
or U16185 (N_16185,N_15556,N_15517);
nand U16186 (N_16186,N_15665,N_15617);
or U16187 (N_16187,N_15380,N_15310);
xor U16188 (N_16188,N_15095,N_15450);
nor U16189 (N_16189,N_15110,N_15551);
xnor U16190 (N_16190,N_15424,N_15305);
nand U16191 (N_16191,N_15206,N_15576);
xnor U16192 (N_16192,N_15006,N_15683);
or U16193 (N_16193,N_15586,N_15905);
nor U16194 (N_16194,N_15630,N_15927);
xnor U16195 (N_16195,N_15889,N_15570);
and U16196 (N_16196,N_15505,N_15217);
nor U16197 (N_16197,N_15454,N_15818);
nor U16198 (N_16198,N_15226,N_15789);
nand U16199 (N_16199,N_15624,N_15819);
and U16200 (N_16200,N_15622,N_15409);
and U16201 (N_16201,N_15013,N_15571);
xnor U16202 (N_16202,N_15733,N_15320);
or U16203 (N_16203,N_15572,N_15267);
xor U16204 (N_16204,N_15040,N_15000);
xor U16205 (N_16205,N_15863,N_15666);
xor U16206 (N_16206,N_15599,N_15117);
nor U16207 (N_16207,N_15752,N_15264);
xnor U16208 (N_16208,N_15851,N_15906);
xnor U16209 (N_16209,N_15259,N_15119);
and U16210 (N_16210,N_15523,N_15604);
nand U16211 (N_16211,N_15018,N_15726);
or U16212 (N_16212,N_15946,N_15084);
nand U16213 (N_16213,N_15416,N_15514);
or U16214 (N_16214,N_15258,N_15775);
or U16215 (N_16215,N_15801,N_15315);
nor U16216 (N_16216,N_15400,N_15725);
xor U16217 (N_16217,N_15427,N_15949);
nor U16218 (N_16218,N_15357,N_15023);
and U16219 (N_16219,N_15482,N_15577);
nor U16220 (N_16220,N_15167,N_15560);
xor U16221 (N_16221,N_15044,N_15620);
nor U16222 (N_16222,N_15707,N_15967);
nor U16223 (N_16223,N_15243,N_15541);
xor U16224 (N_16224,N_15185,N_15673);
or U16225 (N_16225,N_15592,N_15772);
nor U16226 (N_16226,N_15147,N_15515);
xor U16227 (N_16227,N_15228,N_15512);
nor U16228 (N_16228,N_15171,N_15712);
nand U16229 (N_16229,N_15078,N_15169);
nand U16230 (N_16230,N_15837,N_15421);
xor U16231 (N_16231,N_15936,N_15536);
xnor U16232 (N_16232,N_15983,N_15723);
xnor U16233 (N_16233,N_15304,N_15068);
nor U16234 (N_16234,N_15866,N_15116);
nor U16235 (N_16235,N_15494,N_15921);
nand U16236 (N_16236,N_15030,N_15976);
xnor U16237 (N_16237,N_15191,N_15113);
or U16238 (N_16238,N_15115,N_15689);
xnor U16239 (N_16239,N_15038,N_15152);
or U16240 (N_16240,N_15887,N_15636);
nand U16241 (N_16241,N_15224,N_15958);
and U16242 (N_16242,N_15825,N_15151);
nor U16243 (N_16243,N_15914,N_15272);
or U16244 (N_16244,N_15827,N_15656);
nand U16245 (N_16245,N_15298,N_15658);
nor U16246 (N_16246,N_15491,N_15359);
or U16247 (N_16247,N_15254,N_15674);
and U16248 (N_16248,N_15742,N_15504);
and U16249 (N_16249,N_15842,N_15821);
nor U16250 (N_16250,N_15162,N_15498);
or U16251 (N_16251,N_15082,N_15343);
and U16252 (N_16252,N_15862,N_15229);
or U16253 (N_16253,N_15286,N_15193);
xor U16254 (N_16254,N_15516,N_15908);
nor U16255 (N_16255,N_15054,N_15727);
xor U16256 (N_16256,N_15090,N_15247);
xnor U16257 (N_16257,N_15785,N_15470);
nand U16258 (N_16258,N_15478,N_15759);
nor U16259 (N_16259,N_15061,N_15975);
and U16260 (N_16260,N_15506,N_15181);
and U16261 (N_16261,N_15311,N_15174);
xnor U16262 (N_16262,N_15525,N_15667);
nand U16263 (N_16263,N_15456,N_15710);
xor U16264 (N_16264,N_15756,N_15642);
nand U16265 (N_16265,N_15912,N_15843);
or U16266 (N_16266,N_15007,N_15065);
xnor U16267 (N_16267,N_15164,N_15275);
nand U16268 (N_16268,N_15649,N_15916);
and U16269 (N_16269,N_15306,N_15964);
xnor U16270 (N_16270,N_15559,N_15355);
nor U16271 (N_16271,N_15569,N_15778);
xnor U16272 (N_16272,N_15497,N_15668);
nand U16273 (N_16273,N_15769,N_15751);
or U16274 (N_16274,N_15632,N_15075);
and U16275 (N_16275,N_15749,N_15670);
or U16276 (N_16276,N_15145,N_15438);
xor U16277 (N_16277,N_15386,N_15993);
xnor U16278 (N_16278,N_15324,N_15398);
or U16279 (N_16279,N_15817,N_15755);
nor U16280 (N_16280,N_15813,N_15621);
and U16281 (N_16281,N_15950,N_15510);
xor U16282 (N_16282,N_15814,N_15131);
nand U16283 (N_16283,N_15852,N_15786);
nand U16284 (N_16284,N_15529,N_15815);
or U16285 (N_16285,N_15276,N_15329);
xor U16286 (N_16286,N_15100,N_15221);
and U16287 (N_16287,N_15022,N_15165);
or U16288 (N_16288,N_15952,N_15784);
xor U16289 (N_16289,N_15526,N_15738);
and U16290 (N_16290,N_15522,N_15657);
nor U16291 (N_16291,N_15564,N_15836);
or U16292 (N_16292,N_15647,N_15200);
and U16293 (N_16293,N_15754,N_15841);
nand U16294 (N_16294,N_15042,N_15350);
nand U16295 (N_16295,N_15015,N_15773);
or U16296 (N_16296,N_15287,N_15208);
nand U16297 (N_16297,N_15702,N_15730);
and U16298 (N_16298,N_15161,N_15291);
or U16299 (N_16299,N_15362,N_15063);
xor U16300 (N_16300,N_15469,N_15025);
or U16301 (N_16301,N_15846,N_15168);
nor U16302 (N_16302,N_15770,N_15748);
nand U16303 (N_16303,N_15209,N_15242);
or U16304 (N_16304,N_15653,N_15679);
nand U16305 (N_16305,N_15459,N_15688);
nor U16306 (N_16306,N_15376,N_15233);
xnor U16307 (N_16307,N_15587,N_15447);
and U16308 (N_16308,N_15368,N_15045);
and U16309 (N_16309,N_15464,N_15779);
nor U16310 (N_16310,N_15473,N_15872);
and U16311 (N_16311,N_15261,N_15441);
nor U16312 (N_16312,N_15750,N_15309);
and U16313 (N_16313,N_15886,N_15940);
or U16314 (N_16314,N_15704,N_15824);
or U16315 (N_16315,N_15299,N_15777);
nand U16316 (N_16316,N_15429,N_15902);
xor U16317 (N_16317,N_15939,N_15070);
nand U16318 (N_16318,N_15705,N_15831);
or U16319 (N_16319,N_15337,N_15270);
or U16320 (N_16320,N_15133,N_15745);
and U16321 (N_16321,N_15431,N_15616);
and U16322 (N_16322,N_15001,N_15137);
xor U16323 (N_16323,N_15978,N_15568);
nor U16324 (N_16324,N_15177,N_15351);
nor U16325 (N_16325,N_15646,N_15294);
xor U16326 (N_16326,N_15080,N_15487);
xnor U16327 (N_16327,N_15308,N_15741);
xor U16328 (N_16328,N_15323,N_15660);
and U16329 (N_16329,N_15289,N_15971);
or U16330 (N_16330,N_15026,N_15783);
nor U16331 (N_16331,N_15249,N_15184);
or U16332 (N_16332,N_15567,N_15011);
nand U16333 (N_16333,N_15524,N_15806);
and U16334 (N_16334,N_15812,N_15159);
nor U16335 (N_16335,N_15349,N_15428);
nand U16336 (N_16336,N_15060,N_15135);
or U16337 (N_16337,N_15031,N_15283);
and U16338 (N_16338,N_15461,N_15645);
xor U16339 (N_16339,N_15141,N_15430);
nor U16340 (N_16340,N_15816,N_15389);
and U16341 (N_16341,N_15002,N_15677);
nand U16342 (N_16342,N_15445,N_15605);
nand U16343 (N_16343,N_15890,N_15232);
nand U16344 (N_16344,N_15111,N_15074);
xor U16345 (N_16345,N_15881,N_15848);
nor U16346 (N_16346,N_15893,N_15328);
xnor U16347 (N_16347,N_15105,N_15325);
nand U16348 (N_16348,N_15455,N_15901);
or U16349 (N_16349,N_15029,N_15614);
or U16350 (N_16350,N_15387,N_15005);
and U16351 (N_16351,N_15189,N_15367);
nor U16352 (N_16352,N_15680,N_15303);
xor U16353 (N_16353,N_15590,N_15059);
or U16354 (N_16354,N_15440,N_15255);
nor U16355 (N_16355,N_15053,N_15537);
nand U16356 (N_16356,N_15891,N_15332);
nor U16357 (N_16357,N_15077,N_15736);
and U16358 (N_16358,N_15610,N_15716);
or U16359 (N_16359,N_15046,N_15019);
or U16360 (N_16360,N_15458,N_15969);
nand U16361 (N_16361,N_15062,N_15508);
xor U16362 (N_16362,N_15507,N_15477);
and U16363 (N_16363,N_15929,N_15589);
and U16364 (N_16364,N_15994,N_15981);
nor U16365 (N_16365,N_15546,N_15425);
xor U16366 (N_16366,N_15640,N_15363);
nand U16367 (N_16367,N_15701,N_15016);
nor U16368 (N_16368,N_15835,N_15318);
or U16369 (N_16369,N_15935,N_15527);
nand U16370 (N_16370,N_15925,N_15148);
nand U16371 (N_16371,N_15988,N_15444);
nand U16372 (N_16372,N_15187,N_15003);
or U16373 (N_16373,N_15032,N_15951);
or U16374 (N_16374,N_15502,N_15853);
xnor U16375 (N_16375,N_15112,N_15453);
xor U16376 (N_16376,N_15780,N_15550);
or U16377 (N_16377,N_15319,N_15607);
nand U16378 (N_16378,N_15338,N_15923);
nor U16379 (N_16379,N_15661,N_15593);
xnor U16380 (N_16380,N_15014,N_15468);
or U16381 (N_16381,N_15492,N_15462);
xor U16382 (N_16382,N_15911,N_15388);
and U16383 (N_16383,N_15757,N_15521);
and U16384 (N_16384,N_15039,N_15041);
and U16385 (N_16385,N_15238,N_15760);
nor U16386 (N_16386,N_15302,N_15158);
nand U16387 (N_16387,N_15446,N_15896);
xnor U16388 (N_16388,N_15176,N_15959);
and U16389 (N_16389,N_15295,N_15713);
nand U16390 (N_16390,N_15580,N_15340);
nand U16391 (N_16391,N_15917,N_15600);
nor U16392 (N_16392,N_15840,N_15531);
nor U16393 (N_16393,N_15601,N_15260);
nand U16394 (N_16394,N_15997,N_15698);
or U16395 (N_16395,N_15122,N_15612);
nand U16396 (N_16396,N_15140,N_15503);
nor U16397 (N_16397,N_15374,N_15296);
and U16398 (N_16398,N_15573,N_15083);
or U16399 (N_16399,N_15246,N_15776);
and U16400 (N_16400,N_15519,N_15880);
and U16401 (N_16401,N_15403,N_15966);
nand U16402 (N_16402,N_15269,N_15544);
nand U16403 (N_16403,N_15037,N_15879);
nand U16404 (N_16404,N_15845,N_15196);
and U16405 (N_16405,N_15142,N_15692);
and U16406 (N_16406,N_15004,N_15982);
xnor U16407 (N_16407,N_15822,N_15919);
or U16408 (N_16408,N_15800,N_15915);
nor U16409 (N_16409,N_15534,N_15720);
and U16410 (N_16410,N_15265,N_15407);
and U16411 (N_16411,N_15583,N_15451);
xnor U16412 (N_16412,N_15999,N_15085);
or U16413 (N_16413,N_15984,N_15207);
nor U16414 (N_16414,N_15180,N_15699);
nor U16415 (N_16415,N_15102,N_15341);
xor U16416 (N_16416,N_15114,N_15288);
nand U16417 (N_16417,N_15027,N_15336);
nor U16418 (N_16418,N_15766,N_15092);
xnor U16419 (N_16419,N_15390,N_15972);
or U16420 (N_16420,N_15231,N_15098);
nand U16421 (N_16421,N_15449,N_15417);
xor U16422 (N_16422,N_15838,N_15354);
or U16423 (N_16423,N_15711,N_15606);
and U16424 (N_16424,N_15241,N_15937);
and U16425 (N_16425,N_15480,N_15643);
and U16426 (N_16426,N_15634,N_15662);
and U16427 (N_16427,N_15139,N_15052);
or U16428 (N_16428,N_15104,N_15479);
nor U16429 (N_16429,N_15888,N_15552);
nand U16430 (N_16430,N_15979,N_15352);
xor U16431 (N_16431,N_15758,N_15874);
nand U16432 (N_16432,N_15198,N_15244);
and U16433 (N_16433,N_15684,N_15987);
nor U16434 (N_16434,N_15644,N_15036);
and U16435 (N_16435,N_15722,N_15252);
xnor U16436 (N_16436,N_15574,N_15072);
xnor U16437 (N_16437,N_15992,N_15419);
nor U16438 (N_16438,N_15485,N_15434);
nand U16439 (N_16439,N_15664,N_15475);
nor U16440 (N_16440,N_15300,N_15839);
or U16441 (N_16441,N_15530,N_15381);
and U16442 (N_16442,N_15809,N_15154);
and U16443 (N_16443,N_15539,N_15582);
or U16444 (N_16444,N_15944,N_15804);
and U16445 (N_16445,N_15810,N_15875);
xor U16446 (N_16446,N_15202,N_15204);
and U16447 (N_16447,N_15365,N_15143);
nand U16448 (N_16448,N_15173,N_15918);
nand U16449 (N_16449,N_15496,N_15913);
and U16450 (N_16450,N_15250,N_15271);
nand U16451 (N_16451,N_15619,N_15071);
and U16452 (N_16452,N_15179,N_15706);
or U16453 (N_16453,N_15563,N_15963);
nand U16454 (N_16454,N_15860,N_15928);
or U16455 (N_16455,N_15795,N_15290);
nor U16456 (N_16456,N_15714,N_15215);
and U16457 (N_16457,N_15618,N_15467);
xor U16458 (N_16458,N_15739,N_15830);
nor U16459 (N_16459,N_15753,N_15222);
or U16460 (N_16460,N_15476,N_15557);
nand U16461 (N_16461,N_15826,N_15511);
nand U16462 (N_16462,N_15868,N_15064);
xor U16463 (N_16463,N_15820,N_15873);
xor U16464 (N_16464,N_15379,N_15864);
xnor U16465 (N_16465,N_15542,N_15107);
nand U16466 (N_16466,N_15857,N_15907);
xnor U16467 (N_16467,N_15292,N_15237);
nand U16468 (N_16468,N_15094,N_15894);
and U16469 (N_16469,N_15371,N_15124);
xnor U16470 (N_16470,N_15128,N_15930);
and U16471 (N_16471,N_15854,N_15638);
and U16472 (N_16472,N_15481,N_15195);
nor U16473 (N_16473,N_15415,N_15268);
nor U16474 (N_16474,N_15321,N_15669);
nand U16475 (N_16475,N_15746,N_15737);
xnor U16476 (N_16476,N_15437,N_15166);
nor U16477 (N_16477,N_15900,N_15549);
nand U16478 (N_16478,N_15493,N_15499);
nand U16479 (N_16479,N_15613,N_15279);
xnor U16480 (N_16480,N_15681,N_15028);
nor U16481 (N_16481,N_15833,N_15190);
nand U16482 (N_16482,N_15948,N_15126);
nor U16483 (N_16483,N_15346,N_15540);
nor U16484 (N_16484,N_15378,N_15322);
xnor U16485 (N_16485,N_15728,N_15285);
nand U16486 (N_16486,N_15385,N_15798);
or U16487 (N_16487,N_15448,N_15257);
or U16488 (N_16488,N_15829,N_15849);
and U16489 (N_16489,N_15623,N_15277);
nand U16490 (N_16490,N_15103,N_15088);
and U16491 (N_16491,N_15339,N_15990);
nand U16492 (N_16492,N_15782,N_15724);
nor U16493 (N_16493,N_15957,N_15186);
nor U16494 (N_16494,N_15132,N_15220);
nand U16495 (N_16495,N_15899,N_15608);
and U16496 (N_16496,N_15973,N_15697);
and U16497 (N_16497,N_15808,N_15073);
and U16498 (N_16498,N_15597,N_15263);
nor U16499 (N_16499,N_15358,N_15628);
nand U16500 (N_16500,N_15106,N_15213);
or U16501 (N_16501,N_15860,N_15981);
nor U16502 (N_16502,N_15103,N_15365);
xnor U16503 (N_16503,N_15361,N_15008);
xnor U16504 (N_16504,N_15423,N_15588);
xor U16505 (N_16505,N_15126,N_15283);
or U16506 (N_16506,N_15750,N_15133);
or U16507 (N_16507,N_15922,N_15340);
and U16508 (N_16508,N_15222,N_15389);
or U16509 (N_16509,N_15020,N_15876);
xor U16510 (N_16510,N_15092,N_15972);
xor U16511 (N_16511,N_15221,N_15550);
nand U16512 (N_16512,N_15384,N_15289);
nand U16513 (N_16513,N_15556,N_15982);
xnor U16514 (N_16514,N_15439,N_15080);
xnor U16515 (N_16515,N_15748,N_15428);
nand U16516 (N_16516,N_15232,N_15780);
and U16517 (N_16517,N_15489,N_15669);
and U16518 (N_16518,N_15057,N_15472);
and U16519 (N_16519,N_15927,N_15884);
or U16520 (N_16520,N_15251,N_15171);
and U16521 (N_16521,N_15661,N_15084);
nand U16522 (N_16522,N_15100,N_15138);
nor U16523 (N_16523,N_15895,N_15608);
nand U16524 (N_16524,N_15549,N_15361);
and U16525 (N_16525,N_15696,N_15026);
nand U16526 (N_16526,N_15002,N_15653);
nand U16527 (N_16527,N_15546,N_15378);
nor U16528 (N_16528,N_15920,N_15918);
nand U16529 (N_16529,N_15410,N_15915);
nand U16530 (N_16530,N_15088,N_15535);
nand U16531 (N_16531,N_15253,N_15965);
and U16532 (N_16532,N_15502,N_15885);
or U16533 (N_16533,N_15820,N_15035);
and U16534 (N_16534,N_15099,N_15384);
nand U16535 (N_16535,N_15432,N_15900);
nor U16536 (N_16536,N_15358,N_15079);
or U16537 (N_16537,N_15214,N_15011);
or U16538 (N_16538,N_15716,N_15224);
nor U16539 (N_16539,N_15936,N_15047);
nor U16540 (N_16540,N_15078,N_15339);
nor U16541 (N_16541,N_15386,N_15377);
nand U16542 (N_16542,N_15759,N_15040);
nor U16543 (N_16543,N_15808,N_15466);
nor U16544 (N_16544,N_15663,N_15015);
xor U16545 (N_16545,N_15498,N_15494);
nand U16546 (N_16546,N_15986,N_15506);
nor U16547 (N_16547,N_15132,N_15026);
nand U16548 (N_16548,N_15680,N_15192);
nand U16549 (N_16549,N_15448,N_15805);
and U16550 (N_16550,N_15847,N_15066);
nand U16551 (N_16551,N_15813,N_15346);
nor U16552 (N_16552,N_15029,N_15974);
xnor U16553 (N_16553,N_15088,N_15250);
nand U16554 (N_16554,N_15548,N_15491);
and U16555 (N_16555,N_15409,N_15752);
or U16556 (N_16556,N_15842,N_15633);
nor U16557 (N_16557,N_15076,N_15362);
nor U16558 (N_16558,N_15669,N_15054);
nor U16559 (N_16559,N_15589,N_15551);
xnor U16560 (N_16560,N_15022,N_15144);
nand U16561 (N_16561,N_15057,N_15149);
xor U16562 (N_16562,N_15241,N_15986);
xor U16563 (N_16563,N_15659,N_15235);
nor U16564 (N_16564,N_15746,N_15609);
xnor U16565 (N_16565,N_15196,N_15949);
xor U16566 (N_16566,N_15491,N_15345);
or U16567 (N_16567,N_15047,N_15649);
nand U16568 (N_16568,N_15810,N_15488);
nor U16569 (N_16569,N_15440,N_15278);
and U16570 (N_16570,N_15342,N_15921);
nor U16571 (N_16571,N_15038,N_15022);
and U16572 (N_16572,N_15028,N_15286);
and U16573 (N_16573,N_15999,N_15458);
nand U16574 (N_16574,N_15602,N_15725);
nand U16575 (N_16575,N_15077,N_15504);
xor U16576 (N_16576,N_15198,N_15504);
and U16577 (N_16577,N_15231,N_15423);
nand U16578 (N_16578,N_15829,N_15480);
and U16579 (N_16579,N_15570,N_15472);
and U16580 (N_16580,N_15782,N_15558);
or U16581 (N_16581,N_15353,N_15524);
nor U16582 (N_16582,N_15607,N_15993);
nor U16583 (N_16583,N_15756,N_15829);
and U16584 (N_16584,N_15601,N_15558);
xnor U16585 (N_16585,N_15333,N_15713);
nor U16586 (N_16586,N_15833,N_15660);
xnor U16587 (N_16587,N_15108,N_15226);
or U16588 (N_16588,N_15793,N_15003);
or U16589 (N_16589,N_15585,N_15149);
xor U16590 (N_16590,N_15729,N_15561);
nand U16591 (N_16591,N_15179,N_15076);
or U16592 (N_16592,N_15276,N_15107);
and U16593 (N_16593,N_15974,N_15617);
xor U16594 (N_16594,N_15616,N_15079);
or U16595 (N_16595,N_15657,N_15474);
xnor U16596 (N_16596,N_15452,N_15562);
or U16597 (N_16597,N_15311,N_15270);
xnor U16598 (N_16598,N_15026,N_15907);
nor U16599 (N_16599,N_15305,N_15861);
nor U16600 (N_16600,N_15121,N_15343);
xnor U16601 (N_16601,N_15521,N_15085);
nand U16602 (N_16602,N_15018,N_15516);
nand U16603 (N_16603,N_15759,N_15835);
nand U16604 (N_16604,N_15315,N_15378);
or U16605 (N_16605,N_15079,N_15100);
xor U16606 (N_16606,N_15495,N_15885);
nand U16607 (N_16607,N_15999,N_15058);
nor U16608 (N_16608,N_15701,N_15083);
and U16609 (N_16609,N_15017,N_15022);
xnor U16610 (N_16610,N_15572,N_15037);
or U16611 (N_16611,N_15151,N_15535);
nor U16612 (N_16612,N_15816,N_15697);
nand U16613 (N_16613,N_15522,N_15242);
nand U16614 (N_16614,N_15440,N_15573);
nand U16615 (N_16615,N_15079,N_15507);
or U16616 (N_16616,N_15341,N_15733);
nand U16617 (N_16617,N_15759,N_15765);
nand U16618 (N_16618,N_15189,N_15529);
nor U16619 (N_16619,N_15123,N_15268);
or U16620 (N_16620,N_15628,N_15847);
or U16621 (N_16621,N_15687,N_15522);
xnor U16622 (N_16622,N_15246,N_15089);
nand U16623 (N_16623,N_15874,N_15441);
nand U16624 (N_16624,N_15999,N_15690);
xnor U16625 (N_16625,N_15762,N_15149);
or U16626 (N_16626,N_15158,N_15084);
xor U16627 (N_16627,N_15025,N_15131);
or U16628 (N_16628,N_15411,N_15020);
nor U16629 (N_16629,N_15786,N_15067);
and U16630 (N_16630,N_15732,N_15902);
or U16631 (N_16631,N_15696,N_15705);
or U16632 (N_16632,N_15197,N_15917);
or U16633 (N_16633,N_15907,N_15143);
nor U16634 (N_16634,N_15739,N_15984);
xnor U16635 (N_16635,N_15403,N_15640);
nand U16636 (N_16636,N_15757,N_15417);
or U16637 (N_16637,N_15308,N_15850);
and U16638 (N_16638,N_15993,N_15267);
nand U16639 (N_16639,N_15057,N_15844);
nor U16640 (N_16640,N_15799,N_15658);
or U16641 (N_16641,N_15050,N_15756);
xnor U16642 (N_16642,N_15932,N_15727);
nor U16643 (N_16643,N_15333,N_15887);
nor U16644 (N_16644,N_15140,N_15252);
xnor U16645 (N_16645,N_15921,N_15197);
nor U16646 (N_16646,N_15588,N_15094);
or U16647 (N_16647,N_15092,N_15858);
nand U16648 (N_16648,N_15713,N_15140);
xor U16649 (N_16649,N_15131,N_15822);
nand U16650 (N_16650,N_15781,N_15202);
nand U16651 (N_16651,N_15717,N_15237);
and U16652 (N_16652,N_15827,N_15350);
or U16653 (N_16653,N_15323,N_15034);
nor U16654 (N_16654,N_15839,N_15819);
nor U16655 (N_16655,N_15110,N_15707);
nor U16656 (N_16656,N_15092,N_15015);
xor U16657 (N_16657,N_15993,N_15206);
or U16658 (N_16658,N_15162,N_15985);
nor U16659 (N_16659,N_15827,N_15387);
nor U16660 (N_16660,N_15592,N_15797);
nand U16661 (N_16661,N_15120,N_15649);
or U16662 (N_16662,N_15938,N_15976);
nand U16663 (N_16663,N_15803,N_15616);
nor U16664 (N_16664,N_15650,N_15070);
nand U16665 (N_16665,N_15975,N_15292);
or U16666 (N_16666,N_15658,N_15772);
and U16667 (N_16667,N_15671,N_15106);
and U16668 (N_16668,N_15561,N_15800);
xor U16669 (N_16669,N_15822,N_15500);
nand U16670 (N_16670,N_15368,N_15878);
nor U16671 (N_16671,N_15767,N_15707);
nor U16672 (N_16672,N_15645,N_15887);
or U16673 (N_16673,N_15144,N_15740);
or U16674 (N_16674,N_15638,N_15883);
and U16675 (N_16675,N_15832,N_15402);
nand U16676 (N_16676,N_15194,N_15698);
nand U16677 (N_16677,N_15973,N_15710);
or U16678 (N_16678,N_15261,N_15329);
and U16679 (N_16679,N_15231,N_15180);
and U16680 (N_16680,N_15956,N_15620);
and U16681 (N_16681,N_15034,N_15841);
xnor U16682 (N_16682,N_15487,N_15469);
nor U16683 (N_16683,N_15513,N_15845);
nor U16684 (N_16684,N_15353,N_15504);
or U16685 (N_16685,N_15825,N_15806);
nor U16686 (N_16686,N_15128,N_15038);
and U16687 (N_16687,N_15170,N_15021);
and U16688 (N_16688,N_15970,N_15097);
nand U16689 (N_16689,N_15362,N_15991);
xnor U16690 (N_16690,N_15768,N_15916);
or U16691 (N_16691,N_15322,N_15419);
or U16692 (N_16692,N_15329,N_15053);
xor U16693 (N_16693,N_15539,N_15566);
nand U16694 (N_16694,N_15214,N_15889);
xnor U16695 (N_16695,N_15350,N_15097);
and U16696 (N_16696,N_15936,N_15588);
nor U16697 (N_16697,N_15042,N_15705);
nand U16698 (N_16698,N_15219,N_15991);
or U16699 (N_16699,N_15373,N_15030);
xnor U16700 (N_16700,N_15832,N_15972);
nor U16701 (N_16701,N_15871,N_15734);
nor U16702 (N_16702,N_15707,N_15375);
and U16703 (N_16703,N_15856,N_15073);
and U16704 (N_16704,N_15036,N_15112);
or U16705 (N_16705,N_15343,N_15375);
nand U16706 (N_16706,N_15686,N_15790);
nand U16707 (N_16707,N_15378,N_15556);
nor U16708 (N_16708,N_15403,N_15131);
nor U16709 (N_16709,N_15514,N_15132);
nor U16710 (N_16710,N_15045,N_15223);
xor U16711 (N_16711,N_15359,N_15549);
nand U16712 (N_16712,N_15650,N_15951);
xor U16713 (N_16713,N_15759,N_15826);
nand U16714 (N_16714,N_15183,N_15239);
or U16715 (N_16715,N_15138,N_15935);
nor U16716 (N_16716,N_15312,N_15448);
nor U16717 (N_16717,N_15859,N_15662);
xnor U16718 (N_16718,N_15478,N_15550);
xnor U16719 (N_16719,N_15758,N_15614);
or U16720 (N_16720,N_15727,N_15019);
xor U16721 (N_16721,N_15040,N_15154);
or U16722 (N_16722,N_15329,N_15669);
and U16723 (N_16723,N_15952,N_15164);
nand U16724 (N_16724,N_15519,N_15667);
nand U16725 (N_16725,N_15571,N_15476);
or U16726 (N_16726,N_15664,N_15793);
xnor U16727 (N_16727,N_15068,N_15282);
nand U16728 (N_16728,N_15464,N_15201);
nor U16729 (N_16729,N_15069,N_15337);
nand U16730 (N_16730,N_15069,N_15677);
nand U16731 (N_16731,N_15331,N_15056);
nand U16732 (N_16732,N_15065,N_15232);
nand U16733 (N_16733,N_15074,N_15143);
nor U16734 (N_16734,N_15459,N_15245);
and U16735 (N_16735,N_15526,N_15321);
xnor U16736 (N_16736,N_15313,N_15683);
xnor U16737 (N_16737,N_15687,N_15911);
nand U16738 (N_16738,N_15409,N_15988);
nand U16739 (N_16739,N_15241,N_15187);
nor U16740 (N_16740,N_15330,N_15063);
nor U16741 (N_16741,N_15845,N_15987);
or U16742 (N_16742,N_15605,N_15457);
nor U16743 (N_16743,N_15379,N_15415);
or U16744 (N_16744,N_15197,N_15819);
nand U16745 (N_16745,N_15018,N_15827);
and U16746 (N_16746,N_15277,N_15648);
nand U16747 (N_16747,N_15712,N_15668);
nand U16748 (N_16748,N_15982,N_15035);
or U16749 (N_16749,N_15811,N_15453);
or U16750 (N_16750,N_15368,N_15980);
or U16751 (N_16751,N_15018,N_15795);
or U16752 (N_16752,N_15335,N_15419);
nor U16753 (N_16753,N_15149,N_15012);
nand U16754 (N_16754,N_15892,N_15231);
xor U16755 (N_16755,N_15492,N_15012);
xnor U16756 (N_16756,N_15297,N_15010);
xnor U16757 (N_16757,N_15977,N_15299);
or U16758 (N_16758,N_15159,N_15479);
nor U16759 (N_16759,N_15957,N_15714);
nand U16760 (N_16760,N_15833,N_15658);
nand U16761 (N_16761,N_15420,N_15605);
nor U16762 (N_16762,N_15060,N_15101);
nand U16763 (N_16763,N_15689,N_15394);
or U16764 (N_16764,N_15716,N_15089);
nor U16765 (N_16765,N_15236,N_15428);
xnor U16766 (N_16766,N_15242,N_15924);
xnor U16767 (N_16767,N_15463,N_15568);
nand U16768 (N_16768,N_15969,N_15521);
xor U16769 (N_16769,N_15426,N_15132);
nor U16770 (N_16770,N_15175,N_15016);
nand U16771 (N_16771,N_15325,N_15368);
and U16772 (N_16772,N_15094,N_15011);
nand U16773 (N_16773,N_15270,N_15741);
and U16774 (N_16774,N_15077,N_15131);
xnor U16775 (N_16775,N_15381,N_15881);
nor U16776 (N_16776,N_15658,N_15988);
nor U16777 (N_16777,N_15949,N_15126);
and U16778 (N_16778,N_15615,N_15248);
or U16779 (N_16779,N_15706,N_15132);
nand U16780 (N_16780,N_15018,N_15901);
or U16781 (N_16781,N_15226,N_15853);
and U16782 (N_16782,N_15463,N_15827);
xor U16783 (N_16783,N_15760,N_15012);
xor U16784 (N_16784,N_15915,N_15029);
nand U16785 (N_16785,N_15376,N_15399);
nand U16786 (N_16786,N_15128,N_15377);
xor U16787 (N_16787,N_15238,N_15811);
or U16788 (N_16788,N_15973,N_15864);
xor U16789 (N_16789,N_15140,N_15427);
nor U16790 (N_16790,N_15420,N_15834);
nand U16791 (N_16791,N_15295,N_15953);
nand U16792 (N_16792,N_15516,N_15989);
nor U16793 (N_16793,N_15410,N_15821);
or U16794 (N_16794,N_15309,N_15741);
or U16795 (N_16795,N_15724,N_15770);
xnor U16796 (N_16796,N_15469,N_15200);
nand U16797 (N_16797,N_15958,N_15428);
and U16798 (N_16798,N_15840,N_15055);
nand U16799 (N_16799,N_15370,N_15133);
or U16800 (N_16800,N_15352,N_15747);
nor U16801 (N_16801,N_15406,N_15601);
xor U16802 (N_16802,N_15894,N_15102);
nand U16803 (N_16803,N_15127,N_15243);
or U16804 (N_16804,N_15672,N_15847);
xnor U16805 (N_16805,N_15942,N_15020);
xor U16806 (N_16806,N_15287,N_15513);
and U16807 (N_16807,N_15138,N_15980);
or U16808 (N_16808,N_15349,N_15907);
or U16809 (N_16809,N_15344,N_15452);
xnor U16810 (N_16810,N_15639,N_15266);
or U16811 (N_16811,N_15508,N_15183);
nand U16812 (N_16812,N_15444,N_15274);
nor U16813 (N_16813,N_15977,N_15449);
nand U16814 (N_16814,N_15750,N_15396);
xnor U16815 (N_16815,N_15712,N_15755);
nand U16816 (N_16816,N_15979,N_15893);
or U16817 (N_16817,N_15531,N_15862);
xnor U16818 (N_16818,N_15547,N_15441);
or U16819 (N_16819,N_15763,N_15985);
xor U16820 (N_16820,N_15224,N_15983);
nor U16821 (N_16821,N_15362,N_15304);
nor U16822 (N_16822,N_15401,N_15657);
and U16823 (N_16823,N_15213,N_15212);
or U16824 (N_16824,N_15475,N_15846);
nor U16825 (N_16825,N_15869,N_15240);
and U16826 (N_16826,N_15341,N_15232);
xor U16827 (N_16827,N_15946,N_15285);
or U16828 (N_16828,N_15648,N_15481);
xor U16829 (N_16829,N_15958,N_15413);
and U16830 (N_16830,N_15956,N_15668);
and U16831 (N_16831,N_15159,N_15281);
or U16832 (N_16832,N_15206,N_15202);
or U16833 (N_16833,N_15791,N_15581);
or U16834 (N_16834,N_15831,N_15754);
nand U16835 (N_16835,N_15003,N_15845);
nor U16836 (N_16836,N_15784,N_15995);
or U16837 (N_16837,N_15816,N_15984);
nor U16838 (N_16838,N_15322,N_15101);
nand U16839 (N_16839,N_15449,N_15357);
or U16840 (N_16840,N_15159,N_15623);
nand U16841 (N_16841,N_15165,N_15880);
or U16842 (N_16842,N_15387,N_15367);
xor U16843 (N_16843,N_15429,N_15056);
and U16844 (N_16844,N_15036,N_15703);
or U16845 (N_16845,N_15943,N_15271);
nor U16846 (N_16846,N_15755,N_15757);
nor U16847 (N_16847,N_15303,N_15469);
nand U16848 (N_16848,N_15074,N_15736);
and U16849 (N_16849,N_15262,N_15714);
and U16850 (N_16850,N_15763,N_15683);
and U16851 (N_16851,N_15313,N_15014);
or U16852 (N_16852,N_15654,N_15242);
xnor U16853 (N_16853,N_15586,N_15837);
nor U16854 (N_16854,N_15901,N_15908);
nand U16855 (N_16855,N_15416,N_15539);
or U16856 (N_16856,N_15385,N_15574);
and U16857 (N_16857,N_15447,N_15151);
nand U16858 (N_16858,N_15759,N_15982);
and U16859 (N_16859,N_15160,N_15653);
nor U16860 (N_16860,N_15422,N_15816);
nor U16861 (N_16861,N_15265,N_15587);
or U16862 (N_16862,N_15462,N_15958);
nand U16863 (N_16863,N_15735,N_15846);
and U16864 (N_16864,N_15830,N_15538);
nor U16865 (N_16865,N_15602,N_15983);
nor U16866 (N_16866,N_15898,N_15661);
xor U16867 (N_16867,N_15086,N_15230);
nor U16868 (N_16868,N_15769,N_15575);
nand U16869 (N_16869,N_15983,N_15623);
xnor U16870 (N_16870,N_15228,N_15040);
and U16871 (N_16871,N_15098,N_15919);
nor U16872 (N_16872,N_15195,N_15847);
nor U16873 (N_16873,N_15637,N_15359);
nand U16874 (N_16874,N_15768,N_15602);
nand U16875 (N_16875,N_15252,N_15639);
nor U16876 (N_16876,N_15772,N_15757);
nand U16877 (N_16877,N_15824,N_15029);
or U16878 (N_16878,N_15790,N_15285);
xnor U16879 (N_16879,N_15431,N_15036);
nor U16880 (N_16880,N_15797,N_15436);
nand U16881 (N_16881,N_15794,N_15910);
nand U16882 (N_16882,N_15002,N_15007);
nand U16883 (N_16883,N_15250,N_15850);
nand U16884 (N_16884,N_15682,N_15744);
or U16885 (N_16885,N_15663,N_15318);
or U16886 (N_16886,N_15659,N_15056);
nand U16887 (N_16887,N_15922,N_15374);
nand U16888 (N_16888,N_15770,N_15234);
xor U16889 (N_16889,N_15085,N_15867);
nand U16890 (N_16890,N_15731,N_15889);
nor U16891 (N_16891,N_15581,N_15066);
and U16892 (N_16892,N_15947,N_15116);
xor U16893 (N_16893,N_15336,N_15603);
and U16894 (N_16894,N_15507,N_15820);
nand U16895 (N_16895,N_15935,N_15806);
xnor U16896 (N_16896,N_15273,N_15561);
nand U16897 (N_16897,N_15701,N_15106);
nor U16898 (N_16898,N_15505,N_15702);
xor U16899 (N_16899,N_15772,N_15697);
and U16900 (N_16900,N_15795,N_15600);
nand U16901 (N_16901,N_15021,N_15039);
xnor U16902 (N_16902,N_15476,N_15800);
and U16903 (N_16903,N_15056,N_15235);
nand U16904 (N_16904,N_15638,N_15644);
or U16905 (N_16905,N_15344,N_15604);
or U16906 (N_16906,N_15432,N_15096);
or U16907 (N_16907,N_15073,N_15098);
nor U16908 (N_16908,N_15743,N_15683);
nand U16909 (N_16909,N_15588,N_15983);
or U16910 (N_16910,N_15122,N_15522);
or U16911 (N_16911,N_15550,N_15171);
xnor U16912 (N_16912,N_15042,N_15486);
nand U16913 (N_16913,N_15642,N_15088);
nand U16914 (N_16914,N_15689,N_15293);
or U16915 (N_16915,N_15357,N_15617);
xnor U16916 (N_16916,N_15997,N_15583);
and U16917 (N_16917,N_15454,N_15887);
nand U16918 (N_16918,N_15298,N_15011);
and U16919 (N_16919,N_15275,N_15645);
xor U16920 (N_16920,N_15866,N_15218);
and U16921 (N_16921,N_15972,N_15051);
nand U16922 (N_16922,N_15755,N_15223);
xnor U16923 (N_16923,N_15590,N_15659);
nand U16924 (N_16924,N_15496,N_15584);
or U16925 (N_16925,N_15343,N_15629);
nand U16926 (N_16926,N_15464,N_15220);
xnor U16927 (N_16927,N_15624,N_15262);
and U16928 (N_16928,N_15392,N_15738);
nand U16929 (N_16929,N_15674,N_15641);
nand U16930 (N_16930,N_15527,N_15382);
or U16931 (N_16931,N_15950,N_15407);
nand U16932 (N_16932,N_15051,N_15746);
nand U16933 (N_16933,N_15735,N_15643);
or U16934 (N_16934,N_15597,N_15932);
or U16935 (N_16935,N_15658,N_15983);
nand U16936 (N_16936,N_15534,N_15816);
or U16937 (N_16937,N_15441,N_15362);
nor U16938 (N_16938,N_15699,N_15255);
nor U16939 (N_16939,N_15771,N_15799);
nor U16940 (N_16940,N_15074,N_15441);
nand U16941 (N_16941,N_15843,N_15005);
nor U16942 (N_16942,N_15286,N_15957);
nor U16943 (N_16943,N_15763,N_15645);
and U16944 (N_16944,N_15886,N_15871);
and U16945 (N_16945,N_15995,N_15208);
or U16946 (N_16946,N_15486,N_15937);
nor U16947 (N_16947,N_15255,N_15867);
nand U16948 (N_16948,N_15117,N_15209);
xnor U16949 (N_16949,N_15165,N_15839);
nor U16950 (N_16950,N_15038,N_15163);
nor U16951 (N_16951,N_15320,N_15926);
and U16952 (N_16952,N_15052,N_15711);
nand U16953 (N_16953,N_15799,N_15928);
or U16954 (N_16954,N_15621,N_15272);
nand U16955 (N_16955,N_15179,N_15070);
or U16956 (N_16956,N_15835,N_15118);
nand U16957 (N_16957,N_15038,N_15767);
xnor U16958 (N_16958,N_15812,N_15208);
nor U16959 (N_16959,N_15929,N_15800);
nand U16960 (N_16960,N_15467,N_15719);
xnor U16961 (N_16961,N_15682,N_15064);
and U16962 (N_16962,N_15603,N_15571);
nand U16963 (N_16963,N_15666,N_15465);
and U16964 (N_16964,N_15026,N_15526);
nor U16965 (N_16965,N_15018,N_15898);
and U16966 (N_16966,N_15044,N_15262);
xnor U16967 (N_16967,N_15672,N_15324);
nor U16968 (N_16968,N_15164,N_15220);
xnor U16969 (N_16969,N_15712,N_15886);
nor U16970 (N_16970,N_15459,N_15527);
xnor U16971 (N_16971,N_15060,N_15962);
nor U16972 (N_16972,N_15145,N_15888);
xnor U16973 (N_16973,N_15088,N_15438);
nand U16974 (N_16974,N_15973,N_15935);
or U16975 (N_16975,N_15848,N_15516);
and U16976 (N_16976,N_15777,N_15996);
or U16977 (N_16977,N_15540,N_15020);
xor U16978 (N_16978,N_15982,N_15684);
or U16979 (N_16979,N_15189,N_15084);
xor U16980 (N_16980,N_15091,N_15158);
nor U16981 (N_16981,N_15079,N_15591);
nand U16982 (N_16982,N_15634,N_15565);
or U16983 (N_16983,N_15418,N_15429);
and U16984 (N_16984,N_15998,N_15660);
xor U16985 (N_16985,N_15268,N_15820);
nor U16986 (N_16986,N_15659,N_15194);
nand U16987 (N_16987,N_15019,N_15504);
and U16988 (N_16988,N_15988,N_15967);
nor U16989 (N_16989,N_15933,N_15099);
and U16990 (N_16990,N_15755,N_15435);
or U16991 (N_16991,N_15160,N_15355);
or U16992 (N_16992,N_15128,N_15034);
xnor U16993 (N_16993,N_15993,N_15766);
and U16994 (N_16994,N_15643,N_15326);
nor U16995 (N_16995,N_15645,N_15399);
and U16996 (N_16996,N_15165,N_15904);
xnor U16997 (N_16997,N_15270,N_15251);
xnor U16998 (N_16998,N_15427,N_15297);
nor U16999 (N_16999,N_15983,N_15637);
xor U17000 (N_17000,N_16836,N_16175);
and U17001 (N_17001,N_16472,N_16545);
xor U17002 (N_17002,N_16172,N_16881);
nor U17003 (N_17003,N_16916,N_16627);
nand U17004 (N_17004,N_16827,N_16796);
and U17005 (N_17005,N_16416,N_16092);
or U17006 (N_17006,N_16270,N_16862);
nand U17007 (N_17007,N_16927,N_16804);
nand U17008 (N_17008,N_16769,N_16753);
and U17009 (N_17009,N_16053,N_16737);
and U17010 (N_17010,N_16992,N_16693);
nor U17011 (N_17011,N_16157,N_16715);
nor U17012 (N_17012,N_16022,N_16949);
nand U17013 (N_17013,N_16406,N_16631);
or U17014 (N_17014,N_16476,N_16512);
nand U17015 (N_17015,N_16444,N_16784);
and U17016 (N_17016,N_16371,N_16634);
nand U17017 (N_17017,N_16780,N_16125);
xnor U17018 (N_17018,N_16642,N_16317);
and U17019 (N_17019,N_16541,N_16695);
or U17020 (N_17020,N_16795,N_16523);
nand U17021 (N_17021,N_16132,N_16121);
or U17022 (N_17022,N_16391,N_16962);
nor U17023 (N_17023,N_16341,N_16837);
or U17024 (N_17024,N_16577,N_16338);
and U17025 (N_17025,N_16483,N_16783);
or U17026 (N_17026,N_16449,N_16332);
xor U17027 (N_17027,N_16787,N_16032);
xnor U17028 (N_17028,N_16785,N_16115);
nor U17029 (N_17029,N_16537,N_16832);
or U17030 (N_17030,N_16180,N_16249);
or U17031 (N_17031,N_16434,N_16245);
nand U17032 (N_17032,N_16812,N_16575);
nor U17033 (N_17033,N_16681,N_16716);
nor U17034 (N_17034,N_16727,N_16357);
or U17035 (N_17035,N_16899,N_16387);
xnor U17036 (N_17036,N_16898,N_16935);
xor U17037 (N_17037,N_16581,N_16934);
nor U17038 (N_17038,N_16134,N_16010);
xnor U17039 (N_17039,N_16845,N_16509);
xor U17040 (N_17040,N_16858,N_16603);
and U17041 (N_17041,N_16493,N_16351);
or U17042 (N_17042,N_16422,N_16446);
xor U17043 (N_17043,N_16637,N_16551);
nand U17044 (N_17044,N_16869,N_16366);
nand U17045 (N_17045,N_16739,N_16518);
or U17046 (N_17046,N_16432,N_16177);
or U17047 (N_17047,N_16385,N_16722);
or U17048 (N_17048,N_16275,N_16081);
xor U17049 (N_17049,N_16638,N_16356);
or U17050 (N_17050,N_16808,N_16141);
and U17051 (N_17051,N_16209,N_16268);
nor U17052 (N_17052,N_16571,N_16654);
nand U17053 (N_17053,N_16570,N_16191);
or U17054 (N_17054,N_16254,N_16590);
nor U17055 (N_17055,N_16677,N_16643);
nor U17056 (N_17056,N_16520,N_16706);
nor U17057 (N_17057,N_16398,N_16792);
xor U17058 (N_17058,N_16324,N_16563);
nand U17059 (N_17059,N_16798,N_16516);
nor U17060 (N_17060,N_16376,N_16912);
xor U17061 (N_17061,N_16770,N_16131);
xor U17062 (N_17062,N_16861,N_16276);
xor U17063 (N_17063,N_16743,N_16610);
nor U17064 (N_17064,N_16136,N_16891);
xor U17065 (N_17065,N_16561,N_16670);
xor U17066 (N_17066,N_16467,N_16182);
nor U17067 (N_17067,N_16764,N_16781);
and U17068 (N_17068,N_16207,N_16395);
nor U17069 (N_17069,N_16421,N_16198);
and U17070 (N_17070,N_16223,N_16860);
xnor U17071 (N_17071,N_16128,N_16194);
nor U17072 (N_17072,N_16224,N_16025);
nand U17073 (N_17073,N_16246,N_16323);
and U17074 (N_17074,N_16761,N_16041);
nor U17075 (N_17075,N_16419,N_16777);
and U17076 (N_17076,N_16502,N_16913);
nand U17077 (N_17077,N_16863,N_16088);
nor U17078 (N_17078,N_16091,N_16400);
xor U17079 (N_17079,N_16242,N_16353);
nand U17080 (N_17080,N_16187,N_16925);
nor U17081 (N_17081,N_16468,N_16280);
or U17082 (N_17082,N_16622,N_16582);
nor U17083 (N_17083,N_16601,N_16261);
or U17084 (N_17084,N_16847,N_16953);
nor U17085 (N_17085,N_16647,N_16973);
nor U17086 (N_17086,N_16469,N_16386);
xnor U17087 (N_17087,N_16217,N_16308);
xor U17088 (N_17088,N_16407,N_16384);
xor U17089 (N_17089,N_16750,N_16564);
xor U17090 (N_17090,N_16604,N_16124);
xor U17091 (N_17091,N_16515,N_16184);
nand U17092 (N_17092,N_16746,N_16623);
xnor U17093 (N_17093,N_16758,N_16521);
and U17094 (N_17094,N_16077,N_16440);
nor U17095 (N_17095,N_16201,N_16807);
nand U17096 (N_17096,N_16292,N_16215);
nand U17097 (N_17097,N_16890,N_16596);
or U17098 (N_17098,N_16549,N_16287);
or U17099 (N_17099,N_16733,N_16969);
xnor U17100 (N_17100,N_16165,N_16649);
xnor U17101 (N_17101,N_16364,N_16546);
nand U17102 (N_17102,N_16170,N_16282);
nand U17103 (N_17103,N_16848,N_16679);
nor U17104 (N_17104,N_16797,N_16240);
or U17105 (N_17105,N_16116,N_16361);
and U17106 (N_17106,N_16877,N_16105);
xor U17107 (N_17107,N_16085,N_16882);
and U17108 (N_17108,N_16906,N_16316);
nand U17109 (N_17109,N_16613,N_16894);
nor U17110 (N_17110,N_16293,N_16760);
or U17111 (N_17111,N_16667,N_16218);
or U17112 (N_17112,N_16803,N_16955);
nor U17113 (N_17113,N_16352,N_16363);
nand U17114 (N_17114,N_16956,N_16045);
or U17115 (N_17115,N_16993,N_16489);
and U17116 (N_17116,N_16745,N_16196);
nand U17117 (N_17117,N_16931,N_16004);
nand U17118 (N_17118,N_16097,N_16701);
xor U17119 (N_17119,N_16021,N_16872);
or U17120 (N_17120,N_16926,N_16311);
nand U17121 (N_17121,N_16548,N_16148);
or U17122 (N_17122,N_16763,N_16011);
or U17123 (N_17123,N_16833,N_16789);
nor U17124 (N_17124,N_16979,N_16768);
nand U17125 (N_17125,N_16174,N_16854);
nor U17126 (N_17126,N_16988,N_16164);
xor U17127 (N_17127,N_16943,N_16598);
and U17128 (N_17128,N_16285,N_16806);
or U17129 (N_17129,N_16463,N_16216);
nand U17130 (N_17130,N_16040,N_16110);
xor U17131 (N_17131,N_16936,N_16016);
or U17132 (N_17132,N_16714,N_16122);
or U17133 (N_17133,N_16436,N_16241);
xnor U17134 (N_17134,N_16542,N_16661);
xor U17135 (N_17135,N_16248,N_16402);
nor U17136 (N_17136,N_16584,N_16726);
or U17137 (N_17137,N_16100,N_16648);
nand U17138 (N_17138,N_16461,N_16659);
nor U17139 (N_17139,N_16058,N_16499);
or U17140 (N_17140,N_16056,N_16220);
and U17141 (N_17141,N_16297,N_16072);
xor U17142 (N_17142,N_16809,N_16388);
nand U17143 (N_17143,N_16871,N_16347);
or U17144 (N_17144,N_16612,N_16756);
xnor U17145 (N_17145,N_16123,N_16686);
nor U17146 (N_17146,N_16015,N_16178);
nand U17147 (N_17147,N_16909,N_16828);
or U17148 (N_17148,N_16409,N_16961);
nor U17149 (N_17149,N_16660,N_16901);
or U17150 (N_17150,N_16873,N_16405);
or U17151 (N_17151,N_16445,N_16288);
and U17152 (N_17152,N_16102,N_16491);
nor U17153 (N_17153,N_16080,N_16732);
xor U17154 (N_17154,N_16908,N_16597);
xnor U17155 (N_17155,N_16876,N_16083);
xnor U17156 (N_17156,N_16206,N_16645);
nor U17157 (N_17157,N_16569,N_16013);
and U17158 (N_17158,N_16629,N_16382);
nor U17159 (N_17159,N_16046,N_16576);
xor U17160 (N_17160,N_16999,N_16555);
xnor U17161 (N_17161,N_16204,N_16298);
xnor U17162 (N_17162,N_16572,N_16062);
or U17163 (N_17163,N_16984,N_16458);
nor U17164 (N_17164,N_16525,N_16920);
nor U17165 (N_17165,N_16967,N_16651);
or U17166 (N_17166,N_16104,N_16778);
nor U17167 (N_17167,N_16118,N_16611);
nor U17168 (N_17168,N_16676,N_16754);
and U17169 (N_17169,N_16336,N_16031);
nor U17170 (N_17170,N_16766,N_16375);
xnor U17171 (N_17171,N_16673,N_16782);
nor U17172 (N_17172,N_16420,N_16857);
or U17173 (N_17173,N_16921,N_16154);
nor U17174 (N_17174,N_16729,N_16239);
nor U17175 (N_17175,N_16138,N_16001);
nor U17176 (N_17176,N_16600,N_16079);
or U17177 (N_17177,N_16109,N_16635);
or U17178 (N_17178,N_16163,N_16482);
xnor U17179 (N_17179,N_16199,N_16625);
nand U17180 (N_17180,N_16399,N_16313);
and U17181 (N_17181,N_16672,N_16291);
and U17182 (N_17182,N_16008,N_16579);
nor U17183 (N_17183,N_16543,N_16552);
nor U17184 (N_17184,N_16284,N_16488);
nor U17185 (N_17185,N_16390,N_16996);
nand U17186 (N_17186,N_16724,N_16960);
xor U17187 (N_17187,N_16617,N_16773);
and U17188 (N_17188,N_16588,N_16533);
nand U17189 (N_17189,N_16306,N_16302);
or U17190 (N_17190,N_16107,N_16067);
nand U17191 (N_17191,N_16428,N_16158);
or U17192 (N_17192,N_16071,N_16964);
xor U17193 (N_17193,N_16933,N_16595);
and U17194 (N_17194,N_16817,N_16179);
xor U17195 (N_17195,N_16972,N_16559);
or U17196 (N_17196,N_16139,N_16208);
or U17197 (N_17197,N_16707,N_16719);
nor U17198 (N_17198,N_16879,N_16700);
nor U17199 (N_17199,N_16819,N_16678);
nand U17200 (N_17200,N_16294,N_16279);
nand U17201 (N_17201,N_16012,N_16007);
or U17202 (N_17202,N_16917,N_16839);
nor U17203 (N_17203,N_16003,N_16277);
and U17204 (N_17204,N_16456,N_16583);
nor U17205 (N_17205,N_16404,N_16619);
and U17206 (N_17206,N_16959,N_16663);
nor U17207 (N_17207,N_16038,N_16334);
nor U17208 (N_17208,N_16259,N_16029);
or U17209 (N_17209,N_16915,N_16704);
xnor U17210 (N_17210,N_16900,N_16143);
and U17211 (N_17211,N_16705,N_16903);
xnor U17212 (N_17212,N_16103,N_16566);
nand U17213 (N_17213,N_16337,N_16618);
or U17214 (N_17214,N_16066,N_16286);
xor U17215 (N_17215,N_16599,N_16723);
nand U17216 (N_17216,N_16821,N_16851);
xnor U17217 (N_17217,N_16197,N_16522);
nand U17218 (N_17218,N_16813,N_16466);
and U17219 (N_17219,N_16048,N_16980);
or U17220 (N_17220,N_16084,N_16271);
nor U17221 (N_17221,N_16859,N_16310);
nand U17222 (N_17222,N_16593,N_16236);
nand U17223 (N_17223,N_16650,N_16687);
nor U17224 (N_17224,N_16305,N_16602);
xor U17225 (N_17225,N_16547,N_16800);
nand U17226 (N_17226,N_16843,N_16195);
or U17227 (N_17227,N_16986,N_16145);
nand U17228 (N_17228,N_16811,N_16691);
and U17229 (N_17229,N_16896,N_16892);
nor U17230 (N_17230,N_16168,N_16633);
and U17231 (N_17231,N_16354,N_16429);
nor U17232 (N_17232,N_16089,N_16640);
xor U17233 (N_17233,N_16978,N_16414);
and U17234 (N_17234,N_16529,N_16674);
or U17235 (N_17235,N_16653,N_16300);
or U17236 (N_17236,N_16093,N_16607);
nand U17237 (N_17237,N_16658,N_16322);
and U17238 (N_17238,N_16856,N_16689);
and U17239 (N_17239,N_16159,N_16692);
or U17240 (N_17240,N_16940,N_16558);
nand U17241 (N_17241,N_16269,N_16675);
xor U17242 (N_17242,N_16477,N_16063);
nand U17243 (N_17243,N_16911,N_16776);
xnor U17244 (N_17244,N_16233,N_16929);
nand U17245 (N_17245,N_16744,N_16481);
nand U17246 (N_17246,N_16169,N_16668);
nand U17247 (N_17247,N_16887,N_16771);
nand U17248 (N_17248,N_16329,N_16786);
and U17249 (N_17249,N_16137,N_16874);
nor U17250 (N_17250,N_16225,N_16709);
and U17251 (N_17251,N_16496,N_16574);
nand U17252 (N_17252,N_16055,N_16460);
nor U17253 (N_17253,N_16788,N_16304);
and U17254 (N_17254,N_16765,N_16479);
and U17255 (N_17255,N_16680,N_16203);
or U17256 (N_17256,N_16235,N_16365);
xnor U17257 (N_17257,N_16227,N_16262);
xor U17258 (N_17258,N_16315,N_16657);
and U17259 (N_17259,N_16902,N_16530);
or U17260 (N_17260,N_16202,N_16487);
and U17261 (N_17261,N_16970,N_16822);
nor U17262 (N_17262,N_16866,N_16303);
nand U17263 (N_17263,N_16928,N_16826);
and U17264 (N_17264,N_16741,N_16738);
nand U17265 (N_17265,N_16824,N_16345);
nor U17266 (N_17266,N_16205,N_16578);
xnor U17267 (N_17267,N_16621,N_16005);
nand U17268 (N_17268,N_16507,N_16907);
or U17269 (N_17269,N_16646,N_16325);
xor U17270 (N_17270,N_16888,N_16794);
or U17271 (N_17271,N_16231,N_16247);
and U17272 (N_17272,N_16362,N_16255);
nand U17273 (N_17273,N_16162,N_16717);
nor U17274 (N_17274,N_16568,N_16752);
nor U17275 (N_17275,N_16396,N_16251);
nor U17276 (N_17276,N_16181,N_16922);
xnor U17277 (N_17277,N_16731,N_16553);
and U17278 (N_17278,N_16885,N_16096);
nand U17279 (N_17279,N_16266,N_16265);
xnor U17280 (N_17280,N_16358,N_16470);
nand U17281 (N_17281,N_16020,N_16439);
xor U17282 (N_17282,N_16868,N_16014);
nand U17283 (N_17283,N_16447,N_16526);
nor U17284 (N_17284,N_16319,N_16968);
or U17285 (N_17285,N_16682,N_16283);
and U17286 (N_17286,N_16383,N_16531);
nor U17287 (N_17287,N_16260,N_16135);
nor U17288 (N_17288,N_16052,N_16026);
nand U17289 (N_17289,N_16703,N_16171);
xor U17290 (N_17290,N_16702,N_16000);
or U17291 (N_17291,N_16699,N_16513);
nor U17292 (N_17292,N_16560,N_16173);
nor U17293 (N_17293,N_16278,N_16937);
nand U17294 (N_17294,N_16229,N_16485);
xnor U17295 (N_17295,N_16274,N_16985);
or U17296 (N_17296,N_16453,N_16186);
nor U17297 (N_17297,N_16348,N_16728);
and U17298 (N_17298,N_16114,N_16327);
nor U17299 (N_17299,N_16594,N_16591);
or U17300 (N_17300,N_16587,N_16867);
xor U17301 (N_17301,N_16910,N_16688);
nand U17302 (N_17302,N_16842,N_16636);
xor U17303 (N_17303,N_16430,N_16111);
or U17304 (N_17304,N_16987,N_16814);
xnor U17305 (N_17305,N_16256,N_16721);
xor U17306 (N_17306,N_16257,N_16698);
nand U17307 (N_17307,N_16374,N_16024);
xor U17308 (N_17308,N_16144,N_16639);
nand U17309 (N_17309,N_16608,N_16090);
or U17310 (N_17310,N_16027,N_16994);
or U17311 (N_17311,N_16497,N_16065);
or U17312 (N_17312,N_16219,N_16825);
nor U17313 (N_17313,N_16142,N_16585);
and U17314 (N_17314,N_16425,N_16870);
or U17315 (N_17315,N_16050,N_16448);
and U17316 (N_17316,N_16340,N_16036);
nand U17317 (N_17317,N_16947,N_16018);
or U17318 (N_17318,N_16441,N_16944);
xor U17319 (N_17319,N_16464,N_16343);
nor U17320 (N_17320,N_16393,N_16975);
nand U17321 (N_17321,N_16480,N_16438);
nand U17322 (N_17322,N_16685,N_16991);
nor U17323 (N_17323,N_16711,N_16289);
xnor U17324 (N_17324,N_16370,N_16401);
and U17325 (N_17325,N_16150,N_16326);
nand U17326 (N_17326,N_16989,N_16818);
nand U17327 (N_17327,N_16212,N_16147);
nand U17328 (N_17328,N_16054,N_16829);
xnor U17329 (N_17329,N_16963,N_16210);
nand U17330 (N_17330,N_16117,N_16410);
xnor U17331 (N_17331,N_16495,N_16697);
nand U17332 (N_17332,N_16296,N_16995);
nor U17333 (N_17333,N_16958,N_16492);
and U17334 (N_17334,N_16751,N_16234);
and U17335 (N_17335,N_16043,N_16415);
xnor U17336 (N_17336,N_16849,N_16889);
xor U17337 (N_17337,N_16330,N_16632);
or U17338 (N_17338,N_16474,N_16539);
xor U17339 (N_17339,N_16919,N_16006);
nor U17340 (N_17340,N_16793,N_16309);
nor U17341 (N_17341,N_16450,N_16321);
nand U17342 (N_17342,N_16683,N_16748);
nand U17343 (N_17343,N_16883,N_16380);
or U17344 (N_17344,N_16226,N_16238);
xnor U17345 (N_17345,N_16258,N_16562);
nand U17346 (N_17346,N_16267,N_16615);
xnor U17347 (N_17347,N_16880,N_16228);
and U17348 (N_17348,N_16759,N_16853);
nand U17349 (N_17349,N_16835,N_16662);
nand U17350 (N_17350,N_16830,N_16342);
nand U17351 (N_17351,N_16802,N_16424);
nand U17352 (N_17352,N_16630,N_16451);
nor U17353 (N_17353,N_16433,N_16965);
or U17354 (N_17354,N_16166,N_16816);
nor U17355 (N_17355,N_16427,N_16185);
nand U17356 (N_17356,N_16127,N_16360);
nand U17357 (N_17357,N_16408,N_16801);
xor U17358 (N_17358,N_16455,N_16734);
and U17359 (N_17359,N_16126,N_16775);
and U17360 (N_17360,N_16740,N_16914);
nor U17361 (N_17361,N_16534,N_16767);
or U17362 (N_17362,N_16221,N_16047);
nand U17363 (N_17363,N_16799,N_16389);
or U17364 (N_17364,N_16156,N_16815);
nand U17365 (N_17365,N_16684,N_16418);
nor U17366 (N_17366,N_16951,N_16503);
and U17367 (N_17367,N_16544,N_16098);
nor U17368 (N_17368,N_16443,N_16772);
or U17369 (N_17369,N_16606,N_16344);
or U17370 (N_17370,N_16214,N_16243);
and U17371 (N_17371,N_16982,N_16550);
and U17372 (N_17372,N_16791,N_16060);
nor U17373 (N_17373,N_16078,N_16459);
nor U17374 (N_17374,N_16412,N_16379);
and U17375 (N_17375,N_16666,N_16997);
or U17376 (N_17376,N_16932,N_16397);
nor U17377 (N_17377,N_16101,N_16211);
or U17378 (N_17378,N_16718,N_16656);
nor U17379 (N_17379,N_16253,N_16230);
and U17380 (N_17380,N_16974,N_16712);
or U17381 (N_17381,N_16002,N_16232);
xor U17382 (N_17382,N_16517,N_16328);
and U17383 (N_17383,N_16130,N_16318);
nand U17384 (N_17384,N_16017,N_16841);
xor U17385 (N_17385,N_16314,N_16536);
or U17386 (N_17386,N_16998,N_16435);
and U17387 (N_17387,N_16494,N_16565);
nor U17388 (N_17388,N_16805,N_16167);
nand U17389 (N_17389,N_16950,N_16977);
and U17390 (N_17390,N_16349,N_16696);
nor U17391 (N_17391,N_16957,N_16592);
or U17392 (N_17392,N_16510,N_16381);
xor U17393 (N_17393,N_16075,N_16628);
xnor U17394 (N_17394,N_16884,N_16735);
and U17395 (N_17395,N_16664,N_16264);
nor U17396 (N_17396,N_16690,N_16244);
nor U17397 (N_17397,N_16411,N_16140);
xor U17398 (N_17398,N_16501,N_16665);
or U17399 (N_17399,N_16034,N_16059);
nor U17400 (N_17400,N_16064,N_16426);
nand U17401 (N_17401,N_16367,N_16971);
nand U17402 (N_17402,N_16535,N_16009);
and U17403 (N_17403,N_16616,N_16878);
and U17404 (N_17404,N_16082,N_16373);
xnor U17405 (N_17405,N_16457,N_16073);
and U17406 (N_17406,N_16834,N_16473);
xnor U17407 (N_17407,N_16042,N_16966);
xor U17408 (N_17408,N_16213,N_16790);
xor U17409 (N_17409,N_16146,N_16442);
nand U17410 (N_17410,N_16200,N_16312);
nor U17411 (N_17411,N_16838,N_16035);
and U17412 (N_17412,N_16307,N_16755);
xnor U17413 (N_17413,N_16061,N_16762);
or U17414 (N_17414,N_16129,N_16589);
or U17415 (N_17415,N_16567,N_16850);
and U17416 (N_17416,N_16624,N_16295);
xor U17417 (N_17417,N_16413,N_16188);
or U17418 (N_17418,N_16049,N_16272);
nand U17419 (N_17419,N_16160,N_16720);
nand U17420 (N_17420,N_16694,N_16671);
xnor U17421 (N_17421,N_16051,N_16301);
or U17422 (N_17422,N_16532,N_16133);
nand U17423 (N_17423,N_16644,N_16475);
xnor U17424 (N_17424,N_16840,N_16923);
xor U17425 (N_17425,N_16070,N_16946);
xor U17426 (N_17426,N_16320,N_16904);
and U17427 (N_17427,N_16190,N_16151);
and U17428 (N_17428,N_16019,N_16193);
xnor U17429 (N_17429,N_16176,N_16844);
nor U17430 (N_17430,N_16189,N_16981);
or U17431 (N_17431,N_16948,N_16846);
and U17432 (N_17432,N_16508,N_16895);
nand U17433 (N_17433,N_16641,N_16465);
nand U17434 (N_17434,N_16037,N_16368);
or U17435 (N_17435,N_16511,N_16823);
xnor U17436 (N_17436,N_16945,N_16852);
nand U17437 (N_17437,N_16939,N_16030);
xnor U17438 (N_17438,N_16586,N_16669);
xor U17439 (N_17439,N_16237,N_16941);
nand U17440 (N_17440,N_16346,N_16620);
nor U17441 (N_17441,N_16153,N_16897);
nor U17442 (N_17442,N_16954,N_16486);
or U17443 (N_17443,N_16905,N_16614);
and U17444 (N_17444,N_16730,N_16120);
and U17445 (N_17445,N_16655,N_16335);
xnor U17446 (N_17446,N_16222,N_16355);
nand U17447 (N_17447,N_16099,N_16865);
nor U17448 (N_17448,N_16527,N_16263);
xor U17449 (N_17449,N_16273,N_16506);
and U17450 (N_17450,N_16454,N_16192);
nor U17451 (N_17451,N_16039,N_16757);
or U17452 (N_17452,N_16113,N_16417);
nor U17453 (N_17453,N_16094,N_16875);
and U17454 (N_17454,N_16106,N_16252);
nor U17455 (N_17455,N_16299,N_16749);
nor U17456 (N_17456,N_16095,N_16076);
xnor U17457 (N_17457,N_16983,N_16990);
nor U17458 (N_17458,N_16924,N_16023);
xnor U17459 (N_17459,N_16779,N_16573);
nor U17460 (N_17460,N_16423,N_16514);
or U17461 (N_17461,N_16250,N_16952);
and U17462 (N_17462,N_16074,N_16725);
nor U17463 (N_17463,N_16976,N_16033);
nor U17464 (N_17464,N_16044,N_16930);
nor U17465 (N_17465,N_16333,N_16339);
xor U17466 (N_17466,N_16708,N_16736);
or U17467 (N_17467,N_16161,N_16528);
nor U17468 (N_17468,N_16069,N_16938);
or U17469 (N_17469,N_16372,N_16112);
and U17470 (N_17470,N_16462,N_16498);
nand U17471 (N_17471,N_16152,N_16331);
xor U17472 (N_17472,N_16377,N_16392);
xnor U17473 (N_17473,N_16504,N_16554);
nand U17474 (N_17474,N_16810,N_16713);
nor U17475 (N_17475,N_16556,N_16057);
nor U17476 (N_17476,N_16359,N_16710);
or U17477 (N_17477,N_16918,N_16942);
and U17478 (N_17478,N_16864,N_16369);
and U17479 (N_17479,N_16538,N_16500);
and U17480 (N_17480,N_16403,N_16484);
or U17481 (N_17481,N_16281,N_16028);
nor U17482 (N_17482,N_16478,N_16831);
nand U17483 (N_17483,N_16452,N_16855);
and U17484 (N_17484,N_16437,N_16290);
nand U17485 (N_17485,N_16519,N_16087);
nand U17486 (N_17486,N_16490,N_16394);
and U17487 (N_17487,N_16471,N_16068);
xnor U17488 (N_17488,N_16086,N_16886);
and U17489 (N_17489,N_16605,N_16183);
nand U17490 (N_17490,N_16626,N_16149);
and U17491 (N_17491,N_16524,N_16505);
xor U17492 (N_17492,N_16609,N_16557);
nor U17493 (N_17493,N_16431,N_16820);
or U17494 (N_17494,N_16155,N_16108);
or U17495 (N_17495,N_16893,N_16119);
or U17496 (N_17496,N_16580,N_16742);
nor U17497 (N_17497,N_16774,N_16747);
nor U17498 (N_17498,N_16652,N_16378);
nand U17499 (N_17499,N_16540,N_16350);
nor U17500 (N_17500,N_16154,N_16319);
nor U17501 (N_17501,N_16694,N_16153);
or U17502 (N_17502,N_16522,N_16155);
nor U17503 (N_17503,N_16784,N_16473);
nand U17504 (N_17504,N_16271,N_16193);
or U17505 (N_17505,N_16190,N_16150);
or U17506 (N_17506,N_16734,N_16922);
or U17507 (N_17507,N_16414,N_16595);
nand U17508 (N_17508,N_16203,N_16968);
nand U17509 (N_17509,N_16872,N_16853);
and U17510 (N_17510,N_16721,N_16191);
or U17511 (N_17511,N_16643,N_16654);
nor U17512 (N_17512,N_16172,N_16491);
nand U17513 (N_17513,N_16705,N_16928);
nor U17514 (N_17514,N_16869,N_16311);
xnor U17515 (N_17515,N_16937,N_16589);
xor U17516 (N_17516,N_16340,N_16270);
nand U17517 (N_17517,N_16798,N_16544);
and U17518 (N_17518,N_16403,N_16701);
nor U17519 (N_17519,N_16734,N_16489);
or U17520 (N_17520,N_16331,N_16082);
xnor U17521 (N_17521,N_16853,N_16835);
or U17522 (N_17522,N_16112,N_16958);
nand U17523 (N_17523,N_16643,N_16610);
and U17524 (N_17524,N_16870,N_16658);
nor U17525 (N_17525,N_16461,N_16613);
and U17526 (N_17526,N_16774,N_16756);
and U17527 (N_17527,N_16588,N_16205);
xor U17528 (N_17528,N_16740,N_16467);
or U17529 (N_17529,N_16407,N_16091);
and U17530 (N_17530,N_16686,N_16337);
or U17531 (N_17531,N_16772,N_16883);
nor U17532 (N_17532,N_16332,N_16924);
or U17533 (N_17533,N_16976,N_16544);
nand U17534 (N_17534,N_16925,N_16381);
nor U17535 (N_17535,N_16815,N_16761);
nor U17536 (N_17536,N_16884,N_16039);
xor U17537 (N_17537,N_16160,N_16208);
or U17538 (N_17538,N_16667,N_16521);
and U17539 (N_17539,N_16836,N_16485);
xnor U17540 (N_17540,N_16583,N_16367);
and U17541 (N_17541,N_16569,N_16270);
xnor U17542 (N_17542,N_16904,N_16850);
or U17543 (N_17543,N_16266,N_16436);
and U17544 (N_17544,N_16617,N_16798);
nor U17545 (N_17545,N_16620,N_16841);
and U17546 (N_17546,N_16107,N_16867);
xor U17547 (N_17547,N_16143,N_16881);
nand U17548 (N_17548,N_16659,N_16316);
or U17549 (N_17549,N_16449,N_16378);
xor U17550 (N_17550,N_16483,N_16652);
xnor U17551 (N_17551,N_16615,N_16147);
nor U17552 (N_17552,N_16527,N_16342);
or U17553 (N_17553,N_16098,N_16570);
or U17554 (N_17554,N_16460,N_16021);
or U17555 (N_17555,N_16539,N_16196);
nand U17556 (N_17556,N_16868,N_16655);
nand U17557 (N_17557,N_16726,N_16234);
or U17558 (N_17558,N_16248,N_16647);
nor U17559 (N_17559,N_16908,N_16795);
nor U17560 (N_17560,N_16741,N_16104);
nand U17561 (N_17561,N_16486,N_16743);
or U17562 (N_17562,N_16946,N_16789);
nand U17563 (N_17563,N_16543,N_16898);
xnor U17564 (N_17564,N_16597,N_16666);
nand U17565 (N_17565,N_16813,N_16033);
and U17566 (N_17566,N_16596,N_16699);
and U17567 (N_17567,N_16477,N_16069);
xor U17568 (N_17568,N_16433,N_16207);
nor U17569 (N_17569,N_16676,N_16763);
xnor U17570 (N_17570,N_16900,N_16344);
nor U17571 (N_17571,N_16715,N_16778);
xnor U17572 (N_17572,N_16948,N_16161);
xor U17573 (N_17573,N_16877,N_16886);
or U17574 (N_17574,N_16123,N_16291);
or U17575 (N_17575,N_16205,N_16674);
and U17576 (N_17576,N_16271,N_16073);
and U17577 (N_17577,N_16203,N_16420);
nand U17578 (N_17578,N_16191,N_16938);
xor U17579 (N_17579,N_16696,N_16528);
nand U17580 (N_17580,N_16314,N_16148);
nand U17581 (N_17581,N_16096,N_16829);
xor U17582 (N_17582,N_16045,N_16367);
nand U17583 (N_17583,N_16911,N_16231);
xnor U17584 (N_17584,N_16299,N_16369);
or U17585 (N_17585,N_16942,N_16912);
or U17586 (N_17586,N_16050,N_16727);
or U17587 (N_17587,N_16072,N_16466);
or U17588 (N_17588,N_16370,N_16916);
nand U17589 (N_17589,N_16845,N_16798);
and U17590 (N_17590,N_16112,N_16270);
and U17591 (N_17591,N_16322,N_16662);
nand U17592 (N_17592,N_16443,N_16580);
or U17593 (N_17593,N_16541,N_16080);
xnor U17594 (N_17594,N_16606,N_16033);
nand U17595 (N_17595,N_16153,N_16677);
nor U17596 (N_17596,N_16211,N_16188);
nand U17597 (N_17597,N_16189,N_16181);
nor U17598 (N_17598,N_16399,N_16757);
nor U17599 (N_17599,N_16407,N_16778);
and U17600 (N_17600,N_16987,N_16190);
nand U17601 (N_17601,N_16901,N_16875);
and U17602 (N_17602,N_16251,N_16813);
xor U17603 (N_17603,N_16757,N_16315);
nand U17604 (N_17604,N_16540,N_16255);
nand U17605 (N_17605,N_16942,N_16887);
or U17606 (N_17606,N_16195,N_16140);
xor U17607 (N_17607,N_16058,N_16237);
or U17608 (N_17608,N_16370,N_16193);
nor U17609 (N_17609,N_16653,N_16986);
and U17610 (N_17610,N_16364,N_16304);
nor U17611 (N_17611,N_16246,N_16430);
or U17612 (N_17612,N_16416,N_16012);
and U17613 (N_17613,N_16446,N_16861);
nor U17614 (N_17614,N_16739,N_16361);
nor U17615 (N_17615,N_16036,N_16341);
or U17616 (N_17616,N_16812,N_16849);
nand U17617 (N_17617,N_16274,N_16823);
nor U17618 (N_17618,N_16323,N_16619);
nand U17619 (N_17619,N_16963,N_16570);
nand U17620 (N_17620,N_16741,N_16685);
xnor U17621 (N_17621,N_16532,N_16747);
xnor U17622 (N_17622,N_16126,N_16320);
nand U17623 (N_17623,N_16056,N_16836);
nor U17624 (N_17624,N_16443,N_16805);
nor U17625 (N_17625,N_16419,N_16044);
nor U17626 (N_17626,N_16905,N_16124);
xnor U17627 (N_17627,N_16289,N_16394);
nand U17628 (N_17628,N_16957,N_16632);
xnor U17629 (N_17629,N_16604,N_16125);
nor U17630 (N_17630,N_16374,N_16318);
or U17631 (N_17631,N_16469,N_16290);
and U17632 (N_17632,N_16067,N_16475);
nor U17633 (N_17633,N_16333,N_16662);
xor U17634 (N_17634,N_16879,N_16190);
or U17635 (N_17635,N_16421,N_16355);
xnor U17636 (N_17636,N_16855,N_16253);
nor U17637 (N_17637,N_16430,N_16168);
or U17638 (N_17638,N_16844,N_16334);
nor U17639 (N_17639,N_16432,N_16875);
nor U17640 (N_17640,N_16248,N_16209);
nor U17641 (N_17641,N_16331,N_16460);
or U17642 (N_17642,N_16798,N_16185);
xor U17643 (N_17643,N_16714,N_16824);
or U17644 (N_17644,N_16098,N_16611);
xnor U17645 (N_17645,N_16310,N_16325);
nand U17646 (N_17646,N_16362,N_16886);
xnor U17647 (N_17647,N_16811,N_16295);
xor U17648 (N_17648,N_16740,N_16040);
and U17649 (N_17649,N_16343,N_16993);
and U17650 (N_17650,N_16206,N_16416);
nand U17651 (N_17651,N_16617,N_16348);
or U17652 (N_17652,N_16351,N_16416);
nand U17653 (N_17653,N_16272,N_16547);
xor U17654 (N_17654,N_16109,N_16713);
nand U17655 (N_17655,N_16300,N_16382);
xor U17656 (N_17656,N_16417,N_16221);
nand U17657 (N_17657,N_16060,N_16710);
nor U17658 (N_17658,N_16060,N_16243);
nor U17659 (N_17659,N_16937,N_16176);
and U17660 (N_17660,N_16067,N_16996);
and U17661 (N_17661,N_16798,N_16702);
nor U17662 (N_17662,N_16522,N_16627);
nor U17663 (N_17663,N_16667,N_16049);
or U17664 (N_17664,N_16959,N_16999);
or U17665 (N_17665,N_16532,N_16613);
xnor U17666 (N_17666,N_16026,N_16908);
and U17667 (N_17667,N_16186,N_16468);
or U17668 (N_17668,N_16380,N_16972);
and U17669 (N_17669,N_16941,N_16940);
and U17670 (N_17670,N_16025,N_16986);
xnor U17671 (N_17671,N_16565,N_16416);
or U17672 (N_17672,N_16220,N_16988);
xor U17673 (N_17673,N_16127,N_16982);
or U17674 (N_17674,N_16649,N_16176);
or U17675 (N_17675,N_16088,N_16930);
nand U17676 (N_17676,N_16409,N_16040);
and U17677 (N_17677,N_16767,N_16857);
xnor U17678 (N_17678,N_16910,N_16489);
nand U17679 (N_17679,N_16762,N_16429);
or U17680 (N_17680,N_16506,N_16950);
and U17681 (N_17681,N_16667,N_16819);
and U17682 (N_17682,N_16283,N_16299);
and U17683 (N_17683,N_16003,N_16988);
nor U17684 (N_17684,N_16199,N_16534);
or U17685 (N_17685,N_16047,N_16373);
and U17686 (N_17686,N_16720,N_16688);
nor U17687 (N_17687,N_16347,N_16301);
or U17688 (N_17688,N_16628,N_16539);
xnor U17689 (N_17689,N_16931,N_16970);
nor U17690 (N_17690,N_16122,N_16180);
and U17691 (N_17691,N_16142,N_16846);
xor U17692 (N_17692,N_16584,N_16613);
nor U17693 (N_17693,N_16811,N_16681);
and U17694 (N_17694,N_16797,N_16475);
or U17695 (N_17695,N_16256,N_16029);
nor U17696 (N_17696,N_16774,N_16908);
xor U17697 (N_17697,N_16870,N_16163);
nor U17698 (N_17698,N_16522,N_16593);
nand U17699 (N_17699,N_16462,N_16614);
and U17700 (N_17700,N_16603,N_16953);
nor U17701 (N_17701,N_16697,N_16093);
and U17702 (N_17702,N_16254,N_16733);
or U17703 (N_17703,N_16988,N_16432);
nand U17704 (N_17704,N_16664,N_16535);
and U17705 (N_17705,N_16790,N_16496);
and U17706 (N_17706,N_16960,N_16039);
or U17707 (N_17707,N_16076,N_16118);
xor U17708 (N_17708,N_16448,N_16165);
or U17709 (N_17709,N_16432,N_16827);
xor U17710 (N_17710,N_16887,N_16176);
xor U17711 (N_17711,N_16306,N_16046);
xnor U17712 (N_17712,N_16043,N_16607);
nand U17713 (N_17713,N_16490,N_16721);
or U17714 (N_17714,N_16893,N_16638);
xor U17715 (N_17715,N_16682,N_16209);
nor U17716 (N_17716,N_16541,N_16713);
and U17717 (N_17717,N_16764,N_16838);
nand U17718 (N_17718,N_16705,N_16484);
nor U17719 (N_17719,N_16831,N_16878);
nand U17720 (N_17720,N_16199,N_16819);
nor U17721 (N_17721,N_16742,N_16290);
nand U17722 (N_17722,N_16349,N_16377);
or U17723 (N_17723,N_16671,N_16303);
nand U17724 (N_17724,N_16719,N_16534);
or U17725 (N_17725,N_16404,N_16756);
nand U17726 (N_17726,N_16360,N_16952);
xnor U17727 (N_17727,N_16654,N_16838);
nor U17728 (N_17728,N_16090,N_16943);
nand U17729 (N_17729,N_16161,N_16013);
nand U17730 (N_17730,N_16654,N_16362);
and U17731 (N_17731,N_16287,N_16887);
nand U17732 (N_17732,N_16128,N_16653);
xnor U17733 (N_17733,N_16953,N_16363);
xor U17734 (N_17734,N_16523,N_16604);
or U17735 (N_17735,N_16298,N_16369);
and U17736 (N_17736,N_16575,N_16838);
xnor U17737 (N_17737,N_16421,N_16115);
and U17738 (N_17738,N_16049,N_16654);
nand U17739 (N_17739,N_16286,N_16551);
nand U17740 (N_17740,N_16416,N_16159);
xnor U17741 (N_17741,N_16357,N_16176);
or U17742 (N_17742,N_16424,N_16784);
nand U17743 (N_17743,N_16548,N_16768);
xnor U17744 (N_17744,N_16032,N_16731);
and U17745 (N_17745,N_16030,N_16936);
nand U17746 (N_17746,N_16973,N_16190);
xnor U17747 (N_17747,N_16618,N_16379);
or U17748 (N_17748,N_16198,N_16971);
nor U17749 (N_17749,N_16958,N_16961);
and U17750 (N_17750,N_16072,N_16024);
xor U17751 (N_17751,N_16910,N_16904);
and U17752 (N_17752,N_16118,N_16868);
or U17753 (N_17753,N_16943,N_16817);
and U17754 (N_17754,N_16892,N_16195);
nor U17755 (N_17755,N_16802,N_16525);
or U17756 (N_17756,N_16243,N_16205);
or U17757 (N_17757,N_16756,N_16565);
or U17758 (N_17758,N_16631,N_16041);
nand U17759 (N_17759,N_16026,N_16171);
and U17760 (N_17760,N_16828,N_16572);
xor U17761 (N_17761,N_16534,N_16911);
nor U17762 (N_17762,N_16339,N_16517);
nor U17763 (N_17763,N_16435,N_16257);
nor U17764 (N_17764,N_16909,N_16374);
xnor U17765 (N_17765,N_16518,N_16126);
nand U17766 (N_17766,N_16954,N_16998);
and U17767 (N_17767,N_16720,N_16936);
nor U17768 (N_17768,N_16065,N_16117);
nor U17769 (N_17769,N_16222,N_16646);
xor U17770 (N_17770,N_16856,N_16780);
and U17771 (N_17771,N_16292,N_16030);
and U17772 (N_17772,N_16330,N_16236);
or U17773 (N_17773,N_16576,N_16573);
or U17774 (N_17774,N_16031,N_16963);
and U17775 (N_17775,N_16423,N_16441);
nand U17776 (N_17776,N_16779,N_16297);
and U17777 (N_17777,N_16628,N_16746);
and U17778 (N_17778,N_16896,N_16157);
xor U17779 (N_17779,N_16896,N_16498);
xor U17780 (N_17780,N_16710,N_16314);
and U17781 (N_17781,N_16647,N_16834);
or U17782 (N_17782,N_16649,N_16377);
nand U17783 (N_17783,N_16210,N_16240);
nand U17784 (N_17784,N_16060,N_16095);
or U17785 (N_17785,N_16631,N_16829);
or U17786 (N_17786,N_16770,N_16362);
nand U17787 (N_17787,N_16928,N_16845);
xor U17788 (N_17788,N_16831,N_16538);
xnor U17789 (N_17789,N_16955,N_16288);
or U17790 (N_17790,N_16051,N_16930);
nand U17791 (N_17791,N_16368,N_16191);
xor U17792 (N_17792,N_16462,N_16362);
or U17793 (N_17793,N_16497,N_16598);
or U17794 (N_17794,N_16860,N_16714);
or U17795 (N_17795,N_16453,N_16119);
and U17796 (N_17796,N_16992,N_16261);
and U17797 (N_17797,N_16112,N_16238);
or U17798 (N_17798,N_16407,N_16633);
xor U17799 (N_17799,N_16553,N_16001);
or U17800 (N_17800,N_16784,N_16007);
and U17801 (N_17801,N_16638,N_16541);
or U17802 (N_17802,N_16806,N_16112);
or U17803 (N_17803,N_16892,N_16306);
xor U17804 (N_17804,N_16558,N_16882);
or U17805 (N_17805,N_16156,N_16122);
and U17806 (N_17806,N_16280,N_16068);
and U17807 (N_17807,N_16056,N_16182);
and U17808 (N_17808,N_16388,N_16972);
nand U17809 (N_17809,N_16954,N_16099);
nor U17810 (N_17810,N_16494,N_16894);
nand U17811 (N_17811,N_16692,N_16179);
nand U17812 (N_17812,N_16600,N_16407);
nand U17813 (N_17813,N_16886,N_16907);
nor U17814 (N_17814,N_16815,N_16599);
nand U17815 (N_17815,N_16265,N_16535);
xor U17816 (N_17816,N_16305,N_16187);
nand U17817 (N_17817,N_16703,N_16264);
nor U17818 (N_17818,N_16131,N_16418);
nand U17819 (N_17819,N_16074,N_16721);
nor U17820 (N_17820,N_16469,N_16137);
nor U17821 (N_17821,N_16923,N_16967);
nor U17822 (N_17822,N_16957,N_16424);
xnor U17823 (N_17823,N_16768,N_16121);
and U17824 (N_17824,N_16829,N_16842);
and U17825 (N_17825,N_16118,N_16047);
nor U17826 (N_17826,N_16430,N_16304);
or U17827 (N_17827,N_16712,N_16588);
and U17828 (N_17828,N_16141,N_16544);
xnor U17829 (N_17829,N_16301,N_16140);
or U17830 (N_17830,N_16060,N_16472);
xnor U17831 (N_17831,N_16641,N_16829);
and U17832 (N_17832,N_16549,N_16621);
and U17833 (N_17833,N_16236,N_16374);
or U17834 (N_17834,N_16285,N_16503);
or U17835 (N_17835,N_16843,N_16334);
nand U17836 (N_17836,N_16605,N_16490);
xor U17837 (N_17837,N_16890,N_16874);
or U17838 (N_17838,N_16142,N_16054);
nand U17839 (N_17839,N_16674,N_16320);
or U17840 (N_17840,N_16546,N_16813);
xnor U17841 (N_17841,N_16028,N_16589);
and U17842 (N_17842,N_16471,N_16330);
nand U17843 (N_17843,N_16074,N_16339);
nand U17844 (N_17844,N_16615,N_16006);
xnor U17845 (N_17845,N_16640,N_16415);
nor U17846 (N_17846,N_16774,N_16785);
nor U17847 (N_17847,N_16675,N_16963);
and U17848 (N_17848,N_16084,N_16805);
nor U17849 (N_17849,N_16776,N_16169);
xor U17850 (N_17850,N_16968,N_16550);
or U17851 (N_17851,N_16972,N_16293);
nor U17852 (N_17852,N_16057,N_16827);
nand U17853 (N_17853,N_16657,N_16462);
and U17854 (N_17854,N_16074,N_16293);
or U17855 (N_17855,N_16349,N_16776);
and U17856 (N_17856,N_16071,N_16490);
and U17857 (N_17857,N_16993,N_16596);
xor U17858 (N_17858,N_16101,N_16910);
or U17859 (N_17859,N_16526,N_16666);
and U17860 (N_17860,N_16186,N_16888);
or U17861 (N_17861,N_16807,N_16583);
nand U17862 (N_17862,N_16382,N_16573);
and U17863 (N_17863,N_16122,N_16292);
and U17864 (N_17864,N_16749,N_16139);
and U17865 (N_17865,N_16254,N_16666);
nand U17866 (N_17866,N_16410,N_16092);
nand U17867 (N_17867,N_16767,N_16148);
nor U17868 (N_17868,N_16316,N_16895);
nor U17869 (N_17869,N_16759,N_16002);
xor U17870 (N_17870,N_16828,N_16773);
xnor U17871 (N_17871,N_16172,N_16560);
or U17872 (N_17872,N_16938,N_16074);
xor U17873 (N_17873,N_16451,N_16197);
xnor U17874 (N_17874,N_16291,N_16406);
nor U17875 (N_17875,N_16858,N_16083);
or U17876 (N_17876,N_16915,N_16995);
or U17877 (N_17877,N_16641,N_16905);
nand U17878 (N_17878,N_16681,N_16942);
nor U17879 (N_17879,N_16416,N_16890);
and U17880 (N_17880,N_16579,N_16812);
nor U17881 (N_17881,N_16962,N_16845);
xnor U17882 (N_17882,N_16193,N_16403);
nor U17883 (N_17883,N_16919,N_16411);
xor U17884 (N_17884,N_16833,N_16640);
nand U17885 (N_17885,N_16488,N_16108);
and U17886 (N_17886,N_16997,N_16058);
nand U17887 (N_17887,N_16956,N_16553);
nand U17888 (N_17888,N_16954,N_16675);
or U17889 (N_17889,N_16688,N_16843);
nand U17890 (N_17890,N_16799,N_16155);
and U17891 (N_17891,N_16729,N_16741);
nand U17892 (N_17892,N_16836,N_16660);
xor U17893 (N_17893,N_16633,N_16804);
nor U17894 (N_17894,N_16827,N_16681);
and U17895 (N_17895,N_16451,N_16356);
or U17896 (N_17896,N_16586,N_16096);
nand U17897 (N_17897,N_16852,N_16880);
or U17898 (N_17898,N_16944,N_16030);
or U17899 (N_17899,N_16333,N_16366);
and U17900 (N_17900,N_16063,N_16594);
nor U17901 (N_17901,N_16505,N_16653);
or U17902 (N_17902,N_16847,N_16608);
or U17903 (N_17903,N_16745,N_16889);
nand U17904 (N_17904,N_16197,N_16190);
xor U17905 (N_17905,N_16216,N_16308);
nand U17906 (N_17906,N_16629,N_16033);
and U17907 (N_17907,N_16433,N_16808);
xnor U17908 (N_17908,N_16763,N_16286);
xnor U17909 (N_17909,N_16910,N_16021);
xnor U17910 (N_17910,N_16014,N_16938);
xnor U17911 (N_17911,N_16042,N_16199);
and U17912 (N_17912,N_16307,N_16398);
and U17913 (N_17913,N_16076,N_16084);
and U17914 (N_17914,N_16295,N_16581);
and U17915 (N_17915,N_16002,N_16117);
nor U17916 (N_17916,N_16300,N_16930);
nand U17917 (N_17917,N_16593,N_16206);
or U17918 (N_17918,N_16537,N_16283);
nand U17919 (N_17919,N_16531,N_16984);
xnor U17920 (N_17920,N_16137,N_16550);
xnor U17921 (N_17921,N_16816,N_16148);
or U17922 (N_17922,N_16926,N_16387);
nor U17923 (N_17923,N_16625,N_16989);
xor U17924 (N_17924,N_16848,N_16469);
or U17925 (N_17925,N_16586,N_16499);
and U17926 (N_17926,N_16975,N_16071);
xor U17927 (N_17927,N_16600,N_16496);
xnor U17928 (N_17928,N_16489,N_16869);
xor U17929 (N_17929,N_16944,N_16804);
xor U17930 (N_17930,N_16260,N_16015);
nor U17931 (N_17931,N_16318,N_16377);
and U17932 (N_17932,N_16224,N_16274);
xnor U17933 (N_17933,N_16633,N_16215);
xnor U17934 (N_17934,N_16903,N_16813);
nor U17935 (N_17935,N_16196,N_16952);
nand U17936 (N_17936,N_16191,N_16754);
and U17937 (N_17937,N_16889,N_16037);
nor U17938 (N_17938,N_16079,N_16687);
nand U17939 (N_17939,N_16644,N_16637);
or U17940 (N_17940,N_16249,N_16403);
and U17941 (N_17941,N_16375,N_16156);
and U17942 (N_17942,N_16612,N_16563);
nor U17943 (N_17943,N_16814,N_16044);
or U17944 (N_17944,N_16250,N_16493);
or U17945 (N_17945,N_16489,N_16466);
nor U17946 (N_17946,N_16922,N_16367);
and U17947 (N_17947,N_16670,N_16326);
nor U17948 (N_17948,N_16737,N_16574);
xor U17949 (N_17949,N_16079,N_16019);
nor U17950 (N_17950,N_16927,N_16386);
nand U17951 (N_17951,N_16330,N_16258);
or U17952 (N_17952,N_16507,N_16900);
nand U17953 (N_17953,N_16993,N_16148);
nor U17954 (N_17954,N_16299,N_16290);
or U17955 (N_17955,N_16325,N_16224);
nand U17956 (N_17956,N_16428,N_16049);
xor U17957 (N_17957,N_16191,N_16886);
nor U17958 (N_17958,N_16927,N_16123);
xnor U17959 (N_17959,N_16078,N_16417);
xnor U17960 (N_17960,N_16108,N_16999);
and U17961 (N_17961,N_16708,N_16931);
or U17962 (N_17962,N_16931,N_16402);
and U17963 (N_17963,N_16646,N_16606);
or U17964 (N_17964,N_16834,N_16298);
and U17965 (N_17965,N_16642,N_16790);
nor U17966 (N_17966,N_16899,N_16039);
xor U17967 (N_17967,N_16749,N_16955);
or U17968 (N_17968,N_16997,N_16062);
nand U17969 (N_17969,N_16394,N_16485);
nor U17970 (N_17970,N_16455,N_16259);
xor U17971 (N_17971,N_16784,N_16820);
nand U17972 (N_17972,N_16983,N_16475);
and U17973 (N_17973,N_16816,N_16929);
xnor U17974 (N_17974,N_16057,N_16357);
and U17975 (N_17975,N_16897,N_16316);
xnor U17976 (N_17976,N_16285,N_16445);
or U17977 (N_17977,N_16932,N_16757);
xor U17978 (N_17978,N_16177,N_16866);
nand U17979 (N_17979,N_16338,N_16623);
nor U17980 (N_17980,N_16144,N_16169);
and U17981 (N_17981,N_16091,N_16037);
xnor U17982 (N_17982,N_16889,N_16634);
xor U17983 (N_17983,N_16389,N_16208);
or U17984 (N_17984,N_16768,N_16080);
and U17985 (N_17985,N_16499,N_16471);
nor U17986 (N_17986,N_16076,N_16454);
xor U17987 (N_17987,N_16652,N_16650);
or U17988 (N_17988,N_16977,N_16289);
nor U17989 (N_17989,N_16756,N_16096);
nand U17990 (N_17990,N_16782,N_16688);
nand U17991 (N_17991,N_16450,N_16170);
or U17992 (N_17992,N_16258,N_16732);
nand U17993 (N_17993,N_16225,N_16432);
nand U17994 (N_17994,N_16705,N_16671);
xnor U17995 (N_17995,N_16577,N_16141);
or U17996 (N_17996,N_16837,N_16993);
or U17997 (N_17997,N_16214,N_16733);
and U17998 (N_17998,N_16806,N_16086);
nor U17999 (N_17999,N_16967,N_16867);
nor U18000 (N_18000,N_17681,N_17631);
nand U18001 (N_18001,N_17876,N_17419);
nand U18002 (N_18002,N_17174,N_17399);
or U18003 (N_18003,N_17221,N_17806);
nand U18004 (N_18004,N_17683,N_17616);
and U18005 (N_18005,N_17461,N_17216);
xnor U18006 (N_18006,N_17226,N_17818);
nand U18007 (N_18007,N_17252,N_17220);
nand U18008 (N_18008,N_17290,N_17870);
nor U18009 (N_18009,N_17327,N_17843);
and U18010 (N_18010,N_17707,N_17502);
nor U18011 (N_18011,N_17137,N_17739);
or U18012 (N_18012,N_17863,N_17073);
and U18013 (N_18013,N_17810,N_17005);
nand U18014 (N_18014,N_17271,N_17170);
xnor U18015 (N_18015,N_17288,N_17506);
nor U18016 (N_18016,N_17504,N_17183);
and U18017 (N_18017,N_17319,N_17841);
and U18018 (N_18018,N_17454,N_17425);
nand U18019 (N_18019,N_17516,N_17686);
or U18020 (N_18020,N_17565,N_17108);
or U18021 (N_18021,N_17572,N_17006);
xnor U18022 (N_18022,N_17374,N_17385);
and U18023 (N_18023,N_17154,N_17110);
or U18024 (N_18024,N_17519,N_17898);
xor U18025 (N_18025,N_17725,N_17963);
xnor U18026 (N_18026,N_17028,N_17178);
and U18027 (N_18027,N_17797,N_17266);
nand U18028 (N_18028,N_17250,N_17321);
or U18029 (N_18029,N_17705,N_17396);
and U18030 (N_18030,N_17689,N_17901);
nand U18031 (N_18031,N_17404,N_17851);
nor U18032 (N_18032,N_17625,N_17621);
nand U18033 (N_18033,N_17258,N_17105);
and U18034 (N_18034,N_17150,N_17534);
or U18035 (N_18035,N_17801,N_17121);
nand U18036 (N_18036,N_17302,N_17596);
xor U18037 (N_18037,N_17004,N_17791);
and U18038 (N_18038,N_17222,N_17790);
nor U18039 (N_18039,N_17094,N_17256);
nand U18040 (N_18040,N_17085,N_17612);
nor U18041 (N_18041,N_17556,N_17403);
and U18042 (N_18042,N_17915,N_17693);
nand U18043 (N_18043,N_17649,N_17280);
nor U18044 (N_18044,N_17091,N_17832);
xor U18045 (N_18045,N_17335,N_17058);
xnor U18046 (N_18046,N_17601,N_17977);
and U18047 (N_18047,N_17279,N_17249);
xor U18048 (N_18048,N_17914,N_17561);
or U18049 (N_18049,N_17918,N_17270);
and U18050 (N_18050,N_17162,N_17934);
nor U18051 (N_18051,N_17262,N_17694);
or U18052 (N_18052,N_17051,N_17439);
and U18053 (N_18053,N_17200,N_17084);
xnor U18054 (N_18054,N_17466,N_17517);
nand U18055 (N_18055,N_17940,N_17524);
or U18056 (N_18056,N_17124,N_17779);
nor U18057 (N_18057,N_17053,N_17584);
and U18058 (N_18058,N_17937,N_17985);
or U18059 (N_18059,N_17230,N_17599);
nor U18060 (N_18060,N_17752,N_17749);
and U18061 (N_18061,N_17254,N_17484);
nand U18062 (N_18062,N_17392,N_17549);
nand U18063 (N_18063,N_17669,N_17225);
or U18064 (N_18064,N_17278,N_17962);
or U18065 (N_18065,N_17113,N_17792);
nand U18066 (N_18066,N_17629,N_17630);
and U18067 (N_18067,N_17045,N_17957);
or U18068 (N_18068,N_17337,N_17718);
nor U18069 (N_18069,N_17386,N_17345);
nor U18070 (N_18070,N_17182,N_17435);
or U18071 (N_18071,N_17470,N_17858);
or U18072 (N_18072,N_17195,N_17646);
or U18073 (N_18073,N_17219,N_17798);
or U18074 (N_18074,N_17507,N_17023);
nor U18075 (N_18075,N_17925,N_17207);
nor U18076 (N_18076,N_17706,N_17933);
and U18077 (N_18077,N_17776,N_17164);
or U18078 (N_18078,N_17363,N_17981);
nand U18079 (N_18079,N_17034,N_17365);
xor U18080 (N_18080,N_17414,N_17037);
nand U18081 (N_18081,N_17447,N_17871);
xor U18082 (N_18082,N_17587,N_17734);
or U18083 (N_18083,N_17093,N_17632);
nor U18084 (N_18084,N_17515,N_17623);
xor U18085 (N_18085,N_17443,N_17078);
xnor U18086 (N_18086,N_17410,N_17188);
xnor U18087 (N_18087,N_17163,N_17911);
xnor U18088 (N_18088,N_17316,N_17635);
xnor U18089 (N_18089,N_17029,N_17009);
xor U18090 (N_18090,N_17213,N_17741);
and U18091 (N_18091,N_17203,N_17800);
nand U18092 (N_18092,N_17010,N_17943);
nand U18093 (N_18093,N_17438,N_17149);
xnor U18094 (N_18094,N_17532,N_17611);
nand U18095 (N_18095,N_17261,N_17833);
xnor U18096 (N_18096,N_17969,N_17950);
and U18097 (N_18097,N_17661,N_17910);
xor U18098 (N_18098,N_17186,N_17824);
or U18099 (N_18099,N_17952,N_17793);
nand U18100 (N_18100,N_17092,N_17882);
nand U18101 (N_18101,N_17300,N_17521);
or U18102 (N_18102,N_17684,N_17083);
or U18103 (N_18103,N_17936,N_17309);
xnor U18104 (N_18104,N_17433,N_17486);
nor U18105 (N_18105,N_17239,N_17756);
xnor U18106 (N_18106,N_17273,N_17112);
nand U18107 (N_18107,N_17274,N_17059);
nor U18108 (N_18108,N_17566,N_17780);
nor U18109 (N_18109,N_17986,N_17859);
and U18110 (N_18110,N_17628,N_17269);
xnor U18111 (N_18111,N_17732,N_17487);
or U18112 (N_18112,N_17807,N_17357);
nand U18113 (N_18113,N_17452,N_17054);
or U18114 (N_18114,N_17692,N_17451);
nor U18115 (N_18115,N_17930,N_17272);
or U18116 (N_18116,N_17971,N_17991);
xnor U18117 (N_18117,N_17238,N_17980);
and U18118 (N_18118,N_17724,N_17445);
and U18119 (N_18119,N_17458,N_17899);
and U18120 (N_18120,N_17146,N_17785);
and U18121 (N_18121,N_17227,N_17488);
or U18122 (N_18122,N_17232,N_17497);
and U18123 (N_18123,N_17430,N_17064);
xor U18124 (N_18124,N_17949,N_17248);
nor U18125 (N_18125,N_17554,N_17493);
nor U18126 (N_18126,N_17578,N_17420);
or U18127 (N_18127,N_17535,N_17241);
and U18128 (N_18128,N_17883,N_17573);
and U18129 (N_18129,N_17546,N_17842);
nand U18130 (N_18130,N_17398,N_17602);
nand U18131 (N_18131,N_17089,N_17804);
or U18132 (N_18132,N_17994,N_17953);
and U18133 (N_18133,N_17942,N_17772);
and U18134 (N_18134,N_17900,N_17234);
and U18135 (N_18135,N_17153,N_17904);
or U18136 (N_18136,N_17434,N_17728);
nor U18137 (N_18137,N_17555,N_17846);
and U18138 (N_18138,N_17831,N_17086);
nor U18139 (N_18139,N_17537,N_17614);
xnor U18140 (N_18140,N_17944,N_17464);
nand U18141 (N_18141,N_17680,N_17235);
or U18142 (N_18142,N_17654,N_17324);
or U18143 (N_18143,N_17326,N_17378);
or U18144 (N_18144,N_17559,N_17784);
nand U18145 (N_18145,N_17973,N_17066);
nor U18146 (N_18146,N_17591,N_17125);
or U18147 (N_18147,N_17191,N_17036);
xnor U18148 (N_18148,N_17929,N_17893);
xor U18149 (N_18149,N_17020,N_17039);
nand U18150 (N_18150,N_17140,N_17723);
xor U18151 (N_18151,N_17536,N_17197);
or U18152 (N_18152,N_17878,N_17165);
or U18153 (N_18153,N_17096,N_17827);
and U18154 (N_18154,N_17527,N_17212);
or U18155 (N_18155,N_17325,N_17312);
and U18156 (N_18156,N_17022,N_17283);
xnor U18157 (N_18157,N_17938,N_17617);
nand U18158 (N_18158,N_17716,N_17839);
nor U18159 (N_18159,N_17619,N_17127);
nor U18160 (N_18160,N_17017,N_17947);
nand U18161 (N_18161,N_17729,N_17173);
and U18162 (N_18162,N_17874,N_17627);
and U18163 (N_18163,N_17922,N_17012);
xor U18164 (N_18164,N_17463,N_17877);
nand U18165 (N_18165,N_17961,N_17913);
nand U18166 (N_18166,N_17301,N_17677);
xor U18167 (N_18167,N_17315,N_17525);
nor U18168 (N_18168,N_17416,N_17553);
nand U18169 (N_18169,N_17330,N_17364);
xor U18170 (N_18170,N_17354,N_17287);
nand U18171 (N_18171,N_17881,N_17989);
or U18172 (N_18172,N_17755,N_17067);
xnor U18173 (N_18173,N_17282,N_17655);
or U18174 (N_18174,N_17016,N_17286);
xor U18175 (N_18175,N_17820,N_17634);
xor U18176 (N_18176,N_17808,N_17215);
and U18177 (N_18177,N_17342,N_17129);
xnor U18178 (N_18178,N_17822,N_17490);
or U18179 (N_18179,N_17512,N_17926);
and U18180 (N_18180,N_17594,N_17424);
and U18181 (N_18181,N_17508,N_17708);
and U18182 (N_18182,N_17637,N_17277);
xor U18183 (N_18183,N_17794,N_17068);
and U18184 (N_18184,N_17581,N_17263);
xor U18185 (N_18185,N_17069,N_17640);
or U18186 (N_18186,N_17155,N_17123);
xnor U18187 (N_18187,N_17698,N_17401);
or U18188 (N_18188,N_17509,N_17742);
or U18189 (N_18189,N_17606,N_17769);
and U18190 (N_18190,N_17803,N_17551);
nand U18191 (N_18191,N_17823,N_17854);
or U18192 (N_18192,N_17079,N_17787);
nand U18193 (N_18193,N_17495,N_17855);
nor U18194 (N_18194,N_17848,N_17771);
or U18195 (N_18195,N_17082,N_17361);
and U18196 (N_18196,N_17528,N_17142);
nor U18197 (N_18197,N_17648,N_17193);
xnor U18198 (N_18198,N_17147,N_17131);
and U18199 (N_18199,N_17442,N_17117);
and U18200 (N_18200,N_17021,N_17715);
nand U18201 (N_18201,N_17428,N_17558);
nand U18202 (N_18202,N_17418,N_17838);
or U18203 (N_18203,N_17987,N_17025);
xnor U18204 (N_18204,N_17189,N_17429);
or U18205 (N_18205,N_17908,N_17690);
nor U18206 (N_18206,N_17008,N_17935);
or U18207 (N_18207,N_17002,N_17709);
nand U18208 (N_18208,N_17738,N_17688);
xnor U18209 (N_18209,N_17967,N_17620);
nand U18210 (N_18210,N_17449,N_17895);
nand U18211 (N_18211,N_17257,N_17687);
and U18212 (N_18212,N_17115,N_17358);
nor U18213 (N_18213,N_17691,N_17745);
xor U18214 (N_18214,N_17604,N_17329);
and U18215 (N_18215,N_17380,N_17003);
nand U18216 (N_18216,N_17931,N_17349);
nor U18217 (N_18217,N_17338,N_17607);
and U18218 (N_18218,N_17600,N_17879);
nor U18219 (N_18219,N_17662,N_17526);
and U18220 (N_18220,N_17144,N_17579);
or U18221 (N_18221,N_17367,N_17520);
or U18222 (N_18222,N_17886,N_17245);
nand U18223 (N_18223,N_17332,N_17633);
and U18224 (N_18224,N_17917,N_17339);
nand U18225 (N_18225,N_17647,N_17198);
nand U18226 (N_18226,N_17264,N_17436);
nor U18227 (N_18227,N_17641,N_17666);
or U18228 (N_18228,N_17141,N_17043);
xnor U18229 (N_18229,N_17701,N_17783);
and U18230 (N_18230,N_17869,N_17544);
or U18231 (N_18231,N_17597,N_17313);
and U18232 (N_18232,N_17668,N_17122);
xnor U18233 (N_18233,N_17076,N_17494);
nand U18234 (N_18234,N_17095,N_17097);
xnor U18235 (N_18235,N_17390,N_17446);
nor U18236 (N_18236,N_17158,N_17478);
nand U18237 (N_18237,N_17695,N_17441);
or U18238 (N_18238,N_17968,N_17626);
or U18239 (N_18239,N_17356,N_17765);
nor U18240 (N_18240,N_17906,N_17440);
or U18241 (N_18241,N_17202,N_17866);
nor U18242 (N_18242,N_17482,N_17460);
or U18243 (N_18243,N_17362,N_17897);
or U18244 (N_18244,N_17595,N_17956);
and U18245 (N_18245,N_17295,N_17618);
and U18246 (N_18246,N_17422,N_17829);
and U18247 (N_18247,N_17903,N_17575);
nor U18248 (N_18248,N_17861,N_17767);
and U18249 (N_18249,N_17727,N_17860);
or U18250 (N_18250,N_17642,N_17714);
nor U18251 (N_18251,N_17702,N_17975);
and U18252 (N_18252,N_17027,N_17624);
nand U18253 (N_18253,N_17169,N_17958);
nor U18254 (N_18254,N_17653,N_17498);
or U18255 (N_18255,N_17570,N_17387);
xor U18256 (N_18256,N_17291,N_17761);
nor U18257 (N_18257,N_17161,N_17214);
or U18258 (N_18258,N_17294,N_17360);
or U18259 (N_18259,N_17366,N_17622);
nor U18260 (N_18260,N_17699,N_17993);
and U18261 (N_18261,N_17444,N_17204);
nor U18262 (N_18262,N_17781,N_17795);
xor U18263 (N_18263,N_17340,N_17585);
nor U18264 (N_18264,N_17945,N_17685);
and U18265 (N_18265,N_17676,N_17032);
xnor U18266 (N_18266,N_17919,N_17696);
and U18267 (N_18267,N_17412,N_17799);
nor U18268 (N_18268,N_17737,N_17758);
xor U18269 (N_18269,N_17101,N_17306);
nor U18270 (N_18270,N_17821,N_17583);
xnor U18271 (N_18271,N_17061,N_17237);
nor U18272 (N_18272,N_17377,N_17181);
nor U18273 (N_18273,N_17087,N_17284);
or U18274 (N_18274,N_17176,N_17875);
and U18275 (N_18275,N_17015,N_17996);
and U18276 (N_18276,N_17166,N_17768);
nand U18277 (N_18277,N_17231,N_17334);
nor U18278 (N_18278,N_17501,N_17638);
and U18279 (N_18279,N_17921,N_17746);
xor U18280 (N_18280,N_17046,N_17305);
or U18281 (N_18281,N_17351,N_17529);
and U18282 (N_18282,N_17580,N_17133);
and U18283 (N_18283,N_17988,N_17011);
or U18284 (N_18284,N_17134,N_17373);
or U18285 (N_18285,N_17948,N_17151);
nand U18286 (N_18286,N_17598,N_17102);
nor U18287 (N_18287,N_17884,N_17159);
or U18288 (N_18288,N_17605,N_17719);
or U18289 (N_18289,N_17703,N_17001);
or U18290 (N_18290,N_17236,N_17090);
nand U18291 (N_18291,N_17786,N_17530);
nand U18292 (N_18292,N_17480,N_17109);
or U18293 (N_18293,N_17052,N_17965);
nand U18294 (N_18294,N_17639,N_17432);
nor U18295 (N_18295,N_17671,N_17397);
nor U18296 (N_18296,N_17609,N_17750);
nor U18297 (N_18297,N_17887,N_17156);
xnor U18298 (N_18298,N_17849,N_17588);
nor U18299 (N_18299,N_17383,N_17762);
and U18300 (N_18300,N_17782,N_17205);
nor U18301 (N_18301,N_17130,N_17311);
or U18302 (N_18302,N_17909,N_17187);
xnor U18303 (N_18303,N_17531,N_17834);
nor U18304 (N_18304,N_17050,N_17888);
and U18305 (N_18305,N_17700,N_17984);
and U18306 (N_18306,N_17116,N_17569);
nand U18307 (N_18307,N_17976,N_17244);
xor U18308 (N_18308,N_17491,N_17513);
nand U18309 (N_18309,N_17457,N_17468);
nand U18310 (N_18310,N_17119,N_17070);
and U18311 (N_18311,N_17242,N_17711);
nand U18312 (N_18312,N_17353,N_17348);
or U18313 (N_18313,N_17307,N_17522);
nand U18314 (N_18314,N_17243,N_17056);
xor U18315 (N_18315,N_17297,N_17160);
xor U18316 (N_18316,N_17099,N_17731);
nand U18317 (N_18317,N_17920,N_17577);
xor U18318 (N_18318,N_17114,N_17891);
and U18319 (N_18319,N_17643,N_17489);
nand U18320 (N_18320,N_17907,N_17928);
nand U18321 (N_18321,N_17582,N_17927);
xor U18322 (N_18322,N_17759,N_17548);
and U18323 (N_18323,N_17405,N_17845);
and U18324 (N_18324,N_17148,N_17409);
nor U18325 (N_18325,N_17813,N_17774);
nand U18326 (N_18326,N_17320,N_17000);
and U18327 (N_18327,N_17276,N_17175);
and U18328 (N_18328,N_17228,N_17932);
nand U18329 (N_18329,N_17744,N_17199);
xnor U18330 (N_18330,N_17865,N_17310);
nor U18331 (N_18331,N_17645,N_17479);
and U18332 (N_18332,N_17659,N_17168);
and U18333 (N_18333,N_17518,N_17304);
and U18334 (N_18334,N_17350,N_17812);
xor U18335 (N_18335,N_17568,N_17179);
nand U18336 (N_18336,N_17080,N_17343);
or U18337 (N_18337,N_17916,N_17024);
or U18338 (N_18338,N_17071,N_17788);
nand U18339 (N_18339,N_17376,N_17474);
nor U18340 (N_18340,N_17035,N_17657);
and U18341 (N_18341,N_17471,N_17802);
nor U18342 (N_18342,N_17152,N_17902);
and U18343 (N_18343,N_17816,N_17275);
nor U18344 (N_18344,N_17281,N_17352);
nor U18345 (N_18345,N_17636,N_17736);
xnor U18346 (N_18346,N_17103,N_17789);
xnor U18347 (N_18347,N_17955,N_17379);
or U18348 (N_18348,N_17062,N_17825);
nor U18349 (N_18349,N_17088,N_17892);
nand U18350 (N_18350,N_17293,N_17757);
nor U18351 (N_18351,N_17992,N_17044);
or U18352 (N_18352,N_17074,N_17978);
or U18353 (N_18353,N_17472,N_17206);
and U18354 (N_18354,N_17453,N_17815);
nand U18355 (N_18355,N_17562,N_17475);
nand U18356 (N_18356,N_17960,N_17394);
and U18357 (N_18357,N_17372,N_17658);
and U18358 (N_18358,N_17924,N_17201);
nor U18359 (N_18359,N_17533,N_17217);
xor U18360 (N_18360,N_17259,N_17145);
or U18361 (N_18361,N_17013,N_17857);
nor U18362 (N_18362,N_17055,N_17550);
xnor U18363 (N_18363,N_17682,N_17826);
nand U18364 (N_18364,N_17185,N_17672);
xnor U18365 (N_18365,N_17042,N_17292);
xor U18366 (N_18366,N_17972,N_17072);
nand U18367 (N_18367,N_17836,N_17754);
xor U18368 (N_18368,N_17941,N_17722);
nor U18369 (N_18369,N_17448,N_17964);
or U18370 (N_18370,N_17697,N_17308);
nor U18371 (N_18371,N_17844,N_17346);
nand U18372 (N_18372,N_17862,N_17511);
xnor U18373 (N_18373,N_17406,N_17065);
nor U18374 (N_18374,N_17048,N_17819);
xnor U18375 (N_18375,N_17031,N_17835);
nor U18376 (N_18376,N_17979,N_17171);
nor U18377 (N_18377,N_17660,N_17328);
and U18378 (N_18378,N_17426,N_17999);
and U18379 (N_18379,N_17450,N_17650);
xnor U18380 (N_18380,N_17740,N_17375);
nand U18381 (N_18381,N_17959,N_17564);
nor U18382 (N_18382,N_17223,N_17733);
nand U18383 (N_18383,N_17856,N_17111);
nor U18384 (N_18384,N_17775,N_17995);
and U18385 (N_18385,N_17407,N_17603);
nand U18386 (N_18386,N_17251,N_17384);
and U18387 (N_18387,N_17500,N_17492);
nor U18388 (N_18388,N_17411,N_17665);
xor U18389 (N_18389,N_17211,N_17382);
and U18390 (N_18390,N_17743,N_17853);
nand U18391 (N_18391,N_17018,N_17077);
nand U18392 (N_18392,N_17388,N_17208);
nand U18393 (N_18393,N_17030,N_17905);
xnor U18394 (N_18394,N_17608,N_17864);
or U18395 (N_18395,N_17717,N_17260);
nand U18396 (N_18396,N_17196,N_17408);
or U18397 (N_18397,N_17100,N_17773);
xor U18398 (N_18398,N_17210,N_17563);
and U18399 (N_18399,N_17423,N_17098);
xor U18400 (N_18400,N_17852,N_17610);
or U18401 (N_18401,N_17370,N_17104);
nor U18402 (N_18402,N_17184,N_17341);
xor U18403 (N_18403,N_17644,N_17766);
nand U18404 (N_18404,N_17303,N_17298);
or U18405 (N_18405,N_17721,N_17106);
nand U18406 (N_18406,N_17355,N_17557);
or U18407 (N_18407,N_17253,N_17730);
and U18408 (N_18408,N_17867,N_17007);
nor U18409 (N_18409,N_17126,N_17889);
and U18410 (N_18410,N_17229,N_17437);
or U18411 (N_18411,N_17651,N_17267);
and U18412 (N_18412,N_17847,N_17393);
or U18413 (N_18413,N_17510,N_17136);
xor U18414 (N_18414,N_17514,N_17760);
nand U18415 (N_18415,N_17499,N_17763);
or U18416 (N_18416,N_17811,N_17710);
xnor U18417 (N_18417,N_17966,N_17167);
nand U18418 (N_18418,N_17983,N_17413);
xnor U18419 (N_18419,N_17539,N_17545);
nand U18420 (N_18420,N_17224,N_17040);
nor U18421 (N_18421,N_17974,N_17574);
and U18422 (N_18422,N_17485,N_17026);
and U18423 (N_18423,N_17391,N_17369);
xor U18424 (N_18424,N_17496,N_17190);
or U18425 (N_18425,N_17246,N_17139);
xor U18426 (N_18426,N_17057,N_17336);
xnor U18427 (N_18427,N_17047,N_17828);
or U18428 (N_18428,N_17778,N_17523);
xnor U18429 (N_18429,N_17753,N_17840);
or U18430 (N_18430,N_17589,N_17194);
nor U18431 (N_18431,N_17667,N_17268);
or U18432 (N_18432,N_17415,N_17299);
xor U18433 (N_18433,N_17664,N_17997);
and U18434 (N_18434,N_17255,N_17467);
xor U18435 (N_18435,N_17247,N_17371);
nor U18436 (N_18436,N_17417,N_17896);
and U18437 (N_18437,N_17982,N_17322);
nand U18438 (N_18438,N_17567,N_17233);
xnor U18439 (N_18439,N_17590,N_17873);
xnor U18440 (N_18440,N_17720,N_17770);
and U18441 (N_18441,N_17192,N_17713);
xor U18442 (N_18442,N_17033,N_17177);
nand U18443 (N_18443,N_17389,N_17837);
and U18444 (N_18444,N_17613,N_17049);
xnor U18445 (N_18445,N_17970,N_17751);
nand U18446 (N_18446,N_17586,N_17400);
nand U18447 (N_18447,N_17483,N_17323);
nand U18448 (N_18448,N_17885,N_17041);
or U18449 (N_18449,N_17359,N_17265);
xor U18450 (N_18450,N_17890,N_17395);
nand U18451 (N_18451,N_17764,N_17455);
and U18452 (N_18452,N_17704,N_17285);
nand U18453 (N_18453,N_17135,N_17998);
nand U18454 (N_18454,N_17473,N_17850);
nand U18455 (N_18455,N_17538,N_17314);
nand U18456 (N_18456,N_17663,N_17817);
nor U18457 (N_18457,N_17465,N_17209);
or U18458 (N_18458,N_17075,N_17540);
nor U18459 (N_18459,N_17317,N_17576);
or U18460 (N_18460,N_17289,N_17063);
and U18461 (N_18461,N_17592,N_17431);
nand U18462 (N_18462,N_17128,N_17615);
xnor U18463 (N_18463,N_17954,N_17469);
xnor U18464 (N_18464,N_17456,N_17240);
nor U18465 (N_18465,N_17543,N_17038);
nand U18466 (N_18466,N_17796,N_17333);
nor U18467 (N_18467,N_17296,N_17318);
and U18468 (N_18468,N_17726,N_17132);
or U18469 (N_18469,N_17678,N_17560);
nand U18470 (N_18470,N_17748,N_17481);
nor U18471 (N_18471,N_17459,N_17939);
nand U18472 (N_18472,N_17172,N_17107);
nor U18473 (N_18473,N_17673,N_17675);
nor U18474 (N_18474,N_17138,N_17868);
nand U18475 (N_18475,N_17923,N_17462);
nor U18476 (N_18476,N_17344,N_17180);
nand U18477 (N_18477,N_17674,N_17571);
nand U18478 (N_18478,N_17541,N_17652);
or U18479 (N_18479,N_17477,N_17990);
xor U18480 (N_18480,N_17946,N_17912);
xor U18481 (N_18481,N_17381,N_17747);
xor U18482 (N_18482,N_17670,N_17157);
and U18483 (N_18483,N_17872,N_17019);
or U18484 (N_18484,N_17331,N_17118);
xor U18485 (N_18485,N_17805,N_17120);
and U18486 (N_18486,N_17476,N_17542);
nand U18487 (N_18487,N_17547,N_17368);
xor U18488 (N_18488,N_17014,N_17503);
xnor U18489 (N_18489,N_17830,N_17777);
nor U18490 (N_18490,N_17814,N_17060);
nand U18491 (N_18491,N_17809,N_17552);
and U18492 (N_18492,N_17712,N_17402);
or U18493 (N_18493,N_17656,N_17593);
nand U18494 (N_18494,N_17505,N_17421);
or U18495 (N_18495,N_17951,N_17081);
or U18496 (N_18496,N_17347,N_17880);
nand U18497 (N_18497,N_17735,N_17679);
or U18498 (N_18498,N_17894,N_17218);
and U18499 (N_18499,N_17427,N_17143);
and U18500 (N_18500,N_17110,N_17081);
xor U18501 (N_18501,N_17193,N_17476);
nor U18502 (N_18502,N_17522,N_17219);
nand U18503 (N_18503,N_17345,N_17012);
nor U18504 (N_18504,N_17788,N_17294);
nand U18505 (N_18505,N_17188,N_17286);
nor U18506 (N_18506,N_17884,N_17158);
or U18507 (N_18507,N_17484,N_17892);
and U18508 (N_18508,N_17554,N_17583);
nand U18509 (N_18509,N_17802,N_17248);
nand U18510 (N_18510,N_17489,N_17819);
nor U18511 (N_18511,N_17977,N_17966);
nand U18512 (N_18512,N_17829,N_17208);
xnor U18513 (N_18513,N_17319,N_17232);
or U18514 (N_18514,N_17866,N_17681);
or U18515 (N_18515,N_17619,N_17568);
and U18516 (N_18516,N_17871,N_17996);
nor U18517 (N_18517,N_17092,N_17810);
nor U18518 (N_18518,N_17967,N_17297);
xnor U18519 (N_18519,N_17657,N_17951);
or U18520 (N_18520,N_17128,N_17838);
nor U18521 (N_18521,N_17566,N_17183);
and U18522 (N_18522,N_17817,N_17753);
nor U18523 (N_18523,N_17291,N_17860);
nor U18524 (N_18524,N_17769,N_17786);
or U18525 (N_18525,N_17608,N_17471);
nor U18526 (N_18526,N_17037,N_17509);
and U18527 (N_18527,N_17980,N_17621);
nor U18528 (N_18528,N_17282,N_17323);
nand U18529 (N_18529,N_17472,N_17034);
nor U18530 (N_18530,N_17388,N_17884);
nor U18531 (N_18531,N_17158,N_17275);
nand U18532 (N_18532,N_17927,N_17038);
nand U18533 (N_18533,N_17157,N_17253);
nor U18534 (N_18534,N_17417,N_17864);
and U18535 (N_18535,N_17579,N_17541);
nor U18536 (N_18536,N_17487,N_17070);
xnor U18537 (N_18537,N_17093,N_17408);
nand U18538 (N_18538,N_17596,N_17252);
nor U18539 (N_18539,N_17603,N_17282);
or U18540 (N_18540,N_17681,N_17648);
and U18541 (N_18541,N_17673,N_17658);
or U18542 (N_18542,N_17512,N_17675);
or U18543 (N_18543,N_17615,N_17675);
nand U18544 (N_18544,N_17045,N_17518);
nor U18545 (N_18545,N_17066,N_17341);
or U18546 (N_18546,N_17452,N_17323);
nand U18547 (N_18547,N_17001,N_17288);
nand U18548 (N_18548,N_17986,N_17076);
or U18549 (N_18549,N_17847,N_17690);
nand U18550 (N_18550,N_17057,N_17490);
and U18551 (N_18551,N_17249,N_17429);
nand U18552 (N_18552,N_17857,N_17581);
xnor U18553 (N_18553,N_17459,N_17616);
nor U18554 (N_18554,N_17515,N_17777);
or U18555 (N_18555,N_17202,N_17134);
or U18556 (N_18556,N_17335,N_17498);
and U18557 (N_18557,N_17732,N_17837);
nor U18558 (N_18558,N_17720,N_17960);
and U18559 (N_18559,N_17394,N_17169);
or U18560 (N_18560,N_17921,N_17975);
and U18561 (N_18561,N_17729,N_17949);
or U18562 (N_18562,N_17488,N_17180);
nand U18563 (N_18563,N_17453,N_17606);
xor U18564 (N_18564,N_17337,N_17110);
nand U18565 (N_18565,N_17181,N_17908);
and U18566 (N_18566,N_17351,N_17554);
nand U18567 (N_18567,N_17018,N_17950);
nand U18568 (N_18568,N_17231,N_17970);
or U18569 (N_18569,N_17452,N_17868);
or U18570 (N_18570,N_17433,N_17095);
or U18571 (N_18571,N_17198,N_17235);
or U18572 (N_18572,N_17238,N_17863);
and U18573 (N_18573,N_17051,N_17109);
nand U18574 (N_18574,N_17906,N_17913);
xnor U18575 (N_18575,N_17477,N_17431);
or U18576 (N_18576,N_17233,N_17495);
and U18577 (N_18577,N_17933,N_17183);
nor U18578 (N_18578,N_17809,N_17037);
and U18579 (N_18579,N_17798,N_17008);
nand U18580 (N_18580,N_17506,N_17355);
or U18581 (N_18581,N_17885,N_17405);
and U18582 (N_18582,N_17299,N_17144);
nor U18583 (N_18583,N_17783,N_17798);
or U18584 (N_18584,N_17430,N_17985);
and U18585 (N_18585,N_17088,N_17632);
and U18586 (N_18586,N_17773,N_17537);
nor U18587 (N_18587,N_17905,N_17431);
or U18588 (N_18588,N_17775,N_17781);
and U18589 (N_18589,N_17053,N_17028);
or U18590 (N_18590,N_17597,N_17232);
xnor U18591 (N_18591,N_17069,N_17394);
nand U18592 (N_18592,N_17081,N_17754);
nand U18593 (N_18593,N_17516,N_17224);
or U18594 (N_18594,N_17737,N_17657);
and U18595 (N_18595,N_17505,N_17017);
xor U18596 (N_18596,N_17085,N_17773);
nand U18597 (N_18597,N_17661,N_17850);
and U18598 (N_18598,N_17352,N_17233);
xor U18599 (N_18599,N_17947,N_17230);
nor U18600 (N_18600,N_17183,N_17690);
xor U18601 (N_18601,N_17691,N_17088);
xnor U18602 (N_18602,N_17754,N_17011);
nand U18603 (N_18603,N_17599,N_17837);
and U18604 (N_18604,N_17961,N_17726);
nor U18605 (N_18605,N_17628,N_17479);
and U18606 (N_18606,N_17365,N_17122);
xor U18607 (N_18607,N_17493,N_17927);
or U18608 (N_18608,N_17490,N_17819);
or U18609 (N_18609,N_17677,N_17947);
and U18610 (N_18610,N_17613,N_17283);
xnor U18611 (N_18611,N_17645,N_17309);
or U18612 (N_18612,N_17377,N_17303);
and U18613 (N_18613,N_17114,N_17870);
and U18614 (N_18614,N_17484,N_17552);
xor U18615 (N_18615,N_17526,N_17784);
nand U18616 (N_18616,N_17776,N_17397);
and U18617 (N_18617,N_17042,N_17642);
nand U18618 (N_18618,N_17376,N_17978);
or U18619 (N_18619,N_17832,N_17864);
nor U18620 (N_18620,N_17920,N_17038);
xnor U18621 (N_18621,N_17415,N_17927);
nand U18622 (N_18622,N_17240,N_17198);
nor U18623 (N_18623,N_17797,N_17062);
and U18624 (N_18624,N_17857,N_17237);
nand U18625 (N_18625,N_17168,N_17899);
nor U18626 (N_18626,N_17289,N_17306);
xnor U18627 (N_18627,N_17679,N_17372);
xor U18628 (N_18628,N_17557,N_17793);
nor U18629 (N_18629,N_17798,N_17452);
xor U18630 (N_18630,N_17254,N_17073);
and U18631 (N_18631,N_17683,N_17507);
and U18632 (N_18632,N_17106,N_17037);
and U18633 (N_18633,N_17011,N_17422);
xor U18634 (N_18634,N_17696,N_17707);
xor U18635 (N_18635,N_17829,N_17047);
nand U18636 (N_18636,N_17416,N_17825);
nor U18637 (N_18637,N_17142,N_17839);
and U18638 (N_18638,N_17577,N_17459);
or U18639 (N_18639,N_17761,N_17135);
nor U18640 (N_18640,N_17017,N_17704);
nand U18641 (N_18641,N_17647,N_17965);
and U18642 (N_18642,N_17666,N_17456);
and U18643 (N_18643,N_17294,N_17009);
nand U18644 (N_18644,N_17897,N_17272);
xor U18645 (N_18645,N_17895,N_17521);
and U18646 (N_18646,N_17327,N_17465);
nor U18647 (N_18647,N_17226,N_17739);
nand U18648 (N_18648,N_17454,N_17311);
nor U18649 (N_18649,N_17456,N_17255);
or U18650 (N_18650,N_17097,N_17454);
nand U18651 (N_18651,N_17995,N_17361);
xor U18652 (N_18652,N_17783,N_17852);
or U18653 (N_18653,N_17257,N_17173);
nor U18654 (N_18654,N_17675,N_17411);
and U18655 (N_18655,N_17859,N_17079);
nand U18656 (N_18656,N_17103,N_17599);
xor U18657 (N_18657,N_17536,N_17266);
or U18658 (N_18658,N_17367,N_17564);
nand U18659 (N_18659,N_17878,N_17550);
and U18660 (N_18660,N_17624,N_17236);
xor U18661 (N_18661,N_17723,N_17993);
or U18662 (N_18662,N_17260,N_17032);
nand U18663 (N_18663,N_17865,N_17147);
nor U18664 (N_18664,N_17112,N_17340);
nand U18665 (N_18665,N_17815,N_17049);
nor U18666 (N_18666,N_17015,N_17754);
or U18667 (N_18667,N_17335,N_17635);
or U18668 (N_18668,N_17261,N_17119);
nand U18669 (N_18669,N_17089,N_17279);
xnor U18670 (N_18670,N_17624,N_17240);
and U18671 (N_18671,N_17822,N_17593);
nand U18672 (N_18672,N_17032,N_17137);
or U18673 (N_18673,N_17696,N_17490);
nor U18674 (N_18674,N_17827,N_17442);
and U18675 (N_18675,N_17500,N_17202);
nor U18676 (N_18676,N_17027,N_17901);
xnor U18677 (N_18677,N_17677,N_17273);
xnor U18678 (N_18678,N_17006,N_17425);
nand U18679 (N_18679,N_17493,N_17028);
and U18680 (N_18680,N_17090,N_17797);
or U18681 (N_18681,N_17250,N_17795);
nor U18682 (N_18682,N_17009,N_17383);
nand U18683 (N_18683,N_17334,N_17061);
xor U18684 (N_18684,N_17799,N_17903);
and U18685 (N_18685,N_17796,N_17659);
xnor U18686 (N_18686,N_17826,N_17081);
or U18687 (N_18687,N_17294,N_17957);
nor U18688 (N_18688,N_17491,N_17831);
and U18689 (N_18689,N_17296,N_17300);
or U18690 (N_18690,N_17818,N_17018);
and U18691 (N_18691,N_17878,N_17108);
and U18692 (N_18692,N_17903,N_17560);
nand U18693 (N_18693,N_17719,N_17057);
nor U18694 (N_18694,N_17041,N_17468);
or U18695 (N_18695,N_17035,N_17492);
and U18696 (N_18696,N_17738,N_17515);
nand U18697 (N_18697,N_17225,N_17903);
and U18698 (N_18698,N_17446,N_17332);
nand U18699 (N_18699,N_17082,N_17569);
xor U18700 (N_18700,N_17321,N_17295);
nor U18701 (N_18701,N_17422,N_17824);
nor U18702 (N_18702,N_17339,N_17005);
xor U18703 (N_18703,N_17472,N_17748);
nor U18704 (N_18704,N_17317,N_17701);
or U18705 (N_18705,N_17782,N_17555);
xor U18706 (N_18706,N_17619,N_17564);
and U18707 (N_18707,N_17648,N_17258);
and U18708 (N_18708,N_17975,N_17509);
nor U18709 (N_18709,N_17897,N_17254);
or U18710 (N_18710,N_17966,N_17169);
or U18711 (N_18711,N_17164,N_17017);
nor U18712 (N_18712,N_17881,N_17715);
or U18713 (N_18713,N_17498,N_17190);
nand U18714 (N_18714,N_17153,N_17266);
or U18715 (N_18715,N_17413,N_17870);
and U18716 (N_18716,N_17604,N_17261);
xor U18717 (N_18717,N_17483,N_17518);
xor U18718 (N_18718,N_17628,N_17255);
nand U18719 (N_18719,N_17028,N_17943);
nand U18720 (N_18720,N_17149,N_17758);
xnor U18721 (N_18721,N_17798,N_17794);
nand U18722 (N_18722,N_17831,N_17275);
or U18723 (N_18723,N_17015,N_17803);
or U18724 (N_18724,N_17554,N_17440);
and U18725 (N_18725,N_17405,N_17469);
nor U18726 (N_18726,N_17576,N_17010);
nand U18727 (N_18727,N_17864,N_17743);
nor U18728 (N_18728,N_17561,N_17777);
nand U18729 (N_18729,N_17350,N_17664);
nand U18730 (N_18730,N_17874,N_17770);
and U18731 (N_18731,N_17017,N_17988);
nand U18732 (N_18732,N_17361,N_17278);
nand U18733 (N_18733,N_17046,N_17641);
nand U18734 (N_18734,N_17112,N_17428);
xor U18735 (N_18735,N_17226,N_17960);
and U18736 (N_18736,N_17280,N_17663);
nor U18737 (N_18737,N_17308,N_17258);
xnor U18738 (N_18738,N_17286,N_17468);
and U18739 (N_18739,N_17339,N_17974);
nor U18740 (N_18740,N_17498,N_17766);
xor U18741 (N_18741,N_17716,N_17295);
xor U18742 (N_18742,N_17774,N_17246);
xor U18743 (N_18743,N_17502,N_17091);
nand U18744 (N_18744,N_17755,N_17219);
nand U18745 (N_18745,N_17812,N_17936);
or U18746 (N_18746,N_17695,N_17995);
and U18747 (N_18747,N_17754,N_17974);
nand U18748 (N_18748,N_17904,N_17167);
or U18749 (N_18749,N_17572,N_17299);
or U18750 (N_18750,N_17450,N_17694);
nor U18751 (N_18751,N_17968,N_17254);
or U18752 (N_18752,N_17377,N_17193);
and U18753 (N_18753,N_17736,N_17312);
nand U18754 (N_18754,N_17548,N_17589);
xnor U18755 (N_18755,N_17833,N_17841);
or U18756 (N_18756,N_17453,N_17491);
and U18757 (N_18757,N_17684,N_17757);
or U18758 (N_18758,N_17379,N_17160);
or U18759 (N_18759,N_17252,N_17436);
or U18760 (N_18760,N_17912,N_17368);
xnor U18761 (N_18761,N_17171,N_17958);
and U18762 (N_18762,N_17317,N_17201);
xnor U18763 (N_18763,N_17038,N_17402);
and U18764 (N_18764,N_17182,N_17217);
nand U18765 (N_18765,N_17707,N_17249);
and U18766 (N_18766,N_17295,N_17820);
and U18767 (N_18767,N_17487,N_17406);
xnor U18768 (N_18768,N_17500,N_17055);
or U18769 (N_18769,N_17177,N_17476);
nor U18770 (N_18770,N_17813,N_17108);
or U18771 (N_18771,N_17546,N_17861);
or U18772 (N_18772,N_17854,N_17900);
nor U18773 (N_18773,N_17305,N_17819);
nand U18774 (N_18774,N_17186,N_17455);
or U18775 (N_18775,N_17756,N_17042);
xor U18776 (N_18776,N_17802,N_17540);
and U18777 (N_18777,N_17807,N_17643);
and U18778 (N_18778,N_17343,N_17671);
xor U18779 (N_18779,N_17767,N_17456);
and U18780 (N_18780,N_17485,N_17532);
nor U18781 (N_18781,N_17821,N_17658);
xnor U18782 (N_18782,N_17661,N_17567);
xor U18783 (N_18783,N_17739,N_17095);
and U18784 (N_18784,N_17274,N_17454);
nor U18785 (N_18785,N_17957,N_17394);
nor U18786 (N_18786,N_17308,N_17266);
nor U18787 (N_18787,N_17888,N_17157);
and U18788 (N_18788,N_17249,N_17360);
nand U18789 (N_18789,N_17341,N_17672);
nor U18790 (N_18790,N_17702,N_17718);
and U18791 (N_18791,N_17669,N_17654);
or U18792 (N_18792,N_17563,N_17847);
and U18793 (N_18793,N_17706,N_17458);
nand U18794 (N_18794,N_17436,N_17656);
nor U18795 (N_18795,N_17323,N_17291);
nor U18796 (N_18796,N_17617,N_17657);
xnor U18797 (N_18797,N_17945,N_17850);
and U18798 (N_18798,N_17546,N_17370);
nand U18799 (N_18799,N_17969,N_17112);
xnor U18800 (N_18800,N_17091,N_17416);
nand U18801 (N_18801,N_17154,N_17397);
and U18802 (N_18802,N_17826,N_17058);
nand U18803 (N_18803,N_17639,N_17816);
xnor U18804 (N_18804,N_17834,N_17074);
nand U18805 (N_18805,N_17720,N_17840);
or U18806 (N_18806,N_17165,N_17159);
nand U18807 (N_18807,N_17480,N_17558);
and U18808 (N_18808,N_17108,N_17900);
nor U18809 (N_18809,N_17528,N_17503);
nand U18810 (N_18810,N_17761,N_17467);
nor U18811 (N_18811,N_17840,N_17668);
xor U18812 (N_18812,N_17140,N_17004);
xnor U18813 (N_18813,N_17364,N_17913);
and U18814 (N_18814,N_17345,N_17681);
and U18815 (N_18815,N_17693,N_17337);
xnor U18816 (N_18816,N_17833,N_17120);
or U18817 (N_18817,N_17853,N_17892);
nor U18818 (N_18818,N_17784,N_17192);
or U18819 (N_18819,N_17449,N_17046);
or U18820 (N_18820,N_17736,N_17233);
xnor U18821 (N_18821,N_17744,N_17241);
and U18822 (N_18822,N_17365,N_17863);
or U18823 (N_18823,N_17751,N_17146);
and U18824 (N_18824,N_17689,N_17548);
xor U18825 (N_18825,N_17867,N_17381);
nand U18826 (N_18826,N_17131,N_17053);
or U18827 (N_18827,N_17862,N_17004);
nor U18828 (N_18828,N_17611,N_17538);
nand U18829 (N_18829,N_17496,N_17935);
xor U18830 (N_18830,N_17039,N_17128);
or U18831 (N_18831,N_17038,N_17707);
nor U18832 (N_18832,N_17648,N_17989);
nor U18833 (N_18833,N_17254,N_17428);
or U18834 (N_18834,N_17446,N_17780);
xnor U18835 (N_18835,N_17122,N_17688);
nor U18836 (N_18836,N_17347,N_17728);
nand U18837 (N_18837,N_17002,N_17645);
nand U18838 (N_18838,N_17519,N_17066);
xor U18839 (N_18839,N_17074,N_17704);
nand U18840 (N_18840,N_17075,N_17656);
xnor U18841 (N_18841,N_17366,N_17617);
or U18842 (N_18842,N_17076,N_17685);
or U18843 (N_18843,N_17242,N_17108);
and U18844 (N_18844,N_17055,N_17150);
and U18845 (N_18845,N_17458,N_17821);
or U18846 (N_18846,N_17964,N_17380);
and U18847 (N_18847,N_17288,N_17500);
nor U18848 (N_18848,N_17862,N_17412);
xnor U18849 (N_18849,N_17319,N_17825);
xor U18850 (N_18850,N_17271,N_17494);
xnor U18851 (N_18851,N_17351,N_17520);
and U18852 (N_18852,N_17578,N_17706);
nand U18853 (N_18853,N_17079,N_17936);
xor U18854 (N_18854,N_17081,N_17678);
nand U18855 (N_18855,N_17867,N_17109);
nand U18856 (N_18856,N_17174,N_17830);
nor U18857 (N_18857,N_17487,N_17606);
nor U18858 (N_18858,N_17689,N_17713);
nand U18859 (N_18859,N_17852,N_17493);
xnor U18860 (N_18860,N_17855,N_17569);
or U18861 (N_18861,N_17734,N_17946);
or U18862 (N_18862,N_17841,N_17272);
or U18863 (N_18863,N_17452,N_17222);
and U18864 (N_18864,N_17722,N_17795);
nand U18865 (N_18865,N_17169,N_17611);
or U18866 (N_18866,N_17839,N_17786);
nand U18867 (N_18867,N_17104,N_17525);
or U18868 (N_18868,N_17380,N_17928);
xnor U18869 (N_18869,N_17488,N_17125);
xor U18870 (N_18870,N_17518,N_17116);
xnor U18871 (N_18871,N_17746,N_17494);
and U18872 (N_18872,N_17417,N_17418);
nand U18873 (N_18873,N_17578,N_17313);
nand U18874 (N_18874,N_17732,N_17933);
or U18875 (N_18875,N_17993,N_17930);
and U18876 (N_18876,N_17120,N_17188);
and U18877 (N_18877,N_17318,N_17362);
nand U18878 (N_18878,N_17089,N_17021);
xnor U18879 (N_18879,N_17317,N_17497);
and U18880 (N_18880,N_17886,N_17202);
nor U18881 (N_18881,N_17693,N_17381);
and U18882 (N_18882,N_17226,N_17157);
xnor U18883 (N_18883,N_17763,N_17077);
nor U18884 (N_18884,N_17981,N_17023);
nand U18885 (N_18885,N_17783,N_17723);
xor U18886 (N_18886,N_17312,N_17902);
nand U18887 (N_18887,N_17463,N_17375);
and U18888 (N_18888,N_17621,N_17971);
xor U18889 (N_18889,N_17882,N_17258);
or U18890 (N_18890,N_17511,N_17496);
and U18891 (N_18891,N_17035,N_17063);
nor U18892 (N_18892,N_17779,N_17984);
xor U18893 (N_18893,N_17928,N_17599);
nor U18894 (N_18894,N_17924,N_17846);
or U18895 (N_18895,N_17510,N_17461);
xnor U18896 (N_18896,N_17808,N_17444);
nand U18897 (N_18897,N_17631,N_17156);
or U18898 (N_18898,N_17933,N_17858);
and U18899 (N_18899,N_17392,N_17038);
xor U18900 (N_18900,N_17081,N_17922);
or U18901 (N_18901,N_17617,N_17028);
nor U18902 (N_18902,N_17764,N_17296);
nor U18903 (N_18903,N_17220,N_17981);
and U18904 (N_18904,N_17356,N_17163);
nor U18905 (N_18905,N_17067,N_17554);
nand U18906 (N_18906,N_17187,N_17386);
nand U18907 (N_18907,N_17641,N_17644);
nand U18908 (N_18908,N_17027,N_17411);
or U18909 (N_18909,N_17563,N_17403);
nor U18910 (N_18910,N_17186,N_17233);
nand U18911 (N_18911,N_17719,N_17991);
nand U18912 (N_18912,N_17937,N_17808);
and U18913 (N_18913,N_17556,N_17357);
nand U18914 (N_18914,N_17042,N_17964);
nor U18915 (N_18915,N_17392,N_17582);
nand U18916 (N_18916,N_17114,N_17811);
nor U18917 (N_18917,N_17768,N_17347);
and U18918 (N_18918,N_17788,N_17957);
nand U18919 (N_18919,N_17605,N_17442);
nor U18920 (N_18920,N_17964,N_17426);
xnor U18921 (N_18921,N_17974,N_17119);
or U18922 (N_18922,N_17200,N_17157);
xor U18923 (N_18923,N_17411,N_17431);
and U18924 (N_18924,N_17354,N_17826);
xnor U18925 (N_18925,N_17619,N_17332);
nor U18926 (N_18926,N_17983,N_17145);
nand U18927 (N_18927,N_17056,N_17973);
nand U18928 (N_18928,N_17600,N_17886);
and U18929 (N_18929,N_17138,N_17030);
and U18930 (N_18930,N_17438,N_17600);
nand U18931 (N_18931,N_17373,N_17322);
and U18932 (N_18932,N_17866,N_17754);
xnor U18933 (N_18933,N_17327,N_17684);
nand U18934 (N_18934,N_17668,N_17833);
nand U18935 (N_18935,N_17210,N_17679);
and U18936 (N_18936,N_17514,N_17291);
xor U18937 (N_18937,N_17747,N_17610);
nor U18938 (N_18938,N_17763,N_17571);
nor U18939 (N_18939,N_17202,N_17620);
or U18940 (N_18940,N_17703,N_17654);
nor U18941 (N_18941,N_17398,N_17765);
xor U18942 (N_18942,N_17499,N_17851);
xnor U18943 (N_18943,N_17857,N_17824);
and U18944 (N_18944,N_17791,N_17237);
nand U18945 (N_18945,N_17489,N_17003);
nand U18946 (N_18946,N_17403,N_17148);
or U18947 (N_18947,N_17778,N_17777);
xnor U18948 (N_18948,N_17977,N_17378);
nand U18949 (N_18949,N_17538,N_17641);
or U18950 (N_18950,N_17995,N_17387);
nand U18951 (N_18951,N_17041,N_17676);
or U18952 (N_18952,N_17704,N_17366);
xor U18953 (N_18953,N_17870,N_17184);
or U18954 (N_18954,N_17087,N_17189);
xnor U18955 (N_18955,N_17207,N_17571);
nor U18956 (N_18956,N_17899,N_17923);
or U18957 (N_18957,N_17490,N_17478);
nor U18958 (N_18958,N_17806,N_17699);
nor U18959 (N_18959,N_17223,N_17697);
xor U18960 (N_18960,N_17453,N_17154);
nor U18961 (N_18961,N_17273,N_17808);
or U18962 (N_18962,N_17497,N_17815);
nor U18963 (N_18963,N_17437,N_17467);
xnor U18964 (N_18964,N_17300,N_17156);
nand U18965 (N_18965,N_17474,N_17745);
or U18966 (N_18966,N_17060,N_17079);
or U18967 (N_18967,N_17197,N_17173);
nor U18968 (N_18968,N_17395,N_17490);
nor U18969 (N_18969,N_17769,N_17584);
xor U18970 (N_18970,N_17051,N_17412);
nor U18971 (N_18971,N_17381,N_17640);
nand U18972 (N_18972,N_17302,N_17485);
nand U18973 (N_18973,N_17427,N_17137);
or U18974 (N_18974,N_17586,N_17348);
or U18975 (N_18975,N_17600,N_17213);
and U18976 (N_18976,N_17073,N_17344);
nand U18977 (N_18977,N_17761,N_17155);
or U18978 (N_18978,N_17833,N_17907);
or U18979 (N_18979,N_17040,N_17394);
nand U18980 (N_18980,N_17470,N_17274);
nand U18981 (N_18981,N_17045,N_17482);
nand U18982 (N_18982,N_17532,N_17388);
nor U18983 (N_18983,N_17656,N_17108);
xor U18984 (N_18984,N_17539,N_17110);
or U18985 (N_18985,N_17439,N_17731);
or U18986 (N_18986,N_17075,N_17699);
xor U18987 (N_18987,N_17323,N_17290);
nand U18988 (N_18988,N_17685,N_17124);
nand U18989 (N_18989,N_17318,N_17655);
nor U18990 (N_18990,N_17652,N_17292);
or U18991 (N_18991,N_17065,N_17397);
and U18992 (N_18992,N_17076,N_17936);
nand U18993 (N_18993,N_17239,N_17463);
and U18994 (N_18994,N_17407,N_17769);
xnor U18995 (N_18995,N_17148,N_17464);
xnor U18996 (N_18996,N_17256,N_17905);
and U18997 (N_18997,N_17448,N_17048);
nor U18998 (N_18998,N_17465,N_17818);
and U18999 (N_18999,N_17853,N_17032);
nand U19000 (N_19000,N_18152,N_18846);
or U19001 (N_19001,N_18867,N_18068);
and U19002 (N_19002,N_18914,N_18140);
xnor U19003 (N_19003,N_18711,N_18721);
or U19004 (N_19004,N_18714,N_18266);
nor U19005 (N_19005,N_18813,N_18079);
or U19006 (N_19006,N_18248,N_18179);
nor U19007 (N_19007,N_18506,N_18476);
or U19008 (N_19008,N_18393,N_18116);
nand U19009 (N_19009,N_18906,N_18467);
and U19010 (N_19010,N_18960,N_18427);
xnor U19011 (N_19011,N_18433,N_18866);
xnor U19012 (N_19012,N_18600,N_18363);
nand U19013 (N_19013,N_18730,N_18466);
xnor U19014 (N_19014,N_18579,N_18539);
xnor U19015 (N_19015,N_18536,N_18135);
nor U19016 (N_19016,N_18608,N_18702);
and U19017 (N_19017,N_18159,N_18840);
xor U19018 (N_19018,N_18122,N_18346);
nor U19019 (N_19019,N_18250,N_18035);
nor U19020 (N_19020,N_18665,N_18145);
and U19021 (N_19021,N_18304,N_18217);
and U19022 (N_19022,N_18580,N_18954);
nor U19023 (N_19023,N_18861,N_18676);
and U19024 (N_19024,N_18596,N_18207);
and U19025 (N_19025,N_18057,N_18432);
nand U19026 (N_19026,N_18184,N_18471);
nand U19027 (N_19027,N_18630,N_18383);
and U19028 (N_19028,N_18055,N_18519);
and U19029 (N_19029,N_18123,N_18104);
nor U19030 (N_19030,N_18913,N_18884);
and U19031 (N_19031,N_18288,N_18237);
nand U19032 (N_19032,N_18321,N_18933);
xor U19033 (N_19033,N_18921,N_18934);
or U19034 (N_19034,N_18632,N_18703);
xor U19035 (N_19035,N_18053,N_18768);
and U19036 (N_19036,N_18518,N_18688);
or U19037 (N_19037,N_18149,N_18949);
nand U19038 (N_19038,N_18917,N_18710);
xor U19039 (N_19039,N_18113,N_18107);
or U19040 (N_19040,N_18182,N_18190);
nand U19041 (N_19041,N_18621,N_18064);
xor U19042 (N_19042,N_18005,N_18357);
or U19043 (N_19043,N_18114,N_18628);
xor U19044 (N_19044,N_18388,N_18426);
or U19045 (N_19045,N_18749,N_18661);
nor U19046 (N_19046,N_18338,N_18213);
xor U19047 (N_19047,N_18351,N_18110);
xor U19048 (N_19048,N_18429,N_18627);
nand U19049 (N_19049,N_18886,N_18294);
or U19050 (N_19050,N_18374,N_18824);
or U19051 (N_19051,N_18946,N_18958);
or U19052 (N_19052,N_18814,N_18095);
or U19053 (N_19053,N_18000,N_18125);
or U19054 (N_19054,N_18137,N_18260);
and U19055 (N_19055,N_18574,N_18236);
xor U19056 (N_19056,N_18528,N_18924);
nand U19057 (N_19057,N_18722,N_18882);
nor U19058 (N_19058,N_18832,N_18075);
nor U19059 (N_19059,N_18619,N_18708);
nand U19060 (N_19060,N_18955,N_18747);
nor U19061 (N_19061,N_18558,N_18133);
nand U19062 (N_19062,N_18512,N_18333);
and U19063 (N_19063,N_18436,N_18717);
nor U19064 (N_19064,N_18398,N_18218);
nand U19065 (N_19065,N_18381,N_18533);
nand U19066 (N_19066,N_18119,N_18617);
nor U19067 (N_19067,N_18166,N_18061);
or U19068 (N_19068,N_18508,N_18146);
xor U19069 (N_19069,N_18953,N_18431);
and U19070 (N_19070,N_18441,N_18544);
nor U19071 (N_19071,N_18698,N_18736);
nand U19072 (N_19072,N_18550,N_18775);
or U19073 (N_19073,N_18977,N_18912);
nor U19074 (N_19074,N_18607,N_18058);
or U19075 (N_19075,N_18578,N_18738);
xor U19076 (N_19076,N_18451,N_18496);
nand U19077 (N_19077,N_18888,N_18935);
nand U19078 (N_19078,N_18943,N_18648);
and U19079 (N_19079,N_18989,N_18595);
nand U19080 (N_19080,N_18662,N_18167);
and U19081 (N_19081,N_18894,N_18087);
or U19082 (N_19082,N_18985,N_18102);
and U19083 (N_19083,N_18754,N_18234);
and U19084 (N_19084,N_18868,N_18379);
nand U19085 (N_19085,N_18594,N_18660);
and U19086 (N_19086,N_18643,N_18928);
nand U19087 (N_19087,N_18664,N_18671);
nand U19088 (N_19088,N_18575,N_18838);
nor U19089 (N_19089,N_18270,N_18313);
nand U19090 (N_19090,N_18988,N_18926);
xnor U19091 (N_19091,N_18175,N_18981);
nand U19092 (N_19092,N_18879,N_18870);
xnor U19093 (N_19093,N_18434,N_18931);
xnor U19094 (N_19094,N_18446,N_18899);
nor U19095 (N_19095,N_18654,N_18147);
and U19096 (N_19096,N_18240,N_18060);
or U19097 (N_19097,N_18718,N_18878);
and U19098 (N_19098,N_18601,N_18535);
nand U19099 (N_19099,N_18825,N_18138);
or U19100 (N_19100,N_18997,N_18983);
and U19101 (N_19101,N_18547,N_18587);
or U19102 (N_19102,N_18039,N_18844);
or U19103 (N_19103,N_18514,N_18850);
nor U19104 (N_19104,N_18895,N_18111);
nor U19105 (N_19105,N_18545,N_18872);
xnor U19106 (N_19106,N_18097,N_18416);
nand U19107 (N_19107,N_18479,N_18742);
and U19108 (N_19108,N_18078,N_18130);
xor U19109 (N_19109,N_18475,N_18284);
nor U19110 (N_19110,N_18833,N_18085);
and U19111 (N_19111,N_18724,N_18827);
or U19112 (N_19112,N_18455,N_18625);
or U19113 (N_19113,N_18999,N_18344);
nand U19114 (N_19114,N_18076,N_18158);
nand U19115 (N_19115,N_18837,N_18776);
xnor U19116 (N_19116,N_18219,N_18740);
or U19117 (N_19117,N_18232,N_18705);
and U19118 (N_19118,N_18561,N_18945);
and U19119 (N_19119,N_18382,N_18750);
or U19120 (N_19120,N_18155,N_18864);
nor U19121 (N_19121,N_18081,N_18369);
nor U19122 (N_19122,N_18975,N_18719);
nor U19123 (N_19123,N_18598,N_18020);
and U19124 (N_19124,N_18731,N_18101);
or U19125 (N_19125,N_18969,N_18787);
nand U19126 (N_19126,N_18187,N_18817);
nor U19127 (N_19127,N_18340,N_18525);
nor U19128 (N_19128,N_18809,N_18729);
nand U19129 (N_19129,N_18847,N_18021);
nand U19130 (N_19130,N_18411,N_18973);
and U19131 (N_19131,N_18229,N_18571);
xnor U19132 (N_19132,N_18568,N_18329);
or U19133 (N_19133,N_18936,N_18073);
xor U19134 (N_19134,N_18728,N_18212);
and U19135 (N_19135,N_18353,N_18994);
nand U19136 (N_19136,N_18741,N_18406);
xnor U19137 (N_19137,N_18693,N_18942);
xor U19138 (N_19138,N_18515,N_18077);
nand U19139 (N_19139,N_18883,N_18919);
or U19140 (N_19140,N_18183,N_18551);
xnor U19141 (N_19141,N_18689,N_18759);
and U19142 (N_19142,N_18366,N_18745);
nand U19143 (N_19143,N_18385,N_18018);
and U19144 (N_19144,N_18652,N_18490);
xor U19145 (N_19145,N_18129,N_18339);
and U19146 (N_19146,N_18238,N_18979);
nand U19147 (N_19147,N_18770,N_18161);
xnor U19148 (N_19148,N_18541,N_18410);
and U19149 (N_19149,N_18940,N_18634);
and U19150 (N_19150,N_18450,N_18573);
xor U19151 (N_19151,N_18589,N_18700);
nor U19152 (N_19152,N_18247,N_18143);
nand U19153 (N_19153,N_18725,N_18562);
xnor U19154 (N_19154,N_18891,N_18836);
and U19155 (N_19155,N_18224,N_18144);
and U19156 (N_19156,N_18922,N_18364);
and U19157 (N_19157,N_18042,N_18791);
xnor U19158 (N_19158,N_18413,N_18713);
or U19159 (N_19159,N_18696,N_18126);
nor U19160 (N_19160,N_18811,N_18164);
nor U19161 (N_19161,N_18963,N_18666);
or U19162 (N_19162,N_18509,N_18249);
nor U19163 (N_19163,N_18204,N_18865);
nor U19164 (N_19164,N_18786,N_18602);
xnor U19165 (N_19165,N_18362,N_18358);
nor U19166 (N_19166,N_18459,N_18656);
nand U19167 (N_19167,N_18819,N_18905);
or U19168 (N_19168,N_18045,N_18692);
and U19169 (N_19169,N_18323,N_18485);
xor U19170 (N_19170,N_18559,N_18510);
nor U19171 (N_19171,N_18324,N_18390);
xor U19172 (N_19172,N_18604,N_18992);
and U19173 (N_19173,N_18881,N_18877);
xnor U19174 (N_19174,N_18089,N_18059);
nor U19175 (N_19175,N_18769,N_18428);
or U19176 (N_19176,N_18456,N_18845);
nand U19177 (N_19177,N_18549,N_18762);
xnor U19178 (N_19178,N_18556,N_18370);
xor U19179 (N_19179,N_18520,N_18307);
or U19180 (N_19180,N_18258,N_18253);
nor U19181 (N_19181,N_18707,N_18373);
nor U19182 (N_19182,N_18778,N_18056);
nor U19183 (N_19183,N_18835,N_18136);
xor U19184 (N_19184,N_18501,N_18030);
or U19185 (N_19185,N_18488,N_18016);
nand U19186 (N_19186,N_18334,N_18690);
and U19187 (N_19187,N_18640,N_18567);
xor U19188 (N_19188,N_18848,N_18153);
nand U19189 (N_19189,N_18022,N_18156);
nor U19190 (N_19190,N_18169,N_18291);
nand U19191 (N_19191,N_18522,N_18440);
nand U19192 (N_19192,N_18618,N_18537);
nor U19193 (N_19193,N_18189,N_18025);
and U19194 (N_19194,N_18597,N_18442);
and U19195 (N_19195,N_18534,N_18265);
xor U19196 (N_19196,N_18091,N_18215);
or U19197 (N_19197,N_18771,N_18259);
nand U19198 (N_19198,N_18117,N_18317);
or U19199 (N_19199,N_18548,N_18585);
and U19200 (N_19200,N_18804,N_18829);
or U19201 (N_19201,N_18910,N_18008);
and U19202 (N_19202,N_18629,N_18243);
nand U19203 (N_19203,N_18916,N_18326);
and U19204 (N_19204,N_18447,N_18854);
xnor U19205 (N_19205,N_18487,N_18435);
xnor U19206 (N_19206,N_18088,N_18380);
nor U19207 (N_19207,N_18191,N_18320);
nor U19208 (N_19208,N_18150,N_18929);
or U19209 (N_19209,N_18576,N_18686);
xnor U19210 (N_19210,N_18869,N_18735);
nor U19211 (N_19211,N_18785,N_18503);
xnor U19212 (N_19212,N_18843,N_18430);
xor U19213 (N_19213,N_18802,N_18423);
and U19214 (N_19214,N_18287,N_18492);
nand U19215 (N_19215,N_18277,N_18310);
or U19216 (N_19216,N_18401,N_18659);
nor U19217 (N_19217,N_18743,N_18974);
or U19218 (N_19218,N_18566,N_18887);
and U19219 (N_19219,N_18474,N_18641);
or U19220 (N_19220,N_18332,N_18186);
or U19221 (N_19221,N_18460,N_18746);
nor U19222 (N_19222,N_18026,N_18908);
nand U19223 (N_19223,N_18684,N_18970);
xor U19224 (N_19224,N_18511,N_18472);
xnor U19225 (N_19225,N_18653,N_18674);
nand U19226 (N_19226,N_18599,N_18180);
nor U19227 (N_19227,N_18706,N_18695);
xor U19228 (N_19228,N_18051,N_18495);
nor U19229 (N_19229,N_18546,N_18124);
or U19230 (N_19230,N_18790,N_18203);
and U19231 (N_19231,N_18414,N_18484);
nand U19232 (N_19232,N_18726,N_18202);
nor U19233 (N_19233,N_18048,N_18192);
and U19234 (N_19234,N_18314,N_18221);
or U19235 (N_19235,N_18360,N_18614);
nand U19236 (N_19236,N_18134,N_18682);
and U19237 (N_19237,N_18343,N_18583);
nor U19238 (N_19238,N_18925,N_18372);
and U19239 (N_19239,N_18327,N_18386);
or U19240 (N_19240,N_18408,N_18831);
xor U19241 (N_19241,N_18763,N_18049);
nand U19242 (N_19242,N_18720,N_18465);
nor U19243 (N_19243,N_18828,N_18815);
nor U19244 (N_19244,N_18683,N_18067);
nor U19245 (N_19245,N_18712,N_18084);
or U19246 (N_19246,N_18415,N_18966);
nor U19247 (N_19247,N_18563,N_18670);
or U19248 (N_19248,N_18489,N_18148);
or U19249 (N_19249,N_18392,N_18131);
xnor U19250 (N_19250,N_18311,N_18685);
nand U19251 (N_19251,N_18593,N_18118);
or U19252 (N_19252,N_18753,N_18792);
xor U19253 (N_19253,N_18855,N_18011);
nor U19254 (N_19254,N_18054,N_18090);
or U19255 (N_19255,N_18109,N_18673);
nand U19256 (N_19256,N_18283,N_18803);
or U19257 (N_19257,N_18289,N_18890);
or U19258 (N_19258,N_18453,N_18739);
nand U19259 (N_19259,N_18069,N_18875);
nand U19260 (N_19260,N_18391,N_18160);
nand U19261 (N_19261,N_18115,N_18610);
nor U19262 (N_19262,N_18444,N_18419);
and U19263 (N_19263,N_18330,N_18454);
or U19264 (N_19264,N_18093,N_18893);
xor U19265 (N_19265,N_18529,N_18478);
nor U19266 (N_19266,N_18246,N_18469);
xnor U19267 (N_19267,N_18959,N_18553);
nor U19268 (N_19268,N_18230,N_18798);
nor U19269 (N_19269,N_18603,N_18586);
nand U19270 (N_19270,N_18157,N_18760);
or U19271 (N_19271,N_18151,N_18498);
or U19272 (N_19272,N_18278,N_18582);
and U19273 (N_19273,N_18376,N_18863);
nand U19274 (N_19274,N_18033,N_18038);
nor U19275 (N_19275,N_18178,N_18062);
and U19276 (N_19276,N_18691,N_18231);
nand U19277 (N_19277,N_18470,N_18588);
nand U19278 (N_19278,N_18306,N_18396);
or U19279 (N_19279,N_18612,N_18907);
or U19280 (N_19280,N_18504,N_18675);
xor U19281 (N_19281,N_18402,N_18687);
and U19282 (N_19282,N_18560,N_18421);
or U19283 (N_19283,N_18188,N_18106);
and U19284 (N_19284,N_18611,N_18464);
and U19285 (N_19285,N_18852,N_18672);
or U19286 (N_19286,N_18354,N_18772);
xnor U19287 (N_19287,N_18968,N_18400);
nor U19288 (N_19288,N_18856,N_18245);
or U19289 (N_19289,N_18302,N_18208);
or U19290 (N_19290,N_18816,N_18028);
nand U19291 (N_19291,N_18513,N_18885);
and U19292 (N_19292,N_18375,N_18063);
nor U19293 (N_19293,N_18807,N_18318);
and U19294 (N_19294,N_18173,N_18951);
and U19295 (N_19295,N_18262,N_18701);
xnor U19296 (N_19296,N_18909,N_18923);
nor U19297 (N_19297,N_18801,N_18244);
or U19298 (N_19298,N_18932,N_18663);
and U19299 (N_19299,N_18378,N_18995);
or U19300 (N_19300,N_18029,N_18859);
or U19301 (N_19301,N_18737,N_18577);
or U19302 (N_19302,N_18716,N_18538);
and U19303 (N_19303,N_18046,N_18920);
or U19304 (N_19304,N_18261,N_18540);
xnor U19305 (N_19305,N_18987,N_18609);
or U19306 (N_19306,N_18002,N_18633);
nand U19307 (N_19307,N_18336,N_18225);
or U19308 (N_19308,N_18437,N_18233);
nor U19309 (N_19309,N_18036,N_18649);
nor U19310 (N_19310,N_18425,N_18473);
or U19311 (N_19311,N_18482,N_18680);
and U19312 (N_19312,N_18342,N_18194);
xnor U19313 (N_19313,N_18004,N_18279);
or U19314 (N_19314,N_18499,N_18412);
and U19315 (N_19315,N_18468,N_18715);
xnor U19316 (N_19316,N_18001,N_18239);
nand U19317 (N_19317,N_18781,N_18751);
nor U19318 (N_19318,N_18918,N_18991);
nor U19319 (N_19319,N_18849,N_18552);
and U19320 (N_19320,N_18842,N_18555);
and U19321 (N_19321,N_18210,N_18993);
nor U19322 (N_19322,N_18198,N_18316);
xnor U19323 (N_19323,N_18530,N_18622);
nand U19324 (N_19324,N_18403,N_18581);
nor U19325 (N_19325,N_18226,N_18584);
nand U19326 (N_19326,N_18037,N_18500);
or U19327 (N_19327,N_18174,N_18368);
nor U19328 (N_19328,N_18650,N_18857);
nor U19329 (N_19329,N_18105,N_18290);
and U19330 (N_19330,N_18214,N_18862);
xor U19331 (N_19331,N_18789,N_18570);
or U19332 (N_19332,N_18681,N_18624);
nor U19333 (N_19333,N_18024,N_18003);
or U19334 (N_19334,N_18911,N_18027);
or U19335 (N_19335,N_18723,N_18154);
nand U19336 (N_19336,N_18784,N_18616);
and U19337 (N_19337,N_18377,N_18295);
xor U19338 (N_19338,N_18752,N_18980);
nand U19339 (N_19339,N_18978,N_18761);
xor U19340 (N_19340,N_18971,N_18438);
xor U19341 (N_19341,N_18205,N_18309);
nor U19342 (N_19342,N_18766,N_18590);
nor U19343 (N_19343,N_18502,N_18669);
or U19344 (N_19344,N_18276,N_18420);
or U19345 (N_19345,N_18193,N_18812);
or U19346 (N_19346,N_18361,N_18252);
nand U19347 (N_19347,N_18565,N_18255);
nor U19348 (N_19348,N_18904,N_18086);
xnor U19349 (N_19349,N_18325,N_18543);
nor U19350 (N_19350,N_18418,N_18635);
nand U19351 (N_19351,N_18795,N_18070);
or U19352 (N_19352,N_18898,N_18834);
or U19353 (N_19353,N_18315,N_18505);
and U19354 (N_19354,N_18301,N_18976);
nor U19355 (N_19355,N_18507,N_18794);
nor U19356 (N_19356,N_18774,N_18986);
xor U19357 (N_19357,N_18439,N_18962);
and U19358 (N_19358,N_18092,N_18032);
xor U19359 (N_19359,N_18860,N_18200);
xor U19360 (N_19360,N_18312,N_18196);
nor U19361 (N_19361,N_18658,N_18052);
nand U19362 (N_19362,N_18554,N_18462);
or U19363 (N_19363,N_18275,N_18010);
or U19364 (N_19364,N_18162,N_18572);
nand U19365 (N_19365,N_18172,N_18083);
nor U19366 (N_19366,N_18494,N_18251);
or U19367 (N_19367,N_18235,N_18096);
nor U19368 (N_19368,N_18939,N_18044);
nor U19369 (N_19369,N_18915,N_18254);
xor U19370 (N_19370,N_18477,N_18965);
and U19371 (N_19371,N_18532,N_18493);
and U19372 (N_19372,N_18796,N_18072);
and U19373 (N_19373,N_18263,N_18269);
nand U19374 (N_19374,N_18637,N_18697);
nand U19375 (N_19375,N_18734,N_18103);
and U19376 (N_19376,N_18367,N_18756);
nand U19377 (N_19377,N_18080,N_18165);
xnor U19378 (N_19378,N_18564,N_18331);
nor U19379 (N_19379,N_18220,N_18181);
nand U19380 (N_19380,N_18041,N_18389);
and U19381 (N_19381,N_18043,N_18941);
nor U19382 (N_19382,N_18195,N_18349);
nand U19383 (N_19383,N_18808,N_18098);
nor U19384 (N_19384,N_18897,N_18788);
xnor U19385 (N_19385,N_18206,N_18930);
or U19386 (N_19386,N_18542,N_18557);
nor U19387 (N_19387,N_18800,N_18121);
and U19388 (N_19388,N_18591,N_18355);
nand U19389 (N_19389,N_18066,N_18889);
or U19390 (N_19390,N_18605,N_18359);
nand U19391 (N_19391,N_18405,N_18944);
xor U19392 (N_19392,N_18938,N_18461);
nor U19393 (N_19393,N_18211,N_18839);
or U19394 (N_19394,N_18733,N_18704);
and U19395 (N_19395,N_18384,N_18242);
and U19396 (N_19396,N_18082,N_18452);
nand U19397 (N_19397,N_18957,N_18758);
and U19398 (N_19398,N_18448,N_18282);
xnor U19399 (N_19399,N_18806,N_18352);
nand U19400 (N_19400,N_18345,N_18679);
and U19401 (N_19401,N_18657,N_18727);
nor U19402 (N_19402,N_18748,N_18257);
or U19403 (N_19403,N_18142,N_18015);
nor U19404 (N_19404,N_18006,N_18777);
xnor U19405 (N_19405,N_18858,N_18371);
xnor U19406 (N_19406,N_18303,N_18099);
nor U19407 (N_19407,N_18201,N_18606);
or U19408 (N_19408,N_18399,N_18222);
or U19409 (N_19409,N_18335,N_18480);
nor U19410 (N_19410,N_18779,N_18132);
or U19411 (N_19411,N_18851,N_18620);
and U19412 (N_19412,N_18782,N_18171);
and U19413 (N_19413,N_18409,N_18964);
or U19414 (N_19414,N_18014,N_18636);
or U19415 (N_19415,N_18216,N_18443);
or U19416 (N_19416,N_18521,N_18516);
nor U19417 (N_19417,N_18292,N_18972);
nand U19418 (N_19418,N_18365,N_18163);
nor U19419 (N_19419,N_18286,N_18638);
or U19420 (N_19420,N_18651,N_18818);
or U19421 (N_19421,N_18424,N_18677);
xnor U19422 (N_19422,N_18463,N_18871);
and U19423 (N_19423,N_18271,N_18694);
or U19424 (N_19424,N_18780,N_18170);
and U19425 (N_19425,N_18830,N_18387);
nand U19426 (N_19426,N_18139,N_18876);
nand U19427 (N_19427,N_18305,N_18199);
and U19428 (N_19428,N_18937,N_18094);
xor U19429 (N_19429,N_18322,N_18655);
nand U19430 (N_19430,N_18668,N_18645);
xor U19431 (N_19431,N_18281,N_18826);
nor U19432 (N_19432,N_18407,N_18982);
or U19433 (N_19433,N_18280,N_18527);
or U19434 (N_19434,N_18892,N_18793);
or U19435 (N_19435,N_18497,N_18961);
or U19436 (N_19436,N_18017,N_18209);
nor U19437 (N_19437,N_18990,N_18296);
or U19438 (N_19438,N_18293,N_18642);
xor U19439 (N_19439,N_18639,N_18013);
and U19440 (N_19440,N_18267,N_18822);
and U19441 (N_19441,N_18458,N_18264);
nand U19442 (N_19442,N_18950,N_18732);
xor U19443 (N_19443,N_18397,N_18023);
nor U19444 (N_19444,N_18647,N_18967);
nor U19445 (N_19445,N_18457,N_18873);
and U19446 (N_19446,N_18394,N_18228);
and U19447 (N_19447,N_18341,N_18308);
nand U19448 (N_19448,N_18273,N_18422);
nand U19449 (N_19449,N_18256,N_18823);
nand U19450 (N_19450,N_18128,N_18517);
nor U19451 (N_19451,N_18483,N_18297);
or U19452 (N_19452,N_18065,N_18007);
nand U19453 (N_19453,N_18757,N_18896);
and U19454 (N_19454,N_18031,N_18404);
nor U19455 (N_19455,N_18100,N_18185);
and U19456 (N_19456,N_18034,N_18523);
nor U19457 (N_19457,N_18012,N_18613);
xnor U19458 (N_19458,N_18040,N_18678);
nand U19459 (N_19459,N_18120,N_18900);
xor U19460 (N_19460,N_18821,N_18947);
nand U19461 (N_19461,N_18347,N_18699);
xor U19462 (N_19462,N_18764,N_18773);
nand U19463 (N_19463,N_18952,N_18623);
xor U19464 (N_19464,N_18272,N_18481);
nor U19465 (N_19465,N_18927,N_18644);
or U19466 (N_19466,N_18298,N_18141);
nor U19467 (N_19467,N_18984,N_18274);
xnor U19468 (N_19468,N_18880,N_18112);
and U19469 (N_19469,N_18783,N_18319);
xor U19470 (N_19470,N_18009,N_18874);
and U19471 (N_19471,N_18299,N_18531);
nor U19472 (N_19472,N_18998,N_18903);
or U19473 (N_19473,N_18449,N_18799);
xnor U19474 (N_19474,N_18417,N_18071);
nor U19475 (N_19475,N_18395,N_18074);
nor U19476 (N_19476,N_18300,N_18853);
or U19477 (N_19477,N_18901,N_18646);
and U19478 (N_19478,N_18667,N_18176);
nor U19479 (N_19479,N_18820,N_18356);
xor U19480 (N_19480,N_18765,N_18197);
nand U19481 (N_19481,N_18223,N_18127);
nand U19482 (N_19482,N_18350,N_18268);
nand U19483 (N_19483,N_18241,N_18755);
and U19484 (N_19484,N_18337,N_18524);
nand U19485 (N_19485,N_18177,N_18797);
nor U19486 (N_19486,N_18050,N_18956);
or U19487 (N_19487,N_18709,N_18486);
xnor U19488 (N_19488,N_18810,N_18626);
or U19489 (N_19489,N_18227,N_18805);
nor U19490 (N_19490,N_18445,N_18902);
nor U19491 (N_19491,N_18491,N_18108);
and U19492 (N_19492,N_18948,N_18019);
nor U19493 (N_19493,N_18996,N_18767);
and U19494 (N_19494,N_18569,N_18047);
xnor U19495 (N_19495,N_18328,N_18348);
nand U19496 (N_19496,N_18285,N_18744);
and U19497 (N_19497,N_18615,N_18841);
xor U19498 (N_19498,N_18631,N_18168);
xor U19499 (N_19499,N_18526,N_18592);
and U19500 (N_19500,N_18784,N_18073);
or U19501 (N_19501,N_18018,N_18659);
xnor U19502 (N_19502,N_18880,N_18499);
or U19503 (N_19503,N_18713,N_18328);
or U19504 (N_19504,N_18433,N_18298);
or U19505 (N_19505,N_18045,N_18730);
nor U19506 (N_19506,N_18057,N_18136);
and U19507 (N_19507,N_18229,N_18143);
or U19508 (N_19508,N_18135,N_18193);
xor U19509 (N_19509,N_18443,N_18460);
and U19510 (N_19510,N_18704,N_18498);
nor U19511 (N_19511,N_18136,N_18998);
or U19512 (N_19512,N_18228,N_18490);
nand U19513 (N_19513,N_18176,N_18063);
nor U19514 (N_19514,N_18245,N_18464);
and U19515 (N_19515,N_18333,N_18010);
nor U19516 (N_19516,N_18129,N_18776);
xnor U19517 (N_19517,N_18134,N_18533);
nor U19518 (N_19518,N_18244,N_18565);
nor U19519 (N_19519,N_18460,N_18083);
xnor U19520 (N_19520,N_18631,N_18392);
xor U19521 (N_19521,N_18221,N_18615);
and U19522 (N_19522,N_18309,N_18690);
xor U19523 (N_19523,N_18271,N_18968);
nand U19524 (N_19524,N_18451,N_18986);
nor U19525 (N_19525,N_18708,N_18763);
xor U19526 (N_19526,N_18147,N_18453);
xor U19527 (N_19527,N_18481,N_18458);
or U19528 (N_19528,N_18274,N_18395);
xor U19529 (N_19529,N_18837,N_18498);
or U19530 (N_19530,N_18859,N_18601);
nor U19531 (N_19531,N_18635,N_18770);
nor U19532 (N_19532,N_18976,N_18219);
nor U19533 (N_19533,N_18769,N_18133);
nor U19534 (N_19534,N_18785,N_18287);
and U19535 (N_19535,N_18521,N_18906);
nor U19536 (N_19536,N_18444,N_18521);
or U19537 (N_19537,N_18566,N_18973);
nor U19538 (N_19538,N_18806,N_18557);
nand U19539 (N_19539,N_18173,N_18106);
nor U19540 (N_19540,N_18655,N_18288);
and U19541 (N_19541,N_18387,N_18312);
or U19542 (N_19542,N_18526,N_18123);
nand U19543 (N_19543,N_18346,N_18139);
xor U19544 (N_19544,N_18067,N_18251);
and U19545 (N_19545,N_18591,N_18114);
nand U19546 (N_19546,N_18982,N_18828);
or U19547 (N_19547,N_18734,N_18547);
and U19548 (N_19548,N_18337,N_18628);
xor U19549 (N_19549,N_18720,N_18212);
and U19550 (N_19550,N_18070,N_18980);
or U19551 (N_19551,N_18475,N_18772);
nor U19552 (N_19552,N_18633,N_18977);
and U19553 (N_19553,N_18002,N_18604);
and U19554 (N_19554,N_18505,N_18379);
nor U19555 (N_19555,N_18211,N_18249);
nor U19556 (N_19556,N_18335,N_18746);
or U19557 (N_19557,N_18789,N_18153);
or U19558 (N_19558,N_18054,N_18988);
and U19559 (N_19559,N_18493,N_18142);
nor U19560 (N_19560,N_18406,N_18286);
nand U19561 (N_19561,N_18417,N_18685);
and U19562 (N_19562,N_18599,N_18426);
xnor U19563 (N_19563,N_18327,N_18111);
xor U19564 (N_19564,N_18451,N_18372);
nand U19565 (N_19565,N_18032,N_18784);
or U19566 (N_19566,N_18014,N_18095);
nand U19567 (N_19567,N_18691,N_18071);
nand U19568 (N_19568,N_18905,N_18681);
nand U19569 (N_19569,N_18839,N_18424);
xnor U19570 (N_19570,N_18212,N_18523);
xnor U19571 (N_19571,N_18006,N_18790);
or U19572 (N_19572,N_18575,N_18565);
nand U19573 (N_19573,N_18012,N_18867);
or U19574 (N_19574,N_18091,N_18257);
xor U19575 (N_19575,N_18343,N_18782);
or U19576 (N_19576,N_18349,N_18326);
nor U19577 (N_19577,N_18694,N_18259);
or U19578 (N_19578,N_18210,N_18262);
nor U19579 (N_19579,N_18819,N_18693);
or U19580 (N_19580,N_18139,N_18052);
xnor U19581 (N_19581,N_18932,N_18651);
and U19582 (N_19582,N_18153,N_18350);
nor U19583 (N_19583,N_18946,N_18989);
nand U19584 (N_19584,N_18298,N_18983);
and U19585 (N_19585,N_18991,N_18655);
and U19586 (N_19586,N_18050,N_18904);
nand U19587 (N_19587,N_18950,N_18582);
and U19588 (N_19588,N_18591,N_18041);
xor U19589 (N_19589,N_18095,N_18534);
and U19590 (N_19590,N_18781,N_18547);
nor U19591 (N_19591,N_18404,N_18680);
nand U19592 (N_19592,N_18843,N_18490);
and U19593 (N_19593,N_18389,N_18393);
nor U19594 (N_19594,N_18180,N_18016);
or U19595 (N_19595,N_18545,N_18076);
nor U19596 (N_19596,N_18531,N_18330);
xnor U19597 (N_19597,N_18287,N_18577);
or U19598 (N_19598,N_18547,N_18766);
nand U19599 (N_19599,N_18446,N_18630);
xor U19600 (N_19600,N_18856,N_18747);
and U19601 (N_19601,N_18138,N_18286);
xor U19602 (N_19602,N_18369,N_18124);
xnor U19603 (N_19603,N_18774,N_18631);
xnor U19604 (N_19604,N_18270,N_18464);
nor U19605 (N_19605,N_18310,N_18032);
nand U19606 (N_19606,N_18552,N_18693);
or U19607 (N_19607,N_18886,N_18885);
nand U19608 (N_19608,N_18699,N_18757);
nand U19609 (N_19609,N_18143,N_18810);
or U19610 (N_19610,N_18565,N_18021);
or U19611 (N_19611,N_18874,N_18687);
or U19612 (N_19612,N_18336,N_18062);
and U19613 (N_19613,N_18545,N_18029);
xor U19614 (N_19614,N_18481,N_18161);
xnor U19615 (N_19615,N_18499,N_18229);
nor U19616 (N_19616,N_18134,N_18935);
or U19617 (N_19617,N_18693,N_18438);
or U19618 (N_19618,N_18808,N_18058);
xor U19619 (N_19619,N_18264,N_18958);
xnor U19620 (N_19620,N_18880,N_18400);
nand U19621 (N_19621,N_18599,N_18360);
nor U19622 (N_19622,N_18977,N_18452);
or U19623 (N_19623,N_18070,N_18583);
xnor U19624 (N_19624,N_18302,N_18305);
or U19625 (N_19625,N_18488,N_18324);
xnor U19626 (N_19626,N_18979,N_18146);
nor U19627 (N_19627,N_18740,N_18619);
nand U19628 (N_19628,N_18335,N_18084);
or U19629 (N_19629,N_18782,N_18864);
or U19630 (N_19630,N_18298,N_18138);
nor U19631 (N_19631,N_18389,N_18829);
and U19632 (N_19632,N_18989,N_18067);
nor U19633 (N_19633,N_18276,N_18934);
nor U19634 (N_19634,N_18236,N_18578);
and U19635 (N_19635,N_18411,N_18853);
nor U19636 (N_19636,N_18927,N_18181);
and U19637 (N_19637,N_18506,N_18395);
or U19638 (N_19638,N_18364,N_18342);
xnor U19639 (N_19639,N_18538,N_18638);
and U19640 (N_19640,N_18714,N_18235);
and U19641 (N_19641,N_18177,N_18323);
and U19642 (N_19642,N_18552,N_18493);
nand U19643 (N_19643,N_18459,N_18079);
nand U19644 (N_19644,N_18745,N_18356);
or U19645 (N_19645,N_18320,N_18518);
xor U19646 (N_19646,N_18298,N_18176);
xnor U19647 (N_19647,N_18823,N_18874);
nand U19648 (N_19648,N_18004,N_18085);
or U19649 (N_19649,N_18039,N_18568);
and U19650 (N_19650,N_18768,N_18273);
or U19651 (N_19651,N_18806,N_18511);
or U19652 (N_19652,N_18150,N_18407);
nand U19653 (N_19653,N_18720,N_18541);
or U19654 (N_19654,N_18940,N_18694);
xnor U19655 (N_19655,N_18560,N_18102);
and U19656 (N_19656,N_18111,N_18495);
nor U19657 (N_19657,N_18528,N_18907);
and U19658 (N_19658,N_18360,N_18505);
or U19659 (N_19659,N_18105,N_18563);
xnor U19660 (N_19660,N_18029,N_18475);
or U19661 (N_19661,N_18724,N_18421);
nor U19662 (N_19662,N_18347,N_18442);
and U19663 (N_19663,N_18538,N_18456);
nor U19664 (N_19664,N_18173,N_18217);
nand U19665 (N_19665,N_18280,N_18998);
and U19666 (N_19666,N_18119,N_18566);
and U19667 (N_19667,N_18603,N_18264);
nor U19668 (N_19668,N_18916,N_18879);
nor U19669 (N_19669,N_18088,N_18664);
nand U19670 (N_19670,N_18074,N_18253);
nor U19671 (N_19671,N_18533,N_18926);
xnor U19672 (N_19672,N_18235,N_18782);
nand U19673 (N_19673,N_18851,N_18727);
or U19674 (N_19674,N_18669,N_18767);
nor U19675 (N_19675,N_18474,N_18447);
or U19676 (N_19676,N_18478,N_18219);
and U19677 (N_19677,N_18475,N_18036);
and U19678 (N_19678,N_18691,N_18789);
and U19679 (N_19679,N_18780,N_18882);
nor U19680 (N_19680,N_18177,N_18916);
nand U19681 (N_19681,N_18327,N_18507);
or U19682 (N_19682,N_18337,N_18110);
xnor U19683 (N_19683,N_18694,N_18941);
xor U19684 (N_19684,N_18267,N_18790);
or U19685 (N_19685,N_18263,N_18548);
xnor U19686 (N_19686,N_18994,N_18723);
nand U19687 (N_19687,N_18387,N_18187);
and U19688 (N_19688,N_18609,N_18068);
nand U19689 (N_19689,N_18092,N_18204);
or U19690 (N_19690,N_18967,N_18368);
or U19691 (N_19691,N_18076,N_18560);
and U19692 (N_19692,N_18809,N_18356);
nor U19693 (N_19693,N_18884,N_18420);
and U19694 (N_19694,N_18427,N_18724);
or U19695 (N_19695,N_18460,N_18728);
and U19696 (N_19696,N_18305,N_18112);
nor U19697 (N_19697,N_18394,N_18978);
xor U19698 (N_19698,N_18395,N_18730);
and U19699 (N_19699,N_18025,N_18178);
or U19700 (N_19700,N_18482,N_18821);
nand U19701 (N_19701,N_18758,N_18958);
and U19702 (N_19702,N_18680,N_18240);
nand U19703 (N_19703,N_18067,N_18951);
and U19704 (N_19704,N_18059,N_18959);
nor U19705 (N_19705,N_18284,N_18929);
and U19706 (N_19706,N_18009,N_18007);
and U19707 (N_19707,N_18289,N_18877);
or U19708 (N_19708,N_18491,N_18557);
and U19709 (N_19709,N_18894,N_18116);
or U19710 (N_19710,N_18764,N_18753);
nor U19711 (N_19711,N_18529,N_18255);
nor U19712 (N_19712,N_18269,N_18643);
nor U19713 (N_19713,N_18541,N_18897);
and U19714 (N_19714,N_18793,N_18330);
or U19715 (N_19715,N_18193,N_18349);
nand U19716 (N_19716,N_18707,N_18914);
xor U19717 (N_19717,N_18804,N_18784);
xor U19718 (N_19718,N_18490,N_18684);
or U19719 (N_19719,N_18899,N_18385);
nand U19720 (N_19720,N_18327,N_18165);
and U19721 (N_19721,N_18515,N_18217);
or U19722 (N_19722,N_18083,N_18297);
or U19723 (N_19723,N_18849,N_18567);
nor U19724 (N_19724,N_18960,N_18972);
and U19725 (N_19725,N_18044,N_18652);
nor U19726 (N_19726,N_18973,N_18339);
and U19727 (N_19727,N_18319,N_18933);
nand U19728 (N_19728,N_18183,N_18723);
xnor U19729 (N_19729,N_18920,N_18866);
xnor U19730 (N_19730,N_18123,N_18514);
nor U19731 (N_19731,N_18423,N_18771);
and U19732 (N_19732,N_18263,N_18623);
nand U19733 (N_19733,N_18281,N_18443);
xor U19734 (N_19734,N_18268,N_18112);
xnor U19735 (N_19735,N_18559,N_18842);
or U19736 (N_19736,N_18039,N_18204);
nand U19737 (N_19737,N_18360,N_18079);
or U19738 (N_19738,N_18307,N_18917);
and U19739 (N_19739,N_18404,N_18916);
or U19740 (N_19740,N_18105,N_18835);
xnor U19741 (N_19741,N_18077,N_18074);
nor U19742 (N_19742,N_18574,N_18768);
or U19743 (N_19743,N_18498,N_18131);
nor U19744 (N_19744,N_18058,N_18919);
and U19745 (N_19745,N_18508,N_18052);
nand U19746 (N_19746,N_18227,N_18830);
nand U19747 (N_19747,N_18502,N_18837);
nand U19748 (N_19748,N_18131,N_18226);
nor U19749 (N_19749,N_18907,N_18891);
xor U19750 (N_19750,N_18814,N_18697);
xnor U19751 (N_19751,N_18272,N_18361);
or U19752 (N_19752,N_18107,N_18294);
xor U19753 (N_19753,N_18138,N_18873);
xnor U19754 (N_19754,N_18660,N_18242);
xnor U19755 (N_19755,N_18341,N_18713);
or U19756 (N_19756,N_18535,N_18349);
nand U19757 (N_19757,N_18647,N_18316);
nand U19758 (N_19758,N_18178,N_18988);
or U19759 (N_19759,N_18408,N_18421);
and U19760 (N_19760,N_18269,N_18503);
or U19761 (N_19761,N_18794,N_18269);
xnor U19762 (N_19762,N_18010,N_18706);
or U19763 (N_19763,N_18839,N_18419);
or U19764 (N_19764,N_18154,N_18510);
or U19765 (N_19765,N_18065,N_18016);
nand U19766 (N_19766,N_18122,N_18553);
nor U19767 (N_19767,N_18854,N_18822);
nand U19768 (N_19768,N_18641,N_18784);
xor U19769 (N_19769,N_18590,N_18293);
nand U19770 (N_19770,N_18501,N_18605);
and U19771 (N_19771,N_18543,N_18780);
nand U19772 (N_19772,N_18941,N_18172);
xnor U19773 (N_19773,N_18247,N_18193);
or U19774 (N_19774,N_18834,N_18860);
xor U19775 (N_19775,N_18263,N_18248);
and U19776 (N_19776,N_18879,N_18060);
xnor U19777 (N_19777,N_18441,N_18760);
xnor U19778 (N_19778,N_18221,N_18520);
xor U19779 (N_19779,N_18941,N_18268);
nand U19780 (N_19780,N_18925,N_18508);
or U19781 (N_19781,N_18519,N_18092);
or U19782 (N_19782,N_18740,N_18554);
nor U19783 (N_19783,N_18286,N_18150);
nor U19784 (N_19784,N_18516,N_18273);
nand U19785 (N_19785,N_18145,N_18441);
nand U19786 (N_19786,N_18965,N_18998);
xor U19787 (N_19787,N_18982,N_18587);
nor U19788 (N_19788,N_18718,N_18224);
nor U19789 (N_19789,N_18685,N_18004);
and U19790 (N_19790,N_18703,N_18943);
and U19791 (N_19791,N_18165,N_18281);
and U19792 (N_19792,N_18434,N_18213);
nand U19793 (N_19793,N_18490,N_18332);
nand U19794 (N_19794,N_18211,N_18154);
or U19795 (N_19795,N_18831,N_18626);
nor U19796 (N_19796,N_18309,N_18416);
nor U19797 (N_19797,N_18938,N_18063);
nor U19798 (N_19798,N_18258,N_18532);
and U19799 (N_19799,N_18466,N_18078);
or U19800 (N_19800,N_18513,N_18311);
or U19801 (N_19801,N_18578,N_18667);
nand U19802 (N_19802,N_18582,N_18637);
nand U19803 (N_19803,N_18091,N_18847);
and U19804 (N_19804,N_18494,N_18035);
or U19805 (N_19805,N_18039,N_18631);
xor U19806 (N_19806,N_18799,N_18266);
nand U19807 (N_19807,N_18414,N_18388);
nor U19808 (N_19808,N_18247,N_18165);
nand U19809 (N_19809,N_18567,N_18405);
xnor U19810 (N_19810,N_18289,N_18889);
or U19811 (N_19811,N_18059,N_18153);
and U19812 (N_19812,N_18578,N_18717);
nor U19813 (N_19813,N_18445,N_18046);
nand U19814 (N_19814,N_18315,N_18974);
nor U19815 (N_19815,N_18268,N_18271);
xnor U19816 (N_19816,N_18453,N_18151);
nand U19817 (N_19817,N_18654,N_18310);
xnor U19818 (N_19818,N_18440,N_18657);
nand U19819 (N_19819,N_18527,N_18474);
or U19820 (N_19820,N_18883,N_18148);
nor U19821 (N_19821,N_18147,N_18571);
xnor U19822 (N_19822,N_18397,N_18314);
nand U19823 (N_19823,N_18704,N_18985);
nor U19824 (N_19824,N_18700,N_18889);
xor U19825 (N_19825,N_18112,N_18608);
xor U19826 (N_19826,N_18499,N_18146);
or U19827 (N_19827,N_18784,N_18098);
xnor U19828 (N_19828,N_18061,N_18446);
nand U19829 (N_19829,N_18845,N_18074);
and U19830 (N_19830,N_18404,N_18892);
or U19831 (N_19831,N_18215,N_18500);
nor U19832 (N_19832,N_18697,N_18163);
nor U19833 (N_19833,N_18129,N_18918);
and U19834 (N_19834,N_18762,N_18081);
and U19835 (N_19835,N_18445,N_18928);
or U19836 (N_19836,N_18308,N_18788);
xnor U19837 (N_19837,N_18935,N_18709);
nand U19838 (N_19838,N_18184,N_18230);
nor U19839 (N_19839,N_18549,N_18916);
nand U19840 (N_19840,N_18347,N_18969);
xnor U19841 (N_19841,N_18371,N_18173);
nand U19842 (N_19842,N_18601,N_18776);
or U19843 (N_19843,N_18143,N_18636);
and U19844 (N_19844,N_18452,N_18428);
nor U19845 (N_19845,N_18220,N_18594);
or U19846 (N_19846,N_18837,N_18241);
nand U19847 (N_19847,N_18108,N_18349);
and U19848 (N_19848,N_18139,N_18063);
xor U19849 (N_19849,N_18635,N_18786);
xnor U19850 (N_19850,N_18589,N_18249);
or U19851 (N_19851,N_18642,N_18832);
and U19852 (N_19852,N_18565,N_18757);
nor U19853 (N_19853,N_18614,N_18634);
or U19854 (N_19854,N_18356,N_18421);
nand U19855 (N_19855,N_18826,N_18357);
or U19856 (N_19856,N_18598,N_18234);
or U19857 (N_19857,N_18218,N_18764);
or U19858 (N_19858,N_18355,N_18722);
or U19859 (N_19859,N_18013,N_18005);
and U19860 (N_19860,N_18087,N_18049);
xnor U19861 (N_19861,N_18662,N_18676);
xor U19862 (N_19862,N_18718,N_18286);
or U19863 (N_19863,N_18589,N_18210);
and U19864 (N_19864,N_18978,N_18609);
or U19865 (N_19865,N_18598,N_18198);
nand U19866 (N_19866,N_18544,N_18624);
nand U19867 (N_19867,N_18771,N_18396);
nand U19868 (N_19868,N_18920,N_18493);
xor U19869 (N_19869,N_18813,N_18898);
xnor U19870 (N_19870,N_18661,N_18644);
xnor U19871 (N_19871,N_18142,N_18388);
xnor U19872 (N_19872,N_18586,N_18280);
nor U19873 (N_19873,N_18378,N_18565);
xor U19874 (N_19874,N_18790,N_18723);
or U19875 (N_19875,N_18041,N_18970);
nor U19876 (N_19876,N_18137,N_18125);
nand U19877 (N_19877,N_18002,N_18314);
or U19878 (N_19878,N_18311,N_18059);
nand U19879 (N_19879,N_18936,N_18179);
or U19880 (N_19880,N_18246,N_18014);
xnor U19881 (N_19881,N_18317,N_18372);
and U19882 (N_19882,N_18606,N_18846);
xor U19883 (N_19883,N_18823,N_18470);
or U19884 (N_19884,N_18153,N_18660);
nand U19885 (N_19885,N_18346,N_18102);
xor U19886 (N_19886,N_18846,N_18695);
and U19887 (N_19887,N_18403,N_18807);
and U19888 (N_19888,N_18001,N_18500);
and U19889 (N_19889,N_18648,N_18757);
nand U19890 (N_19890,N_18390,N_18601);
or U19891 (N_19891,N_18497,N_18693);
nand U19892 (N_19892,N_18141,N_18922);
and U19893 (N_19893,N_18657,N_18333);
nor U19894 (N_19894,N_18882,N_18470);
nand U19895 (N_19895,N_18391,N_18499);
nand U19896 (N_19896,N_18700,N_18270);
or U19897 (N_19897,N_18416,N_18183);
and U19898 (N_19898,N_18023,N_18591);
nor U19899 (N_19899,N_18580,N_18645);
and U19900 (N_19900,N_18869,N_18487);
or U19901 (N_19901,N_18372,N_18723);
or U19902 (N_19902,N_18704,N_18022);
and U19903 (N_19903,N_18224,N_18591);
or U19904 (N_19904,N_18392,N_18273);
or U19905 (N_19905,N_18038,N_18822);
and U19906 (N_19906,N_18962,N_18893);
nor U19907 (N_19907,N_18344,N_18319);
nand U19908 (N_19908,N_18518,N_18637);
nand U19909 (N_19909,N_18424,N_18998);
xnor U19910 (N_19910,N_18321,N_18651);
nand U19911 (N_19911,N_18554,N_18141);
nor U19912 (N_19912,N_18573,N_18402);
nand U19913 (N_19913,N_18821,N_18455);
nor U19914 (N_19914,N_18016,N_18116);
nand U19915 (N_19915,N_18694,N_18000);
xnor U19916 (N_19916,N_18171,N_18691);
and U19917 (N_19917,N_18288,N_18701);
nor U19918 (N_19918,N_18724,N_18765);
or U19919 (N_19919,N_18325,N_18570);
or U19920 (N_19920,N_18612,N_18021);
nand U19921 (N_19921,N_18433,N_18088);
or U19922 (N_19922,N_18357,N_18720);
nand U19923 (N_19923,N_18381,N_18400);
xor U19924 (N_19924,N_18754,N_18954);
nand U19925 (N_19925,N_18495,N_18384);
xnor U19926 (N_19926,N_18935,N_18391);
and U19927 (N_19927,N_18753,N_18897);
xor U19928 (N_19928,N_18892,N_18623);
or U19929 (N_19929,N_18159,N_18765);
nor U19930 (N_19930,N_18811,N_18162);
nand U19931 (N_19931,N_18315,N_18792);
nand U19932 (N_19932,N_18987,N_18751);
or U19933 (N_19933,N_18383,N_18604);
and U19934 (N_19934,N_18623,N_18540);
nor U19935 (N_19935,N_18127,N_18485);
and U19936 (N_19936,N_18550,N_18025);
and U19937 (N_19937,N_18538,N_18561);
nand U19938 (N_19938,N_18842,N_18787);
nand U19939 (N_19939,N_18228,N_18269);
or U19940 (N_19940,N_18643,N_18836);
nand U19941 (N_19941,N_18993,N_18457);
and U19942 (N_19942,N_18998,N_18354);
nor U19943 (N_19943,N_18334,N_18659);
or U19944 (N_19944,N_18451,N_18139);
or U19945 (N_19945,N_18915,N_18540);
nand U19946 (N_19946,N_18609,N_18524);
nor U19947 (N_19947,N_18720,N_18448);
nor U19948 (N_19948,N_18254,N_18677);
and U19949 (N_19949,N_18915,N_18193);
xnor U19950 (N_19950,N_18441,N_18564);
and U19951 (N_19951,N_18002,N_18546);
xnor U19952 (N_19952,N_18934,N_18554);
or U19953 (N_19953,N_18455,N_18277);
xor U19954 (N_19954,N_18467,N_18571);
xnor U19955 (N_19955,N_18408,N_18164);
nor U19956 (N_19956,N_18423,N_18609);
or U19957 (N_19957,N_18331,N_18231);
nand U19958 (N_19958,N_18955,N_18119);
nor U19959 (N_19959,N_18140,N_18114);
xnor U19960 (N_19960,N_18428,N_18269);
nor U19961 (N_19961,N_18441,N_18509);
or U19962 (N_19962,N_18977,N_18187);
xnor U19963 (N_19963,N_18509,N_18596);
or U19964 (N_19964,N_18312,N_18372);
xnor U19965 (N_19965,N_18329,N_18017);
and U19966 (N_19966,N_18586,N_18324);
or U19967 (N_19967,N_18059,N_18363);
xnor U19968 (N_19968,N_18628,N_18816);
and U19969 (N_19969,N_18694,N_18266);
nor U19970 (N_19970,N_18334,N_18388);
xnor U19971 (N_19971,N_18030,N_18113);
nor U19972 (N_19972,N_18697,N_18288);
or U19973 (N_19973,N_18460,N_18085);
or U19974 (N_19974,N_18821,N_18946);
nand U19975 (N_19975,N_18781,N_18506);
xor U19976 (N_19976,N_18809,N_18009);
xor U19977 (N_19977,N_18453,N_18397);
nand U19978 (N_19978,N_18139,N_18495);
nor U19979 (N_19979,N_18904,N_18675);
xnor U19980 (N_19980,N_18810,N_18877);
and U19981 (N_19981,N_18490,N_18399);
nor U19982 (N_19982,N_18823,N_18491);
or U19983 (N_19983,N_18864,N_18660);
or U19984 (N_19984,N_18035,N_18582);
and U19985 (N_19985,N_18556,N_18876);
xnor U19986 (N_19986,N_18789,N_18338);
nand U19987 (N_19987,N_18651,N_18878);
or U19988 (N_19988,N_18510,N_18985);
nand U19989 (N_19989,N_18234,N_18833);
or U19990 (N_19990,N_18223,N_18433);
and U19991 (N_19991,N_18793,N_18558);
nand U19992 (N_19992,N_18881,N_18296);
nand U19993 (N_19993,N_18595,N_18101);
and U19994 (N_19994,N_18735,N_18666);
nor U19995 (N_19995,N_18905,N_18087);
nand U19996 (N_19996,N_18090,N_18295);
nor U19997 (N_19997,N_18213,N_18069);
xnor U19998 (N_19998,N_18578,N_18851);
xor U19999 (N_19999,N_18934,N_18731);
nand U20000 (N_20000,N_19820,N_19171);
or U20001 (N_20001,N_19695,N_19004);
xnor U20002 (N_20002,N_19288,N_19808);
and U20003 (N_20003,N_19365,N_19603);
nor U20004 (N_20004,N_19879,N_19095);
xor U20005 (N_20005,N_19576,N_19577);
nor U20006 (N_20006,N_19940,N_19180);
and U20007 (N_20007,N_19671,N_19342);
and U20008 (N_20008,N_19875,N_19587);
nand U20009 (N_20009,N_19255,N_19588);
nor U20010 (N_20010,N_19298,N_19832);
nor U20011 (N_20011,N_19308,N_19607);
nand U20012 (N_20012,N_19640,N_19903);
xor U20013 (N_20013,N_19391,N_19211);
xnor U20014 (N_20014,N_19685,N_19407);
nor U20015 (N_20015,N_19451,N_19977);
xnor U20016 (N_20016,N_19434,N_19793);
and U20017 (N_20017,N_19060,N_19559);
xor U20018 (N_20018,N_19411,N_19684);
and U20019 (N_20019,N_19333,N_19268);
xnor U20020 (N_20020,N_19639,N_19030);
or U20021 (N_20021,N_19872,N_19345);
and U20022 (N_20022,N_19387,N_19353);
and U20023 (N_20023,N_19601,N_19259);
nand U20024 (N_20024,N_19652,N_19773);
and U20025 (N_20025,N_19711,N_19961);
and U20026 (N_20026,N_19332,N_19074);
and U20027 (N_20027,N_19433,N_19683);
nand U20028 (N_20028,N_19924,N_19141);
xnor U20029 (N_20029,N_19462,N_19878);
xor U20030 (N_20030,N_19756,N_19835);
or U20031 (N_20031,N_19973,N_19656);
xor U20032 (N_20032,N_19529,N_19312);
nor U20033 (N_20033,N_19173,N_19057);
nand U20034 (N_20034,N_19943,N_19783);
nand U20035 (N_20035,N_19976,N_19406);
nand U20036 (N_20036,N_19599,N_19665);
nand U20037 (N_20037,N_19472,N_19292);
or U20038 (N_20038,N_19625,N_19690);
nor U20039 (N_20039,N_19956,N_19351);
nand U20040 (N_20040,N_19612,N_19539);
nand U20041 (N_20041,N_19889,N_19618);
nor U20042 (N_20042,N_19944,N_19410);
or U20043 (N_20043,N_19987,N_19922);
xnor U20044 (N_20044,N_19465,N_19809);
and U20045 (N_20045,N_19494,N_19150);
nor U20046 (N_20046,N_19957,N_19827);
nand U20047 (N_20047,N_19281,N_19771);
or U20048 (N_20048,N_19525,N_19646);
and U20049 (N_20049,N_19311,N_19779);
and U20050 (N_20050,N_19796,N_19048);
nor U20051 (N_20051,N_19081,N_19517);
xor U20052 (N_20052,N_19191,N_19340);
or U20053 (N_20053,N_19269,N_19226);
and U20054 (N_20054,N_19923,N_19825);
xor U20055 (N_20055,N_19833,N_19675);
xnor U20056 (N_20056,N_19421,N_19329);
or U20057 (N_20057,N_19915,N_19155);
nand U20058 (N_20058,N_19196,N_19495);
nor U20059 (N_20059,N_19129,N_19642);
xor U20060 (N_20060,N_19659,N_19500);
xor U20061 (N_20061,N_19737,N_19159);
nor U20062 (N_20062,N_19454,N_19181);
xor U20063 (N_20063,N_19749,N_19726);
xnor U20064 (N_20064,N_19860,N_19846);
xnor U20065 (N_20065,N_19845,N_19664);
nor U20066 (N_20066,N_19810,N_19381);
nor U20067 (N_20067,N_19869,N_19934);
nor U20068 (N_20068,N_19105,N_19997);
nand U20069 (N_20069,N_19611,N_19724);
or U20070 (N_20070,N_19775,N_19578);
or U20071 (N_20071,N_19859,N_19140);
nor U20072 (N_20072,N_19346,N_19350);
xor U20073 (N_20073,N_19195,N_19532);
xnor U20074 (N_20074,N_19236,N_19026);
nor U20075 (N_20075,N_19948,N_19398);
or U20076 (N_20076,N_19101,N_19955);
and U20077 (N_20077,N_19117,N_19349);
nand U20078 (N_20078,N_19186,N_19044);
or U20079 (N_20079,N_19297,N_19723);
nor U20080 (N_20080,N_19914,N_19718);
nand U20081 (N_20081,N_19187,N_19228);
nor U20082 (N_20082,N_19457,N_19324);
and U20083 (N_20083,N_19466,N_19999);
or U20084 (N_20084,N_19676,N_19490);
and U20085 (N_20085,N_19772,N_19207);
nand U20086 (N_20086,N_19686,N_19609);
nor U20087 (N_20087,N_19289,N_19029);
or U20088 (N_20088,N_19214,N_19250);
nand U20089 (N_20089,N_19082,N_19784);
xor U20090 (N_20090,N_19931,N_19476);
xnor U20091 (N_20091,N_19864,N_19215);
and U20092 (N_20092,N_19307,N_19232);
or U20093 (N_20093,N_19036,N_19927);
and U20094 (N_20094,N_19261,N_19326);
and U20095 (N_20095,N_19224,N_19636);
or U20096 (N_20096,N_19005,N_19011);
nand U20097 (N_20097,N_19699,N_19156);
nand U20098 (N_20098,N_19870,N_19902);
nand U20099 (N_20099,N_19777,N_19506);
xnor U20100 (N_20100,N_19189,N_19192);
nor U20101 (N_20101,N_19469,N_19803);
nor U20102 (N_20102,N_19774,N_19418);
nor U20103 (N_20103,N_19020,N_19453);
nor U20104 (N_20104,N_19897,N_19496);
xnor U20105 (N_20105,N_19507,N_19364);
nand U20106 (N_20106,N_19790,N_19648);
xor U20107 (N_20107,N_19780,N_19763);
and U20108 (N_20108,N_19691,N_19840);
xor U20109 (N_20109,N_19730,N_19965);
or U20110 (N_20110,N_19358,N_19000);
xnor U20111 (N_20111,N_19304,N_19866);
nand U20112 (N_20112,N_19092,N_19982);
xnor U20113 (N_20113,N_19834,N_19217);
nor U20114 (N_20114,N_19432,N_19574);
nand U20115 (N_20115,N_19899,N_19714);
nor U20116 (N_20116,N_19641,N_19637);
xor U20117 (N_20117,N_19753,N_19460);
nand U20118 (N_20118,N_19971,N_19594);
and U20119 (N_20119,N_19791,N_19645);
nor U20120 (N_20120,N_19331,N_19850);
or U20121 (N_20121,N_19185,N_19152);
xnor U20122 (N_20122,N_19049,N_19626);
or U20123 (N_20123,N_19527,N_19100);
xnor U20124 (N_20124,N_19830,N_19284);
or U20125 (N_20125,N_19585,N_19119);
or U20126 (N_20126,N_19919,N_19814);
and U20127 (N_20127,N_19440,N_19857);
nor U20128 (N_20128,N_19168,N_19447);
and U20129 (N_20129,N_19019,N_19680);
nor U20130 (N_20130,N_19430,N_19888);
nand U20131 (N_20131,N_19498,N_19868);
nor U20132 (N_20132,N_19776,N_19689);
xnor U20133 (N_20133,N_19727,N_19424);
and U20134 (N_20134,N_19535,N_19522);
or U20135 (N_20135,N_19627,N_19589);
and U20136 (N_20136,N_19437,N_19426);
nand U20137 (N_20137,N_19383,N_19681);
nand U20138 (N_20138,N_19120,N_19677);
and U20139 (N_20139,N_19634,N_19041);
or U20140 (N_20140,N_19423,N_19974);
nor U20141 (N_20141,N_19414,N_19293);
and U20142 (N_20142,N_19070,N_19372);
xnor U20143 (N_20143,N_19144,N_19134);
or U20144 (N_20144,N_19415,N_19564);
nor U20145 (N_20145,N_19488,N_19438);
xor U20146 (N_20146,N_19028,N_19463);
and U20147 (N_20147,N_19752,N_19039);
and U20148 (N_20148,N_19738,N_19993);
or U20149 (N_20149,N_19499,N_19382);
nor U20150 (N_20150,N_19706,N_19988);
nor U20151 (N_20151,N_19761,N_19524);
nand U20152 (N_20152,N_19533,N_19658);
or U20153 (N_20153,N_19170,N_19911);
xnor U20154 (N_20154,N_19205,N_19076);
nand U20155 (N_20155,N_19489,N_19768);
and U20156 (N_20156,N_19201,N_19059);
nand U20157 (N_20157,N_19317,N_19449);
nand U20158 (N_20158,N_19190,N_19528);
and U20159 (N_20159,N_19595,N_19565);
nor U20160 (N_20160,N_19265,N_19256);
and U20161 (N_20161,N_19286,N_19045);
xnor U20162 (N_20162,N_19184,N_19571);
nor U20163 (N_20163,N_19649,N_19876);
nor U20164 (N_20164,N_19344,N_19767);
or U20165 (N_20165,N_19778,N_19492);
xor U20166 (N_20166,N_19886,N_19693);
and U20167 (N_20167,N_19073,N_19586);
or U20168 (N_20168,N_19741,N_19538);
or U20169 (N_20169,N_19669,N_19303);
nor U20170 (N_20170,N_19994,N_19946);
and U20171 (N_20171,N_19839,N_19550);
nand U20172 (N_20172,N_19202,N_19253);
xnor U20173 (N_20173,N_19003,N_19952);
nor U20174 (N_20174,N_19133,N_19836);
xor U20175 (N_20175,N_19580,N_19031);
xnor U20176 (N_20176,N_19852,N_19657);
xnor U20177 (N_20177,N_19816,N_19408);
and U20178 (N_20178,N_19127,N_19318);
or U20179 (N_20179,N_19428,N_19285);
and U20180 (N_20180,N_19592,N_19557);
nor U20181 (N_20181,N_19234,N_19313);
and U20182 (N_20182,N_19483,N_19480);
nand U20183 (N_20183,N_19166,N_19046);
and U20184 (N_20184,N_19021,N_19194);
nand U20185 (N_20185,N_19370,N_19497);
nand U20186 (N_20186,N_19275,N_19853);
and U20187 (N_20187,N_19824,N_19015);
nor U20188 (N_20188,N_19945,N_19422);
nor U20189 (N_20189,N_19023,N_19481);
and U20190 (N_20190,N_19037,N_19396);
and U20191 (N_20191,N_19980,N_19139);
or U20192 (N_20192,N_19047,N_19416);
xnor U20193 (N_20193,N_19376,N_19663);
and U20194 (N_20194,N_19673,N_19950);
or U20195 (N_20195,N_19598,N_19176);
nand U20196 (N_20196,N_19717,N_19131);
or U20197 (N_20197,N_19198,N_19471);
nand U20198 (N_20198,N_19963,N_19958);
or U20199 (N_20199,N_19062,N_19251);
and U20200 (N_20200,N_19633,N_19065);
and U20201 (N_20201,N_19622,N_19504);
or U20202 (N_20202,N_19066,N_19766);
nor U20203 (N_20203,N_19068,N_19855);
nand U20204 (N_20204,N_19179,N_19002);
xor U20205 (N_20205,N_19355,N_19912);
xor U20206 (N_20206,N_19951,N_19709);
and U20207 (N_20207,N_19838,N_19802);
xor U20208 (N_20208,N_19368,N_19010);
nor U20209 (N_20209,N_19485,N_19754);
nor U20210 (N_20210,N_19896,N_19223);
or U20211 (N_20211,N_19321,N_19518);
or U20212 (N_20212,N_19847,N_19510);
and U20213 (N_20213,N_19990,N_19918);
xnor U20214 (N_20214,N_19443,N_19509);
or U20215 (N_20215,N_19932,N_19162);
xnor U20216 (N_20216,N_19404,N_19731);
xnor U20217 (N_20217,N_19165,N_19747);
xnor U20218 (N_20218,N_19556,N_19482);
and U20219 (N_20219,N_19380,N_19083);
nand U20220 (N_20220,N_19635,N_19632);
nand U20221 (N_20221,N_19064,N_19096);
or U20222 (N_20222,N_19540,N_19969);
nand U20223 (N_20223,N_19456,N_19939);
nor U20224 (N_20224,N_19319,N_19757);
nor U20225 (N_20225,N_19904,N_19962);
nor U20226 (N_20226,N_19605,N_19563);
and U20227 (N_20227,N_19008,N_19093);
nand U20228 (N_20228,N_19937,N_19992);
and U20229 (N_20229,N_19638,N_19474);
nor U20230 (N_20230,N_19475,N_19617);
or U20231 (N_20231,N_19821,N_19792);
or U20232 (N_20232,N_19526,N_19405);
nand U20233 (N_20233,N_19051,N_19579);
nor U20234 (N_20234,N_19241,N_19862);
and U20235 (N_20235,N_19341,N_19245);
and U20236 (N_20236,N_19826,N_19890);
nand U20237 (N_20237,N_19278,N_19998);
nand U20238 (N_20238,N_19042,N_19549);
nand U20239 (N_20239,N_19644,N_19570);
nor U20240 (N_20240,N_19177,N_19666);
nor U20241 (N_20241,N_19104,N_19544);
xnor U20242 (N_20242,N_19745,N_19620);
nand U20243 (N_20243,N_19043,N_19335);
and U20244 (N_20244,N_19450,N_19735);
xor U20245 (N_20245,N_19569,N_19392);
or U20246 (N_20246,N_19995,N_19744);
nand U20247 (N_20247,N_19885,N_19197);
or U20248 (N_20248,N_19694,N_19258);
and U20249 (N_20249,N_19295,N_19328);
or U20250 (N_20250,N_19327,N_19271);
nand U20251 (N_20251,N_19390,N_19551);
or U20252 (N_20252,N_19097,N_19800);
nor U20253 (N_20253,N_19698,N_19722);
xnor U20254 (N_20254,N_19893,N_19877);
or U20255 (N_20255,N_19545,N_19696);
and U20256 (N_20256,N_19079,N_19356);
nor U20257 (N_20257,N_19283,N_19486);
or U20258 (N_20258,N_19983,N_19027);
and U20259 (N_20259,N_19464,N_19736);
or U20260 (N_20260,N_19600,N_19759);
xnor U20261 (N_20261,N_19025,N_19291);
or U20262 (N_20262,N_19032,N_19334);
nand U20263 (N_20263,N_19098,N_19263);
nand U20264 (N_20264,N_19145,N_19616);
nor U20265 (N_20265,N_19901,N_19262);
or U20266 (N_20266,N_19455,N_19220);
nand U20267 (N_20267,N_19523,N_19970);
and U20268 (N_20268,N_19908,N_19913);
and U20269 (N_20269,N_19831,N_19050);
nor U20270 (N_20270,N_19764,N_19209);
or U20271 (N_20271,N_19887,N_19512);
or U20272 (N_20272,N_19363,N_19541);
xor U20273 (N_20273,N_19608,N_19403);
xnor U20274 (N_20274,N_19861,N_19389);
nor U20275 (N_20275,N_19158,N_19765);
and U20276 (N_20276,N_19906,N_19084);
or U20277 (N_20277,N_19339,N_19536);
nand U20278 (N_20278,N_19781,N_19558);
nor U20279 (N_20279,N_19619,N_19397);
or U20280 (N_20280,N_19959,N_19703);
nand U20281 (N_20281,N_19441,N_19732);
or U20282 (N_20282,N_19935,N_19841);
xor U20283 (N_20283,N_19981,N_19146);
and U20284 (N_20284,N_19280,N_19966);
nor U20285 (N_20285,N_19360,N_19909);
nand U20286 (N_20286,N_19697,N_19077);
xnor U20287 (N_20287,N_19710,N_19290);
nor U20288 (N_20288,N_19199,N_19247);
xor U20289 (N_20289,N_19124,N_19222);
nand U20290 (N_20290,N_19725,N_19844);
and U20291 (N_20291,N_19055,N_19530);
xor U20292 (N_20292,N_19301,N_19229);
nor U20293 (N_20293,N_19034,N_19933);
xnor U20294 (N_20294,N_19679,N_19798);
or U20295 (N_20295,N_19881,N_19548);
or U20296 (N_20296,N_19604,N_19277);
or U20297 (N_20297,N_19056,N_19322);
nor U20298 (N_20298,N_19110,N_19760);
xor U20299 (N_20299,N_19367,N_19797);
nand U20300 (N_20300,N_19954,N_19273);
or U20301 (N_20301,N_19085,N_19435);
xnor U20302 (N_20302,N_19248,N_19299);
and U20303 (N_20303,N_19149,N_19115);
nor U20304 (N_20304,N_19856,N_19660);
nor U20305 (N_20305,N_19871,N_19508);
nand U20306 (N_20306,N_19964,N_19947);
and U20307 (N_20307,N_19305,N_19514);
and U20308 (N_20308,N_19148,N_19702);
nand U20309 (N_20309,N_19038,N_19593);
nand U20310 (N_20310,N_19910,N_19806);
nor U20311 (N_20311,N_19921,N_19114);
and U20312 (N_20312,N_19748,N_19596);
or U20313 (N_20313,N_19621,N_19366);
or U20314 (N_20314,N_19606,N_19431);
or U20315 (N_20315,N_19459,N_19385);
or U20316 (N_20316,N_19087,N_19552);
nor U20317 (N_20317,N_19058,N_19054);
or U20318 (N_20318,N_19624,N_19672);
or U20319 (N_20319,N_19078,N_19799);
or U20320 (N_20320,N_19602,N_19704);
or U20321 (N_20321,N_19720,N_19033);
or U20322 (N_20322,N_19427,N_19795);
or U20323 (N_20323,N_19707,N_19178);
or U20324 (N_20324,N_19219,N_19701);
and U20325 (N_20325,N_19719,N_19547);
and U20326 (N_20326,N_19941,N_19337);
and U20327 (N_20327,N_19928,N_19022);
and U20328 (N_20328,N_19183,N_19505);
nor U20329 (N_20329,N_19819,N_19487);
nor U20330 (N_20330,N_19244,N_19172);
xor U20331 (N_20331,N_19786,N_19828);
nor U20332 (N_20332,N_19531,N_19984);
nand U20333 (N_20333,N_19746,N_19436);
or U20334 (N_20334,N_19743,N_19788);
nand U20335 (N_20335,N_19823,N_19972);
xor U20336 (N_20336,N_19560,N_19789);
and U20337 (N_20337,N_19213,N_19597);
xnor U20338 (N_20338,N_19402,N_19705);
nor U20339 (N_20339,N_19154,N_19001);
nor U20340 (N_20340,N_19478,N_19583);
and U20341 (N_20341,N_19369,N_19409);
nor U20342 (N_20342,N_19543,N_19296);
nor U20343 (N_20343,N_19968,N_19667);
nand U20344 (N_20344,N_19413,N_19257);
and U20345 (N_20345,N_19929,N_19384);
nor U20346 (N_20346,N_19713,N_19315);
nand U20347 (N_20347,N_19160,N_19949);
or U20348 (N_20348,N_19700,N_19442);
and U20349 (N_20349,N_19135,N_19534);
and U20350 (N_20350,N_19867,N_19762);
and U20351 (N_20351,N_19287,N_19212);
xnor U20352 (N_20352,N_19661,N_19237);
and U20353 (N_20353,N_19208,N_19581);
xor U20354 (N_20354,N_19960,N_19357);
nand U20355 (N_20355,N_19916,N_19643);
nand U20356 (N_20356,N_19310,N_19264);
or U20357 (N_20357,N_19818,N_19573);
nor U20358 (N_20358,N_19647,N_19006);
nand U20359 (N_20359,N_19446,N_19515);
xor U20360 (N_20360,N_19206,N_19132);
nor U20361 (N_20361,N_19467,N_19118);
nor U20362 (N_20362,N_19582,N_19254);
nand U20363 (N_20363,N_19650,N_19069);
nor U20364 (N_20364,N_19425,N_19572);
and U20365 (N_20365,N_19246,N_19142);
xor U20366 (N_20366,N_19352,N_19610);
or U20367 (N_20367,N_19204,N_19343);
and U20368 (N_20368,N_19138,N_19323);
xor U20369 (N_20369,N_19468,N_19815);
nand U20370 (N_20370,N_19546,N_19182);
nand U20371 (N_20371,N_19294,N_19188);
nor U20372 (N_20372,N_19614,N_19668);
nand U20373 (N_20373,N_19272,N_19979);
nor U20374 (N_20374,N_19123,N_19121);
and U20375 (N_20375,N_19018,N_19309);
nor U20376 (N_20376,N_19394,N_19444);
nand U20377 (N_20377,N_19143,N_19099);
nor U20378 (N_20378,N_19225,N_19883);
xnor U20379 (N_20379,N_19655,N_19942);
xor U20380 (N_20380,N_19270,N_19874);
and U20381 (N_20381,N_19109,N_19674);
xor U20382 (N_20382,N_19537,N_19053);
nand U20383 (N_20383,N_19067,N_19300);
nor U20384 (N_20384,N_19898,N_19016);
xnor U20385 (N_20385,N_19362,N_19623);
or U20386 (N_20386,N_19811,N_19112);
nor U20387 (N_20387,N_19511,N_19439);
xnor U20388 (N_20388,N_19107,N_19233);
and U20389 (N_20389,N_19061,N_19375);
nand U20390 (N_20390,N_19210,N_19203);
nor U20391 (N_20391,N_19785,N_19395);
or U20392 (N_20392,N_19715,N_19477);
or U20393 (N_20393,N_19473,N_19555);
and U20394 (N_20394,N_19266,N_19348);
xor U20395 (N_20395,N_19071,N_19420);
nor U20396 (N_20396,N_19801,N_19917);
nor U20397 (N_20397,N_19721,N_19651);
nor U20398 (N_20398,N_19519,N_19111);
nand U20399 (N_20399,N_19063,N_19035);
nor U20400 (N_20400,N_19843,N_19920);
and U20401 (N_20401,N_19895,N_19670);
xnor U20402 (N_20402,N_19386,N_19848);
nor U20403 (N_20403,N_19448,N_19267);
nand U20404 (N_20404,N_19314,N_19822);
nand U20405 (N_20405,N_19812,N_19967);
and U20406 (N_20406,N_19193,N_19106);
nand U20407 (N_20407,N_19491,N_19770);
nand U20408 (N_20408,N_19520,N_19086);
and U20409 (N_20409,N_19130,N_19751);
or U20410 (N_20410,N_19938,N_19227);
nand U20411 (N_20411,N_19975,N_19758);
and U20412 (N_20412,N_19175,N_19470);
nor U20413 (N_20413,N_19230,N_19240);
and U20414 (N_20414,N_19678,N_19513);
nor U20415 (N_20415,N_19122,N_19837);
xnor U20416 (N_20416,N_19553,N_19040);
xor U20417 (N_20417,N_19854,N_19052);
nand U20418 (N_20418,N_19167,N_19359);
nand U20419 (N_20419,N_19782,N_19399);
or U20420 (N_20420,N_19169,N_19249);
xnor U20421 (N_20421,N_19014,N_19484);
nand U20422 (N_20422,N_19930,N_19989);
nand U20423 (N_20423,N_19007,N_19379);
nand U20424 (N_20424,N_19401,N_19502);
nor U20425 (N_20425,N_19371,N_19089);
nand U20426 (N_20426,N_19075,N_19103);
and U20427 (N_20427,N_19147,N_19017);
nand U20428 (N_20428,N_19174,N_19137);
and U20429 (N_20429,N_19688,N_19996);
and U20430 (N_20430,N_19161,N_19242);
xnor U20431 (N_20431,N_19562,N_19412);
xnor U20432 (N_20432,N_19126,N_19164);
or U20433 (N_20433,N_19687,N_19692);
or U20434 (N_20434,N_19728,N_19128);
nor U20435 (N_20435,N_19012,N_19094);
nand U20436 (N_20436,N_19231,N_19306);
nand U20437 (N_20437,N_19566,N_19716);
nand U20438 (N_20438,N_19884,N_19088);
nor U20439 (N_20439,N_19009,N_19794);
nand U20440 (N_20440,N_19252,N_19378);
xnor U20441 (N_20441,N_19157,N_19336);
nand U20442 (N_20442,N_19458,N_19892);
nand U20443 (N_20443,N_19151,N_19316);
or U20444 (N_20444,N_19108,N_19804);
nand U20445 (N_20445,N_19153,N_19393);
nor U20446 (N_20446,N_19863,N_19953);
and U20447 (N_20447,N_19080,N_19136);
and U20448 (N_20448,N_19813,N_19493);
nor U20449 (N_20449,N_19842,N_19873);
nand U20450 (N_20450,N_19417,N_19712);
xor U20451 (N_20451,N_19260,N_19851);
nor U20452 (N_20452,N_19388,N_19739);
and U20453 (N_20453,N_19653,N_19373);
or U20454 (N_20454,N_19554,N_19628);
xor U20455 (N_20455,N_19091,N_19239);
nor U20456 (N_20456,N_19429,N_19200);
and U20457 (N_20457,N_19013,N_19361);
nor U20458 (N_20458,N_19102,N_19907);
nand U20459 (N_20459,N_19805,N_19750);
and U20460 (N_20460,N_19561,N_19461);
or U20461 (N_20461,N_19354,N_19116);
nor U20462 (N_20462,N_19880,N_19279);
and U20463 (N_20463,N_19445,N_19787);
nand U20464 (N_20464,N_19320,N_19905);
and U20465 (N_20465,N_19024,N_19567);
nor U20466 (N_20466,N_19936,N_19733);
nor U20467 (N_20467,N_19991,N_19891);
or U20468 (N_20468,N_19817,N_19986);
nand U20469 (N_20469,N_19542,N_19734);
nor U20470 (N_20470,N_19925,N_19330);
or U20471 (N_20471,N_19682,N_19829);
or U20472 (N_20472,N_19613,N_19274);
nand U20473 (N_20473,N_19708,N_19568);
nor U20474 (N_20474,N_19374,N_19629);
xnor U20475 (N_20475,N_19419,N_19479);
nand U20476 (N_20476,N_19377,N_19325);
and U20477 (N_20477,N_19894,N_19882);
nor U20478 (N_20478,N_19113,N_19163);
or U20479 (N_20479,N_19243,N_19926);
and U20480 (N_20480,N_19221,N_19858);
xnor U20481 (N_20481,N_19865,N_19740);
and U20482 (N_20482,N_19985,N_19516);
nand U20483 (N_20483,N_19400,N_19090);
nor U20484 (N_20484,N_19347,N_19662);
nand U20485 (N_20485,N_19584,N_19978);
or U20486 (N_20486,N_19769,N_19590);
xor U20487 (N_20487,N_19521,N_19742);
or U20488 (N_20488,N_19235,N_19631);
nand U20489 (N_20489,N_19503,N_19900);
nand U20490 (N_20490,N_19591,N_19216);
nor U20491 (N_20491,N_19630,N_19125);
nand U20492 (N_20492,N_19654,N_19575);
xor U20493 (N_20493,N_19501,N_19338);
or U20494 (N_20494,N_19755,N_19615);
and U20495 (N_20495,N_19302,N_19849);
xor U20496 (N_20496,N_19072,N_19807);
and U20497 (N_20497,N_19218,N_19729);
or U20498 (N_20498,N_19282,N_19276);
xor U20499 (N_20499,N_19238,N_19452);
and U20500 (N_20500,N_19942,N_19285);
or U20501 (N_20501,N_19804,N_19906);
nand U20502 (N_20502,N_19220,N_19795);
and U20503 (N_20503,N_19060,N_19499);
nand U20504 (N_20504,N_19528,N_19088);
nor U20505 (N_20505,N_19483,N_19801);
and U20506 (N_20506,N_19414,N_19271);
and U20507 (N_20507,N_19922,N_19610);
xor U20508 (N_20508,N_19921,N_19528);
nor U20509 (N_20509,N_19148,N_19962);
nand U20510 (N_20510,N_19709,N_19765);
xnor U20511 (N_20511,N_19105,N_19592);
xnor U20512 (N_20512,N_19873,N_19768);
or U20513 (N_20513,N_19136,N_19801);
and U20514 (N_20514,N_19479,N_19636);
xnor U20515 (N_20515,N_19694,N_19002);
nand U20516 (N_20516,N_19450,N_19376);
xnor U20517 (N_20517,N_19091,N_19590);
nor U20518 (N_20518,N_19687,N_19536);
or U20519 (N_20519,N_19455,N_19521);
and U20520 (N_20520,N_19211,N_19536);
and U20521 (N_20521,N_19821,N_19016);
and U20522 (N_20522,N_19808,N_19737);
nor U20523 (N_20523,N_19358,N_19139);
and U20524 (N_20524,N_19122,N_19063);
or U20525 (N_20525,N_19930,N_19702);
xnor U20526 (N_20526,N_19319,N_19711);
or U20527 (N_20527,N_19367,N_19662);
nor U20528 (N_20528,N_19841,N_19165);
xor U20529 (N_20529,N_19071,N_19351);
and U20530 (N_20530,N_19682,N_19083);
and U20531 (N_20531,N_19258,N_19016);
nand U20532 (N_20532,N_19247,N_19867);
nor U20533 (N_20533,N_19445,N_19500);
or U20534 (N_20534,N_19874,N_19722);
nand U20535 (N_20535,N_19809,N_19996);
or U20536 (N_20536,N_19246,N_19495);
nor U20537 (N_20537,N_19953,N_19307);
nor U20538 (N_20538,N_19746,N_19739);
or U20539 (N_20539,N_19308,N_19658);
and U20540 (N_20540,N_19457,N_19361);
xor U20541 (N_20541,N_19533,N_19173);
nor U20542 (N_20542,N_19039,N_19135);
nor U20543 (N_20543,N_19740,N_19080);
nor U20544 (N_20544,N_19223,N_19937);
nand U20545 (N_20545,N_19110,N_19856);
and U20546 (N_20546,N_19893,N_19277);
or U20547 (N_20547,N_19199,N_19139);
and U20548 (N_20548,N_19144,N_19986);
xor U20549 (N_20549,N_19613,N_19169);
nand U20550 (N_20550,N_19310,N_19917);
nand U20551 (N_20551,N_19599,N_19384);
nor U20552 (N_20552,N_19468,N_19153);
nor U20553 (N_20553,N_19976,N_19140);
or U20554 (N_20554,N_19464,N_19134);
or U20555 (N_20555,N_19393,N_19523);
and U20556 (N_20556,N_19457,N_19407);
and U20557 (N_20557,N_19529,N_19141);
xor U20558 (N_20558,N_19145,N_19165);
and U20559 (N_20559,N_19080,N_19420);
nor U20560 (N_20560,N_19849,N_19074);
or U20561 (N_20561,N_19095,N_19085);
or U20562 (N_20562,N_19890,N_19559);
or U20563 (N_20563,N_19452,N_19894);
nand U20564 (N_20564,N_19150,N_19716);
and U20565 (N_20565,N_19645,N_19279);
xor U20566 (N_20566,N_19462,N_19095);
nor U20567 (N_20567,N_19900,N_19617);
and U20568 (N_20568,N_19095,N_19826);
nand U20569 (N_20569,N_19322,N_19966);
nand U20570 (N_20570,N_19034,N_19631);
and U20571 (N_20571,N_19608,N_19829);
nand U20572 (N_20572,N_19986,N_19565);
xnor U20573 (N_20573,N_19137,N_19290);
or U20574 (N_20574,N_19625,N_19148);
xor U20575 (N_20575,N_19282,N_19238);
nand U20576 (N_20576,N_19239,N_19352);
nand U20577 (N_20577,N_19637,N_19460);
and U20578 (N_20578,N_19480,N_19788);
nand U20579 (N_20579,N_19429,N_19341);
nand U20580 (N_20580,N_19119,N_19804);
xor U20581 (N_20581,N_19724,N_19555);
nor U20582 (N_20582,N_19006,N_19738);
nor U20583 (N_20583,N_19882,N_19014);
or U20584 (N_20584,N_19057,N_19577);
and U20585 (N_20585,N_19376,N_19074);
or U20586 (N_20586,N_19477,N_19590);
nand U20587 (N_20587,N_19194,N_19947);
or U20588 (N_20588,N_19202,N_19446);
or U20589 (N_20589,N_19639,N_19923);
nor U20590 (N_20590,N_19759,N_19554);
and U20591 (N_20591,N_19372,N_19514);
xnor U20592 (N_20592,N_19954,N_19939);
or U20593 (N_20593,N_19712,N_19500);
nand U20594 (N_20594,N_19731,N_19744);
xor U20595 (N_20595,N_19517,N_19149);
xor U20596 (N_20596,N_19119,N_19124);
nor U20597 (N_20597,N_19680,N_19883);
nand U20598 (N_20598,N_19728,N_19954);
and U20599 (N_20599,N_19831,N_19383);
and U20600 (N_20600,N_19572,N_19961);
xor U20601 (N_20601,N_19636,N_19910);
or U20602 (N_20602,N_19906,N_19708);
nor U20603 (N_20603,N_19375,N_19251);
or U20604 (N_20604,N_19022,N_19198);
nor U20605 (N_20605,N_19723,N_19755);
nor U20606 (N_20606,N_19683,N_19014);
or U20607 (N_20607,N_19308,N_19528);
nand U20608 (N_20608,N_19189,N_19525);
nor U20609 (N_20609,N_19005,N_19494);
nand U20610 (N_20610,N_19381,N_19674);
xor U20611 (N_20611,N_19693,N_19390);
and U20612 (N_20612,N_19023,N_19549);
or U20613 (N_20613,N_19886,N_19043);
nor U20614 (N_20614,N_19043,N_19801);
nand U20615 (N_20615,N_19070,N_19388);
nor U20616 (N_20616,N_19220,N_19282);
nand U20617 (N_20617,N_19768,N_19791);
and U20618 (N_20618,N_19097,N_19493);
xor U20619 (N_20619,N_19238,N_19376);
nand U20620 (N_20620,N_19417,N_19992);
and U20621 (N_20621,N_19799,N_19253);
xnor U20622 (N_20622,N_19565,N_19568);
nand U20623 (N_20623,N_19617,N_19313);
nor U20624 (N_20624,N_19636,N_19714);
or U20625 (N_20625,N_19402,N_19009);
or U20626 (N_20626,N_19888,N_19184);
nor U20627 (N_20627,N_19564,N_19493);
nor U20628 (N_20628,N_19757,N_19949);
xnor U20629 (N_20629,N_19572,N_19965);
nor U20630 (N_20630,N_19145,N_19079);
xnor U20631 (N_20631,N_19831,N_19536);
xnor U20632 (N_20632,N_19511,N_19217);
or U20633 (N_20633,N_19185,N_19527);
xor U20634 (N_20634,N_19511,N_19901);
nand U20635 (N_20635,N_19236,N_19709);
nor U20636 (N_20636,N_19502,N_19767);
nor U20637 (N_20637,N_19427,N_19660);
nand U20638 (N_20638,N_19565,N_19470);
nor U20639 (N_20639,N_19844,N_19305);
and U20640 (N_20640,N_19455,N_19791);
nor U20641 (N_20641,N_19293,N_19769);
nand U20642 (N_20642,N_19142,N_19275);
xnor U20643 (N_20643,N_19431,N_19332);
or U20644 (N_20644,N_19456,N_19034);
and U20645 (N_20645,N_19350,N_19134);
nand U20646 (N_20646,N_19030,N_19576);
or U20647 (N_20647,N_19081,N_19127);
nand U20648 (N_20648,N_19219,N_19949);
nand U20649 (N_20649,N_19780,N_19535);
xor U20650 (N_20650,N_19892,N_19694);
nor U20651 (N_20651,N_19766,N_19921);
or U20652 (N_20652,N_19670,N_19245);
xor U20653 (N_20653,N_19979,N_19639);
nor U20654 (N_20654,N_19838,N_19774);
nand U20655 (N_20655,N_19490,N_19855);
xor U20656 (N_20656,N_19714,N_19120);
nor U20657 (N_20657,N_19482,N_19017);
xor U20658 (N_20658,N_19786,N_19111);
nand U20659 (N_20659,N_19681,N_19107);
xnor U20660 (N_20660,N_19408,N_19308);
and U20661 (N_20661,N_19994,N_19716);
nor U20662 (N_20662,N_19844,N_19028);
nor U20663 (N_20663,N_19950,N_19010);
nor U20664 (N_20664,N_19180,N_19785);
or U20665 (N_20665,N_19803,N_19189);
nand U20666 (N_20666,N_19550,N_19504);
and U20667 (N_20667,N_19313,N_19591);
and U20668 (N_20668,N_19677,N_19524);
and U20669 (N_20669,N_19732,N_19521);
or U20670 (N_20670,N_19320,N_19935);
or U20671 (N_20671,N_19631,N_19314);
nand U20672 (N_20672,N_19112,N_19086);
nor U20673 (N_20673,N_19344,N_19419);
and U20674 (N_20674,N_19051,N_19787);
nor U20675 (N_20675,N_19397,N_19277);
and U20676 (N_20676,N_19148,N_19633);
and U20677 (N_20677,N_19151,N_19932);
and U20678 (N_20678,N_19104,N_19331);
nand U20679 (N_20679,N_19094,N_19892);
and U20680 (N_20680,N_19810,N_19184);
xnor U20681 (N_20681,N_19224,N_19062);
or U20682 (N_20682,N_19650,N_19176);
nand U20683 (N_20683,N_19205,N_19391);
nor U20684 (N_20684,N_19926,N_19577);
nor U20685 (N_20685,N_19054,N_19831);
or U20686 (N_20686,N_19822,N_19060);
or U20687 (N_20687,N_19080,N_19644);
or U20688 (N_20688,N_19497,N_19329);
xnor U20689 (N_20689,N_19704,N_19184);
nand U20690 (N_20690,N_19075,N_19878);
xnor U20691 (N_20691,N_19057,N_19059);
nand U20692 (N_20692,N_19947,N_19866);
or U20693 (N_20693,N_19882,N_19488);
xnor U20694 (N_20694,N_19833,N_19357);
nand U20695 (N_20695,N_19369,N_19264);
nor U20696 (N_20696,N_19988,N_19546);
nor U20697 (N_20697,N_19673,N_19946);
xnor U20698 (N_20698,N_19531,N_19639);
nor U20699 (N_20699,N_19670,N_19393);
nor U20700 (N_20700,N_19006,N_19245);
nor U20701 (N_20701,N_19715,N_19428);
xnor U20702 (N_20702,N_19993,N_19678);
nor U20703 (N_20703,N_19408,N_19806);
xnor U20704 (N_20704,N_19926,N_19542);
or U20705 (N_20705,N_19035,N_19174);
nand U20706 (N_20706,N_19587,N_19895);
or U20707 (N_20707,N_19637,N_19471);
and U20708 (N_20708,N_19355,N_19229);
nor U20709 (N_20709,N_19976,N_19128);
nor U20710 (N_20710,N_19051,N_19374);
xor U20711 (N_20711,N_19563,N_19224);
nand U20712 (N_20712,N_19756,N_19932);
xor U20713 (N_20713,N_19229,N_19058);
nand U20714 (N_20714,N_19043,N_19014);
nand U20715 (N_20715,N_19972,N_19392);
and U20716 (N_20716,N_19926,N_19483);
nand U20717 (N_20717,N_19100,N_19494);
nand U20718 (N_20718,N_19323,N_19435);
and U20719 (N_20719,N_19537,N_19244);
and U20720 (N_20720,N_19807,N_19098);
xor U20721 (N_20721,N_19139,N_19561);
and U20722 (N_20722,N_19711,N_19983);
xnor U20723 (N_20723,N_19233,N_19139);
nor U20724 (N_20724,N_19381,N_19270);
nand U20725 (N_20725,N_19629,N_19471);
nand U20726 (N_20726,N_19915,N_19593);
and U20727 (N_20727,N_19126,N_19697);
nor U20728 (N_20728,N_19349,N_19514);
and U20729 (N_20729,N_19129,N_19166);
and U20730 (N_20730,N_19684,N_19831);
xnor U20731 (N_20731,N_19064,N_19870);
nor U20732 (N_20732,N_19005,N_19332);
xor U20733 (N_20733,N_19775,N_19659);
nand U20734 (N_20734,N_19136,N_19908);
nand U20735 (N_20735,N_19641,N_19436);
or U20736 (N_20736,N_19959,N_19267);
or U20737 (N_20737,N_19441,N_19911);
and U20738 (N_20738,N_19337,N_19407);
nand U20739 (N_20739,N_19623,N_19191);
and U20740 (N_20740,N_19140,N_19384);
or U20741 (N_20741,N_19804,N_19714);
nand U20742 (N_20742,N_19753,N_19278);
xor U20743 (N_20743,N_19626,N_19569);
and U20744 (N_20744,N_19505,N_19596);
xnor U20745 (N_20745,N_19560,N_19708);
and U20746 (N_20746,N_19968,N_19406);
nor U20747 (N_20747,N_19368,N_19342);
nor U20748 (N_20748,N_19514,N_19839);
and U20749 (N_20749,N_19254,N_19422);
nor U20750 (N_20750,N_19637,N_19894);
and U20751 (N_20751,N_19189,N_19952);
xnor U20752 (N_20752,N_19517,N_19993);
and U20753 (N_20753,N_19796,N_19814);
nand U20754 (N_20754,N_19681,N_19621);
xnor U20755 (N_20755,N_19872,N_19357);
nand U20756 (N_20756,N_19545,N_19641);
and U20757 (N_20757,N_19859,N_19917);
nand U20758 (N_20758,N_19800,N_19776);
nand U20759 (N_20759,N_19541,N_19729);
nor U20760 (N_20760,N_19729,N_19644);
xnor U20761 (N_20761,N_19501,N_19158);
and U20762 (N_20762,N_19876,N_19309);
nand U20763 (N_20763,N_19862,N_19473);
and U20764 (N_20764,N_19779,N_19093);
xor U20765 (N_20765,N_19084,N_19193);
nand U20766 (N_20766,N_19643,N_19554);
xor U20767 (N_20767,N_19355,N_19091);
and U20768 (N_20768,N_19882,N_19001);
or U20769 (N_20769,N_19571,N_19498);
nand U20770 (N_20770,N_19480,N_19298);
xnor U20771 (N_20771,N_19795,N_19888);
or U20772 (N_20772,N_19227,N_19621);
or U20773 (N_20773,N_19824,N_19911);
nor U20774 (N_20774,N_19093,N_19298);
nor U20775 (N_20775,N_19334,N_19538);
nand U20776 (N_20776,N_19293,N_19134);
and U20777 (N_20777,N_19355,N_19781);
nand U20778 (N_20778,N_19569,N_19239);
and U20779 (N_20779,N_19399,N_19012);
nand U20780 (N_20780,N_19624,N_19997);
xor U20781 (N_20781,N_19420,N_19504);
or U20782 (N_20782,N_19944,N_19368);
nand U20783 (N_20783,N_19144,N_19063);
xnor U20784 (N_20784,N_19741,N_19687);
or U20785 (N_20785,N_19973,N_19892);
or U20786 (N_20786,N_19522,N_19778);
nand U20787 (N_20787,N_19425,N_19641);
and U20788 (N_20788,N_19453,N_19758);
nand U20789 (N_20789,N_19476,N_19937);
and U20790 (N_20790,N_19770,N_19284);
nor U20791 (N_20791,N_19202,N_19163);
nor U20792 (N_20792,N_19362,N_19435);
nor U20793 (N_20793,N_19046,N_19485);
and U20794 (N_20794,N_19358,N_19418);
and U20795 (N_20795,N_19285,N_19912);
xnor U20796 (N_20796,N_19576,N_19414);
nor U20797 (N_20797,N_19966,N_19257);
nand U20798 (N_20798,N_19937,N_19770);
nand U20799 (N_20799,N_19196,N_19729);
or U20800 (N_20800,N_19105,N_19366);
and U20801 (N_20801,N_19782,N_19029);
nand U20802 (N_20802,N_19020,N_19081);
nor U20803 (N_20803,N_19966,N_19049);
nand U20804 (N_20804,N_19597,N_19751);
xor U20805 (N_20805,N_19052,N_19566);
nor U20806 (N_20806,N_19019,N_19351);
or U20807 (N_20807,N_19552,N_19050);
xnor U20808 (N_20808,N_19003,N_19610);
nand U20809 (N_20809,N_19731,N_19194);
or U20810 (N_20810,N_19290,N_19802);
xnor U20811 (N_20811,N_19054,N_19173);
nand U20812 (N_20812,N_19794,N_19744);
or U20813 (N_20813,N_19905,N_19397);
or U20814 (N_20814,N_19096,N_19218);
and U20815 (N_20815,N_19230,N_19285);
nor U20816 (N_20816,N_19654,N_19947);
and U20817 (N_20817,N_19459,N_19678);
nor U20818 (N_20818,N_19668,N_19365);
nor U20819 (N_20819,N_19207,N_19503);
xor U20820 (N_20820,N_19671,N_19443);
nor U20821 (N_20821,N_19632,N_19899);
and U20822 (N_20822,N_19588,N_19544);
xnor U20823 (N_20823,N_19700,N_19514);
xor U20824 (N_20824,N_19711,N_19698);
nor U20825 (N_20825,N_19145,N_19840);
xor U20826 (N_20826,N_19824,N_19300);
or U20827 (N_20827,N_19066,N_19047);
nand U20828 (N_20828,N_19626,N_19903);
or U20829 (N_20829,N_19879,N_19373);
xnor U20830 (N_20830,N_19596,N_19209);
or U20831 (N_20831,N_19280,N_19012);
nand U20832 (N_20832,N_19759,N_19527);
xor U20833 (N_20833,N_19669,N_19654);
and U20834 (N_20834,N_19768,N_19197);
nand U20835 (N_20835,N_19833,N_19007);
xnor U20836 (N_20836,N_19940,N_19233);
or U20837 (N_20837,N_19762,N_19754);
xor U20838 (N_20838,N_19989,N_19835);
nand U20839 (N_20839,N_19982,N_19794);
nand U20840 (N_20840,N_19315,N_19001);
nor U20841 (N_20841,N_19468,N_19694);
or U20842 (N_20842,N_19619,N_19013);
nor U20843 (N_20843,N_19936,N_19330);
or U20844 (N_20844,N_19321,N_19909);
xor U20845 (N_20845,N_19999,N_19090);
or U20846 (N_20846,N_19880,N_19559);
xor U20847 (N_20847,N_19830,N_19778);
and U20848 (N_20848,N_19098,N_19899);
and U20849 (N_20849,N_19620,N_19265);
and U20850 (N_20850,N_19181,N_19922);
nand U20851 (N_20851,N_19217,N_19009);
nor U20852 (N_20852,N_19957,N_19636);
nor U20853 (N_20853,N_19005,N_19876);
xor U20854 (N_20854,N_19268,N_19594);
nand U20855 (N_20855,N_19456,N_19336);
and U20856 (N_20856,N_19040,N_19016);
nand U20857 (N_20857,N_19489,N_19754);
nor U20858 (N_20858,N_19061,N_19081);
xnor U20859 (N_20859,N_19460,N_19376);
nor U20860 (N_20860,N_19730,N_19139);
xor U20861 (N_20861,N_19119,N_19532);
and U20862 (N_20862,N_19326,N_19259);
nor U20863 (N_20863,N_19297,N_19015);
and U20864 (N_20864,N_19349,N_19059);
or U20865 (N_20865,N_19111,N_19041);
or U20866 (N_20866,N_19425,N_19865);
nand U20867 (N_20867,N_19122,N_19180);
nand U20868 (N_20868,N_19469,N_19008);
nand U20869 (N_20869,N_19613,N_19995);
or U20870 (N_20870,N_19807,N_19960);
nor U20871 (N_20871,N_19306,N_19822);
or U20872 (N_20872,N_19678,N_19026);
and U20873 (N_20873,N_19163,N_19523);
xnor U20874 (N_20874,N_19845,N_19263);
and U20875 (N_20875,N_19778,N_19380);
nand U20876 (N_20876,N_19638,N_19492);
nand U20877 (N_20877,N_19068,N_19367);
nor U20878 (N_20878,N_19984,N_19528);
or U20879 (N_20879,N_19016,N_19096);
nand U20880 (N_20880,N_19038,N_19941);
nor U20881 (N_20881,N_19797,N_19016);
or U20882 (N_20882,N_19677,N_19943);
nor U20883 (N_20883,N_19106,N_19631);
or U20884 (N_20884,N_19813,N_19225);
or U20885 (N_20885,N_19587,N_19987);
and U20886 (N_20886,N_19717,N_19573);
nand U20887 (N_20887,N_19923,N_19291);
nand U20888 (N_20888,N_19168,N_19951);
xnor U20889 (N_20889,N_19796,N_19265);
nand U20890 (N_20890,N_19624,N_19385);
nand U20891 (N_20891,N_19104,N_19598);
nand U20892 (N_20892,N_19637,N_19087);
and U20893 (N_20893,N_19490,N_19864);
nand U20894 (N_20894,N_19598,N_19809);
or U20895 (N_20895,N_19919,N_19452);
and U20896 (N_20896,N_19294,N_19768);
or U20897 (N_20897,N_19613,N_19437);
and U20898 (N_20898,N_19984,N_19718);
or U20899 (N_20899,N_19990,N_19871);
nand U20900 (N_20900,N_19891,N_19849);
nor U20901 (N_20901,N_19712,N_19208);
nand U20902 (N_20902,N_19949,N_19249);
xor U20903 (N_20903,N_19774,N_19456);
and U20904 (N_20904,N_19108,N_19868);
and U20905 (N_20905,N_19536,N_19220);
or U20906 (N_20906,N_19835,N_19912);
xnor U20907 (N_20907,N_19437,N_19655);
nand U20908 (N_20908,N_19655,N_19623);
xor U20909 (N_20909,N_19111,N_19067);
and U20910 (N_20910,N_19012,N_19361);
nor U20911 (N_20911,N_19092,N_19808);
or U20912 (N_20912,N_19507,N_19105);
nor U20913 (N_20913,N_19900,N_19613);
or U20914 (N_20914,N_19129,N_19340);
xnor U20915 (N_20915,N_19541,N_19396);
nand U20916 (N_20916,N_19699,N_19858);
nand U20917 (N_20917,N_19484,N_19385);
or U20918 (N_20918,N_19232,N_19727);
nand U20919 (N_20919,N_19494,N_19591);
nor U20920 (N_20920,N_19435,N_19567);
xor U20921 (N_20921,N_19073,N_19677);
xnor U20922 (N_20922,N_19729,N_19789);
and U20923 (N_20923,N_19374,N_19843);
nand U20924 (N_20924,N_19069,N_19531);
xor U20925 (N_20925,N_19959,N_19883);
xnor U20926 (N_20926,N_19375,N_19941);
xnor U20927 (N_20927,N_19711,N_19661);
nand U20928 (N_20928,N_19477,N_19208);
xnor U20929 (N_20929,N_19657,N_19465);
nand U20930 (N_20930,N_19978,N_19706);
xor U20931 (N_20931,N_19356,N_19005);
xnor U20932 (N_20932,N_19830,N_19607);
xnor U20933 (N_20933,N_19537,N_19731);
xnor U20934 (N_20934,N_19263,N_19015);
nor U20935 (N_20935,N_19999,N_19050);
nand U20936 (N_20936,N_19476,N_19587);
or U20937 (N_20937,N_19030,N_19607);
xor U20938 (N_20938,N_19516,N_19512);
or U20939 (N_20939,N_19839,N_19167);
and U20940 (N_20940,N_19453,N_19481);
or U20941 (N_20941,N_19630,N_19727);
nand U20942 (N_20942,N_19901,N_19950);
or U20943 (N_20943,N_19983,N_19523);
nand U20944 (N_20944,N_19343,N_19463);
or U20945 (N_20945,N_19081,N_19060);
nor U20946 (N_20946,N_19459,N_19554);
or U20947 (N_20947,N_19581,N_19152);
nand U20948 (N_20948,N_19310,N_19291);
and U20949 (N_20949,N_19231,N_19107);
nand U20950 (N_20950,N_19708,N_19086);
and U20951 (N_20951,N_19717,N_19740);
nand U20952 (N_20952,N_19140,N_19415);
or U20953 (N_20953,N_19703,N_19209);
and U20954 (N_20954,N_19980,N_19199);
and U20955 (N_20955,N_19152,N_19834);
and U20956 (N_20956,N_19528,N_19037);
nor U20957 (N_20957,N_19850,N_19036);
or U20958 (N_20958,N_19058,N_19359);
and U20959 (N_20959,N_19847,N_19243);
and U20960 (N_20960,N_19812,N_19332);
or U20961 (N_20961,N_19112,N_19696);
or U20962 (N_20962,N_19250,N_19427);
nor U20963 (N_20963,N_19762,N_19785);
xnor U20964 (N_20964,N_19341,N_19163);
xnor U20965 (N_20965,N_19667,N_19171);
or U20966 (N_20966,N_19999,N_19740);
or U20967 (N_20967,N_19685,N_19054);
nand U20968 (N_20968,N_19534,N_19109);
nor U20969 (N_20969,N_19074,N_19552);
or U20970 (N_20970,N_19719,N_19176);
nor U20971 (N_20971,N_19025,N_19500);
or U20972 (N_20972,N_19080,N_19116);
xnor U20973 (N_20973,N_19779,N_19983);
and U20974 (N_20974,N_19853,N_19335);
xnor U20975 (N_20975,N_19511,N_19756);
or U20976 (N_20976,N_19894,N_19942);
nand U20977 (N_20977,N_19311,N_19668);
nor U20978 (N_20978,N_19166,N_19636);
nand U20979 (N_20979,N_19469,N_19525);
xnor U20980 (N_20980,N_19504,N_19525);
or U20981 (N_20981,N_19895,N_19015);
xnor U20982 (N_20982,N_19772,N_19591);
or U20983 (N_20983,N_19355,N_19024);
and U20984 (N_20984,N_19583,N_19879);
and U20985 (N_20985,N_19160,N_19230);
and U20986 (N_20986,N_19202,N_19994);
and U20987 (N_20987,N_19628,N_19710);
nor U20988 (N_20988,N_19203,N_19037);
nand U20989 (N_20989,N_19480,N_19447);
nand U20990 (N_20990,N_19765,N_19467);
and U20991 (N_20991,N_19064,N_19083);
nand U20992 (N_20992,N_19913,N_19637);
and U20993 (N_20993,N_19453,N_19036);
or U20994 (N_20994,N_19849,N_19686);
nand U20995 (N_20995,N_19633,N_19194);
xnor U20996 (N_20996,N_19128,N_19291);
xor U20997 (N_20997,N_19217,N_19896);
nor U20998 (N_20998,N_19457,N_19247);
nand U20999 (N_20999,N_19799,N_19506);
nand U21000 (N_21000,N_20548,N_20567);
or U21001 (N_21001,N_20996,N_20038);
or U21002 (N_21002,N_20336,N_20977);
nor U21003 (N_21003,N_20769,N_20077);
or U21004 (N_21004,N_20464,N_20684);
or U21005 (N_21005,N_20795,N_20507);
nor U21006 (N_21006,N_20687,N_20782);
nand U21007 (N_21007,N_20579,N_20185);
or U21008 (N_21008,N_20367,N_20810);
xor U21009 (N_21009,N_20377,N_20941);
or U21010 (N_21010,N_20732,N_20125);
and U21011 (N_21011,N_20521,N_20851);
xnor U21012 (N_21012,N_20334,N_20702);
nor U21013 (N_21013,N_20499,N_20707);
nand U21014 (N_21014,N_20302,N_20820);
xnor U21015 (N_21015,N_20823,N_20969);
nor U21016 (N_21016,N_20379,N_20117);
xnor U21017 (N_21017,N_20994,N_20455);
nand U21018 (N_21018,N_20469,N_20554);
nand U21019 (N_21019,N_20420,N_20271);
or U21020 (N_21020,N_20793,N_20405);
xor U21021 (N_21021,N_20090,N_20219);
nand U21022 (N_21022,N_20743,N_20354);
xnor U21023 (N_21023,N_20510,N_20605);
or U21024 (N_21024,N_20116,N_20791);
nand U21025 (N_21025,N_20467,N_20488);
nor U21026 (N_21026,N_20589,N_20410);
nor U21027 (N_21027,N_20040,N_20056);
nand U21028 (N_21028,N_20193,N_20588);
nor U21029 (N_21029,N_20217,N_20475);
nor U21030 (N_21030,N_20574,N_20950);
or U21031 (N_21031,N_20258,N_20955);
or U21032 (N_21032,N_20847,N_20321);
and U21033 (N_21033,N_20300,N_20696);
nor U21034 (N_21034,N_20345,N_20122);
nor U21035 (N_21035,N_20834,N_20858);
and U21036 (N_21036,N_20067,N_20179);
nand U21037 (N_21037,N_20546,N_20590);
nor U21038 (N_21038,N_20340,N_20569);
nor U21039 (N_21039,N_20197,N_20722);
and U21040 (N_21040,N_20211,N_20873);
nand U21041 (N_21041,N_20493,N_20031);
and U21042 (N_21042,N_20511,N_20451);
nand U21043 (N_21043,N_20747,N_20572);
and U21044 (N_21044,N_20752,N_20233);
nand U21045 (N_21045,N_20418,N_20290);
and U21046 (N_21046,N_20070,N_20541);
xnor U21047 (N_21047,N_20656,N_20638);
or U21048 (N_21048,N_20839,N_20838);
and U21049 (N_21049,N_20074,N_20210);
xor U21050 (N_21050,N_20937,N_20706);
xnor U21051 (N_21051,N_20194,N_20093);
xor U21052 (N_21052,N_20331,N_20815);
nand U21053 (N_21053,N_20852,N_20776);
and U21054 (N_21054,N_20880,N_20928);
xnor U21055 (N_21055,N_20957,N_20781);
nand U21056 (N_21056,N_20974,N_20514);
nand U21057 (N_21057,N_20787,N_20057);
or U21058 (N_21058,N_20814,N_20385);
nand U21059 (N_21059,N_20693,N_20021);
and U21060 (N_21060,N_20384,N_20727);
xor U21061 (N_21061,N_20654,N_20601);
xnor U21062 (N_21062,N_20421,N_20319);
nand U21063 (N_21063,N_20476,N_20890);
and U21064 (N_21064,N_20128,N_20137);
nor U21065 (N_21065,N_20984,N_20886);
nor U21066 (N_21066,N_20450,N_20208);
xnor U21067 (N_21067,N_20425,N_20084);
xnor U21068 (N_21068,N_20049,N_20351);
xor U21069 (N_21069,N_20762,N_20527);
nor U21070 (N_21070,N_20529,N_20655);
nor U21071 (N_21071,N_20353,N_20885);
or U21072 (N_21072,N_20131,N_20364);
nor U21073 (N_21073,N_20501,N_20399);
xnor U21074 (N_21074,N_20494,N_20323);
nand U21075 (N_21075,N_20066,N_20254);
and U21076 (N_21076,N_20136,N_20901);
and U21077 (N_21077,N_20689,N_20540);
or U21078 (N_21078,N_20036,N_20698);
or U21079 (N_21079,N_20802,N_20874);
and U21080 (N_21080,N_20539,N_20436);
and U21081 (N_21081,N_20155,N_20573);
and U21082 (N_21082,N_20631,N_20526);
nand U21083 (N_21083,N_20267,N_20101);
and U21084 (N_21084,N_20860,N_20387);
nor U21085 (N_21085,N_20224,N_20045);
nor U21086 (N_21086,N_20766,N_20803);
nor U21087 (N_21087,N_20604,N_20568);
nor U21088 (N_21088,N_20456,N_20606);
xor U21089 (N_21089,N_20979,N_20751);
and U21090 (N_21090,N_20821,N_20327);
nand U21091 (N_21091,N_20800,N_20054);
and U21092 (N_21092,N_20047,N_20010);
and U21093 (N_21093,N_20775,N_20593);
or U21094 (N_21094,N_20028,N_20893);
and U21095 (N_21095,N_20404,N_20383);
nor U21096 (N_21096,N_20866,N_20665);
nor U21097 (N_21097,N_20152,N_20492);
and U21098 (N_21098,N_20431,N_20390);
nor U21099 (N_21099,N_20489,N_20059);
nor U21100 (N_21100,N_20462,N_20356);
xor U21101 (N_21101,N_20855,N_20711);
or U21102 (N_21102,N_20582,N_20615);
xor U21103 (N_21103,N_20720,N_20647);
nand U21104 (N_21104,N_20556,N_20204);
or U21105 (N_21105,N_20205,N_20177);
xor U21106 (N_21106,N_20448,N_20234);
or U21107 (N_21107,N_20934,N_20898);
and U21108 (N_21108,N_20381,N_20069);
nand U21109 (N_21109,N_20403,N_20457);
and U21110 (N_21110,N_20350,N_20240);
or U21111 (N_21111,N_20299,N_20932);
xor U21112 (N_21112,N_20679,N_20400);
nand U21113 (N_21113,N_20484,N_20549);
nand U21114 (N_21114,N_20491,N_20704);
nand U21115 (N_21115,N_20854,N_20623);
nand U21116 (N_21116,N_20006,N_20325);
xor U21117 (N_21117,N_20639,N_20285);
and U21118 (N_21118,N_20226,N_20044);
and U21119 (N_21119,N_20829,N_20482);
or U21120 (N_21120,N_20481,N_20386);
xor U21121 (N_21121,N_20102,N_20833);
or U21122 (N_21122,N_20915,N_20329);
and U21123 (N_21123,N_20107,N_20894);
or U21124 (N_21124,N_20311,N_20471);
or U21125 (N_21125,N_20146,N_20876);
and U21126 (N_21126,N_20912,N_20002);
or U21127 (N_21127,N_20767,N_20788);
and U21128 (N_21128,N_20671,N_20628);
or U21129 (N_21129,N_20291,N_20250);
xnor U21130 (N_21130,N_20328,N_20630);
nand U21131 (N_21131,N_20434,N_20342);
nand U21132 (N_21132,N_20598,N_20595);
xnor U21133 (N_21133,N_20423,N_20921);
nor U21134 (N_21134,N_20175,N_20729);
and U21135 (N_21135,N_20280,N_20708);
nand U21136 (N_21136,N_20092,N_20440);
nor U21137 (N_21137,N_20472,N_20053);
and U21138 (N_21138,N_20426,N_20566);
or U21139 (N_21139,N_20278,N_20292);
xnor U21140 (N_21140,N_20113,N_20786);
nand U21141 (N_21141,N_20919,N_20458);
nor U21142 (N_21142,N_20758,N_20168);
and U21143 (N_21143,N_20065,N_20121);
nand U21144 (N_21144,N_20214,N_20227);
or U21145 (N_21145,N_20678,N_20139);
xor U21146 (N_21146,N_20799,N_20369);
and U21147 (N_21147,N_20402,N_20145);
nand U21148 (N_21148,N_20252,N_20463);
nor U21149 (N_21149,N_20936,N_20277);
nor U21150 (N_21150,N_20674,N_20599);
or U21151 (N_21151,N_20393,N_20642);
or U21152 (N_21152,N_20373,N_20570);
or U21153 (N_21153,N_20024,N_20719);
or U21154 (N_21154,N_20844,N_20009);
nand U21155 (N_21155,N_20718,N_20673);
nor U21156 (N_21156,N_20602,N_20923);
nand U21157 (N_21157,N_20668,N_20878);
and U21158 (N_21158,N_20963,N_20949);
or U21159 (N_21159,N_20683,N_20978);
or U21160 (N_21160,N_20441,N_20358);
nand U21161 (N_21161,N_20999,N_20862);
nor U21162 (N_21162,N_20413,N_20594);
xor U21163 (N_21163,N_20407,N_20315);
and U21164 (N_21164,N_20600,N_20512);
xor U21165 (N_21165,N_20138,N_20657);
and U21166 (N_21166,N_20041,N_20135);
and U21167 (N_21167,N_20749,N_20253);
or U21168 (N_21168,N_20777,N_20812);
xnor U21169 (N_21169,N_20391,N_20691);
and U21170 (N_21170,N_20836,N_20734);
or U21171 (N_21171,N_20938,N_20905);
and U21172 (N_21172,N_20757,N_20889);
and U21173 (N_21173,N_20621,N_20150);
nand U21174 (N_21174,N_20430,N_20536);
nor U21175 (N_21175,N_20946,N_20360);
and U21176 (N_21176,N_20105,N_20365);
xor U21177 (N_21177,N_20653,N_20617);
or U21178 (N_21178,N_20465,N_20592);
nand U21179 (N_21179,N_20586,N_20332);
xnor U21180 (N_21180,N_20305,N_20337);
nor U21181 (N_21181,N_20532,N_20910);
or U21182 (N_21182,N_20538,N_20948);
nand U21183 (N_21183,N_20738,N_20147);
or U21184 (N_21184,N_20951,N_20826);
xnor U21185 (N_21185,N_20148,N_20761);
or U21186 (N_21186,N_20991,N_20731);
and U21187 (N_21187,N_20447,N_20075);
or U21188 (N_21188,N_20318,N_20944);
and U21189 (N_21189,N_20008,N_20670);
nor U21190 (N_21190,N_20875,N_20026);
nor U21191 (N_21191,N_20099,N_20163);
xnor U21192 (N_21192,N_20203,N_20658);
xnor U21193 (N_21193,N_20760,N_20675);
or U21194 (N_21194,N_20518,N_20645);
xnor U21195 (N_21195,N_20239,N_20713);
nor U21196 (N_21196,N_20106,N_20611);
nand U21197 (N_21197,N_20189,N_20230);
or U21198 (N_21198,N_20524,N_20322);
and U21199 (N_21199,N_20841,N_20634);
and U21200 (N_21200,N_20587,N_20603);
nor U21201 (N_21201,N_20162,N_20324);
nand U21202 (N_21202,N_20000,N_20772);
nor U21203 (N_21203,N_20966,N_20157);
nor U21204 (N_21204,N_20238,N_20103);
nor U21205 (N_21205,N_20953,N_20068);
or U21206 (N_21206,N_20971,N_20312);
nand U21207 (N_21207,N_20716,N_20335);
nand U21208 (N_21208,N_20914,N_20112);
or U21209 (N_21209,N_20468,N_20133);
or U21210 (N_21210,N_20520,N_20871);
xor U21211 (N_21211,N_20735,N_20960);
or U21212 (N_21212,N_20308,N_20543);
or U21213 (N_21213,N_20055,N_20073);
xnor U21214 (N_21214,N_20114,N_20768);
and U21215 (N_21215,N_20362,N_20161);
xor U21216 (N_21216,N_20246,N_20924);
nor U21217 (N_21217,N_20637,N_20376);
nand U21218 (N_21218,N_20187,N_20550);
xor U21219 (N_21219,N_20840,N_20895);
nor U21220 (N_21220,N_20109,N_20681);
and U21221 (N_21221,N_20142,N_20382);
nand U21222 (N_21222,N_20745,N_20268);
or U21223 (N_21223,N_20251,N_20730);
and U21224 (N_21224,N_20771,N_20432);
nor U21225 (N_21225,N_20740,N_20712);
nor U21226 (N_21226,N_20141,N_20857);
or U21227 (N_21227,N_20537,N_20888);
nand U21228 (N_21228,N_20863,N_20326);
nand U21229 (N_21229,N_20906,N_20629);
xnor U21230 (N_21230,N_20181,N_20294);
nand U21231 (N_21231,N_20095,N_20877);
xor U21232 (N_21232,N_20632,N_20682);
and U21233 (N_21233,N_20723,N_20371);
nor U21234 (N_21234,N_20968,N_20108);
nor U21235 (N_21235,N_20378,N_20981);
nor U21236 (N_21236,N_20506,N_20037);
or U21237 (N_21237,N_20939,N_20029);
nand U21238 (N_21238,N_20174,N_20742);
nor U21239 (N_21239,N_20864,N_20257);
or U21240 (N_21240,N_20933,N_20052);
nor U21241 (N_21241,N_20990,N_20962);
nor U21242 (N_21242,N_20433,N_20165);
nand U21243 (N_21243,N_20437,N_20050);
xnor U21244 (N_21244,N_20832,N_20296);
or U21245 (N_21245,N_20827,N_20307);
or U21246 (N_21246,N_20746,N_20245);
xnor U21247 (N_21247,N_20728,N_20672);
or U21248 (N_21248,N_20930,N_20553);
nand U21249 (N_21249,N_20361,N_20725);
nor U21250 (N_21250,N_20288,N_20581);
and U21251 (N_21251,N_20273,N_20804);
and U21252 (N_21252,N_20453,N_20947);
and U21253 (N_21253,N_20709,N_20229);
xnor U21254 (N_21254,N_20422,N_20835);
nand U21255 (N_21255,N_20692,N_20072);
and U21256 (N_21256,N_20993,N_20209);
or U21257 (N_21257,N_20446,N_20438);
nand U21258 (N_21258,N_20564,N_20313);
nor U21259 (N_21259,N_20794,N_20191);
xnor U21260 (N_21260,N_20242,N_20366);
xnor U21261 (N_21261,N_20547,N_20881);
or U21262 (N_21262,N_20259,N_20007);
xnor U21263 (N_21263,N_20184,N_20908);
nor U21264 (N_21264,N_20750,N_20223);
nor U21265 (N_21265,N_20435,N_20417);
and U21266 (N_21266,N_20079,N_20487);
nand U21267 (N_21267,N_20132,N_20640);
and U21268 (N_21268,N_20186,N_20355);
xor U21269 (N_21269,N_20477,N_20096);
xnor U21270 (N_21270,N_20452,N_20005);
or U21271 (N_21271,N_20973,N_20669);
nand U21272 (N_21272,N_20779,N_20967);
xor U21273 (N_21273,N_20166,N_20975);
or U21274 (N_21274,N_20498,N_20119);
xor U21275 (N_21275,N_20091,N_20347);
or U21276 (N_21276,N_20945,N_20571);
nor U21277 (N_21277,N_20522,N_20503);
xor U21278 (N_21278,N_20918,N_20062);
xor U21279 (N_21279,N_20202,N_20648);
and U21280 (N_21280,N_20517,N_20688);
nor U21281 (N_21281,N_20170,N_20797);
nand U21282 (N_21282,N_20169,N_20626);
xnor U21283 (N_21283,N_20160,N_20882);
and U21284 (N_21284,N_20561,N_20126);
or U21285 (N_21285,N_20042,N_20011);
nor U21286 (N_21286,N_20256,N_20035);
nand U21287 (N_21287,N_20609,N_20085);
and U21288 (N_21288,N_20001,N_20215);
and U21289 (N_21289,N_20198,N_20306);
nand U21290 (N_21290,N_20904,N_20232);
and U21291 (N_21291,N_20935,N_20736);
nor U21292 (N_21292,N_20111,N_20123);
nand U21293 (N_21293,N_20352,N_20992);
nand U21294 (N_21294,N_20544,N_20884);
or U21295 (N_21295,N_20705,N_20490);
xor U21296 (N_21296,N_20545,N_20798);
and U21297 (N_21297,N_20333,N_20183);
xor U21298 (N_21298,N_20172,N_20644);
and U21299 (N_21299,N_20428,N_20221);
xor U21300 (N_21300,N_20869,N_20703);
nand U21301 (N_21301,N_20865,N_20509);
nor U21302 (N_21302,N_20392,N_20811);
nand U21303 (N_21303,N_20666,N_20015);
and U21304 (N_21304,N_20954,N_20756);
xor U21305 (N_21305,N_20287,N_20585);
nor U21306 (N_21306,N_20303,N_20618);
nor U21307 (N_21307,N_20228,N_20359);
or U21308 (N_21308,N_20429,N_20159);
and U21309 (N_21309,N_20427,N_20997);
xnor U21310 (N_21310,N_20530,N_20043);
and U21311 (N_21311,N_20710,N_20976);
or U21312 (N_21312,N_20190,N_20098);
xor U21313 (N_21313,N_20927,N_20374);
nor U21314 (N_21314,N_20231,N_20260);
or U21315 (N_21315,N_20624,N_20531);
or U21316 (N_21316,N_20528,N_20870);
and U21317 (N_21317,N_20416,N_20902);
or U21318 (N_21318,N_20770,N_20596);
xor U21319 (N_21319,N_20619,N_20555);
and U21320 (N_21320,N_20891,N_20911);
or U21321 (N_21321,N_20580,N_20282);
nor U21322 (N_21322,N_20081,N_20479);
nor U21323 (N_21323,N_20087,N_20717);
xnor U21324 (N_21324,N_20807,N_20643);
nor U21325 (N_21325,N_20459,N_20398);
nand U21326 (N_21326,N_20620,N_20442);
xor U21327 (N_21327,N_20523,N_20357);
nor U21328 (N_21328,N_20241,N_20200);
or U21329 (N_21329,N_20505,N_20726);
or U21330 (N_21330,N_20247,N_20316);
xor U21331 (N_21331,N_20995,N_20088);
nor U21332 (N_21332,N_20922,N_20789);
nor U21333 (N_21333,N_20304,N_20542);
nand U21334 (N_21334,N_20926,N_20032);
nand U21335 (N_21335,N_20301,N_20310);
nand U21336 (N_21336,N_20389,N_20014);
nand U21337 (N_21337,N_20896,N_20480);
nand U21338 (N_21338,N_20048,N_20780);
and U21339 (N_21339,N_20641,N_20213);
and U21340 (N_21340,N_20064,N_20083);
nand U21341 (N_21341,N_20218,N_20485);
and U21342 (N_21342,N_20412,N_20676);
nand U21343 (N_21343,N_20608,N_20220);
and U21344 (N_21344,N_20023,N_20627);
nor U21345 (N_21345,N_20461,N_20843);
and U21346 (N_21346,N_20424,N_20754);
xor U21347 (N_21347,N_20249,N_20578);
and U21348 (N_21348,N_20338,N_20983);
nor U21349 (N_21349,N_20497,N_20610);
and U21350 (N_21350,N_20646,N_20764);
nand U21351 (N_21351,N_20279,N_20243);
nand U21352 (N_21352,N_20261,N_20685);
xor U21353 (N_21353,N_20346,N_20677);
xnor U21354 (N_21354,N_20842,N_20636);
xnor U21355 (N_21355,N_20818,N_20167);
xor U21356 (N_21356,N_20397,N_20956);
nand U21357 (N_21357,N_20225,N_20774);
xor U21358 (N_21358,N_20828,N_20845);
nor U21359 (N_21359,N_20649,N_20275);
and U21360 (N_21360,N_20368,N_20831);
or U21361 (N_21361,N_20853,N_20130);
nor U21362 (N_21362,N_20755,N_20408);
xnor U21363 (N_21363,N_20100,N_20003);
nor U21364 (N_21364,N_20721,N_20034);
nor U21365 (N_21365,N_20349,N_20824);
nor U21366 (N_21366,N_20583,N_20460);
or U21367 (N_21367,N_20917,N_20659);
and U21368 (N_21368,N_20748,N_20801);
nor U21369 (N_21369,N_20591,N_20439);
and U21370 (N_21370,N_20790,N_20110);
xor U21371 (N_21371,N_20662,N_20796);
and U21372 (N_21372,N_20124,N_20076);
or U21373 (N_21373,N_20201,N_20018);
nor U21374 (N_21374,N_20173,N_20715);
xnor U21375 (N_21375,N_20785,N_20848);
nand U21376 (N_21376,N_20348,N_20019);
nor U21377 (N_21377,N_20030,N_20650);
and U21378 (N_21378,N_20664,N_20892);
xnor U21379 (N_21379,N_20396,N_20080);
nand U21380 (N_21380,N_20900,N_20633);
xnor U21381 (N_21381,N_20017,N_20565);
xor U21382 (N_21382,N_20196,N_20989);
or U21383 (N_21383,N_20986,N_20699);
nor U21384 (N_21384,N_20533,N_20502);
xor U21385 (N_21385,N_20741,N_20613);
or U21386 (N_21386,N_20444,N_20559);
and U21387 (N_21387,N_20089,N_20262);
xnor U21388 (N_21388,N_20134,N_20737);
or U21389 (N_21389,N_20525,N_20972);
nor U21390 (N_21390,N_20816,N_20856);
or U21391 (N_21391,N_20394,N_20560);
nand U21392 (N_21392,N_20701,N_20140);
and U21393 (N_21393,N_20474,N_20033);
or U21394 (N_21394,N_20320,N_20663);
nand U21395 (N_21395,N_20607,N_20411);
or U21396 (N_21396,N_20817,N_20519);
nand U21397 (N_21397,N_20899,N_20276);
nand U21398 (N_21398,N_20920,N_20317);
nor U21399 (N_21399,N_20552,N_20942);
or U21400 (N_21400,N_20151,N_20199);
nor U21401 (N_21401,N_20809,N_20058);
nand U21402 (N_21402,N_20071,N_20515);
or U21403 (N_21403,N_20808,N_20763);
nor U21404 (N_21404,N_20255,N_20206);
or U21405 (N_21405,N_20516,N_20913);
and U21406 (N_21406,N_20907,N_20562);
xor U21407 (N_21407,N_20867,N_20264);
nor U21408 (N_21408,N_20660,N_20805);
nor U21409 (N_21409,N_20212,N_20861);
xnor U21410 (N_21410,N_20998,N_20961);
or U21411 (N_21411,N_20295,N_20284);
and U21412 (N_21412,N_20222,N_20272);
xor U21413 (N_21413,N_20143,N_20178);
nand U21414 (N_21414,N_20158,N_20897);
xnor U21415 (N_21415,N_20825,N_20192);
nor U21416 (N_21416,N_20931,N_20207);
nand U21417 (N_21417,N_20289,N_20164);
nand U21418 (N_21418,N_20120,N_20822);
or U21419 (N_21419,N_20753,N_20409);
and U21420 (N_21420,N_20739,N_20557);
xor U21421 (N_21421,N_20925,N_20176);
xor U21422 (N_21422,N_20104,N_20270);
nand U21423 (N_21423,N_20597,N_20235);
and U21424 (N_21424,N_20694,N_20063);
or U21425 (N_21425,N_20180,N_20286);
nand U21426 (N_21426,N_20443,N_20266);
xnor U21427 (N_21427,N_20395,N_20470);
nor U21428 (N_21428,N_20614,N_20248);
and U21429 (N_21429,N_20445,N_20985);
and U21430 (N_21430,N_20171,N_20269);
or U21431 (N_21431,N_20265,N_20958);
and U21432 (N_21432,N_20020,N_20388);
nand U21433 (N_21433,N_20733,N_20773);
xnor U21434 (N_21434,N_20027,N_20830);
xnor U21435 (N_21435,N_20535,N_20483);
nor U21436 (N_21436,N_20375,N_20667);
or U21437 (N_21437,N_20850,N_20622);
or U21438 (N_21438,N_20144,N_20903);
or U21439 (N_21439,N_20883,N_20466);
xor U21440 (N_21440,N_20980,N_20274);
or U21441 (N_21441,N_20082,N_20401);
nor U21442 (N_21442,N_20298,N_20486);
and U21443 (N_21443,N_20236,N_20652);
nand U21444 (N_21444,N_20025,N_20330);
nand U21445 (N_21445,N_20341,N_20577);
nand U21446 (N_21446,N_20988,N_20419);
nor U21447 (N_21447,N_20118,N_20495);
or U21448 (N_21448,N_20806,N_20868);
nand U21449 (N_21449,N_20690,N_20478);
xor U21450 (N_21450,N_20952,N_20454);
or U21451 (N_21451,N_20061,N_20013);
nor U21452 (N_21452,N_20612,N_20625);
or U21453 (N_21453,N_20778,N_20149);
or U21454 (N_21454,N_20513,N_20887);
nor U21455 (N_21455,N_20339,N_20022);
nor U21456 (N_21456,N_20046,N_20859);
and U21457 (N_21457,N_20680,N_20714);
and U21458 (N_21458,N_20344,N_20837);
or U21459 (N_21459,N_20982,N_20616);
and U21460 (N_21460,N_20415,N_20724);
nor U21461 (N_21461,N_20959,N_20263);
and U21462 (N_21462,N_20651,N_20759);
and U21463 (N_21463,N_20813,N_20216);
or U21464 (N_21464,N_20872,N_20293);
nand U21465 (N_21465,N_20765,N_20970);
and U21466 (N_21466,N_20244,N_20094);
and U21467 (N_21467,N_20584,N_20473);
or U21468 (N_21468,N_20363,N_20558);
or U21469 (N_21469,N_20695,N_20188);
nand U21470 (N_21470,N_20012,N_20406);
xor U21471 (N_21471,N_20496,N_20661);
nand U21472 (N_21472,N_20156,N_20060);
or U21473 (N_21473,N_20154,N_20504);
xnor U21474 (N_21474,N_20575,N_20283);
or U21475 (N_21475,N_20127,N_20879);
or U21476 (N_21476,N_20635,N_20309);
or U21477 (N_21477,N_20792,N_20097);
xor U21478 (N_21478,N_20004,N_20929);
nand U21479 (N_21479,N_20964,N_20697);
or U21480 (N_21480,N_20370,N_20297);
nor U21481 (N_21481,N_20237,N_20700);
xor U21482 (N_21482,N_20576,N_20051);
nand U21483 (N_21483,N_20372,N_20551);
xor U21484 (N_21484,N_20909,N_20449);
and U21485 (N_21485,N_20500,N_20534);
and U21486 (N_21486,N_20314,N_20849);
xor U21487 (N_21487,N_20039,N_20115);
nand U21488 (N_21488,N_20016,N_20078);
or U21489 (N_21489,N_20783,N_20129);
or U21490 (N_21490,N_20744,N_20281);
xor U21491 (N_21491,N_20343,N_20940);
xnor U21492 (N_21492,N_20508,N_20846);
nor U21493 (N_21493,N_20987,N_20086);
nand U21494 (N_21494,N_20943,N_20563);
nor U21495 (N_21495,N_20686,N_20414);
or U21496 (N_21496,N_20965,N_20380);
nand U21497 (N_21497,N_20784,N_20916);
nand U21498 (N_21498,N_20819,N_20153);
nand U21499 (N_21499,N_20195,N_20182);
nand U21500 (N_21500,N_20688,N_20027);
xor U21501 (N_21501,N_20768,N_20159);
or U21502 (N_21502,N_20865,N_20733);
or U21503 (N_21503,N_20971,N_20456);
xor U21504 (N_21504,N_20079,N_20492);
nor U21505 (N_21505,N_20552,N_20436);
nor U21506 (N_21506,N_20711,N_20863);
or U21507 (N_21507,N_20221,N_20929);
nor U21508 (N_21508,N_20564,N_20255);
or U21509 (N_21509,N_20593,N_20925);
and U21510 (N_21510,N_20484,N_20495);
nor U21511 (N_21511,N_20153,N_20706);
or U21512 (N_21512,N_20159,N_20319);
or U21513 (N_21513,N_20085,N_20280);
nor U21514 (N_21514,N_20403,N_20459);
or U21515 (N_21515,N_20937,N_20272);
and U21516 (N_21516,N_20020,N_20060);
xor U21517 (N_21517,N_20885,N_20981);
nand U21518 (N_21518,N_20623,N_20771);
xnor U21519 (N_21519,N_20099,N_20602);
nand U21520 (N_21520,N_20747,N_20897);
and U21521 (N_21521,N_20270,N_20872);
or U21522 (N_21522,N_20986,N_20889);
nor U21523 (N_21523,N_20208,N_20875);
and U21524 (N_21524,N_20792,N_20861);
nor U21525 (N_21525,N_20013,N_20771);
xor U21526 (N_21526,N_20852,N_20727);
or U21527 (N_21527,N_20487,N_20442);
and U21528 (N_21528,N_20311,N_20787);
nand U21529 (N_21529,N_20189,N_20978);
or U21530 (N_21530,N_20399,N_20370);
and U21531 (N_21531,N_20925,N_20012);
xnor U21532 (N_21532,N_20844,N_20296);
and U21533 (N_21533,N_20932,N_20884);
xor U21534 (N_21534,N_20113,N_20007);
nand U21535 (N_21535,N_20946,N_20351);
nand U21536 (N_21536,N_20472,N_20400);
xor U21537 (N_21537,N_20564,N_20208);
xor U21538 (N_21538,N_20467,N_20198);
xnor U21539 (N_21539,N_20042,N_20858);
or U21540 (N_21540,N_20493,N_20355);
nand U21541 (N_21541,N_20150,N_20365);
or U21542 (N_21542,N_20895,N_20040);
nand U21543 (N_21543,N_20501,N_20353);
nand U21544 (N_21544,N_20586,N_20612);
nand U21545 (N_21545,N_20022,N_20810);
or U21546 (N_21546,N_20642,N_20683);
nand U21547 (N_21547,N_20549,N_20724);
nand U21548 (N_21548,N_20326,N_20717);
and U21549 (N_21549,N_20761,N_20450);
nor U21550 (N_21550,N_20683,N_20811);
nand U21551 (N_21551,N_20161,N_20235);
or U21552 (N_21552,N_20083,N_20764);
or U21553 (N_21553,N_20913,N_20281);
or U21554 (N_21554,N_20295,N_20828);
nor U21555 (N_21555,N_20112,N_20123);
or U21556 (N_21556,N_20784,N_20030);
nand U21557 (N_21557,N_20796,N_20769);
nor U21558 (N_21558,N_20050,N_20665);
and U21559 (N_21559,N_20974,N_20680);
or U21560 (N_21560,N_20924,N_20737);
and U21561 (N_21561,N_20640,N_20030);
xor U21562 (N_21562,N_20539,N_20038);
nand U21563 (N_21563,N_20842,N_20918);
and U21564 (N_21564,N_20489,N_20699);
xnor U21565 (N_21565,N_20272,N_20675);
xor U21566 (N_21566,N_20248,N_20899);
xor U21567 (N_21567,N_20915,N_20062);
xor U21568 (N_21568,N_20661,N_20985);
and U21569 (N_21569,N_20150,N_20573);
nand U21570 (N_21570,N_20557,N_20105);
and U21571 (N_21571,N_20014,N_20010);
xnor U21572 (N_21572,N_20817,N_20923);
xnor U21573 (N_21573,N_20927,N_20359);
or U21574 (N_21574,N_20127,N_20003);
or U21575 (N_21575,N_20038,N_20055);
nor U21576 (N_21576,N_20160,N_20665);
nor U21577 (N_21577,N_20454,N_20534);
or U21578 (N_21578,N_20061,N_20182);
or U21579 (N_21579,N_20086,N_20615);
xnor U21580 (N_21580,N_20717,N_20460);
or U21581 (N_21581,N_20197,N_20209);
nand U21582 (N_21582,N_20001,N_20288);
or U21583 (N_21583,N_20752,N_20503);
or U21584 (N_21584,N_20226,N_20443);
and U21585 (N_21585,N_20921,N_20816);
and U21586 (N_21586,N_20875,N_20870);
and U21587 (N_21587,N_20666,N_20517);
xor U21588 (N_21588,N_20914,N_20674);
nor U21589 (N_21589,N_20194,N_20844);
nor U21590 (N_21590,N_20301,N_20592);
or U21591 (N_21591,N_20367,N_20168);
and U21592 (N_21592,N_20305,N_20153);
xor U21593 (N_21593,N_20204,N_20552);
xor U21594 (N_21594,N_20775,N_20926);
and U21595 (N_21595,N_20070,N_20420);
nand U21596 (N_21596,N_20010,N_20644);
xnor U21597 (N_21597,N_20669,N_20881);
xnor U21598 (N_21598,N_20747,N_20685);
xor U21599 (N_21599,N_20631,N_20150);
nor U21600 (N_21600,N_20475,N_20747);
or U21601 (N_21601,N_20959,N_20245);
xnor U21602 (N_21602,N_20289,N_20591);
or U21603 (N_21603,N_20459,N_20222);
or U21604 (N_21604,N_20095,N_20675);
nand U21605 (N_21605,N_20593,N_20245);
or U21606 (N_21606,N_20135,N_20204);
and U21607 (N_21607,N_20656,N_20508);
or U21608 (N_21608,N_20549,N_20730);
nand U21609 (N_21609,N_20185,N_20201);
xnor U21610 (N_21610,N_20577,N_20217);
and U21611 (N_21611,N_20023,N_20895);
or U21612 (N_21612,N_20783,N_20179);
or U21613 (N_21613,N_20915,N_20174);
or U21614 (N_21614,N_20822,N_20856);
nor U21615 (N_21615,N_20324,N_20635);
xnor U21616 (N_21616,N_20803,N_20708);
xor U21617 (N_21617,N_20446,N_20933);
nor U21618 (N_21618,N_20318,N_20728);
nor U21619 (N_21619,N_20222,N_20718);
xor U21620 (N_21620,N_20000,N_20144);
nor U21621 (N_21621,N_20474,N_20839);
nand U21622 (N_21622,N_20505,N_20395);
and U21623 (N_21623,N_20591,N_20139);
xnor U21624 (N_21624,N_20978,N_20404);
nor U21625 (N_21625,N_20500,N_20241);
nand U21626 (N_21626,N_20335,N_20167);
and U21627 (N_21627,N_20060,N_20043);
nor U21628 (N_21628,N_20112,N_20423);
and U21629 (N_21629,N_20825,N_20931);
nor U21630 (N_21630,N_20906,N_20333);
nor U21631 (N_21631,N_20165,N_20466);
xor U21632 (N_21632,N_20370,N_20832);
or U21633 (N_21633,N_20769,N_20531);
nand U21634 (N_21634,N_20419,N_20616);
and U21635 (N_21635,N_20335,N_20816);
nand U21636 (N_21636,N_20746,N_20765);
xor U21637 (N_21637,N_20592,N_20345);
and U21638 (N_21638,N_20783,N_20361);
or U21639 (N_21639,N_20042,N_20110);
and U21640 (N_21640,N_20767,N_20921);
nand U21641 (N_21641,N_20664,N_20632);
xnor U21642 (N_21642,N_20147,N_20768);
and U21643 (N_21643,N_20520,N_20609);
or U21644 (N_21644,N_20452,N_20668);
nor U21645 (N_21645,N_20529,N_20028);
and U21646 (N_21646,N_20508,N_20676);
nor U21647 (N_21647,N_20195,N_20933);
nand U21648 (N_21648,N_20636,N_20491);
and U21649 (N_21649,N_20818,N_20808);
and U21650 (N_21650,N_20240,N_20207);
and U21651 (N_21651,N_20048,N_20495);
and U21652 (N_21652,N_20774,N_20802);
or U21653 (N_21653,N_20230,N_20961);
nand U21654 (N_21654,N_20057,N_20952);
xor U21655 (N_21655,N_20947,N_20518);
and U21656 (N_21656,N_20495,N_20866);
nor U21657 (N_21657,N_20008,N_20912);
or U21658 (N_21658,N_20702,N_20659);
and U21659 (N_21659,N_20367,N_20067);
nor U21660 (N_21660,N_20744,N_20978);
and U21661 (N_21661,N_20998,N_20337);
xnor U21662 (N_21662,N_20791,N_20761);
and U21663 (N_21663,N_20038,N_20550);
or U21664 (N_21664,N_20297,N_20411);
and U21665 (N_21665,N_20527,N_20004);
and U21666 (N_21666,N_20473,N_20996);
nor U21667 (N_21667,N_20969,N_20055);
and U21668 (N_21668,N_20424,N_20284);
nand U21669 (N_21669,N_20322,N_20561);
or U21670 (N_21670,N_20973,N_20105);
nand U21671 (N_21671,N_20743,N_20738);
or U21672 (N_21672,N_20271,N_20943);
and U21673 (N_21673,N_20262,N_20942);
nand U21674 (N_21674,N_20957,N_20303);
and U21675 (N_21675,N_20762,N_20047);
xor U21676 (N_21676,N_20148,N_20136);
or U21677 (N_21677,N_20337,N_20527);
and U21678 (N_21678,N_20662,N_20989);
xor U21679 (N_21679,N_20309,N_20611);
or U21680 (N_21680,N_20563,N_20783);
nand U21681 (N_21681,N_20679,N_20654);
nand U21682 (N_21682,N_20224,N_20884);
or U21683 (N_21683,N_20363,N_20335);
nor U21684 (N_21684,N_20680,N_20313);
xor U21685 (N_21685,N_20463,N_20508);
nor U21686 (N_21686,N_20525,N_20935);
nand U21687 (N_21687,N_20603,N_20495);
xor U21688 (N_21688,N_20565,N_20896);
and U21689 (N_21689,N_20963,N_20593);
or U21690 (N_21690,N_20284,N_20534);
nor U21691 (N_21691,N_20886,N_20791);
and U21692 (N_21692,N_20806,N_20750);
and U21693 (N_21693,N_20429,N_20358);
nor U21694 (N_21694,N_20426,N_20099);
nor U21695 (N_21695,N_20220,N_20329);
and U21696 (N_21696,N_20994,N_20947);
nand U21697 (N_21697,N_20899,N_20868);
xnor U21698 (N_21698,N_20312,N_20354);
or U21699 (N_21699,N_20930,N_20925);
or U21700 (N_21700,N_20407,N_20782);
xor U21701 (N_21701,N_20059,N_20200);
nand U21702 (N_21702,N_20526,N_20900);
nand U21703 (N_21703,N_20755,N_20051);
xor U21704 (N_21704,N_20127,N_20932);
nor U21705 (N_21705,N_20889,N_20771);
nand U21706 (N_21706,N_20084,N_20732);
nor U21707 (N_21707,N_20990,N_20745);
and U21708 (N_21708,N_20508,N_20501);
and U21709 (N_21709,N_20684,N_20882);
or U21710 (N_21710,N_20046,N_20766);
or U21711 (N_21711,N_20532,N_20390);
nand U21712 (N_21712,N_20336,N_20746);
nor U21713 (N_21713,N_20531,N_20674);
or U21714 (N_21714,N_20764,N_20261);
nor U21715 (N_21715,N_20621,N_20726);
or U21716 (N_21716,N_20152,N_20089);
xnor U21717 (N_21717,N_20476,N_20426);
xnor U21718 (N_21718,N_20974,N_20865);
or U21719 (N_21719,N_20392,N_20213);
or U21720 (N_21720,N_20336,N_20973);
and U21721 (N_21721,N_20878,N_20227);
nand U21722 (N_21722,N_20606,N_20243);
or U21723 (N_21723,N_20018,N_20459);
nand U21724 (N_21724,N_20851,N_20259);
and U21725 (N_21725,N_20578,N_20867);
and U21726 (N_21726,N_20372,N_20053);
nor U21727 (N_21727,N_20887,N_20201);
and U21728 (N_21728,N_20250,N_20020);
nor U21729 (N_21729,N_20056,N_20542);
nor U21730 (N_21730,N_20272,N_20687);
nor U21731 (N_21731,N_20639,N_20565);
nor U21732 (N_21732,N_20585,N_20411);
and U21733 (N_21733,N_20843,N_20605);
nor U21734 (N_21734,N_20864,N_20070);
nand U21735 (N_21735,N_20060,N_20077);
xnor U21736 (N_21736,N_20676,N_20525);
xor U21737 (N_21737,N_20281,N_20984);
and U21738 (N_21738,N_20071,N_20250);
nor U21739 (N_21739,N_20864,N_20097);
or U21740 (N_21740,N_20590,N_20377);
nor U21741 (N_21741,N_20681,N_20175);
nand U21742 (N_21742,N_20111,N_20545);
xor U21743 (N_21743,N_20162,N_20545);
xnor U21744 (N_21744,N_20050,N_20508);
and U21745 (N_21745,N_20870,N_20307);
nor U21746 (N_21746,N_20253,N_20177);
nor U21747 (N_21747,N_20068,N_20954);
nand U21748 (N_21748,N_20225,N_20021);
xnor U21749 (N_21749,N_20664,N_20450);
or U21750 (N_21750,N_20052,N_20199);
nand U21751 (N_21751,N_20085,N_20441);
nand U21752 (N_21752,N_20356,N_20975);
or U21753 (N_21753,N_20902,N_20608);
nor U21754 (N_21754,N_20975,N_20174);
nand U21755 (N_21755,N_20641,N_20462);
xor U21756 (N_21756,N_20596,N_20009);
nand U21757 (N_21757,N_20657,N_20664);
or U21758 (N_21758,N_20988,N_20334);
xnor U21759 (N_21759,N_20599,N_20829);
nand U21760 (N_21760,N_20899,N_20528);
and U21761 (N_21761,N_20994,N_20507);
nand U21762 (N_21762,N_20302,N_20087);
nand U21763 (N_21763,N_20175,N_20130);
xnor U21764 (N_21764,N_20688,N_20362);
and U21765 (N_21765,N_20412,N_20347);
or U21766 (N_21766,N_20764,N_20961);
and U21767 (N_21767,N_20074,N_20816);
and U21768 (N_21768,N_20439,N_20253);
nand U21769 (N_21769,N_20545,N_20144);
nor U21770 (N_21770,N_20756,N_20584);
nor U21771 (N_21771,N_20005,N_20682);
and U21772 (N_21772,N_20238,N_20388);
nor U21773 (N_21773,N_20943,N_20065);
or U21774 (N_21774,N_20656,N_20465);
and U21775 (N_21775,N_20168,N_20745);
xor U21776 (N_21776,N_20823,N_20393);
or U21777 (N_21777,N_20007,N_20379);
and U21778 (N_21778,N_20151,N_20186);
and U21779 (N_21779,N_20213,N_20324);
and U21780 (N_21780,N_20618,N_20447);
xnor U21781 (N_21781,N_20946,N_20288);
xor U21782 (N_21782,N_20270,N_20940);
and U21783 (N_21783,N_20996,N_20166);
and U21784 (N_21784,N_20738,N_20753);
nor U21785 (N_21785,N_20222,N_20805);
xnor U21786 (N_21786,N_20223,N_20135);
or U21787 (N_21787,N_20299,N_20712);
and U21788 (N_21788,N_20267,N_20740);
and U21789 (N_21789,N_20351,N_20506);
xor U21790 (N_21790,N_20117,N_20533);
or U21791 (N_21791,N_20851,N_20195);
nor U21792 (N_21792,N_20559,N_20673);
or U21793 (N_21793,N_20019,N_20075);
or U21794 (N_21794,N_20842,N_20714);
or U21795 (N_21795,N_20137,N_20030);
or U21796 (N_21796,N_20658,N_20785);
xor U21797 (N_21797,N_20265,N_20493);
nor U21798 (N_21798,N_20057,N_20402);
nor U21799 (N_21799,N_20027,N_20070);
nor U21800 (N_21800,N_20877,N_20051);
xnor U21801 (N_21801,N_20805,N_20615);
nor U21802 (N_21802,N_20492,N_20122);
nand U21803 (N_21803,N_20977,N_20993);
xor U21804 (N_21804,N_20102,N_20059);
and U21805 (N_21805,N_20276,N_20976);
nand U21806 (N_21806,N_20774,N_20201);
or U21807 (N_21807,N_20881,N_20697);
or U21808 (N_21808,N_20649,N_20635);
and U21809 (N_21809,N_20474,N_20457);
and U21810 (N_21810,N_20651,N_20111);
and U21811 (N_21811,N_20632,N_20934);
and U21812 (N_21812,N_20739,N_20730);
nand U21813 (N_21813,N_20340,N_20306);
or U21814 (N_21814,N_20106,N_20757);
and U21815 (N_21815,N_20299,N_20972);
nor U21816 (N_21816,N_20631,N_20499);
and U21817 (N_21817,N_20486,N_20671);
nor U21818 (N_21818,N_20676,N_20938);
nor U21819 (N_21819,N_20520,N_20996);
xnor U21820 (N_21820,N_20738,N_20024);
and U21821 (N_21821,N_20263,N_20716);
nand U21822 (N_21822,N_20925,N_20765);
nor U21823 (N_21823,N_20175,N_20600);
nor U21824 (N_21824,N_20832,N_20474);
nand U21825 (N_21825,N_20567,N_20933);
nor U21826 (N_21826,N_20273,N_20178);
nor U21827 (N_21827,N_20145,N_20135);
nor U21828 (N_21828,N_20163,N_20749);
nor U21829 (N_21829,N_20156,N_20342);
and U21830 (N_21830,N_20289,N_20658);
or U21831 (N_21831,N_20572,N_20047);
nor U21832 (N_21832,N_20487,N_20871);
nand U21833 (N_21833,N_20923,N_20257);
or U21834 (N_21834,N_20980,N_20397);
and U21835 (N_21835,N_20349,N_20304);
or U21836 (N_21836,N_20985,N_20356);
nand U21837 (N_21837,N_20087,N_20704);
or U21838 (N_21838,N_20609,N_20692);
and U21839 (N_21839,N_20989,N_20500);
or U21840 (N_21840,N_20507,N_20103);
nand U21841 (N_21841,N_20753,N_20863);
and U21842 (N_21842,N_20101,N_20289);
xor U21843 (N_21843,N_20331,N_20883);
nor U21844 (N_21844,N_20383,N_20625);
and U21845 (N_21845,N_20634,N_20191);
or U21846 (N_21846,N_20230,N_20620);
xnor U21847 (N_21847,N_20871,N_20317);
and U21848 (N_21848,N_20507,N_20991);
nand U21849 (N_21849,N_20151,N_20581);
nand U21850 (N_21850,N_20744,N_20487);
and U21851 (N_21851,N_20722,N_20716);
nand U21852 (N_21852,N_20636,N_20137);
xor U21853 (N_21853,N_20213,N_20173);
nor U21854 (N_21854,N_20867,N_20267);
or U21855 (N_21855,N_20028,N_20422);
xor U21856 (N_21856,N_20083,N_20994);
xnor U21857 (N_21857,N_20093,N_20853);
or U21858 (N_21858,N_20077,N_20251);
and U21859 (N_21859,N_20240,N_20081);
and U21860 (N_21860,N_20860,N_20887);
and U21861 (N_21861,N_20197,N_20570);
or U21862 (N_21862,N_20606,N_20607);
xor U21863 (N_21863,N_20298,N_20557);
nor U21864 (N_21864,N_20616,N_20114);
xor U21865 (N_21865,N_20850,N_20489);
or U21866 (N_21866,N_20239,N_20952);
nand U21867 (N_21867,N_20104,N_20116);
nand U21868 (N_21868,N_20967,N_20213);
nor U21869 (N_21869,N_20041,N_20008);
nand U21870 (N_21870,N_20859,N_20321);
and U21871 (N_21871,N_20558,N_20042);
and U21872 (N_21872,N_20642,N_20415);
xor U21873 (N_21873,N_20908,N_20317);
xor U21874 (N_21874,N_20070,N_20898);
nor U21875 (N_21875,N_20872,N_20014);
nor U21876 (N_21876,N_20643,N_20064);
and U21877 (N_21877,N_20033,N_20792);
xnor U21878 (N_21878,N_20609,N_20989);
and U21879 (N_21879,N_20270,N_20032);
xnor U21880 (N_21880,N_20546,N_20210);
xor U21881 (N_21881,N_20399,N_20561);
xor U21882 (N_21882,N_20196,N_20928);
and U21883 (N_21883,N_20121,N_20961);
and U21884 (N_21884,N_20484,N_20325);
and U21885 (N_21885,N_20462,N_20029);
nor U21886 (N_21886,N_20915,N_20655);
xor U21887 (N_21887,N_20079,N_20889);
xor U21888 (N_21888,N_20772,N_20324);
and U21889 (N_21889,N_20842,N_20113);
xnor U21890 (N_21890,N_20446,N_20010);
nand U21891 (N_21891,N_20208,N_20510);
nand U21892 (N_21892,N_20880,N_20881);
nand U21893 (N_21893,N_20179,N_20072);
nor U21894 (N_21894,N_20467,N_20678);
or U21895 (N_21895,N_20421,N_20140);
nor U21896 (N_21896,N_20921,N_20701);
and U21897 (N_21897,N_20623,N_20885);
or U21898 (N_21898,N_20704,N_20412);
xnor U21899 (N_21899,N_20721,N_20664);
nand U21900 (N_21900,N_20040,N_20561);
xnor U21901 (N_21901,N_20763,N_20454);
or U21902 (N_21902,N_20419,N_20697);
and U21903 (N_21903,N_20619,N_20024);
nor U21904 (N_21904,N_20474,N_20899);
xor U21905 (N_21905,N_20795,N_20154);
and U21906 (N_21906,N_20031,N_20396);
nand U21907 (N_21907,N_20095,N_20199);
nor U21908 (N_21908,N_20201,N_20044);
nor U21909 (N_21909,N_20298,N_20311);
or U21910 (N_21910,N_20068,N_20222);
xnor U21911 (N_21911,N_20269,N_20668);
xor U21912 (N_21912,N_20861,N_20291);
or U21913 (N_21913,N_20056,N_20544);
or U21914 (N_21914,N_20700,N_20363);
nor U21915 (N_21915,N_20953,N_20066);
nor U21916 (N_21916,N_20181,N_20449);
xnor U21917 (N_21917,N_20036,N_20167);
nand U21918 (N_21918,N_20783,N_20809);
xnor U21919 (N_21919,N_20376,N_20813);
and U21920 (N_21920,N_20215,N_20245);
nor U21921 (N_21921,N_20782,N_20109);
nor U21922 (N_21922,N_20065,N_20401);
and U21923 (N_21923,N_20099,N_20324);
and U21924 (N_21924,N_20326,N_20394);
xor U21925 (N_21925,N_20526,N_20989);
xor U21926 (N_21926,N_20940,N_20919);
or U21927 (N_21927,N_20503,N_20760);
nor U21928 (N_21928,N_20390,N_20568);
nand U21929 (N_21929,N_20636,N_20939);
nor U21930 (N_21930,N_20386,N_20331);
or U21931 (N_21931,N_20235,N_20560);
or U21932 (N_21932,N_20673,N_20289);
and U21933 (N_21933,N_20253,N_20655);
nand U21934 (N_21934,N_20845,N_20559);
xnor U21935 (N_21935,N_20390,N_20198);
and U21936 (N_21936,N_20544,N_20665);
nand U21937 (N_21937,N_20528,N_20263);
xnor U21938 (N_21938,N_20243,N_20179);
and U21939 (N_21939,N_20516,N_20669);
or U21940 (N_21940,N_20732,N_20150);
nand U21941 (N_21941,N_20994,N_20515);
nand U21942 (N_21942,N_20962,N_20850);
or U21943 (N_21943,N_20096,N_20593);
nor U21944 (N_21944,N_20789,N_20036);
and U21945 (N_21945,N_20372,N_20562);
and U21946 (N_21946,N_20058,N_20244);
or U21947 (N_21947,N_20714,N_20764);
or U21948 (N_21948,N_20486,N_20707);
xor U21949 (N_21949,N_20182,N_20933);
or U21950 (N_21950,N_20115,N_20145);
nand U21951 (N_21951,N_20090,N_20757);
nor U21952 (N_21952,N_20214,N_20889);
or U21953 (N_21953,N_20941,N_20386);
nor U21954 (N_21954,N_20439,N_20751);
and U21955 (N_21955,N_20416,N_20349);
or U21956 (N_21956,N_20545,N_20212);
nand U21957 (N_21957,N_20183,N_20638);
or U21958 (N_21958,N_20520,N_20354);
nand U21959 (N_21959,N_20181,N_20127);
and U21960 (N_21960,N_20966,N_20206);
nor U21961 (N_21961,N_20472,N_20964);
nand U21962 (N_21962,N_20236,N_20744);
or U21963 (N_21963,N_20237,N_20303);
and U21964 (N_21964,N_20589,N_20725);
xnor U21965 (N_21965,N_20790,N_20425);
nor U21966 (N_21966,N_20039,N_20828);
nor U21967 (N_21967,N_20390,N_20700);
and U21968 (N_21968,N_20058,N_20465);
nand U21969 (N_21969,N_20597,N_20916);
nor U21970 (N_21970,N_20069,N_20127);
or U21971 (N_21971,N_20431,N_20881);
nand U21972 (N_21972,N_20092,N_20659);
xnor U21973 (N_21973,N_20572,N_20505);
and U21974 (N_21974,N_20512,N_20255);
and U21975 (N_21975,N_20960,N_20939);
or U21976 (N_21976,N_20843,N_20196);
nand U21977 (N_21977,N_20728,N_20463);
or U21978 (N_21978,N_20618,N_20185);
nand U21979 (N_21979,N_20200,N_20840);
nand U21980 (N_21980,N_20921,N_20740);
xor U21981 (N_21981,N_20008,N_20580);
xnor U21982 (N_21982,N_20268,N_20178);
and U21983 (N_21983,N_20687,N_20453);
nand U21984 (N_21984,N_20074,N_20373);
nor U21985 (N_21985,N_20860,N_20444);
nand U21986 (N_21986,N_20929,N_20682);
xnor U21987 (N_21987,N_20266,N_20678);
nand U21988 (N_21988,N_20348,N_20399);
xor U21989 (N_21989,N_20943,N_20448);
or U21990 (N_21990,N_20479,N_20815);
nor U21991 (N_21991,N_20313,N_20476);
nand U21992 (N_21992,N_20215,N_20621);
or U21993 (N_21993,N_20803,N_20787);
xnor U21994 (N_21994,N_20239,N_20769);
nand U21995 (N_21995,N_20805,N_20207);
nand U21996 (N_21996,N_20503,N_20687);
nand U21997 (N_21997,N_20856,N_20178);
nand U21998 (N_21998,N_20509,N_20744);
or U21999 (N_21999,N_20322,N_20908);
nand U22000 (N_22000,N_21718,N_21515);
xnor U22001 (N_22001,N_21141,N_21335);
nand U22002 (N_22002,N_21761,N_21380);
xnor U22003 (N_22003,N_21442,N_21531);
and U22004 (N_22004,N_21259,N_21486);
or U22005 (N_22005,N_21524,N_21615);
or U22006 (N_22006,N_21426,N_21365);
and U22007 (N_22007,N_21988,N_21474);
nand U22008 (N_22008,N_21996,N_21928);
and U22009 (N_22009,N_21063,N_21134);
and U22010 (N_22010,N_21030,N_21495);
and U22011 (N_22011,N_21060,N_21088);
nand U22012 (N_22012,N_21298,N_21168);
nor U22013 (N_22013,N_21385,N_21744);
xnor U22014 (N_22014,N_21084,N_21845);
and U22015 (N_22015,N_21910,N_21956);
nand U22016 (N_22016,N_21086,N_21350);
and U22017 (N_22017,N_21596,N_21138);
nand U22018 (N_22018,N_21483,N_21042);
nand U22019 (N_22019,N_21386,N_21758);
xnor U22020 (N_22020,N_21831,N_21711);
nand U22021 (N_22021,N_21942,N_21287);
or U22022 (N_22022,N_21919,N_21931);
nand U22023 (N_22023,N_21684,N_21820);
nor U22024 (N_22024,N_21713,N_21962);
nor U22025 (N_22025,N_21303,N_21308);
or U22026 (N_22026,N_21485,N_21267);
nand U22027 (N_22027,N_21216,N_21767);
nor U22028 (N_22028,N_21853,N_21858);
or U22029 (N_22029,N_21302,N_21887);
xor U22030 (N_22030,N_21059,N_21791);
nand U22031 (N_22031,N_21582,N_21462);
or U22032 (N_22032,N_21629,N_21904);
or U22033 (N_22033,N_21435,N_21850);
xor U22034 (N_22034,N_21561,N_21207);
or U22035 (N_22035,N_21292,N_21448);
or U22036 (N_22036,N_21158,N_21519);
nor U22037 (N_22037,N_21508,N_21450);
and U22038 (N_22038,N_21983,N_21768);
or U22039 (N_22039,N_21021,N_21129);
nand U22040 (N_22040,N_21798,N_21098);
nor U22041 (N_22041,N_21563,N_21861);
nor U22042 (N_22042,N_21407,N_21116);
nor U22043 (N_22043,N_21955,N_21149);
and U22044 (N_22044,N_21081,N_21449);
or U22045 (N_22045,N_21429,N_21248);
nor U22046 (N_22046,N_21225,N_21566);
xor U22047 (N_22047,N_21576,N_21991);
or U22048 (N_22048,N_21705,N_21899);
xor U22049 (N_22049,N_21943,N_21927);
or U22050 (N_22050,N_21505,N_21218);
xnor U22051 (N_22051,N_21989,N_21388);
or U22052 (N_22052,N_21265,N_21987);
nand U22053 (N_22053,N_21630,N_21359);
nor U22054 (N_22054,N_21215,N_21314);
or U22055 (N_22055,N_21725,N_21854);
xnor U22056 (N_22056,N_21840,N_21774);
nor U22057 (N_22057,N_21530,N_21310);
or U22058 (N_22058,N_21214,N_21393);
and U22059 (N_22059,N_21280,N_21620);
nand U22060 (N_22060,N_21644,N_21010);
xor U22061 (N_22061,N_21476,N_21006);
xnor U22062 (N_22062,N_21747,N_21307);
nand U22063 (N_22063,N_21982,N_21814);
and U22064 (N_22064,N_21281,N_21704);
and U22065 (N_22065,N_21464,N_21222);
nand U22066 (N_22066,N_21169,N_21183);
nor U22067 (N_22067,N_21773,N_21522);
nor U22068 (N_22068,N_21258,N_21616);
nor U22069 (N_22069,N_21201,N_21889);
or U22070 (N_22070,N_21130,N_21080);
and U22071 (N_22071,N_21839,N_21806);
nand U22072 (N_22072,N_21184,N_21502);
and U22073 (N_22073,N_21602,N_21613);
nand U22074 (N_22074,N_21859,N_21998);
nor U22075 (N_22075,N_21673,N_21078);
xor U22076 (N_22076,N_21750,N_21586);
nor U22077 (N_22077,N_21631,N_21945);
nor U22078 (N_22078,N_21004,N_21875);
or U22079 (N_22079,N_21735,N_21396);
xnor U22080 (N_22080,N_21319,N_21473);
nand U22081 (N_22081,N_21066,N_21901);
and U22082 (N_22082,N_21651,N_21491);
and U22083 (N_22083,N_21572,N_21173);
nor U22084 (N_22084,N_21667,N_21848);
nor U22085 (N_22085,N_21097,N_21900);
xor U22086 (N_22086,N_21120,N_21946);
nand U22087 (N_22087,N_21057,N_21961);
xnor U22088 (N_22088,N_21855,N_21997);
or U22089 (N_22089,N_21344,N_21096);
nor U22090 (N_22090,N_21489,N_21568);
nor U22091 (N_22091,N_21699,N_21133);
nand U22092 (N_22092,N_21271,N_21441);
nand U22093 (N_22093,N_21706,N_21804);
and U22094 (N_22094,N_21465,N_21234);
nor U22095 (N_22095,N_21870,N_21577);
xor U22096 (N_22096,N_21322,N_21019);
or U22097 (N_22097,N_21581,N_21769);
and U22098 (N_22098,N_21005,N_21023);
or U22099 (N_22099,N_21682,N_21075);
nor U22100 (N_22100,N_21438,N_21797);
nand U22101 (N_22101,N_21406,N_21578);
nor U22102 (N_22102,N_21600,N_21695);
nor U22103 (N_22103,N_21389,N_21362);
or U22104 (N_22104,N_21847,N_21580);
nor U22105 (N_22105,N_21147,N_21364);
nor U22106 (N_22106,N_21224,N_21748);
nand U22107 (N_22107,N_21492,N_21082);
xnor U22108 (N_22108,N_21049,N_21941);
nand U22109 (N_22109,N_21148,N_21377);
and U22110 (N_22110,N_21624,N_21361);
and U22111 (N_22111,N_21356,N_21893);
and U22112 (N_22112,N_21410,N_21331);
xnor U22113 (N_22113,N_21151,N_21549);
and U22114 (N_22114,N_21205,N_21683);
nor U22115 (N_22115,N_21822,N_21570);
nand U22116 (N_22116,N_21497,N_21881);
or U22117 (N_22117,N_21805,N_21771);
and U22118 (N_22118,N_21488,N_21069);
nor U22119 (N_22119,N_21228,N_21587);
or U22120 (N_22120,N_21918,N_21415);
xnor U22121 (N_22121,N_21609,N_21527);
nor U22122 (N_22122,N_21295,N_21584);
nor U22123 (N_22123,N_21702,N_21990);
nand U22124 (N_22124,N_21249,N_21874);
nor U22125 (N_22125,N_21413,N_21643);
nor U22126 (N_22126,N_21073,N_21440);
or U22127 (N_22127,N_21679,N_21812);
nor U22128 (N_22128,N_21455,N_21716);
nor U22129 (N_22129,N_21313,N_21504);
xor U22130 (N_22130,N_21425,N_21551);
and U22131 (N_22131,N_21018,N_21334);
nand U22132 (N_22132,N_21035,N_21293);
nand U22133 (N_22133,N_21211,N_21039);
nand U22134 (N_22134,N_21968,N_21015);
or U22135 (N_22135,N_21276,N_21866);
nand U22136 (N_22136,N_21724,N_21903);
nand U22137 (N_22137,N_21008,N_21227);
xnor U22138 (N_22138,N_21418,N_21503);
and U22139 (N_22139,N_21783,N_21112);
or U22140 (N_22140,N_21601,N_21826);
and U22141 (N_22141,N_21051,N_21756);
nor U22142 (N_22142,N_21381,N_21432);
xnor U22143 (N_22143,N_21034,N_21040);
or U22144 (N_22144,N_21178,N_21970);
and U22145 (N_22145,N_21548,N_21604);
nor U22146 (N_22146,N_21871,N_21852);
xnor U22147 (N_22147,N_21730,N_21779);
and U22148 (N_22148,N_21647,N_21443);
or U22149 (N_22149,N_21339,N_21099);
and U22150 (N_22150,N_21213,N_21496);
and U22151 (N_22151,N_21430,N_21083);
and U22152 (N_22152,N_21275,N_21501);
nor U22153 (N_22153,N_21772,N_21226);
nor U22154 (N_22154,N_21204,N_21564);
and U22155 (N_22155,N_21456,N_21740);
nand U22156 (N_22156,N_21318,N_21846);
and U22157 (N_22157,N_21938,N_21793);
nand U22158 (N_22158,N_21424,N_21958);
or U22159 (N_22159,N_21786,N_21646);
nand U22160 (N_22160,N_21825,N_21177);
nor U22161 (N_22161,N_21967,N_21268);
nor U22162 (N_22162,N_21614,N_21709);
nand U22163 (N_22163,N_21995,N_21939);
and U22164 (N_22164,N_21033,N_21074);
nor U22165 (N_22165,N_21865,N_21746);
or U22166 (N_22166,N_21710,N_21403);
xnor U22167 (N_22167,N_21002,N_21460);
or U22168 (N_22168,N_21165,N_21011);
xor U22169 (N_22169,N_21001,N_21144);
nor U22170 (N_22170,N_21431,N_21209);
nor U22171 (N_22171,N_21934,N_21680);
nand U22172 (N_22172,N_21762,N_21553);
xnor U22173 (N_22173,N_21729,N_21072);
nor U22174 (N_22174,N_21022,N_21003);
nand U22175 (N_22175,N_21171,N_21575);
and U22176 (N_22176,N_21583,N_21017);
or U22177 (N_22177,N_21664,N_21283);
or U22178 (N_22178,N_21367,N_21662);
nand U22179 (N_22179,N_21212,N_21890);
xor U22180 (N_22180,N_21045,N_21411);
or U22181 (N_22181,N_21546,N_21597);
xnor U22182 (N_22182,N_21787,N_21252);
nand U22183 (N_22183,N_21885,N_21542);
nor U22184 (N_22184,N_21844,N_21694);
nor U22185 (N_22185,N_21020,N_21944);
and U22186 (N_22186,N_21196,N_21693);
or U22187 (N_22187,N_21880,N_21284);
or U22188 (N_22188,N_21816,N_21079);
xnor U22189 (N_22189,N_21969,N_21437);
xnor U22190 (N_22190,N_21463,N_21327);
nor U22191 (N_22191,N_21077,N_21291);
and U22192 (N_22192,N_21154,N_21778);
or U22193 (N_22193,N_21398,N_21980);
and U22194 (N_22194,N_21330,N_21898);
and U22195 (N_22195,N_21338,N_21780);
nand U22196 (N_22196,N_21557,N_21626);
or U22197 (N_22197,N_21357,N_21421);
and U22198 (N_22198,N_21832,N_21311);
or U22199 (N_22199,N_21813,N_21482);
xor U22200 (N_22200,N_21690,N_21558);
nand U22201 (N_22201,N_21156,N_21883);
nor U22202 (N_22202,N_21608,N_21223);
and U22203 (N_22203,N_21119,N_21766);
or U22204 (N_22204,N_21959,N_21652);
xor U22205 (N_22205,N_21366,N_21041);
xnor U22206 (N_22206,N_21288,N_21061);
or U22207 (N_22207,N_21470,N_21529);
and U22208 (N_22208,N_21765,N_21187);
nand U22209 (N_22209,N_21164,N_21741);
xnor U22210 (N_22210,N_21979,N_21838);
nand U22211 (N_22211,N_21315,N_21737);
and U22212 (N_22212,N_21777,N_21500);
xnor U22213 (N_22213,N_21126,N_21255);
and U22214 (N_22214,N_21416,N_21137);
or U22215 (N_22215,N_21090,N_21146);
and U22216 (N_22216,N_21957,N_21534);
nand U22217 (N_22217,N_21487,N_21627);
xnor U22218 (N_22218,N_21043,N_21317);
nand U22219 (N_22219,N_21867,N_21118);
xnor U22220 (N_22220,N_21573,N_21949);
and U22221 (N_22221,N_21922,N_21068);
nor U22222 (N_22222,N_21236,N_21301);
nand U22223 (N_22223,N_21562,N_21947);
or U22224 (N_22224,N_21404,N_21790);
or U22225 (N_22225,N_21469,N_21677);
nor U22226 (N_22226,N_21610,N_21185);
and U22227 (N_22227,N_21902,N_21985);
or U22228 (N_22228,N_21738,N_21794);
and U22229 (N_22229,N_21712,N_21749);
nand U22230 (N_22230,N_21210,N_21325);
and U22231 (N_22231,N_21321,N_21160);
nor U22232 (N_22232,N_21000,N_21190);
nand U22233 (N_22233,N_21672,N_21188);
or U22234 (N_22234,N_21194,N_21521);
nand U22235 (N_22235,N_21166,N_21815);
nand U22236 (N_22236,N_21451,N_21197);
or U22237 (N_22237,N_21402,N_21309);
nor U22238 (N_22238,N_21954,N_21191);
xor U22239 (N_22239,N_21262,N_21810);
nand U22240 (N_22240,N_21447,N_21481);
nand U22241 (N_22241,N_21828,N_21506);
and U22242 (N_22242,N_21665,N_21466);
nand U22243 (N_22243,N_21897,N_21100);
or U22244 (N_22244,N_21294,N_21930);
nor U22245 (N_22245,N_21528,N_21490);
nand U22246 (N_22246,N_21419,N_21670);
and U22247 (N_22247,N_21297,N_21924);
xor U22248 (N_22248,N_21976,N_21175);
nand U22249 (N_22249,N_21127,N_21688);
nand U22250 (N_22250,N_21278,N_21660);
xor U22251 (N_22251,N_21697,N_21550);
nor U22252 (N_22252,N_21089,N_21478);
or U22253 (N_22253,N_21849,N_21370);
xnor U22254 (N_22254,N_21556,N_21895);
nor U22255 (N_22255,N_21532,N_21101);
nand U22256 (N_22256,N_21544,N_21993);
and U22257 (N_22257,N_21621,N_21172);
or U22258 (N_22258,N_21541,N_21540);
nand U22259 (N_22259,N_21841,N_21727);
or U22260 (N_22260,N_21369,N_21567);
or U22261 (N_22261,N_21868,N_21108);
xnor U22262 (N_22262,N_21428,N_21842);
xnor U22263 (N_22263,N_21819,N_21594);
and U22264 (N_22264,N_21378,N_21263);
nand U22265 (N_22265,N_21676,N_21799);
xor U22266 (N_22266,N_21111,N_21731);
and U22267 (N_22267,N_21843,N_21827);
xnor U22268 (N_22268,N_21739,N_21390);
xnor U22269 (N_22269,N_21498,N_21675);
nand U22270 (N_22270,N_21065,N_21289);
nand U22271 (N_22271,N_21760,N_21299);
or U22272 (N_22272,N_21170,N_21221);
or U22273 (N_22273,N_21669,N_21208);
or U22274 (N_22274,N_21121,N_21346);
nand U22275 (N_22275,N_21994,N_21836);
nand U22276 (N_22276,N_21494,N_21102);
xor U22277 (N_22277,N_21666,N_21510);
or U22278 (N_22278,N_21547,N_21445);
nor U22279 (N_22279,N_21543,N_21878);
or U22280 (N_22280,N_21016,N_21131);
nor U22281 (N_22281,N_21714,N_21717);
nand U22282 (N_22282,N_21349,N_21351);
nand U22283 (N_22283,N_21745,N_21231);
or U22284 (N_22284,N_21135,N_21094);
nor U22285 (N_22285,N_21353,N_21408);
nor U22286 (N_22286,N_21638,N_21220);
nand U22287 (N_22287,N_21818,N_21243);
nand U22288 (N_22288,N_21142,N_21400);
xor U22289 (N_22289,N_21181,N_21873);
nand U22290 (N_22290,N_21981,N_21296);
or U22291 (N_22291,N_21571,N_21340);
xor U22292 (N_22292,N_21992,N_21862);
nor U22293 (N_22293,N_21452,N_21833);
nor U22294 (N_22294,N_21085,N_21513);
xor U22295 (N_22295,N_21246,N_21368);
and U22296 (N_22296,N_21189,N_21908);
or U22297 (N_22297,N_21517,N_21117);
nand U22298 (N_22298,N_21233,N_21764);
nor U22299 (N_22299,N_21835,N_21305);
and U22300 (N_22300,N_21807,N_21701);
nor U22301 (N_22301,N_21726,N_21374);
and U22302 (N_22302,N_21105,N_21417);
xnor U22303 (N_22303,N_21555,N_21590);
or U22304 (N_22304,N_21113,N_21789);
or U22305 (N_22305,N_21434,N_21014);
or U22306 (N_22306,N_21054,N_21024);
or U22307 (N_22307,N_21755,N_21678);
nand U22308 (N_22308,N_21395,N_21484);
or U22309 (N_22309,N_21480,N_21387);
nand U22310 (N_22310,N_21625,N_21559);
nand U22311 (N_22311,N_21607,N_21264);
nor U22312 (N_22312,N_21312,N_21723);
and U22313 (N_22313,N_21087,N_21458);
or U22314 (N_22314,N_21752,N_21921);
and U22315 (N_22315,N_21459,N_21479);
or U22316 (N_22316,N_21892,N_21384);
or U22317 (N_22317,N_21115,N_21538);
xnor U22318 (N_22318,N_21800,N_21106);
and U22319 (N_22319,N_21341,N_21273);
xnor U22320 (N_22320,N_21592,N_21457);
xor U22321 (N_22321,N_21689,N_21446);
nand U22322 (N_22322,N_21007,N_21122);
nor U22323 (N_22323,N_21427,N_21070);
and U22324 (N_22324,N_21091,N_21863);
or U22325 (N_22325,N_21525,N_21326);
nand U22326 (N_22326,N_21235,N_21076);
xor U22327 (N_22327,N_21145,N_21055);
and U22328 (N_22328,N_21948,N_21320);
and U22329 (N_22329,N_21230,N_21238);
nand U22330 (N_22330,N_21661,N_21645);
and U22331 (N_22331,N_21972,N_21894);
nor U22332 (N_22332,N_21656,N_21179);
nand U22333 (N_22333,N_21788,N_21648);
nor U22334 (N_22334,N_21046,N_21044);
nor U22335 (N_22335,N_21668,N_21692);
nor U22336 (N_22336,N_21195,N_21728);
or U22337 (N_22337,N_21250,N_21244);
nand U22338 (N_22338,N_21781,N_21036);
nor U22339 (N_22339,N_21067,N_21256);
nor U22340 (N_22340,N_21879,N_21260);
xor U22341 (N_22341,N_21143,N_21823);
nand U22342 (N_22342,N_21593,N_21423);
xnor U22343 (N_22343,N_21512,N_21038);
xnor U22344 (N_22344,N_21891,N_21926);
and U22345 (N_22345,N_21591,N_21655);
nor U22346 (N_22346,N_21757,N_21304);
or U22347 (N_22347,N_21439,N_21639);
or U22348 (N_22348,N_21654,N_21588);
or U22349 (N_22349,N_21025,N_21792);
or U22350 (N_22350,N_21518,N_21200);
xnor U22351 (N_22351,N_21554,N_21342);
xnor U22352 (N_22352,N_21623,N_21619);
or U22353 (N_22353,N_21092,N_21569);
xnor U22354 (N_22354,N_21920,N_21093);
and U22355 (N_22355,N_21152,N_21720);
or U22356 (N_22356,N_21733,N_21708);
xnor U22357 (N_22357,N_21539,N_21056);
nor U22358 (N_22358,N_21401,N_21526);
xnor U22359 (N_22359,N_21270,N_21493);
and U22360 (N_22360,N_21633,N_21964);
nand U22361 (N_22361,N_21912,N_21963);
or U22362 (N_22362,N_21770,N_21649);
nor U22363 (N_22363,N_21808,N_21742);
nand U22364 (N_22364,N_21420,N_21743);
and U22365 (N_22365,N_21950,N_21192);
nor U22366 (N_22366,N_21472,N_21240);
nor U22367 (N_22367,N_21477,N_21139);
nand U22368 (N_22368,N_21932,N_21132);
and U22369 (N_22369,N_21953,N_21906);
or U22370 (N_22370,N_21632,N_21336);
xor U22371 (N_22371,N_21155,N_21971);
or U22372 (N_22372,N_21343,N_21009);
nor U22373 (N_22373,N_21376,N_21329);
nand U22374 (N_22374,N_21817,N_21261);
xor U22375 (N_22375,N_21373,N_21659);
nand U22376 (N_22376,N_21785,N_21560);
and U22377 (N_22377,N_21124,N_21383);
xnor U22378 (N_22378,N_21685,N_21161);
xnor U22379 (N_22379,N_21691,N_21203);
or U22380 (N_22380,N_21872,N_21719);
or U22381 (N_22381,N_21186,N_21877);
or U22382 (N_22382,N_21123,N_21707);
nor U22383 (N_22383,N_21290,N_21860);
or U22384 (N_22384,N_21657,N_21925);
or U22385 (N_22385,N_21153,N_21611);
xnor U22386 (N_22386,N_21888,N_21612);
xor U22387 (N_22387,N_21409,N_21811);
or U22388 (N_22388,N_21219,N_21461);
and U22389 (N_22389,N_21382,N_21174);
nand U22390 (N_22390,N_21606,N_21864);
and U22391 (N_22391,N_21360,N_21937);
and U22392 (N_22392,N_21681,N_21300);
nor U22393 (N_22393,N_21975,N_21199);
and U22394 (N_22394,N_21869,N_21973);
xnor U22395 (N_22395,N_21809,N_21715);
nor U22396 (N_22396,N_21444,N_21722);
nor U22397 (N_22397,N_21795,N_21574);
nand U22398 (N_22398,N_21436,N_21274);
xor U22399 (N_22399,N_21414,N_21372);
nand U22400 (N_22400,N_21150,N_21514);
and U22401 (N_22401,N_21251,N_21266);
or U22402 (N_22402,N_21277,N_21279);
and U22403 (N_22403,N_21348,N_21110);
nand U22404 (N_22404,N_21978,N_21617);
nor U22405 (N_22405,N_21984,N_21935);
and U22406 (N_22406,N_21062,N_21037);
xor U22407 (N_22407,N_21700,N_21876);
and U22408 (N_22408,N_21965,N_21915);
or U22409 (N_22409,N_21333,N_21658);
and U22410 (N_22410,N_21782,N_21650);
xnor U22411 (N_22411,N_21851,N_21585);
or U22412 (N_22412,N_21242,N_21687);
xnor U22413 (N_22413,N_21337,N_21751);
nor U22414 (N_22414,N_21703,N_21167);
nand U22415 (N_22415,N_21802,N_21986);
and U22416 (N_22416,N_21837,N_21285);
nand U22417 (N_22417,N_21058,N_21397);
nor U22418 (N_22418,N_21775,N_21732);
xor U22419 (N_22419,N_21829,N_21052);
xor U22420 (N_22420,N_21974,N_21050);
nor U22421 (N_22421,N_21999,N_21951);
xnor U22422 (N_22422,N_21405,N_21162);
or U22423 (N_22423,N_21537,N_21157);
xor U22424 (N_22424,N_21128,N_21371);
or U22425 (N_22425,N_21332,N_21640);
nand U22426 (N_22426,N_21229,N_21394);
nand U22427 (N_22427,N_21392,N_21721);
nand U22428 (N_22428,N_21286,N_21929);
xor U22429 (N_22429,N_21114,N_21509);
xor U22430 (N_22430,N_21104,N_21355);
and U22431 (N_22431,N_21412,N_21422);
and U22432 (N_22432,N_21966,N_21907);
xnor U22433 (N_22433,N_21671,N_21159);
and U22434 (N_22434,N_21622,N_21511);
nor U22435 (N_22435,N_21923,N_21535);
nor U22436 (N_22436,N_21977,N_21598);
xor U22437 (N_22437,N_21952,N_21032);
xnor U22438 (N_22438,N_21579,N_21834);
xnor U22439 (N_22439,N_21821,N_21830);
xnor U22440 (N_22440,N_21026,N_21140);
and U22441 (N_22441,N_21565,N_21523);
nand U22442 (N_22442,N_21109,N_21107);
nand U22443 (N_22443,N_21824,N_21595);
nand U22444 (N_22444,N_21734,N_21674);
nand U22445 (N_22445,N_21763,N_21347);
nand U22446 (N_22446,N_21467,N_21391);
or U22447 (N_22447,N_21642,N_21217);
nor U22448 (N_22448,N_21801,N_21375);
nand U22449 (N_22449,N_21198,N_21323);
nand U22450 (N_22450,N_21796,N_21636);
nand U22451 (N_22451,N_21202,N_21247);
or U22452 (N_22452,N_21499,N_21916);
or U22453 (N_22453,N_21545,N_21125);
xor U22454 (N_22454,N_21363,N_21886);
and U22455 (N_22455,N_21206,N_21237);
nor U22456 (N_22456,N_21882,N_21905);
and U22457 (N_22457,N_21776,N_21533);
nand U22458 (N_22458,N_21618,N_21064);
and U22459 (N_22459,N_21603,N_21232);
nor U22460 (N_22460,N_21507,N_21029);
and U22461 (N_22461,N_21031,N_21940);
or U22462 (N_22462,N_21163,N_21917);
xnor U22463 (N_22463,N_21027,N_21759);
or U22464 (N_22464,N_21784,N_21552);
nor U22465 (N_22465,N_21245,N_21433);
nor U22466 (N_22466,N_21663,N_21896);
xor U22467 (N_22467,N_21071,N_21637);
and U22468 (N_22468,N_21328,N_21698);
nor U22469 (N_22469,N_21911,N_21933);
xor U22470 (N_22470,N_21182,N_21269);
nand U22471 (N_22471,N_21012,N_21653);
nand U22472 (N_22472,N_21628,N_21345);
nand U22473 (N_22473,N_21354,N_21536);
and U22474 (N_22474,N_21358,N_21399);
nor U22475 (N_22475,N_21475,N_21180);
nand U22476 (N_22476,N_21282,N_21754);
and U22477 (N_22477,N_21176,N_21641);
xor U22478 (N_22478,N_21913,N_21599);
or U22479 (N_22479,N_21316,N_21635);
xor U22480 (N_22480,N_21803,N_21960);
nand U22481 (N_22481,N_21095,N_21028);
nand U22482 (N_22482,N_21324,N_21468);
nor U22483 (N_22483,N_21241,N_21453);
nand U22484 (N_22484,N_21053,N_21634);
or U22485 (N_22485,N_21272,N_21753);
or U22486 (N_22486,N_21589,N_21239);
nor U22487 (N_22487,N_21047,N_21352);
and U22488 (N_22488,N_21516,N_21013);
and U22489 (N_22489,N_21696,N_21306);
or U22490 (N_22490,N_21257,N_21253);
nand U22491 (N_22491,N_21254,N_21856);
and U22492 (N_22492,N_21471,N_21379);
xnor U22493 (N_22493,N_21936,N_21520);
nor U22494 (N_22494,N_21857,N_21686);
and U22495 (N_22495,N_21914,N_21454);
and U22496 (N_22496,N_21193,N_21884);
or U22497 (N_22497,N_21048,N_21736);
and U22498 (N_22498,N_21136,N_21605);
or U22499 (N_22499,N_21909,N_21103);
nand U22500 (N_22500,N_21576,N_21756);
nor U22501 (N_22501,N_21729,N_21519);
nor U22502 (N_22502,N_21796,N_21813);
or U22503 (N_22503,N_21353,N_21470);
xor U22504 (N_22504,N_21912,N_21326);
nand U22505 (N_22505,N_21543,N_21903);
and U22506 (N_22506,N_21333,N_21029);
nand U22507 (N_22507,N_21621,N_21362);
nand U22508 (N_22508,N_21008,N_21007);
and U22509 (N_22509,N_21407,N_21396);
nor U22510 (N_22510,N_21098,N_21075);
nor U22511 (N_22511,N_21654,N_21979);
or U22512 (N_22512,N_21421,N_21022);
xnor U22513 (N_22513,N_21823,N_21285);
and U22514 (N_22514,N_21882,N_21187);
xnor U22515 (N_22515,N_21803,N_21273);
nor U22516 (N_22516,N_21035,N_21216);
or U22517 (N_22517,N_21445,N_21347);
xor U22518 (N_22518,N_21026,N_21782);
or U22519 (N_22519,N_21802,N_21638);
or U22520 (N_22520,N_21692,N_21784);
nor U22521 (N_22521,N_21461,N_21393);
xnor U22522 (N_22522,N_21873,N_21524);
nand U22523 (N_22523,N_21348,N_21182);
nand U22524 (N_22524,N_21502,N_21144);
xor U22525 (N_22525,N_21122,N_21478);
and U22526 (N_22526,N_21378,N_21108);
xnor U22527 (N_22527,N_21521,N_21921);
nor U22528 (N_22528,N_21297,N_21186);
and U22529 (N_22529,N_21704,N_21817);
or U22530 (N_22530,N_21760,N_21469);
and U22531 (N_22531,N_21807,N_21430);
nand U22532 (N_22532,N_21985,N_21131);
nor U22533 (N_22533,N_21915,N_21676);
and U22534 (N_22534,N_21839,N_21548);
xor U22535 (N_22535,N_21569,N_21585);
xor U22536 (N_22536,N_21346,N_21090);
nor U22537 (N_22537,N_21992,N_21407);
xor U22538 (N_22538,N_21406,N_21822);
nor U22539 (N_22539,N_21213,N_21661);
nor U22540 (N_22540,N_21007,N_21325);
nand U22541 (N_22541,N_21526,N_21386);
and U22542 (N_22542,N_21462,N_21595);
xnor U22543 (N_22543,N_21655,N_21516);
or U22544 (N_22544,N_21314,N_21770);
nor U22545 (N_22545,N_21202,N_21677);
or U22546 (N_22546,N_21059,N_21631);
xnor U22547 (N_22547,N_21270,N_21479);
xnor U22548 (N_22548,N_21737,N_21453);
nor U22549 (N_22549,N_21801,N_21178);
or U22550 (N_22550,N_21208,N_21673);
nor U22551 (N_22551,N_21299,N_21375);
nand U22552 (N_22552,N_21108,N_21331);
nand U22553 (N_22553,N_21259,N_21834);
nor U22554 (N_22554,N_21508,N_21067);
xor U22555 (N_22555,N_21262,N_21483);
nor U22556 (N_22556,N_21806,N_21038);
nor U22557 (N_22557,N_21137,N_21544);
and U22558 (N_22558,N_21357,N_21114);
or U22559 (N_22559,N_21346,N_21430);
nand U22560 (N_22560,N_21829,N_21445);
or U22561 (N_22561,N_21762,N_21494);
or U22562 (N_22562,N_21949,N_21562);
xnor U22563 (N_22563,N_21052,N_21733);
nor U22564 (N_22564,N_21146,N_21522);
nor U22565 (N_22565,N_21673,N_21658);
nor U22566 (N_22566,N_21282,N_21527);
or U22567 (N_22567,N_21448,N_21752);
or U22568 (N_22568,N_21828,N_21145);
nor U22569 (N_22569,N_21559,N_21866);
or U22570 (N_22570,N_21648,N_21852);
or U22571 (N_22571,N_21941,N_21285);
or U22572 (N_22572,N_21233,N_21254);
nand U22573 (N_22573,N_21358,N_21325);
and U22574 (N_22574,N_21561,N_21141);
nand U22575 (N_22575,N_21403,N_21511);
nand U22576 (N_22576,N_21718,N_21417);
or U22577 (N_22577,N_21438,N_21115);
nand U22578 (N_22578,N_21592,N_21576);
nor U22579 (N_22579,N_21264,N_21998);
and U22580 (N_22580,N_21831,N_21453);
nor U22581 (N_22581,N_21554,N_21568);
xnor U22582 (N_22582,N_21559,N_21969);
or U22583 (N_22583,N_21600,N_21195);
nor U22584 (N_22584,N_21887,N_21280);
nor U22585 (N_22585,N_21611,N_21647);
xnor U22586 (N_22586,N_21601,N_21117);
or U22587 (N_22587,N_21847,N_21379);
xnor U22588 (N_22588,N_21558,N_21847);
or U22589 (N_22589,N_21545,N_21578);
xnor U22590 (N_22590,N_21045,N_21464);
and U22591 (N_22591,N_21976,N_21002);
nand U22592 (N_22592,N_21849,N_21695);
xnor U22593 (N_22593,N_21037,N_21664);
nand U22594 (N_22594,N_21713,N_21705);
and U22595 (N_22595,N_21147,N_21896);
or U22596 (N_22596,N_21051,N_21052);
nor U22597 (N_22597,N_21880,N_21167);
xnor U22598 (N_22598,N_21309,N_21537);
and U22599 (N_22599,N_21304,N_21516);
xor U22600 (N_22600,N_21138,N_21813);
xnor U22601 (N_22601,N_21882,N_21684);
xor U22602 (N_22602,N_21306,N_21081);
nor U22603 (N_22603,N_21339,N_21596);
xor U22604 (N_22604,N_21703,N_21261);
and U22605 (N_22605,N_21829,N_21567);
xnor U22606 (N_22606,N_21735,N_21650);
and U22607 (N_22607,N_21209,N_21624);
and U22608 (N_22608,N_21157,N_21735);
and U22609 (N_22609,N_21323,N_21713);
and U22610 (N_22610,N_21694,N_21325);
nor U22611 (N_22611,N_21107,N_21219);
and U22612 (N_22612,N_21104,N_21631);
nand U22613 (N_22613,N_21086,N_21261);
nor U22614 (N_22614,N_21108,N_21237);
nor U22615 (N_22615,N_21147,N_21263);
and U22616 (N_22616,N_21249,N_21756);
or U22617 (N_22617,N_21365,N_21301);
or U22618 (N_22618,N_21966,N_21067);
nor U22619 (N_22619,N_21459,N_21004);
nand U22620 (N_22620,N_21470,N_21550);
nand U22621 (N_22621,N_21125,N_21496);
nand U22622 (N_22622,N_21374,N_21133);
or U22623 (N_22623,N_21930,N_21602);
or U22624 (N_22624,N_21835,N_21575);
or U22625 (N_22625,N_21700,N_21585);
or U22626 (N_22626,N_21031,N_21334);
nor U22627 (N_22627,N_21414,N_21829);
and U22628 (N_22628,N_21660,N_21860);
nor U22629 (N_22629,N_21954,N_21037);
nand U22630 (N_22630,N_21686,N_21932);
nand U22631 (N_22631,N_21669,N_21992);
and U22632 (N_22632,N_21133,N_21211);
xnor U22633 (N_22633,N_21933,N_21312);
nand U22634 (N_22634,N_21631,N_21967);
or U22635 (N_22635,N_21998,N_21719);
and U22636 (N_22636,N_21353,N_21305);
nand U22637 (N_22637,N_21969,N_21986);
xnor U22638 (N_22638,N_21403,N_21753);
or U22639 (N_22639,N_21361,N_21682);
and U22640 (N_22640,N_21957,N_21187);
and U22641 (N_22641,N_21364,N_21047);
and U22642 (N_22642,N_21930,N_21151);
xor U22643 (N_22643,N_21244,N_21906);
or U22644 (N_22644,N_21692,N_21843);
and U22645 (N_22645,N_21122,N_21305);
nand U22646 (N_22646,N_21686,N_21579);
or U22647 (N_22647,N_21964,N_21463);
and U22648 (N_22648,N_21270,N_21097);
nand U22649 (N_22649,N_21984,N_21581);
and U22650 (N_22650,N_21226,N_21858);
and U22651 (N_22651,N_21653,N_21059);
xnor U22652 (N_22652,N_21385,N_21969);
xor U22653 (N_22653,N_21277,N_21242);
nand U22654 (N_22654,N_21493,N_21318);
nor U22655 (N_22655,N_21584,N_21858);
or U22656 (N_22656,N_21323,N_21843);
xor U22657 (N_22657,N_21582,N_21333);
nor U22658 (N_22658,N_21218,N_21193);
nor U22659 (N_22659,N_21628,N_21072);
nand U22660 (N_22660,N_21229,N_21952);
or U22661 (N_22661,N_21326,N_21826);
xnor U22662 (N_22662,N_21669,N_21295);
or U22663 (N_22663,N_21979,N_21803);
nand U22664 (N_22664,N_21485,N_21356);
nor U22665 (N_22665,N_21888,N_21851);
and U22666 (N_22666,N_21574,N_21029);
nor U22667 (N_22667,N_21915,N_21754);
and U22668 (N_22668,N_21674,N_21505);
xnor U22669 (N_22669,N_21969,N_21389);
nor U22670 (N_22670,N_21534,N_21737);
xnor U22671 (N_22671,N_21228,N_21980);
xnor U22672 (N_22672,N_21301,N_21726);
nand U22673 (N_22673,N_21241,N_21371);
or U22674 (N_22674,N_21998,N_21593);
nand U22675 (N_22675,N_21272,N_21734);
or U22676 (N_22676,N_21063,N_21782);
and U22677 (N_22677,N_21613,N_21773);
or U22678 (N_22678,N_21625,N_21742);
xnor U22679 (N_22679,N_21229,N_21667);
nand U22680 (N_22680,N_21618,N_21930);
nor U22681 (N_22681,N_21749,N_21829);
and U22682 (N_22682,N_21492,N_21342);
xnor U22683 (N_22683,N_21043,N_21250);
or U22684 (N_22684,N_21609,N_21200);
or U22685 (N_22685,N_21856,N_21764);
and U22686 (N_22686,N_21022,N_21269);
nor U22687 (N_22687,N_21922,N_21536);
and U22688 (N_22688,N_21572,N_21017);
nor U22689 (N_22689,N_21754,N_21597);
nand U22690 (N_22690,N_21971,N_21309);
and U22691 (N_22691,N_21271,N_21639);
and U22692 (N_22692,N_21217,N_21816);
xnor U22693 (N_22693,N_21175,N_21285);
or U22694 (N_22694,N_21311,N_21165);
nor U22695 (N_22695,N_21651,N_21383);
nand U22696 (N_22696,N_21837,N_21319);
or U22697 (N_22697,N_21454,N_21628);
and U22698 (N_22698,N_21248,N_21232);
nand U22699 (N_22699,N_21244,N_21399);
and U22700 (N_22700,N_21571,N_21859);
or U22701 (N_22701,N_21161,N_21956);
and U22702 (N_22702,N_21175,N_21071);
and U22703 (N_22703,N_21667,N_21405);
nor U22704 (N_22704,N_21172,N_21939);
xor U22705 (N_22705,N_21619,N_21900);
and U22706 (N_22706,N_21229,N_21712);
and U22707 (N_22707,N_21445,N_21802);
nand U22708 (N_22708,N_21343,N_21720);
nand U22709 (N_22709,N_21982,N_21708);
nor U22710 (N_22710,N_21147,N_21005);
nor U22711 (N_22711,N_21401,N_21373);
xor U22712 (N_22712,N_21065,N_21886);
and U22713 (N_22713,N_21065,N_21937);
and U22714 (N_22714,N_21368,N_21405);
nand U22715 (N_22715,N_21086,N_21069);
nand U22716 (N_22716,N_21626,N_21433);
nand U22717 (N_22717,N_21385,N_21274);
nor U22718 (N_22718,N_21607,N_21711);
or U22719 (N_22719,N_21357,N_21131);
nand U22720 (N_22720,N_21466,N_21610);
nand U22721 (N_22721,N_21851,N_21572);
or U22722 (N_22722,N_21344,N_21286);
and U22723 (N_22723,N_21502,N_21053);
xnor U22724 (N_22724,N_21563,N_21256);
or U22725 (N_22725,N_21488,N_21358);
nand U22726 (N_22726,N_21562,N_21590);
and U22727 (N_22727,N_21654,N_21164);
and U22728 (N_22728,N_21337,N_21840);
xnor U22729 (N_22729,N_21365,N_21775);
xor U22730 (N_22730,N_21963,N_21855);
nand U22731 (N_22731,N_21315,N_21269);
nor U22732 (N_22732,N_21858,N_21631);
xnor U22733 (N_22733,N_21086,N_21504);
nand U22734 (N_22734,N_21880,N_21495);
xor U22735 (N_22735,N_21452,N_21127);
nor U22736 (N_22736,N_21428,N_21675);
xnor U22737 (N_22737,N_21146,N_21355);
xor U22738 (N_22738,N_21011,N_21463);
xnor U22739 (N_22739,N_21428,N_21136);
and U22740 (N_22740,N_21768,N_21567);
nand U22741 (N_22741,N_21551,N_21209);
and U22742 (N_22742,N_21770,N_21935);
or U22743 (N_22743,N_21935,N_21998);
and U22744 (N_22744,N_21588,N_21227);
nor U22745 (N_22745,N_21481,N_21125);
nor U22746 (N_22746,N_21597,N_21902);
nor U22747 (N_22747,N_21708,N_21316);
nand U22748 (N_22748,N_21585,N_21557);
or U22749 (N_22749,N_21841,N_21922);
xnor U22750 (N_22750,N_21269,N_21505);
or U22751 (N_22751,N_21888,N_21932);
nand U22752 (N_22752,N_21371,N_21321);
or U22753 (N_22753,N_21376,N_21425);
or U22754 (N_22754,N_21650,N_21222);
nand U22755 (N_22755,N_21968,N_21475);
and U22756 (N_22756,N_21273,N_21723);
nor U22757 (N_22757,N_21493,N_21758);
or U22758 (N_22758,N_21448,N_21422);
nor U22759 (N_22759,N_21538,N_21511);
or U22760 (N_22760,N_21137,N_21951);
nand U22761 (N_22761,N_21055,N_21893);
nor U22762 (N_22762,N_21926,N_21734);
nand U22763 (N_22763,N_21842,N_21432);
xnor U22764 (N_22764,N_21440,N_21333);
and U22765 (N_22765,N_21365,N_21790);
xor U22766 (N_22766,N_21963,N_21001);
or U22767 (N_22767,N_21843,N_21330);
xnor U22768 (N_22768,N_21141,N_21726);
xnor U22769 (N_22769,N_21704,N_21205);
xor U22770 (N_22770,N_21555,N_21814);
nand U22771 (N_22771,N_21669,N_21626);
xnor U22772 (N_22772,N_21710,N_21815);
or U22773 (N_22773,N_21735,N_21145);
nor U22774 (N_22774,N_21401,N_21789);
and U22775 (N_22775,N_21762,N_21595);
nor U22776 (N_22776,N_21404,N_21295);
nor U22777 (N_22777,N_21538,N_21727);
nor U22778 (N_22778,N_21060,N_21092);
nand U22779 (N_22779,N_21995,N_21242);
nand U22780 (N_22780,N_21277,N_21083);
nor U22781 (N_22781,N_21679,N_21078);
xor U22782 (N_22782,N_21658,N_21315);
nor U22783 (N_22783,N_21944,N_21100);
nand U22784 (N_22784,N_21620,N_21857);
or U22785 (N_22785,N_21053,N_21281);
xnor U22786 (N_22786,N_21119,N_21513);
nor U22787 (N_22787,N_21358,N_21570);
nand U22788 (N_22788,N_21788,N_21808);
nor U22789 (N_22789,N_21468,N_21881);
xor U22790 (N_22790,N_21289,N_21838);
nand U22791 (N_22791,N_21964,N_21647);
nor U22792 (N_22792,N_21657,N_21521);
nor U22793 (N_22793,N_21565,N_21838);
xnor U22794 (N_22794,N_21471,N_21834);
xor U22795 (N_22795,N_21734,N_21415);
or U22796 (N_22796,N_21647,N_21896);
nor U22797 (N_22797,N_21174,N_21985);
nand U22798 (N_22798,N_21568,N_21024);
and U22799 (N_22799,N_21287,N_21676);
nand U22800 (N_22800,N_21135,N_21579);
nor U22801 (N_22801,N_21994,N_21846);
or U22802 (N_22802,N_21998,N_21713);
or U22803 (N_22803,N_21019,N_21041);
nor U22804 (N_22804,N_21119,N_21148);
xor U22805 (N_22805,N_21524,N_21893);
or U22806 (N_22806,N_21786,N_21268);
or U22807 (N_22807,N_21060,N_21489);
or U22808 (N_22808,N_21867,N_21369);
and U22809 (N_22809,N_21309,N_21944);
and U22810 (N_22810,N_21196,N_21291);
xor U22811 (N_22811,N_21768,N_21949);
nor U22812 (N_22812,N_21537,N_21885);
or U22813 (N_22813,N_21369,N_21301);
or U22814 (N_22814,N_21448,N_21789);
xnor U22815 (N_22815,N_21272,N_21319);
or U22816 (N_22816,N_21352,N_21496);
or U22817 (N_22817,N_21890,N_21789);
xor U22818 (N_22818,N_21589,N_21208);
nand U22819 (N_22819,N_21690,N_21092);
and U22820 (N_22820,N_21245,N_21738);
nand U22821 (N_22821,N_21610,N_21609);
and U22822 (N_22822,N_21570,N_21963);
or U22823 (N_22823,N_21909,N_21530);
nand U22824 (N_22824,N_21357,N_21988);
nor U22825 (N_22825,N_21865,N_21354);
and U22826 (N_22826,N_21344,N_21425);
or U22827 (N_22827,N_21012,N_21497);
nand U22828 (N_22828,N_21474,N_21747);
xnor U22829 (N_22829,N_21859,N_21673);
nand U22830 (N_22830,N_21023,N_21759);
xor U22831 (N_22831,N_21143,N_21633);
and U22832 (N_22832,N_21479,N_21884);
xor U22833 (N_22833,N_21301,N_21272);
nor U22834 (N_22834,N_21522,N_21748);
xor U22835 (N_22835,N_21209,N_21631);
nand U22836 (N_22836,N_21306,N_21592);
or U22837 (N_22837,N_21743,N_21544);
nand U22838 (N_22838,N_21557,N_21737);
xnor U22839 (N_22839,N_21389,N_21597);
nor U22840 (N_22840,N_21326,N_21883);
or U22841 (N_22841,N_21544,N_21067);
nand U22842 (N_22842,N_21394,N_21711);
or U22843 (N_22843,N_21958,N_21202);
and U22844 (N_22844,N_21870,N_21536);
or U22845 (N_22845,N_21915,N_21506);
and U22846 (N_22846,N_21786,N_21086);
xnor U22847 (N_22847,N_21501,N_21817);
xor U22848 (N_22848,N_21514,N_21731);
nor U22849 (N_22849,N_21378,N_21864);
or U22850 (N_22850,N_21086,N_21197);
xnor U22851 (N_22851,N_21764,N_21374);
and U22852 (N_22852,N_21672,N_21349);
nand U22853 (N_22853,N_21546,N_21027);
or U22854 (N_22854,N_21789,N_21018);
xnor U22855 (N_22855,N_21244,N_21217);
nor U22856 (N_22856,N_21078,N_21136);
nand U22857 (N_22857,N_21298,N_21465);
nand U22858 (N_22858,N_21297,N_21603);
nand U22859 (N_22859,N_21968,N_21099);
or U22860 (N_22860,N_21582,N_21655);
nor U22861 (N_22861,N_21542,N_21216);
and U22862 (N_22862,N_21253,N_21591);
nor U22863 (N_22863,N_21536,N_21806);
or U22864 (N_22864,N_21693,N_21229);
or U22865 (N_22865,N_21084,N_21193);
or U22866 (N_22866,N_21325,N_21434);
nand U22867 (N_22867,N_21801,N_21231);
xor U22868 (N_22868,N_21019,N_21867);
and U22869 (N_22869,N_21290,N_21414);
or U22870 (N_22870,N_21899,N_21764);
xor U22871 (N_22871,N_21487,N_21229);
xnor U22872 (N_22872,N_21952,N_21271);
nand U22873 (N_22873,N_21894,N_21671);
xnor U22874 (N_22874,N_21716,N_21722);
or U22875 (N_22875,N_21515,N_21205);
or U22876 (N_22876,N_21575,N_21068);
and U22877 (N_22877,N_21769,N_21207);
and U22878 (N_22878,N_21640,N_21546);
nand U22879 (N_22879,N_21198,N_21261);
nor U22880 (N_22880,N_21026,N_21584);
nor U22881 (N_22881,N_21225,N_21746);
nor U22882 (N_22882,N_21168,N_21336);
and U22883 (N_22883,N_21425,N_21538);
xor U22884 (N_22884,N_21215,N_21660);
xnor U22885 (N_22885,N_21636,N_21329);
or U22886 (N_22886,N_21296,N_21554);
nand U22887 (N_22887,N_21654,N_21132);
xor U22888 (N_22888,N_21336,N_21516);
nor U22889 (N_22889,N_21171,N_21207);
nor U22890 (N_22890,N_21855,N_21760);
xor U22891 (N_22891,N_21424,N_21634);
nor U22892 (N_22892,N_21495,N_21924);
nand U22893 (N_22893,N_21471,N_21264);
or U22894 (N_22894,N_21147,N_21170);
nand U22895 (N_22895,N_21997,N_21069);
xor U22896 (N_22896,N_21476,N_21849);
or U22897 (N_22897,N_21621,N_21525);
or U22898 (N_22898,N_21964,N_21671);
xnor U22899 (N_22899,N_21787,N_21703);
nand U22900 (N_22900,N_21596,N_21796);
and U22901 (N_22901,N_21659,N_21606);
or U22902 (N_22902,N_21021,N_21058);
nor U22903 (N_22903,N_21741,N_21188);
or U22904 (N_22904,N_21581,N_21125);
xnor U22905 (N_22905,N_21890,N_21548);
nor U22906 (N_22906,N_21968,N_21342);
and U22907 (N_22907,N_21313,N_21247);
or U22908 (N_22908,N_21916,N_21399);
and U22909 (N_22909,N_21870,N_21927);
and U22910 (N_22910,N_21902,N_21862);
nor U22911 (N_22911,N_21168,N_21655);
and U22912 (N_22912,N_21085,N_21378);
xor U22913 (N_22913,N_21873,N_21929);
nand U22914 (N_22914,N_21019,N_21721);
xor U22915 (N_22915,N_21035,N_21619);
or U22916 (N_22916,N_21221,N_21465);
or U22917 (N_22917,N_21173,N_21973);
nor U22918 (N_22918,N_21943,N_21102);
or U22919 (N_22919,N_21118,N_21678);
and U22920 (N_22920,N_21602,N_21407);
xnor U22921 (N_22921,N_21413,N_21156);
nor U22922 (N_22922,N_21605,N_21907);
or U22923 (N_22923,N_21693,N_21592);
and U22924 (N_22924,N_21428,N_21159);
nand U22925 (N_22925,N_21923,N_21837);
and U22926 (N_22926,N_21462,N_21542);
and U22927 (N_22927,N_21693,N_21826);
nor U22928 (N_22928,N_21024,N_21753);
nor U22929 (N_22929,N_21926,N_21915);
and U22930 (N_22930,N_21063,N_21632);
xnor U22931 (N_22931,N_21568,N_21152);
nand U22932 (N_22932,N_21376,N_21946);
nand U22933 (N_22933,N_21709,N_21928);
and U22934 (N_22934,N_21077,N_21164);
nor U22935 (N_22935,N_21203,N_21585);
and U22936 (N_22936,N_21702,N_21152);
and U22937 (N_22937,N_21484,N_21102);
nand U22938 (N_22938,N_21645,N_21615);
and U22939 (N_22939,N_21910,N_21124);
or U22940 (N_22940,N_21422,N_21906);
or U22941 (N_22941,N_21208,N_21345);
nor U22942 (N_22942,N_21369,N_21924);
and U22943 (N_22943,N_21800,N_21644);
nand U22944 (N_22944,N_21106,N_21779);
or U22945 (N_22945,N_21760,N_21890);
nor U22946 (N_22946,N_21793,N_21456);
or U22947 (N_22947,N_21103,N_21047);
nor U22948 (N_22948,N_21801,N_21426);
or U22949 (N_22949,N_21758,N_21183);
or U22950 (N_22950,N_21564,N_21173);
xnor U22951 (N_22951,N_21321,N_21420);
nor U22952 (N_22952,N_21376,N_21418);
nand U22953 (N_22953,N_21855,N_21906);
or U22954 (N_22954,N_21654,N_21150);
and U22955 (N_22955,N_21182,N_21638);
xor U22956 (N_22956,N_21034,N_21495);
or U22957 (N_22957,N_21145,N_21399);
nor U22958 (N_22958,N_21506,N_21003);
xor U22959 (N_22959,N_21446,N_21764);
and U22960 (N_22960,N_21755,N_21712);
xnor U22961 (N_22961,N_21209,N_21076);
nor U22962 (N_22962,N_21241,N_21294);
and U22963 (N_22963,N_21611,N_21794);
or U22964 (N_22964,N_21008,N_21571);
nand U22965 (N_22965,N_21839,N_21342);
or U22966 (N_22966,N_21729,N_21580);
and U22967 (N_22967,N_21275,N_21716);
nor U22968 (N_22968,N_21801,N_21098);
and U22969 (N_22969,N_21217,N_21799);
or U22970 (N_22970,N_21118,N_21950);
and U22971 (N_22971,N_21155,N_21482);
nand U22972 (N_22972,N_21224,N_21327);
xor U22973 (N_22973,N_21703,N_21598);
or U22974 (N_22974,N_21401,N_21313);
xor U22975 (N_22975,N_21955,N_21962);
xor U22976 (N_22976,N_21128,N_21523);
and U22977 (N_22977,N_21817,N_21235);
and U22978 (N_22978,N_21832,N_21433);
xnor U22979 (N_22979,N_21089,N_21338);
nand U22980 (N_22980,N_21656,N_21385);
and U22981 (N_22981,N_21109,N_21129);
xor U22982 (N_22982,N_21786,N_21891);
and U22983 (N_22983,N_21892,N_21049);
nor U22984 (N_22984,N_21017,N_21829);
and U22985 (N_22985,N_21942,N_21939);
nor U22986 (N_22986,N_21774,N_21008);
xnor U22987 (N_22987,N_21734,N_21043);
or U22988 (N_22988,N_21406,N_21844);
or U22989 (N_22989,N_21827,N_21080);
nor U22990 (N_22990,N_21248,N_21017);
nor U22991 (N_22991,N_21026,N_21955);
or U22992 (N_22992,N_21274,N_21826);
nor U22993 (N_22993,N_21239,N_21712);
nand U22994 (N_22994,N_21532,N_21214);
and U22995 (N_22995,N_21884,N_21093);
nand U22996 (N_22996,N_21051,N_21603);
nand U22997 (N_22997,N_21101,N_21489);
or U22998 (N_22998,N_21297,N_21457);
xor U22999 (N_22999,N_21940,N_21712);
or U23000 (N_23000,N_22370,N_22963);
nand U23001 (N_23001,N_22396,N_22414);
xnor U23002 (N_23002,N_22031,N_22090);
and U23003 (N_23003,N_22186,N_22210);
and U23004 (N_23004,N_22857,N_22206);
and U23005 (N_23005,N_22127,N_22093);
and U23006 (N_23006,N_22136,N_22696);
or U23007 (N_23007,N_22431,N_22767);
nand U23008 (N_23008,N_22001,N_22873);
or U23009 (N_23009,N_22656,N_22713);
nand U23010 (N_23010,N_22759,N_22267);
nor U23011 (N_23011,N_22260,N_22983);
or U23012 (N_23012,N_22307,N_22363);
nor U23013 (N_23013,N_22649,N_22567);
or U23014 (N_23014,N_22705,N_22073);
and U23015 (N_23015,N_22992,N_22464);
nor U23016 (N_23016,N_22999,N_22636);
xnor U23017 (N_23017,N_22651,N_22671);
or U23018 (N_23018,N_22087,N_22768);
nor U23019 (N_23019,N_22848,N_22965);
and U23020 (N_23020,N_22347,N_22766);
or U23021 (N_23021,N_22381,N_22786);
and U23022 (N_23022,N_22161,N_22410);
or U23023 (N_23023,N_22368,N_22351);
nor U23024 (N_23024,N_22187,N_22874);
or U23025 (N_23025,N_22703,N_22392);
or U23026 (N_23026,N_22015,N_22379);
nand U23027 (N_23027,N_22164,N_22064);
nor U23028 (N_23028,N_22434,N_22994);
xor U23029 (N_23029,N_22466,N_22953);
and U23030 (N_23030,N_22911,N_22721);
and U23031 (N_23031,N_22035,N_22739);
and U23032 (N_23032,N_22184,N_22674);
and U23033 (N_23033,N_22909,N_22350);
and U23034 (N_23034,N_22938,N_22074);
nor U23035 (N_23035,N_22476,N_22216);
xor U23036 (N_23036,N_22812,N_22889);
nor U23037 (N_23037,N_22398,N_22844);
xnor U23038 (N_23038,N_22185,N_22592);
nand U23039 (N_23039,N_22927,N_22198);
xnor U23040 (N_23040,N_22383,N_22153);
nand U23041 (N_23041,N_22457,N_22319);
nor U23042 (N_23042,N_22838,N_22180);
and U23043 (N_23043,N_22227,N_22795);
nand U23044 (N_23044,N_22566,N_22724);
nand U23045 (N_23045,N_22700,N_22339);
xnor U23046 (N_23046,N_22106,N_22968);
xor U23047 (N_23047,N_22715,N_22317);
xor U23048 (N_23048,N_22482,N_22799);
or U23049 (N_23049,N_22560,N_22254);
or U23050 (N_23050,N_22104,N_22382);
nor U23051 (N_23051,N_22896,N_22587);
xnor U23052 (N_23052,N_22808,N_22862);
nand U23053 (N_23053,N_22833,N_22331);
nor U23054 (N_23054,N_22039,N_22130);
xnor U23055 (N_23055,N_22509,N_22883);
nor U23056 (N_23056,N_22418,N_22310);
xnor U23057 (N_23057,N_22367,N_22289);
and U23058 (N_23058,N_22910,N_22668);
nor U23059 (N_23059,N_22459,N_22046);
xor U23060 (N_23060,N_22283,N_22754);
xnor U23061 (N_23061,N_22109,N_22977);
nand U23062 (N_23062,N_22384,N_22607);
xnor U23063 (N_23063,N_22040,N_22286);
and U23064 (N_23064,N_22913,N_22742);
nand U23065 (N_23065,N_22866,N_22257);
xnor U23066 (N_23066,N_22010,N_22438);
xor U23067 (N_23067,N_22669,N_22270);
xor U23068 (N_23068,N_22121,N_22652);
nor U23069 (N_23069,N_22232,N_22547);
or U23070 (N_23070,N_22655,N_22624);
nor U23071 (N_23071,N_22784,N_22043);
nand U23072 (N_23072,N_22507,N_22411);
and U23073 (N_23073,N_22262,N_22579);
nand U23074 (N_23074,N_22907,N_22247);
and U23075 (N_23075,N_22013,N_22203);
nand U23076 (N_23076,N_22179,N_22020);
nand U23077 (N_23077,N_22847,N_22234);
or U23078 (N_23078,N_22901,N_22060);
nor U23079 (N_23079,N_22924,N_22058);
xor U23080 (N_23080,N_22231,N_22535);
xnor U23081 (N_23081,N_22026,N_22108);
nor U23082 (N_23082,N_22630,N_22248);
nor U23083 (N_23083,N_22814,N_22226);
nor U23084 (N_23084,N_22555,N_22923);
xnor U23085 (N_23085,N_22008,N_22191);
and U23086 (N_23086,N_22449,N_22735);
nor U23087 (N_23087,N_22024,N_22794);
and U23088 (N_23088,N_22675,N_22285);
nand U23089 (N_23089,N_22325,N_22877);
xnor U23090 (N_23090,N_22036,N_22249);
and U23091 (N_23091,N_22855,N_22710);
nor U23092 (N_23092,N_22214,N_22810);
xor U23093 (N_23093,N_22068,N_22236);
nand U23094 (N_23094,N_22773,N_22460);
and U23095 (N_23095,N_22830,N_22959);
nor U23096 (N_23096,N_22564,N_22229);
and U23097 (N_23097,N_22776,N_22346);
nand U23098 (N_23098,N_22215,N_22276);
xor U23099 (N_23099,N_22619,N_22540);
nor U23100 (N_23100,N_22912,N_22683);
and U23101 (N_23101,N_22193,N_22801);
and U23102 (N_23102,N_22691,N_22686);
nor U23103 (N_23103,N_22103,N_22741);
or U23104 (N_23104,N_22320,N_22097);
nor U23105 (N_23105,N_22712,N_22296);
nor U23106 (N_23106,N_22006,N_22306);
or U23107 (N_23107,N_22168,N_22771);
nand U23108 (N_23108,N_22205,N_22644);
and U23109 (N_23109,N_22360,N_22358);
nor U23110 (N_23110,N_22561,N_22932);
nand U23111 (N_23111,N_22688,N_22281);
nand U23112 (N_23112,N_22080,N_22760);
nand U23113 (N_23113,N_22979,N_22167);
nand U23114 (N_23114,N_22195,N_22850);
and U23115 (N_23115,N_22775,N_22643);
nand U23116 (N_23116,N_22872,N_22666);
nor U23117 (N_23117,N_22718,N_22878);
or U23118 (N_23118,N_22077,N_22621);
or U23119 (N_23119,N_22305,N_22991);
xor U23120 (N_23120,N_22982,N_22615);
and U23121 (N_23121,N_22625,N_22072);
nor U23122 (N_23122,N_22242,N_22494);
and U23123 (N_23123,N_22985,N_22793);
or U23124 (N_23124,N_22403,N_22559);
nor U23125 (N_23125,N_22616,N_22415);
or U23126 (N_23126,N_22056,N_22879);
or U23127 (N_23127,N_22327,N_22653);
xor U23128 (N_23128,N_22817,N_22419);
and U23129 (N_23129,N_22960,N_22421);
xor U23130 (N_23130,N_22397,N_22785);
or U23131 (N_23131,N_22684,N_22119);
xnor U23132 (N_23132,N_22638,N_22528);
and U23133 (N_23133,N_22554,N_22552);
nor U23134 (N_23134,N_22445,N_22011);
or U23135 (N_23135,N_22563,N_22828);
and U23136 (N_23136,N_22311,N_22033);
nand U23137 (N_23137,N_22526,N_22943);
or U23138 (N_23138,N_22192,N_22551);
or U23139 (N_23139,N_22882,N_22014);
nor U23140 (N_23140,N_22996,N_22299);
and U23141 (N_23141,N_22536,N_22219);
xnor U23142 (N_23142,N_22030,N_22098);
nand U23143 (N_23143,N_22617,N_22291);
or U23144 (N_23144,N_22832,N_22629);
xor U23145 (N_23145,N_22394,N_22697);
nand U23146 (N_23146,N_22321,N_22524);
nand U23147 (N_23147,N_22545,N_22333);
or U23148 (N_23148,N_22980,N_22730);
nor U23149 (N_23149,N_22239,N_22870);
nand U23150 (N_23150,N_22679,N_22264);
or U23151 (N_23151,N_22677,N_22726);
nor U23152 (N_23152,N_22542,N_22986);
xnor U23153 (N_23153,N_22399,N_22225);
or U23154 (N_23154,N_22637,N_22322);
xor U23155 (N_23155,N_22701,N_22208);
nand U23156 (N_23156,N_22544,N_22894);
xor U23157 (N_23157,N_22940,N_22261);
and U23158 (N_23158,N_22978,N_22600);
and U23159 (N_23159,N_22790,N_22173);
and U23160 (N_23160,N_22070,N_22114);
nor U23161 (N_23161,N_22928,N_22869);
nand U23162 (N_23162,N_22608,N_22361);
or U23163 (N_23163,N_22471,N_22251);
nand U23164 (N_23164,N_22217,N_22211);
xor U23165 (N_23165,N_22865,N_22473);
xor U23166 (N_23166,N_22300,N_22484);
nor U23167 (N_23167,N_22720,N_22271);
nand U23168 (N_23168,N_22355,N_22533);
nor U23169 (N_23169,N_22606,N_22377);
xor U23170 (N_23170,N_22425,N_22572);
and U23171 (N_23171,N_22266,N_22273);
or U23172 (N_23172,N_22681,N_22084);
nand U23173 (N_23173,N_22244,N_22452);
xor U23174 (N_23174,N_22420,N_22532);
or U23175 (N_23175,N_22915,N_22349);
xor U23176 (N_23176,N_22102,N_22038);
or U23177 (N_23177,N_22824,N_22086);
nand U23178 (N_23178,N_22171,N_22576);
nand U23179 (N_23179,N_22632,N_22821);
xnor U23180 (N_23180,N_22791,N_22788);
and U23181 (N_23181,N_22424,N_22843);
or U23182 (N_23182,N_22849,N_22825);
nand U23183 (N_23183,N_22504,N_22100);
nor U23184 (N_23184,N_22258,N_22069);
or U23185 (N_23185,N_22378,N_22054);
nor U23186 (N_23186,N_22190,N_22277);
nor U23187 (N_23187,N_22096,N_22336);
or U23188 (N_23188,N_22151,N_22479);
nor U23189 (N_23189,N_22406,N_22057);
nand U23190 (N_23190,N_22642,N_22240);
nand U23191 (N_23191,N_22495,N_22517);
nor U23192 (N_23192,N_22920,N_22380);
or U23193 (N_23193,N_22498,N_22160);
or U23194 (N_23194,N_22212,N_22856);
and U23195 (N_23195,N_22423,N_22166);
nand U23196 (N_23196,N_22172,N_22835);
or U23197 (N_23197,N_22998,N_22597);
nand U23198 (N_23198,N_22340,N_22680);
nand U23199 (N_23199,N_22993,N_22816);
nand U23200 (N_23200,N_22772,N_22255);
xnor U23201 (N_23201,N_22548,N_22950);
nand U23202 (N_23202,N_22780,N_22512);
nand U23203 (N_23203,N_22763,N_22593);
xnor U23204 (N_23204,N_22891,N_22961);
or U23205 (N_23205,N_22954,N_22525);
or U23206 (N_23206,N_22238,N_22111);
and U23207 (N_23207,N_22826,N_22292);
nor U23208 (N_23208,N_22926,N_22221);
or U23209 (N_23209,N_22553,N_22188);
or U23210 (N_23210,N_22189,N_22487);
and U23211 (N_23211,N_22076,N_22122);
or U23212 (N_23212,N_22156,N_22018);
xor U23213 (N_23213,N_22400,N_22521);
and U23214 (N_23214,N_22141,N_22829);
xnor U23215 (N_23215,N_22515,N_22357);
nor U23216 (N_23216,N_22751,N_22142);
nor U23217 (N_23217,N_22749,N_22967);
and U23218 (N_23218,N_22520,N_22888);
xor U23219 (N_23219,N_22485,N_22138);
nor U23220 (N_23220,N_22246,N_22746);
nand U23221 (N_23221,N_22622,N_22032);
xor U23222 (N_23222,N_22113,N_22628);
nand U23223 (N_23223,N_22342,N_22385);
and U23224 (N_23224,N_22009,N_22748);
xnor U23225 (N_23225,N_22634,N_22448);
or U23226 (N_23226,N_22078,N_22519);
xor U23227 (N_23227,N_22887,N_22609);
or U23228 (N_23228,N_22029,N_22472);
or U23229 (N_23229,N_22204,N_22750);
and U23230 (N_23230,N_22695,N_22233);
xor U23231 (N_23231,N_22401,N_22662);
xnor U23232 (N_23232,N_22989,N_22842);
and U23233 (N_23233,N_22729,N_22152);
xor U23234 (N_23234,N_22369,N_22470);
nand U23235 (N_23235,N_22618,N_22129);
and U23236 (N_23236,N_22302,N_22478);
nor U23237 (N_23237,N_22981,N_22324);
nand U23238 (N_23238,N_22755,N_22667);
nor U23239 (N_23239,N_22962,N_22620);
nor U23240 (N_23240,N_22335,N_22326);
nand U23241 (N_23241,N_22209,N_22605);
xnor U23242 (N_23242,N_22025,N_22241);
xor U23243 (N_23243,N_22427,N_22177);
nand U23244 (N_23244,N_22687,N_22163);
or U23245 (N_23245,N_22997,N_22259);
nand U23246 (N_23246,N_22491,N_22287);
and U23247 (N_23247,N_22461,N_22933);
nor U23248 (N_23248,N_22575,N_22885);
and U23249 (N_23249,N_22481,N_22207);
nand U23250 (N_23250,N_22412,N_22770);
nor U23251 (N_23251,N_22016,N_22301);
xor U23252 (N_23252,N_22139,N_22725);
and U23253 (N_23253,N_22947,N_22178);
and U23254 (N_23254,N_22774,N_22316);
or U23255 (N_23255,N_22493,N_22557);
nand U23256 (N_23256,N_22274,N_22441);
nand U23257 (N_23257,N_22343,N_22514);
nor U23258 (N_23258,N_22792,N_22456);
nand U23259 (N_23259,N_22511,N_22131);
nand U23260 (N_23260,N_22182,N_22904);
nand U23261 (N_23261,N_22323,N_22717);
nor U23262 (N_23262,N_22871,N_22465);
xor U23263 (N_23263,N_22603,N_22577);
xnor U23264 (N_23264,N_22099,N_22762);
or U23265 (N_23265,N_22462,N_22948);
or U23266 (N_23266,N_22447,N_22732);
and U23267 (N_23267,N_22580,N_22846);
or U23268 (N_23268,N_22585,N_22574);
or U23269 (N_23269,N_22454,N_22995);
xor U23270 (N_23270,N_22143,N_22081);
nand U23271 (N_23271,N_22467,N_22646);
xor U23272 (N_23272,N_22796,N_22516);
xor U23273 (N_23273,N_22777,N_22416);
nor U23274 (N_23274,N_22974,N_22731);
nand U23275 (N_23275,N_22807,N_22641);
nor U23276 (N_23276,N_22132,N_22003);
nand U23277 (N_23277,N_22635,N_22365);
nor U23278 (N_23278,N_22558,N_22451);
and U23279 (N_23279,N_22845,N_22089);
xnor U23280 (N_23280,N_22312,N_22529);
xnor U23281 (N_23281,N_22645,N_22437);
or U23282 (N_23282,N_22329,N_22711);
nor U23283 (N_23283,N_22602,N_22303);
nand U23284 (N_23284,N_22530,N_22657);
or U23285 (N_23285,N_22126,N_22155);
and U23286 (N_23286,N_22738,N_22659);
nor U23287 (N_23287,N_22123,N_22027);
nand U23288 (N_23288,N_22714,N_22578);
nand U23289 (N_23289,N_22744,N_22395);
xnor U23290 (N_23290,N_22988,N_22658);
and U23291 (N_23291,N_22028,N_22964);
xor U23292 (N_23292,N_22391,N_22150);
or U23293 (N_23293,N_22408,N_22931);
and U23294 (N_23294,N_22094,N_22144);
xor U23295 (N_23295,N_22702,N_22747);
xor U23296 (N_23296,N_22941,N_22263);
xnor U23297 (N_23297,N_22275,N_22699);
xnor U23298 (N_23298,N_22868,N_22269);
xor U23299 (N_23299,N_22047,N_22764);
nand U23300 (N_23300,N_22146,N_22704);
nand U23301 (N_23301,N_22145,N_22468);
and U23302 (N_23302,N_22463,N_22531);
nor U23303 (N_23303,N_22815,N_22095);
and U23304 (N_23304,N_22134,N_22065);
xor U23305 (N_23305,N_22405,N_22886);
nor U23306 (N_23306,N_22042,N_22908);
nand U23307 (N_23307,N_22804,N_22958);
xnor U23308 (N_23308,N_22213,N_22112);
nand U23309 (N_23309,N_22693,N_22348);
and U23310 (N_23310,N_22728,N_22413);
nor U23311 (N_23311,N_22949,N_22951);
and U23312 (N_23312,N_22435,N_22797);
nor U23313 (N_23313,N_22475,N_22522);
and U23314 (N_23314,N_22389,N_22716);
or U23315 (N_23315,N_22176,N_22082);
nand U23316 (N_23316,N_22256,N_22137);
xnor U23317 (N_23317,N_22497,N_22012);
xnor U23318 (N_23318,N_22672,N_22839);
and U23319 (N_23319,N_22061,N_22297);
and U23320 (N_23320,N_22194,N_22929);
nand U23321 (N_23321,N_22598,N_22243);
or U23322 (N_23322,N_22085,N_22279);
or U23323 (N_23323,N_22477,N_22053);
xnor U23324 (N_23324,N_22737,N_22903);
nand U23325 (N_23325,N_22854,N_22823);
or U23326 (N_23326,N_22133,N_22694);
or U23327 (N_23327,N_22573,N_22809);
and U23328 (N_23328,N_22811,N_22633);
xor U23329 (N_23329,N_22976,N_22892);
nor U23330 (N_23330,N_22984,N_22366);
nor U23331 (N_23331,N_22957,N_22935);
nor U23332 (N_23332,N_22059,N_22353);
xnor U23333 (N_23333,N_22362,N_22092);
xor U23334 (N_23334,N_22761,N_22304);
nand U23335 (N_23335,N_22613,N_22181);
or U23336 (N_23336,N_22157,N_22050);
nor U23337 (N_23337,N_22987,N_22590);
xnor U23338 (N_23338,N_22594,N_22990);
nor U23339 (N_23339,N_22083,N_22373);
xnor U23340 (N_23340,N_22752,N_22818);
nor U23341 (N_23341,N_22149,N_22591);
and U23342 (N_23342,N_22510,N_22546);
xnor U23343 (N_23343,N_22228,N_22805);
xnor U23344 (N_23344,N_22062,N_22110);
nor U23345 (N_23345,N_22402,N_22734);
or U23346 (N_23346,N_22867,N_22428);
nand U23347 (N_23347,N_22334,N_22864);
and U23348 (N_23348,N_22019,N_22282);
or U23349 (N_23349,N_22115,N_22944);
xnor U23350 (N_23350,N_22541,N_22650);
nor U23351 (N_23351,N_22822,N_22197);
xor U23352 (N_23352,N_22690,N_22937);
nand U23353 (N_23353,N_22075,N_22543);
or U23354 (N_23354,N_22158,N_22364);
nand U23355 (N_23355,N_22798,N_22387);
nand U23356 (N_23356,N_22819,N_22202);
nor U23357 (N_23357,N_22930,N_22945);
nand U23358 (N_23358,N_22740,N_22709);
or U23359 (N_23359,N_22806,N_22841);
and U23360 (N_23360,N_22736,N_22480);
nand U23361 (N_23361,N_22309,N_22765);
and U23362 (N_23362,N_22200,N_22523);
nand U23363 (N_23363,N_22527,N_22660);
nand U23364 (N_23364,N_22165,N_22569);
and U23365 (N_23365,N_22921,N_22422);
or U23366 (N_23366,N_22169,N_22128);
or U23367 (N_23367,N_22631,N_22469);
or U23368 (N_23368,N_22670,N_22582);
nand U23369 (N_23369,N_22884,N_22439);
and U23370 (N_23370,N_22022,N_22827);
or U23371 (N_23371,N_22781,N_22837);
xor U23372 (N_23372,N_22925,N_22583);
xnor U23373 (N_23373,N_22272,N_22237);
nand U23374 (N_23374,N_22021,N_22224);
or U23375 (N_23375,N_22374,N_22639);
nor U23376 (N_23376,N_22290,N_22159);
and U23377 (N_23377,N_22223,N_22154);
or U23378 (N_23378,N_22919,N_22966);
nand U23379 (N_23379,N_22596,N_22895);
xor U23380 (N_23380,N_22971,N_22876);
xor U23381 (N_23381,N_22956,N_22783);
nor U23382 (N_23382,N_22235,N_22860);
and U23383 (N_23383,N_22778,N_22513);
and U23384 (N_23384,N_22492,N_22549);
nor U23385 (N_23385,N_22787,N_22034);
nor U23386 (N_23386,N_22426,N_22175);
and U23387 (N_23387,N_22386,N_22443);
and U23388 (N_23388,N_22442,N_22071);
and U23389 (N_23389,N_22004,N_22678);
nand U23390 (N_23390,N_22091,N_22486);
xnor U23391 (N_23391,N_22952,N_22488);
xnor U23392 (N_23392,N_22851,N_22664);
and U23393 (N_23393,N_22005,N_22922);
or U23394 (N_23394,N_22753,N_22565);
nor U23395 (N_23395,N_22359,N_22455);
or U23396 (N_23396,N_22893,N_22375);
and U23397 (N_23397,N_22496,N_22955);
and U23398 (N_23398,N_22432,N_22313);
and U23399 (N_23399,N_22673,N_22789);
and U23400 (N_23400,N_22682,N_22007);
xnor U23401 (N_23401,N_22328,N_22610);
nor U23402 (N_23402,N_22067,N_22218);
or U23403 (N_23403,N_22648,N_22782);
or U23404 (N_23404,N_22125,N_22390);
or U23405 (N_23405,N_22604,N_22581);
nand U23406 (N_23406,N_22972,N_22429);
and U23407 (N_23407,N_22330,N_22288);
nand U23408 (N_23408,N_22836,N_22483);
xnor U23409 (N_23409,N_22537,N_22852);
nor U23410 (N_23410,N_22404,N_22376);
xor U23411 (N_23411,N_22444,N_22101);
nand U23412 (N_23412,N_22183,N_22199);
or U23413 (N_23413,N_22758,N_22626);
xor U23414 (N_23414,N_22294,N_22332);
nand U23415 (N_23415,N_22708,N_22450);
nor U23416 (N_23416,N_22757,N_22140);
nand U23417 (N_23417,N_22474,N_22733);
nand U23418 (N_23418,N_22105,N_22501);
xnor U23419 (N_23419,N_22393,N_22707);
and U23420 (N_23420,N_22489,N_22352);
xnor U23421 (N_23421,N_22148,N_22875);
and U23422 (N_23422,N_22723,N_22859);
or U23423 (N_23423,N_22174,N_22906);
nor U23424 (N_23424,N_22663,N_22250);
xnor U23425 (N_23425,N_22820,N_22088);
and U23426 (N_23426,N_22041,N_22000);
nand U23427 (N_23427,N_22918,N_22506);
and U23428 (N_23428,N_22490,N_22356);
and U23429 (N_23429,N_22900,N_22905);
xor U23430 (N_23430,N_22409,N_22571);
or U23431 (N_23431,N_22252,N_22135);
or U23432 (N_23432,N_22245,N_22800);
or U23433 (N_23433,N_22124,N_22118);
nand U23434 (N_23434,N_22371,N_22314);
nor U23435 (N_23435,N_22831,N_22858);
nand U23436 (N_23436,N_22665,N_22881);
nor U23437 (N_23437,N_22341,N_22265);
nand U23438 (N_23438,N_22293,N_22916);
and U23439 (N_23439,N_22048,N_22969);
and U23440 (N_23440,N_22813,N_22756);
and U23441 (N_23441,N_22268,N_22942);
and U23442 (N_23442,N_22107,N_22201);
and U23443 (N_23443,N_22280,N_22589);
xnor U23444 (N_23444,N_22162,N_22898);
and U23445 (N_23445,N_22315,N_22970);
or U23446 (N_23446,N_22914,N_22647);
nor U23447 (N_23447,N_22433,N_22051);
and U23448 (N_23448,N_22430,N_22407);
and U23449 (N_23449,N_22345,N_22769);
nor U23450 (N_23450,N_22745,N_22599);
nor U23451 (N_23451,N_22902,N_22354);
or U23452 (N_23452,N_22453,N_22063);
and U23453 (N_23453,N_22840,N_22897);
nor U23454 (N_23454,N_22436,N_22899);
nand U23455 (N_23455,N_22934,N_22337);
nand U23456 (N_23456,N_22505,N_22779);
nor U23457 (N_23457,N_22586,N_22502);
nand U23458 (N_23458,N_22689,N_22508);
xor U23459 (N_23459,N_22037,N_22861);
xnor U23460 (N_23460,N_22803,N_22743);
and U23461 (N_23461,N_22722,N_22939);
xor U23462 (N_23462,N_22147,N_22698);
nor U23463 (N_23463,N_22640,N_22880);
and U23464 (N_23464,N_22117,N_22538);
or U23465 (N_23465,N_22002,N_22890);
xnor U23466 (N_23466,N_22220,N_22562);
nor U23467 (N_23467,N_22055,N_22052);
nor U23468 (N_23468,N_22308,N_22044);
nand U23469 (N_23469,N_22802,N_22556);
or U23470 (N_23470,N_22230,N_22584);
nor U23471 (N_23471,N_22568,N_22372);
xnor U23472 (N_23472,N_22446,N_22116);
nor U23473 (N_23473,N_22253,N_22614);
xor U23474 (N_23474,N_22049,N_22588);
nor U23475 (N_23475,N_22417,N_22298);
nor U23476 (N_23476,N_22222,N_22570);
xor U23477 (N_23477,N_22946,N_22388);
and U23478 (N_23478,N_22503,N_22917);
xnor U23479 (N_23479,N_22627,N_22623);
nor U23480 (N_23480,N_22550,N_22458);
nand U23481 (N_23481,N_22595,N_22499);
nand U23482 (N_23482,N_22685,N_22023);
and U23483 (N_23483,N_22534,N_22196);
and U23484 (N_23484,N_22661,N_22973);
nand U23485 (N_23485,N_22079,N_22719);
and U23486 (N_23486,N_22612,N_22727);
xor U23487 (N_23487,N_22863,N_22066);
nor U23488 (N_23488,N_22120,N_22017);
and U23489 (N_23489,N_22539,N_22975);
nand U23490 (N_23490,N_22654,N_22500);
nor U23491 (N_23491,N_22601,N_22318);
nor U23492 (N_23492,N_22676,N_22936);
or U23493 (N_23493,N_22440,N_22834);
nand U23494 (N_23494,N_22278,N_22706);
nand U23495 (N_23495,N_22170,N_22344);
nand U23496 (N_23496,N_22692,N_22853);
nor U23497 (N_23497,N_22045,N_22338);
xnor U23498 (N_23498,N_22611,N_22295);
nand U23499 (N_23499,N_22284,N_22518);
xnor U23500 (N_23500,N_22662,N_22285);
and U23501 (N_23501,N_22897,N_22519);
nand U23502 (N_23502,N_22739,N_22142);
and U23503 (N_23503,N_22363,N_22298);
xnor U23504 (N_23504,N_22956,N_22863);
and U23505 (N_23505,N_22516,N_22867);
nand U23506 (N_23506,N_22266,N_22207);
and U23507 (N_23507,N_22349,N_22780);
and U23508 (N_23508,N_22679,N_22643);
nand U23509 (N_23509,N_22142,N_22570);
xnor U23510 (N_23510,N_22872,N_22878);
nor U23511 (N_23511,N_22051,N_22530);
nor U23512 (N_23512,N_22326,N_22629);
nand U23513 (N_23513,N_22189,N_22877);
or U23514 (N_23514,N_22833,N_22656);
nor U23515 (N_23515,N_22461,N_22791);
or U23516 (N_23516,N_22259,N_22511);
nor U23517 (N_23517,N_22669,N_22913);
and U23518 (N_23518,N_22088,N_22798);
or U23519 (N_23519,N_22905,N_22765);
and U23520 (N_23520,N_22567,N_22692);
nand U23521 (N_23521,N_22117,N_22600);
nand U23522 (N_23522,N_22719,N_22279);
and U23523 (N_23523,N_22584,N_22259);
and U23524 (N_23524,N_22717,N_22970);
nor U23525 (N_23525,N_22397,N_22420);
and U23526 (N_23526,N_22133,N_22945);
and U23527 (N_23527,N_22783,N_22946);
and U23528 (N_23528,N_22126,N_22342);
xnor U23529 (N_23529,N_22307,N_22512);
xor U23530 (N_23530,N_22678,N_22490);
nor U23531 (N_23531,N_22970,N_22671);
xnor U23532 (N_23532,N_22659,N_22295);
xnor U23533 (N_23533,N_22946,N_22564);
xor U23534 (N_23534,N_22050,N_22310);
xnor U23535 (N_23535,N_22507,N_22069);
or U23536 (N_23536,N_22981,N_22047);
and U23537 (N_23537,N_22324,N_22736);
or U23538 (N_23538,N_22077,N_22024);
nor U23539 (N_23539,N_22733,N_22456);
nand U23540 (N_23540,N_22172,N_22515);
and U23541 (N_23541,N_22098,N_22201);
xor U23542 (N_23542,N_22240,N_22901);
nor U23543 (N_23543,N_22889,N_22368);
xnor U23544 (N_23544,N_22687,N_22849);
nor U23545 (N_23545,N_22971,N_22305);
and U23546 (N_23546,N_22732,N_22430);
nand U23547 (N_23547,N_22172,N_22110);
xnor U23548 (N_23548,N_22760,N_22772);
and U23549 (N_23549,N_22637,N_22839);
nor U23550 (N_23550,N_22916,N_22755);
xor U23551 (N_23551,N_22484,N_22527);
or U23552 (N_23552,N_22879,N_22498);
or U23553 (N_23553,N_22108,N_22917);
or U23554 (N_23554,N_22422,N_22347);
nor U23555 (N_23555,N_22414,N_22065);
nand U23556 (N_23556,N_22962,N_22788);
nor U23557 (N_23557,N_22692,N_22073);
or U23558 (N_23558,N_22583,N_22224);
nand U23559 (N_23559,N_22779,N_22806);
and U23560 (N_23560,N_22548,N_22662);
or U23561 (N_23561,N_22269,N_22205);
or U23562 (N_23562,N_22846,N_22169);
and U23563 (N_23563,N_22350,N_22710);
nor U23564 (N_23564,N_22481,N_22405);
nor U23565 (N_23565,N_22660,N_22501);
nand U23566 (N_23566,N_22407,N_22117);
xnor U23567 (N_23567,N_22734,N_22606);
nand U23568 (N_23568,N_22527,N_22865);
nand U23569 (N_23569,N_22408,N_22539);
and U23570 (N_23570,N_22396,N_22722);
nand U23571 (N_23571,N_22825,N_22045);
nor U23572 (N_23572,N_22395,N_22806);
nand U23573 (N_23573,N_22182,N_22600);
nand U23574 (N_23574,N_22228,N_22626);
nor U23575 (N_23575,N_22881,N_22995);
nand U23576 (N_23576,N_22086,N_22046);
nor U23577 (N_23577,N_22660,N_22537);
nor U23578 (N_23578,N_22719,N_22493);
and U23579 (N_23579,N_22321,N_22393);
or U23580 (N_23580,N_22279,N_22539);
nor U23581 (N_23581,N_22908,N_22181);
nor U23582 (N_23582,N_22801,N_22658);
and U23583 (N_23583,N_22811,N_22345);
or U23584 (N_23584,N_22662,N_22619);
nand U23585 (N_23585,N_22650,N_22008);
nand U23586 (N_23586,N_22733,N_22088);
and U23587 (N_23587,N_22606,N_22311);
and U23588 (N_23588,N_22230,N_22213);
or U23589 (N_23589,N_22117,N_22071);
nand U23590 (N_23590,N_22770,N_22001);
or U23591 (N_23591,N_22451,N_22634);
xor U23592 (N_23592,N_22010,N_22392);
and U23593 (N_23593,N_22700,N_22873);
xnor U23594 (N_23594,N_22662,N_22256);
and U23595 (N_23595,N_22276,N_22643);
or U23596 (N_23596,N_22365,N_22268);
and U23597 (N_23597,N_22195,N_22151);
or U23598 (N_23598,N_22729,N_22691);
nor U23599 (N_23599,N_22115,N_22334);
and U23600 (N_23600,N_22103,N_22724);
nand U23601 (N_23601,N_22172,N_22020);
nand U23602 (N_23602,N_22460,N_22320);
and U23603 (N_23603,N_22400,N_22315);
and U23604 (N_23604,N_22322,N_22420);
nor U23605 (N_23605,N_22476,N_22798);
nand U23606 (N_23606,N_22257,N_22182);
and U23607 (N_23607,N_22288,N_22197);
nor U23608 (N_23608,N_22527,N_22026);
xor U23609 (N_23609,N_22175,N_22296);
xor U23610 (N_23610,N_22370,N_22086);
nor U23611 (N_23611,N_22051,N_22934);
nand U23612 (N_23612,N_22379,N_22460);
nor U23613 (N_23613,N_22256,N_22653);
nor U23614 (N_23614,N_22341,N_22187);
nand U23615 (N_23615,N_22391,N_22197);
nor U23616 (N_23616,N_22092,N_22540);
xnor U23617 (N_23617,N_22868,N_22905);
or U23618 (N_23618,N_22389,N_22983);
xnor U23619 (N_23619,N_22689,N_22470);
or U23620 (N_23620,N_22396,N_22091);
and U23621 (N_23621,N_22044,N_22615);
and U23622 (N_23622,N_22690,N_22141);
nor U23623 (N_23623,N_22718,N_22871);
nand U23624 (N_23624,N_22913,N_22310);
or U23625 (N_23625,N_22463,N_22042);
and U23626 (N_23626,N_22342,N_22789);
xnor U23627 (N_23627,N_22421,N_22089);
or U23628 (N_23628,N_22977,N_22063);
or U23629 (N_23629,N_22706,N_22334);
and U23630 (N_23630,N_22863,N_22406);
or U23631 (N_23631,N_22233,N_22131);
nor U23632 (N_23632,N_22488,N_22320);
nor U23633 (N_23633,N_22323,N_22720);
and U23634 (N_23634,N_22579,N_22498);
and U23635 (N_23635,N_22660,N_22980);
nand U23636 (N_23636,N_22418,N_22318);
or U23637 (N_23637,N_22769,N_22379);
or U23638 (N_23638,N_22412,N_22234);
or U23639 (N_23639,N_22669,N_22726);
nor U23640 (N_23640,N_22296,N_22260);
or U23641 (N_23641,N_22917,N_22128);
and U23642 (N_23642,N_22330,N_22378);
xor U23643 (N_23643,N_22028,N_22405);
or U23644 (N_23644,N_22114,N_22322);
and U23645 (N_23645,N_22796,N_22317);
nor U23646 (N_23646,N_22532,N_22446);
nand U23647 (N_23647,N_22210,N_22288);
and U23648 (N_23648,N_22769,N_22533);
nand U23649 (N_23649,N_22264,N_22641);
and U23650 (N_23650,N_22362,N_22790);
or U23651 (N_23651,N_22449,N_22703);
nand U23652 (N_23652,N_22856,N_22120);
and U23653 (N_23653,N_22739,N_22547);
xnor U23654 (N_23654,N_22894,N_22695);
or U23655 (N_23655,N_22495,N_22221);
or U23656 (N_23656,N_22649,N_22170);
or U23657 (N_23657,N_22543,N_22200);
xor U23658 (N_23658,N_22091,N_22732);
nor U23659 (N_23659,N_22187,N_22709);
xor U23660 (N_23660,N_22641,N_22945);
nand U23661 (N_23661,N_22772,N_22161);
nand U23662 (N_23662,N_22810,N_22499);
nand U23663 (N_23663,N_22502,N_22211);
or U23664 (N_23664,N_22098,N_22037);
and U23665 (N_23665,N_22535,N_22704);
xnor U23666 (N_23666,N_22857,N_22630);
and U23667 (N_23667,N_22823,N_22564);
xor U23668 (N_23668,N_22498,N_22857);
and U23669 (N_23669,N_22078,N_22343);
and U23670 (N_23670,N_22387,N_22392);
xor U23671 (N_23671,N_22956,N_22724);
or U23672 (N_23672,N_22748,N_22293);
xnor U23673 (N_23673,N_22870,N_22079);
nor U23674 (N_23674,N_22573,N_22630);
xor U23675 (N_23675,N_22928,N_22550);
and U23676 (N_23676,N_22065,N_22433);
xnor U23677 (N_23677,N_22992,N_22371);
xnor U23678 (N_23678,N_22341,N_22122);
or U23679 (N_23679,N_22889,N_22535);
nor U23680 (N_23680,N_22305,N_22742);
nor U23681 (N_23681,N_22994,N_22706);
nor U23682 (N_23682,N_22266,N_22992);
or U23683 (N_23683,N_22753,N_22429);
or U23684 (N_23684,N_22520,N_22395);
nand U23685 (N_23685,N_22082,N_22525);
nand U23686 (N_23686,N_22806,N_22899);
nand U23687 (N_23687,N_22075,N_22710);
xor U23688 (N_23688,N_22583,N_22174);
xor U23689 (N_23689,N_22132,N_22180);
and U23690 (N_23690,N_22533,N_22151);
nand U23691 (N_23691,N_22010,N_22170);
or U23692 (N_23692,N_22135,N_22254);
nor U23693 (N_23693,N_22616,N_22401);
and U23694 (N_23694,N_22670,N_22354);
xnor U23695 (N_23695,N_22354,N_22930);
and U23696 (N_23696,N_22550,N_22851);
xor U23697 (N_23697,N_22787,N_22036);
and U23698 (N_23698,N_22244,N_22574);
nand U23699 (N_23699,N_22803,N_22028);
nand U23700 (N_23700,N_22600,N_22341);
xor U23701 (N_23701,N_22206,N_22656);
and U23702 (N_23702,N_22541,N_22440);
xor U23703 (N_23703,N_22194,N_22498);
or U23704 (N_23704,N_22870,N_22148);
nand U23705 (N_23705,N_22466,N_22580);
nor U23706 (N_23706,N_22670,N_22858);
or U23707 (N_23707,N_22028,N_22875);
and U23708 (N_23708,N_22406,N_22265);
xnor U23709 (N_23709,N_22267,N_22572);
or U23710 (N_23710,N_22209,N_22147);
xor U23711 (N_23711,N_22163,N_22873);
nor U23712 (N_23712,N_22780,N_22261);
nor U23713 (N_23713,N_22939,N_22241);
nor U23714 (N_23714,N_22601,N_22252);
nand U23715 (N_23715,N_22057,N_22263);
and U23716 (N_23716,N_22168,N_22377);
nor U23717 (N_23717,N_22540,N_22215);
nand U23718 (N_23718,N_22816,N_22377);
or U23719 (N_23719,N_22291,N_22472);
nor U23720 (N_23720,N_22531,N_22254);
and U23721 (N_23721,N_22608,N_22492);
and U23722 (N_23722,N_22478,N_22305);
xnor U23723 (N_23723,N_22255,N_22242);
or U23724 (N_23724,N_22024,N_22651);
or U23725 (N_23725,N_22319,N_22388);
and U23726 (N_23726,N_22779,N_22204);
or U23727 (N_23727,N_22194,N_22744);
xor U23728 (N_23728,N_22064,N_22921);
or U23729 (N_23729,N_22384,N_22590);
nand U23730 (N_23730,N_22885,N_22318);
nand U23731 (N_23731,N_22376,N_22772);
nor U23732 (N_23732,N_22963,N_22617);
nand U23733 (N_23733,N_22793,N_22146);
or U23734 (N_23734,N_22363,N_22230);
xnor U23735 (N_23735,N_22115,N_22491);
nor U23736 (N_23736,N_22587,N_22879);
nand U23737 (N_23737,N_22797,N_22642);
and U23738 (N_23738,N_22490,N_22324);
xor U23739 (N_23739,N_22605,N_22776);
nor U23740 (N_23740,N_22804,N_22993);
nand U23741 (N_23741,N_22428,N_22467);
nor U23742 (N_23742,N_22105,N_22120);
nand U23743 (N_23743,N_22190,N_22523);
nand U23744 (N_23744,N_22302,N_22809);
and U23745 (N_23745,N_22603,N_22600);
nor U23746 (N_23746,N_22967,N_22856);
or U23747 (N_23747,N_22700,N_22389);
or U23748 (N_23748,N_22006,N_22210);
nand U23749 (N_23749,N_22307,N_22833);
or U23750 (N_23750,N_22108,N_22009);
nor U23751 (N_23751,N_22692,N_22079);
nor U23752 (N_23752,N_22834,N_22387);
xnor U23753 (N_23753,N_22698,N_22690);
xor U23754 (N_23754,N_22625,N_22949);
nand U23755 (N_23755,N_22588,N_22148);
nor U23756 (N_23756,N_22975,N_22477);
and U23757 (N_23757,N_22364,N_22555);
nand U23758 (N_23758,N_22365,N_22544);
nand U23759 (N_23759,N_22284,N_22477);
xnor U23760 (N_23760,N_22937,N_22196);
and U23761 (N_23761,N_22265,N_22928);
xor U23762 (N_23762,N_22042,N_22962);
nand U23763 (N_23763,N_22014,N_22493);
and U23764 (N_23764,N_22457,N_22604);
nand U23765 (N_23765,N_22132,N_22733);
nor U23766 (N_23766,N_22254,N_22868);
and U23767 (N_23767,N_22197,N_22999);
nand U23768 (N_23768,N_22167,N_22702);
nand U23769 (N_23769,N_22344,N_22857);
nor U23770 (N_23770,N_22309,N_22840);
or U23771 (N_23771,N_22334,N_22928);
and U23772 (N_23772,N_22006,N_22911);
nor U23773 (N_23773,N_22548,N_22744);
nor U23774 (N_23774,N_22293,N_22869);
xor U23775 (N_23775,N_22472,N_22817);
or U23776 (N_23776,N_22329,N_22595);
nand U23777 (N_23777,N_22909,N_22093);
and U23778 (N_23778,N_22638,N_22231);
or U23779 (N_23779,N_22097,N_22263);
nand U23780 (N_23780,N_22924,N_22540);
nand U23781 (N_23781,N_22688,N_22961);
nand U23782 (N_23782,N_22916,N_22836);
nor U23783 (N_23783,N_22308,N_22796);
or U23784 (N_23784,N_22341,N_22661);
nor U23785 (N_23785,N_22582,N_22002);
nor U23786 (N_23786,N_22458,N_22107);
and U23787 (N_23787,N_22154,N_22891);
or U23788 (N_23788,N_22557,N_22832);
and U23789 (N_23789,N_22310,N_22273);
xnor U23790 (N_23790,N_22107,N_22193);
or U23791 (N_23791,N_22590,N_22884);
and U23792 (N_23792,N_22333,N_22413);
nor U23793 (N_23793,N_22073,N_22745);
nor U23794 (N_23794,N_22915,N_22220);
and U23795 (N_23795,N_22158,N_22925);
nand U23796 (N_23796,N_22896,N_22865);
nand U23797 (N_23797,N_22259,N_22364);
nand U23798 (N_23798,N_22667,N_22231);
xnor U23799 (N_23799,N_22542,N_22783);
or U23800 (N_23800,N_22407,N_22418);
nand U23801 (N_23801,N_22781,N_22650);
or U23802 (N_23802,N_22365,N_22163);
and U23803 (N_23803,N_22290,N_22482);
nor U23804 (N_23804,N_22909,N_22284);
nand U23805 (N_23805,N_22745,N_22854);
or U23806 (N_23806,N_22012,N_22558);
or U23807 (N_23807,N_22365,N_22387);
nor U23808 (N_23808,N_22536,N_22183);
nand U23809 (N_23809,N_22936,N_22129);
xor U23810 (N_23810,N_22047,N_22757);
xor U23811 (N_23811,N_22097,N_22277);
nor U23812 (N_23812,N_22858,N_22527);
xnor U23813 (N_23813,N_22663,N_22728);
nor U23814 (N_23814,N_22443,N_22328);
and U23815 (N_23815,N_22506,N_22710);
xnor U23816 (N_23816,N_22899,N_22189);
or U23817 (N_23817,N_22063,N_22253);
nand U23818 (N_23818,N_22802,N_22442);
xor U23819 (N_23819,N_22404,N_22147);
nand U23820 (N_23820,N_22021,N_22969);
xor U23821 (N_23821,N_22211,N_22303);
xnor U23822 (N_23822,N_22103,N_22566);
and U23823 (N_23823,N_22756,N_22666);
and U23824 (N_23824,N_22671,N_22271);
nor U23825 (N_23825,N_22417,N_22333);
nor U23826 (N_23826,N_22589,N_22104);
nor U23827 (N_23827,N_22472,N_22367);
and U23828 (N_23828,N_22224,N_22848);
xnor U23829 (N_23829,N_22136,N_22021);
or U23830 (N_23830,N_22963,N_22361);
nand U23831 (N_23831,N_22273,N_22922);
nor U23832 (N_23832,N_22654,N_22275);
xor U23833 (N_23833,N_22890,N_22460);
and U23834 (N_23834,N_22851,N_22037);
nor U23835 (N_23835,N_22120,N_22414);
and U23836 (N_23836,N_22920,N_22199);
xnor U23837 (N_23837,N_22378,N_22885);
xor U23838 (N_23838,N_22311,N_22380);
nand U23839 (N_23839,N_22545,N_22682);
xnor U23840 (N_23840,N_22209,N_22658);
nor U23841 (N_23841,N_22504,N_22223);
nand U23842 (N_23842,N_22378,N_22823);
and U23843 (N_23843,N_22151,N_22723);
nand U23844 (N_23844,N_22567,N_22490);
or U23845 (N_23845,N_22324,N_22352);
nor U23846 (N_23846,N_22868,N_22072);
or U23847 (N_23847,N_22359,N_22847);
nor U23848 (N_23848,N_22723,N_22853);
nor U23849 (N_23849,N_22486,N_22406);
or U23850 (N_23850,N_22660,N_22762);
xor U23851 (N_23851,N_22333,N_22896);
xnor U23852 (N_23852,N_22986,N_22425);
nand U23853 (N_23853,N_22434,N_22975);
xor U23854 (N_23854,N_22956,N_22691);
nand U23855 (N_23855,N_22286,N_22752);
and U23856 (N_23856,N_22155,N_22267);
nor U23857 (N_23857,N_22054,N_22213);
xor U23858 (N_23858,N_22564,N_22460);
nor U23859 (N_23859,N_22650,N_22625);
xor U23860 (N_23860,N_22527,N_22749);
or U23861 (N_23861,N_22561,N_22448);
nor U23862 (N_23862,N_22859,N_22019);
and U23863 (N_23863,N_22343,N_22692);
and U23864 (N_23864,N_22597,N_22517);
or U23865 (N_23865,N_22310,N_22103);
and U23866 (N_23866,N_22657,N_22406);
xor U23867 (N_23867,N_22453,N_22849);
nand U23868 (N_23868,N_22440,N_22349);
and U23869 (N_23869,N_22145,N_22749);
nand U23870 (N_23870,N_22109,N_22284);
nand U23871 (N_23871,N_22521,N_22632);
and U23872 (N_23872,N_22151,N_22309);
and U23873 (N_23873,N_22334,N_22078);
nand U23874 (N_23874,N_22723,N_22053);
nor U23875 (N_23875,N_22335,N_22690);
nor U23876 (N_23876,N_22291,N_22059);
nor U23877 (N_23877,N_22817,N_22126);
nor U23878 (N_23878,N_22192,N_22225);
and U23879 (N_23879,N_22739,N_22676);
nand U23880 (N_23880,N_22809,N_22251);
nand U23881 (N_23881,N_22882,N_22177);
nand U23882 (N_23882,N_22402,N_22054);
nor U23883 (N_23883,N_22842,N_22655);
and U23884 (N_23884,N_22731,N_22055);
and U23885 (N_23885,N_22924,N_22301);
xnor U23886 (N_23886,N_22666,N_22534);
or U23887 (N_23887,N_22452,N_22748);
or U23888 (N_23888,N_22253,N_22468);
nand U23889 (N_23889,N_22784,N_22561);
and U23890 (N_23890,N_22112,N_22327);
or U23891 (N_23891,N_22848,N_22096);
or U23892 (N_23892,N_22785,N_22618);
nand U23893 (N_23893,N_22906,N_22305);
nand U23894 (N_23894,N_22820,N_22683);
and U23895 (N_23895,N_22457,N_22514);
xnor U23896 (N_23896,N_22373,N_22118);
xor U23897 (N_23897,N_22429,N_22284);
xor U23898 (N_23898,N_22016,N_22711);
nand U23899 (N_23899,N_22038,N_22794);
and U23900 (N_23900,N_22617,N_22389);
nand U23901 (N_23901,N_22048,N_22888);
xnor U23902 (N_23902,N_22091,N_22251);
or U23903 (N_23903,N_22315,N_22696);
or U23904 (N_23904,N_22496,N_22522);
xor U23905 (N_23905,N_22189,N_22738);
and U23906 (N_23906,N_22405,N_22416);
and U23907 (N_23907,N_22311,N_22678);
xor U23908 (N_23908,N_22887,N_22398);
or U23909 (N_23909,N_22503,N_22863);
and U23910 (N_23910,N_22719,N_22847);
and U23911 (N_23911,N_22816,N_22805);
nor U23912 (N_23912,N_22575,N_22061);
xnor U23913 (N_23913,N_22565,N_22307);
nand U23914 (N_23914,N_22202,N_22927);
and U23915 (N_23915,N_22226,N_22164);
nor U23916 (N_23916,N_22328,N_22638);
nor U23917 (N_23917,N_22755,N_22651);
and U23918 (N_23918,N_22291,N_22657);
and U23919 (N_23919,N_22090,N_22583);
nor U23920 (N_23920,N_22471,N_22503);
xnor U23921 (N_23921,N_22846,N_22441);
xnor U23922 (N_23922,N_22717,N_22949);
and U23923 (N_23923,N_22421,N_22386);
nand U23924 (N_23924,N_22659,N_22655);
and U23925 (N_23925,N_22540,N_22346);
xnor U23926 (N_23926,N_22655,N_22251);
nor U23927 (N_23927,N_22022,N_22409);
or U23928 (N_23928,N_22349,N_22668);
or U23929 (N_23929,N_22535,N_22558);
nand U23930 (N_23930,N_22787,N_22408);
nand U23931 (N_23931,N_22465,N_22460);
nor U23932 (N_23932,N_22698,N_22977);
nand U23933 (N_23933,N_22634,N_22392);
or U23934 (N_23934,N_22697,N_22294);
xor U23935 (N_23935,N_22593,N_22033);
or U23936 (N_23936,N_22890,N_22932);
xnor U23937 (N_23937,N_22747,N_22439);
xnor U23938 (N_23938,N_22293,N_22541);
xor U23939 (N_23939,N_22647,N_22893);
or U23940 (N_23940,N_22238,N_22685);
and U23941 (N_23941,N_22793,N_22720);
xnor U23942 (N_23942,N_22165,N_22207);
and U23943 (N_23943,N_22699,N_22739);
or U23944 (N_23944,N_22504,N_22208);
nor U23945 (N_23945,N_22381,N_22821);
nand U23946 (N_23946,N_22726,N_22079);
nand U23947 (N_23947,N_22708,N_22279);
or U23948 (N_23948,N_22815,N_22612);
nor U23949 (N_23949,N_22907,N_22460);
or U23950 (N_23950,N_22009,N_22538);
and U23951 (N_23951,N_22740,N_22690);
nand U23952 (N_23952,N_22487,N_22315);
nor U23953 (N_23953,N_22958,N_22400);
xnor U23954 (N_23954,N_22135,N_22456);
nand U23955 (N_23955,N_22876,N_22471);
nor U23956 (N_23956,N_22849,N_22771);
nand U23957 (N_23957,N_22441,N_22381);
nor U23958 (N_23958,N_22783,N_22484);
nand U23959 (N_23959,N_22163,N_22564);
xor U23960 (N_23960,N_22621,N_22448);
nand U23961 (N_23961,N_22666,N_22920);
nand U23962 (N_23962,N_22524,N_22908);
nand U23963 (N_23963,N_22312,N_22307);
nand U23964 (N_23964,N_22550,N_22932);
nand U23965 (N_23965,N_22429,N_22305);
and U23966 (N_23966,N_22346,N_22148);
nand U23967 (N_23967,N_22326,N_22631);
xnor U23968 (N_23968,N_22978,N_22360);
and U23969 (N_23969,N_22833,N_22996);
xor U23970 (N_23970,N_22329,N_22864);
nand U23971 (N_23971,N_22727,N_22154);
nor U23972 (N_23972,N_22226,N_22624);
xor U23973 (N_23973,N_22093,N_22533);
or U23974 (N_23974,N_22519,N_22256);
or U23975 (N_23975,N_22553,N_22061);
or U23976 (N_23976,N_22232,N_22904);
nor U23977 (N_23977,N_22350,N_22838);
and U23978 (N_23978,N_22710,N_22089);
xor U23979 (N_23979,N_22438,N_22053);
nand U23980 (N_23980,N_22595,N_22086);
nor U23981 (N_23981,N_22343,N_22094);
or U23982 (N_23982,N_22647,N_22324);
xnor U23983 (N_23983,N_22881,N_22398);
nor U23984 (N_23984,N_22837,N_22610);
and U23985 (N_23985,N_22418,N_22955);
nand U23986 (N_23986,N_22487,N_22138);
xor U23987 (N_23987,N_22656,N_22939);
nor U23988 (N_23988,N_22220,N_22206);
nand U23989 (N_23989,N_22701,N_22070);
and U23990 (N_23990,N_22870,N_22018);
nand U23991 (N_23991,N_22513,N_22686);
and U23992 (N_23992,N_22076,N_22218);
nor U23993 (N_23993,N_22461,N_22581);
and U23994 (N_23994,N_22167,N_22940);
or U23995 (N_23995,N_22258,N_22886);
xor U23996 (N_23996,N_22711,N_22029);
xor U23997 (N_23997,N_22000,N_22524);
nor U23998 (N_23998,N_22908,N_22748);
xnor U23999 (N_23999,N_22778,N_22919);
nor U24000 (N_24000,N_23236,N_23212);
xor U24001 (N_24001,N_23149,N_23086);
and U24002 (N_24002,N_23623,N_23608);
nand U24003 (N_24003,N_23641,N_23787);
nor U24004 (N_24004,N_23851,N_23252);
nand U24005 (N_24005,N_23545,N_23433);
xnor U24006 (N_24006,N_23559,N_23001);
and U24007 (N_24007,N_23510,N_23846);
or U24008 (N_24008,N_23144,N_23082);
and U24009 (N_24009,N_23333,N_23084);
nor U24010 (N_24010,N_23651,N_23513);
and U24011 (N_24011,N_23339,N_23043);
nor U24012 (N_24012,N_23294,N_23492);
or U24013 (N_24013,N_23221,N_23135);
or U24014 (N_24014,N_23749,N_23183);
nand U24015 (N_24015,N_23985,N_23818);
or U24016 (N_24016,N_23401,N_23382);
nor U24017 (N_24017,N_23399,N_23165);
or U24018 (N_24018,N_23599,N_23400);
xnor U24019 (N_24019,N_23189,N_23437);
and U24020 (N_24020,N_23041,N_23298);
nand U24021 (N_24021,N_23882,N_23344);
xor U24022 (N_24022,N_23918,N_23206);
xnor U24023 (N_24023,N_23705,N_23520);
and U24024 (N_24024,N_23604,N_23529);
and U24025 (N_24025,N_23963,N_23774);
nand U24026 (N_24026,N_23569,N_23708);
nand U24027 (N_24027,N_23442,N_23314);
xnor U24028 (N_24028,N_23118,N_23104);
or U24029 (N_24029,N_23226,N_23715);
xor U24030 (N_24030,N_23178,N_23993);
or U24031 (N_24031,N_23887,N_23813);
and U24032 (N_24032,N_23665,N_23776);
nand U24033 (N_24033,N_23688,N_23472);
nand U24034 (N_24034,N_23573,N_23577);
nand U24035 (N_24035,N_23463,N_23826);
nor U24036 (N_24036,N_23151,N_23042);
nor U24037 (N_24037,N_23969,N_23272);
nand U24038 (N_24038,N_23976,N_23578);
nor U24039 (N_24039,N_23532,N_23975);
and U24040 (N_24040,N_23311,N_23678);
nor U24041 (N_24041,N_23110,N_23026);
nand U24042 (N_24042,N_23420,N_23836);
xor U24043 (N_24043,N_23295,N_23340);
xor U24044 (N_24044,N_23824,N_23536);
nand U24045 (N_24045,N_23989,N_23910);
or U24046 (N_24046,N_23177,N_23711);
nand U24047 (N_24047,N_23156,N_23871);
or U24048 (N_24048,N_23157,N_23704);
xor U24049 (N_24049,N_23893,N_23241);
or U24050 (N_24050,N_23673,N_23005);
and U24051 (N_24051,N_23480,N_23025);
nand U24052 (N_24052,N_23927,N_23058);
nand U24053 (N_24053,N_23231,N_23497);
xor U24054 (N_24054,N_23315,N_23753);
or U24055 (N_24055,N_23974,N_23820);
xnor U24056 (N_24056,N_23039,N_23342);
or U24057 (N_24057,N_23421,N_23065);
or U24058 (N_24058,N_23655,N_23676);
xor U24059 (N_24059,N_23318,N_23773);
xnor U24060 (N_24060,N_23331,N_23316);
and U24061 (N_24061,N_23588,N_23972);
nor U24062 (N_24062,N_23343,N_23732);
nand U24063 (N_24063,N_23816,N_23292);
nand U24064 (N_24064,N_23683,N_23855);
and U24065 (N_24065,N_23092,N_23111);
or U24066 (N_24066,N_23878,N_23435);
xnor U24067 (N_24067,N_23658,N_23371);
nor U24068 (N_24068,N_23973,N_23570);
and U24069 (N_24069,N_23150,N_23992);
xor U24070 (N_24070,N_23438,N_23654);
xnor U24071 (N_24071,N_23263,N_23763);
xnor U24072 (N_24072,N_23970,N_23209);
xnor U24073 (N_24073,N_23689,N_23502);
and U24074 (N_24074,N_23495,N_23391);
xnor U24075 (N_24075,N_23684,N_23585);
and U24076 (N_24076,N_23727,N_23982);
and U24077 (N_24077,N_23482,N_23134);
or U24078 (N_24078,N_23304,N_23978);
and U24079 (N_24079,N_23266,N_23739);
nor U24080 (N_24080,N_23936,N_23791);
nand U24081 (N_24081,N_23751,N_23872);
xor U24082 (N_24082,N_23103,N_23056);
nor U24083 (N_24083,N_23358,N_23411);
and U24084 (N_24084,N_23247,N_23580);
nand U24085 (N_24085,N_23067,N_23842);
nand U24086 (N_24086,N_23594,N_23809);
nand U24087 (N_24087,N_23153,N_23913);
xor U24088 (N_24088,N_23938,N_23552);
nor U24089 (N_24089,N_23377,N_23116);
or U24090 (N_24090,N_23019,N_23176);
xnor U24091 (N_24091,N_23376,N_23747);
nand U24092 (N_24092,N_23759,N_23385);
nand U24093 (N_24093,N_23995,N_23243);
and U24094 (N_24094,N_23922,N_23018);
nand U24095 (N_24095,N_23741,N_23662);
or U24096 (N_24096,N_23831,N_23860);
or U24097 (N_24097,N_23550,N_23907);
xor U24098 (N_24098,N_23138,N_23720);
xnor U24099 (N_24099,N_23379,N_23210);
nand U24100 (N_24100,N_23519,N_23187);
nor U24101 (N_24101,N_23485,N_23162);
nor U24102 (N_24102,N_23843,N_23249);
nand U24103 (N_24103,N_23583,N_23903);
or U24104 (N_24104,N_23657,N_23461);
nor U24105 (N_24105,N_23612,N_23561);
or U24106 (N_24106,N_23079,N_23228);
xor U24107 (N_24107,N_23489,N_23862);
xnor U24108 (N_24108,N_23046,N_23631);
nand U24109 (N_24109,N_23650,N_23511);
or U24110 (N_24110,N_23384,N_23539);
nor U24111 (N_24111,N_23548,N_23494);
xor U24112 (N_24112,N_23962,N_23737);
nand U24113 (N_24113,N_23870,N_23251);
and U24114 (N_24114,N_23370,N_23475);
nand U24115 (N_24115,N_23905,N_23589);
or U24116 (N_24116,N_23127,N_23591);
xor U24117 (N_24117,N_23464,N_23537);
xnor U24118 (N_24118,N_23235,N_23839);
and U24119 (N_24119,N_23327,N_23897);
nand U24120 (N_24120,N_23512,N_23131);
nand U24121 (N_24121,N_23467,N_23238);
nor U24122 (N_24122,N_23666,N_23285);
and U24123 (N_24123,N_23509,N_23447);
or U24124 (N_24124,N_23027,N_23731);
nor U24125 (N_24125,N_23788,N_23821);
xnor U24126 (N_24126,N_23011,N_23387);
nand U24127 (N_24127,N_23037,N_23514);
nor U24128 (N_24128,N_23160,N_23598);
or U24129 (N_24129,N_23572,N_23476);
xnor U24130 (N_24130,N_23540,N_23359);
nor U24131 (N_24131,N_23328,N_23671);
xor U24132 (N_24132,N_23863,N_23155);
nand U24133 (N_24133,N_23964,N_23953);
and U24134 (N_24134,N_23639,N_23644);
nor U24135 (N_24135,N_23255,N_23392);
nand U24136 (N_24136,N_23163,N_23636);
xor U24137 (N_24137,N_23909,N_23775);
or U24138 (N_24138,N_23603,N_23045);
and U24139 (N_24139,N_23770,N_23931);
and U24140 (N_24140,N_23023,N_23217);
nor U24141 (N_24141,N_23722,N_23047);
and U24142 (N_24142,N_23253,N_23083);
and U24143 (N_24143,N_23404,N_23817);
or U24144 (N_24144,N_23915,N_23606);
or U24145 (N_24145,N_23319,N_23718);
xnor U24146 (N_24146,N_23560,N_23614);
nand U24147 (N_24147,N_23772,N_23490);
nand U24148 (N_24148,N_23345,N_23670);
or U24149 (N_24149,N_23900,N_23367);
nand U24150 (N_24150,N_23771,N_23672);
nand U24151 (N_24151,N_23054,N_23088);
nand U24152 (N_24152,N_23547,N_23203);
nand U24153 (N_24153,N_23661,N_23431);
and U24154 (N_24154,N_23170,N_23659);
or U24155 (N_24155,N_23957,N_23616);
or U24156 (N_24156,N_23533,N_23745);
or U24157 (N_24157,N_23275,N_23432);
or U24158 (N_24158,N_23262,N_23060);
and U24159 (N_24159,N_23388,N_23694);
and U24160 (N_24160,N_23069,N_23748);
or U24161 (N_24161,N_23136,N_23997);
or U24162 (N_24162,N_23522,N_23287);
xnor U24163 (N_24163,N_23917,N_23814);
nor U24164 (N_24164,N_23626,N_23811);
nand U24165 (N_24165,N_23906,N_23615);
nand U24166 (N_24166,N_23725,N_23258);
nand U24167 (N_24167,N_23126,N_23699);
nor U24168 (N_24168,N_23436,N_23166);
nand U24169 (N_24169,N_23424,N_23764);
nand U24170 (N_24170,N_23955,N_23194);
nor U24171 (N_24171,N_23706,N_23434);
and U24172 (N_24172,N_23714,N_23777);
xor U24173 (N_24173,N_23305,N_23324);
xnor U24174 (N_24174,N_23954,N_23190);
nand U24175 (N_24175,N_23498,N_23015);
nand U24176 (N_24176,N_23460,N_23996);
and U24177 (N_24177,N_23124,N_23197);
xnor U24178 (N_24178,N_23668,N_23968);
or U24179 (N_24179,N_23602,N_23121);
nand U24180 (N_24180,N_23981,N_23419);
xnor U24181 (N_24181,N_23638,N_23402);
xnor U24182 (N_24182,N_23828,N_23161);
or U24183 (N_24183,N_23302,N_23680);
nand U24184 (N_24184,N_23686,N_23040);
nand U24185 (N_24185,N_23526,N_23857);
nor U24186 (N_24186,N_23240,N_23653);
or U24187 (N_24187,N_23102,N_23944);
nor U24188 (N_24188,N_23980,N_23754);
nand U24189 (N_24189,N_23418,N_23806);
nand U24190 (N_24190,N_23428,N_23850);
xor U24191 (N_24191,N_23852,N_23214);
xnor U24192 (N_24192,N_23899,N_23201);
and U24193 (N_24193,N_23458,N_23406);
nand U24194 (N_24194,N_23336,N_23279);
nand U24195 (N_24195,N_23825,N_23876);
or U24196 (N_24196,N_23596,N_23613);
xor U24197 (N_24197,N_23493,N_23234);
nand U24198 (N_24198,N_23713,N_23457);
and U24199 (N_24199,N_23325,N_23780);
and U24200 (N_24200,N_23035,N_23091);
or U24201 (N_24201,N_23914,N_23624);
or U24202 (N_24202,N_23488,N_23164);
xnor U24203 (N_24203,N_23628,N_23273);
or U24204 (N_24204,N_23115,N_23858);
or U24205 (N_24205,N_23622,N_23395);
or U24206 (N_24206,N_23077,N_23191);
nor U24207 (N_24207,N_23276,N_23140);
or U24208 (N_24208,N_23182,N_23592);
nor U24209 (N_24209,N_23994,N_23146);
and U24210 (N_24210,N_23679,N_23028);
and U24211 (N_24211,N_23620,N_23926);
or U24212 (N_24212,N_23733,N_23429);
xnor U24213 (N_24213,N_23089,N_23712);
or U24214 (N_24214,N_23904,N_23167);
and U24215 (N_24215,N_23139,N_23508);
nand U24216 (N_24216,N_23597,N_23426);
nand U24217 (N_24217,N_23632,N_23538);
nand U24218 (N_24218,N_23925,N_23875);
xnor U24219 (N_24219,N_23709,N_23427);
nand U24220 (N_24220,N_23723,N_23270);
xnor U24221 (N_24221,N_23990,N_23372);
or U24222 (N_24222,N_23335,N_23122);
xnor U24223 (N_24223,N_23491,N_23822);
nor U24224 (N_24224,N_23128,N_23987);
nand U24225 (N_24225,N_23055,N_23269);
xor U24226 (N_24226,N_23450,N_23901);
nor U24227 (N_24227,N_23849,N_23796);
and U24228 (N_24228,N_23365,N_23916);
xnor U24229 (N_24229,N_23541,N_23991);
xor U24230 (N_24230,N_23669,N_23074);
xnor U24231 (N_24231,N_23299,N_23087);
and U24232 (N_24232,N_23911,N_23179);
nand U24233 (N_24233,N_23109,N_23186);
nor U24234 (N_24234,N_23934,N_23652);
and U24235 (N_24235,N_23171,N_23282);
nor U24236 (N_24236,N_23677,N_23417);
and U24237 (N_24237,N_23719,N_23756);
nor U24238 (N_24238,N_23507,N_23700);
and U24239 (N_24239,N_23117,N_23451);
and U24240 (N_24240,N_23730,N_23629);
nand U24241 (N_24241,N_23667,N_23147);
and U24242 (N_24242,N_23920,N_23648);
nand U24243 (N_24243,N_23500,N_23114);
nor U24244 (N_24244,N_23172,N_23352);
nor U24245 (N_24245,N_23466,N_23867);
or U24246 (N_24246,N_23674,N_23080);
nor U24247 (N_24247,N_23891,N_23430);
xnor U24248 (N_24248,N_23357,N_23564);
nand U24249 (N_24249,N_23057,N_23169);
nand U24250 (N_24250,N_23568,N_23516);
or U24251 (N_24251,N_23070,N_23329);
and U24252 (N_24252,N_23072,N_23752);
and U24253 (N_24253,N_23396,N_23779);
xnor U24254 (N_24254,N_23601,N_23141);
xnor U24255 (N_24255,N_23798,N_23303);
xor U24256 (N_24256,N_23233,N_23259);
nor U24257 (N_24257,N_23322,N_23154);
nor U24258 (N_24258,N_23260,N_23643);
nor U24259 (N_24259,N_23479,N_23721);
xnor U24260 (N_24260,N_23152,N_23998);
xnor U24261 (N_24261,N_23635,N_23726);
xnor U24262 (N_24262,N_23459,N_23448);
xnor U24263 (N_24263,N_23609,N_23784);
or U24264 (N_24264,N_23293,N_23013);
or U24265 (N_24265,N_23803,N_23120);
xnor U24266 (N_24266,N_23364,N_23530);
or U24267 (N_24267,N_23192,N_23283);
xnor U24268 (N_24268,N_23830,N_23309);
nand U24269 (N_24269,N_23280,N_23943);
xnor U24270 (N_24270,N_23002,N_23804);
nand U24271 (N_24271,N_23697,N_23059);
or U24272 (N_24272,N_23765,N_23525);
nor U24273 (N_24273,N_23185,N_23363);
xor U24274 (N_24274,N_23886,N_23827);
nor U24275 (N_24275,N_23143,N_23261);
nor U24276 (N_24276,N_23563,N_23734);
or U24277 (N_24277,N_23782,N_23310);
and U24278 (N_24278,N_23068,N_23245);
and U24279 (N_24279,N_23647,N_23014);
nand U24280 (N_24280,N_23503,N_23605);
or U24281 (N_24281,N_23884,N_23554);
xnor U24282 (N_24282,N_23574,N_23009);
or U24283 (N_24283,N_23664,N_23724);
nor U24284 (N_24284,N_23693,N_23113);
nor U24285 (N_24285,N_23625,N_23085);
or U24286 (N_24286,N_23254,N_23902);
nand U24287 (N_24287,N_23349,N_23557);
xor U24288 (N_24288,N_23937,N_23394);
and U24289 (N_24289,N_23675,N_23355);
xnor U24290 (N_24290,N_23044,N_23810);
or U24291 (N_24291,N_23755,N_23361);
and U24292 (N_24292,N_23029,N_23956);
nand U24293 (N_24293,N_23337,N_23021);
nand U24294 (N_24294,N_23696,N_23119);
nand U24295 (N_24295,N_23312,N_23685);
nor U24296 (N_24296,N_23835,N_23761);
or U24297 (N_24297,N_23071,N_23617);
nand U24298 (N_24298,N_23880,N_23003);
nand U24299 (N_24299,N_23301,N_23341);
or U24300 (N_24300,N_23941,N_23052);
and U24301 (N_24301,N_23439,N_23215);
nor U24302 (N_24302,N_23208,N_23890);
nor U24303 (N_24303,N_23595,N_23308);
or U24304 (N_24304,N_23610,N_23838);
or U24305 (N_24305,N_23174,N_23033);
or U24306 (N_24306,N_23145,N_23440);
or U24307 (N_24307,N_23840,N_23453);
nand U24308 (N_24308,N_23945,N_23050);
nand U24309 (N_24309,N_23223,N_23017);
or U24310 (N_24310,N_23801,N_23845);
nand U24311 (N_24311,N_23237,N_23584);
and U24312 (N_24312,N_23297,N_23695);
or U24313 (N_24313,N_23123,N_23881);
or U24314 (N_24314,N_23107,N_23767);
and U24315 (N_24315,N_23137,N_23184);
nand U24316 (N_24316,N_23527,N_23004);
xnor U24317 (N_24317,N_23534,N_23959);
xnor U24318 (N_24318,N_23742,N_23330);
nor U24319 (N_24319,N_23378,N_23097);
nand U24320 (N_24320,N_23173,N_23812);
nand U24321 (N_24321,N_23888,N_23290);
nand U24322 (N_24322,N_23100,N_23274);
nand U24323 (N_24323,N_23196,N_23521);
or U24324 (N_24324,N_23542,N_23063);
and U24325 (N_24325,N_23108,N_23618);
nor U24326 (N_24326,N_23866,N_23856);
or U24327 (N_24327,N_23389,N_23928);
xnor U24328 (N_24328,N_23769,N_23353);
and U24329 (N_24329,N_23929,N_23222);
or U24330 (N_24330,N_23038,N_23244);
nor U24331 (N_24331,N_23408,N_23142);
nor U24332 (N_24332,N_23778,N_23032);
or U24333 (N_24333,N_23218,N_23646);
nand U24334 (N_24334,N_23278,N_23794);
nor U24335 (N_24335,N_23877,N_23762);
and U24336 (N_24336,N_23642,N_23474);
and U24337 (N_24337,N_23889,N_23868);
nand U24338 (N_24338,N_23351,N_23300);
nand U24339 (N_24339,N_23374,N_23819);
xor U24340 (N_24340,N_23571,N_23523);
or U24341 (N_24341,N_23861,N_23950);
and U24342 (N_24342,N_23094,N_23397);
nand U24343 (N_24343,N_23579,N_23805);
or U24344 (N_24344,N_23783,N_23455);
nor U24345 (N_24345,N_23932,N_23898);
nand U24346 (N_24346,N_23219,N_23250);
nor U24347 (N_24347,N_23885,N_23213);
nand U24348 (N_24348,N_23795,N_23199);
nor U24349 (N_24349,N_23239,N_23334);
nor U24350 (N_24350,N_23229,N_23180);
xnor U24351 (N_24351,N_23815,N_23487);
nor U24352 (N_24352,N_23832,N_23348);
and U24353 (N_24353,N_23366,N_23874);
xnor U24354 (N_24354,N_23637,N_23942);
xnor U24355 (N_24355,N_23469,N_23586);
or U24356 (N_24356,N_23125,N_23879);
and U24357 (N_24357,N_23531,N_23486);
nand U24358 (N_24358,N_23360,N_23535);
xnor U24359 (N_24359,N_23347,N_23656);
and U24360 (N_24360,N_23073,N_23307);
xnor U24361 (N_24361,N_23132,N_23248);
nand U24362 (N_24362,N_23416,N_23268);
nand U24363 (N_24363,N_23716,N_23061);
and U24364 (N_24364,N_23462,N_23565);
nand U24365 (N_24365,N_23634,N_23649);
nor U24366 (N_24366,N_23528,N_23148);
nor U24367 (N_24367,N_23543,N_23768);
and U24368 (N_24368,N_23744,N_23291);
nor U24369 (N_24369,N_23443,N_23296);
nor U24370 (N_24370,N_23940,N_23967);
nand U24371 (N_24371,N_23785,N_23332);
and U24372 (N_24372,N_23965,N_23284);
or U24373 (N_24373,N_23354,N_23211);
xnor U24374 (N_24374,N_23690,N_23468);
nor U24375 (N_24375,N_23338,N_23205);
nor U24376 (N_24376,N_23952,N_23277);
and U24377 (N_24377,N_23946,N_23381);
and U24378 (N_24378,N_23986,N_23947);
or U24379 (N_24379,N_23415,N_23735);
nor U24380 (N_24380,N_23048,N_23317);
xnor U24381 (N_24381,N_23386,N_23471);
or U24382 (N_24382,N_23707,N_23064);
nor U24383 (N_24383,N_23477,N_23930);
xnor U24384 (N_24384,N_23621,N_23869);
nor U24385 (N_24385,N_23627,N_23256);
or U24386 (N_24386,N_23556,N_23587);
or U24387 (N_24387,N_23757,N_23593);
nor U24388 (N_24388,N_23834,N_23101);
nor U24389 (N_24389,N_23020,N_23633);
and U24390 (N_24390,N_23912,N_23066);
nand U24391 (N_24391,N_23313,N_23413);
and U24392 (N_24392,N_23619,N_23326);
or U24393 (N_24393,N_23076,N_23949);
xnor U24394 (N_24394,N_23198,N_23766);
and U24395 (N_24395,N_23454,N_23112);
nand U24396 (N_24396,N_23224,N_23935);
and U24397 (N_24397,N_23346,N_23220);
or U24398 (N_24398,N_23390,N_23499);
or U24399 (N_24399,N_23130,N_23544);
and U24400 (N_24400,N_23008,N_23106);
or U24401 (N_24401,N_23242,N_23195);
and U24402 (N_24402,N_23750,N_23288);
nand U24403 (N_24403,N_23600,N_23425);
xor U24404 (N_24404,N_23012,N_23193);
and U24405 (N_24405,N_23159,N_23441);
and U24406 (N_24406,N_23181,N_23999);
or U24407 (N_24407,N_23793,N_23216);
nor U24408 (N_24408,N_23865,N_23681);
or U24409 (N_24409,N_23687,N_23034);
or U24410 (N_24410,N_23567,N_23409);
or U24411 (N_24411,N_23504,N_23465);
nor U24412 (N_24412,N_23422,N_23405);
and U24413 (N_24413,N_23743,N_23576);
or U24414 (N_24414,N_23702,N_23844);
nor U24415 (N_24415,N_23546,N_23575);
or U24416 (N_24416,N_23470,N_23383);
nor U24417 (N_24417,N_23175,N_23710);
nor U24418 (N_24418,N_23473,N_23051);
or U24419 (N_24419,N_23663,N_23264);
nand U24420 (N_24420,N_23188,N_23022);
xor U24421 (N_24421,N_23566,N_23892);
nand U24422 (N_24422,N_23007,N_23607);
nor U24423 (N_24423,N_23807,N_23802);
nor U24424 (N_24424,N_23698,N_23873);
xor U24425 (N_24425,N_23407,N_23081);
xnor U24426 (N_24426,N_23016,N_23983);
and U24427 (N_24427,N_23093,N_23919);
and U24428 (N_24428,N_23859,N_23078);
and U24429 (N_24429,N_23854,N_23496);
nor U24430 (N_24430,N_23823,N_23933);
xor U24431 (N_24431,N_23847,N_23611);
xnor U24432 (N_24432,N_23031,N_23728);
or U24433 (N_24433,N_23207,N_23505);
or U24434 (N_24434,N_23232,N_23864);
nor U24435 (N_24435,N_23966,N_23924);
xor U24436 (N_24436,N_23362,N_23090);
or U24437 (N_24437,N_23202,N_23740);
and U24438 (N_24438,N_23797,N_23271);
xor U24439 (N_24439,N_23000,N_23230);
xor U24440 (N_24440,N_23703,N_23691);
xor U24441 (N_24441,N_23129,N_23168);
and U24442 (N_24442,N_23036,N_23062);
nor U24443 (N_24443,N_23133,N_23977);
nand U24444 (N_24444,N_23948,N_23010);
or U24445 (N_24445,N_23030,N_23524);
xnor U24446 (N_24446,N_23760,N_23246);
or U24447 (N_24447,N_23225,N_23738);
nor U24448 (N_24448,N_23590,N_23403);
and U24449 (N_24449,N_23320,N_23414);
nand U24450 (N_24450,N_23848,N_23829);
or U24451 (N_24451,N_23971,N_23800);
xnor U24452 (N_24452,N_23267,N_23380);
xor U24453 (N_24453,N_23896,N_23781);
and U24454 (N_24454,N_23323,N_23356);
xnor U24455 (N_24455,N_23988,N_23501);
nand U24456 (N_24456,N_23444,N_23581);
and U24457 (N_24457,N_23096,N_23321);
and U24458 (N_24458,N_23729,N_23786);
xor U24459 (N_24459,N_23515,N_23369);
nor U24460 (N_24460,N_23049,N_23582);
xor U24461 (N_24461,N_23449,N_23553);
and U24462 (N_24462,N_23053,N_23549);
or U24463 (N_24463,N_23289,N_23640);
or U24464 (N_24464,N_23446,N_23682);
or U24465 (N_24465,N_23939,N_23660);
nor U24466 (N_24466,N_23281,N_23790);
or U24467 (N_24467,N_23837,N_23398);
nor U24468 (N_24468,N_23789,N_23958);
nor U24469 (N_24469,N_23075,N_23257);
or U24470 (N_24470,N_23306,N_23736);
xnor U24471 (N_24471,N_23200,N_23506);
or U24472 (N_24472,N_23895,N_23984);
nand U24473 (N_24473,N_23551,N_23456);
and U24474 (N_24474,N_23923,N_23645);
xnor U24475 (N_24475,N_23951,N_23979);
and U24476 (N_24476,N_23558,N_23746);
xor U24477 (N_24477,N_23227,N_23158);
nor U24478 (N_24478,N_23350,N_23853);
or U24479 (N_24479,N_23908,N_23410);
and U24480 (N_24480,N_23961,N_23701);
xnor U24481 (N_24481,N_23099,N_23562);
and U24482 (N_24482,N_23024,N_23518);
and U24483 (N_24483,N_23373,N_23393);
nor U24484 (N_24484,N_23423,N_23841);
nand U24485 (N_24485,N_23630,N_23921);
nand U24486 (N_24486,N_23105,N_23517);
and U24487 (N_24487,N_23717,N_23960);
or U24488 (N_24488,N_23483,N_23833);
nor U24489 (N_24489,N_23478,N_23095);
nand U24490 (N_24490,N_23758,N_23286);
and U24491 (N_24491,N_23883,N_23808);
nor U24492 (N_24492,N_23265,N_23445);
and U24493 (N_24493,N_23792,N_23484);
nand U24494 (N_24494,N_23555,N_23368);
and U24495 (N_24495,N_23799,N_23481);
nor U24496 (N_24496,N_23006,N_23204);
xnor U24497 (N_24497,N_23375,N_23692);
and U24498 (N_24498,N_23098,N_23412);
xor U24499 (N_24499,N_23452,N_23894);
xor U24500 (N_24500,N_23018,N_23137);
nand U24501 (N_24501,N_23887,N_23648);
or U24502 (N_24502,N_23983,N_23661);
xor U24503 (N_24503,N_23086,N_23012);
or U24504 (N_24504,N_23781,N_23244);
nand U24505 (N_24505,N_23263,N_23598);
or U24506 (N_24506,N_23953,N_23466);
or U24507 (N_24507,N_23339,N_23202);
or U24508 (N_24508,N_23828,N_23776);
and U24509 (N_24509,N_23189,N_23991);
nand U24510 (N_24510,N_23485,N_23148);
and U24511 (N_24511,N_23208,N_23209);
or U24512 (N_24512,N_23957,N_23913);
or U24513 (N_24513,N_23056,N_23902);
xor U24514 (N_24514,N_23338,N_23868);
xnor U24515 (N_24515,N_23135,N_23988);
nor U24516 (N_24516,N_23011,N_23667);
and U24517 (N_24517,N_23017,N_23471);
or U24518 (N_24518,N_23982,N_23163);
nor U24519 (N_24519,N_23783,N_23142);
or U24520 (N_24520,N_23845,N_23407);
nor U24521 (N_24521,N_23076,N_23851);
and U24522 (N_24522,N_23745,N_23559);
or U24523 (N_24523,N_23329,N_23987);
xnor U24524 (N_24524,N_23760,N_23251);
nor U24525 (N_24525,N_23320,N_23192);
nand U24526 (N_24526,N_23967,N_23682);
xnor U24527 (N_24527,N_23239,N_23643);
nand U24528 (N_24528,N_23334,N_23486);
nand U24529 (N_24529,N_23947,N_23498);
and U24530 (N_24530,N_23467,N_23841);
nor U24531 (N_24531,N_23875,N_23039);
or U24532 (N_24532,N_23818,N_23051);
and U24533 (N_24533,N_23158,N_23399);
nor U24534 (N_24534,N_23480,N_23671);
xor U24535 (N_24535,N_23060,N_23432);
nand U24536 (N_24536,N_23220,N_23590);
nand U24537 (N_24537,N_23443,N_23465);
nor U24538 (N_24538,N_23571,N_23683);
or U24539 (N_24539,N_23709,N_23144);
xor U24540 (N_24540,N_23610,N_23775);
nand U24541 (N_24541,N_23699,N_23684);
nor U24542 (N_24542,N_23110,N_23945);
and U24543 (N_24543,N_23188,N_23437);
and U24544 (N_24544,N_23665,N_23695);
xnor U24545 (N_24545,N_23753,N_23375);
nand U24546 (N_24546,N_23913,N_23575);
or U24547 (N_24547,N_23935,N_23660);
or U24548 (N_24548,N_23287,N_23695);
or U24549 (N_24549,N_23427,N_23137);
nor U24550 (N_24550,N_23034,N_23594);
nand U24551 (N_24551,N_23896,N_23220);
nor U24552 (N_24552,N_23238,N_23817);
and U24553 (N_24553,N_23702,N_23925);
nand U24554 (N_24554,N_23324,N_23714);
nand U24555 (N_24555,N_23241,N_23685);
nor U24556 (N_24556,N_23349,N_23786);
and U24557 (N_24557,N_23565,N_23158);
xor U24558 (N_24558,N_23797,N_23147);
or U24559 (N_24559,N_23024,N_23490);
nor U24560 (N_24560,N_23020,N_23383);
and U24561 (N_24561,N_23473,N_23010);
nor U24562 (N_24562,N_23263,N_23816);
xnor U24563 (N_24563,N_23268,N_23863);
xnor U24564 (N_24564,N_23484,N_23983);
nand U24565 (N_24565,N_23560,N_23160);
and U24566 (N_24566,N_23396,N_23072);
nand U24567 (N_24567,N_23402,N_23267);
xor U24568 (N_24568,N_23195,N_23835);
xor U24569 (N_24569,N_23976,N_23845);
and U24570 (N_24570,N_23515,N_23280);
nand U24571 (N_24571,N_23739,N_23876);
or U24572 (N_24572,N_23343,N_23579);
xor U24573 (N_24573,N_23655,N_23912);
nand U24574 (N_24574,N_23044,N_23437);
or U24575 (N_24575,N_23352,N_23096);
nand U24576 (N_24576,N_23988,N_23945);
nor U24577 (N_24577,N_23143,N_23928);
xor U24578 (N_24578,N_23720,N_23052);
nor U24579 (N_24579,N_23015,N_23686);
nand U24580 (N_24580,N_23454,N_23095);
and U24581 (N_24581,N_23451,N_23413);
xor U24582 (N_24582,N_23784,N_23085);
nor U24583 (N_24583,N_23666,N_23646);
and U24584 (N_24584,N_23939,N_23861);
xor U24585 (N_24585,N_23479,N_23598);
nor U24586 (N_24586,N_23941,N_23222);
nand U24587 (N_24587,N_23889,N_23555);
or U24588 (N_24588,N_23035,N_23041);
or U24589 (N_24589,N_23743,N_23608);
or U24590 (N_24590,N_23862,N_23627);
nand U24591 (N_24591,N_23615,N_23652);
xor U24592 (N_24592,N_23656,N_23111);
and U24593 (N_24593,N_23918,N_23605);
nand U24594 (N_24594,N_23025,N_23172);
nor U24595 (N_24595,N_23729,N_23091);
nand U24596 (N_24596,N_23198,N_23021);
xnor U24597 (N_24597,N_23805,N_23430);
and U24598 (N_24598,N_23574,N_23341);
nand U24599 (N_24599,N_23959,N_23805);
and U24600 (N_24600,N_23924,N_23551);
and U24601 (N_24601,N_23049,N_23644);
xor U24602 (N_24602,N_23388,N_23063);
xnor U24603 (N_24603,N_23194,N_23147);
and U24604 (N_24604,N_23943,N_23915);
or U24605 (N_24605,N_23365,N_23360);
and U24606 (N_24606,N_23566,N_23304);
and U24607 (N_24607,N_23425,N_23888);
xor U24608 (N_24608,N_23449,N_23565);
nand U24609 (N_24609,N_23533,N_23766);
xnor U24610 (N_24610,N_23187,N_23796);
xor U24611 (N_24611,N_23458,N_23573);
xor U24612 (N_24612,N_23427,N_23114);
or U24613 (N_24613,N_23546,N_23958);
and U24614 (N_24614,N_23642,N_23680);
and U24615 (N_24615,N_23533,N_23356);
xnor U24616 (N_24616,N_23433,N_23578);
or U24617 (N_24617,N_23492,N_23647);
xnor U24618 (N_24618,N_23894,N_23255);
and U24619 (N_24619,N_23841,N_23532);
or U24620 (N_24620,N_23735,N_23445);
or U24621 (N_24621,N_23473,N_23961);
nor U24622 (N_24622,N_23096,N_23266);
nor U24623 (N_24623,N_23303,N_23180);
and U24624 (N_24624,N_23081,N_23256);
xor U24625 (N_24625,N_23410,N_23366);
or U24626 (N_24626,N_23912,N_23972);
or U24627 (N_24627,N_23826,N_23372);
nor U24628 (N_24628,N_23125,N_23279);
and U24629 (N_24629,N_23610,N_23554);
or U24630 (N_24630,N_23728,N_23184);
xor U24631 (N_24631,N_23848,N_23309);
or U24632 (N_24632,N_23894,N_23106);
nand U24633 (N_24633,N_23193,N_23441);
xnor U24634 (N_24634,N_23132,N_23324);
nor U24635 (N_24635,N_23903,N_23080);
xor U24636 (N_24636,N_23570,N_23946);
and U24637 (N_24637,N_23519,N_23403);
and U24638 (N_24638,N_23701,N_23426);
xnor U24639 (N_24639,N_23573,N_23013);
or U24640 (N_24640,N_23661,N_23830);
or U24641 (N_24641,N_23847,N_23668);
nand U24642 (N_24642,N_23053,N_23199);
nand U24643 (N_24643,N_23078,N_23532);
and U24644 (N_24644,N_23174,N_23161);
nand U24645 (N_24645,N_23865,N_23996);
nand U24646 (N_24646,N_23250,N_23279);
nor U24647 (N_24647,N_23819,N_23317);
xor U24648 (N_24648,N_23253,N_23749);
nand U24649 (N_24649,N_23744,N_23408);
and U24650 (N_24650,N_23590,N_23122);
nand U24651 (N_24651,N_23828,N_23895);
nand U24652 (N_24652,N_23489,N_23134);
nand U24653 (N_24653,N_23109,N_23105);
and U24654 (N_24654,N_23481,N_23540);
xnor U24655 (N_24655,N_23808,N_23299);
xnor U24656 (N_24656,N_23750,N_23912);
xnor U24657 (N_24657,N_23023,N_23573);
or U24658 (N_24658,N_23208,N_23547);
nand U24659 (N_24659,N_23893,N_23524);
nor U24660 (N_24660,N_23922,N_23267);
xnor U24661 (N_24661,N_23385,N_23510);
or U24662 (N_24662,N_23402,N_23080);
nor U24663 (N_24663,N_23213,N_23784);
nor U24664 (N_24664,N_23419,N_23221);
nand U24665 (N_24665,N_23523,N_23558);
nand U24666 (N_24666,N_23391,N_23897);
nand U24667 (N_24667,N_23646,N_23350);
or U24668 (N_24668,N_23193,N_23985);
nor U24669 (N_24669,N_23407,N_23733);
xnor U24670 (N_24670,N_23124,N_23901);
and U24671 (N_24671,N_23495,N_23458);
nand U24672 (N_24672,N_23411,N_23854);
nand U24673 (N_24673,N_23227,N_23319);
and U24674 (N_24674,N_23930,N_23137);
and U24675 (N_24675,N_23485,N_23560);
nor U24676 (N_24676,N_23728,N_23118);
or U24677 (N_24677,N_23694,N_23009);
nand U24678 (N_24678,N_23189,N_23409);
or U24679 (N_24679,N_23607,N_23483);
nand U24680 (N_24680,N_23336,N_23385);
nand U24681 (N_24681,N_23853,N_23981);
nor U24682 (N_24682,N_23528,N_23400);
xnor U24683 (N_24683,N_23578,N_23328);
xnor U24684 (N_24684,N_23109,N_23807);
nor U24685 (N_24685,N_23824,N_23344);
and U24686 (N_24686,N_23667,N_23799);
nor U24687 (N_24687,N_23435,N_23793);
xnor U24688 (N_24688,N_23569,N_23621);
xnor U24689 (N_24689,N_23776,N_23931);
or U24690 (N_24690,N_23568,N_23931);
xor U24691 (N_24691,N_23275,N_23580);
nand U24692 (N_24692,N_23661,N_23006);
xnor U24693 (N_24693,N_23223,N_23541);
nand U24694 (N_24694,N_23203,N_23854);
and U24695 (N_24695,N_23770,N_23929);
nand U24696 (N_24696,N_23596,N_23645);
xnor U24697 (N_24697,N_23406,N_23619);
xnor U24698 (N_24698,N_23945,N_23713);
xor U24699 (N_24699,N_23041,N_23313);
or U24700 (N_24700,N_23709,N_23395);
xor U24701 (N_24701,N_23611,N_23853);
xnor U24702 (N_24702,N_23477,N_23712);
or U24703 (N_24703,N_23120,N_23960);
or U24704 (N_24704,N_23087,N_23253);
xor U24705 (N_24705,N_23844,N_23221);
nand U24706 (N_24706,N_23627,N_23777);
nor U24707 (N_24707,N_23177,N_23750);
or U24708 (N_24708,N_23301,N_23389);
xnor U24709 (N_24709,N_23249,N_23507);
xnor U24710 (N_24710,N_23490,N_23079);
or U24711 (N_24711,N_23922,N_23653);
and U24712 (N_24712,N_23859,N_23434);
and U24713 (N_24713,N_23602,N_23023);
xor U24714 (N_24714,N_23331,N_23643);
xor U24715 (N_24715,N_23312,N_23095);
nor U24716 (N_24716,N_23348,N_23748);
nand U24717 (N_24717,N_23092,N_23492);
and U24718 (N_24718,N_23331,N_23458);
xnor U24719 (N_24719,N_23694,N_23063);
xor U24720 (N_24720,N_23261,N_23856);
nor U24721 (N_24721,N_23835,N_23877);
nand U24722 (N_24722,N_23647,N_23843);
and U24723 (N_24723,N_23317,N_23762);
or U24724 (N_24724,N_23850,N_23722);
nor U24725 (N_24725,N_23209,N_23101);
nor U24726 (N_24726,N_23471,N_23992);
and U24727 (N_24727,N_23863,N_23805);
or U24728 (N_24728,N_23281,N_23935);
or U24729 (N_24729,N_23748,N_23196);
nand U24730 (N_24730,N_23579,N_23934);
nand U24731 (N_24731,N_23514,N_23943);
nand U24732 (N_24732,N_23192,N_23016);
nand U24733 (N_24733,N_23328,N_23403);
nor U24734 (N_24734,N_23352,N_23272);
nor U24735 (N_24735,N_23970,N_23124);
xor U24736 (N_24736,N_23357,N_23384);
nor U24737 (N_24737,N_23062,N_23203);
nor U24738 (N_24738,N_23687,N_23035);
nand U24739 (N_24739,N_23659,N_23606);
or U24740 (N_24740,N_23137,N_23952);
nand U24741 (N_24741,N_23886,N_23946);
nor U24742 (N_24742,N_23657,N_23894);
and U24743 (N_24743,N_23774,N_23855);
or U24744 (N_24744,N_23195,N_23790);
xor U24745 (N_24745,N_23485,N_23130);
or U24746 (N_24746,N_23002,N_23250);
or U24747 (N_24747,N_23751,N_23574);
nor U24748 (N_24748,N_23760,N_23168);
xnor U24749 (N_24749,N_23445,N_23260);
or U24750 (N_24750,N_23690,N_23274);
xor U24751 (N_24751,N_23781,N_23553);
nor U24752 (N_24752,N_23776,N_23291);
nand U24753 (N_24753,N_23248,N_23376);
and U24754 (N_24754,N_23243,N_23996);
nand U24755 (N_24755,N_23337,N_23221);
and U24756 (N_24756,N_23005,N_23924);
or U24757 (N_24757,N_23211,N_23808);
or U24758 (N_24758,N_23063,N_23813);
nand U24759 (N_24759,N_23660,N_23964);
nor U24760 (N_24760,N_23176,N_23131);
xnor U24761 (N_24761,N_23422,N_23955);
or U24762 (N_24762,N_23496,N_23313);
xor U24763 (N_24763,N_23829,N_23240);
nand U24764 (N_24764,N_23983,N_23078);
and U24765 (N_24765,N_23140,N_23744);
nor U24766 (N_24766,N_23656,N_23677);
and U24767 (N_24767,N_23894,N_23670);
or U24768 (N_24768,N_23857,N_23995);
or U24769 (N_24769,N_23712,N_23775);
or U24770 (N_24770,N_23579,N_23450);
nor U24771 (N_24771,N_23459,N_23712);
nor U24772 (N_24772,N_23452,N_23025);
nand U24773 (N_24773,N_23109,N_23567);
nor U24774 (N_24774,N_23864,N_23525);
and U24775 (N_24775,N_23481,N_23746);
or U24776 (N_24776,N_23581,N_23288);
nor U24777 (N_24777,N_23018,N_23498);
or U24778 (N_24778,N_23818,N_23553);
and U24779 (N_24779,N_23073,N_23714);
nor U24780 (N_24780,N_23712,N_23140);
nor U24781 (N_24781,N_23713,N_23740);
or U24782 (N_24782,N_23879,N_23662);
nor U24783 (N_24783,N_23405,N_23077);
and U24784 (N_24784,N_23895,N_23582);
nand U24785 (N_24785,N_23412,N_23135);
or U24786 (N_24786,N_23850,N_23124);
xnor U24787 (N_24787,N_23817,N_23787);
and U24788 (N_24788,N_23376,N_23005);
and U24789 (N_24789,N_23702,N_23326);
xor U24790 (N_24790,N_23763,N_23606);
nand U24791 (N_24791,N_23752,N_23138);
and U24792 (N_24792,N_23033,N_23059);
or U24793 (N_24793,N_23529,N_23003);
and U24794 (N_24794,N_23238,N_23075);
and U24795 (N_24795,N_23798,N_23114);
or U24796 (N_24796,N_23668,N_23171);
nor U24797 (N_24797,N_23132,N_23194);
or U24798 (N_24798,N_23625,N_23299);
or U24799 (N_24799,N_23855,N_23123);
nor U24800 (N_24800,N_23278,N_23427);
or U24801 (N_24801,N_23584,N_23985);
nor U24802 (N_24802,N_23064,N_23615);
and U24803 (N_24803,N_23798,N_23678);
or U24804 (N_24804,N_23198,N_23583);
nor U24805 (N_24805,N_23171,N_23340);
and U24806 (N_24806,N_23489,N_23329);
nand U24807 (N_24807,N_23198,N_23662);
nor U24808 (N_24808,N_23725,N_23102);
xor U24809 (N_24809,N_23366,N_23035);
xnor U24810 (N_24810,N_23454,N_23787);
nand U24811 (N_24811,N_23580,N_23863);
or U24812 (N_24812,N_23242,N_23717);
and U24813 (N_24813,N_23813,N_23156);
and U24814 (N_24814,N_23873,N_23735);
nor U24815 (N_24815,N_23020,N_23793);
and U24816 (N_24816,N_23128,N_23317);
xor U24817 (N_24817,N_23626,N_23434);
nor U24818 (N_24818,N_23475,N_23494);
xor U24819 (N_24819,N_23910,N_23804);
nand U24820 (N_24820,N_23685,N_23891);
or U24821 (N_24821,N_23839,N_23002);
and U24822 (N_24822,N_23263,N_23278);
xor U24823 (N_24823,N_23271,N_23471);
xnor U24824 (N_24824,N_23040,N_23198);
or U24825 (N_24825,N_23357,N_23391);
nor U24826 (N_24826,N_23788,N_23853);
nor U24827 (N_24827,N_23527,N_23795);
xor U24828 (N_24828,N_23087,N_23070);
nand U24829 (N_24829,N_23605,N_23724);
xor U24830 (N_24830,N_23868,N_23539);
nor U24831 (N_24831,N_23224,N_23090);
and U24832 (N_24832,N_23211,N_23192);
and U24833 (N_24833,N_23967,N_23033);
and U24834 (N_24834,N_23564,N_23347);
nor U24835 (N_24835,N_23524,N_23378);
and U24836 (N_24836,N_23487,N_23479);
nor U24837 (N_24837,N_23292,N_23684);
nor U24838 (N_24838,N_23109,N_23059);
xnor U24839 (N_24839,N_23410,N_23050);
nor U24840 (N_24840,N_23791,N_23578);
and U24841 (N_24841,N_23720,N_23348);
nand U24842 (N_24842,N_23188,N_23357);
nand U24843 (N_24843,N_23529,N_23574);
nand U24844 (N_24844,N_23085,N_23572);
and U24845 (N_24845,N_23427,N_23636);
nand U24846 (N_24846,N_23885,N_23279);
nand U24847 (N_24847,N_23899,N_23606);
nor U24848 (N_24848,N_23112,N_23230);
nand U24849 (N_24849,N_23820,N_23528);
and U24850 (N_24850,N_23020,N_23662);
nor U24851 (N_24851,N_23013,N_23507);
and U24852 (N_24852,N_23356,N_23372);
and U24853 (N_24853,N_23209,N_23088);
nand U24854 (N_24854,N_23295,N_23599);
and U24855 (N_24855,N_23904,N_23017);
nand U24856 (N_24856,N_23589,N_23374);
nor U24857 (N_24857,N_23402,N_23423);
xnor U24858 (N_24858,N_23361,N_23474);
nor U24859 (N_24859,N_23879,N_23449);
nand U24860 (N_24860,N_23906,N_23629);
nor U24861 (N_24861,N_23580,N_23838);
nor U24862 (N_24862,N_23512,N_23528);
xor U24863 (N_24863,N_23103,N_23835);
or U24864 (N_24864,N_23188,N_23289);
xor U24865 (N_24865,N_23700,N_23316);
xnor U24866 (N_24866,N_23477,N_23245);
nor U24867 (N_24867,N_23925,N_23690);
nand U24868 (N_24868,N_23177,N_23579);
xnor U24869 (N_24869,N_23005,N_23894);
nor U24870 (N_24870,N_23334,N_23096);
xnor U24871 (N_24871,N_23784,N_23874);
nand U24872 (N_24872,N_23823,N_23370);
and U24873 (N_24873,N_23328,N_23651);
and U24874 (N_24874,N_23046,N_23085);
and U24875 (N_24875,N_23356,N_23085);
nand U24876 (N_24876,N_23691,N_23311);
or U24877 (N_24877,N_23617,N_23842);
nor U24878 (N_24878,N_23085,N_23111);
and U24879 (N_24879,N_23032,N_23529);
xor U24880 (N_24880,N_23086,N_23846);
nand U24881 (N_24881,N_23503,N_23007);
or U24882 (N_24882,N_23898,N_23672);
xnor U24883 (N_24883,N_23700,N_23350);
or U24884 (N_24884,N_23177,N_23134);
and U24885 (N_24885,N_23994,N_23316);
and U24886 (N_24886,N_23676,N_23758);
nand U24887 (N_24887,N_23174,N_23888);
xnor U24888 (N_24888,N_23188,N_23591);
nand U24889 (N_24889,N_23559,N_23106);
or U24890 (N_24890,N_23480,N_23422);
nand U24891 (N_24891,N_23568,N_23993);
xor U24892 (N_24892,N_23212,N_23858);
nor U24893 (N_24893,N_23806,N_23629);
nand U24894 (N_24894,N_23643,N_23449);
nor U24895 (N_24895,N_23075,N_23098);
xor U24896 (N_24896,N_23760,N_23739);
nor U24897 (N_24897,N_23169,N_23317);
and U24898 (N_24898,N_23464,N_23374);
nand U24899 (N_24899,N_23581,N_23582);
nand U24900 (N_24900,N_23496,N_23293);
nor U24901 (N_24901,N_23481,N_23861);
and U24902 (N_24902,N_23303,N_23584);
or U24903 (N_24903,N_23261,N_23114);
or U24904 (N_24904,N_23140,N_23090);
nor U24905 (N_24905,N_23052,N_23243);
and U24906 (N_24906,N_23042,N_23502);
nor U24907 (N_24907,N_23242,N_23167);
and U24908 (N_24908,N_23343,N_23261);
nor U24909 (N_24909,N_23925,N_23317);
nor U24910 (N_24910,N_23962,N_23570);
nand U24911 (N_24911,N_23927,N_23937);
or U24912 (N_24912,N_23187,N_23253);
nand U24913 (N_24913,N_23691,N_23651);
nand U24914 (N_24914,N_23687,N_23550);
nor U24915 (N_24915,N_23981,N_23658);
xnor U24916 (N_24916,N_23410,N_23753);
xnor U24917 (N_24917,N_23868,N_23448);
xor U24918 (N_24918,N_23077,N_23779);
nor U24919 (N_24919,N_23973,N_23450);
xnor U24920 (N_24920,N_23683,N_23228);
xnor U24921 (N_24921,N_23898,N_23934);
or U24922 (N_24922,N_23680,N_23577);
nor U24923 (N_24923,N_23227,N_23582);
nand U24924 (N_24924,N_23793,N_23250);
and U24925 (N_24925,N_23016,N_23358);
and U24926 (N_24926,N_23073,N_23142);
and U24927 (N_24927,N_23756,N_23002);
nor U24928 (N_24928,N_23240,N_23832);
nor U24929 (N_24929,N_23817,N_23759);
nor U24930 (N_24930,N_23229,N_23960);
nor U24931 (N_24931,N_23271,N_23689);
xor U24932 (N_24932,N_23852,N_23756);
and U24933 (N_24933,N_23429,N_23819);
and U24934 (N_24934,N_23555,N_23546);
nor U24935 (N_24935,N_23628,N_23804);
xnor U24936 (N_24936,N_23790,N_23530);
xnor U24937 (N_24937,N_23584,N_23274);
nand U24938 (N_24938,N_23583,N_23325);
or U24939 (N_24939,N_23095,N_23986);
and U24940 (N_24940,N_23158,N_23055);
nand U24941 (N_24941,N_23332,N_23569);
xor U24942 (N_24942,N_23989,N_23018);
or U24943 (N_24943,N_23428,N_23017);
nand U24944 (N_24944,N_23120,N_23245);
xor U24945 (N_24945,N_23603,N_23996);
xnor U24946 (N_24946,N_23710,N_23010);
nand U24947 (N_24947,N_23734,N_23483);
or U24948 (N_24948,N_23498,N_23752);
or U24949 (N_24949,N_23158,N_23213);
nor U24950 (N_24950,N_23574,N_23763);
xor U24951 (N_24951,N_23598,N_23311);
xor U24952 (N_24952,N_23880,N_23365);
or U24953 (N_24953,N_23051,N_23007);
nand U24954 (N_24954,N_23959,N_23498);
xor U24955 (N_24955,N_23353,N_23095);
and U24956 (N_24956,N_23677,N_23545);
nand U24957 (N_24957,N_23891,N_23746);
nand U24958 (N_24958,N_23554,N_23027);
nand U24959 (N_24959,N_23483,N_23676);
nor U24960 (N_24960,N_23263,N_23485);
nor U24961 (N_24961,N_23246,N_23674);
nor U24962 (N_24962,N_23949,N_23851);
nand U24963 (N_24963,N_23013,N_23421);
nand U24964 (N_24964,N_23410,N_23335);
nor U24965 (N_24965,N_23516,N_23864);
or U24966 (N_24966,N_23877,N_23059);
xor U24967 (N_24967,N_23998,N_23247);
nand U24968 (N_24968,N_23414,N_23821);
xor U24969 (N_24969,N_23719,N_23289);
and U24970 (N_24970,N_23789,N_23107);
or U24971 (N_24971,N_23122,N_23117);
or U24972 (N_24972,N_23839,N_23483);
xnor U24973 (N_24973,N_23276,N_23142);
and U24974 (N_24974,N_23904,N_23606);
xnor U24975 (N_24975,N_23213,N_23491);
xor U24976 (N_24976,N_23927,N_23941);
xor U24977 (N_24977,N_23202,N_23433);
and U24978 (N_24978,N_23645,N_23757);
xnor U24979 (N_24979,N_23740,N_23447);
and U24980 (N_24980,N_23893,N_23955);
or U24981 (N_24981,N_23475,N_23176);
nor U24982 (N_24982,N_23203,N_23683);
nand U24983 (N_24983,N_23915,N_23480);
or U24984 (N_24984,N_23854,N_23489);
or U24985 (N_24985,N_23599,N_23905);
and U24986 (N_24986,N_23504,N_23397);
nand U24987 (N_24987,N_23634,N_23111);
nand U24988 (N_24988,N_23090,N_23691);
or U24989 (N_24989,N_23772,N_23595);
xor U24990 (N_24990,N_23574,N_23071);
nor U24991 (N_24991,N_23893,N_23870);
or U24992 (N_24992,N_23030,N_23788);
xnor U24993 (N_24993,N_23264,N_23645);
nand U24994 (N_24994,N_23154,N_23666);
or U24995 (N_24995,N_23872,N_23333);
nor U24996 (N_24996,N_23368,N_23106);
xor U24997 (N_24997,N_23650,N_23255);
xnor U24998 (N_24998,N_23650,N_23923);
xnor U24999 (N_24999,N_23157,N_23270);
xor U25000 (N_25000,N_24255,N_24772);
xor U25001 (N_25001,N_24815,N_24812);
nor U25002 (N_25002,N_24161,N_24220);
and U25003 (N_25003,N_24333,N_24919);
and U25004 (N_25004,N_24711,N_24915);
xnor U25005 (N_25005,N_24501,N_24642);
nand U25006 (N_25006,N_24735,N_24877);
and U25007 (N_25007,N_24669,N_24571);
and U25008 (N_25008,N_24419,N_24310);
and U25009 (N_25009,N_24362,N_24949);
nand U25010 (N_25010,N_24903,N_24613);
nor U25011 (N_25011,N_24562,N_24207);
nand U25012 (N_25012,N_24496,N_24216);
xor U25013 (N_25013,N_24175,N_24533);
nor U25014 (N_25014,N_24058,N_24403);
nand U25015 (N_25015,N_24884,N_24347);
nor U25016 (N_25016,N_24155,N_24345);
xor U25017 (N_25017,N_24371,N_24957);
nor U25018 (N_25018,N_24367,N_24616);
nor U25019 (N_25019,N_24498,N_24311);
and U25020 (N_25020,N_24809,N_24340);
and U25021 (N_25021,N_24726,N_24064);
nand U25022 (N_25022,N_24661,N_24689);
nor U25023 (N_25023,N_24793,N_24757);
and U25024 (N_25024,N_24628,N_24690);
or U25025 (N_25025,N_24872,N_24750);
or U25026 (N_25026,N_24704,N_24331);
nand U25027 (N_25027,N_24684,N_24626);
nor U25028 (N_25028,N_24485,N_24452);
or U25029 (N_25029,N_24062,N_24830);
and U25030 (N_25030,N_24540,N_24154);
nand U25031 (N_25031,N_24699,N_24837);
xnor U25032 (N_25032,N_24682,N_24404);
or U25033 (N_25033,N_24434,N_24094);
and U25034 (N_25034,N_24104,N_24103);
xor U25035 (N_25035,N_24596,N_24924);
nand U25036 (N_25036,N_24388,N_24999);
xnor U25037 (N_25037,N_24017,N_24728);
and U25038 (N_25038,N_24210,N_24226);
nor U25039 (N_25039,N_24379,N_24851);
or U25040 (N_25040,N_24865,N_24260);
and U25041 (N_25041,N_24709,N_24989);
nor U25042 (N_25042,N_24391,N_24576);
nand U25043 (N_25043,N_24927,N_24027);
or U25044 (N_25044,N_24916,N_24363);
nor U25045 (N_25045,N_24636,N_24724);
or U25046 (N_25046,N_24753,N_24836);
nor U25047 (N_25047,N_24779,N_24184);
or U25048 (N_25048,N_24010,N_24209);
or U25049 (N_25049,N_24551,N_24511);
and U25050 (N_25050,N_24171,N_24147);
or U25051 (N_25051,N_24675,N_24022);
xnor U25052 (N_25052,N_24470,N_24464);
and U25053 (N_25053,N_24713,N_24280);
nor U25054 (N_25054,N_24202,N_24433);
nor U25055 (N_25055,N_24276,N_24284);
nor U25056 (N_25056,N_24274,N_24710);
nor U25057 (N_25057,N_24273,N_24931);
xor U25058 (N_25058,N_24194,N_24866);
or U25059 (N_25059,N_24401,N_24494);
xnor U25060 (N_25060,N_24023,N_24467);
xnor U25061 (N_25061,N_24488,N_24799);
nor U25062 (N_25062,N_24900,N_24195);
or U25063 (N_25063,N_24676,N_24878);
xnor U25064 (N_25064,N_24818,N_24248);
and U25065 (N_25065,N_24933,N_24893);
or U25066 (N_25066,N_24290,N_24415);
and U25067 (N_25067,N_24440,N_24688);
nand U25068 (N_25068,N_24460,N_24702);
and U25069 (N_25069,N_24230,N_24905);
nor U25070 (N_25070,N_24083,N_24244);
and U25071 (N_25071,N_24707,N_24126);
and U25072 (N_25072,N_24835,N_24348);
and U25073 (N_25073,N_24431,N_24219);
and U25074 (N_25074,N_24622,N_24887);
xnor U25075 (N_25075,N_24674,N_24639);
nor U25076 (N_25076,N_24538,N_24984);
nor U25077 (N_25077,N_24876,N_24070);
xor U25078 (N_25078,N_24605,N_24518);
xor U25079 (N_25079,N_24937,N_24177);
xnor U25080 (N_25080,N_24664,N_24738);
nor U25081 (N_25081,N_24287,N_24638);
or U25082 (N_25082,N_24162,N_24392);
nor U25083 (N_25083,N_24838,N_24268);
or U25084 (N_25084,N_24473,N_24354);
nand U25085 (N_25085,N_24574,N_24668);
nand U25086 (N_25086,N_24867,N_24257);
and U25087 (N_25087,N_24503,N_24665);
nor U25088 (N_25088,N_24173,N_24071);
nand U25089 (N_25089,N_24625,N_24890);
or U25090 (N_25090,N_24353,N_24030);
and U25091 (N_25091,N_24981,N_24833);
xor U25092 (N_25092,N_24577,N_24124);
xor U25093 (N_25093,N_24962,N_24373);
xor U25094 (N_25094,N_24519,N_24364);
and U25095 (N_25095,N_24293,N_24547);
nand U25096 (N_25096,N_24304,N_24253);
nor U25097 (N_25097,N_24634,N_24493);
nor U25098 (N_25098,N_24250,N_24918);
or U25099 (N_25099,N_24424,N_24108);
or U25100 (N_25100,N_24294,N_24151);
or U25101 (N_25101,N_24059,N_24411);
xor U25102 (N_25102,N_24899,N_24204);
or U25103 (N_25103,N_24040,N_24343);
and U25104 (N_25104,N_24659,N_24015);
xnor U25105 (N_25105,N_24934,N_24529);
or U25106 (N_25106,N_24045,N_24536);
xnor U25107 (N_25107,N_24445,N_24858);
and U25108 (N_25108,N_24930,N_24959);
nand U25109 (N_25109,N_24604,N_24384);
nand U25110 (N_25110,N_24188,N_24249);
xnor U25111 (N_25111,N_24454,N_24881);
nor U25112 (N_25112,N_24901,N_24802);
nor U25113 (N_25113,N_24137,N_24206);
xnor U25114 (N_25114,N_24760,N_24006);
and U25115 (N_25115,N_24050,N_24681);
and U25116 (N_25116,N_24853,N_24176);
nor U25117 (N_25117,N_24745,N_24279);
xnor U25118 (N_25118,N_24546,N_24555);
nand U25119 (N_25119,N_24964,N_24289);
and U25120 (N_25120,N_24465,N_24861);
and U25121 (N_25121,N_24978,N_24283);
or U25122 (N_25122,N_24009,N_24941);
nor U25123 (N_25123,N_24068,N_24559);
or U25124 (N_25124,N_24208,N_24992);
or U25125 (N_25125,N_24840,N_24971);
nand U25126 (N_25126,N_24448,N_24939);
xor U25127 (N_25127,N_24489,N_24338);
or U25128 (N_25128,N_24775,N_24556);
nor U25129 (N_25129,N_24146,N_24589);
nand U25130 (N_25130,N_24116,N_24966);
or U25131 (N_25131,N_24641,N_24599);
nor U25132 (N_25132,N_24839,N_24259);
xnor U25133 (N_25133,N_24048,N_24435);
nor U25134 (N_25134,N_24883,N_24288);
and U25135 (N_25135,N_24197,N_24459);
nor U25136 (N_25136,N_24698,N_24282);
xnor U25137 (N_25137,N_24826,N_24947);
nor U25138 (N_25138,N_24746,N_24951);
xnor U25139 (N_25139,N_24223,N_24317);
or U25140 (N_25140,N_24224,N_24967);
xnor U25141 (N_25141,N_24087,N_24233);
nor U25142 (N_25142,N_24038,N_24213);
nor U25143 (N_25143,N_24337,N_24123);
or U25144 (N_25144,N_24549,N_24850);
nor U25145 (N_25145,N_24456,N_24532);
nor U25146 (N_25146,N_24943,N_24285);
and U25147 (N_25147,N_24160,N_24408);
or U25148 (N_25148,N_24157,N_24381);
or U25149 (N_25149,N_24670,N_24410);
nand U25150 (N_25150,N_24004,N_24222);
nor U25151 (N_25151,N_24841,N_24564);
or U25152 (N_25152,N_24032,N_24522);
nand U25153 (N_25153,N_24380,N_24458);
nand U25154 (N_25154,N_24781,N_24590);
xor U25155 (N_25155,N_24429,N_24619);
and U25156 (N_25156,N_24407,N_24066);
nand U25157 (N_25157,N_24716,N_24142);
xnor U25158 (N_25158,N_24798,N_24139);
xnor U25159 (N_25159,N_24514,N_24028);
or U25160 (N_25160,N_24561,N_24221);
nor U25161 (N_25161,N_24422,N_24394);
or U25162 (N_25162,N_24857,N_24203);
and U25163 (N_25163,N_24717,N_24100);
xor U25164 (N_25164,N_24780,N_24860);
or U25165 (N_25165,N_24786,N_24752);
or U25166 (N_25166,N_24808,N_24648);
nor U25167 (N_25167,N_24683,N_24052);
nor U25168 (N_25168,N_24629,N_24953);
nand U25169 (N_25169,N_24200,N_24671);
nand U25170 (N_25170,N_24272,N_24791);
nor U25171 (N_25171,N_24080,N_24778);
xor U25172 (N_25172,N_24400,N_24056);
nand U25173 (N_25173,N_24266,N_24859);
xor U25174 (N_25174,N_24987,N_24660);
and U25175 (N_25175,N_24092,N_24148);
and U25176 (N_25176,N_24898,N_24495);
and U25177 (N_25177,N_24425,N_24275);
and U25178 (N_25178,N_24531,N_24679);
and U25179 (N_25179,N_24020,N_24358);
and U25180 (N_25180,N_24121,N_24201);
or U25181 (N_25181,N_24913,N_24880);
nor U25182 (N_25182,N_24955,N_24879);
nand U25183 (N_25183,N_24356,N_24297);
and U25184 (N_25184,N_24755,N_24972);
and U25185 (N_25185,N_24906,N_24784);
nand U25186 (N_25186,N_24178,N_24366);
xor U25187 (N_25187,N_24563,N_24041);
and U25188 (N_25188,N_24193,N_24088);
or U25189 (N_25189,N_24412,N_24932);
nand U25190 (N_25190,N_24455,N_24346);
nor U25191 (N_25191,N_24914,N_24097);
nor U25192 (N_25192,N_24695,N_24117);
nor U25193 (N_25193,N_24828,N_24043);
xor U25194 (N_25194,N_24870,N_24397);
and U25195 (N_25195,N_24262,N_24723);
xor U25196 (N_25196,N_24714,N_24766);
xor U25197 (N_25197,N_24462,N_24504);
and U25198 (N_25198,N_24653,N_24269);
or U25199 (N_25199,N_24483,N_24727);
xor U25200 (N_25200,N_24819,N_24073);
or U25201 (N_25201,N_24782,N_24342);
nor U25202 (N_25202,N_24657,N_24801);
nor U25203 (N_25203,N_24385,N_24600);
or U25204 (N_25204,N_24306,N_24457);
xnor U25205 (N_25205,N_24646,N_24891);
or U25206 (N_25206,N_24731,N_24387);
nor U25207 (N_25207,N_24990,N_24963);
nand U25208 (N_25208,N_24180,N_24067);
nand U25209 (N_25209,N_24003,N_24140);
xnor U25210 (N_25210,N_24278,N_24444);
or U25211 (N_25211,N_24921,N_24813);
and U25212 (N_25212,N_24803,N_24476);
nand U25213 (N_25213,N_24973,N_24994);
xor U25214 (N_25214,N_24189,N_24008);
nor U25215 (N_25215,N_24446,N_24982);
xnor U25216 (N_25216,N_24521,N_24398);
and U25217 (N_25217,N_24976,N_24512);
xor U25218 (N_25218,N_24243,N_24820);
nor U25219 (N_25219,N_24693,N_24748);
and U25220 (N_25220,N_24548,N_24302);
xnor U25221 (N_25221,N_24908,N_24795);
or U25222 (N_25222,N_24888,N_24938);
and U25223 (N_25223,N_24621,N_24214);
nor U25224 (N_25224,N_24399,N_24960);
nor U25225 (N_25225,N_24520,N_24946);
nor U25226 (N_25226,N_24036,N_24437);
xnor U25227 (N_25227,N_24507,N_24237);
nor U25228 (N_25228,N_24854,N_24570);
nor U25229 (N_25229,N_24736,N_24814);
nor U25230 (N_25230,N_24120,N_24252);
xor U25231 (N_25231,N_24261,N_24607);
or U25232 (N_25232,N_24614,N_24316);
and U25233 (N_25233,N_24078,N_24113);
or U25234 (N_25234,N_24300,N_24390);
nor U25235 (N_25235,N_24807,N_24344);
and U25236 (N_25236,N_24002,N_24430);
nor U25237 (N_25237,N_24701,N_24005);
or U25238 (N_25238,N_24560,N_24740);
nand U25239 (N_25239,N_24131,N_24537);
and U25240 (N_25240,N_24796,N_24361);
nand U25241 (N_25241,N_24662,N_24090);
nor U25242 (N_25242,N_24321,N_24831);
nand U25243 (N_25243,N_24703,N_24935);
xor U25244 (N_25244,N_24771,N_24086);
and U25245 (N_25245,N_24185,N_24119);
nor U25246 (N_25246,N_24240,N_24527);
or U25247 (N_25247,N_24238,N_24744);
nand U25248 (N_25248,N_24631,N_24319);
and U25249 (N_25249,N_24061,N_24940);
nand U25250 (N_25250,N_24788,N_24925);
xnor U25251 (N_25251,N_24095,N_24085);
and U25252 (N_25252,N_24827,N_24484);
nand U25253 (N_25253,N_24011,N_24152);
xor U25254 (N_25254,N_24132,N_24842);
nand U25255 (N_25255,N_24334,N_24609);
and U25256 (N_25256,N_24133,N_24725);
nand U25257 (N_25257,N_24948,N_24797);
and U25258 (N_25258,N_24479,N_24414);
and U25259 (N_25259,N_24658,N_24125);
xor U25260 (N_25260,N_24697,N_24322);
and U25261 (N_25261,N_24182,N_24037);
nand U25262 (N_25262,N_24477,N_24107);
nand U25263 (N_25263,N_24649,N_24583);
nor U25264 (N_25264,N_24428,N_24330);
and U25265 (N_25265,N_24307,N_24318);
nand U25266 (N_25266,N_24911,N_24482);
xor U25267 (N_25267,N_24236,N_24234);
nand U25268 (N_25268,N_24928,N_24118);
nand U25269 (N_25269,N_24747,N_24524);
and U25270 (N_25270,N_24611,N_24598);
nor U25271 (N_25271,N_24910,N_24375);
and U25272 (N_25272,N_24051,N_24301);
and U25273 (N_25273,N_24773,N_24063);
nor U25274 (N_25274,N_24663,N_24922);
and U25275 (N_25275,N_24436,N_24060);
nor U25276 (N_25276,N_24141,N_24296);
and U25277 (N_25277,N_24499,N_24303);
xor U25278 (N_25278,N_24591,N_24416);
nor U25279 (N_25279,N_24144,N_24834);
nand U25280 (N_25280,N_24315,N_24582);
xor U25281 (N_25281,N_24926,N_24557);
and U25282 (N_25282,N_24190,N_24323);
or U25283 (N_25283,N_24065,N_24308);
and U25284 (N_25284,N_24763,N_24706);
nand U25285 (N_25285,N_24917,N_24875);
or U25286 (N_25286,N_24128,N_24115);
xnor U25287 (N_25287,N_24349,N_24822);
nand U25288 (N_25288,N_24516,N_24767);
nand U25289 (N_25289,N_24652,N_24324);
nor U25290 (N_25290,N_24047,N_24535);
or U25291 (N_25291,N_24515,N_24647);
nand U25292 (N_25292,N_24046,N_24565);
xnor U25293 (N_25293,N_24072,N_24602);
or U25294 (N_25294,N_24667,N_24135);
nor U25295 (N_25295,N_24534,N_24192);
xnor U25296 (N_25296,N_24566,N_24286);
and U25297 (N_25297,N_24016,N_24843);
xnor U25298 (N_25298,N_24627,N_24776);
nand U25299 (N_25299,N_24687,N_24215);
nand U25300 (N_25300,N_24320,N_24774);
or U25301 (N_25301,N_24376,N_24904);
xor U25302 (N_25302,N_24228,N_24894);
xnor U25303 (N_25303,N_24313,N_24034);
and U25304 (N_25304,N_24965,N_24474);
nand U25305 (N_25305,N_24632,N_24014);
nor U25306 (N_25306,N_24920,N_24800);
and U25307 (N_25307,N_24035,N_24762);
or U25308 (N_25308,N_24977,N_24374);
or U25309 (N_25309,N_24239,N_24143);
and U25310 (N_25310,N_24174,N_24885);
xor U25311 (N_25311,N_24271,N_24623);
and U25312 (N_25312,N_24134,N_24985);
nand U25313 (N_25313,N_24805,N_24587);
nand U25314 (N_25314,N_24427,N_24874);
and U25315 (N_25315,N_24804,N_24829);
and U25316 (N_25316,N_24359,N_24018);
and U25317 (N_25317,N_24886,N_24787);
or U25318 (N_25318,N_24021,N_24069);
nand U25319 (N_25319,N_24712,N_24569);
nand U25320 (N_25320,N_24449,N_24929);
nor U25321 (N_25321,N_24907,N_24677);
nor U25322 (N_25322,N_24205,N_24673);
xor U25323 (N_25323,N_24497,N_24383);
and U25324 (N_25324,N_24864,N_24370);
and U25325 (N_25325,N_24783,N_24823);
or U25326 (N_25326,N_24305,N_24769);
nor U25327 (N_25327,N_24856,N_24298);
or U25328 (N_25328,N_24453,N_24756);
nand U25329 (N_25329,N_24227,N_24246);
nor U25330 (N_25330,N_24594,N_24149);
or U25331 (N_25331,N_24475,N_24732);
nor U25332 (N_25332,N_24360,N_24247);
xor U25333 (N_25333,N_24656,N_24486);
nor U25334 (N_25334,N_24281,N_24572);
or U25335 (N_25335,N_24265,N_24742);
or U25336 (N_25336,N_24352,N_24158);
nand U25337 (N_25337,N_24517,N_24655);
nand U25338 (N_25338,N_24395,N_24029);
nor U25339 (N_25339,N_24196,N_24974);
and U25340 (N_25340,N_24089,N_24770);
nand U25341 (N_25341,N_24743,N_24761);
and U25342 (N_25342,N_24912,N_24077);
nor U25343 (N_25343,N_24442,N_24871);
nand U25344 (N_25344,N_24217,N_24355);
and U25345 (N_25345,N_24382,N_24007);
and U25346 (N_25346,N_24764,N_24490);
nand U25347 (N_25347,N_24944,N_24525);
xor U25348 (N_25348,N_24645,N_24506);
nor U25349 (N_25349,N_24789,N_24277);
nor U25350 (N_25350,N_24686,N_24393);
xor U25351 (N_25351,N_24491,N_24705);
nor U25352 (N_25352,N_24954,N_24024);
xnor U25353 (N_25353,N_24580,N_24420);
and U25354 (N_25354,N_24644,N_24413);
and U25355 (N_25355,N_24451,N_24620);
or U25356 (N_25356,N_24509,N_24463);
nor U25357 (N_25357,N_24765,N_24544);
or U25358 (N_25358,N_24811,N_24057);
and U25359 (N_25359,N_24172,N_24150);
xnor U25360 (N_25360,N_24084,N_24292);
and U25361 (N_25361,N_24426,N_24610);
or U25362 (N_25362,N_24542,N_24241);
nor U25363 (N_25363,N_24167,N_24633);
nand U25364 (N_25364,N_24708,N_24526);
xor U25365 (N_25365,N_24295,N_24291);
nand U25366 (N_25366,N_24970,N_24183);
nor U25367 (N_25367,N_24543,N_24405);
nor U25368 (N_25368,N_24896,N_24105);
nor U25369 (N_25369,N_24096,N_24979);
xor U25370 (N_25370,N_24573,N_24862);
or U25371 (N_25371,N_24326,N_24471);
nor U25372 (N_25372,N_24492,N_24528);
or U25373 (N_25373,N_24868,N_24044);
or U25374 (N_25374,N_24466,N_24720);
nand U25375 (N_25375,N_24335,N_24700);
or U25376 (N_25376,N_24166,N_24054);
nor U25377 (N_25377,N_24164,N_24545);
nor U25378 (N_25378,N_24986,N_24612);
nor U25379 (N_25379,N_24396,N_24618);
and U25380 (N_25380,N_24350,N_24079);
or U25381 (N_25381,N_24696,N_24505);
nand U25382 (N_25382,N_24443,N_24242);
and U25383 (N_25383,N_24579,N_24357);
xnor U25384 (N_25384,N_24502,N_24439);
or U25385 (N_25385,N_24026,N_24575);
nor U25386 (N_25386,N_24988,N_24950);
nand U25387 (N_25387,N_24075,N_24558);
nor U25388 (N_25388,N_24211,N_24539);
xor U25389 (N_25389,N_24314,N_24733);
nand U25390 (N_25390,N_24768,N_24637);
nand U25391 (N_25391,N_24258,N_24235);
nor U25392 (N_25392,N_24777,N_24329);
or U25393 (N_25393,N_24692,N_24165);
or U25394 (N_25394,N_24759,N_24968);
or U25395 (N_25395,N_24187,N_24309);
nand U25396 (N_25396,N_24640,N_24191);
and U25397 (N_25397,N_24997,N_24472);
nor U25398 (N_25398,N_24650,N_24111);
xnor U25399 (N_25399,N_24055,N_24601);
nand U25400 (N_25400,N_24341,N_24130);
and U25401 (N_25401,N_24127,N_24550);
or U25402 (N_25402,N_24098,N_24816);
and U25403 (N_25403,N_24721,N_24554);
xnor U25404 (N_25404,N_24500,N_24312);
or U25405 (N_25405,N_24678,N_24945);
nor U25406 (N_25406,N_24270,N_24824);
or U25407 (N_25407,N_24995,N_24372);
nor U25408 (N_25408,N_24481,N_24909);
and U25409 (N_25409,N_24179,N_24597);
nand U25410 (N_25410,N_24849,N_24672);
or U25411 (N_25411,N_24794,N_24012);
nor U25412 (N_25412,N_24169,N_24848);
xor U25413 (N_25413,N_24680,N_24351);
and U25414 (N_25414,N_24325,N_24122);
and U25415 (N_25415,N_24106,N_24145);
or U25416 (N_25416,N_24336,N_24074);
nor U25417 (N_25417,N_24758,N_24212);
xor U25418 (N_25418,N_24588,N_24734);
xor U25419 (N_25419,N_24956,N_24754);
and U25420 (N_25420,N_24168,N_24961);
nand U25421 (N_25421,N_24643,N_24417);
xnor U25422 (N_25422,N_24181,N_24846);
nor U25423 (N_25423,N_24617,N_24751);
and U25424 (N_25424,N_24513,N_24469);
nor U25425 (N_25425,N_24983,N_24654);
nor U25426 (N_25426,N_24153,N_24790);
nor U25427 (N_25427,N_24792,N_24694);
nor U25428 (N_25428,N_24651,N_24447);
and U25429 (N_25429,N_24892,N_24581);
xnor U25430 (N_25430,N_24718,N_24895);
xor U25431 (N_25431,N_24615,N_24869);
nor U25432 (N_25432,N_24019,N_24741);
nor U25433 (N_25433,N_24510,N_24592);
xnor U25434 (N_25434,N_24975,N_24993);
nor U25435 (N_25435,N_24389,N_24586);
nand U25436 (N_25436,N_24508,N_24093);
or U25437 (N_25437,N_24749,N_24635);
nor U25438 (N_25438,N_24267,N_24832);
nand U25439 (N_25439,N_24980,N_24578);
nand U25440 (N_25440,N_24845,N_24541);
or U25441 (N_25441,N_24402,N_24081);
xnor U25442 (N_25442,N_24377,N_24902);
nand U25443 (N_25443,N_24722,N_24112);
or U25444 (N_25444,N_24873,N_24685);
nor U25445 (N_25445,N_24369,N_24882);
or U25446 (N_25446,N_24737,N_24998);
or U25447 (N_25447,N_24339,N_24432);
nand U25448 (N_25448,N_24739,N_24608);
or U25449 (N_25449,N_24606,N_24102);
xnor U25450 (N_25450,N_24378,N_24039);
and U25451 (N_25451,N_24299,N_24821);
nor U25452 (N_25452,N_24263,N_24855);
xor U25453 (N_25453,N_24245,N_24368);
nand U25454 (N_25454,N_24421,N_24110);
nand U25455 (N_25455,N_24365,N_24952);
nor U25456 (N_25456,N_24198,N_24552);
nand U25457 (N_25457,N_24114,N_24593);
xnor U25458 (N_25458,N_24225,N_24785);
nor U25459 (N_25459,N_24327,N_24082);
nor U25460 (N_25460,N_24715,N_24441);
xnor U25461 (N_25461,N_24042,N_24825);
nand U25462 (N_25462,N_24256,N_24076);
or U25463 (N_25463,N_24889,N_24691);
nor U25464 (N_25464,N_24170,N_24199);
nor U25465 (N_25465,N_24136,N_24186);
and U25466 (N_25466,N_24418,N_24033);
or U25467 (N_25467,N_24897,N_24109);
xnor U25468 (N_25468,N_24129,N_24480);
and U25469 (N_25469,N_24478,N_24806);
and U25470 (N_25470,N_24996,N_24923);
nor U25471 (N_25471,N_24729,N_24231);
xnor U25472 (N_25472,N_24852,N_24468);
nor U25473 (N_25473,N_24138,N_24817);
or U25474 (N_25474,N_24232,N_24719);
nand U25475 (N_25475,N_24218,N_24958);
and U25476 (N_25476,N_24001,N_24438);
xor U25477 (N_25477,N_24406,N_24530);
and U25478 (N_25478,N_24091,N_24666);
or U25479 (N_25479,N_24101,N_24450);
or U25480 (N_25480,N_24523,N_24053);
and U25481 (N_25481,N_24156,N_24844);
xor U25482 (N_25482,N_24585,N_24584);
nor U25483 (N_25483,N_24423,N_24386);
and U25484 (N_25484,N_24847,N_24603);
or U25485 (N_25485,N_24332,N_24159);
and U25486 (N_25486,N_24487,N_24595);
nor U25487 (N_25487,N_24553,N_24461);
or U25488 (N_25488,N_24624,N_24229);
or U25489 (N_25489,N_24264,N_24031);
nor U25490 (N_25490,N_24969,N_24025);
nand U25491 (N_25491,N_24863,N_24099);
nand U25492 (N_25492,N_24000,N_24730);
nor U25493 (N_25493,N_24936,N_24810);
or U25494 (N_25494,N_24630,N_24163);
and U25495 (N_25495,N_24409,N_24049);
nand U25496 (N_25496,N_24251,N_24567);
or U25497 (N_25497,N_24328,N_24254);
nand U25498 (N_25498,N_24991,N_24568);
xor U25499 (N_25499,N_24942,N_24013);
nor U25500 (N_25500,N_24445,N_24498);
nand U25501 (N_25501,N_24492,N_24273);
or U25502 (N_25502,N_24557,N_24116);
and U25503 (N_25503,N_24666,N_24184);
nor U25504 (N_25504,N_24682,N_24341);
nor U25505 (N_25505,N_24218,N_24733);
nor U25506 (N_25506,N_24138,N_24010);
xor U25507 (N_25507,N_24937,N_24393);
nor U25508 (N_25508,N_24179,N_24067);
and U25509 (N_25509,N_24470,N_24644);
nor U25510 (N_25510,N_24688,N_24835);
xnor U25511 (N_25511,N_24389,N_24528);
nor U25512 (N_25512,N_24722,N_24977);
or U25513 (N_25513,N_24353,N_24726);
nor U25514 (N_25514,N_24635,N_24399);
or U25515 (N_25515,N_24226,N_24813);
xor U25516 (N_25516,N_24240,N_24701);
xor U25517 (N_25517,N_24420,N_24016);
or U25518 (N_25518,N_24341,N_24541);
nor U25519 (N_25519,N_24506,N_24515);
xnor U25520 (N_25520,N_24119,N_24557);
nor U25521 (N_25521,N_24607,N_24485);
or U25522 (N_25522,N_24615,N_24589);
or U25523 (N_25523,N_24170,N_24897);
and U25524 (N_25524,N_24473,N_24840);
or U25525 (N_25525,N_24927,N_24364);
or U25526 (N_25526,N_24666,N_24984);
xor U25527 (N_25527,N_24110,N_24303);
or U25528 (N_25528,N_24162,N_24469);
or U25529 (N_25529,N_24431,N_24376);
or U25530 (N_25530,N_24697,N_24792);
or U25531 (N_25531,N_24407,N_24222);
nand U25532 (N_25532,N_24687,N_24840);
and U25533 (N_25533,N_24641,N_24782);
or U25534 (N_25534,N_24353,N_24082);
and U25535 (N_25535,N_24300,N_24183);
or U25536 (N_25536,N_24373,N_24273);
and U25537 (N_25537,N_24399,N_24276);
xor U25538 (N_25538,N_24829,N_24542);
xnor U25539 (N_25539,N_24738,N_24147);
nor U25540 (N_25540,N_24517,N_24234);
xor U25541 (N_25541,N_24572,N_24765);
nor U25542 (N_25542,N_24953,N_24074);
xor U25543 (N_25543,N_24620,N_24447);
nor U25544 (N_25544,N_24225,N_24839);
nand U25545 (N_25545,N_24013,N_24312);
xnor U25546 (N_25546,N_24657,N_24237);
xor U25547 (N_25547,N_24179,N_24546);
nand U25548 (N_25548,N_24616,N_24486);
nor U25549 (N_25549,N_24038,N_24638);
and U25550 (N_25550,N_24084,N_24737);
nand U25551 (N_25551,N_24459,N_24055);
nand U25552 (N_25552,N_24072,N_24062);
nor U25553 (N_25553,N_24030,N_24823);
nand U25554 (N_25554,N_24170,N_24172);
nand U25555 (N_25555,N_24674,N_24379);
xor U25556 (N_25556,N_24341,N_24756);
nor U25557 (N_25557,N_24140,N_24554);
nor U25558 (N_25558,N_24519,N_24523);
and U25559 (N_25559,N_24078,N_24991);
or U25560 (N_25560,N_24186,N_24662);
and U25561 (N_25561,N_24419,N_24981);
or U25562 (N_25562,N_24951,N_24501);
and U25563 (N_25563,N_24203,N_24123);
nand U25564 (N_25564,N_24876,N_24136);
xnor U25565 (N_25565,N_24845,N_24130);
and U25566 (N_25566,N_24019,N_24127);
xnor U25567 (N_25567,N_24585,N_24721);
nor U25568 (N_25568,N_24777,N_24105);
nand U25569 (N_25569,N_24849,N_24697);
xnor U25570 (N_25570,N_24487,N_24922);
nor U25571 (N_25571,N_24663,N_24492);
nor U25572 (N_25572,N_24435,N_24103);
nor U25573 (N_25573,N_24649,N_24015);
nor U25574 (N_25574,N_24309,N_24147);
and U25575 (N_25575,N_24875,N_24829);
nand U25576 (N_25576,N_24168,N_24481);
nand U25577 (N_25577,N_24489,N_24411);
or U25578 (N_25578,N_24859,N_24824);
and U25579 (N_25579,N_24066,N_24821);
and U25580 (N_25580,N_24641,N_24767);
xor U25581 (N_25581,N_24309,N_24828);
nand U25582 (N_25582,N_24531,N_24383);
or U25583 (N_25583,N_24217,N_24318);
nor U25584 (N_25584,N_24232,N_24809);
and U25585 (N_25585,N_24383,N_24382);
nor U25586 (N_25586,N_24721,N_24124);
nand U25587 (N_25587,N_24831,N_24364);
and U25588 (N_25588,N_24250,N_24890);
nand U25589 (N_25589,N_24749,N_24846);
and U25590 (N_25590,N_24330,N_24319);
and U25591 (N_25591,N_24706,N_24392);
or U25592 (N_25592,N_24130,N_24796);
nor U25593 (N_25593,N_24865,N_24870);
or U25594 (N_25594,N_24484,N_24767);
or U25595 (N_25595,N_24703,N_24257);
or U25596 (N_25596,N_24447,N_24863);
nor U25597 (N_25597,N_24723,N_24188);
nand U25598 (N_25598,N_24932,N_24757);
or U25599 (N_25599,N_24826,N_24543);
nand U25600 (N_25600,N_24004,N_24530);
xor U25601 (N_25601,N_24801,N_24525);
and U25602 (N_25602,N_24229,N_24641);
nand U25603 (N_25603,N_24721,N_24331);
or U25604 (N_25604,N_24789,N_24253);
nand U25605 (N_25605,N_24081,N_24371);
nor U25606 (N_25606,N_24787,N_24699);
or U25607 (N_25607,N_24316,N_24309);
nand U25608 (N_25608,N_24835,N_24398);
xor U25609 (N_25609,N_24168,N_24076);
nand U25610 (N_25610,N_24459,N_24649);
or U25611 (N_25611,N_24109,N_24586);
or U25612 (N_25612,N_24325,N_24918);
nor U25613 (N_25613,N_24326,N_24797);
xor U25614 (N_25614,N_24661,N_24138);
xor U25615 (N_25615,N_24108,N_24703);
xnor U25616 (N_25616,N_24911,N_24812);
xor U25617 (N_25617,N_24972,N_24962);
xnor U25618 (N_25618,N_24814,N_24301);
xnor U25619 (N_25619,N_24481,N_24043);
or U25620 (N_25620,N_24511,N_24872);
or U25621 (N_25621,N_24917,N_24354);
xor U25622 (N_25622,N_24401,N_24002);
and U25623 (N_25623,N_24393,N_24262);
nand U25624 (N_25624,N_24188,N_24520);
and U25625 (N_25625,N_24304,N_24432);
xnor U25626 (N_25626,N_24627,N_24369);
or U25627 (N_25627,N_24133,N_24328);
nand U25628 (N_25628,N_24808,N_24601);
or U25629 (N_25629,N_24592,N_24359);
or U25630 (N_25630,N_24237,N_24652);
nand U25631 (N_25631,N_24438,N_24317);
xnor U25632 (N_25632,N_24772,N_24481);
or U25633 (N_25633,N_24772,N_24474);
and U25634 (N_25634,N_24174,N_24638);
nand U25635 (N_25635,N_24501,N_24066);
nand U25636 (N_25636,N_24951,N_24273);
nor U25637 (N_25637,N_24651,N_24086);
nor U25638 (N_25638,N_24495,N_24261);
xor U25639 (N_25639,N_24401,N_24391);
nand U25640 (N_25640,N_24457,N_24360);
nor U25641 (N_25641,N_24239,N_24707);
and U25642 (N_25642,N_24200,N_24292);
xor U25643 (N_25643,N_24811,N_24111);
nand U25644 (N_25644,N_24409,N_24820);
or U25645 (N_25645,N_24990,N_24740);
and U25646 (N_25646,N_24878,N_24931);
and U25647 (N_25647,N_24909,N_24876);
xor U25648 (N_25648,N_24500,N_24564);
nand U25649 (N_25649,N_24106,N_24163);
nand U25650 (N_25650,N_24613,N_24624);
nand U25651 (N_25651,N_24505,N_24634);
nand U25652 (N_25652,N_24749,N_24796);
nand U25653 (N_25653,N_24386,N_24629);
nor U25654 (N_25654,N_24944,N_24360);
nand U25655 (N_25655,N_24343,N_24062);
nor U25656 (N_25656,N_24022,N_24892);
nor U25657 (N_25657,N_24670,N_24203);
or U25658 (N_25658,N_24129,N_24021);
nand U25659 (N_25659,N_24232,N_24931);
and U25660 (N_25660,N_24416,N_24901);
xnor U25661 (N_25661,N_24950,N_24803);
nor U25662 (N_25662,N_24607,N_24302);
and U25663 (N_25663,N_24690,N_24853);
nor U25664 (N_25664,N_24872,N_24915);
and U25665 (N_25665,N_24376,N_24776);
and U25666 (N_25666,N_24038,N_24307);
and U25667 (N_25667,N_24808,N_24479);
or U25668 (N_25668,N_24911,N_24225);
nand U25669 (N_25669,N_24548,N_24564);
and U25670 (N_25670,N_24362,N_24750);
nand U25671 (N_25671,N_24658,N_24278);
xor U25672 (N_25672,N_24475,N_24768);
xor U25673 (N_25673,N_24077,N_24148);
nor U25674 (N_25674,N_24390,N_24942);
and U25675 (N_25675,N_24241,N_24685);
or U25676 (N_25676,N_24121,N_24111);
or U25677 (N_25677,N_24885,N_24953);
or U25678 (N_25678,N_24282,N_24083);
or U25679 (N_25679,N_24575,N_24539);
nor U25680 (N_25680,N_24437,N_24279);
and U25681 (N_25681,N_24535,N_24734);
nand U25682 (N_25682,N_24086,N_24461);
nand U25683 (N_25683,N_24378,N_24943);
xnor U25684 (N_25684,N_24738,N_24142);
and U25685 (N_25685,N_24868,N_24828);
xnor U25686 (N_25686,N_24359,N_24155);
xnor U25687 (N_25687,N_24009,N_24564);
xnor U25688 (N_25688,N_24469,N_24391);
xnor U25689 (N_25689,N_24852,N_24174);
xnor U25690 (N_25690,N_24829,N_24785);
xnor U25691 (N_25691,N_24075,N_24529);
and U25692 (N_25692,N_24115,N_24813);
or U25693 (N_25693,N_24844,N_24148);
nor U25694 (N_25694,N_24661,N_24854);
nor U25695 (N_25695,N_24319,N_24883);
nor U25696 (N_25696,N_24330,N_24719);
nor U25697 (N_25697,N_24741,N_24626);
or U25698 (N_25698,N_24809,N_24374);
nor U25699 (N_25699,N_24401,N_24981);
xnor U25700 (N_25700,N_24326,N_24651);
and U25701 (N_25701,N_24812,N_24225);
nand U25702 (N_25702,N_24378,N_24577);
and U25703 (N_25703,N_24175,N_24551);
and U25704 (N_25704,N_24379,N_24904);
nand U25705 (N_25705,N_24705,N_24227);
xor U25706 (N_25706,N_24455,N_24342);
nor U25707 (N_25707,N_24757,N_24949);
xnor U25708 (N_25708,N_24544,N_24392);
xor U25709 (N_25709,N_24220,N_24150);
nand U25710 (N_25710,N_24295,N_24283);
nor U25711 (N_25711,N_24215,N_24720);
and U25712 (N_25712,N_24073,N_24637);
nand U25713 (N_25713,N_24971,N_24009);
or U25714 (N_25714,N_24509,N_24189);
nand U25715 (N_25715,N_24845,N_24204);
xnor U25716 (N_25716,N_24405,N_24362);
nor U25717 (N_25717,N_24597,N_24486);
and U25718 (N_25718,N_24724,N_24457);
or U25719 (N_25719,N_24803,N_24926);
xnor U25720 (N_25720,N_24017,N_24912);
or U25721 (N_25721,N_24989,N_24628);
nand U25722 (N_25722,N_24454,N_24955);
nand U25723 (N_25723,N_24993,N_24205);
xnor U25724 (N_25724,N_24364,N_24922);
or U25725 (N_25725,N_24636,N_24056);
nand U25726 (N_25726,N_24196,N_24916);
or U25727 (N_25727,N_24950,N_24349);
nor U25728 (N_25728,N_24676,N_24842);
nor U25729 (N_25729,N_24369,N_24648);
nor U25730 (N_25730,N_24459,N_24300);
xnor U25731 (N_25731,N_24977,N_24913);
xor U25732 (N_25732,N_24981,N_24662);
or U25733 (N_25733,N_24562,N_24178);
and U25734 (N_25734,N_24255,N_24406);
or U25735 (N_25735,N_24937,N_24206);
nor U25736 (N_25736,N_24778,N_24102);
nor U25737 (N_25737,N_24708,N_24505);
xnor U25738 (N_25738,N_24606,N_24084);
nor U25739 (N_25739,N_24487,N_24813);
nand U25740 (N_25740,N_24003,N_24485);
nand U25741 (N_25741,N_24956,N_24304);
xor U25742 (N_25742,N_24575,N_24284);
and U25743 (N_25743,N_24045,N_24095);
xor U25744 (N_25744,N_24715,N_24775);
and U25745 (N_25745,N_24805,N_24323);
or U25746 (N_25746,N_24179,N_24480);
or U25747 (N_25747,N_24682,N_24843);
xor U25748 (N_25748,N_24570,N_24535);
or U25749 (N_25749,N_24010,N_24410);
or U25750 (N_25750,N_24099,N_24445);
nor U25751 (N_25751,N_24301,N_24204);
nor U25752 (N_25752,N_24514,N_24340);
nor U25753 (N_25753,N_24300,N_24570);
xor U25754 (N_25754,N_24624,N_24433);
and U25755 (N_25755,N_24078,N_24585);
nand U25756 (N_25756,N_24924,N_24334);
nor U25757 (N_25757,N_24684,N_24475);
xnor U25758 (N_25758,N_24710,N_24586);
and U25759 (N_25759,N_24576,N_24533);
and U25760 (N_25760,N_24416,N_24015);
and U25761 (N_25761,N_24626,N_24507);
or U25762 (N_25762,N_24114,N_24643);
nand U25763 (N_25763,N_24057,N_24841);
nand U25764 (N_25764,N_24130,N_24318);
or U25765 (N_25765,N_24771,N_24979);
nor U25766 (N_25766,N_24609,N_24196);
xor U25767 (N_25767,N_24117,N_24594);
nand U25768 (N_25768,N_24330,N_24463);
nand U25769 (N_25769,N_24127,N_24248);
nand U25770 (N_25770,N_24294,N_24049);
and U25771 (N_25771,N_24878,N_24548);
nand U25772 (N_25772,N_24685,N_24957);
or U25773 (N_25773,N_24172,N_24183);
nor U25774 (N_25774,N_24723,N_24877);
nand U25775 (N_25775,N_24206,N_24550);
or U25776 (N_25776,N_24962,N_24516);
xor U25777 (N_25777,N_24966,N_24262);
nand U25778 (N_25778,N_24540,N_24954);
nand U25779 (N_25779,N_24746,N_24924);
nand U25780 (N_25780,N_24903,N_24880);
nor U25781 (N_25781,N_24006,N_24064);
xor U25782 (N_25782,N_24487,N_24623);
nand U25783 (N_25783,N_24467,N_24198);
xnor U25784 (N_25784,N_24101,N_24996);
or U25785 (N_25785,N_24202,N_24270);
nand U25786 (N_25786,N_24539,N_24364);
xor U25787 (N_25787,N_24775,N_24709);
nor U25788 (N_25788,N_24162,N_24892);
xnor U25789 (N_25789,N_24640,N_24498);
or U25790 (N_25790,N_24258,N_24435);
or U25791 (N_25791,N_24464,N_24150);
or U25792 (N_25792,N_24072,N_24143);
xor U25793 (N_25793,N_24372,N_24721);
nand U25794 (N_25794,N_24355,N_24232);
and U25795 (N_25795,N_24630,N_24351);
nand U25796 (N_25796,N_24815,N_24687);
and U25797 (N_25797,N_24360,N_24037);
and U25798 (N_25798,N_24564,N_24561);
or U25799 (N_25799,N_24245,N_24680);
nand U25800 (N_25800,N_24988,N_24532);
and U25801 (N_25801,N_24352,N_24879);
nand U25802 (N_25802,N_24838,N_24663);
or U25803 (N_25803,N_24893,N_24304);
nand U25804 (N_25804,N_24981,N_24128);
and U25805 (N_25805,N_24259,N_24097);
and U25806 (N_25806,N_24980,N_24620);
nor U25807 (N_25807,N_24794,N_24390);
and U25808 (N_25808,N_24930,N_24286);
and U25809 (N_25809,N_24369,N_24875);
nand U25810 (N_25810,N_24342,N_24079);
nor U25811 (N_25811,N_24799,N_24849);
nor U25812 (N_25812,N_24970,N_24367);
xor U25813 (N_25813,N_24489,N_24100);
nor U25814 (N_25814,N_24728,N_24680);
xor U25815 (N_25815,N_24410,N_24642);
nor U25816 (N_25816,N_24138,N_24439);
and U25817 (N_25817,N_24018,N_24834);
nand U25818 (N_25818,N_24033,N_24809);
nor U25819 (N_25819,N_24767,N_24747);
and U25820 (N_25820,N_24664,N_24873);
nor U25821 (N_25821,N_24151,N_24767);
nand U25822 (N_25822,N_24178,N_24714);
or U25823 (N_25823,N_24739,N_24849);
nor U25824 (N_25824,N_24430,N_24648);
and U25825 (N_25825,N_24519,N_24200);
and U25826 (N_25826,N_24464,N_24298);
nand U25827 (N_25827,N_24144,N_24556);
and U25828 (N_25828,N_24539,N_24793);
nand U25829 (N_25829,N_24015,N_24851);
nand U25830 (N_25830,N_24692,N_24302);
or U25831 (N_25831,N_24845,N_24446);
xor U25832 (N_25832,N_24806,N_24573);
xor U25833 (N_25833,N_24735,N_24057);
or U25834 (N_25834,N_24297,N_24559);
and U25835 (N_25835,N_24890,N_24866);
nand U25836 (N_25836,N_24123,N_24576);
or U25837 (N_25837,N_24634,N_24965);
nor U25838 (N_25838,N_24375,N_24924);
xnor U25839 (N_25839,N_24911,N_24712);
nor U25840 (N_25840,N_24725,N_24517);
nor U25841 (N_25841,N_24540,N_24414);
xor U25842 (N_25842,N_24018,N_24151);
nand U25843 (N_25843,N_24106,N_24395);
or U25844 (N_25844,N_24771,N_24695);
and U25845 (N_25845,N_24604,N_24112);
xor U25846 (N_25846,N_24028,N_24616);
nand U25847 (N_25847,N_24348,N_24783);
and U25848 (N_25848,N_24678,N_24476);
xnor U25849 (N_25849,N_24328,N_24572);
nor U25850 (N_25850,N_24011,N_24105);
xnor U25851 (N_25851,N_24729,N_24978);
or U25852 (N_25852,N_24510,N_24974);
nand U25853 (N_25853,N_24971,N_24713);
nand U25854 (N_25854,N_24306,N_24358);
and U25855 (N_25855,N_24835,N_24261);
and U25856 (N_25856,N_24718,N_24949);
or U25857 (N_25857,N_24857,N_24576);
nor U25858 (N_25858,N_24385,N_24752);
nor U25859 (N_25859,N_24182,N_24228);
xor U25860 (N_25860,N_24913,N_24495);
xor U25861 (N_25861,N_24735,N_24081);
nand U25862 (N_25862,N_24587,N_24686);
nor U25863 (N_25863,N_24722,N_24885);
xnor U25864 (N_25864,N_24680,N_24175);
nand U25865 (N_25865,N_24017,N_24574);
or U25866 (N_25866,N_24539,N_24231);
nand U25867 (N_25867,N_24597,N_24421);
xor U25868 (N_25868,N_24548,N_24883);
xor U25869 (N_25869,N_24704,N_24461);
xor U25870 (N_25870,N_24063,N_24672);
nor U25871 (N_25871,N_24780,N_24709);
or U25872 (N_25872,N_24839,N_24070);
nand U25873 (N_25873,N_24276,N_24085);
or U25874 (N_25874,N_24991,N_24607);
and U25875 (N_25875,N_24152,N_24236);
xnor U25876 (N_25876,N_24946,N_24004);
or U25877 (N_25877,N_24147,N_24671);
nand U25878 (N_25878,N_24163,N_24236);
nand U25879 (N_25879,N_24861,N_24876);
xnor U25880 (N_25880,N_24208,N_24998);
and U25881 (N_25881,N_24237,N_24738);
xor U25882 (N_25882,N_24939,N_24076);
and U25883 (N_25883,N_24595,N_24861);
or U25884 (N_25884,N_24375,N_24142);
xnor U25885 (N_25885,N_24317,N_24923);
or U25886 (N_25886,N_24686,N_24649);
nor U25887 (N_25887,N_24729,N_24010);
xor U25888 (N_25888,N_24049,N_24899);
or U25889 (N_25889,N_24435,N_24544);
or U25890 (N_25890,N_24284,N_24883);
nor U25891 (N_25891,N_24121,N_24139);
nor U25892 (N_25892,N_24615,N_24926);
xor U25893 (N_25893,N_24154,N_24894);
nand U25894 (N_25894,N_24824,N_24437);
nand U25895 (N_25895,N_24181,N_24765);
and U25896 (N_25896,N_24639,N_24148);
xnor U25897 (N_25897,N_24916,N_24764);
nor U25898 (N_25898,N_24752,N_24659);
nand U25899 (N_25899,N_24337,N_24755);
nor U25900 (N_25900,N_24535,N_24691);
nor U25901 (N_25901,N_24535,N_24297);
or U25902 (N_25902,N_24686,N_24222);
nand U25903 (N_25903,N_24381,N_24461);
nor U25904 (N_25904,N_24596,N_24517);
or U25905 (N_25905,N_24705,N_24203);
or U25906 (N_25906,N_24520,N_24680);
and U25907 (N_25907,N_24925,N_24583);
nand U25908 (N_25908,N_24253,N_24483);
nand U25909 (N_25909,N_24879,N_24724);
xnor U25910 (N_25910,N_24830,N_24099);
nand U25911 (N_25911,N_24683,N_24055);
or U25912 (N_25912,N_24488,N_24391);
xnor U25913 (N_25913,N_24780,N_24662);
xnor U25914 (N_25914,N_24465,N_24601);
and U25915 (N_25915,N_24826,N_24325);
nor U25916 (N_25916,N_24656,N_24491);
nor U25917 (N_25917,N_24790,N_24774);
nor U25918 (N_25918,N_24857,N_24922);
and U25919 (N_25919,N_24447,N_24134);
nand U25920 (N_25920,N_24073,N_24576);
xor U25921 (N_25921,N_24612,N_24357);
xnor U25922 (N_25922,N_24639,N_24532);
and U25923 (N_25923,N_24086,N_24720);
or U25924 (N_25924,N_24645,N_24823);
or U25925 (N_25925,N_24714,N_24559);
xnor U25926 (N_25926,N_24716,N_24200);
xor U25927 (N_25927,N_24827,N_24630);
or U25928 (N_25928,N_24798,N_24102);
and U25929 (N_25929,N_24709,N_24559);
nor U25930 (N_25930,N_24241,N_24607);
nand U25931 (N_25931,N_24765,N_24828);
and U25932 (N_25932,N_24718,N_24424);
or U25933 (N_25933,N_24788,N_24364);
nor U25934 (N_25934,N_24351,N_24531);
nor U25935 (N_25935,N_24797,N_24089);
or U25936 (N_25936,N_24953,N_24517);
xnor U25937 (N_25937,N_24148,N_24346);
or U25938 (N_25938,N_24923,N_24373);
nand U25939 (N_25939,N_24795,N_24040);
nor U25940 (N_25940,N_24628,N_24663);
or U25941 (N_25941,N_24447,N_24322);
and U25942 (N_25942,N_24389,N_24143);
and U25943 (N_25943,N_24310,N_24235);
or U25944 (N_25944,N_24220,N_24012);
and U25945 (N_25945,N_24637,N_24931);
and U25946 (N_25946,N_24685,N_24460);
nor U25947 (N_25947,N_24532,N_24187);
nor U25948 (N_25948,N_24606,N_24386);
xor U25949 (N_25949,N_24366,N_24869);
nor U25950 (N_25950,N_24813,N_24024);
nor U25951 (N_25951,N_24406,N_24597);
xor U25952 (N_25952,N_24497,N_24636);
nor U25953 (N_25953,N_24859,N_24484);
and U25954 (N_25954,N_24728,N_24899);
nor U25955 (N_25955,N_24208,N_24638);
and U25956 (N_25956,N_24204,N_24989);
or U25957 (N_25957,N_24657,N_24624);
xor U25958 (N_25958,N_24016,N_24492);
nand U25959 (N_25959,N_24031,N_24929);
or U25960 (N_25960,N_24735,N_24460);
or U25961 (N_25961,N_24314,N_24703);
and U25962 (N_25962,N_24163,N_24871);
xnor U25963 (N_25963,N_24598,N_24351);
nand U25964 (N_25964,N_24712,N_24164);
xor U25965 (N_25965,N_24727,N_24211);
and U25966 (N_25966,N_24902,N_24199);
and U25967 (N_25967,N_24588,N_24062);
nor U25968 (N_25968,N_24754,N_24268);
or U25969 (N_25969,N_24844,N_24894);
and U25970 (N_25970,N_24289,N_24404);
nor U25971 (N_25971,N_24379,N_24877);
and U25972 (N_25972,N_24631,N_24321);
nand U25973 (N_25973,N_24954,N_24812);
and U25974 (N_25974,N_24618,N_24622);
xnor U25975 (N_25975,N_24596,N_24563);
nor U25976 (N_25976,N_24200,N_24123);
nand U25977 (N_25977,N_24512,N_24528);
nor U25978 (N_25978,N_24458,N_24335);
and U25979 (N_25979,N_24467,N_24424);
and U25980 (N_25980,N_24829,N_24989);
xor U25981 (N_25981,N_24725,N_24553);
and U25982 (N_25982,N_24441,N_24308);
nor U25983 (N_25983,N_24475,N_24738);
and U25984 (N_25984,N_24941,N_24262);
xor U25985 (N_25985,N_24919,N_24191);
and U25986 (N_25986,N_24937,N_24615);
nand U25987 (N_25987,N_24034,N_24879);
nand U25988 (N_25988,N_24985,N_24593);
or U25989 (N_25989,N_24324,N_24068);
nor U25990 (N_25990,N_24858,N_24713);
or U25991 (N_25991,N_24133,N_24910);
nor U25992 (N_25992,N_24680,N_24589);
nand U25993 (N_25993,N_24786,N_24381);
nor U25994 (N_25994,N_24948,N_24572);
and U25995 (N_25995,N_24858,N_24332);
nor U25996 (N_25996,N_24787,N_24979);
or U25997 (N_25997,N_24216,N_24099);
and U25998 (N_25998,N_24722,N_24504);
nor U25999 (N_25999,N_24193,N_24013);
xor U26000 (N_26000,N_25960,N_25011);
nor U26001 (N_26001,N_25119,N_25566);
nor U26002 (N_26002,N_25242,N_25238);
or U26003 (N_26003,N_25070,N_25902);
nor U26004 (N_26004,N_25776,N_25355);
nand U26005 (N_26005,N_25321,N_25615);
nand U26006 (N_26006,N_25704,N_25648);
xor U26007 (N_26007,N_25244,N_25398);
nor U26008 (N_26008,N_25548,N_25609);
and U26009 (N_26009,N_25970,N_25120);
xnor U26010 (N_26010,N_25488,N_25212);
or U26011 (N_26011,N_25807,N_25980);
nand U26012 (N_26012,N_25599,N_25264);
xor U26013 (N_26013,N_25876,N_25809);
or U26014 (N_26014,N_25605,N_25381);
xnor U26015 (N_26015,N_25383,N_25183);
or U26016 (N_26016,N_25944,N_25639);
xor U26017 (N_26017,N_25029,N_25695);
or U26018 (N_26018,N_25565,N_25144);
nand U26019 (N_26019,N_25991,N_25797);
and U26020 (N_26020,N_25401,N_25514);
xnor U26021 (N_26021,N_25533,N_25719);
nand U26022 (N_26022,N_25554,N_25839);
and U26023 (N_26023,N_25400,N_25028);
nand U26024 (N_26024,N_25095,N_25058);
or U26025 (N_26025,N_25055,N_25754);
nand U26026 (N_26026,N_25301,N_25893);
xor U26027 (N_26027,N_25252,N_25228);
and U26028 (N_26028,N_25319,N_25056);
nor U26029 (N_26029,N_25414,N_25691);
xnor U26030 (N_26030,N_25993,N_25663);
nor U26031 (N_26031,N_25077,N_25142);
or U26032 (N_26032,N_25758,N_25971);
xnor U26033 (N_26033,N_25637,N_25521);
or U26034 (N_26034,N_25715,N_25764);
or U26035 (N_26035,N_25102,N_25498);
nor U26036 (N_26036,N_25847,N_25946);
nand U26037 (N_26037,N_25898,N_25841);
nand U26038 (N_26038,N_25802,N_25277);
xnor U26039 (N_26039,N_25878,N_25812);
nor U26040 (N_26040,N_25374,N_25757);
or U26041 (N_26041,N_25517,N_25805);
nor U26042 (N_26042,N_25061,N_25240);
nand U26043 (N_26043,N_25372,N_25487);
xor U26044 (N_26044,N_25750,N_25798);
nand U26045 (N_26045,N_25771,N_25344);
xnor U26046 (N_26046,N_25849,N_25935);
or U26047 (N_26047,N_25094,N_25018);
nor U26048 (N_26048,N_25528,N_25774);
nand U26049 (N_26049,N_25207,N_25957);
or U26050 (N_26050,N_25818,N_25641);
nand U26051 (N_26051,N_25230,N_25469);
nor U26052 (N_26052,N_25112,N_25416);
and U26053 (N_26053,N_25836,N_25689);
and U26054 (N_26054,N_25138,N_25622);
nand U26055 (N_26055,N_25089,N_25241);
nand U26056 (N_26056,N_25567,N_25146);
or U26057 (N_26057,N_25200,N_25043);
or U26058 (N_26058,N_25871,N_25880);
or U26059 (N_26059,N_25668,N_25698);
nand U26060 (N_26060,N_25940,N_25642);
and U26061 (N_26061,N_25122,N_25198);
nand U26062 (N_26062,N_25678,N_25752);
nand U26063 (N_26063,N_25900,N_25889);
nand U26064 (N_26064,N_25644,N_25125);
and U26065 (N_26065,N_25779,N_25643);
xnor U26066 (N_26066,N_25101,N_25432);
and U26067 (N_26067,N_25187,N_25934);
nor U26068 (N_26068,N_25324,N_25051);
xnor U26069 (N_26069,N_25965,N_25068);
and U26070 (N_26070,N_25604,N_25938);
or U26071 (N_26071,N_25099,N_25368);
nand U26072 (N_26072,N_25652,N_25822);
or U26073 (N_26073,N_25843,N_25558);
xnor U26074 (N_26074,N_25922,N_25888);
nand U26075 (N_26075,N_25925,N_25071);
and U26076 (N_26076,N_25526,N_25306);
nand U26077 (N_26077,N_25134,N_25366);
nor U26078 (N_26078,N_25202,N_25196);
nand U26079 (N_26079,N_25979,N_25059);
and U26080 (N_26080,N_25882,N_25072);
or U26081 (N_26081,N_25015,N_25420);
xor U26082 (N_26082,N_25687,N_25740);
nor U26083 (N_26083,N_25865,N_25166);
or U26084 (N_26084,N_25515,N_25601);
nor U26085 (N_26085,N_25378,N_25586);
nor U26086 (N_26086,N_25794,N_25217);
nor U26087 (N_26087,N_25821,N_25098);
or U26088 (N_26088,N_25780,N_25547);
nand U26089 (N_26089,N_25218,N_25382);
nor U26090 (N_26090,N_25860,N_25305);
xnor U26091 (N_26091,N_25781,N_25247);
nand U26092 (N_26092,N_25271,N_25295);
nor U26093 (N_26093,N_25275,N_25943);
and U26094 (N_26094,N_25906,N_25039);
or U26095 (N_26095,N_25760,N_25429);
nand U26096 (N_26096,N_25079,N_25551);
or U26097 (N_26097,N_25158,N_25457);
nor U26098 (N_26098,N_25160,N_25103);
xor U26099 (N_26099,N_25769,N_25861);
xor U26100 (N_26100,N_25937,N_25623);
nor U26101 (N_26101,N_25872,N_25336);
and U26102 (N_26102,N_25220,N_25048);
and U26103 (N_26103,N_25359,N_25670);
nor U26104 (N_26104,N_25667,N_25694);
and U26105 (N_26105,N_25193,N_25743);
xnor U26106 (N_26106,N_25826,N_25279);
nand U26107 (N_26107,N_25507,N_25294);
and U26108 (N_26108,N_25895,N_25522);
or U26109 (N_26109,N_25097,N_25563);
xnor U26110 (N_26110,N_25360,N_25133);
nor U26111 (N_26111,N_25076,N_25789);
or U26112 (N_26112,N_25536,N_25284);
nand U26113 (N_26113,N_25140,N_25655);
nand U26114 (N_26114,N_25243,N_25427);
or U26115 (N_26115,N_25830,N_25574);
and U26116 (N_26116,N_25475,N_25621);
nand U26117 (N_26117,N_25856,N_25405);
or U26118 (N_26118,N_25185,N_25811);
and U26119 (N_26119,N_25316,N_25369);
xnor U26120 (N_26120,N_25389,N_25082);
xnor U26121 (N_26121,N_25659,N_25763);
nor U26122 (N_26122,N_25364,N_25555);
nand U26123 (N_26123,N_25920,N_25176);
xor U26124 (N_26124,N_25000,N_25025);
xnor U26125 (N_26125,N_25741,N_25542);
and U26126 (N_26126,N_25523,N_25494);
nor U26127 (N_26127,N_25292,N_25014);
or U26128 (N_26128,N_25057,N_25988);
xor U26129 (N_26129,N_25091,N_25245);
or U26130 (N_26130,N_25022,N_25788);
and U26131 (N_26131,N_25385,N_25896);
xor U26132 (N_26132,N_25041,N_25434);
nand U26133 (N_26133,N_25341,N_25145);
or U26134 (N_26134,N_25603,N_25040);
nor U26135 (N_26135,N_25147,N_25984);
or U26136 (N_26136,N_25996,N_25908);
or U26137 (N_26137,N_25869,N_25411);
or U26138 (N_26138,N_25538,N_25038);
and U26139 (N_26139,N_25393,N_25660);
nand U26140 (N_26140,N_25465,N_25339);
and U26141 (N_26141,N_25711,N_25417);
nor U26142 (N_26142,N_25897,N_25624);
nor U26143 (N_26143,N_25657,N_25249);
and U26144 (N_26144,N_25092,N_25229);
xnor U26145 (N_26145,N_25472,N_25831);
nor U26146 (N_26146,N_25474,N_25402);
or U26147 (N_26147,N_25491,N_25801);
and U26148 (N_26148,N_25253,N_25181);
xnor U26149 (N_26149,N_25458,N_25795);
nand U26150 (N_26150,N_25633,N_25701);
xnor U26151 (N_26151,N_25718,N_25783);
nand U26152 (N_26152,N_25867,N_25912);
xnor U26153 (N_26153,N_25832,N_25111);
xnor U26154 (N_26154,N_25310,N_25032);
nor U26155 (N_26155,N_25157,N_25464);
or U26156 (N_26156,N_25915,N_25325);
xnor U26157 (N_26157,N_25251,N_25917);
xor U26158 (N_26158,N_25269,N_25972);
xor U26159 (N_26159,N_25820,N_25323);
and U26160 (N_26160,N_25738,N_25167);
nand U26161 (N_26161,N_25923,N_25594);
or U26162 (N_26162,N_25118,N_25209);
or U26163 (N_26163,N_25153,N_25645);
nand U26164 (N_26164,N_25775,N_25404);
or U26165 (N_26165,N_25840,N_25449);
or U26166 (N_26166,N_25141,N_25026);
xor U26167 (N_26167,N_25328,N_25909);
xor U26168 (N_26168,N_25233,N_25737);
nor U26169 (N_26169,N_25451,N_25108);
nor U26170 (N_26170,N_25312,N_25785);
and U26171 (N_26171,N_25197,N_25685);
nor U26172 (N_26172,N_25512,N_25595);
xnor U26173 (N_26173,N_25591,N_25833);
or U26174 (N_26174,N_25213,N_25553);
nor U26175 (N_26175,N_25579,N_25280);
xnor U26176 (N_26176,N_25023,N_25858);
and U26177 (N_26177,N_25790,N_25778);
or U26178 (N_26178,N_25592,N_25390);
nand U26179 (N_26179,N_25463,N_25675);
xor U26180 (N_26180,N_25263,N_25161);
nand U26181 (N_26181,N_25356,N_25413);
nor U26182 (N_26182,N_25471,N_25438);
and U26183 (N_26183,N_25504,N_25268);
or U26184 (N_26184,N_25619,N_25851);
or U26185 (N_26185,N_25949,N_25124);
xnor U26186 (N_26186,N_25992,N_25786);
xor U26187 (N_26187,N_25215,N_25884);
nor U26188 (N_26188,N_25186,N_25274);
nor U26189 (N_26189,N_25834,N_25367);
nand U26190 (N_26190,N_25007,N_25823);
or U26191 (N_26191,N_25700,N_25005);
xor U26192 (N_26192,N_25723,N_25673);
and U26193 (N_26193,N_25501,N_25045);
nor U26194 (N_26194,N_25162,N_25201);
nor U26195 (N_26195,N_25482,N_25674);
and U26196 (N_26196,N_25583,N_25837);
or U26197 (N_26197,N_25534,N_25881);
nor U26198 (N_26198,N_25379,N_25327);
nor U26199 (N_26199,N_25531,N_25455);
nor U26200 (N_26200,N_25034,N_25762);
nand U26201 (N_26201,N_25969,N_25748);
nor U26202 (N_26202,N_25540,N_25532);
nand U26203 (N_26203,N_25496,N_25054);
xor U26204 (N_26204,N_25206,N_25165);
xnor U26205 (N_26205,N_25293,N_25721);
nand U26206 (N_26206,N_25440,N_25891);
xor U26207 (N_26207,N_25787,N_25857);
nand U26208 (N_26208,N_25707,N_25333);
nor U26209 (N_26209,N_25497,N_25191);
or U26210 (N_26210,N_25044,N_25669);
nand U26211 (N_26211,N_25903,N_25887);
and U26212 (N_26212,N_25357,N_25733);
nor U26213 (N_26213,N_25791,N_25572);
nand U26214 (N_26214,N_25924,N_25656);
xnor U26215 (N_26215,N_25964,N_25928);
or U26216 (N_26216,N_25063,N_25956);
xnor U26217 (N_26217,N_25137,N_25977);
nor U26218 (N_26218,N_25047,N_25330);
or U26219 (N_26219,N_25990,N_25478);
nor U26220 (N_26220,N_25425,N_25350);
xor U26221 (N_26221,N_25725,N_25877);
nor U26222 (N_26222,N_25329,N_25454);
nand U26223 (N_26223,N_25744,N_25428);
or U26224 (N_26224,N_25033,N_25384);
and U26225 (N_26225,N_25508,N_25998);
or U26226 (N_26226,N_25223,N_25128);
and U26227 (N_26227,N_25117,N_25362);
nor U26228 (N_26228,N_25300,N_25625);
and U26229 (N_26229,N_25661,N_25278);
xnor U26230 (N_26230,N_25431,N_25049);
nand U26231 (N_26231,N_25611,N_25864);
nand U26232 (N_26232,N_25708,N_25211);
and U26233 (N_26233,N_25870,N_25921);
nor U26234 (N_26234,N_25311,N_25665);
and U26235 (N_26235,N_25951,N_25234);
xnor U26236 (N_26236,N_25947,N_25009);
xor U26237 (N_26237,N_25983,N_25835);
nand U26238 (N_26238,N_25712,N_25890);
or U26239 (N_26239,N_25502,N_25746);
xor U26240 (N_26240,N_25347,N_25545);
or U26241 (N_26241,N_25456,N_25679);
and U26242 (N_26242,N_25237,N_25338);
xor U26243 (N_26243,N_25816,N_25845);
xor U26244 (N_26244,N_25224,N_25395);
and U26245 (N_26245,N_25804,N_25466);
and U26246 (N_26246,N_25424,N_25216);
xor U26247 (N_26247,N_25672,N_25426);
and U26248 (N_26248,N_25168,N_25495);
nand U26249 (N_26249,N_25352,N_25334);
or U26250 (N_26250,N_25219,N_25799);
nor U26251 (N_26251,N_25894,N_25267);
xnor U26252 (N_26252,N_25999,N_25062);
or U26253 (N_26253,N_25690,N_25069);
or U26254 (N_26254,N_25568,N_25730);
nand U26255 (N_26255,N_25444,N_25800);
nor U26256 (N_26256,N_25608,N_25927);
xor U26257 (N_26257,N_25735,N_25706);
and U26258 (N_26258,N_25527,N_25606);
nor U26259 (N_26259,N_25885,N_25021);
nand U26260 (N_26260,N_25114,N_25083);
xnor U26261 (N_26261,N_25745,N_25596);
or U26262 (N_26262,N_25868,N_25346);
xnor U26263 (N_26263,N_25130,N_25647);
nand U26264 (N_26264,N_25259,N_25654);
and U26265 (N_26265,N_25408,N_25598);
and U26266 (N_26266,N_25358,N_25948);
nand U26267 (N_26267,N_25905,N_25607);
nand U26268 (N_26268,N_25559,N_25520);
or U26269 (N_26269,N_25418,N_25462);
nor U26270 (N_26270,N_25129,N_25602);
nand U26271 (N_26271,N_25696,N_25180);
nor U26272 (N_26272,N_25664,N_25035);
and U26273 (N_26273,N_25172,N_25945);
xor U26274 (N_26274,N_25087,N_25262);
nand U26275 (N_26275,N_25467,N_25001);
or U26276 (N_26276,N_25331,N_25376);
or U26277 (N_26277,N_25406,N_25461);
and U26278 (N_26278,N_25227,N_25982);
xor U26279 (N_26279,N_25577,N_25739);
nand U26280 (N_26280,N_25989,N_25164);
and U26281 (N_26281,N_25322,N_25838);
nand U26282 (N_26282,N_25883,N_25853);
and U26283 (N_26283,N_25081,N_25828);
nand U26284 (N_26284,N_25027,N_25939);
xor U26285 (N_26285,N_25096,N_25453);
nor U26286 (N_26286,N_25636,N_25729);
nor U26287 (N_26287,N_25473,N_25631);
nor U26288 (N_26288,N_25017,N_25203);
nor U26289 (N_26289,N_25010,N_25286);
or U26290 (N_26290,N_25480,N_25627);
or U26291 (N_26291,N_25616,N_25135);
and U26292 (N_26292,N_25289,N_25825);
and U26293 (N_26293,N_25377,N_25582);
and U26294 (N_26294,N_25152,N_25699);
xor U26295 (N_26295,N_25530,N_25634);
xnor U26296 (N_26296,N_25650,N_25584);
nor U26297 (N_26297,N_25195,N_25772);
or U26298 (N_26298,N_25653,N_25182);
and U26299 (N_26299,N_25315,N_25214);
or U26300 (N_26300,N_25297,N_25354);
and U26301 (N_26301,N_25481,N_25387);
and U26302 (N_26302,N_25476,N_25728);
or U26303 (N_26303,N_25874,N_25447);
or U26304 (N_26304,N_25978,N_25163);
or U26305 (N_26305,N_25593,N_25535);
and U26306 (N_26306,N_25550,N_25318);
xor U26307 (N_26307,N_25012,N_25225);
xnor U26308 (N_26308,N_25302,N_25681);
xnor U26309 (N_26309,N_25516,N_25235);
nand U26310 (N_26310,N_25067,N_25248);
or U26311 (N_26311,N_25793,N_25204);
nand U26312 (N_26312,N_25985,N_25784);
or U26313 (N_26313,N_25986,N_25873);
nand U26314 (N_26314,N_25987,N_25485);
nor U26315 (N_26315,N_25640,N_25886);
xnor U26316 (N_26316,N_25105,N_25848);
xnor U26317 (N_26317,N_25899,N_25423);
nor U26318 (N_26318,N_25852,N_25720);
nand U26319 (N_26319,N_25933,N_25862);
nor U26320 (N_26320,N_25952,N_25020);
xnor U26321 (N_26321,N_25510,N_25468);
nor U26322 (N_26322,N_25570,N_25086);
and U26323 (N_26323,N_25314,N_25953);
nor U26324 (N_26324,N_25340,N_25499);
or U26325 (N_26325,N_25177,N_25765);
nand U26326 (N_26326,N_25918,N_25265);
and U26327 (N_26327,N_25460,N_25742);
nor U26328 (N_26328,N_25109,N_25846);
nor U26329 (N_26329,N_25179,N_25332);
nand U26330 (N_26330,N_25518,N_25002);
and U26331 (N_26331,N_25194,N_25030);
or U26332 (N_26332,N_25052,N_25004);
xor U26333 (N_26333,N_25148,N_25630);
xor U26334 (N_26334,N_25932,N_25208);
nand U26335 (N_26335,N_25132,N_25492);
or U26336 (N_26336,N_25815,N_25806);
and U26337 (N_26337,N_25036,N_25391);
or U26338 (N_26338,N_25854,N_25388);
or U26339 (N_26339,N_25226,N_25863);
nor U26340 (N_26340,N_25756,N_25326);
nor U26341 (N_26341,N_25403,N_25930);
nor U26342 (N_26342,N_25065,N_25610);
xnor U26343 (N_26343,N_25250,N_25632);
and U26344 (N_26344,N_25666,N_25261);
xnor U26345 (N_26345,N_25174,N_25587);
or U26346 (N_26346,N_25459,N_25581);
xor U26347 (N_26347,N_25942,N_25844);
nor U26348 (N_26348,N_25290,N_25671);
and U26349 (N_26349,N_25175,N_25717);
nand U26350 (N_26350,N_25088,N_25692);
nand U26351 (N_26351,N_25307,N_25139);
nor U26352 (N_26352,N_25770,N_25747);
and U26353 (N_26353,N_25500,N_25173);
and U26354 (N_26354,N_25371,N_25452);
nor U26355 (N_26355,N_25967,N_25154);
nand U26356 (N_26356,N_25936,N_25131);
nand U26357 (N_26357,N_25529,N_25926);
xnor U26358 (N_26358,N_25370,N_25337);
or U26359 (N_26359,N_25450,N_25159);
or U26360 (N_26360,N_25722,N_25635);
nor U26361 (N_26361,N_25808,N_25777);
xnor U26362 (N_26362,N_25430,N_25693);
or U26363 (N_26363,N_25024,N_25973);
xnor U26364 (N_26364,N_25490,N_25824);
and U26365 (N_26365,N_25127,N_25571);
nand U26366 (N_26366,N_25629,N_25997);
xnor U26367 (N_26367,N_25031,N_25188);
and U26368 (N_26368,N_25073,N_25819);
nor U26369 (N_26369,N_25110,N_25597);
xnor U26370 (N_26370,N_25184,N_25626);
nor U26371 (N_26371,N_25954,N_25576);
or U26372 (N_26372,N_25589,N_25239);
or U26373 (N_26373,N_25178,N_25074);
or U26374 (N_26374,N_25435,N_25304);
and U26375 (N_26375,N_25879,N_25910);
nor U26376 (N_26376,N_25386,N_25966);
and U26377 (N_26377,N_25755,N_25676);
nand U26378 (N_26378,N_25751,N_25136);
xnor U26379 (N_26379,N_25976,N_25731);
nand U26380 (N_26380,N_25658,N_25422);
xor U26381 (N_26381,N_25901,N_25761);
xnor U26382 (N_26382,N_25291,N_25552);
xor U26383 (N_26383,N_25697,N_25008);
xor U26384 (N_26384,N_25270,N_25232);
and U26385 (N_26385,N_25156,N_25486);
nor U26386 (N_26386,N_25974,N_25782);
nand U26387 (N_26387,N_25614,N_25524);
xor U26388 (N_26388,N_25439,N_25392);
nor U26389 (N_26389,N_25084,N_25037);
or U26390 (N_26390,N_25506,N_25573);
or U26391 (N_26391,N_25931,N_25813);
or U26392 (N_26392,N_25859,N_25962);
nor U26393 (N_26393,N_25913,N_25702);
nand U26394 (N_26394,N_25189,N_25349);
xor U26395 (N_26395,N_25246,N_25365);
or U26396 (N_26396,N_25409,N_25221);
and U26397 (N_26397,N_25569,N_25662);
or U26398 (N_26398,N_25298,N_25236);
and U26399 (N_26399,N_25150,N_25817);
or U26400 (N_26400,N_25561,N_25546);
or U26401 (N_26401,N_25638,N_25309);
xnor U26402 (N_26402,N_25003,N_25600);
or U26403 (N_26403,N_25519,N_25308);
or U26404 (N_26404,N_25911,N_25727);
and U26405 (N_26405,N_25726,N_25539);
and U26406 (N_26406,N_25285,N_25543);
nor U26407 (N_26407,N_25116,N_25281);
xnor U26408 (N_26408,N_25149,N_25399);
nand U26409 (N_26409,N_25053,N_25335);
or U26410 (N_26410,N_25171,N_25710);
xnor U26411 (N_26411,N_25904,N_25078);
or U26412 (N_26412,N_25705,N_25375);
xnor U26413 (N_26413,N_25829,N_25866);
and U26414 (N_26414,N_25688,N_25724);
nand U26415 (N_26415,N_25317,N_25433);
nand U26416 (N_26416,N_25963,N_25994);
xnor U26417 (N_26417,N_25525,N_25544);
xnor U26418 (N_26418,N_25415,N_25505);
xor U26419 (N_26419,N_25907,N_25677);
or U26420 (N_26420,N_25282,N_25210);
and U26421 (N_26421,N_25231,N_25950);
or U26422 (N_26422,N_25541,N_25580);
xnor U26423 (N_26423,N_25090,N_25564);
nor U26424 (N_26424,N_25155,N_25320);
nand U26425 (N_26425,N_25714,N_25276);
and U26426 (N_26426,N_25303,N_25773);
and U26427 (N_26427,N_25397,N_25477);
or U26428 (N_26428,N_25736,N_25407);
nor U26429 (N_26429,N_25995,N_25919);
xnor U26430 (N_26430,N_25222,N_25511);
nor U26431 (N_26431,N_25732,N_25578);
nand U26432 (N_26432,N_25590,N_25855);
or U26433 (N_26433,N_25588,N_25272);
nor U26434 (N_26434,N_25814,N_25351);
xor U26435 (N_26435,N_25503,N_25562);
or U26436 (N_26436,N_25684,N_25850);
nand U26437 (N_26437,N_25169,N_25767);
or U26438 (N_26438,N_25646,N_25620);
nand U26439 (N_26439,N_25556,N_25394);
or U26440 (N_26440,N_25941,N_25313);
and U26441 (N_26441,N_25445,N_25205);
nand U26442 (N_26442,N_25190,N_25709);
xor U26443 (N_26443,N_25575,N_25019);
and U26444 (N_26444,N_25343,N_25651);
or U26445 (N_26445,N_25256,N_25493);
and U26446 (N_26446,N_25064,N_25716);
xnor U26447 (N_26447,N_25273,N_25121);
and U26448 (N_26448,N_25106,N_25151);
xnor U26449 (N_26449,N_25050,N_25585);
nor U26450 (N_26450,N_25443,N_25113);
or U26451 (N_26451,N_25628,N_25649);
and U26452 (N_26452,N_25016,N_25255);
xor U26453 (N_26453,N_25703,N_25192);
xor U26454 (N_26454,N_25916,N_25373);
nor U26455 (N_26455,N_25353,N_25613);
or U26456 (N_26456,N_25686,N_25479);
nand U26457 (N_26457,N_25442,N_25075);
and U26458 (N_26458,N_25810,N_25959);
and U26459 (N_26459,N_25080,N_25557);
xor U26460 (N_26460,N_25126,N_25955);
or U26461 (N_26461,N_25342,N_25803);
nor U26462 (N_26462,N_25143,N_25266);
xnor U26463 (N_26463,N_25296,N_25446);
and U26464 (N_26464,N_25489,N_25958);
or U26465 (N_26465,N_25170,N_25470);
xnor U26466 (N_26466,N_25042,N_25345);
nor U26467 (N_26467,N_25412,N_25260);
nor U26468 (N_26468,N_25396,N_25199);
and U26469 (N_26469,N_25560,N_25448);
and U26470 (N_26470,N_25100,N_25753);
and U26471 (N_26471,N_25682,N_25361);
and U26472 (N_26472,N_25419,N_25875);
nand U26473 (N_26473,N_25914,N_25013);
and U26474 (N_26474,N_25617,N_25441);
nand U26475 (N_26475,N_25254,N_25680);
or U26476 (N_26476,N_25968,N_25975);
or U26477 (N_26477,N_25484,N_25060);
xnor U26478 (N_26478,N_25827,N_25749);
or U26479 (N_26479,N_25618,N_25104);
nand U26480 (N_26480,N_25288,N_25796);
nor U26481 (N_26481,N_25549,N_25085);
xnor U26482 (N_26482,N_25107,N_25299);
and U26483 (N_26483,N_25436,N_25046);
nand U26484 (N_26484,N_25115,N_25483);
xnor U26485 (N_26485,N_25792,N_25612);
nor U26486 (N_26486,N_25421,N_25981);
xnor U26487 (N_26487,N_25509,N_25283);
xor U26488 (N_26488,N_25842,N_25892);
nand U26489 (N_26489,N_25768,N_25006);
nand U26490 (N_26490,N_25713,N_25380);
or U26491 (N_26491,N_25766,N_25363);
and U26492 (N_26492,N_25093,N_25759);
or U26493 (N_26493,N_25961,N_25437);
nor U26494 (N_26494,N_25257,N_25410);
and U26495 (N_26495,N_25066,N_25537);
xnor U26496 (N_26496,N_25348,N_25683);
nand U26497 (N_26497,N_25287,N_25929);
nand U26498 (N_26498,N_25734,N_25513);
or U26499 (N_26499,N_25258,N_25123);
xnor U26500 (N_26500,N_25879,N_25146);
xor U26501 (N_26501,N_25580,N_25546);
nand U26502 (N_26502,N_25804,N_25070);
nor U26503 (N_26503,N_25736,N_25447);
or U26504 (N_26504,N_25702,N_25190);
nor U26505 (N_26505,N_25998,N_25856);
or U26506 (N_26506,N_25481,N_25139);
nand U26507 (N_26507,N_25086,N_25313);
xor U26508 (N_26508,N_25215,N_25706);
or U26509 (N_26509,N_25181,N_25024);
nand U26510 (N_26510,N_25171,N_25836);
nand U26511 (N_26511,N_25945,N_25411);
nand U26512 (N_26512,N_25820,N_25354);
or U26513 (N_26513,N_25899,N_25644);
nand U26514 (N_26514,N_25293,N_25732);
or U26515 (N_26515,N_25253,N_25302);
nand U26516 (N_26516,N_25218,N_25984);
xor U26517 (N_26517,N_25989,N_25452);
nand U26518 (N_26518,N_25664,N_25582);
or U26519 (N_26519,N_25366,N_25185);
and U26520 (N_26520,N_25770,N_25504);
xor U26521 (N_26521,N_25016,N_25541);
or U26522 (N_26522,N_25566,N_25942);
or U26523 (N_26523,N_25587,N_25084);
xor U26524 (N_26524,N_25319,N_25165);
xnor U26525 (N_26525,N_25356,N_25114);
or U26526 (N_26526,N_25790,N_25900);
nand U26527 (N_26527,N_25075,N_25538);
xnor U26528 (N_26528,N_25580,N_25797);
nand U26529 (N_26529,N_25861,N_25095);
or U26530 (N_26530,N_25555,N_25293);
xor U26531 (N_26531,N_25618,N_25118);
nor U26532 (N_26532,N_25821,N_25679);
nand U26533 (N_26533,N_25872,N_25961);
nand U26534 (N_26534,N_25647,N_25151);
nor U26535 (N_26535,N_25740,N_25552);
or U26536 (N_26536,N_25236,N_25808);
and U26537 (N_26537,N_25436,N_25133);
nand U26538 (N_26538,N_25205,N_25048);
and U26539 (N_26539,N_25941,N_25769);
nor U26540 (N_26540,N_25938,N_25306);
nand U26541 (N_26541,N_25743,N_25050);
and U26542 (N_26542,N_25055,N_25342);
or U26543 (N_26543,N_25247,N_25380);
and U26544 (N_26544,N_25077,N_25105);
nor U26545 (N_26545,N_25909,N_25256);
xor U26546 (N_26546,N_25231,N_25175);
and U26547 (N_26547,N_25156,N_25880);
nand U26548 (N_26548,N_25667,N_25355);
and U26549 (N_26549,N_25957,N_25058);
xnor U26550 (N_26550,N_25796,N_25133);
nor U26551 (N_26551,N_25193,N_25535);
or U26552 (N_26552,N_25490,N_25489);
nor U26553 (N_26553,N_25522,N_25871);
nor U26554 (N_26554,N_25964,N_25976);
nor U26555 (N_26555,N_25302,N_25528);
nor U26556 (N_26556,N_25511,N_25676);
xnor U26557 (N_26557,N_25847,N_25430);
nand U26558 (N_26558,N_25500,N_25857);
and U26559 (N_26559,N_25923,N_25799);
or U26560 (N_26560,N_25618,N_25977);
nor U26561 (N_26561,N_25564,N_25141);
nand U26562 (N_26562,N_25630,N_25051);
nor U26563 (N_26563,N_25982,N_25334);
or U26564 (N_26564,N_25772,N_25932);
xor U26565 (N_26565,N_25589,N_25625);
and U26566 (N_26566,N_25610,N_25373);
nand U26567 (N_26567,N_25009,N_25489);
xnor U26568 (N_26568,N_25235,N_25796);
or U26569 (N_26569,N_25830,N_25589);
or U26570 (N_26570,N_25798,N_25613);
and U26571 (N_26571,N_25941,N_25940);
xor U26572 (N_26572,N_25306,N_25077);
nand U26573 (N_26573,N_25881,N_25268);
nand U26574 (N_26574,N_25050,N_25834);
nor U26575 (N_26575,N_25272,N_25059);
xor U26576 (N_26576,N_25934,N_25938);
nand U26577 (N_26577,N_25528,N_25973);
and U26578 (N_26578,N_25193,N_25704);
xor U26579 (N_26579,N_25126,N_25434);
or U26580 (N_26580,N_25569,N_25659);
and U26581 (N_26581,N_25639,N_25880);
and U26582 (N_26582,N_25722,N_25590);
or U26583 (N_26583,N_25369,N_25847);
or U26584 (N_26584,N_25043,N_25211);
xnor U26585 (N_26585,N_25406,N_25272);
nor U26586 (N_26586,N_25585,N_25247);
nor U26587 (N_26587,N_25892,N_25423);
xor U26588 (N_26588,N_25500,N_25098);
and U26589 (N_26589,N_25091,N_25793);
nor U26590 (N_26590,N_25437,N_25495);
nand U26591 (N_26591,N_25649,N_25690);
nor U26592 (N_26592,N_25780,N_25779);
xor U26593 (N_26593,N_25423,N_25967);
and U26594 (N_26594,N_25848,N_25795);
nand U26595 (N_26595,N_25709,N_25459);
nand U26596 (N_26596,N_25045,N_25373);
nor U26597 (N_26597,N_25631,N_25033);
or U26598 (N_26598,N_25304,N_25128);
nor U26599 (N_26599,N_25292,N_25617);
or U26600 (N_26600,N_25695,N_25879);
xnor U26601 (N_26601,N_25958,N_25904);
or U26602 (N_26602,N_25083,N_25601);
and U26603 (N_26603,N_25279,N_25950);
nand U26604 (N_26604,N_25025,N_25737);
and U26605 (N_26605,N_25165,N_25955);
or U26606 (N_26606,N_25899,N_25770);
nand U26607 (N_26607,N_25999,N_25609);
and U26608 (N_26608,N_25483,N_25475);
or U26609 (N_26609,N_25916,N_25914);
nor U26610 (N_26610,N_25194,N_25441);
and U26611 (N_26611,N_25124,N_25848);
and U26612 (N_26612,N_25725,N_25314);
nand U26613 (N_26613,N_25327,N_25371);
nand U26614 (N_26614,N_25464,N_25351);
xor U26615 (N_26615,N_25879,N_25200);
nand U26616 (N_26616,N_25012,N_25823);
nor U26617 (N_26617,N_25517,N_25786);
or U26618 (N_26618,N_25014,N_25114);
nand U26619 (N_26619,N_25023,N_25976);
nor U26620 (N_26620,N_25201,N_25235);
xor U26621 (N_26621,N_25886,N_25519);
nand U26622 (N_26622,N_25110,N_25086);
xnor U26623 (N_26623,N_25291,N_25372);
xnor U26624 (N_26624,N_25733,N_25888);
xor U26625 (N_26625,N_25555,N_25409);
and U26626 (N_26626,N_25031,N_25027);
and U26627 (N_26627,N_25325,N_25932);
or U26628 (N_26628,N_25170,N_25394);
nor U26629 (N_26629,N_25206,N_25397);
or U26630 (N_26630,N_25804,N_25268);
and U26631 (N_26631,N_25706,N_25095);
or U26632 (N_26632,N_25567,N_25126);
and U26633 (N_26633,N_25296,N_25280);
nor U26634 (N_26634,N_25139,N_25009);
nand U26635 (N_26635,N_25166,N_25107);
xor U26636 (N_26636,N_25602,N_25090);
nor U26637 (N_26637,N_25737,N_25586);
xor U26638 (N_26638,N_25303,N_25026);
and U26639 (N_26639,N_25230,N_25698);
nand U26640 (N_26640,N_25994,N_25607);
or U26641 (N_26641,N_25782,N_25548);
nor U26642 (N_26642,N_25737,N_25882);
nand U26643 (N_26643,N_25771,N_25755);
and U26644 (N_26644,N_25031,N_25605);
xor U26645 (N_26645,N_25568,N_25589);
or U26646 (N_26646,N_25705,N_25486);
xnor U26647 (N_26647,N_25113,N_25842);
and U26648 (N_26648,N_25444,N_25447);
and U26649 (N_26649,N_25048,N_25884);
nand U26650 (N_26650,N_25686,N_25467);
or U26651 (N_26651,N_25429,N_25701);
nor U26652 (N_26652,N_25653,N_25732);
or U26653 (N_26653,N_25762,N_25557);
nand U26654 (N_26654,N_25762,N_25392);
nor U26655 (N_26655,N_25461,N_25641);
or U26656 (N_26656,N_25340,N_25983);
or U26657 (N_26657,N_25726,N_25584);
nand U26658 (N_26658,N_25104,N_25815);
or U26659 (N_26659,N_25948,N_25910);
nand U26660 (N_26660,N_25745,N_25365);
xnor U26661 (N_26661,N_25874,N_25225);
or U26662 (N_26662,N_25439,N_25282);
xor U26663 (N_26663,N_25236,N_25949);
nand U26664 (N_26664,N_25264,N_25296);
nor U26665 (N_26665,N_25120,N_25395);
nor U26666 (N_26666,N_25897,N_25039);
nor U26667 (N_26667,N_25196,N_25181);
or U26668 (N_26668,N_25104,N_25453);
or U26669 (N_26669,N_25882,N_25896);
xor U26670 (N_26670,N_25291,N_25460);
xnor U26671 (N_26671,N_25356,N_25181);
nor U26672 (N_26672,N_25240,N_25368);
xor U26673 (N_26673,N_25714,N_25904);
xor U26674 (N_26674,N_25877,N_25420);
nor U26675 (N_26675,N_25332,N_25054);
xnor U26676 (N_26676,N_25634,N_25048);
nand U26677 (N_26677,N_25724,N_25455);
or U26678 (N_26678,N_25916,N_25159);
nand U26679 (N_26679,N_25063,N_25179);
nor U26680 (N_26680,N_25749,N_25722);
or U26681 (N_26681,N_25417,N_25567);
and U26682 (N_26682,N_25183,N_25150);
nor U26683 (N_26683,N_25514,N_25094);
or U26684 (N_26684,N_25657,N_25504);
nor U26685 (N_26685,N_25157,N_25263);
xnor U26686 (N_26686,N_25085,N_25348);
and U26687 (N_26687,N_25092,N_25158);
or U26688 (N_26688,N_25813,N_25771);
xnor U26689 (N_26689,N_25078,N_25331);
nor U26690 (N_26690,N_25450,N_25012);
xnor U26691 (N_26691,N_25733,N_25823);
or U26692 (N_26692,N_25334,N_25029);
xor U26693 (N_26693,N_25695,N_25000);
and U26694 (N_26694,N_25086,N_25254);
and U26695 (N_26695,N_25378,N_25304);
or U26696 (N_26696,N_25073,N_25249);
or U26697 (N_26697,N_25449,N_25908);
xor U26698 (N_26698,N_25635,N_25868);
or U26699 (N_26699,N_25349,N_25515);
xor U26700 (N_26700,N_25362,N_25717);
xnor U26701 (N_26701,N_25015,N_25319);
nand U26702 (N_26702,N_25838,N_25522);
xnor U26703 (N_26703,N_25706,N_25894);
nand U26704 (N_26704,N_25246,N_25139);
nor U26705 (N_26705,N_25810,N_25039);
xnor U26706 (N_26706,N_25698,N_25688);
nand U26707 (N_26707,N_25542,N_25708);
xor U26708 (N_26708,N_25174,N_25999);
nor U26709 (N_26709,N_25561,N_25279);
and U26710 (N_26710,N_25446,N_25557);
nor U26711 (N_26711,N_25118,N_25900);
and U26712 (N_26712,N_25807,N_25173);
nand U26713 (N_26713,N_25033,N_25055);
and U26714 (N_26714,N_25353,N_25494);
nand U26715 (N_26715,N_25168,N_25266);
nor U26716 (N_26716,N_25582,N_25595);
nand U26717 (N_26717,N_25857,N_25832);
nand U26718 (N_26718,N_25287,N_25646);
nor U26719 (N_26719,N_25957,N_25909);
nand U26720 (N_26720,N_25891,N_25676);
nor U26721 (N_26721,N_25287,N_25700);
nand U26722 (N_26722,N_25566,N_25116);
nor U26723 (N_26723,N_25050,N_25097);
nor U26724 (N_26724,N_25316,N_25313);
and U26725 (N_26725,N_25791,N_25913);
and U26726 (N_26726,N_25794,N_25019);
nor U26727 (N_26727,N_25179,N_25151);
nand U26728 (N_26728,N_25766,N_25070);
and U26729 (N_26729,N_25203,N_25372);
xor U26730 (N_26730,N_25293,N_25711);
nand U26731 (N_26731,N_25271,N_25904);
nand U26732 (N_26732,N_25794,N_25149);
xnor U26733 (N_26733,N_25072,N_25348);
nand U26734 (N_26734,N_25737,N_25601);
xor U26735 (N_26735,N_25103,N_25618);
or U26736 (N_26736,N_25625,N_25798);
xor U26737 (N_26737,N_25920,N_25130);
xor U26738 (N_26738,N_25436,N_25410);
nand U26739 (N_26739,N_25713,N_25360);
nor U26740 (N_26740,N_25899,N_25848);
xor U26741 (N_26741,N_25424,N_25518);
or U26742 (N_26742,N_25814,N_25514);
nand U26743 (N_26743,N_25021,N_25357);
xor U26744 (N_26744,N_25891,N_25947);
or U26745 (N_26745,N_25173,N_25345);
nor U26746 (N_26746,N_25968,N_25155);
and U26747 (N_26747,N_25049,N_25655);
nor U26748 (N_26748,N_25944,N_25935);
nand U26749 (N_26749,N_25261,N_25926);
xor U26750 (N_26750,N_25892,N_25196);
nand U26751 (N_26751,N_25038,N_25905);
or U26752 (N_26752,N_25984,N_25712);
xor U26753 (N_26753,N_25616,N_25819);
or U26754 (N_26754,N_25977,N_25971);
nor U26755 (N_26755,N_25434,N_25287);
xnor U26756 (N_26756,N_25492,N_25646);
and U26757 (N_26757,N_25207,N_25132);
or U26758 (N_26758,N_25425,N_25724);
nand U26759 (N_26759,N_25947,N_25188);
and U26760 (N_26760,N_25414,N_25519);
and U26761 (N_26761,N_25747,N_25407);
nand U26762 (N_26762,N_25380,N_25524);
nand U26763 (N_26763,N_25839,N_25163);
nand U26764 (N_26764,N_25120,N_25787);
xnor U26765 (N_26765,N_25191,N_25935);
and U26766 (N_26766,N_25831,N_25409);
nand U26767 (N_26767,N_25898,N_25066);
nand U26768 (N_26768,N_25262,N_25436);
xor U26769 (N_26769,N_25799,N_25738);
and U26770 (N_26770,N_25364,N_25942);
or U26771 (N_26771,N_25768,N_25432);
or U26772 (N_26772,N_25399,N_25641);
or U26773 (N_26773,N_25085,N_25694);
and U26774 (N_26774,N_25727,N_25415);
and U26775 (N_26775,N_25153,N_25391);
nor U26776 (N_26776,N_25564,N_25272);
nor U26777 (N_26777,N_25391,N_25260);
nor U26778 (N_26778,N_25828,N_25276);
and U26779 (N_26779,N_25602,N_25672);
and U26780 (N_26780,N_25032,N_25655);
xnor U26781 (N_26781,N_25822,N_25916);
or U26782 (N_26782,N_25936,N_25747);
or U26783 (N_26783,N_25049,N_25260);
xor U26784 (N_26784,N_25734,N_25030);
xor U26785 (N_26785,N_25306,N_25660);
and U26786 (N_26786,N_25126,N_25529);
or U26787 (N_26787,N_25294,N_25178);
xor U26788 (N_26788,N_25597,N_25710);
nor U26789 (N_26789,N_25654,N_25082);
nor U26790 (N_26790,N_25371,N_25830);
and U26791 (N_26791,N_25197,N_25840);
nand U26792 (N_26792,N_25528,N_25827);
nand U26793 (N_26793,N_25723,N_25566);
nand U26794 (N_26794,N_25026,N_25030);
and U26795 (N_26795,N_25163,N_25285);
xor U26796 (N_26796,N_25021,N_25350);
or U26797 (N_26797,N_25159,N_25392);
xor U26798 (N_26798,N_25490,N_25076);
nor U26799 (N_26799,N_25089,N_25808);
nand U26800 (N_26800,N_25838,N_25288);
and U26801 (N_26801,N_25647,N_25369);
nor U26802 (N_26802,N_25211,N_25736);
nand U26803 (N_26803,N_25625,N_25822);
xnor U26804 (N_26804,N_25751,N_25407);
xor U26805 (N_26805,N_25988,N_25344);
nor U26806 (N_26806,N_25882,N_25132);
nor U26807 (N_26807,N_25963,N_25645);
or U26808 (N_26808,N_25766,N_25802);
xor U26809 (N_26809,N_25106,N_25248);
nand U26810 (N_26810,N_25495,N_25486);
xor U26811 (N_26811,N_25122,N_25639);
nand U26812 (N_26812,N_25093,N_25009);
or U26813 (N_26813,N_25918,N_25058);
nand U26814 (N_26814,N_25921,N_25226);
or U26815 (N_26815,N_25299,N_25250);
or U26816 (N_26816,N_25754,N_25017);
or U26817 (N_26817,N_25591,N_25939);
xor U26818 (N_26818,N_25031,N_25374);
nand U26819 (N_26819,N_25065,N_25995);
and U26820 (N_26820,N_25500,N_25001);
xor U26821 (N_26821,N_25557,N_25559);
nand U26822 (N_26822,N_25790,N_25795);
nand U26823 (N_26823,N_25203,N_25857);
nand U26824 (N_26824,N_25106,N_25487);
xnor U26825 (N_26825,N_25308,N_25802);
or U26826 (N_26826,N_25543,N_25738);
nand U26827 (N_26827,N_25289,N_25041);
nand U26828 (N_26828,N_25550,N_25536);
and U26829 (N_26829,N_25970,N_25728);
or U26830 (N_26830,N_25138,N_25472);
nand U26831 (N_26831,N_25944,N_25869);
or U26832 (N_26832,N_25443,N_25549);
or U26833 (N_26833,N_25401,N_25626);
and U26834 (N_26834,N_25459,N_25367);
nor U26835 (N_26835,N_25433,N_25120);
and U26836 (N_26836,N_25663,N_25233);
xnor U26837 (N_26837,N_25413,N_25367);
nor U26838 (N_26838,N_25602,N_25686);
nor U26839 (N_26839,N_25084,N_25832);
and U26840 (N_26840,N_25359,N_25798);
and U26841 (N_26841,N_25570,N_25696);
and U26842 (N_26842,N_25990,N_25115);
or U26843 (N_26843,N_25481,N_25797);
xnor U26844 (N_26844,N_25932,N_25782);
nor U26845 (N_26845,N_25219,N_25284);
and U26846 (N_26846,N_25276,N_25114);
and U26847 (N_26847,N_25179,N_25923);
nor U26848 (N_26848,N_25760,N_25954);
and U26849 (N_26849,N_25109,N_25049);
nand U26850 (N_26850,N_25794,N_25462);
nand U26851 (N_26851,N_25614,N_25477);
and U26852 (N_26852,N_25701,N_25079);
nor U26853 (N_26853,N_25431,N_25242);
nand U26854 (N_26854,N_25825,N_25067);
or U26855 (N_26855,N_25269,N_25119);
or U26856 (N_26856,N_25353,N_25374);
xnor U26857 (N_26857,N_25733,N_25783);
nor U26858 (N_26858,N_25723,N_25951);
and U26859 (N_26859,N_25526,N_25740);
xor U26860 (N_26860,N_25967,N_25266);
nand U26861 (N_26861,N_25469,N_25358);
nand U26862 (N_26862,N_25961,N_25935);
nor U26863 (N_26863,N_25609,N_25163);
xor U26864 (N_26864,N_25510,N_25840);
xnor U26865 (N_26865,N_25816,N_25791);
nand U26866 (N_26866,N_25085,N_25448);
nand U26867 (N_26867,N_25924,N_25098);
and U26868 (N_26868,N_25834,N_25423);
or U26869 (N_26869,N_25853,N_25000);
xnor U26870 (N_26870,N_25421,N_25002);
and U26871 (N_26871,N_25177,N_25758);
xnor U26872 (N_26872,N_25080,N_25102);
or U26873 (N_26873,N_25323,N_25905);
nand U26874 (N_26874,N_25260,N_25896);
or U26875 (N_26875,N_25770,N_25575);
and U26876 (N_26876,N_25879,N_25823);
nand U26877 (N_26877,N_25294,N_25286);
nand U26878 (N_26878,N_25132,N_25596);
nand U26879 (N_26879,N_25383,N_25889);
and U26880 (N_26880,N_25258,N_25344);
or U26881 (N_26881,N_25686,N_25031);
nand U26882 (N_26882,N_25298,N_25492);
and U26883 (N_26883,N_25407,N_25929);
and U26884 (N_26884,N_25371,N_25920);
and U26885 (N_26885,N_25496,N_25112);
and U26886 (N_26886,N_25282,N_25801);
xor U26887 (N_26887,N_25233,N_25633);
and U26888 (N_26888,N_25112,N_25841);
and U26889 (N_26889,N_25717,N_25893);
xnor U26890 (N_26890,N_25142,N_25877);
xor U26891 (N_26891,N_25969,N_25778);
xnor U26892 (N_26892,N_25327,N_25275);
and U26893 (N_26893,N_25769,N_25110);
nand U26894 (N_26894,N_25053,N_25421);
nor U26895 (N_26895,N_25485,N_25049);
nor U26896 (N_26896,N_25432,N_25078);
nor U26897 (N_26897,N_25899,N_25133);
xor U26898 (N_26898,N_25944,N_25724);
nand U26899 (N_26899,N_25282,N_25167);
nor U26900 (N_26900,N_25821,N_25378);
nand U26901 (N_26901,N_25616,N_25922);
nand U26902 (N_26902,N_25730,N_25937);
nor U26903 (N_26903,N_25755,N_25899);
or U26904 (N_26904,N_25597,N_25695);
nand U26905 (N_26905,N_25187,N_25440);
nand U26906 (N_26906,N_25773,N_25222);
nand U26907 (N_26907,N_25013,N_25147);
xor U26908 (N_26908,N_25121,N_25447);
nor U26909 (N_26909,N_25794,N_25688);
xnor U26910 (N_26910,N_25172,N_25411);
nand U26911 (N_26911,N_25395,N_25962);
nand U26912 (N_26912,N_25012,N_25539);
or U26913 (N_26913,N_25665,N_25816);
and U26914 (N_26914,N_25549,N_25272);
xor U26915 (N_26915,N_25919,N_25422);
and U26916 (N_26916,N_25074,N_25761);
nor U26917 (N_26917,N_25341,N_25254);
nand U26918 (N_26918,N_25354,N_25996);
and U26919 (N_26919,N_25762,N_25828);
or U26920 (N_26920,N_25438,N_25059);
nor U26921 (N_26921,N_25324,N_25954);
and U26922 (N_26922,N_25383,N_25077);
xor U26923 (N_26923,N_25475,N_25904);
or U26924 (N_26924,N_25056,N_25300);
and U26925 (N_26925,N_25469,N_25741);
or U26926 (N_26926,N_25297,N_25413);
or U26927 (N_26927,N_25817,N_25836);
nand U26928 (N_26928,N_25912,N_25159);
nand U26929 (N_26929,N_25828,N_25368);
xor U26930 (N_26930,N_25891,N_25222);
nor U26931 (N_26931,N_25052,N_25211);
and U26932 (N_26932,N_25326,N_25962);
nor U26933 (N_26933,N_25973,N_25926);
nor U26934 (N_26934,N_25952,N_25036);
or U26935 (N_26935,N_25666,N_25479);
nor U26936 (N_26936,N_25640,N_25115);
nand U26937 (N_26937,N_25099,N_25948);
nor U26938 (N_26938,N_25121,N_25176);
nor U26939 (N_26939,N_25348,N_25007);
nor U26940 (N_26940,N_25298,N_25016);
xor U26941 (N_26941,N_25487,N_25387);
xnor U26942 (N_26942,N_25016,N_25348);
xor U26943 (N_26943,N_25874,N_25072);
or U26944 (N_26944,N_25607,N_25332);
nor U26945 (N_26945,N_25047,N_25754);
xor U26946 (N_26946,N_25709,N_25656);
and U26947 (N_26947,N_25450,N_25393);
or U26948 (N_26948,N_25238,N_25207);
nand U26949 (N_26949,N_25641,N_25932);
nand U26950 (N_26950,N_25125,N_25706);
or U26951 (N_26951,N_25872,N_25784);
nand U26952 (N_26952,N_25286,N_25856);
and U26953 (N_26953,N_25629,N_25227);
or U26954 (N_26954,N_25908,N_25780);
nor U26955 (N_26955,N_25199,N_25620);
xor U26956 (N_26956,N_25683,N_25432);
or U26957 (N_26957,N_25854,N_25077);
nor U26958 (N_26958,N_25544,N_25492);
or U26959 (N_26959,N_25094,N_25507);
nor U26960 (N_26960,N_25188,N_25575);
and U26961 (N_26961,N_25902,N_25315);
and U26962 (N_26962,N_25290,N_25782);
nand U26963 (N_26963,N_25969,N_25600);
or U26964 (N_26964,N_25269,N_25191);
nand U26965 (N_26965,N_25694,N_25514);
and U26966 (N_26966,N_25161,N_25979);
nand U26967 (N_26967,N_25987,N_25289);
or U26968 (N_26968,N_25868,N_25584);
nor U26969 (N_26969,N_25211,N_25452);
nand U26970 (N_26970,N_25528,N_25186);
nand U26971 (N_26971,N_25290,N_25388);
and U26972 (N_26972,N_25913,N_25157);
or U26973 (N_26973,N_25039,N_25557);
and U26974 (N_26974,N_25235,N_25749);
xor U26975 (N_26975,N_25859,N_25746);
or U26976 (N_26976,N_25262,N_25879);
or U26977 (N_26977,N_25043,N_25362);
nand U26978 (N_26978,N_25320,N_25775);
nor U26979 (N_26979,N_25026,N_25146);
xnor U26980 (N_26980,N_25304,N_25075);
and U26981 (N_26981,N_25984,N_25491);
and U26982 (N_26982,N_25761,N_25101);
nand U26983 (N_26983,N_25870,N_25174);
nand U26984 (N_26984,N_25846,N_25996);
nand U26985 (N_26985,N_25780,N_25137);
and U26986 (N_26986,N_25036,N_25931);
nand U26987 (N_26987,N_25379,N_25661);
or U26988 (N_26988,N_25590,N_25685);
xor U26989 (N_26989,N_25614,N_25485);
xnor U26990 (N_26990,N_25549,N_25308);
nor U26991 (N_26991,N_25512,N_25588);
and U26992 (N_26992,N_25741,N_25023);
and U26993 (N_26993,N_25492,N_25285);
nor U26994 (N_26994,N_25403,N_25231);
and U26995 (N_26995,N_25849,N_25031);
nor U26996 (N_26996,N_25329,N_25356);
nor U26997 (N_26997,N_25616,N_25296);
xor U26998 (N_26998,N_25872,N_25245);
or U26999 (N_26999,N_25878,N_25942);
nor U27000 (N_27000,N_26121,N_26799);
nand U27001 (N_27001,N_26399,N_26979);
nand U27002 (N_27002,N_26343,N_26998);
and U27003 (N_27003,N_26018,N_26826);
and U27004 (N_27004,N_26909,N_26734);
and U27005 (N_27005,N_26823,N_26810);
nor U27006 (N_27006,N_26987,N_26394);
or U27007 (N_27007,N_26054,N_26337);
xnor U27008 (N_27008,N_26384,N_26746);
nand U27009 (N_27009,N_26002,N_26800);
or U27010 (N_27010,N_26463,N_26190);
nor U27011 (N_27011,N_26038,N_26499);
and U27012 (N_27012,N_26392,N_26700);
and U27013 (N_27013,N_26378,N_26990);
nor U27014 (N_27014,N_26162,N_26620);
nor U27015 (N_27015,N_26003,N_26593);
and U27016 (N_27016,N_26505,N_26094);
xnor U27017 (N_27017,N_26296,N_26495);
nand U27018 (N_27018,N_26250,N_26970);
and U27019 (N_27019,N_26313,N_26782);
xor U27020 (N_27020,N_26994,N_26325);
xnor U27021 (N_27021,N_26039,N_26637);
or U27022 (N_27022,N_26662,N_26778);
or U27023 (N_27023,N_26284,N_26073);
nor U27024 (N_27024,N_26780,N_26572);
and U27025 (N_27025,N_26940,N_26923);
nand U27026 (N_27026,N_26096,N_26207);
and U27027 (N_27027,N_26693,N_26506);
or U27028 (N_27028,N_26651,N_26988);
xnor U27029 (N_27029,N_26084,N_26975);
or U27030 (N_27030,N_26544,N_26008);
and U27031 (N_27031,N_26777,N_26640);
nand U27032 (N_27032,N_26441,N_26959);
and U27033 (N_27033,N_26992,N_26231);
nand U27034 (N_27034,N_26426,N_26206);
nor U27035 (N_27035,N_26043,N_26108);
nand U27036 (N_27036,N_26045,N_26772);
nand U27037 (N_27037,N_26664,N_26254);
xor U27038 (N_27038,N_26635,N_26501);
or U27039 (N_27039,N_26532,N_26654);
nand U27040 (N_27040,N_26419,N_26739);
and U27041 (N_27041,N_26571,N_26014);
nand U27042 (N_27042,N_26007,N_26321);
and U27043 (N_27043,N_26704,N_26276);
nor U27044 (N_27044,N_26576,N_26416);
nor U27045 (N_27045,N_26268,N_26507);
and U27046 (N_27046,N_26359,N_26971);
and U27047 (N_27047,N_26630,N_26251);
and U27048 (N_27048,N_26633,N_26607);
nand U27049 (N_27049,N_26997,N_26290);
nand U27050 (N_27050,N_26615,N_26143);
nand U27051 (N_27051,N_26281,N_26036);
nand U27052 (N_27052,N_26145,N_26801);
nor U27053 (N_27053,N_26921,N_26027);
and U27054 (N_27054,N_26591,N_26172);
nor U27055 (N_27055,N_26346,N_26831);
and U27056 (N_27056,N_26872,N_26361);
nor U27057 (N_27057,N_26454,N_26993);
nor U27058 (N_27058,N_26918,N_26811);
nand U27059 (N_27059,N_26118,N_26585);
and U27060 (N_27060,N_26461,N_26851);
nand U27061 (N_27061,N_26349,N_26522);
nor U27062 (N_27062,N_26016,N_26983);
or U27063 (N_27063,N_26294,N_26698);
xnor U27064 (N_27064,N_26056,N_26030);
nor U27065 (N_27065,N_26087,N_26862);
nand U27066 (N_27066,N_26791,N_26414);
or U27067 (N_27067,N_26147,N_26041);
nor U27068 (N_27068,N_26053,N_26853);
nor U27069 (N_27069,N_26995,N_26098);
or U27070 (N_27070,N_26525,N_26339);
nor U27071 (N_27071,N_26939,N_26345);
and U27072 (N_27072,N_26164,N_26974);
or U27073 (N_27073,N_26740,N_26064);
nand U27074 (N_27074,N_26083,N_26534);
or U27075 (N_27075,N_26655,N_26735);
or U27076 (N_27076,N_26813,N_26082);
xnor U27077 (N_27077,N_26199,N_26095);
or U27078 (N_27078,N_26459,N_26964);
or U27079 (N_27079,N_26197,N_26864);
and U27080 (N_27080,N_26561,N_26881);
and U27081 (N_27081,N_26308,N_26950);
nor U27082 (N_27082,N_26338,N_26890);
nor U27083 (N_27083,N_26418,N_26049);
and U27084 (N_27084,N_26491,N_26265);
nor U27085 (N_27085,N_26893,N_26867);
and U27086 (N_27086,N_26672,N_26882);
nand U27087 (N_27087,N_26099,N_26636);
or U27088 (N_27088,N_26606,N_26747);
nor U27089 (N_27089,N_26031,N_26383);
nor U27090 (N_27090,N_26898,N_26784);
nor U27091 (N_27091,N_26945,N_26932);
nor U27092 (N_27092,N_26960,N_26942);
or U27093 (N_27093,N_26330,N_26627);
or U27094 (N_27094,N_26171,N_26194);
xnor U27095 (N_27095,N_26165,N_26671);
xnor U27096 (N_27096,N_26827,N_26825);
nor U27097 (N_27097,N_26114,N_26293);
nor U27098 (N_27098,N_26388,N_26497);
or U27099 (N_27099,N_26173,N_26931);
and U27100 (N_27100,N_26363,N_26248);
nand U27101 (N_27101,N_26528,N_26978);
xnor U27102 (N_27102,N_26322,N_26445);
xnor U27103 (N_27103,N_26598,N_26315);
nand U27104 (N_27104,N_26227,N_26884);
nand U27105 (N_27105,N_26277,N_26547);
nand U27106 (N_27106,N_26260,N_26480);
and U27107 (N_27107,N_26299,N_26798);
xor U27108 (N_27108,N_26174,N_26665);
nand U27109 (N_27109,N_26870,N_26077);
or U27110 (N_27110,N_26437,N_26060);
nor U27111 (N_27111,N_26889,N_26582);
nand U27112 (N_27112,N_26409,N_26543);
and U27113 (N_27113,N_26262,N_26692);
or U27114 (N_27114,N_26267,N_26368);
and U27115 (N_27115,N_26317,N_26223);
nand U27116 (N_27116,N_26424,N_26812);
nor U27117 (N_27117,N_26765,N_26047);
nand U27118 (N_27118,N_26433,N_26580);
nand U27119 (N_27119,N_26006,N_26233);
nand U27120 (N_27120,N_26217,N_26050);
xnor U27121 (N_27121,N_26727,N_26972);
nor U27122 (N_27122,N_26624,N_26819);
and U27123 (N_27123,N_26604,N_26449);
xor U27124 (N_27124,N_26494,N_26177);
or U27125 (N_27125,N_26849,N_26843);
or U27126 (N_27126,N_26367,N_26726);
or U27127 (N_27127,N_26020,N_26518);
nor U27128 (N_27128,N_26485,N_26496);
and U27129 (N_27129,N_26963,N_26523);
nor U27130 (N_27130,N_26478,N_26569);
and U27131 (N_27131,N_26808,N_26913);
nor U27132 (N_27132,N_26832,N_26677);
nor U27133 (N_27133,N_26237,N_26781);
and U27134 (N_27134,N_26824,N_26906);
and U27135 (N_27135,N_26420,N_26895);
xnor U27136 (N_27136,N_26958,N_26065);
nor U27137 (N_27137,N_26151,N_26148);
nand U27138 (N_27138,N_26529,N_26253);
or U27139 (N_27139,N_26481,N_26645);
nand U27140 (N_27140,N_26841,N_26980);
and U27141 (N_27141,N_26548,N_26466);
nand U27142 (N_27142,N_26405,N_26751);
and U27143 (N_27143,N_26689,N_26400);
and U27144 (N_27144,N_26075,N_26435);
nor U27145 (N_27145,N_26397,N_26925);
or U27146 (N_27146,N_26512,N_26549);
and U27147 (N_27147,N_26951,N_26009);
or U27148 (N_27148,N_26771,N_26842);
xnor U27149 (N_27149,N_26103,N_26275);
or U27150 (N_27150,N_26896,N_26219);
and U27151 (N_27151,N_26563,N_26152);
and U27152 (N_27152,N_26017,N_26089);
nor U27153 (N_27153,N_26464,N_26484);
nor U27154 (N_27154,N_26473,N_26888);
and U27155 (N_27155,N_26858,N_26019);
or U27156 (N_27156,N_26912,N_26848);
and U27157 (N_27157,N_26709,N_26954);
nand U27158 (N_27158,N_26395,N_26364);
and U27159 (N_27159,N_26001,N_26042);
and U27160 (N_27160,N_26957,N_26266);
xnor U27161 (N_27161,N_26865,N_26252);
or U27162 (N_27162,N_26144,N_26465);
nand U27163 (N_27163,N_26292,N_26193);
nand U27164 (N_27164,N_26136,N_26188);
xor U27165 (N_27165,N_26638,N_26897);
or U27166 (N_27166,N_26490,N_26869);
nor U27167 (N_27167,N_26369,N_26117);
nand U27168 (N_27168,N_26428,N_26458);
or U27169 (N_27169,N_26632,N_26794);
nor U27170 (N_27170,N_26234,N_26178);
xor U27171 (N_27171,N_26646,N_26900);
nor U27172 (N_27172,N_26025,N_26657);
xor U27173 (N_27173,N_26021,N_26163);
nor U27174 (N_27174,N_26844,N_26436);
nand U27175 (N_27175,N_26937,N_26820);
xnor U27176 (N_27176,N_26180,N_26430);
xor U27177 (N_27177,N_26792,N_26817);
or U27178 (N_27178,N_26470,N_26264);
and U27179 (N_27179,N_26667,N_26822);
xor U27180 (N_27180,N_26026,N_26192);
nand U27181 (N_27181,N_26129,N_26878);
and U27182 (N_27182,N_26269,N_26943);
or U27183 (N_27183,N_26080,N_26996);
nor U27184 (N_27184,N_26535,N_26779);
and U27185 (N_27185,N_26130,N_26695);
and U27186 (N_27186,N_26214,N_26894);
nand U27187 (N_27187,N_26815,N_26258);
nand U27188 (N_27188,N_26175,N_26010);
or U27189 (N_27189,N_26776,N_26707);
nor U27190 (N_27190,N_26456,N_26614);
xnor U27191 (N_27191,N_26289,N_26472);
nor U27192 (N_27192,N_26209,N_26752);
xnor U27193 (N_27193,N_26644,N_26564);
nand U27194 (N_27194,N_26750,N_26855);
or U27195 (N_27195,N_26375,N_26722);
nand U27196 (N_27196,N_26719,N_26319);
xnor U27197 (N_27197,N_26568,N_26052);
and U27198 (N_27198,N_26279,N_26067);
or U27199 (N_27199,N_26347,N_26935);
nand U27200 (N_27200,N_26304,N_26559);
nand U27201 (N_27201,N_26922,N_26215);
nor U27202 (N_27202,N_26566,N_26300);
nor U27203 (N_27203,N_26573,N_26956);
nor U27204 (N_27204,N_26168,N_26723);
and U27205 (N_27205,N_26631,N_26324);
nand U27206 (N_27206,N_26809,N_26204);
nand U27207 (N_27207,N_26986,N_26142);
or U27208 (N_27208,N_26259,N_26111);
or U27209 (N_27209,N_26977,N_26946);
xor U27210 (N_27210,N_26874,N_26115);
or U27211 (N_27211,N_26063,N_26000);
and U27212 (N_27212,N_26270,N_26981);
nand U27213 (N_27213,N_26678,N_26055);
nand U27214 (N_27214,N_26790,N_26594);
xnor U27215 (N_27215,N_26123,N_26297);
and U27216 (N_27216,N_26710,N_26805);
nand U27217 (N_27217,N_26545,N_26157);
and U27218 (N_27218,N_26828,N_26852);
and U27219 (N_27219,N_26429,N_26492);
and U27220 (N_27220,N_26229,N_26032);
or U27221 (N_27221,N_26840,N_26061);
or U27222 (N_27222,N_26616,N_26482);
nand U27223 (N_27223,N_26350,N_26447);
xnor U27224 (N_27224,N_26533,N_26460);
nor U27225 (N_27225,N_26797,N_26057);
nand U27226 (N_27226,N_26814,N_26124);
nand U27227 (N_27227,N_26579,N_26539);
and U27228 (N_27228,N_26316,N_26452);
nor U27229 (N_27229,N_26326,N_26351);
or U27230 (N_27230,N_26581,N_26647);
and U27231 (N_27231,N_26728,N_26149);
xnor U27232 (N_27232,N_26372,N_26242);
nand U27233 (N_27233,N_26112,N_26493);
nand U27234 (N_27234,N_26955,N_26167);
or U27235 (N_27235,N_26622,N_26743);
xnor U27236 (N_27236,N_26915,N_26333);
and U27237 (N_27237,N_26845,N_26176);
or U27238 (N_27238,N_26415,N_26516);
or U27239 (N_27239,N_26285,N_26288);
or U27240 (N_27240,N_26933,N_26877);
nand U27241 (N_27241,N_26969,N_26666);
nand U27242 (N_27242,N_26202,N_26211);
nand U27243 (N_27243,N_26243,N_26421);
nand U27244 (N_27244,N_26521,N_26451);
nand U27245 (N_27245,N_26859,N_26068);
xnor U27246 (N_27246,N_26754,N_26629);
nand U27247 (N_27247,N_26530,N_26610);
or U27248 (N_27248,N_26929,N_26757);
nor U27249 (N_27249,N_26287,N_26531);
nor U27250 (N_27250,N_26307,N_26408);
xor U27251 (N_27251,N_26450,N_26748);
or U27252 (N_27252,N_26406,N_26770);
and U27253 (N_27253,N_26365,N_26675);
xnor U27254 (N_27254,N_26366,N_26391);
or U27255 (N_27255,N_26232,N_26682);
or U27256 (N_27256,N_26737,N_26697);
nand U27257 (N_27257,N_26833,N_26663);
nor U27258 (N_27258,N_26965,N_26122);
and U27259 (N_27259,N_26600,N_26515);
nor U27260 (N_27260,N_26551,N_26905);
nand U27261 (N_27261,N_26320,N_26928);
nor U27262 (N_27262,N_26186,N_26847);
and U27263 (N_27263,N_26101,N_26690);
nor U27264 (N_27264,N_26658,N_26352);
nand U27265 (N_27265,N_26440,N_26866);
xor U27266 (N_27266,N_26595,N_26224);
nor U27267 (N_27267,N_26078,N_26802);
and U27268 (N_27268,N_26371,N_26538);
xor U27269 (N_27269,N_26725,N_26328);
nor U27270 (N_27270,N_26498,N_26871);
nand U27271 (N_27271,N_26015,N_26305);
nor U27272 (N_27272,N_26901,N_26179);
and U27273 (N_27273,N_26362,N_26789);
nor U27274 (N_27274,N_26863,N_26736);
nand U27275 (N_27275,N_26731,N_26717);
or U27276 (N_27276,N_26850,N_26856);
or U27277 (N_27277,N_26113,N_26837);
xor U27278 (N_27278,N_26886,N_26588);
and U27279 (N_27279,N_26713,N_26514);
or U27280 (N_27280,N_26357,N_26413);
or U27281 (N_27281,N_26768,N_26303);
nor U27282 (N_27282,N_26033,N_26344);
or U27283 (N_27283,N_26887,N_26196);
nor U27284 (N_27284,N_26376,N_26386);
and U27285 (N_27285,N_26029,N_26608);
or U27286 (N_27286,N_26230,N_26240);
nand U27287 (N_27287,N_26170,N_26938);
nand U27288 (N_27288,N_26448,N_26774);
and U27289 (N_27289,N_26022,N_26907);
and U27290 (N_27290,N_26011,N_26334);
xnor U27291 (N_27291,N_26541,N_26125);
xor U27292 (N_27292,N_26261,N_26040);
xnor U27293 (N_27293,N_26035,N_26836);
xnor U27294 (N_27294,N_26318,N_26072);
or U27295 (N_27295,N_26721,N_26562);
or U27296 (N_27296,N_26314,N_26634);
and U27297 (N_27297,N_26902,N_26769);
or U27298 (N_27298,N_26210,N_26685);
or U27299 (N_27299,N_26469,N_26968);
nand U27300 (N_27300,N_26093,N_26583);
and U27301 (N_27301,N_26236,N_26028);
xnor U27302 (N_27302,N_26427,N_26653);
or U27303 (N_27303,N_26596,N_26537);
xnor U27304 (N_27304,N_26701,N_26720);
and U27305 (N_27305,N_26764,N_26401);
nor U27306 (N_27306,N_26412,N_26132);
or U27307 (N_27307,N_26892,N_26927);
or U27308 (N_27308,N_26348,N_26185);
and U27309 (N_27309,N_26609,N_26434);
or U27310 (N_27310,N_26329,N_26846);
and U27311 (N_27311,N_26422,N_26390);
or U27312 (N_27312,N_26904,N_26676);
nor U27313 (N_27313,N_26854,N_26355);
xnor U27314 (N_27314,N_26309,N_26228);
xor U27315 (N_27315,N_26468,N_26669);
nor U27316 (N_27316,N_26088,N_26500);
or U27317 (N_27317,N_26138,N_26706);
nand U27318 (N_27318,N_26105,N_26191);
nor U27319 (N_27319,N_26807,N_26340);
nand U27320 (N_27320,N_26659,N_26310);
nor U27321 (N_27321,N_26763,N_26526);
nand U27322 (N_27322,N_26628,N_26166);
and U27323 (N_27323,N_26389,N_26949);
or U27324 (N_27324,N_26218,N_26181);
nor U27325 (N_27325,N_26652,N_26396);
xnor U27326 (N_27326,N_26702,N_26916);
or U27327 (N_27327,N_26756,N_26431);
nor U27328 (N_27328,N_26271,N_26999);
nor U27329 (N_27329,N_26302,N_26953);
nor U27330 (N_27330,N_26574,N_26220);
nor U27331 (N_27331,N_26195,N_26160);
and U27332 (N_27332,N_26730,N_26131);
xnor U27333 (N_27333,N_26161,N_26785);
and U27334 (N_27334,N_26829,N_26656);
nor U27335 (N_27335,N_26476,N_26982);
or U27336 (N_27336,N_26804,N_26203);
and U27337 (N_27337,N_26183,N_26618);
xnor U27338 (N_27338,N_26444,N_26051);
and U27339 (N_27339,N_26660,N_26411);
or U27340 (N_27340,N_26552,N_26453);
or U27341 (N_27341,N_26967,N_26557);
or U27342 (N_27342,N_26718,N_26037);
nor U27343 (N_27343,N_26883,N_26914);
and U27344 (N_27344,N_26467,N_26201);
xor U27345 (N_27345,N_26398,N_26247);
nor U27346 (N_27346,N_26621,N_26489);
and U27347 (N_27347,N_26891,N_26838);
nor U27348 (N_27348,N_26205,N_26642);
or U27349 (N_27349,N_26934,N_26356);
xnor U27350 (N_27350,N_26327,N_26246);
or U27351 (N_27351,N_26648,N_26835);
nor U27352 (N_27352,N_26159,N_26079);
or U27353 (N_27353,N_26373,N_26586);
nor U27354 (N_27354,N_26128,N_26044);
xor U27355 (N_27355,N_26238,N_26775);
nor U27356 (N_27356,N_26336,N_26013);
and U27357 (N_27357,N_26773,N_26911);
nand U27358 (N_27358,N_26565,N_26962);
and U27359 (N_27359,N_26936,N_26255);
xor U27360 (N_27360,N_26189,N_26603);
nor U27361 (N_27361,N_26857,N_26423);
xnor U27362 (N_27362,N_26708,N_26274);
xnor U27363 (N_27363,N_26137,N_26738);
nor U27364 (N_27364,N_26716,N_26919);
nand U27365 (N_27365,N_26680,N_26385);
and U27366 (N_27366,N_26705,N_26374);
nor U27367 (N_27367,N_26712,N_26612);
nor U27368 (N_27368,N_26244,N_26926);
or U27369 (N_27369,N_26759,N_26787);
and U27370 (N_27370,N_26225,N_26074);
or U27371 (N_27371,N_26554,N_26379);
xnor U27372 (N_27372,N_26263,N_26553);
nand U27373 (N_27373,N_26208,N_26158);
xnor U27374 (N_27374,N_26085,N_26387);
and U27375 (N_27375,N_26517,N_26023);
nor U27376 (N_27376,N_26245,N_26331);
and U27377 (N_27377,N_26104,N_26504);
or U27378 (N_27378,N_26976,N_26597);
or U27379 (N_27379,N_26860,N_26475);
or U27380 (N_27380,N_26749,N_26873);
and U27381 (N_27381,N_26353,N_26555);
xor U27382 (N_27382,N_26839,N_26679);
nand U27383 (N_27383,N_26681,N_26097);
or U27384 (N_27384,N_26182,N_26417);
nand U27385 (N_27385,N_26908,N_26024);
xor U27386 (N_27386,N_26989,N_26584);
nand U27387 (N_27387,N_26885,N_26141);
nand U27388 (N_27388,N_26687,N_26298);
nand U27389 (N_27389,N_26221,N_26443);
xnor U27390 (N_27390,N_26917,N_26486);
and U27391 (N_27391,N_26688,N_26510);
nor U27392 (N_27392,N_26438,N_26715);
or U27393 (N_27393,N_26393,N_26575);
nor U27394 (N_27394,N_26133,N_26046);
nor U27395 (N_27395,N_26536,N_26868);
and U27396 (N_27396,N_26380,N_26503);
or U27397 (N_27397,N_26762,N_26169);
nand U27398 (N_27398,N_26272,N_26156);
nand U27399 (N_27399,N_26599,N_26004);
nand U27400 (N_27400,N_26381,N_26623);
and U27401 (N_27401,N_26944,N_26187);
and U27402 (N_27402,N_26425,N_26455);
or U27403 (N_27403,N_26273,N_26342);
xor U27404 (N_27404,N_26542,N_26081);
or U27405 (N_27405,N_26601,N_26879);
nand U27406 (N_27406,N_26724,N_26941);
nor U27407 (N_27407,N_26442,N_26410);
xor U27408 (N_27408,N_26402,N_26483);
nand U27409 (N_27409,N_26341,N_26966);
and U27410 (N_27410,N_26479,N_26200);
and U27411 (N_27411,N_26661,N_26650);
xnor U27412 (N_27412,N_26558,N_26834);
or U27413 (N_27413,N_26069,N_26760);
or U27414 (N_27414,N_26090,N_26474);
and U27415 (N_27415,N_26509,N_26875);
nand U27416 (N_27416,N_26511,N_26107);
xor U27417 (N_27417,N_26457,N_26034);
xnor U27418 (N_27418,N_26519,N_26761);
xor U27419 (N_27419,N_26732,N_26184);
nand U27420 (N_27420,N_26283,N_26556);
nor U27421 (N_27421,N_26668,N_26973);
nor U27422 (N_27422,N_26793,N_26012);
or U27423 (N_27423,N_26745,N_26527);
or U27424 (N_27424,N_26106,N_26110);
xnor U27425 (N_27425,N_26788,N_26135);
xor U27426 (N_27426,N_26439,N_26370);
nor U27427 (N_27427,N_26241,N_26880);
xor U27428 (N_27428,N_26592,N_26477);
nor U27429 (N_27429,N_26153,N_26696);
nand U27430 (N_27430,N_26126,N_26674);
nor U27431 (N_27431,N_26109,N_26140);
xor U27432 (N_27432,N_26767,N_26783);
nor U27433 (N_27433,N_26567,N_26861);
nand U27434 (N_27434,N_26335,N_26766);
and U27435 (N_27435,N_26404,N_26733);
nand U27436 (N_27436,N_26513,N_26432);
or U27437 (N_27437,N_26048,N_26590);
or U27438 (N_27438,N_26991,N_26116);
xor U27439 (N_27439,N_26301,N_26487);
or U27440 (N_27440,N_26282,N_26714);
nor U27441 (N_27441,N_26213,N_26382);
nor U27442 (N_27442,N_26146,N_26686);
nand U27443 (N_27443,N_26086,N_26605);
nor U27444 (N_27444,N_26059,N_26625);
nand U27445 (N_27445,N_26311,N_26930);
and U27446 (N_27446,N_26786,N_26280);
or U27447 (N_27447,N_26816,N_26360);
and U27448 (N_27448,N_26619,N_26684);
or U27449 (N_27449,N_26741,N_26058);
nor U27450 (N_27450,N_26235,N_26471);
and U27451 (N_27451,N_26703,N_26119);
or U27452 (N_27452,N_26673,N_26520);
or U27453 (N_27453,N_26639,N_26617);
and U27454 (N_27454,N_26198,N_26257);
nand U27455 (N_27455,N_26649,N_26589);
and U27456 (N_27456,N_26323,N_26212);
or U27457 (N_27457,N_26796,N_26699);
or U27458 (N_27458,N_26092,N_26755);
nor U27459 (N_27459,N_26462,N_26062);
xnor U27460 (N_27460,N_26070,N_26952);
xor U27461 (N_27461,N_26602,N_26570);
nand U27462 (N_27462,N_26403,N_26226);
and U27463 (N_27463,N_26312,N_26278);
and U27464 (N_27464,N_26694,N_26611);
nand U27465 (N_27465,N_26005,N_26100);
xnor U27466 (N_27466,N_26560,N_26358);
nand U27467 (N_27467,N_26291,N_26550);
xnor U27468 (N_27468,N_26134,N_26803);
nand U27469 (N_27469,N_26222,N_26377);
xnor U27470 (N_27470,N_26076,N_26744);
or U27471 (N_27471,N_26578,N_26150);
nor U27472 (N_27472,N_26753,N_26758);
nor U27473 (N_27473,N_26577,N_26670);
or U27474 (N_27474,N_26643,N_26154);
xor U27475 (N_27475,N_26139,N_26830);
nor U27476 (N_27476,N_26332,N_26540);
xnor U27477 (N_27477,N_26354,N_26502);
nor U27478 (N_27478,N_26729,N_26249);
nor U27479 (N_27479,N_26985,N_26524);
xor U27480 (N_27480,N_26691,N_26071);
or U27481 (N_27481,N_26806,N_26711);
and U27482 (N_27482,N_26910,N_26961);
or U27483 (N_27483,N_26984,N_26306);
and U27484 (N_27484,N_26286,N_26947);
or U27485 (N_27485,N_26818,N_26488);
or U27486 (N_27486,N_26256,N_26876);
and U27487 (N_27487,N_26066,N_26239);
nand U27488 (N_27488,N_26795,N_26641);
or U27489 (N_27489,N_26903,N_26091);
nor U27490 (N_27490,N_26127,N_26920);
and U27491 (N_27491,N_26546,N_26587);
nor U27492 (N_27492,N_26613,N_26899);
nand U27493 (N_27493,N_26821,N_26216);
and U27494 (N_27494,N_26948,N_26683);
xnor U27495 (N_27495,N_26407,N_26295);
and U27496 (N_27496,N_26742,N_26446);
or U27497 (N_27497,N_26508,N_26102);
nand U27498 (N_27498,N_26120,N_26626);
nand U27499 (N_27499,N_26155,N_26924);
and U27500 (N_27500,N_26206,N_26543);
nor U27501 (N_27501,N_26605,N_26571);
or U27502 (N_27502,N_26801,N_26482);
nand U27503 (N_27503,N_26381,N_26634);
and U27504 (N_27504,N_26447,N_26750);
and U27505 (N_27505,N_26538,N_26353);
nand U27506 (N_27506,N_26975,N_26010);
nor U27507 (N_27507,N_26554,N_26954);
nor U27508 (N_27508,N_26622,N_26385);
or U27509 (N_27509,N_26717,N_26513);
nand U27510 (N_27510,N_26440,N_26790);
and U27511 (N_27511,N_26314,N_26779);
or U27512 (N_27512,N_26658,N_26842);
or U27513 (N_27513,N_26712,N_26160);
or U27514 (N_27514,N_26854,N_26220);
and U27515 (N_27515,N_26727,N_26710);
or U27516 (N_27516,N_26452,N_26646);
nor U27517 (N_27517,N_26486,N_26551);
nand U27518 (N_27518,N_26733,N_26973);
xor U27519 (N_27519,N_26122,N_26483);
nor U27520 (N_27520,N_26709,N_26728);
and U27521 (N_27521,N_26800,N_26896);
nand U27522 (N_27522,N_26040,N_26475);
or U27523 (N_27523,N_26421,N_26843);
xnor U27524 (N_27524,N_26162,N_26366);
or U27525 (N_27525,N_26556,N_26133);
nand U27526 (N_27526,N_26670,N_26048);
and U27527 (N_27527,N_26470,N_26867);
or U27528 (N_27528,N_26847,N_26126);
and U27529 (N_27529,N_26613,N_26809);
nor U27530 (N_27530,N_26575,N_26853);
xor U27531 (N_27531,N_26832,N_26424);
or U27532 (N_27532,N_26448,N_26603);
and U27533 (N_27533,N_26871,N_26882);
and U27534 (N_27534,N_26501,N_26517);
nor U27535 (N_27535,N_26097,N_26600);
and U27536 (N_27536,N_26555,N_26941);
xnor U27537 (N_27537,N_26170,N_26913);
and U27538 (N_27538,N_26859,N_26780);
and U27539 (N_27539,N_26959,N_26081);
xnor U27540 (N_27540,N_26032,N_26627);
and U27541 (N_27541,N_26453,N_26332);
nand U27542 (N_27542,N_26756,N_26588);
nor U27543 (N_27543,N_26148,N_26110);
or U27544 (N_27544,N_26462,N_26278);
xor U27545 (N_27545,N_26214,N_26686);
nand U27546 (N_27546,N_26234,N_26737);
xor U27547 (N_27547,N_26971,N_26970);
nand U27548 (N_27548,N_26389,N_26669);
or U27549 (N_27549,N_26079,N_26648);
nand U27550 (N_27550,N_26290,N_26949);
xnor U27551 (N_27551,N_26051,N_26100);
nor U27552 (N_27552,N_26197,N_26411);
nand U27553 (N_27553,N_26250,N_26101);
nor U27554 (N_27554,N_26911,N_26393);
nand U27555 (N_27555,N_26502,N_26145);
nand U27556 (N_27556,N_26638,N_26620);
xor U27557 (N_27557,N_26895,N_26469);
xnor U27558 (N_27558,N_26658,N_26851);
xnor U27559 (N_27559,N_26094,N_26639);
xnor U27560 (N_27560,N_26946,N_26357);
and U27561 (N_27561,N_26016,N_26579);
nor U27562 (N_27562,N_26077,N_26788);
xor U27563 (N_27563,N_26879,N_26444);
nor U27564 (N_27564,N_26982,N_26536);
nor U27565 (N_27565,N_26475,N_26324);
or U27566 (N_27566,N_26996,N_26237);
or U27567 (N_27567,N_26545,N_26368);
and U27568 (N_27568,N_26632,N_26864);
or U27569 (N_27569,N_26654,N_26901);
xor U27570 (N_27570,N_26935,N_26115);
or U27571 (N_27571,N_26911,N_26934);
nand U27572 (N_27572,N_26088,N_26292);
and U27573 (N_27573,N_26094,N_26973);
and U27574 (N_27574,N_26443,N_26652);
xnor U27575 (N_27575,N_26039,N_26275);
nand U27576 (N_27576,N_26797,N_26554);
or U27577 (N_27577,N_26098,N_26740);
nand U27578 (N_27578,N_26466,N_26708);
nand U27579 (N_27579,N_26987,N_26806);
nand U27580 (N_27580,N_26219,N_26694);
nand U27581 (N_27581,N_26384,N_26804);
and U27582 (N_27582,N_26664,N_26258);
xnor U27583 (N_27583,N_26537,N_26109);
and U27584 (N_27584,N_26383,N_26993);
nor U27585 (N_27585,N_26510,N_26593);
xnor U27586 (N_27586,N_26654,N_26737);
or U27587 (N_27587,N_26957,N_26027);
nor U27588 (N_27588,N_26552,N_26146);
or U27589 (N_27589,N_26455,N_26466);
nor U27590 (N_27590,N_26695,N_26056);
and U27591 (N_27591,N_26968,N_26828);
or U27592 (N_27592,N_26163,N_26248);
xor U27593 (N_27593,N_26674,N_26128);
nand U27594 (N_27594,N_26522,N_26710);
xor U27595 (N_27595,N_26702,N_26347);
or U27596 (N_27596,N_26381,N_26385);
or U27597 (N_27597,N_26109,N_26359);
xnor U27598 (N_27598,N_26014,N_26460);
nand U27599 (N_27599,N_26108,N_26178);
nand U27600 (N_27600,N_26065,N_26756);
or U27601 (N_27601,N_26314,N_26121);
nand U27602 (N_27602,N_26363,N_26813);
nor U27603 (N_27603,N_26475,N_26004);
xnor U27604 (N_27604,N_26808,N_26414);
xor U27605 (N_27605,N_26827,N_26586);
or U27606 (N_27606,N_26687,N_26400);
or U27607 (N_27607,N_26884,N_26557);
nand U27608 (N_27608,N_26349,N_26754);
nor U27609 (N_27609,N_26913,N_26569);
xor U27610 (N_27610,N_26527,N_26558);
or U27611 (N_27611,N_26865,N_26524);
nor U27612 (N_27612,N_26158,N_26492);
xnor U27613 (N_27613,N_26961,N_26359);
and U27614 (N_27614,N_26747,N_26874);
or U27615 (N_27615,N_26859,N_26197);
nand U27616 (N_27616,N_26613,N_26058);
xor U27617 (N_27617,N_26783,N_26958);
nand U27618 (N_27618,N_26122,N_26989);
nand U27619 (N_27619,N_26566,N_26273);
or U27620 (N_27620,N_26958,N_26589);
nor U27621 (N_27621,N_26993,N_26949);
and U27622 (N_27622,N_26883,N_26270);
and U27623 (N_27623,N_26276,N_26171);
or U27624 (N_27624,N_26644,N_26685);
nor U27625 (N_27625,N_26266,N_26289);
xnor U27626 (N_27626,N_26899,N_26477);
and U27627 (N_27627,N_26584,N_26531);
nor U27628 (N_27628,N_26437,N_26328);
or U27629 (N_27629,N_26442,N_26780);
xnor U27630 (N_27630,N_26583,N_26198);
or U27631 (N_27631,N_26048,N_26024);
nand U27632 (N_27632,N_26340,N_26691);
nor U27633 (N_27633,N_26833,N_26518);
nand U27634 (N_27634,N_26546,N_26991);
nor U27635 (N_27635,N_26730,N_26208);
nand U27636 (N_27636,N_26339,N_26955);
xor U27637 (N_27637,N_26298,N_26436);
and U27638 (N_27638,N_26177,N_26576);
xnor U27639 (N_27639,N_26931,N_26726);
nor U27640 (N_27640,N_26016,N_26502);
xnor U27641 (N_27641,N_26016,N_26166);
or U27642 (N_27642,N_26203,N_26049);
and U27643 (N_27643,N_26343,N_26024);
nor U27644 (N_27644,N_26001,N_26009);
nand U27645 (N_27645,N_26970,N_26557);
nand U27646 (N_27646,N_26792,N_26658);
nand U27647 (N_27647,N_26762,N_26121);
nor U27648 (N_27648,N_26187,N_26572);
and U27649 (N_27649,N_26149,N_26704);
and U27650 (N_27650,N_26619,N_26164);
nand U27651 (N_27651,N_26278,N_26786);
and U27652 (N_27652,N_26124,N_26025);
xor U27653 (N_27653,N_26886,N_26973);
or U27654 (N_27654,N_26615,N_26205);
and U27655 (N_27655,N_26325,N_26051);
nor U27656 (N_27656,N_26801,N_26579);
xor U27657 (N_27657,N_26661,N_26332);
or U27658 (N_27658,N_26431,N_26884);
xor U27659 (N_27659,N_26027,N_26528);
and U27660 (N_27660,N_26928,N_26390);
and U27661 (N_27661,N_26480,N_26143);
nor U27662 (N_27662,N_26052,N_26704);
nor U27663 (N_27663,N_26257,N_26154);
or U27664 (N_27664,N_26973,N_26735);
nor U27665 (N_27665,N_26581,N_26717);
and U27666 (N_27666,N_26214,N_26714);
nand U27667 (N_27667,N_26314,N_26089);
and U27668 (N_27668,N_26325,N_26601);
and U27669 (N_27669,N_26795,N_26949);
nor U27670 (N_27670,N_26991,N_26874);
nor U27671 (N_27671,N_26249,N_26996);
or U27672 (N_27672,N_26539,N_26761);
or U27673 (N_27673,N_26516,N_26679);
and U27674 (N_27674,N_26311,N_26965);
nor U27675 (N_27675,N_26440,N_26678);
xor U27676 (N_27676,N_26739,N_26115);
nand U27677 (N_27677,N_26400,N_26398);
or U27678 (N_27678,N_26267,N_26742);
nand U27679 (N_27679,N_26043,N_26468);
or U27680 (N_27680,N_26961,N_26458);
nor U27681 (N_27681,N_26532,N_26960);
and U27682 (N_27682,N_26758,N_26738);
or U27683 (N_27683,N_26252,N_26328);
nor U27684 (N_27684,N_26050,N_26942);
and U27685 (N_27685,N_26075,N_26281);
or U27686 (N_27686,N_26736,N_26183);
nand U27687 (N_27687,N_26146,N_26405);
or U27688 (N_27688,N_26894,N_26743);
xor U27689 (N_27689,N_26830,N_26328);
and U27690 (N_27690,N_26714,N_26350);
and U27691 (N_27691,N_26429,N_26487);
nand U27692 (N_27692,N_26293,N_26977);
nor U27693 (N_27693,N_26835,N_26361);
or U27694 (N_27694,N_26115,N_26718);
and U27695 (N_27695,N_26745,N_26024);
or U27696 (N_27696,N_26329,N_26187);
or U27697 (N_27697,N_26007,N_26816);
xnor U27698 (N_27698,N_26210,N_26771);
and U27699 (N_27699,N_26326,N_26480);
xnor U27700 (N_27700,N_26310,N_26266);
or U27701 (N_27701,N_26606,N_26645);
xnor U27702 (N_27702,N_26674,N_26016);
and U27703 (N_27703,N_26622,N_26442);
nor U27704 (N_27704,N_26369,N_26424);
or U27705 (N_27705,N_26429,N_26716);
nand U27706 (N_27706,N_26942,N_26178);
and U27707 (N_27707,N_26772,N_26829);
nand U27708 (N_27708,N_26794,N_26558);
nand U27709 (N_27709,N_26638,N_26737);
and U27710 (N_27710,N_26145,N_26938);
nor U27711 (N_27711,N_26656,N_26465);
nand U27712 (N_27712,N_26188,N_26139);
xor U27713 (N_27713,N_26445,N_26306);
xor U27714 (N_27714,N_26521,N_26969);
nor U27715 (N_27715,N_26074,N_26548);
nor U27716 (N_27716,N_26412,N_26030);
or U27717 (N_27717,N_26898,N_26113);
xnor U27718 (N_27718,N_26030,N_26874);
nand U27719 (N_27719,N_26759,N_26309);
or U27720 (N_27720,N_26165,N_26301);
nand U27721 (N_27721,N_26350,N_26594);
nor U27722 (N_27722,N_26209,N_26581);
and U27723 (N_27723,N_26241,N_26685);
xnor U27724 (N_27724,N_26515,N_26932);
nand U27725 (N_27725,N_26637,N_26524);
xor U27726 (N_27726,N_26983,N_26745);
xnor U27727 (N_27727,N_26103,N_26325);
and U27728 (N_27728,N_26527,N_26172);
nor U27729 (N_27729,N_26541,N_26180);
nand U27730 (N_27730,N_26375,N_26308);
and U27731 (N_27731,N_26835,N_26692);
xnor U27732 (N_27732,N_26625,N_26905);
xnor U27733 (N_27733,N_26096,N_26735);
and U27734 (N_27734,N_26948,N_26266);
xor U27735 (N_27735,N_26229,N_26935);
or U27736 (N_27736,N_26328,N_26671);
and U27737 (N_27737,N_26720,N_26814);
and U27738 (N_27738,N_26132,N_26778);
nor U27739 (N_27739,N_26630,N_26438);
xnor U27740 (N_27740,N_26487,N_26988);
or U27741 (N_27741,N_26000,N_26487);
xnor U27742 (N_27742,N_26684,N_26065);
nor U27743 (N_27743,N_26177,N_26925);
or U27744 (N_27744,N_26952,N_26046);
or U27745 (N_27745,N_26762,N_26997);
nor U27746 (N_27746,N_26176,N_26372);
or U27747 (N_27747,N_26453,N_26865);
nor U27748 (N_27748,N_26942,N_26662);
or U27749 (N_27749,N_26107,N_26119);
nand U27750 (N_27750,N_26750,N_26291);
and U27751 (N_27751,N_26610,N_26859);
nor U27752 (N_27752,N_26908,N_26693);
or U27753 (N_27753,N_26403,N_26864);
or U27754 (N_27754,N_26370,N_26767);
and U27755 (N_27755,N_26483,N_26960);
or U27756 (N_27756,N_26083,N_26544);
nor U27757 (N_27757,N_26212,N_26674);
nand U27758 (N_27758,N_26051,N_26657);
nor U27759 (N_27759,N_26940,N_26420);
or U27760 (N_27760,N_26711,N_26090);
xnor U27761 (N_27761,N_26268,N_26950);
xnor U27762 (N_27762,N_26514,N_26570);
xor U27763 (N_27763,N_26110,N_26368);
nand U27764 (N_27764,N_26502,N_26819);
nand U27765 (N_27765,N_26827,N_26996);
xnor U27766 (N_27766,N_26112,N_26012);
and U27767 (N_27767,N_26178,N_26240);
nand U27768 (N_27768,N_26305,N_26435);
nor U27769 (N_27769,N_26815,N_26029);
nand U27770 (N_27770,N_26399,N_26816);
or U27771 (N_27771,N_26929,N_26976);
and U27772 (N_27772,N_26324,N_26778);
or U27773 (N_27773,N_26201,N_26081);
xnor U27774 (N_27774,N_26164,N_26191);
or U27775 (N_27775,N_26037,N_26875);
and U27776 (N_27776,N_26642,N_26922);
xnor U27777 (N_27777,N_26574,N_26987);
or U27778 (N_27778,N_26920,N_26975);
nand U27779 (N_27779,N_26461,N_26546);
and U27780 (N_27780,N_26559,N_26589);
and U27781 (N_27781,N_26103,N_26223);
nand U27782 (N_27782,N_26380,N_26471);
and U27783 (N_27783,N_26419,N_26735);
nand U27784 (N_27784,N_26293,N_26889);
xor U27785 (N_27785,N_26628,N_26044);
nor U27786 (N_27786,N_26918,N_26533);
xnor U27787 (N_27787,N_26245,N_26156);
nand U27788 (N_27788,N_26394,N_26517);
nand U27789 (N_27789,N_26125,N_26800);
nor U27790 (N_27790,N_26556,N_26538);
or U27791 (N_27791,N_26798,N_26523);
nor U27792 (N_27792,N_26164,N_26438);
xor U27793 (N_27793,N_26135,N_26987);
xor U27794 (N_27794,N_26325,N_26529);
xor U27795 (N_27795,N_26895,N_26417);
xor U27796 (N_27796,N_26228,N_26163);
xor U27797 (N_27797,N_26883,N_26676);
nor U27798 (N_27798,N_26196,N_26808);
nor U27799 (N_27799,N_26256,N_26927);
nand U27800 (N_27800,N_26648,N_26159);
xnor U27801 (N_27801,N_26082,N_26794);
nor U27802 (N_27802,N_26375,N_26221);
and U27803 (N_27803,N_26853,N_26078);
and U27804 (N_27804,N_26683,N_26309);
nor U27805 (N_27805,N_26995,N_26373);
or U27806 (N_27806,N_26279,N_26986);
nor U27807 (N_27807,N_26195,N_26497);
or U27808 (N_27808,N_26917,N_26436);
or U27809 (N_27809,N_26915,N_26581);
nand U27810 (N_27810,N_26385,N_26638);
or U27811 (N_27811,N_26509,N_26098);
xor U27812 (N_27812,N_26334,N_26611);
or U27813 (N_27813,N_26301,N_26011);
nor U27814 (N_27814,N_26284,N_26879);
nor U27815 (N_27815,N_26411,N_26198);
and U27816 (N_27816,N_26799,N_26368);
nand U27817 (N_27817,N_26363,N_26507);
and U27818 (N_27818,N_26316,N_26300);
and U27819 (N_27819,N_26977,N_26621);
and U27820 (N_27820,N_26159,N_26607);
nand U27821 (N_27821,N_26103,N_26751);
nand U27822 (N_27822,N_26527,N_26733);
xnor U27823 (N_27823,N_26889,N_26968);
xor U27824 (N_27824,N_26484,N_26553);
nand U27825 (N_27825,N_26115,N_26847);
nand U27826 (N_27826,N_26217,N_26539);
and U27827 (N_27827,N_26549,N_26065);
and U27828 (N_27828,N_26453,N_26723);
and U27829 (N_27829,N_26685,N_26206);
nor U27830 (N_27830,N_26708,N_26425);
nor U27831 (N_27831,N_26629,N_26899);
nand U27832 (N_27832,N_26008,N_26951);
nor U27833 (N_27833,N_26680,N_26740);
nor U27834 (N_27834,N_26630,N_26820);
or U27835 (N_27835,N_26565,N_26235);
xnor U27836 (N_27836,N_26710,N_26783);
nor U27837 (N_27837,N_26150,N_26035);
or U27838 (N_27838,N_26695,N_26190);
nand U27839 (N_27839,N_26946,N_26345);
and U27840 (N_27840,N_26235,N_26768);
or U27841 (N_27841,N_26534,N_26313);
or U27842 (N_27842,N_26536,N_26128);
nor U27843 (N_27843,N_26797,N_26880);
xor U27844 (N_27844,N_26053,N_26000);
xor U27845 (N_27845,N_26634,N_26484);
and U27846 (N_27846,N_26546,N_26650);
nor U27847 (N_27847,N_26679,N_26774);
xnor U27848 (N_27848,N_26847,N_26254);
or U27849 (N_27849,N_26885,N_26144);
nor U27850 (N_27850,N_26190,N_26209);
nor U27851 (N_27851,N_26187,N_26052);
or U27852 (N_27852,N_26043,N_26021);
and U27853 (N_27853,N_26948,N_26098);
nand U27854 (N_27854,N_26765,N_26058);
or U27855 (N_27855,N_26679,N_26472);
nand U27856 (N_27856,N_26279,N_26089);
xnor U27857 (N_27857,N_26383,N_26667);
nor U27858 (N_27858,N_26161,N_26232);
nor U27859 (N_27859,N_26640,N_26372);
nand U27860 (N_27860,N_26223,N_26137);
or U27861 (N_27861,N_26045,N_26758);
nand U27862 (N_27862,N_26842,N_26123);
xnor U27863 (N_27863,N_26190,N_26120);
nor U27864 (N_27864,N_26520,N_26804);
nand U27865 (N_27865,N_26989,N_26704);
and U27866 (N_27866,N_26686,N_26175);
nand U27867 (N_27867,N_26115,N_26661);
or U27868 (N_27868,N_26431,N_26921);
or U27869 (N_27869,N_26675,N_26583);
xnor U27870 (N_27870,N_26923,N_26347);
nor U27871 (N_27871,N_26032,N_26061);
nor U27872 (N_27872,N_26103,N_26557);
or U27873 (N_27873,N_26576,N_26071);
nand U27874 (N_27874,N_26630,N_26187);
xor U27875 (N_27875,N_26566,N_26744);
and U27876 (N_27876,N_26469,N_26364);
or U27877 (N_27877,N_26150,N_26017);
nor U27878 (N_27878,N_26971,N_26884);
or U27879 (N_27879,N_26699,N_26769);
nor U27880 (N_27880,N_26732,N_26307);
or U27881 (N_27881,N_26758,N_26219);
nor U27882 (N_27882,N_26101,N_26872);
nand U27883 (N_27883,N_26882,N_26233);
xor U27884 (N_27884,N_26153,N_26811);
and U27885 (N_27885,N_26702,N_26994);
nor U27886 (N_27886,N_26493,N_26528);
nor U27887 (N_27887,N_26001,N_26582);
nor U27888 (N_27888,N_26593,N_26700);
and U27889 (N_27889,N_26548,N_26957);
nand U27890 (N_27890,N_26766,N_26049);
and U27891 (N_27891,N_26464,N_26065);
xor U27892 (N_27892,N_26863,N_26506);
nor U27893 (N_27893,N_26982,N_26983);
nor U27894 (N_27894,N_26137,N_26678);
and U27895 (N_27895,N_26624,N_26606);
xnor U27896 (N_27896,N_26680,N_26271);
xnor U27897 (N_27897,N_26991,N_26814);
nor U27898 (N_27898,N_26300,N_26687);
xor U27899 (N_27899,N_26141,N_26907);
and U27900 (N_27900,N_26567,N_26686);
nor U27901 (N_27901,N_26711,N_26634);
xor U27902 (N_27902,N_26181,N_26109);
and U27903 (N_27903,N_26633,N_26528);
nand U27904 (N_27904,N_26388,N_26102);
or U27905 (N_27905,N_26329,N_26422);
nand U27906 (N_27906,N_26666,N_26972);
or U27907 (N_27907,N_26684,N_26193);
nand U27908 (N_27908,N_26319,N_26705);
nand U27909 (N_27909,N_26715,N_26994);
xor U27910 (N_27910,N_26555,N_26601);
or U27911 (N_27911,N_26126,N_26407);
xor U27912 (N_27912,N_26889,N_26687);
xor U27913 (N_27913,N_26851,N_26674);
and U27914 (N_27914,N_26125,N_26667);
or U27915 (N_27915,N_26706,N_26589);
and U27916 (N_27916,N_26324,N_26137);
nor U27917 (N_27917,N_26379,N_26360);
and U27918 (N_27918,N_26768,N_26358);
xor U27919 (N_27919,N_26244,N_26791);
xor U27920 (N_27920,N_26941,N_26096);
nand U27921 (N_27921,N_26151,N_26212);
nor U27922 (N_27922,N_26987,N_26116);
xor U27923 (N_27923,N_26620,N_26323);
nor U27924 (N_27924,N_26939,N_26858);
and U27925 (N_27925,N_26822,N_26701);
nand U27926 (N_27926,N_26013,N_26358);
and U27927 (N_27927,N_26447,N_26435);
and U27928 (N_27928,N_26663,N_26049);
nand U27929 (N_27929,N_26398,N_26760);
xnor U27930 (N_27930,N_26189,N_26448);
nor U27931 (N_27931,N_26054,N_26357);
nor U27932 (N_27932,N_26727,N_26888);
nand U27933 (N_27933,N_26337,N_26971);
and U27934 (N_27934,N_26928,N_26735);
xnor U27935 (N_27935,N_26781,N_26494);
and U27936 (N_27936,N_26926,N_26429);
or U27937 (N_27937,N_26345,N_26033);
nand U27938 (N_27938,N_26202,N_26499);
nand U27939 (N_27939,N_26692,N_26120);
nor U27940 (N_27940,N_26426,N_26695);
nand U27941 (N_27941,N_26671,N_26725);
or U27942 (N_27942,N_26374,N_26677);
and U27943 (N_27943,N_26857,N_26552);
and U27944 (N_27944,N_26331,N_26822);
and U27945 (N_27945,N_26660,N_26500);
and U27946 (N_27946,N_26367,N_26174);
xor U27947 (N_27947,N_26893,N_26180);
and U27948 (N_27948,N_26371,N_26576);
xnor U27949 (N_27949,N_26136,N_26893);
nand U27950 (N_27950,N_26379,N_26884);
xor U27951 (N_27951,N_26031,N_26093);
nand U27952 (N_27952,N_26499,N_26514);
nor U27953 (N_27953,N_26627,N_26231);
nand U27954 (N_27954,N_26356,N_26754);
or U27955 (N_27955,N_26345,N_26331);
nor U27956 (N_27956,N_26008,N_26253);
xor U27957 (N_27957,N_26756,N_26464);
nor U27958 (N_27958,N_26020,N_26675);
or U27959 (N_27959,N_26671,N_26705);
xnor U27960 (N_27960,N_26935,N_26252);
nand U27961 (N_27961,N_26397,N_26848);
nor U27962 (N_27962,N_26546,N_26574);
or U27963 (N_27963,N_26225,N_26537);
xor U27964 (N_27964,N_26613,N_26850);
or U27965 (N_27965,N_26589,N_26835);
nand U27966 (N_27966,N_26558,N_26302);
nand U27967 (N_27967,N_26419,N_26307);
nand U27968 (N_27968,N_26617,N_26387);
nand U27969 (N_27969,N_26978,N_26600);
nand U27970 (N_27970,N_26808,N_26630);
nand U27971 (N_27971,N_26643,N_26672);
and U27972 (N_27972,N_26388,N_26771);
nand U27973 (N_27973,N_26870,N_26851);
xnor U27974 (N_27974,N_26779,N_26798);
and U27975 (N_27975,N_26609,N_26181);
nand U27976 (N_27976,N_26387,N_26824);
nand U27977 (N_27977,N_26523,N_26284);
or U27978 (N_27978,N_26110,N_26553);
nor U27979 (N_27979,N_26826,N_26121);
nor U27980 (N_27980,N_26774,N_26226);
and U27981 (N_27981,N_26553,N_26901);
nor U27982 (N_27982,N_26542,N_26782);
xor U27983 (N_27983,N_26558,N_26218);
nand U27984 (N_27984,N_26790,N_26653);
xnor U27985 (N_27985,N_26904,N_26539);
nand U27986 (N_27986,N_26835,N_26127);
and U27987 (N_27987,N_26999,N_26055);
nand U27988 (N_27988,N_26936,N_26729);
nor U27989 (N_27989,N_26604,N_26112);
nor U27990 (N_27990,N_26854,N_26781);
or U27991 (N_27991,N_26576,N_26650);
nor U27992 (N_27992,N_26837,N_26975);
and U27993 (N_27993,N_26626,N_26541);
or U27994 (N_27994,N_26214,N_26874);
xor U27995 (N_27995,N_26587,N_26702);
or U27996 (N_27996,N_26695,N_26358);
nor U27997 (N_27997,N_26053,N_26698);
or U27998 (N_27998,N_26687,N_26838);
nand U27999 (N_27999,N_26807,N_26649);
nor U28000 (N_28000,N_27939,N_27045);
xor U28001 (N_28001,N_27798,N_27853);
nand U28002 (N_28002,N_27890,N_27543);
nand U28003 (N_28003,N_27788,N_27781);
and U28004 (N_28004,N_27176,N_27080);
or U28005 (N_28005,N_27714,N_27018);
xnor U28006 (N_28006,N_27331,N_27048);
nand U28007 (N_28007,N_27932,N_27568);
xnor U28008 (N_28008,N_27907,N_27068);
nand U28009 (N_28009,N_27782,N_27883);
xnor U28010 (N_28010,N_27409,N_27200);
nor U28011 (N_28011,N_27854,N_27450);
or U28012 (N_28012,N_27737,N_27953);
or U28013 (N_28013,N_27758,N_27575);
nor U28014 (N_28014,N_27770,N_27909);
and U28015 (N_28015,N_27712,N_27401);
nor U28016 (N_28016,N_27898,N_27221);
and U28017 (N_28017,N_27374,N_27121);
and U28018 (N_28018,N_27003,N_27505);
nand U28019 (N_28019,N_27387,N_27475);
nand U28020 (N_28020,N_27943,N_27369);
and U28021 (N_28021,N_27704,N_27750);
or U28022 (N_28022,N_27654,N_27915);
and U28023 (N_28023,N_27825,N_27922);
nand U28024 (N_28024,N_27168,N_27302);
and U28025 (N_28025,N_27926,N_27095);
or U28026 (N_28026,N_27655,N_27673);
xor U28027 (N_28027,N_27887,N_27545);
nand U28028 (N_28028,N_27860,N_27267);
nand U28029 (N_28029,N_27604,N_27960);
or U28030 (N_28030,N_27482,N_27456);
xor U28031 (N_28031,N_27611,N_27992);
xor U28032 (N_28032,N_27415,N_27993);
and U28033 (N_28033,N_27495,N_27977);
xnor U28034 (N_28034,N_27928,N_27541);
xnor U28035 (N_28035,N_27754,N_27265);
nand U28036 (N_28036,N_27914,N_27317);
xor U28037 (N_28037,N_27372,N_27343);
and U28038 (N_28038,N_27063,N_27247);
nand U28039 (N_28039,N_27175,N_27715);
and U28040 (N_28040,N_27602,N_27612);
xnor U28041 (N_28041,N_27817,N_27732);
or U28042 (N_28042,N_27674,N_27620);
or U28043 (N_28043,N_27901,N_27531);
nand U28044 (N_28044,N_27766,N_27806);
or U28045 (N_28045,N_27157,N_27085);
xor U28046 (N_28046,N_27234,N_27272);
and U28047 (N_28047,N_27945,N_27038);
or U28048 (N_28048,N_27181,N_27039);
nand U28049 (N_28049,N_27882,N_27739);
nand U28050 (N_28050,N_27240,N_27903);
and U28051 (N_28051,N_27174,N_27357);
nand U28052 (N_28052,N_27985,N_27550);
and U28053 (N_28053,N_27815,N_27949);
and U28054 (N_28054,N_27707,N_27869);
nor U28055 (N_28055,N_27561,N_27078);
nor U28056 (N_28056,N_27161,N_27461);
xnor U28057 (N_28057,N_27666,N_27278);
xnor U28058 (N_28058,N_27609,N_27800);
nand U28059 (N_28059,N_27678,N_27165);
xor U28060 (N_28060,N_27173,N_27919);
and U28061 (N_28061,N_27978,N_27785);
nor U28062 (N_28062,N_27148,N_27041);
or U28063 (N_28063,N_27417,N_27700);
or U28064 (N_28064,N_27558,N_27793);
and U28065 (N_28065,N_27208,N_27976);
nand U28066 (N_28066,N_27347,N_27320);
nor U28067 (N_28067,N_27486,N_27341);
nor U28068 (N_28068,N_27649,N_27044);
and U28069 (N_28069,N_27728,N_27017);
xor U28070 (N_28070,N_27287,N_27182);
nand U28071 (N_28071,N_27462,N_27711);
or U28072 (N_28072,N_27996,N_27507);
xor U28073 (N_28073,N_27002,N_27937);
or U28074 (N_28074,N_27281,N_27745);
nor U28075 (N_28075,N_27713,N_27315);
xor U28076 (N_28076,N_27878,N_27523);
and U28077 (N_28077,N_27593,N_27941);
nand U28078 (N_28078,N_27336,N_27553);
and U28079 (N_28079,N_27662,N_27004);
or U28080 (N_28080,N_27251,N_27185);
or U28081 (N_28081,N_27399,N_27016);
or U28082 (N_28082,N_27438,N_27188);
nor U28083 (N_28083,N_27963,N_27282);
nand U28084 (N_28084,N_27015,N_27013);
xor U28085 (N_28085,N_27073,N_27660);
nor U28086 (N_28086,N_27093,N_27010);
and U28087 (N_28087,N_27625,N_27327);
and U28088 (N_28088,N_27260,N_27413);
or U28089 (N_28089,N_27857,N_27856);
and U28090 (N_28090,N_27082,N_27615);
nor U28091 (N_28091,N_27009,N_27502);
nand U28092 (N_28092,N_27385,N_27508);
or U28093 (N_28093,N_27458,N_27355);
nand U28094 (N_28094,N_27443,N_27418);
and U28095 (N_28095,N_27743,N_27844);
xnor U28096 (N_28096,N_27735,N_27218);
or U28097 (N_28097,N_27293,N_27171);
nor U28098 (N_28098,N_27153,N_27988);
nand U28099 (N_28099,N_27052,N_27307);
or U28100 (N_28100,N_27868,N_27872);
and U28101 (N_28101,N_27366,N_27407);
and U28102 (N_28102,N_27742,N_27924);
or U28103 (N_28103,N_27566,N_27079);
or U28104 (N_28104,N_27757,N_27353);
nor U28105 (N_28105,N_27773,N_27744);
nand U28106 (N_28106,N_27452,N_27334);
and U28107 (N_28107,N_27330,N_27771);
xor U28108 (N_28108,N_27422,N_27416);
nor U28109 (N_28109,N_27227,N_27464);
xnor U28110 (N_28110,N_27472,N_27727);
xor U28111 (N_28111,N_27821,N_27720);
or U28112 (N_28112,N_27528,N_27444);
and U28113 (N_28113,N_27177,N_27668);
nand U28114 (N_28114,N_27491,N_27554);
nand U28115 (N_28115,N_27709,N_27775);
or U28116 (N_28116,N_27573,N_27367);
nand U28117 (N_28117,N_27511,N_27803);
xor U28118 (N_28118,N_27540,N_27467);
xor U28119 (N_28119,N_27364,N_27269);
or U28120 (N_28120,N_27768,N_27042);
or U28121 (N_28121,N_27968,N_27314);
nor U28122 (N_28122,N_27998,N_27235);
and U28123 (N_28123,N_27751,N_27930);
nand U28124 (N_28124,N_27101,N_27537);
and U28125 (N_28125,N_27586,N_27627);
or U28126 (N_28126,N_27647,N_27783);
and U28127 (N_28127,N_27091,N_27884);
or U28128 (N_28128,N_27279,N_27097);
and U28129 (N_28129,N_27466,N_27498);
or U28130 (N_28130,N_27510,N_27397);
nand U28131 (N_28131,N_27517,N_27414);
nand U28132 (N_28132,N_27250,N_27948);
or U28133 (N_28133,N_27769,N_27661);
nand U28134 (N_28134,N_27832,N_27274);
and U28135 (N_28135,N_27453,N_27525);
and U28136 (N_28136,N_27552,N_27628);
xnor U28137 (N_28137,N_27187,N_27618);
nor U28138 (N_28138,N_27394,N_27633);
nand U28139 (N_28139,N_27186,N_27062);
nor U28140 (N_28140,N_27970,N_27198);
xnor U28141 (N_28141,N_27889,N_27641);
xor U28142 (N_28142,N_27130,N_27156);
nor U28143 (N_28143,N_27827,N_27858);
nand U28144 (N_28144,N_27956,N_27258);
or U28145 (N_28145,N_27448,N_27952);
or U28146 (N_28146,N_27885,N_27576);
and U28147 (N_28147,N_27131,N_27636);
xnor U28148 (N_28148,N_27296,N_27546);
and U28149 (N_28149,N_27373,N_27904);
and U28150 (N_28150,N_27690,N_27066);
nand U28151 (N_28151,N_27995,N_27057);
nand U28152 (N_28152,N_27110,N_27332);
nor U28153 (N_28153,N_27731,N_27719);
and U28154 (N_28154,N_27426,N_27835);
xnor U28155 (N_28155,N_27425,N_27925);
and U28156 (N_28156,N_27534,N_27172);
or U28157 (N_28157,N_27194,N_27337);
and U28158 (N_28158,N_27350,N_27864);
or U28159 (N_28159,N_27492,N_27434);
nor U28160 (N_28160,N_27268,N_27913);
nand U28161 (N_28161,N_27934,N_27244);
xor U28162 (N_28162,N_27624,N_27379);
xnor U28163 (N_28163,N_27684,N_27454);
nor U28164 (N_28164,N_27395,N_27894);
nand U28165 (N_28165,N_27280,N_27096);
nand U28166 (N_28166,N_27642,N_27469);
nand U28167 (N_28167,N_27441,N_27820);
nand U28168 (N_28168,N_27051,N_27643);
nand U28169 (N_28169,N_27271,N_27759);
and U28170 (N_28170,N_27430,N_27484);
nand U28171 (N_28171,N_27478,N_27532);
xnor U28172 (N_28172,N_27529,N_27402);
and U28173 (N_28173,N_27973,N_27962);
or U28174 (N_28174,N_27906,N_27329);
xnor U28175 (N_28175,N_27587,N_27762);
xnor U28176 (N_28176,N_27236,N_27111);
or U28177 (N_28177,N_27946,N_27982);
nand U28178 (N_28178,N_27286,N_27632);
or U28179 (N_28179,N_27163,N_27046);
xor U28180 (N_28180,N_27238,N_27304);
nor U28181 (N_28181,N_27435,N_27630);
xnor U28182 (N_28182,N_27513,N_27951);
nor U28183 (N_28183,N_27254,N_27622);
nor U28184 (N_28184,N_27359,N_27109);
xnor U28185 (N_28185,N_27411,N_27140);
xnor U28186 (N_28186,N_27311,N_27839);
nand U28187 (N_28187,N_27665,N_27935);
or U28188 (N_28188,N_27382,N_27623);
nand U28189 (N_28189,N_27030,N_27207);
xnor U28190 (N_28190,N_27617,N_27473);
xnor U28191 (N_28191,N_27261,N_27999);
or U28192 (N_28192,N_27072,N_27303);
and U28193 (N_28193,N_27792,N_27210);
and U28194 (N_28194,N_27734,N_27285);
or U28195 (N_28195,N_27710,N_27626);
or U28196 (N_28196,N_27445,N_27145);
xnor U28197 (N_28197,N_27862,N_27460);
nor U28198 (N_28198,N_27746,N_27001);
nand U28199 (N_28199,N_27212,N_27058);
or U28200 (N_28200,N_27309,N_27895);
nor U28201 (N_28201,N_27967,N_27432);
nand U28202 (N_28202,N_27138,N_27122);
or U28203 (N_28203,N_27392,N_27794);
or U28204 (N_28204,N_27102,N_27346);
nand U28205 (N_28205,N_27607,N_27826);
nor U28206 (N_28206,N_27160,N_27824);
xor U28207 (N_28207,N_27539,N_27169);
or U28208 (N_28208,N_27405,N_27049);
xnor U28209 (N_28209,N_27283,N_27656);
or U28210 (N_28210,N_27237,N_27075);
xor U28211 (N_28211,N_27214,N_27689);
xnor U28212 (N_28212,N_27777,N_27648);
and U28213 (N_28213,N_27503,N_27692);
or U28214 (N_28214,N_27362,N_27779);
and U28215 (N_28215,N_27500,N_27352);
nand U28216 (N_28216,N_27383,N_27390);
nand U28217 (N_28217,N_27112,N_27270);
xnor U28218 (N_28218,N_27084,N_27032);
nor U28219 (N_28219,N_27446,N_27518);
or U28220 (N_28220,N_27108,N_27089);
or U28221 (N_28221,N_27128,N_27989);
xnor U28222 (N_28222,N_27652,N_27375);
or U28223 (N_28223,N_27955,N_27809);
xor U28224 (N_28224,N_27231,N_27581);
or U28225 (N_28225,N_27664,N_27578);
nor U28226 (N_28226,N_27106,N_27598);
nor U28227 (N_28227,N_27196,N_27986);
or U28228 (N_28228,N_27780,N_27691);
or U28229 (N_28229,N_27321,N_27871);
or U28230 (N_28230,N_27548,N_27787);
nor U28231 (N_28231,N_27682,N_27899);
and U28232 (N_28232,N_27892,N_27594);
and U28233 (N_28233,N_27388,N_27468);
or U28234 (N_28234,N_27429,N_27603);
or U28235 (N_28235,N_27905,N_27569);
nor U28236 (N_28236,N_27127,N_27216);
xor U28237 (N_28237,N_27964,N_27812);
nor U28238 (N_28238,N_27202,N_27076);
and U28239 (N_28239,N_27848,N_27813);
xor U28240 (N_28240,N_27683,N_27908);
nand U28241 (N_28241,N_27902,N_27220);
or U28242 (N_28242,N_27376,N_27893);
nor U28243 (N_28243,N_27301,N_27377);
or U28244 (N_28244,N_27933,N_27248);
and U28245 (N_28245,N_27802,N_27938);
and U28246 (N_28246,N_27556,N_27760);
nand U28247 (N_28247,N_27487,N_27339);
xor U28248 (N_28248,N_27144,N_27805);
or U28249 (N_28249,N_27671,N_27358);
nand U28250 (N_28250,N_27459,N_27465);
nor U28251 (N_28251,N_27645,N_27447);
nand U28252 (N_28252,N_27687,N_27677);
or U28253 (N_28253,N_27947,N_27319);
or U28254 (N_28254,N_27597,N_27778);
and U28255 (N_28255,N_27808,N_27288);
nor U28256 (N_28256,N_27233,N_27136);
or U28257 (N_28257,N_27991,N_27829);
nor U28258 (N_28258,N_27035,N_27873);
xnor U28259 (N_28259,N_27092,N_27669);
xor U28260 (N_28260,N_27098,N_27496);
and U28261 (N_28261,N_27463,N_27980);
nor U28262 (N_28262,N_27506,N_27940);
and U28263 (N_28263,N_27033,N_27206);
nor U28264 (N_28264,N_27349,N_27497);
nand U28265 (N_28265,N_27920,N_27555);
nor U28266 (N_28266,N_27549,N_27847);
nor U28267 (N_28267,N_27736,N_27455);
nand U28268 (N_28268,N_27114,N_27026);
and U28269 (N_28269,N_27470,N_27562);
and U28270 (N_28270,N_27036,N_27961);
xor U28271 (N_28271,N_27149,N_27326);
xor U28272 (N_28272,N_27535,N_27584);
xor U28273 (N_28273,N_27698,N_27776);
and U28274 (N_28274,N_27277,N_27954);
nand U28275 (N_28275,N_27514,N_27253);
xnor U28276 (N_28276,N_27201,N_27107);
nor U28277 (N_28277,N_27480,N_27705);
nor U28278 (N_28278,N_27542,N_27120);
nand U28279 (N_28279,N_27818,N_27983);
nand U28280 (N_28280,N_27255,N_27154);
nand U28281 (N_28281,N_27807,N_27629);
or U28282 (N_28282,N_27834,N_27313);
and U28283 (N_28283,N_27262,N_27040);
or U28284 (N_28284,N_27867,N_27512);
or U28285 (N_28285,N_27990,N_27170);
or U28286 (N_28286,N_27918,N_27393);
xor U28287 (N_28287,N_27944,N_27765);
xnor U28288 (N_28288,N_27816,N_27230);
and U28289 (N_28289,N_27583,N_27333);
or U28290 (N_28290,N_27706,N_27547);
nor U28291 (N_28291,N_27850,N_27494);
nor U28292 (N_28292,N_27229,N_27588);
and U28293 (N_28293,N_27398,N_27205);
and U28294 (N_28294,N_27067,N_27657);
or U28295 (N_28295,N_27224,N_27697);
or U28296 (N_28296,N_27384,N_27008);
xnor U28297 (N_28297,N_27142,N_27876);
and U28298 (N_28298,N_27299,N_27113);
and U28299 (N_28299,N_27410,N_27972);
xor U28300 (N_28300,N_27029,N_27158);
nand U28301 (N_28301,N_27371,N_27595);
and U28302 (N_28302,N_27166,N_27263);
nor U28303 (N_28303,N_27232,N_27191);
nor U28304 (N_28304,N_27276,N_27135);
nand U28305 (N_28305,N_27533,N_27436);
nand U28306 (N_28306,N_27476,N_27675);
nand U28307 (N_28307,N_27701,N_27099);
or U28308 (N_28308,N_27184,N_27021);
and U28309 (N_28309,N_27141,N_27911);
nor U28310 (N_28310,N_27859,N_27014);
and U28311 (N_28311,N_27761,N_27994);
or U28312 (N_28312,N_27064,N_27318);
nor U28313 (N_28313,N_27572,N_27822);
nand U28314 (N_28314,N_27381,N_27764);
or U28315 (N_28315,N_27784,N_27659);
xnor U28316 (N_28316,N_27753,N_27335);
nor U28317 (N_28317,N_27239,N_27755);
xor U28318 (N_28318,N_27223,N_27747);
nor U28319 (N_28319,N_27054,N_27152);
nor U28320 (N_28320,N_27564,N_27351);
xnor U28321 (N_28321,N_27378,N_27228);
nor U28322 (N_28322,N_27580,N_27969);
nor U28323 (N_28323,N_27348,N_27104);
xnor U28324 (N_28324,N_27047,N_27577);
nor U28325 (N_28325,N_27077,N_27891);
xor U28326 (N_28326,N_27126,N_27300);
nand U28327 (N_28327,N_27199,N_27100);
nor U28328 (N_28328,N_27427,N_27338);
nand U28329 (N_28329,N_27243,N_27959);
xor U28330 (N_28330,N_27601,N_27178);
nand U28331 (N_28331,N_27910,N_27217);
or U28332 (N_28332,N_27192,N_27193);
xnor U28333 (N_28333,N_27289,N_27471);
xor U28334 (N_28334,N_27738,N_27756);
and U28335 (N_28335,N_27290,N_27676);
nor U28336 (N_28336,N_27197,N_27143);
nand U28337 (N_28337,N_27879,N_27219);
or U28338 (N_28338,N_27493,N_27479);
xnor U28339 (N_28339,N_27846,N_27167);
nand U28340 (N_28340,N_27000,N_27565);
nor U28341 (N_28341,N_27183,N_27294);
nand U28342 (N_28342,N_27490,N_27504);
and U28343 (N_28343,N_27356,N_27195);
nor U28344 (N_28344,N_27725,N_27249);
nor U28345 (N_28345,N_27987,N_27406);
nor U28346 (N_28346,N_27519,N_27589);
nand U28347 (N_28347,N_27119,N_27722);
nor U28348 (N_28348,N_27020,N_27312);
and U28349 (N_28349,N_27437,N_27424);
or U28350 (N_28350,N_27179,N_27037);
xor U28351 (N_28351,N_27069,N_27396);
and U28352 (N_28352,N_27592,N_27801);
nand U28353 (N_28353,N_27796,N_27966);
nand U28354 (N_28354,N_27567,N_27638);
nor U28355 (N_28355,N_27866,N_27209);
xor U28356 (N_28356,N_27881,N_27726);
nor U28357 (N_28357,N_27133,N_27488);
and U28358 (N_28358,N_27342,N_27830);
nor U28359 (N_28359,N_27070,N_27551);
xor U28360 (N_28360,N_27767,N_27965);
nand U28361 (N_28361,N_27189,N_27022);
nand U28362 (N_28362,N_27386,N_27081);
or U28363 (N_28363,N_27526,N_27132);
nor U28364 (N_28364,N_27103,N_27012);
xor U28365 (N_28365,N_27521,N_27874);
xor U28366 (N_28366,N_27570,N_27646);
or U28367 (N_28367,N_27516,N_27115);
xor U28368 (N_28368,N_27354,N_27789);
and U28369 (N_28369,N_27599,N_27291);
or U28370 (N_28370,N_27631,N_27699);
nand U28371 (N_28371,N_27852,N_27440);
nor U28372 (N_28372,N_27086,N_27831);
nor U28373 (N_28373,N_27489,N_27752);
xnor U28374 (N_28374,N_27865,N_27150);
nor U28375 (N_28375,N_27616,N_27729);
xnor U28376 (N_28376,N_27688,N_27345);
and U28377 (N_28377,N_27083,N_27975);
and U28378 (N_28378,N_27074,N_27324);
nand U28379 (N_28379,N_27134,N_27538);
nor U28380 (N_28380,N_27888,N_27929);
nor U28381 (N_28381,N_27403,N_27703);
and U28382 (N_28382,N_27749,N_27368);
nor U28383 (N_28383,N_27635,N_27256);
xor U28384 (N_28384,N_27105,N_27590);
nor U28385 (N_28385,N_27716,N_27733);
and U28386 (N_28386,N_27608,N_27053);
xnor U28387 (N_28387,N_27637,N_27043);
or U28388 (N_28388,N_27028,N_27997);
or U28389 (N_28389,N_27557,N_27833);
and U28390 (N_28390,N_27912,N_27428);
and U28391 (N_28391,N_27950,N_27419);
or U28392 (N_28392,N_27527,N_27451);
or U28393 (N_28393,N_27843,N_27841);
nor U28394 (N_28394,N_27522,N_27011);
nand U28395 (N_28395,N_27060,N_27059);
xor U28396 (N_28396,N_27360,N_27563);
nor U28397 (N_28397,N_27591,N_27921);
xor U28398 (N_28398,N_27071,N_27686);
and U28399 (N_28399,N_27836,N_27306);
and U28400 (N_28400,N_27204,N_27582);
nor U28401 (N_28401,N_27804,N_27971);
nand U28402 (N_28402,N_27147,N_27389);
nor U28403 (N_28403,N_27875,N_27663);
xor U28404 (N_28404,N_27159,N_27730);
nor U28405 (N_28405,N_27571,N_27694);
nor U28406 (N_28406,N_27442,N_27006);
nand U28407 (N_28407,N_27509,N_27408);
or U28408 (N_28408,N_27241,N_27845);
nor U28409 (N_28409,N_27896,N_27958);
xor U28410 (N_28410,N_27837,N_27325);
xor U28411 (N_28411,N_27786,N_27984);
or U28412 (N_28412,N_27298,N_27087);
and U28413 (N_28413,N_27328,N_27748);
xor U28414 (N_28414,N_27880,N_27672);
nor U28415 (N_28415,N_27252,N_27257);
and U28416 (N_28416,N_27681,N_27763);
or U28417 (N_28417,N_27203,N_27931);
nor U28418 (N_28418,N_27284,N_27721);
nor U28419 (N_28419,N_27055,N_27499);
or U28420 (N_28420,N_27151,N_27667);
nand U28421 (N_28421,N_27579,N_27520);
and U28422 (N_28422,N_27606,N_27363);
and U28423 (N_28423,N_27162,N_27530);
nand U28424 (N_28424,N_27421,N_27146);
nor U28425 (N_28425,N_27790,N_27840);
or U28426 (N_28426,N_27246,N_27477);
or U28427 (N_28427,N_27025,N_27118);
nand U28428 (N_28428,N_27483,N_27155);
and U28429 (N_28429,N_27024,N_27639);
xnor U28430 (N_28430,N_27842,N_27365);
and U28431 (N_28431,N_27861,N_27619);
xor U28432 (N_28432,N_27180,N_27400);
nand U28433 (N_28433,N_27094,N_27670);
nor U28434 (N_28434,N_27129,N_27685);
and U28435 (N_28435,N_27559,N_27050);
nand U28436 (N_28436,N_27693,N_27897);
xor U28437 (N_28437,N_27774,N_27695);
or U28438 (N_28438,N_27264,N_27596);
or U28439 (N_28439,N_27702,N_27927);
nand U28440 (N_28440,N_27658,N_27851);
nor U28441 (N_28441,N_27226,N_27340);
xnor U28442 (N_28442,N_27870,N_27772);
or U28443 (N_28443,N_27090,N_27485);
xor U28444 (N_28444,N_27536,N_27245);
nor U28445 (N_28445,N_27651,N_27797);
or U28446 (N_28446,N_27420,N_27810);
and U28447 (N_28447,N_27275,N_27917);
nor U28448 (N_28448,N_27423,N_27723);
xnor U28449 (N_28449,N_27560,N_27457);
nand U28450 (N_28450,N_27116,N_27923);
nor U28451 (N_28451,N_27323,N_27653);
nor U28452 (N_28452,N_27791,N_27297);
and U28453 (N_28453,N_27474,N_27125);
nor U28454 (N_28454,N_27679,N_27164);
nand U28455 (N_28455,N_27310,N_27005);
or U28456 (N_28456,N_27273,N_27799);
nor U28457 (N_28457,N_27741,N_27123);
and U28458 (N_28458,N_27811,N_27088);
or U28459 (N_28459,N_27370,N_27190);
nor U28460 (N_28460,N_27708,N_27322);
nand U28461 (N_28461,N_27585,N_27814);
or U28462 (N_28462,N_27621,N_27974);
or U28463 (N_28463,N_27717,N_27724);
xnor U28464 (N_28464,N_27061,N_27431);
xnor U28465 (N_28465,N_27942,N_27439);
or U28466 (N_28466,N_27819,N_27524);
and U28467 (N_28467,N_27404,N_27877);
or U28468 (N_28468,N_27242,N_27696);
and U28469 (N_28469,N_27900,N_27316);
xor U28470 (N_28470,N_27031,N_27718);
xor U28471 (N_28471,N_27211,N_27215);
and U28472 (N_28472,N_27740,N_27574);
xnor U28473 (N_28473,N_27614,N_27515);
or U28474 (N_28474,N_27650,N_27027);
xnor U28475 (N_28475,N_27344,N_27613);
and U28476 (N_28476,N_27137,N_27886);
nand U28477 (N_28477,N_27916,N_27380);
or U28478 (N_28478,N_27644,N_27544);
nor U28479 (N_28479,N_27391,N_27863);
xor U28480 (N_28480,N_27225,N_27019);
nand U28481 (N_28481,N_27481,N_27065);
nand U28482 (N_28482,N_27259,N_27305);
nor U28483 (N_28483,N_27433,N_27266);
nor U28484 (N_28484,N_27023,N_27605);
nor U28485 (N_28485,N_27823,N_27412);
and U28486 (N_28486,N_27034,N_27828);
nor U28487 (N_28487,N_27979,N_27634);
nor U28488 (N_28488,N_27640,N_27007);
and U28489 (N_28489,N_27849,N_27361);
nor U28490 (N_28490,N_27295,N_27117);
xor U28491 (N_28491,N_27957,N_27292);
or U28492 (N_28492,N_27501,N_27838);
nand U28493 (N_28493,N_27981,N_27222);
nand U28494 (N_28494,N_27139,N_27600);
and U28495 (N_28495,N_27795,N_27936);
and U28496 (N_28496,N_27124,N_27213);
xnor U28497 (N_28497,N_27308,N_27680);
nand U28498 (N_28498,N_27855,N_27610);
xor U28499 (N_28499,N_27056,N_27449);
xnor U28500 (N_28500,N_27140,N_27783);
and U28501 (N_28501,N_27568,N_27021);
and U28502 (N_28502,N_27029,N_27384);
xor U28503 (N_28503,N_27519,N_27066);
and U28504 (N_28504,N_27305,N_27705);
and U28505 (N_28505,N_27854,N_27510);
nand U28506 (N_28506,N_27953,N_27732);
and U28507 (N_28507,N_27227,N_27216);
xnor U28508 (N_28508,N_27999,N_27563);
and U28509 (N_28509,N_27653,N_27031);
nand U28510 (N_28510,N_27602,N_27930);
xor U28511 (N_28511,N_27600,N_27882);
xnor U28512 (N_28512,N_27815,N_27701);
nand U28513 (N_28513,N_27539,N_27981);
or U28514 (N_28514,N_27835,N_27793);
or U28515 (N_28515,N_27439,N_27434);
nor U28516 (N_28516,N_27413,N_27086);
nand U28517 (N_28517,N_27864,N_27161);
nand U28518 (N_28518,N_27834,N_27725);
and U28519 (N_28519,N_27763,N_27757);
xnor U28520 (N_28520,N_27352,N_27700);
nor U28521 (N_28521,N_27829,N_27341);
or U28522 (N_28522,N_27768,N_27122);
nor U28523 (N_28523,N_27864,N_27599);
nand U28524 (N_28524,N_27587,N_27978);
or U28525 (N_28525,N_27839,N_27341);
or U28526 (N_28526,N_27593,N_27383);
nor U28527 (N_28527,N_27571,N_27922);
and U28528 (N_28528,N_27704,N_27463);
nand U28529 (N_28529,N_27067,N_27431);
nand U28530 (N_28530,N_27397,N_27013);
and U28531 (N_28531,N_27963,N_27719);
or U28532 (N_28532,N_27414,N_27320);
nor U28533 (N_28533,N_27888,N_27913);
xor U28534 (N_28534,N_27235,N_27611);
and U28535 (N_28535,N_27467,N_27196);
or U28536 (N_28536,N_27938,N_27296);
nand U28537 (N_28537,N_27001,N_27903);
nor U28538 (N_28538,N_27905,N_27295);
nand U28539 (N_28539,N_27211,N_27826);
nor U28540 (N_28540,N_27646,N_27194);
and U28541 (N_28541,N_27581,N_27778);
nand U28542 (N_28542,N_27773,N_27993);
xor U28543 (N_28543,N_27122,N_27480);
xnor U28544 (N_28544,N_27115,N_27735);
nand U28545 (N_28545,N_27813,N_27757);
nor U28546 (N_28546,N_27010,N_27419);
or U28547 (N_28547,N_27318,N_27363);
xnor U28548 (N_28548,N_27840,N_27974);
or U28549 (N_28549,N_27271,N_27037);
or U28550 (N_28550,N_27730,N_27128);
or U28551 (N_28551,N_27528,N_27018);
nand U28552 (N_28552,N_27979,N_27332);
nor U28553 (N_28553,N_27477,N_27258);
nand U28554 (N_28554,N_27932,N_27803);
xnor U28555 (N_28555,N_27014,N_27244);
nor U28556 (N_28556,N_27536,N_27220);
or U28557 (N_28557,N_27827,N_27921);
or U28558 (N_28558,N_27897,N_27467);
or U28559 (N_28559,N_27532,N_27134);
or U28560 (N_28560,N_27935,N_27670);
nand U28561 (N_28561,N_27652,N_27216);
nand U28562 (N_28562,N_27510,N_27903);
or U28563 (N_28563,N_27729,N_27144);
or U28564 (N_28564,N_27540,N_27840);
and U28565 (N_28565,N_27600,N_27288);
and U28566 (N_28566,N_27979,N_27964);
nor U28567 (N_28567,N_27768,N_27262);
nand U28568 (N_28568,N_27932,N_27786);
or U28569 (N_28569,N_27044,N_27642);
or U28570 (N_28570,N_27866,N_27254);
and U28571 (N_28571,N_27756,N_27882);
nand U28572 (N_28572,N_27767,N_27094);
xnor U28573 (N_28573,N_27073,N_27546);
or U28574 (N_28574,N_27065,N_27170);
or U28575 (N_28575,N_27806,N_27987);
xor U28576 (N_28576,N_27019,N_27129);
and U28577 (N_28577,N_27998,N_27130);
or U28578 (N_28578,N_27460,N_27974);
xor U28579 (N_28579,N_27183,N_27340);
or U28580 (N_28580,N_27062,N_27151);
nor U28581 (N_28581,N_27142,N_27368);
nor U28582 (N_28582,N_27738,N_27438);
and U28583 (N_28583,N_27579,N_27405);
and U28584 (N_28584,N_27268,N_27367);
xnor U28585 (N_28585,N_27950,N_27811);
nand U28586 (N_28586,N_27232,N_27773);
nand U28587 (N_28587,N_27422,N_27189);
nand U28588 (N_28588,N_27829,N_27234);
nand U28589 (N_28589,N_27171,N_27454);
or U28590 (N_28590,N_27874,N_27553);
nand U28591 (N_28591,N_27132,N_27760);
nand U28592 (N_28592,N_27569,N_27314);
and U28593 (N_28593,N_27549,N_27812);
and U28594 (N_28594,N_27585,N_27553);
or U28595 (N_28595,N_27306,N_27208);
and U28596 (N_28596,N_27510,N_27174);
nor U28597 (N_28597,N_27252,N_27059);
and U28598 (N_28598,N_27561,N_27745);
xor U28599 (N_28599,N_27697,N_27889);
and U28600 (N_28600,N_27426,N_27598);
and U28601 (N_28601,N_27085,N_27631);
nand U28602 (N_28602,N_27542,N_27650);
or U28603 (N_28603,N_27836,N_27192);
or U28604 (N_28604,N_27983,N_27820);
nor U28605 (N_28605,N_27709,N_27483);
or U28606 (N_28606,N_27911,N_27172);
nor U28607 (N_28607,N_27820,N_27675);
nand U28608 (N_28608,N_27257,N_27957);
nor U28609 (N_28609,N_27553,N_27987);
and U28610 (N_28610,N_27140,N_27185);
xor U28611 (N_28611,N_27048,N_27946);
and U28612 (N_28612,N_27908,N_27888);
and U28613 (N_28613,N_27247,N_27610);
and U28614 (N_28614,N_27812,N_27644);
xnor U28615 (N_28615,N_27939,N_27595);
nand U28616 (N_28616,N_27843,N_27018);
or U28617 (N_28617,N_27968,N_27600);
and U28618 (N_28618,N_27987,N_27959);
nor U28619 (N_28619,N_27799,N_27554);
nor U28620 (N_28620,N_27084,N_27097);
or U28621 (N_28621,N_27936,N_27943);
nor U28622 (N_28622,N_27564,N_27590);
nand U28623 (N_28623,N_27158,N_27513);
nor U28624 (N_28624,N_27391,N_27248);
or U28625 (N_28625,N_27343,N_27489);
nand U28626 (N_28626,N_27783,N_27596);
xnor U28627 (N_28627,N_27741,N_27795);
nand U28628 (N_28628,N_27392,N_27077);
nand U28629 (N_28629,N_27652,N_27362);
nor U28630 (N_28630,N_27655,N_27011);
nor U28631 (N_28631,N_27837,N_27537);
and U28632 (N_28632,N_27921,N_27297);
and U28633 (N_28633,N_27890,N_27952);
and U28634 (N_28634,N_27764,N_27118);
xor U28635 (N_28635,N_27722,N_27214);
nand U28636 (N_28636,N_27806,N_27173);
xor U28637 (N_28637,N_27323,N_27573);
nor U28638 (N_28638,N_27077,N_27127);
nor U28639 (N_28639,N_27902,N_27312);
and U28640 (N_28640,N_27146,N_27822);
xor U28641 (N_28641,N_27993,N_27283);
and U28642 (N_28642,N_27131,N_27087);
or U28643 (N_28643,N_27101,N_27363);
nand U28644 (N_28644,N_27013,N_27507);
nor U28645 (N_28645,N_27023,N_27409);
nand U28646 (N_28646,N_27410,N_27076);
nor U28647 (N_28647,N_27214,N_27716);
nor U28648 (N_28648,N_27535,N_27721);
and U28649 (N_28649,N_27589,N_27713);
nand U28650 (N_28650,N_27100,N_27831);
nand U28651 (N_28651,N_27103,N_27567);
nor U28652 (N_28652,N_27366,N_27148);
nor U28653 (N_28653,N_27597,N_27608);
nor U28654 (N_28654,N_27701,N_27547);
and U28655 (N_28655,N_27472,N_27787);
or U28656 (N_28656,N_27900,N_27647);
nor U28657 (N_28657,N_27415,N_27671);
and U28658 (N_28658,N_27579,N_27671);
nor U28659 (N_28659,N_27825,N_27730);
and U28660 (N_28660,N_27802,N_27218);
nor U28661 (N_28661,N_27080,N_27671);
xnor U28662 (N_28662,N_27678,N_27118);
nor U28663 (N_28663,N_27914,N_27308);
nand U28664 (N_28664,N_27762,N_27024);
nand U28665 (N_28665,N_27137,N_27891);
or U28666 (N_28666,N_27278,N_27132);
and U28667 (N_28667,N_27386,N_27118);
nand U28668 (N_28668,N_27375,N_27269);
or U28669 (N_28669,N_27168,N_27049);
nand U28670 (N_28670,N_27785,N_27173);
nor U28671 (N_28671,N_27755,N_27465);
or U28672 (N_28672,N_27072,N_27350);
nor U28673 (N_28673,N_27125,N_27257);
nor U28674 (N_28674,N_27147,N_27410);
nor U28675 (N_28675,N_27287,N_27171);
nor U28676 (N_28676,N_27007,N_27057);
nor U28677 (N_28677,N_27805,N_27217);
and U28678 (N_28678,N_27848,N_27333);
or U28679 (N_28679,N_27206,N_27093);
and U28680 (N_28680,N_27067,N_27267);
nor U28681 (N_28681,N_27037,N_27280);
xor U28682 (N_28682,N_27483,N_27119);
and U28683 (N_28683,N_27097,N_27728);
or U28684 (N_28684,N_27130,N_27630);
or U28685 (N_28685,N_27582,N_27520);
and U28686 (N_28686,N_27255,N_27775);
nor U28687 (N_28687,N_27039,N_27781);
nand U28688 (N_28688,N_27279,N_27035);
xor U28689 (N_28689,N_27703,N_27735);
nand U28690 (N_28690,N_27069,N_27284);
xor U28691 (N_28691,N_27446,N_27544);
and U28692 (N_28692,N_27198,N_27570);
and U28693 (N_28693,N_27283,N_27464);
and U28694 (N_28694,N_27254,N_27321);
xor U28695 (N_28695,N_27063,N_27852);
and U28696 (N_28696,N_27067,N_27403);
nor U28697 (N_28697,N_27812,N_27490);
or U28698 (N_28698,N_27986,N_27634);
and U28699 (N_28699,N_27188,N_27660);
or U28700 (N_28700,N_27835,N_27020);
nor U28701 (N_28701,N_27743,N_27093);
nand U28702 (N_28702,N_27783,N_27014);
xnor U28703 (N_28703,N_27841,N_27603);
nor U28704 (N_28704,N_27056,N_27311);
nor U28705 (N_28705,N_27846,N_27000);
or U28706 (N_28706,N_27687,N_27230);
xor U28707 (N_28707,N_27546,N_27451);
nand U28708 (N_28708,N_27381,N_27515);
and U28709 (N_28709,N_27714,N_27777);
or U28710 (N_28710,N_27040,N_27248);
or U28711 (N_28711,N_27182,N_27252);
and U28712 (N_28712,N_27512,N_27841);
nand U28713 (N_28713,N_27306,N_27582);
nor U28714 (N_28714,N_27598,N_27571);
or U28715 (N_28715,N_27415,N_27948);
xnor U28716 (N_28716,N_27093,N_27879);
xnor U28717 (N_28717,N_27928,N_27004);
xnor U28718 (N_28718,N_27957,N_27532);
or U28719 (N_28719,N_27976,N_27083);
nor U28720 (N_28720,N_27928,N_27862);
nor U28721 (N_28721,N_27924,N_27953);
nor U28722 (N_28722,N_27718,N_27496);
nand U28723 (N_28723,N_27848,N_27449);
xnor U28724 (N_28724,N_27648,N_27956);
xor U28725 (N_28725,N_27525,N_27151);
nand U28726 (N_28726,N_27437,N_27909);
nand U28727 (N_28727,N_27153,N_27203);
and U28728 (N_28728,N_27972,N_27278);
nor U28729 (N_28729,N_27369,N_27046);
nand U28730 (N_28730,N_27219,N_27878);
nand U28731 (N_28731,N_27345,N_27131);
xor U28732 (N_28732,N_27978,N_27700);
nor U28733 (N_28733,N_27672,N_27363);
nor U28734 (N_28734,N_27252,N_27219);
and U28735 (N_28735,N_27899,N_27377);
nand U28736 (N_28736,N_27542,N_27580);
nand U28737 (N_28737,N_27685,N_27817);
nor U28738 (N_28738,N_27022,N_27482);
or U28739 (N_28739,N_27743,N_27381);
or U28740 (N_28740,N_27742,N_27034);
nand U28741 (N_28741,N_27639,N_27099);
nand U28742 (N_28742,N_27440,N_27149);
and U28743 (N_28743,N_27712,N_27101);
nand U28744 (N_28744,N_27602,N_27323);
xnor U28745 (N_28745,N_27600,N_27479);
xnor U28746 (N_28746,N_27915,N_27903);
and U28747 (N_28747,N_27799,N_27108);
xor U28748 (N_28748,N_27323,N_27739);
nor U28749 (N_28749,N_27585,N_27971);
nor U28750 (N_28750,N_27383,N_27677);
and U28751 (N_28751,N_27435,N_27076);
nand U28752 (N_28752,N_27879,N_27943);
nand U28753 (N_28753,N_27086,N_27939);
nor U28754 (N_28754,N_27337,N_27257);
nand U28755 (N_28755,N_27602,N_27190);
and U28756 (N_28756,N_27277,N_27053);
nor U28757 (N_28757,N_27761,N_27544);
nor U28758 (N_28758,N_27693,N_27138);
or U28759 (N_28759,N_27727,N_27845);
xor U28760 (N_28760,N_27229,N_27257);
xnor U28761 (N_28761,N_27214,N_27104);
or U28762 (N_28762,N_27367,N_27502);
nand U28763 (N_28763,N_27375,N_27807);
and U28764 (N_28764,N_27784,N_27727);
nor U28765 (N_28765,N_27559,N_27145);
nor U28766 (N_28766,N_27296,N_27447);
and U28767 (N_28767,N_27218,N_27082);
nor U28768 (N_28768,N_27450,N_27407);
or U28769 (N_28769,N_27779,N_27902);
or U28770 (N_28770,N_27059,N_27689);
or U28771 (N_28771,N_27705,N_27331);
nand U28772 (N_28772,N_27747,N_27875);
or U28773 (N_28773,N_27966,N_27310);
xnor U28774 (N_28774,N_27375,N_27463);
nor U28775 (N_28775,N_27821,N_27199);
nor U28776 (N_28776,N_27000,N_27943);
or U28777 (N_28777,N_27249,N_27728);
nor U28778 (N_28778,N_27062,N_27751);
nand U28779 (N_28779,N_27267,N_27883);
or U28780 (N_28780,N_27835,N_27616);
or U28781 (N_28781,N_27579,N_27580);
and U28782 (N_28782,N_27485,N_27637);
nand U28783 (N_28783,N_27255,N_27039);
or U28784 (N_28784,N_27322,N_27249);
or U28785 (N_28785,N_27455,N_27177);
nand U28786 (N_28786,N_27264,N_27599);
nor U28787 (N_28787,N_27526,N_27263);
xnor U28788 (N_28788,N_27516,N_27691);
nor U28789 (N_28789,N_27209,N_27192);
xor U28790 (N_28790,N_27565,N_27469);
or U28791 (N_28791,N_27508,N_27289);
xor U28792 (N_28792,N_27244,N_27046);
or U28793 (N_28793,N_27563,N_27897);
and U28794 (N_28794,N_27567,N_27922);
and U28795 (N_28795,N_27268,N_27623);
and U28796 (N_28796,N_27073,N_27282);
or U28797 (N_28797,N_27105,N_27163);
nor U28798 (N_28798,N_27182,N_27127);
and U28799 (N_28799,N_27142,N_27839);
and U28800 (N_28800,N_27579,N_27121);
xnor U28801 (N_28801,N_27633,N_27762);
xnor U28802 (N_28802,N_27315,N_27930);
nor U28803 (N_28803,N_27932,N_27453);
and U28804 (N_28804,N_27750,N_27051);
nand U28805 (N_28805,N_27094,N_27737);
or U28806 (N_28806,N_27054,N_27693);
and U28807 (N_28807,N_27112,N_27385);
and U28808 (N_28808,N_27223,N_27347);
nor U28809 (N_28809,N_27631,N_27279);
xor U28810 (N_28810,N_27850,N_27232);
and U28811 (N_28811,N_27806,N_27495);
xor U28812 (N_28812,N_27084,N_27631);
nor U28813 (N_28813,N_27371,N_27803);
or U28814 (N_28814,N_27293,N_27835);
nand U28815 (N_28815,N_27727,N_27717);
and U28816 (N_28816,N_27400,N_27791);
xor U28817 (N_28817,N_27579,N_27807);
nand U28818 (N_28818,N_27860,N_27605);
xnor U28819 (N_28819,N_27768,N_27828);
nor U28820 (N_28820,N_27284,N_27720);
nor U28821 (N_28821,N_27823,N_27249);
or U28822 (N_28822,N_27427,N_27435);
or U28823 (N_28823,N_27199,N_27163);
nand U28824 (N_28824,N_27988,N_27030);
nand U28825 (N_28825,N_27976,N_27091);
or U28826 (N_28826,N_27833,N_27856);
xnor U28827 (N_28827,N_27827,N_27775);
nand U28828 (N_28828,N_27700,N_27254);
or U28829 (N_28829,N_27550,N_27175);
xnor U28830 (N_28830,N_27429,N_27000);
xnor U28831 (N_28831,N_27073,N_27300);
nand U28832 (N_28832,N_27935,N_27139);
xnor U28833 (N_28833,N_27565,N_27724);
or U28834 (N_28834,N_27354,N_27781);
nor U28835 (N_28835,N_27374,N_27867);
or U28836 (N_28836,N_27009,N_27388);
nand U28837 (N_28837,N_27304,N_27539);
nor U28838 (N_28838,N_27760,N_27992);
xnor U28839 (N_28839,N_27327,N_27407);
xor U28840 (N_28840,N_27072,N_27238);
nor U28841 (N_28841,N_27818,N_27183);
and U28842 (N_28842,N_27386,N_27609);
nor U28843 (N_28843,N_27233,N_27076);
and U28844 (N_28844,N_27109,N_27497);
nor U28845 (N_28845,N_27229,N_27705);
xnor U28846 (N_28846,N_27016,N_27289);
nor U28847 (N_28847,N_27097,N_27887);
nand U28848 (N_28848,N_27966,N_27587);
xor U28849 (N_28849,N_27516,N_27803);
nand U28850 (N_28850,N_27615,N_27741);
nand U28851 (N_28851,N_27738,N_27384);
nor U28852 (N_28852,N_27645,N_27557);
nor U28853 (N_28853,N_27950,N_27464);
nor U28854 (N_28854,N_27366,N_27512);
nor U28855 (N_28855,N_27647,N_27638);
and U28856 (N_28856,N_27163,N_27032);
nand U28857 (N_28857,N_27215,N_27440);
or U28858 (N_28858,N_27978,N_27188);
xor U28859 (N_28859,N_27719,N_27181);
xnor U28860 (N_28860,N_27738,N_27895);
nor U28861 (N_28861,N_27851,N_27499);
nand U28862 (N_28862,N_27551,N_27603);
and U28863 (N_28863,N_27847,N_27438);
xor U28864 (N_28864,N_27732,N_27896);
nor U28865 (N_28865,N_27541,N_27713);
or U28866 (N_28866,N_27992,N_27495);
and U28867 (N_28867,N_27007,N_27741);
or U28868 (N_28868,N_27264,N_27552);
or U28869 (N_28869,N_27042,N_27787);
nand U28870 (N_28870,N_27667,N_27920);
or U28871 (N_28871,N_27740,N_27590);
nand U28872 (N_28872,N_27499,N_27317);
nand U28873 (N_28873,N_27929,N_27223);
nor U28874 (N_28874,N_27604,N_27317);
xor U28875 (N_28875,N_27363,N_27447);
and U28876 (N_28876,N_27851,N_27505);
nor U28877 (N_28877,N_27913,N_27938);
xor U28878 (N_28878,N_27046,N_27239);
or U28879 (N_28879,N_27065,N_27508);
or U28880 (N_28880,N_27765,N_27367);
and U28881 (N_28881,N_27048,N_27021);
or U28882 (N_28882,N_27221,N_27132);
or U28883 (N_28883,N_27685,N_27076);
xor U28884 (N_28884,N_27891,N_27701);
or U28885 (N_28885,N_27961,N_27628);
nand U28886 (N_28886,N_27349,N_27106);
or U28887 (N_28887,N_27126,N_27936);
or U28888 (N_28888,N_27073,N_27516);
or U28889 (N_28889,N_27316,N_27517);
or U28890 (N_28890,N_27992,N_27502);
or U28891 (N_28891,N_27602,N_27774);
or U28892 (N_28892,N_27427,N_27507);
nand U28893 (N_28893,N_27535,N_27851);
or U28894 (N_28894,N_27235,N_27362);
xor U28895 (N_28895,N_27933,N_27868);
or U28896 (N_28896,N_27040,N_27709);
or U28897 (N_28897,N_27857,N_27811);
nand U28898 (N_28898,N_27447,N_27710);
or U28899 (N_28899,N_27889,N_27758);
xor U28900 (N_28900,N_27570,N_27132);
nor U28901 (N_28901,N_27194,N_27011);
and U28902 (N_28902,N_27137,N_27469);
nor U28903 (N_28903,N_27828,N_27733);
or U28904 (N_28904,N_27018,N_27504);
and U28905 (N_28905,N_27781,N_27347);
nand U28906 (N_28906,N_27423,N_27017);
and U28907 (N_28907,N_27125,N_27558);
nor U28908 (N_28908,N_27279,N_27370);
or U28909 (N_28909,N_27267,N_27260);
nand U28910 (N_28910,N_27708,N_27914);
nand U28911 (N_28911,N_27014,N_27390);
nand U28912 (N_28912,N_27616,N_27679);
nand U28913 (N_28913,N_27291,N_27798);
xnor U28914 (N_28914,N_27922,N_27470);
and U28915 (N_28915,N_27238,N_27058);
or U28916 (N_28916,N_27710,N_27994);
and U28917 (N_28917,N_27736,N_27789);
or U28918 (N_28918,N_27479,N_27865);
and U28919 (N_28919,N_27277,N_27076);
or U28920 (N_28920,N_27540,N_27307);
xnor U28921 (N_28921,N_27910,N_27875);
nor U28922 (N_28922,N_27701,N_27581);
nor U28923 (N_28923,N_27292,N_27296);
or U28924 (N_28924,N_27999,N_27530);
or U28925 (N_28925,N_27649,N_27628);
xor U28926 (N_28926,N_27062,N_27221);
nand U28927 (N_28927,N_27116,N_27859);
xor U28928 (N_28928,N_27129,N_27672);
and U28929 (N_28929,N_27466,N_27420);
or U28930 (N_28930,N_27586,N_27408);
nand U28931 (N_28931,N_27142,N_27814);
nor U28932 (N_28932,N_27098,N_27033);
nand U28933 (N_28933,N_27535,N_27445);
or U28934 (N_28934,N_27216,N_27837);
or U28935 (N_28935,N_27703,N_27011);
or U28936 (N_28936,N_27024,N_27455);
or U28937 (N_28937,N_27178,N_27916);
and U28938 (N_28938,N_27487,N_27443);
and U28939 (N_28939,N_27344,N_27213);
nand U28940 (N_28940,N_27733,N_27647);
or U28941 (N_28941,N_27289,N_27286);
or U28942 (N_28942,N_27600,N_27910);
xnor U28943 (N_28943,N_27663,N_27789);
nor U28944 (N_28944,N_27514,N_27355);
or U28945 (N_28945,N_27351,N_27299);
xor U28946 (N_28946,N_27675,N_27411);
nand U28947 (N_28947,N_27724,N_27242);
nor U28948 (N_28948,N_27227,N_27237);
nand U28949 (N_28949,N_27304,N_27289);
and U28950 (N_28950,N_27224,N_27903);
nand U28951 (N_28951,N_27677,N_27150);
nand U28952 (N_28952,N_27237,N_27062);
and U28953 (N_28953,N_27118,N_27339);
nand U28954 (N_28954,N_27152,N_27338);
or U28955 (N_28955,N_27212,N_27211);
xnor U28956 (N_28956,N_27016,N_27732);
nor U28957 (N_28957,N_27439,N_27315);
or U28958 (N_28958,N_27697,N_27151);
and U28959 (N_28959,N_27281,N_27336);
nand U28960 (N_28960,N_27395,N_27505);
and U28961 (N_28961,N_27959,N_27301);
nor U28962 (N_28962,N_27775,N_27008);
or U28963 (N_28963,N_27723,N_27247);
xnor U28964 (N_28964,N_27077,N_27388);
xor U28965 (N_28965,N_27125,N_27630);
and U28966 (N_28966,N_27562,N_27112);
nor U28967 (N_28967,N_27527,N_27844);
xnor U28968 (N_28968,N_27996,N_27863);
xor U28969 (N_28969,N_27686,N_27677);
nand U28970 (N_28970,N_27063,N_27363);
nor U28971 (N_28971,N_27289,N_27015);
xnor U28972 (N_28972,N_27987,N_27971);
or U28973 (N_28973,N_27924,N_27872);
and U28974 (N_28974,N_27702,N_27272);
nor U28975 (N_28975,N_27495,N_27279);
xor U28976 (N_28976,N_27624,N_27405);
xnor U28977 (N_28977,N_27342,N_27950);
nand U28978 (N_28978,N_27348,N_27922);
xor U28979 (N_28979,N_27870,N_27894);
nand U28980 (N_28980,N_27382,N_27791);
and U28981 (N_28981,N_27945,N_27144);
or U28982 (N_28982,N_27391,N_27616);
and U28983 (N_28983,N_27489,N_27306);
or U28984 (N_28984,N_27655,N_27029);
xnor U28985 (N_28985,N_27988,N_27786);
or U28986 (N_28986,N_27811,N_27987);
nor U28987 (N_28987,N_27515,N_27326);
or U28988 (N_28988,N_27650,N_27435);
nor U28989 (N_28989,N_27846,N_27965);
and U28990 (N_28990,N_27876,N_27452);
or U28991 (N_28991,N_27519,N_27137);
nor U28992 (N_28992,N_27351,N_27862);
and U28993 (N_28993,N_27509,N_27081);
nor U28994 (N_28994,N_27913,N_27330);
nor U28995 (N_28995,N_27504,N_27979);
nor U28996 (N_28996,N_27867,N_27024);
or U28997 (N_28997,N_27683,N_27868);
nor U28998 (N_28998,N_27882,N_27648);
xnor U28999 (N_28999,N_27867,N_27594);
nor U29000 (N_29000,N_28235,N_28760);
nor U29001 (N_29001,N_28511,N_28953);
xor U29002 (N_29002,N_28335,N_28477);
nor U29003 (N_29003,N_28952,N_28815);
nor U29004 (N_29004,N_28308,N_28174);
xor U29005 (N_29005,N_28980,N_28240);
xnor U29006 (N_29006,N_28364,N_28618);
xnor U29007 (N_29007,N_28877,N_28951);
nand U29008 (N_29008,N_28646,N_28049);
and U29009 (N_29009,N_28725,N_28449);
and U29010 (N_29010,N_28098,N_28237);
and U29011 (N_29011,N_28921,N_28890);
and U29012 (N_29012,N_28816,N_28376);
and U29013 (N_29013,N_28405,N_28132);
and U29014 (N_29014,N_28165,N_28860);
and U29015 (N_29015,N_28221,N_28252);
xor U29016 (N_29016,N_28773,N_28895);
xor U29017 (N_29017,N_28341,N_28406);
xor U29018 (N_29018,N_28798,N_28626);
nor U29019 (N_29019,N_28631,N_28894);
or U29020 (N_29020,N_28995,N_28526);
or U29021 (N_29021,N_28030,N_28923);
xor U29022 (N_29022,N_28647,N_28957);
or U29023 (N_29023,N_28580,N_28474);
nand U29024 (N_29024,N_28400,N_28264);
xnor U29025 (N_29025,N_28115,N_28217);
nand U29026 (N_29026,N_28508,N_28286);
nor U29027 (N_29027,N_28467,N_28485);
and U29028 (N_29028,N_28986,N_28581);
nand U29029 (N_29029,N_28911,N_28463);
and U29030 (N_29030,N_28338,N_28226);
and U29031 (N_29031,N_28686,N_28480);
nor U29032 (N_29032,N_28433,N_28045);
and U29033 (N_29033,N_28799,N_28837);
or U29034 (N_29034,N_28883,N_28590);
or U29035 (N_29035,N_28154,N_28684);
nor U29036 (N_29036,N_28990,N_28993);
and U29037 (N_29037,N_28055,N_28362);
nor U29038 (N_29038,N_28196,N_28231);
xnor U29039 (N_29039,N_28109,N_28788);
nor U29040 (N_29040,N_28705,N_28676);
xnor U29041 (N_29041,N_28718,N_28133);
xor U29042 (N_29042,N_28016,N_28922);
nor U29043 (N_29043,N_28628,N_28600);
nand U29044 (N_29044,N_28092,N_28037);
nor U29045 (N_29045,N_28988,N_28775);
xor U29046 (N_29046,N_28146,N_28163);
or U29047 (N_29047,N_28366,N_28567);
nand U29048 (N_29048,N_28868,N_28932);
or U29049 (N_29049,N_28211,N_28666);
nor U29050 (N_29050,N_28492,N_28562);
nand U29051 (N_29051,N_28658,N_28110);
and U29052 (N_29052,N_28036,N_28248);
nand U29053 (N_29053,N_28404,N_28328);
and U29054 (N_29054,N_28242,N_28206);
and U29055 (N_29055,N_28949,N_28535);
nand U29056 (N_29056,N_28886,N_28593);
and U29057 (N_29057,N_28246,N_28490);
xnor U29058 (N_29058,N_28582,N_28459);
nor U29059 (N_29059,N_28564,N_28357);
and U29060 (N_29060,N_28840,N_28738);
or U29061 (N_29061,N_28101,N_28529);
nand U29062 (N_29062,N_28550,N_28530);
nand U29063 (N_29063,N_28282,N_28822);
nor U29064 (N_29064,N_28586,N_28220);
or U29065 (N_29065,N_28609,N_28315);
nand U29066 (N_29066,N_28538,N_28208);
nand U29067 (N_29067,N_28834,N_28363);
and U29068 (N_29068,N_28108,N_28809);
nor U29069 (N_29069,N_28566,N_28399);
and U29070 (N_29070,N_28097,N_28591);
xor U29071 (N_29071,N_28804,N_28881);
nand U29072 (N_29072,N_28369,N_28352);
and U29073 (N_29073,N_28739,N_28959);
or U29074 (N_29074,N_28380,N_28943);
and U29075 (N_29075,N_28940,N_28519);
nor U29076 (N_29076,N_28428,N_28033);
xnor U29077 (N_29077,N_28408,N_28313);
or U29078 (N_29078,N_28180,N_28325);
nor U29079 (N_29079,N_28546,N_28349);
nor U29080 (N_29080,N_28744,N_28393);
nand U29081 (N_29081,N_28768,N_28861);
nand U29082 (N_29082,N_28501,N_28189);
nor U29083 (N_29083,N_28670,N_28532);
or U29084 (N_29084,N_28625,N_28219);
and U29085 (N_29085,N_28700,N_28446);
or U29086 (N_29086,N_28041,N_28948);
xor U29087 (N_29087,N_28624,N_28149);
xor U29088 (N_29088,N_28355,N_28409);
or U29089 (N_29089,N_28298,N_28391);
and U29090 (N_29090,N_28786,N_28599);
and U29091 (N_29091,N_28426,N_28571);
nand U29092 (N_29092,N_28503,N_28774);
and U29093 (N_29093,N_28724,N_28852);
xnor U29094 (N_29094,N_28120,N_28276);
or U29095 (N_29095,N_28425,N_28152);
and U29096 (N_29096,N_28847,N_28023);
nand U29097 (N_29097,N_28669,N_28392);
nand U29098 (N_29098,N_28175,N_28878);
or U29099 (N_29099,N_28505,N_28401);
nand U29100 (N_29100,N_28765,N_28982);
nor U29101 (N_29101,N_28306,N_28507);
nor U29102 (N_29102,N_28020,N_28899);
or U29103 (N_29103,N_28367,N_28976);
xnor U29104 (N_29104,N_28169,N_28342);
nand U29105 (N_29105,N_28130,N_28227);
or U29106 (N_29106,N_28035,N_28554);
nand U29107 (N_29107,N_28472,N_28632);
nor U29108 (N_29108,N_28673,N_28173);
nand U29109 (N_29109,N_28950,N_28142);
or U29110 (N_29110,N_28360,N_28012);
xor U29111 (N_29111,N_28927,N_28195);
nand U29112 (N_29112,N_28121,N_28859);
and U29113 (N_29113,N_28117,N_28164);
nor U29114 (N_29114,N_28687,N_28509);
or U29115 (N_29115,N_28374,N_28487);
nor U29116 (N_29116,N_28610,N_28300);
and U29117 (N_29117,N_28884,N_28451);
xor U29118 (N_29118,N_28712,N_28692);
and U29119 (N_29119,N_28430,N_28915);
or U29120 (N_29120,N_28569,N_28780);
and U29121 (N_29121,N_28607,N_28332);
or U29122 (N_29122,N_28579,N_28637);
and U29123 (N_29123,N_28821,N_28874);
xor U29124 (N_29124,N_28797,N_28733);
or U29125 (N_29125,N_28551,N_28213);
nor U29126 (N_29126,N_28134,N_28194);
nor U29127 (N_29127,N_28281,N_28722);
or U29128 (N_29128,N_28981,N_28389);
nor U29129 (N_29129,N_28787,N_28057);
nand U29130 (N_29130,N_28261,N_28256);
and U29131 (N_29131,N_28159,N_28061);
xor U29132 (N_29132,N_28064,N_28523);
nand U29133 (N_29133,N_28954,N_28204);
xor U29134 (N_29134,N_28278,N_28207);
or U29135 (N_29135,N_28423,N_28254);
and U29136 (N_29136,N_28751,N_28888);
and U29137 (N_29137,N_28141,N_28065);
or U29138 (N_29138,N_28015,N_28572);
or U29139 (N_29139,N_28277,N_28537);
nand U29140 (N_29140,N_28873,N_28814);
and U29141 (N_29141,N_28462,N_28145);
nor U29142 (N_29142,N_28067,N_28693);
or U29143 (N_29143,N_28148,N_28122);
and U29144 (N_29144,N_28892,N_28914);
or U29145 (N_29145,N_28627,N_28613);
or U29146 (N_29146,N_28489,N_28439);
or U29147 (N_29147,N_28008,N_28191);
and U29148 (N_29148,N_28677,N_28641);
and U29149 (N_29149,N_28728,N_28629);
xor U29150 (N_29150,N_28026,N_28387);
xnor U29151 (N_29151,N_28161,N_28772);
or U29152 (N_29152,N_28536,N_28044);
nor U29153 (N_29153,N_28769,N_28737);
and U29154 (N_29154,N_28573,N_28155);
or U29155 (N_29155,N_28443,N_28214);
or U29156 (N_29156,N_28450,N_28085);
nor U29157 (N_29157,N_28513,N_28455);
nand U29158 (N_29158,N_28650,N_28790);
or U29159 (N_29159,N_28690,N_28688);
nand U29160 (N_29160,N_28001,N_28937);
xnor U29161 (N_29161,N_28568,N_28322);
nor U29162 (N_29162,N_28601,N_28229);
or U29163 (N_29163,N_28233,N_28018);
and U29164 (N_29164,N_28754,N_28828);
nor U29165 (N_29165,N_28386,N_28113);
nor U29166 (N_29166,N_28069,N_28926);
nor U29167 (N_29167,N_28283,N_28448);
nor U29168 (N_29168,N_28946,N_28707);
or U29169 (N_29169,N_28025,N_28654);
nand U29170 (N_29170,N_28063,N_28114);
xor U29171 (N_29171,N_28620,N_28010);
xor U29172 (N_29172,N_28241,N_28694);
xor U29173 (N_29173,N_28397,N_28517);
xor U29174 (N_29174,N_28849,N_28402);
or U29175 (N_29175,N_28305,N_28077);
nor U29176 (N_29176,N_28547,N_28727);
or U29177 (N_29177,N_28955,N_28597);
nor U29178 (N_29178,N_28638,N_28312);
or U29179 (N_29179,N_28831,N_28703);
xor U29180 (N_29180,N_28311,N_28193);
nor U29181 (N_29181,N_28592,N_28603);
xnor U29182 (N_29182,N_28778,N_28333);
nor U29183 (N_29183,N_28717,N_28259);
xor U29184 (N_29184,N_28541,N_28465);
nand U29185 (N_29185,N_28854,N_28350);
nor U29186 (N_29186,N_28839,N_28475);
and U29187 (N_29187,N_28726,N_28781);
nand U29188 (N_29188,N_28906,N_28762);
or U29189 (N_29189,N_28356,N_28617);
nand U29190 (N_29190,N_28909,N_28052);
nor U29191 (N_29191,N_28301,N_28558);
or U29192 (N_29192,N_28583,N_28969);
xnor U29193 (N_29193,N_28095,N_28518);
nor U29194 (N_29194,N_28589,N_28939);
xor U29195 (N_29195,N_28723,N_28904);
or U29196 (N_29196,N_28038,N_28396);
xnor U29197 (N_29197,N_28924,N_28970);
nand U29198 (N_29198,N_28398,N_28087);
nor U29199 (N_29199,N_28758,N_28060);
xor U29200 (N_29200,N_28232,N_28978);
and U29201 (N_29201,N_28343,N_28496);
nand U29202 (N_29202,N_28999,N_28071);
nand U29203 (N_29203,N_28785,N_28295);
or U29204 (N_29204,N_28075,N_28678);
and U29205 (N_29205,N_28263,N_28812);
and U29206 (N_29206,N_28942,N_28099);
nand U29207 (N_29207,N_28292,N_28059);
xor U29208 (N_29208,N_28963,N_28156);
or U29209 (N_29209,N_28671,N_28323);
nor U29210 (N_29210,N_28190,N_28732);
nand U29211 (N_29211,N_28017,N_28789);
or U29212 (N_29212,N_28740,N_28317);
and U29213 (N_29213,N_28046,N_28655);
or U29214 (N_29214,N_28556,N_28716);
nor U29215 (N_29215,N_28351,N_28228);
xor U29216 (N_29216,N_28850,N_28424);
nand U29217 (N_29217,N_28370,N_28106);
nand U29218 (N_29218,N_28466,N_28047);
nor U29219 (N_29219,N_28479,N_28710);
xor U29220 (N_29220,N_28500,N_28050);
xnor U29221 (N_29221,N_28135,N_28808);
or U29222 (N_29222,N_28897,N_28685);
nor U29223 (N_29223,N_28365,N_28652);
and U29224 (N_29224,N_28078,N_28326);
nand U29225 (N_29225,N_28702,N_28329);
xnor U29226 (N_29226,N_28086,N_28889);
xor U29227 (N_29227,N_28810,N_28290);
and U29228 (N_29228,N_28559,N_28137);
nand U29229 (N_29229,N_28731,N_28482);
or U29230 (N_29230,N_28051,N_28497);
nor U29231 (N_29231,N_28696,N_28096);
xnor U29232 (N_29232,N_28805,N_28080);
xor U29233 (N_29233,N_28905,N_28979);
and U29234 (N_29234,N_28486,N_28176);
nand U29235 (N_29235,N_28561,N_28054);
xnor U29236 (N_29236,N_28570,N_28512);
xor U29237 (N_29237,N_28091,N_28994);
or U29238 (N_29238,N_28838,N_28372);
xor U29239 (N_29239,N_28525,N_28975);
and U29240 (N_29240,N_28930,N_28665);
nand U29241 (N_29241,N_28584,N_28014);
and U29242 (N_29242,N_28515,N_28265);
nor U29243 (N_29243,N_28407,N_28913);
xnor U29244 (N_29244,N_28766,N_28210);
nor U29245 (N_29245,N_28960,N_28084);
or U29246 (N_29246,N_28438,N_28461);
and U29247 (N_29247,N_28160,N_28249);
nor U29248 (N_29248,N_28514,N_28378);
nor U29249 (N_29249,N_28247,N_28166);
or U29250 (N_29250,N_28266,N_28179);
and U29251 (N_29251,N_28947,N_28171);
nor U29252 (N_29252,N_28250,N_28623);
nor U29253 (N_29253,N_28985,N_28445);
nand U29254 (N_29254,N_28936,N_28118);
or U29255 (N_29255,N_28661,N_28825);
or U29256 (N_29256,N_28473,N_28288);
xnor U29257 (N_29257,N_28689,N_28403);
xor U29258 (N_29258,N_28876,N_28680);
xnor U29259 (N_29259,N_28845,N_28285);
or U29260 (N_29260,N_28243,N_28000);
nor U29261 (N_29261,N_28444,N_28381);
and U29262 (N_29262,N_28144,N_28644);
xnor U29263 (N_29263,N_28271,N_28698);
and U29264 (N_29264,N_28304,N_28079);
xnor U29265 (N_29265,N_28039,N_28977);
or U29266 (N_29266,N_28792,N_28820);
xnor U29267 (N_29267,N_28824,N_28855);
and U29268 (N_29268,N_28094,N_28262);
nand U29269 (N_29269,N_28280,N_28898);
xor U29270 (N_29270,N_28273,N_28321);
nand U29271 (N_29271,N_28414,N_28663);
and U29272 (N_29272,N_28478,N_28359);
nand U29273 (N_29273,N_28441,N_28076);
xor U29274 (N_29274,N_28901,N_28269);
or U29275 (N_29275,N_28636,N_28320);
and U29276 (N_29276,N_28763,N_28752);
nor U29277 (N_29277,N_28823,N_28245);
and U29278 (N_29278,N_28974,N_28131);
and U29279 (N_29279,N_28761,N_28029);
or U29280 (N_29280,N_28082,N_28973);
nand U29281 (N_29281,N_28183,N_28498);
or U29282 (N_29282,N_28205,N_28056);
nor U29283 (N_29283,N_28848,N_28499);
and U29284 (N_29284,N_28964,N_28314);
nor U29285 (N_29285,N_28345,N_28494);
xnor U29286 (N_29286,N_28434,N_28418);
and U29287 (N_29287,N_28721,N_28996);
nand U29288 (N_29288,N_28293,N_28007);
or U29289 (N_29289,N_28138,N_28100);
nor U29290 (N_29290,N_28560,N_28481);
xor U29291 (N_29291,N_28844,N_28186);
and U29292 (N_29292,N_28125,N_28203);
nand U29293 (N_29293,N_28919,N_28297);
nor U29294 (N_29294,N_28239,N_28882);
nand U29295 (N_29295,N_28234,N_28634);
nand U29296 (N_29296,N_28832,N_28361);
nand U29297 (N_29297,N_28309,N_28531);
xnor U29298 (N_29298,N_28875,N_28377);
nand U29299 (N_29299,N_28124,N_28777);
nor U29300 (N_29300,N_28662,N_28630);
xor U29301 (N_29301,N_28502,N_28136);
xor U29302 (N_29302,N_28967,N_28604);
xor U29303 (N_29303,N_28594,N_28287);
nor U29304 (N_29304,N_28575,N_28188);
nand U29305 (N_29305,N_28682,N_28708);
xor U29306 (N_29306,N_28643,N_28983);
or U29307 (N_29307,N_28826,N_28743);
or U29308 (N_29308,N_28715,N_28436);
nor U29309 (N_29309,N_28938,N_28483);
and U29310 (N_29310,N_28770,N_28817);
nand U29311 (N_29311,N_28388,N_28251);
nand U29312 (N_29312,N_28608,N_28830);
nor U29313 (N_29313,N_28956,N_28918);
nand U29314 (N_29314,N_28656,N_28083);
xor U29315 (N_29315,N_28024,N_28683);
nor U29316 (N_29316,N_28865,N_28453);
xor U29317 (N_29317,N_28544,N_28432);
nand U29318 (N_29318,N_28104,N_28742);
xnor U29319 (N_29319,N_28827,N_28704);
and U29320 (N_29320,N_28435,N_28253);
nand U29321 (N_29321,N_28123,N_28756);
nand U29322 (N_29322,N_28224,N_28454);
nor U29323 (N_29323,N_28074,N_28794);
or U29324 (N_29324,N_28992,N_28371);
xnor U29325 (N_29325,N_28706,N_28040);
and U29326 (N_29326,N_28013,N_28611);
xnor U29327 (N_29327,N_28697,N_28533);
and U29328 (N_29328,N_28294,N_28642);
nand U29329 (N_29329,N_28495,N_28578);
and U29330 (N_29330,N_28931,N_28548);
or U29331 (N_29331,N_28182,N_28750);
or U29332 (N_29332,N_28070,N_28019);
nor U29333 (N_29333,N_28925,N_28150);
or U29334 (N_29334,N_28339,N_28928);
nand U29335 (N_29335,N_28653,N_28504);
xor U29336 (N_29336,N_28555,N_28218);
or U29337 (N_29337,N_28011,N_28172);
nand U29338 (N_29338,N_28659,N_28354);
and U29339 (N_29339,N_28310,N_28934);
nor U29340 (N_29340,N_28319,N_28456);
xnor U29341 (N_29341,N_28192,N_28119);
xnor U29342 (N_29342,N_28028,N_28212);
or U29343 (N_29343,N_28900,N_28053);
nand U29344 (N_29344,N_28128,N_28917);
nor U29345 (N_29345,N_28991,N_28962);
nor U29346 (N_29346,N_28307,N_28185);
or U29347 (N_29347,N_28574,N_28540);
or U29348 (N_29348,N_28089,N_28651);
and U29349 (N_29349,N_28720,N_28471);
nor U29350 (N_29350,N_28958,N_28419);
or U29351 (N_29351,N_28896,N_28639);
nand U29352 (N_29352,N_28116,N_28622);
and U29353 (N_29353,N_28764,N_28880);
xor U29354 (N_29354,N_28800,N_28126);
nand U29355 (N_29355,N_28714,N_28961);
xnor U29356 (N_29356,N_28545,N_28421);
nor U29357 (N_29357,N_28891,N_28072);
or U29358 (N_29358,N_28158,N_28612);
xor U29359 (N_29359,N_28379,N_28524);
nor U29360 (N_29360,N_28563,N_28199);
nor U29361 (N_29361,N_28616,N_28806);
and U29362 (N_29362,N_28635,N_28516);
or U29363 (N_29363,N_28695,N_28713);
nand U29364 (N_29364,N_28843,N_28468);
or U29365 (N_29365,N_28476,N_28565);
nand U29366 (N_29366,N_28989,N_28268);
xnor U29367 (N_29367,N_28879,N_28457);
nand U29368 (N_29368,N_28157,N_28729);
xor U29369 (N_29369,N_28440,N_28140);
xor U29370 (N_29370,N_28929,N_28701);
xnor U29371 (N_29371,N_28216,N_28331);
and U29372 (N_29372,N_28767,N_28527);
nand U29373 (N_29373,N_28674,N_28225);
and U29374 (N_29374,N_28577,N_28759);
and U29375 (N_29375,N_28184,N_28933);
nand U29376 (N_29376,N_28867,N_28022);
nand U29377 (N_29377,N_28941,N_28337);
or U29378 (N_29378,N_28452,N_28006);
or U29379 (N_29379,N_28803,N_28284);
nand U29380 (N_29380,N_28887,N_28966);
and U29381 (N_29381,N_28042,N_28347);
and U29382 (N_29382,N_28836,N_28147);
nor U29383 (N_29383,N_28021,N_28935);
xnor U29384 (N_29384,N_28416,N_28302);
xnor U29385 (N_29385,N_28330,N_28987);
nand U29386 (N_29386,N_28944,N_28353);
nand U29387 (N_29387,N_28068,N_28749);
nor U29388 (N_29388,N_28143,N_28753);
and U29389 (N_29389,N_28711,N_28105);
nand U29390 (N_29390,N_28139,N_28862);
nand U29391 (N_29391,N_28422,N_28869);
nor U29392 (N_29392,N_28296,N_28699);
xor U29393 (N_29393,N_28383,N_28410);
and U29394 (N_29394,N_28543,N_28818);
and U29395 (N_29395,N_28734,N_28346);
or U29396 (N_29396,N_28833,N_28829);
nor U29397 (N_29397,N_28649,N_28793);
and U29398 (N_29398,N_28972,N_28534);
and U29399 (N_29399,N_28334,N_28093);
or U29400 (N_29400,N_28741,N_28984);
and U29401 (N_29401,N_28073,N_28003);
and U29402 (N_29402,N_28458,N_28779);
or U29403 (N_29403,N_28062,N_28178);
nor U29404 (N_29404,N_28776,N_28111);
nand U29405 (N_29405,N_28162,N_28316);
xnor U29406 (N_29406,N_28851,N_28893);
and U29407 (N_29407,N_28864,N_28447);
and U29408 (N_29408,N_28522,N_28437);
nand U29409 (N_29409,N_28034,N_28088);
xnor U29410 (N_29410,N_28675,N_28598);
xnor U29411 (N_29411,N_28260,N_28464);
xnor U29412 (N_29412,N_28596,N_28553);
and U29413 (N_29413,N_28412,N_28427);
and U29414 (N_29414,N_28757,N_28846);
nand U29415 (N_29415,N_28771,N_28382);
xor U29416 (N_29416,N_28920,N_28784);
nand U29417 (N_29417,N_28127,N_28585);
xor U29418 (N_29418,N_28619,N_28657);
nor U29419 (N_29419,N_28384,N_28858);
or U29420 (N_29420,N_28557,N_28375);
or U29421 (N_29421,N_28151,N_28222);
nor U29422 (N_29422,N_28856,N_28506);
and U29423 (N_29423,N_28358,N_28746);
nor U29424 (N_29424,N_28009,N_28303);
or U29425 (N_29425,N_28614,N_28730);
and U29426 (N_29426,N_28719,N_28167);
nand U29427 (N_29427,N_28198,N_28912);
xor U29428 (N_29428,N_28411,N_28648);
and U29429 (N_29429,N_28745,N_28348);
nor U29430 (N_29430,N_28595,N_28257);
nand U29431 (N_29431,N_28417,N_28275);
and U29432 (N_29432,N_28863,N_28813);
nand U29433 (N_29433,N_28395,N_28202);
xnor U29434 (N_29434,N_28420,N_28197);
nor U29435 (N_29435,N_28602,N_28606);
and U29436 (N_29436,N_28299,N_28289);
xnor U29437 (N_29437,N_28027,N_28153);
and U29438 (N_29438,N_28819,N_28679);
nor U29439 (N_29439,N_28004,N_28736);
xor U29440 (N_29440,N_28968,N_28279);
and U29441 (N_29441,N_28031,N_28442);
or U29442 (N_29442,N_28549,N_28493);
nor U29443 (N_29443,N_28802,N_28870);
nand U29444 (N_29444,N_28291,N_28431);
nor U29445 (N_29445,N_28633,N_28587);
or U29446 (N_29446,N_28521,N_28528);
or U29447 (N_29447,N_28200,N_28230);
nand U29448 (N_29448,N_28336,N_28645);
nor U29449 (N_29449,N_28841,N_28005);
xnor U29450 (N_29450,N_28998,N_28238);
xor U29451 (N_29451,N_28783,N_28112);
nor U29452 (N_29452,N_28236,N_28491);
and U29453 (N_29453,N_28469,N_28910);
nor U29454 (N_29454,N_28885,N_28324);
and U29455 (N_29455,N_28916,N_28103);
nor U29456 (N_29456,N_28415,N_28735);
nand U29457 (N_29457,N_28667,N_28460);
nor U29458 (N_29458,N_28058,N_28621);
nand U29459 (N_29459,N_28215,N_28871);
nor U29460 (N_29460,N_28640,N_28660);
or U29461 (N_29461,N_28842,N_28681);
nor U29462 (N_29462,N_28510,N_28748);
xor U29463 (N_29463,N_28201,N_28187);
and U29464 (N_29464,N_28664,N_28107);
nor U29465 (N_29465,N_28177,N_28903);
xor U29466 (N_29466,N_28945,N_28997);
nand U29467 (N_29467,N_28747,N_28672);
or U29468 (N_29468,N_28066,N_28908);
nor U29469 (N_29469,N_28866,N_28796);
nand U29470 (N_29470,N_28258,N_28327);
and U29471 (N_29471,N_28782,N_28413);
or U29472 (N_29472,N_28791,N_28090);
and U29473 (N_29473,N_28394,N_28102);
or U29474 (N_29474,N_28971,N_28032);
nor U29475 (N_29475,N_28255,N_28129);
or U29476 (N_29476,N_28605,N_28709);
xor U29477 (N_29477,N_28539,N_28835);
xor U29478 (N_29478,N_28081,N_28223);
and U29479 (N_29479,N_28853,N_28429);
xnor U29480 (N_29480,N_28168,N_28043);
nand U29481 (N_29481,N_28668,N_28048);
and U29482 (N_29482,N_28576,N_28181);
nor U29483 (N_29483,N_28344,N_28002);
and U29484 (N_29484,N_28552,N_28857);
or U29485 (N_29485,N_28520,N_28318);
or U29486 (N_29486,N_28615,N_28872);
or U29487 (N_29487,N_28691,N_28368);
xor U29488 (N_29488,N_28588,N_28755);
or U29489 (N_29489,N_28244,N_28385);
or U29490 (N_29490,N_28272,N_28274);
nor U29491 (N_29491,N_28801,N_28270);
and U29492 (N_29492,N_28902,N_28170);
and U29493 (N_29493,N_28390,N_28795);
nor U29494 (N_29494,N_28811,N_28340);
nand U29495 (N_29495,N_28470,N_28373);
and U29496 (N_29496,N_28965,N_28267);
or U29497 (N_29497,N_28488,N_28542);
nand U29498 (N_29498,N_28209,N_28807);
nand U29499 (N_29499,N_28484,N_28907);
nand U29500 (N_29500,N_28095,N_28441);
nor U29501 (N_29501,N_28477,N_28821);
or U29502 (N_29502,N_28108,N_28959);
nand U29503 (N_29503,N_28915,N_28733);
nand U29504 (N_29504,N_28485,N_28025);
nor U29505 (N_29505,N_28715,N_28424);
nand U29506 (N_29506,N_28385,N_28185);
nand U29507 (N_29507,N_28245,N_28612);
xor U29508 (N_29508,N_28433,N_28004);
or U29509 (N_29509,N_28517,N_28192);
and U29510 (N_29510,N_28975,N_28899);
nor U29511 (N_29511,N_28588,N_28357);
nand U29512 (N_29512,N_28898,N_28466);
xnor U29513 (N_29513,N_28844,N_28943);
xnor U29514 (N_29514,N_28996,N_28930);
nor U29515 (N_29515,N_28840,N_28466);
xnor U29516 (N_29516,N_28230,N_28219);
xnor U29517 (N_29517,N_28988,N_28264);
nand U29518 (N_29518,N_28929,N_28293);
nor U29519 (N_29519,N_28278,N_28907);
xnor U29520 (N_29520,N_28444,N_28887);
xnor U29521 (N_29521,N_28037,N_28300);
or U29522 (N_29522,N_28201,N_28841);
nor U29523 (N_29523,N_28200,N_28608);
nand U29524 (N_29524,N_28412,N_28706);
xor U29525 (N_29525,N_28296,N_28997);
or U29526 (N_29526,N_28243,N_28612);
or U29527 (N_29527,N_28322,N_28815);
or U29528 (N_29528,N_28472,N_28848);
or U29529 (N_29529,N_28749,N_28476);
nor U29530 (N_29530,N_28239,N_28563);
and U29531 (N_29531,N_28480,N_28038);
and U29532 (N_29532,N_28816,N_28736);
and U29533 (N_29533,N_28400,N_28093);
xor U29534 (N_29534,N_28992,N_28321);
or U29535 (N_29535,N_28318,N_28587);
xor U29536 (N_29536,N_28906,N_28247);
nor U29537 (N_29537,N_28152,N_28961);
nor U29538 (N_29538,N_28432,N_28516);
and U29539 (N_29539,N_28718,N_28413);
nor U29540 (N_29540,N_28502,N_28051);
nand U29541 (N_29541,N_28024,N_28123);
xor U29542 (N_29542,N_28648,N_28271);
nand U29543 (N_29543,N_28814,N_28970);
xnor U29544 (N_29544,N_28049,N_28601);
and U29545 (N_29545,N_28375,N_28676);
xor U29546 (N_29546,N_28003,N_28297);
nand U29547 (N_29547,N_28680,N_28044);
nor U29548 (N_29548,N_28784,N_28896);
or U29549 (N_29549,N_28302,N_28483);
xor U29550 (N_29550,N_28777,N_28960);
xor U29551 (N_29551,N_28137,N_28507);
nand U29552 (N_29552,N_28100,N_28105);
xnor U29553 (N_29553,N_28334,N_28223);
xor U29554 (N_29554,N_28624,N_28847);
and U29555 (N_29555,N_28136,N_28107);
nor U29556 (N_29556,N_28021,N_28740);
and U29557 (N_29557,N_28785,N_28085);
nand U29558 (N_29558,N_28677,N_28920);
or U29559 (N_29559,N_28761,N_28624);
and U29560 (N_29560,N_28683,N_28279);
and U29561 (N_29561,N_28913,N_28185);
or U29562 (N_29562,N_28450,N_28389);
nand U29563 (N_29563,N_28676,N_28429);
or U29564 (N_29564,N_28638,N_28796);
or U29565 (N_29565,N_28293,N_28307);
or U29566 (N_29566,N_28849,N_28316);
nand U29567 (N_29567,N_28416,N_28509);
nor U29568 (N_29568,N_28618,N_28125);
and U29569 (N_29569,N_28571,N_28316);
and U29570 (N_29570,N_28313,N_28177);
or U29571 (N_29571,N_28430,N_28350);
and U29572 (N_29572,N_28329,N_28283);
nor U29573 (N_29573,N_28460,N_28303);
nor U29574 (N_29574,N_28180,N_28294);
and U29575 (N_29575,N_28241,N_28295);
nor U29576 (N_29576,N_28338,N_28201);
and U29577 (N_29577,N_28894,N_28378);
and U29578 (N_29578,N_28179,N_28988);
and U29579 (N_29579,N_28940,N_28945);
nand U29580 (N_29580,N_28264,N_28725);
or U29581 (N_29581,N_28239,N_28452);
or U29582 (N_29582,N_28549,N_28787);
and U29583 (N_29583,N_28905,N_28347);
or U29584 (N_29584,N_28272,N_28995);
or U29585 (N_29585,N_28164,N_28869);
and U29586 (N_29586,N_28131,N_28037);
and U29587 (N_29587,N_28364,N_28109);
xnor U29588 (N_29588,N_28771,N_28909);
xor U29589 (N_29589,N_28511,N_28980);
or U29590 (N_29590,N_28375,N_28286);
nand U29591 (N_29591,N_28705,N_28785);
xnor U29592 (N_29592,N_28283,N_28204);
or U29593 (N_29593,N_28258,N_28768);
nand U29594 (N_29594,N_28737,N_28010);
nand U29595 (N_29595,N_28070,N_28763);
or U29596 (N_29596,N_28792,N_28808);
xnor U29597 (N_29597,N_28504,N_28299);
or U29598 (N_29598,N_28202,N_28786);
or U29599 (N_29599,N_28381,N_28814);
nor U29600 (N_29600,N_28432,N_28985);
or U29601 (N_29601,N_28748,N_28500);
nand U29602 (N_29602,N_28815,N_28155);
nand U29603 (N_29603,N_28684,N_28051);
or U29604 (N_29604,N_28177,N_28238);
or U29605 (N_29605,N_28991,N_28089);
xnor U29606 (N_29606,N_28685,N_28270);
xnor U29607 (N_29607,N_28249,N_28810);
and U29608 (N_29608,N_28869,N_28890);
xnor U29609 (N_29609,N_28377,N_28281);
xor U29610 (N_29610,N_28137,N_28103);
nand U29611 (N_29611,N_28746,N_28372);
nor U29612 (N_29612,N_28058,N_28508);
nand U29613 (N_29613,N_28498,N_28375);
and U29614 (N_29614,N_28836,N_28828);
and U29615 (N_29615,N_28938,N_28528);
nand U29616 (N_29616,N_28201,N_28308);
nand U29617 (N_29617,N_28979,N_28485);
nand U29618 (N_29618,N_28100,N_28924);
or U29619 (N_29619,N_28339,N_28324);
nand U29620 (N_29620,N_28376,N_28418);
or U29621 (N_29621,N_28460,N_28569);
or U29622 (N_29622,N_28871,N_28048);
xnor U29623 (N_29623,N_28281,N_28600);
or U29624 (N_29624,N_28400,N_28772);
nand U29625 (N_29625,N_28198,N_28630);
nand U29626 (N_29626,N_28556,N_28852);
nand U29627 (N_29627,N_28747,N_28954);
xnor U29628 (N_29628,N_28568,N_28649);
nor U29629 (N_29629,N_28693,N_28242);
and U29630 (N_29630,N_28114,N_28612);
nand U29631 (N_29631,N_28419,N_28773);
nand U29632 (N_29632,N_28726,N_28792);
or U29633 (N_29633,N_28256,N_28031);
xor U29634 (N_29634,N_28850,N_28780);
xnor U29635 (N_29635,N_28320,N_28232);
nand U29636 (N_29636,N_28987,N_28534);
xor U29637 (N_29637,N_28760,N_28302);
and U29638 (N_29638,N_28194,N_28664);
nor U29639 (N_29639,N_28461,N_28277);
nand U29640 (N_29640,N_28239,N_28075);
xnor U29641 (N_29641,N_28729,N_28496);
nor U29642 (N_29642,N_28386,N_28429);
xnor U29643 (N_29643,N_28043,N_28276);
nor U29644 (N_29644,N_28811,N_28569);
nor U29645 (N_29645,N_28779,N_28739);
or U29646 (N_29646,N_28792,N_28449);
xor U29647 (N_29647,N_28484,N_28953);
nand U29648 (N_29648,N_28435,N_28601);
or U29649 (N_29649,N_28985,N_28772);
nand U29650 (N_29650,N_28117,N_28273);
or U29651 (N_29651,N_28181,N_28370);
and U29652 (N_29652,N_28292,N_28428);
or U29653 (N_29653,N_28750,N_28953);
xor U29654 (N_29654,N_28350,N_28832);
nand U29655 (N_29655,N_28450,N_28433);
nand U29656 (N_29656,N_28640,N_28983);
xor U29657 (N_29657,N_28290,N_28915);
nor U29658 (N_29658,N_28804,N_28234);
nand U29659 (N_29659,N_28434,N_28092);
nor U29660 (N_29660,N_28789,N_28196);
nand U29661 (N_29661,N_28046,N_28657);
nor U29662 (N_29662,N_28178,N_28598);
and U29663 (N_29663,N_28575,N_28341);
nor U29664 (N_29664,N_28110,N_28441);
xnor U29665 (N_29665,N_28668,N_28453);
and U29666 (N_29666,N_28864,N_28148);
or U29667 (N_29667,N_28666,N_28373);
xor U29668 (N_29668,N_28591,N_28823);
and U29669 (N_29669,N_28331,N_28198);
nand U29670 (N_29670,N_28641,N_28877);
or U29671 (N_29671,N_28647,N_28230);
or U29672 (N_29672,N_28748,N_28508);
and U29673 (N_29673,N_28729,N_28681);
and U29674 (N_29674,N_28839,N_28412);
xor U29675 (N_29675,N_28655,N_28842);
nand U29676 (N_29676,N_28278,N_28914);
and U29677 (N_29677,N_28776,N_28943);
and U29678 (N_29678,N_28943,N_28723);
nor U29679 (N_29679,N_28224,N_28770);
or U29680 (N_29680,N_28043,N_28356);
xnor U29681 (N_29681,N_28961,N_28904);
and U29682 (N_29682,N_28902,N_28750);
nand U29683 (N_29683,N_28246,N_28644);
or U29684 (N_29684,N_28773,N_28475);
nor U29685 (N_29685,N_28890,N_28083);
and U29686 (N_29686,N_28512,N_28636);
and U29687 (N_29687,N_28796,N_28819);
nor U29688 (N_29688,N_28543,N_28789);
xnor U29689 (N_29689,N_28694,N_28831);
xor U29690 (N_29690,N_28066,N_28310);
or U29691 (N_29691,N_28745,N_28620);
xor U29692 (N_29692,N_28519,N_28690);
and U29693 (N_29693,N_28805,N_28694);
and U29694 (N_29694,N_28199,N_28204);
nor U29695 (N_29695,N_28836,N_28660);
and U29696 (N_29696,N_28169,N_28987);
xnor U29697 (N_29697,N_28120,N_28347);
nor U29698 (N_29698,N_28071,N_28125);
and U29699 (N_29699,N_28736,N_28131);
or U29700 (N_29700,N_28651,N_28269);
and U29701 (N_29701,N_28421,N_28758);
nand U29702 (N_29702,N_28995,N_28920);
nor U29703 (N_29703,N_28301,N_28881);
or U29704 (N_29704,N_28462,N_28146);
or U29705 (N_29705,N_28964,N_28416);
xor U29706 (N_29706,N_28722,N_28427);
or U29707 (N_29707,N_28065,N_28639);
xnor U29708 (N_29708,N_28855,N_28957);
or U29709 (N_29709,N_28907,N_28936);
nor U29710 (N_29710,N_28280,N_28079);
or U29711 (N_29711,N_28102,N_28574);
and U29712 (N_29712,N_28287,N_28481);
and U29713 (N_29713,N_28035,N_28244);
or U29714 (N_29714,N_28167,N_28746);
nor U29715 (N_29715,N_28406,N_28164);
xnor U29716 (N_29716,N_28402,N_28222);
nor U29717 (N_29717,N_28168,N_28156);
nand U29718 (N_29718,N_28198,N_28445);
nor U29719 (N_29719,N_28498,N_28532);
xnor U29720 (N_29720,N_28873,N_28029);
nand U29721 (N_29721,N_28493,N_28540);
nor U29722 (N_29722,N_28847,N_28269);
nor U29723 (N_29723,N_28180,N_28103);
or U29724 (N_29724,N_28814,N_28026);
or U29725 (N_29725,N_28798,N_28315);
nor U29726 (N_29726,N_28998,N_28271);
xnor U29727 (N_29727,N_28921,N_28386);
xnor U29728 (N_29728,N_28079,N_28562);
or U29729 (N_29729,N_28028,N_28479);
and U29730 (N_29730,N_28102,N_28673);
nor U29731 (N_29731,N_28437,N_28104);
xnor U29732 (N_29732,N_28001,N_28570);
and U29733 (N_29733,N_28247,N_28447);
xor U29734 (N_29734,N_28648,N_28094);
nand U29735 (N_29735,N_28759,N_28042);
and U29736 (N_29736,N_28830,N_28046);
nor U29737 (N_29737,N_28517,N_28580);
xor U29738 (N_29738,N_28137,N_28915);
or U29739 (N_29739,N_28471,N_28418);
nand U29740 (N_29740,N_28457,N_28459);
nand U29741 (N_29741,N_28603,N_28032);
and U29742 (N_29742,N_28508,N_28962);
and U29743 (N_29743,N_28386,N_28735);
and U29744 (N_29744,N_28875,N_28401);
xor U29745 (N_29745,N_28535,N_28383);
and U29746 (N_29746,N_28094,N_28402);
xnor U29747 (N_29747,N_28176,N_28650);
nand U29748 (N_29748,N_28662,N_28519);
xor U29749 (N_29749,N_28567,N_28333);
or U29750 (N_29750,N_28610,N_28868);
nand U29751 (N_29751,N_28355,N_28915);
or U29752 (N_29752,N_28736,N_28371);
and U29753 (N_29753,N_28189,N_28662);
and U29754 (N_29754,N_28662,N_28213);
nor U29755 (N_29755,N_28903,N_28322);
nor U29756 (N_29756,N_28449,N_28172);
and U29757 (N_29757,N_28165,N_28425);
nor U29758 (N_29758,N_28408,N_28218);
nand U29759 (N_29759,N_28169,N_28291);
nor U29760 (N_29760,N_28862,N_28430);
nor U29761 (N_29761,N_28542,N_28701);
or U29762 (N_29762,N_28200,N_28193);
or U29763 (N_29763,N_28794,N_28851);
xnor U29764 (N_29764,N_28182,N_28409);
nand U29765 (N_29765,N_28017,N_28891);
nor U29766 (N_29766,N_28299,N_28265);
and U29767 (N_29767,N_28159,N_28248);
nand U29768 (N_29768,N_28002,N_28860);
nand U29769 (N_29769,N_28651,N_28422);
and U29770 (N_29770,N_28648,N_28787);
or U29771 (N_29771,N_28089,N_28687);
or U29772 (N_29772,N_28910,N_28523);
or U29773 (N_29773,N_28748,N_28195);
xnor U29774 (N_29774,N_28375,N_28844);
nor U29775 (N_29775,N_28403,N_28911);
nand U29776 (N_29776,N_28894,N_28173);
or U29777 (N_29777,N_28425,N_28404);
xor U29778 (N_29778,N_28101,N_28785);
nor U29779 (N_29779,N_28768,N_28291);
nor U29780 (N_29780,N_28396,N_28447);
xor U29781 (N_29781,N_28091,N_28361);
nand U29782 (N_29782,N_28608,N_28161);
nand U29783 (N_29783,N_28526,N_28224);
nand U29784 (N_29784,N_28863,N_28006);
or U29785 (N_29785,N_28760,N_28081);
nand U29786 (N_29786,N_28870,N_28269);
nor U29787 (N_29787,N_28808,N_28868);
nand U29788 (N_29788,N_28051,N_28058);
and U29789 (N_29789,N_28988,N_28717);
or U29790 (N_29790,N_28144,N_28161);
nand U29791 (N_29791,N_28281,N_28378);
and U29792 (N_29792,N_28430,N_28457);
nand U29793 (N_29793,N_28459,N_28860);
nand U29794 (N_29794,N_28437,N_28059);
nor U29795 (N_29795,N_28360,N_28574);
and U29796 (N_29796,N_28252,N_28965);
nor U29797 (N_29797,N_28602,N_28221);
nand U29798 (N_29798,N_28795,N_28636);
or U29799 (N_29799,N_28719,N_28138);
xor U29800 (N_29800,N_28263,N_28938);
or U29801 (N_29801,N_28964,N_28664);
xnor U29802 (N_29802,N_28219,N_28611);
nand U29803 (N_29803,N_28201,N_28362);
or U29804 (N_29804,N_28267,N_28017);
and U29805 (N_29805,N_28807,N_28015);
nor U29806 (N_29806,N_28015,N_28752);
and U29807 (N_29807,N_28227,N_28777);
or U29808 (N_29808,N_28004,N_28183);
nand U29809 (N_29809,N_28977,N_28314);
nand U29810 (N_29810,N_28218,N_28196);
and U29811 (N_29811,N_28633,N_28896);
and U29812 (N_29812,N_28772,N_28436);
or U29813 (N_29813,N_28171,N_28649);
and U29814 (N_29814,N_28820,N_28323);
and U29815 (N_29815,N_28921,N_28789);
and U29816 (N_29816,N_28299,N_28388);
and U29817 (N_29817,N_28140,N_28035);
xnor U29818 (N_29818,N_28558,N_28862);
or U29819 (N_29819,N_28910,N_28410);
and U29820 (N_29820,N_28709,N_28780);
nand U29821 (N_29821,N_28343,N_28208);
or U29822 (N_29822,N_28236,N_28830);
nand U29823 (N_29823,N_28010,N_28080);
and U29824 (N_29824,N_28827,N_28204);
nor U29825 (N_29825,N_28588,N_28659);
nor U29826 (N_29826,N_28298,N_28877);
nor U29827 (N_29827,N_28548,N_28074);
nor U29828 (N_29828,N_28411,N_28645);
and U29829 (N_29829,N_28351,N_28267);
or U29830 (N_29830,N_28375,N_28236);
xnor U29831 (N_29831,N_28569,N_28675);
nor U29832 (N_29832,N_28043,N_28013);
xnor U29833 (N_29833,N_28843,N_28624);
or U29834 (N_29834,N_28800,N_28877);
nor U29835 (N_29835,N_28278,N_28636);
nor U29836 (N_29836,N_28114,N_28951);
xnor U29837 (N_29837,N_28736,N_28002);
xor U29838 (N_29838,N_28211,N_28784);
and U29839 (N_29839,N_28904,N_28026);
and U29840 (N_29840,N_28331,N_28406);
nor U29841 (N_29841,N_28485,N_28617);
xor U29842 (N_29842,N_28695,N_28538);
or U29843 (N_29843,N_28000,N_28553);
xnor U29844 (N_29844,N_28721,N_28565);
and U29845 (N_29845,N_28948,N_28534);
or U29846 (N_29846,N_28964,N_28028);
xnor U29847 (N_29847,N_28196,N_28226);
nand U29848 (N_29848,N_28434,N_28854);
or U29849 (N_29849,N_28918,N_28763);
and U29850 (N_29850,N_28630,N_28991);
xnor U29851 (N_29851,N_28920,N_28316);
nand U29852 (N_29852,N_28266,N_28692);
or U29853 (N_29853,N_28856,N_28916);
nand U29854 (N_29854,N_28164,N_28706);
nor U29855 (N_29855,N_28379,N_28022);
and U29856 (N_29856,N_28570,N_28205);
and U29857 (N_29857,N_28189,N_28054);
or U29858 (N_29858,N_28680,N_28808);
and U29859 (N_29859,N_28732,N_28267);
xor U29860 (N_29860,N_28219,N_28467);
nor U29861 (N_29861,N_28943,N_28774);
nand U29862 (N_29862,N_28448,N_28161);
nand U29863 (N_29863,N_28119,N_28140);
and U29864 (N_29864,N_28722,N_28541);
and U29865 (N_29865,N_28197,N_28413);
nor U29866 (N_29866,N_28089,N_28092);
nand U29867 (N_29867,N_28474,N_28733);
or U29868 (N_29868,N_28252,N_28313);
or U29869 (N_29869,N_28680,N_28510);
nor U29870 (N_29870,N_28821,N_28503);
and U29871 (N_29871,N_28208,N_28757);
nor U29872 (N_29872,N_28597,N_28516);
nand U29873 (N_29873,N_28954,N_28394);
nand U29874 (N_29874,N_28365,N_28185);
nor U29875 (N_29875,N_28996,N_28048);
and U29876 (N_29876,N_28113,N_28963);
nand U29877 (N_29877,N_28352,N_28629);
or U29878 (N_29878,N_28765,N_28917);
xor U29879 (N_29879,N_28255,N_28952);
nor U29880 (N_29880,N_28504,N_28625);
and U29881 (N_29881,N_28116,N_28292);
xnor U29882 (N_29882,N_28688,N_28676);
or U29883 (N_29883,N_28793,N_28577);
or U29884 (N_29884,N_28903,N_28568);
and U29885 (N_29885,N_28821,N_28783);
nand U29886 (N_29886,N_28143,N_28853);
nand U29887 (N_29887,N_28027,N_28107);
and U29888 (N_29888,N_28519,N_28686);
nand U29889 (N_29889,N_28461,N_28653);
nor U29890 (N_29890,N_28298,N_28507);
nand U29891 (N_29891,N_28232,N_28636);
nand U29892 (N_29892,N_28339,N_28392);
nor U29893 (N_29893,N_28679,N_28537);
or U29894 (N_29894,N_28518,N_28199);
xor U29895 (N_29895,N_28472,N_28518);
or U29896 (N_29896,N_28457,N_28573);
or U29897 (N_29897,N_28758,N_28199);
xnor U29898 (N_29898,N_28168,N_28038);
nand U29899 (N_29899,N_28564,N_28943);
and U29900 (N_29900,N_28241,N_28736);
or U29901 (N_29901,N_28013,N_28562);
or U29902 (N_29902,N_28830,N_28031);
nor U29903 (N_29903,N_28335,N_28842);
nand U29904 (N_29904,N_28320,N_28433);
nand U29905 (N_29905,N_28901,N_28747);
and U29906 (N_29906,N_28302,N_28441);
and U29907 (N_29907,N_28167,N_28711);
nand U29908 (N_29908,N_28488,N_28939);
nor U29909 (N_29909,N_28711,N_28087);
or U29910 (N_29910,N_28819,N_28698);
and U29911 (N_29911,N_28877,N_28263);
or U29912 (N_29912,N_28359,N_28044);
xnor U29913 (N_29913,N_28144,N_28685);
nand U29914 (N_29914,N_28838,N_28005);
nand U29915 (N_29915,N_28759,N_28341);
nand U29916 (N_29916,N_28051,N_28204);
xor U29917 (N_29917,N_28605,N_28853);
nor U29918 (N_29918,N_28366,N_28822);
nor U29919 (N_29919,N_28878,N_28172);
and U29920 (N_29920,N_28387,N_28302);
xnor U29921 (N_29921,N_28793,N_28426);
or U29922 (N_29922,N_28175,N_28534);
or U29923 (N_29923,N_28290,N_28019);
nand U29924 (N_29924,N_28212,N_28597);
nand U29925 (N_29925,N_28271,N_28370);
nand U29926 (N_29926,N_28432,N_28202);
nor U29927 (N_29927,N_28624,N_28138);
nor U29928 (N_29928,N_28641,N_28762);
xor U29929 (N_29929,N_28873,N_28201);
and U29930 (N_29930,N_28180,N_28384);
or U29931 (N_29931,N_28561,N_28586);
or U29932 (N_29932,N_28437,N_28289);
nand U29933 (N_29933,N_28488,N_28139);
xnor U29934 (N_29934,N_28615,N_28462);
xnor U29935 (N_29935,N_28438,N_28883);
and U29936 (N_29936,N_28751,N_28422);
nor U29937 (N_29937,N_28384,N_28096);
nand U29938 (N_29938,N_28117,N_28317);
nand U29939 (N_29939,N_28409,N_28794);
and U29940 (N_29940,N_28088,N_28035);
or U29941 (N_29941,N_28130,N_28438);
and U29942 (N_29942,N_28346,N_28612);
xnor U29943 (N_29943,N_28610,N_28731);
nor U29944 (N_29944,N_28227,N_28885);
xor U29945 (N_29945,N_28248,N_28816);
nand U29946 (N_29946,N_28107,N_28592);
nor U29947 (N_29947,N_28529,N_28684);
and U29948 (N_29948,N_28702,N_28191);
or U29949 (N_29949,N_28078,N_28632);
nand U29950 (N_29950,N_28797,N_28801);
or U29951 (N_29951,N_28852,N_28157);
nor U29952 (N_29952,N_28665,N_28748);
and U29953 (N_29953,N_28143,N_28067);
and U29954 (N_29954,N_28238,N_28976);
or U29955 (N_29955,N_28591,N_28409);
and U29956 (N_29956,N_28592,N_28777);
xnor U29957 (N_29957,N_28023,N_28715);
nand U29958 (N_29958,N_28144,N_28552);
nand U29959 (N_29959,N_28432,N_28471);
nor U29960 (N_29960,N_28940,N_28231);
and U29961 (N_29961,N_28302,N_28753);
and U29962 (N_29962,N_28828,N_28776);
nor U29963 (N_29963,N_28159,N_28648);
nand U29964 (N_29964,N_28185,N_28646);
and U29965 (N_29965,N_28435,N_28370);
nor U29966 (N_29966,N_28097,N_28771);
nor U29967 (N_29967,N_28452,N_28740);
nand U29968 (N_29968,N_28695,N_28087);
and U29969 (N_29969,N_28584,N_28934);
nor U29970 (N_29970,N_28578,N_28557);
nand U29971 (N_29971,N_28305,N_28203);
xor U29972 (N_29972,N_28176,N_28211);
xnor U29973 (N_29973,N_28467,N_28754);
nor U29974 (N_29974,N_28824,N_28413);
nor U29975 (N_29975,N_28056,N_28640);
or U29976 (N_29976,N_28334,N_28677);
nor U29977 (N_29977,N_28101,N_28203);
nor U29978 (N_29978,N_28545,N_28973);
nand U29979 (N_29979,N_28312,N_28213);
xnor U29980 (N_29980,N_28676,N_28072);
xnor U29981 (N_29981,N_28613,N_28884);
and U29982 (N_29982,N_28182,N_28822);
or U29983 (N_29983,N_28860,N_28918);
xor U29984 (N_29984,N_28606,N_28491);
and U29985 (N_29985,N_28382,N_28962);
xnor U29986 (N_29986,N_28993,N_28929);
and U29987 (N_29987,N_28969,N_28476);
nor U29988 (N_29988,N_28291,N_28364);
or U29989 (N_29989,N_28572,N_28964);
or U29990 (N_29990,N_28513,N_28951);
xor U29991 (N_29991,N_28035,N_28032);
nand U29992 (N_29992,N_28915,N_28005);
or U29993 (N_29993,N_28753,N_28391);
nand U29994 (N_29994,N_28454,N_28614);
nor U29995 (N_29995,N_28056,N_28568);
or U29996 (N_29996,N_28839,N_28138);
nor U29997 (N_29997,N_28275,N_28527);
nor U29998 (N_29998,N_28648,N_28210);
nand U29999 (N_29999,N_28270,N_28901);
nor UO_0 (O_0,N_29173,N_29970);
xor UO_1 (O_1,N_29715,N_29703);
xor UO_2 (O_2,N_29522,N_29588);
or UO_3 (O_3,N_29050,N_29199);
or UO_4 (O_4,N_29143,N_29477);
and UO_5 (O_5,N_29462,N_29690);
nand UO_6 (O_6,N_29950,N_29775);
xor UO_7 (O_7,N_29138,N_29790);
xnor UO_8 (O_8,N_29268,N_29293);
or UO_9 (O_9,N_29716,N_29909);
or UO_10 (O_10,N_29398,N_29157);
and UO_11 (O_11,N_29892,N_29174);
and UO_12 (O_12,N_29917,N_29893);
and UO_13 (O_13,N_29793,N_29367);
xnor UO_14 (O_14,N_29567,N_29131);
nand UO_15 (O_15,N_29701,N_29718);
or UO_16 (O_16,N_29440,N_29558);
xnor UO_17 (O_17,N_29724,N_29511);
or UO_18 (O_18,N_29983,N_29415);
or UO_19 (O_19,N_29756,N_29659);
nor UO_20 (O_20,N_29192,N_29359);
or UO_21 (O_21,N_29871,N_29132);
nor UO_22 (O_22,N_29047,N_29602);
and UO_23 (O_23,N_29666,N_29566);
xor UO_24 (O_24,N_29817,N_29673);
nand UO_25 (O_25,N_29176,N_29260);
nor UO_26 (O_26,N_29405,N_29978);
nor UO_27 (O_27,N_29999,N_29127);
and UO_28 (O_28,N_29498,N_29752);
xor UO_29 (O_29,N_29087,N_29510);
nor UO_30 (O_30,N_29934,N_29454);
or UO_31 (O_31,N_29420,N_29707);
and UO_32 (O_32,N_29152,N_29070);
or UO_33 (O_33,N_29646,N_29579);
and UO_34 (O_34,N_29825,N_29942);
nor UO_35 (O_35,N_29532,N_29513);
or UO_36 (O_36,N_29501,N_29534);
nor UO_37 (O_37,N_29166,N_29314);
or UO_38 (O_38,N_29242,N_29134);
or UO_39 (O_39,N_29841,N_29241);
or UO_40 (O_40,N_29280,N_29903);
xor UO_41 (O_41,N_29486,N_29472);
nor UO_42 (O_42,N_29447,N_29966);
nor UO_43 (O_43,N_29740,N_29239);
and UO_44 (O_44,N_29652,N_29044);
xor UO_45 (O_45,N_29717,N_29451);
nand UO_46 (O_46,N_29614,N_29749);
and UO_47 (O_47,N_29834,N_29973);
and UO_48 (O_48,N_29130,N_29880);
nor UO_49 (O_49,N_29720,N_29337);
and UO_50 (O_50,N_29212,N_29678);
nor UO_51 (O_51,N_29040,N_29041);
xnor UO_52 (O_52,N_29581,N_29133);
and UO_53 (O_53,N_29918,N_29531);
xor UO_54 (O_54,N_29615,N_29661);
xor UO_55 (O_55,N_29591,N_29100);
nand UO_56 (O_56,N_29782,N_29453);
nor UO_57 (O_57,N_29304,N_29037);
nand UO_58 (O_58,N_29598,N_29020);
nor UO_59 (O_59,N_29855,N_29623);
nor UO_60 (O_60,N_29524,N_29657);
nand UO_61 (O_61,N_29948,N_29267);
nor UO_62 (O_62,N_29912,N_29866);
and UO_63 (O_63,N_29111,N_29468);
or UO_64 (O_64,N_29504,N_29290);
xnor UO_65 (O_65,N_29497,N_29992);
nand UO_66 (O_66,N_29874,N_29882);
and UO_67 (O_67,N_29021,N_29901);
nand UO_68 (O_68,N_29746,N_29951);
and UO_69 (O_69,N_29119,N_29117);
nand UO_70 (O_70,N_29237,N_29785);
nor UO_71 (O_71,N_29364,N_29265);
or UO_72 (O_72,N_29988,N_29734);
and UO_73 (O_73,N_29272,N_29147);
xor UO_74 (O_74,N_29629,N_29739);
xnor UO_75 (O_75,N_29537,N_29180);
or UO_76 (O_76,N_29528,N_29024);
and UO_77 (O_77,N_29608,N_29484);
nand UO_78 (O_78,N_29234,N_29853);
nor UO_79 (O_79,N_29109,N_29630);
and UO_80 (O_80,N_29419,N_29190);
nor UO_81 (O_81,N_29677,N_29339);
nand UO_82 (O_82,N_29936,N_29676);
xnor UO_83 (O_83,N_29927,N_29075);
or UO_84 (O_84,N_29601,N_29327);
nand UO_85 (O_85,N_29159,N_29023);
xor UO_86 (O_86,N_29164,N_29395);
and UO_87 (O_87,N_29812,N_29307);
nor UO_88 (O_88,N_29654,N_29081);
or UO_89 (O_89,N_29034,N_29953);
xor UO_90 (O_90,N_29368,N_29595);
nand UO_91 (O_91,N_29742,N_29474);
and UO_92 (O_92,N_29637,N_29492);
or UO_93 (O_93,N_29848,N_29162);
xnor UO_94 (O_94,N_29665,N_29198);
nor UO_95 (O_95,N_29895,N_29362);
and UO_96 (O_96,N_29888,N_29064);
xnor UO_97 (O_97,N_29755,N_29252);
nand UO_98 (O_98,N_29305,N_29792);
xnor UO_99 (O_99,N_29672,N_29007);
or UO_100 (O_100,N_29429,N_29799);
or UO_101 (O_101,N_29392,N_29435);
nand UO_102 (O_102,N_29406,N_29128);
nor UO_103 (O_103,N_29827,N_29698);
nand UO_104 (O_104,N_29046,N_29270);
nor UO_105 (O_105,N_29643,N_29886);
xor UO_106 (O_106,N_29771,N_29979);
nand UO_107 (O_107,N_29606,N_29025);
nand UO_108 (O_108,N_29292,N_29923);
and UO_109 (O_109,N_29332,N_29609);
or UO_110 (O_110,N_29674,N_29906);
nor UO_111 (O_111,N_29964,N_29926);
xor UO_112 (O_112,N_29358,N_29471);
xnor UO_113 (O_113,N_29692,N_29165);
and UO_114 (O_114,N_29911,N_29269);
xor UO_115 (O_115,N_29095,N_29053);
and UO_116 (O_116,N_29779,N_29894);
or UO_117 (O_117,N_29865,N_29493);
nor UO_118 (O_118,N_29938,N_29705);
or UO_119 (O_119,N_29441,N_29377);
nor UO_120 (O_120,N_29163,N_29431);
xor UO_121 (O_121,N_29517,N_29306);
nor UO_122 (O_122,N_29660,N_29264);
or UO_123 (O_123,N_29129,N_29092);
xnor UO_124 (O_124,N_29215,N_29640);
xnor UO_125 (O_125,N_29481,N_29899);
nor UO_126 (O_126,N_29506,N_29153);
nand UO_127 (O_127,N_29838,N_29709);
and UO_128 (O_128,N_29846,N_29299);
nor UO_129 (O_129,N_29479,N_29748);
xnor UO_130 (O_130,N_29971,N_29059);
and UO_131 (O_131,N_29571,N_29150);
nor UO_132 (O_132,N_29266,N_29340);
nor UO_133 (O_133,N_29905,N_29250);
or UO_134 (O_134,N_29738,N_29787);
nor UO_135 (O_135,N_29551,N_29283);
or UO_136 (O_136,N_29536,N_29663);
or UO_137 (O_137,N_29777,N_29578);
nand UO_138 (O_138,N_29177,N_29960);
nand UO_139 (O_139,N_29155,N_29586);
nor UO_140 (O_140,N_29937,N_29750);
xnor UO_141 (O_141,N_29671,N_29208);
nand UO_142 (O_142,N_29885,N_29255);
nor UO_143 (O_143,N_29301,N_29388);
and UO_144 (O_144,N_29636,N_29769);
nor UO_145 (O_145,N_29104,N_29074);
or UO_146 (O_146,N_29508,N_29038);
and UO_147 (O_147,N_29699,N_29600);
or UO_148 (O_148,N_29071,N_29488);
and UO_149 (O_149,N_29017,N_29743);
nor UO_150 (O_150,N_29965,N_29554);
xnor UO_151 (O_151,N_29114,N_29689);
nand UO_152 (O_152,N_29030,N_29116);
and UO_153 (O_153,N_29669,N_29085);
nor UO_154 (O_154,N_29353,N_29653);
nand UO_155 (O_155,N_29596,N_29914);
xor UO_156 (O_156,N_29325,N_29010);
nor UO_157 (O_157,N_29655,N_29113);
nor UO_158 (O_158,N_29158,N_29967);
nor UO_159 (O_159,N_29490,N_29712);
and UO_160 (O_160,N_29188,N_29794);
or UO_161 (O_161,N_29930,N_29557);
nor UO_162 (O_162,N_29857,N_29438);
nand UO_163 (O_163,N_29704,N_29137);
and UO_164 (O_164,N_29470,N_29329);
xnor UO_165 (O_165,N_29922,N_29572);
nand UO_166 (O_166,N_29410,N_29338);
or UO_167 (O_167,N_29594,N_29357);
nand UO_168 (O_168,N_29311,N_29144);
nor UO_169 (O_169,N_29804,N_29246);
or UO_170 (O_170,N_29231,N_29390);
nor UO_171 (O_171,N_29284,N_29317);
xnor UO_172 (O_172,N_29887,N_29366);
or UO_173 (O_173,N_29076,N_29754);
and UO_174 (O_174,N_29651,N_29621);
or UO_175 (O_175,N_29184,N_29385);
and UO_176 (O_176,N_29725,N_29422);
and UO_177 (O_177,N_29316,N_29574);
nand UO_178 (O_178,N_29956,N_29428);
nand UO_179 (O_179,N_29816,N_29500);
and UO_180 (O_180,N_29220,N_29618);
xnor UO_181 (O_181,N_29205,N_29530);
nor UO_182 (O_182,N_29919,N_29759);
nand UO_183 (O_183,N_29765,N_29171);
or UO_184 (O_184,N_29226,N_29460);
xor UO_185 (O_185,N_29313,N_29969);
xor UO_186 (O_186,N_29613,N_29943);
and UO_187 (O_187,N_29457,N_29360);
nor UO_188 (O_188,N_29344,N_29788);
nor UO_189 (O_189,N_29962,N_29619);
or UO_190 (O_190,N_29694,N_29802);
nand UO_191 (O_191,N_29624,N_29580);
xnor UO_192 (O_192,N_29032,N_29123);
or UO_193 (O_193,N_29604,N_29945);
nor UO_194 (O_194,N_29328,N_29274);
or UO_195 (O_195,N_29809,N_29638);
or UO_196 (O_196,N_29444,N_29737);
nor UO_197 (O_197,N_29346,N_29256);
nor UO_198 (O_198,N_29741,N_29631);
nor UO_199 (O_199,N_29170,N_29529);
nor UO_200 (O_200,N_29456,N_29278);
xnor UO_201 (O_201,N_29503,N_29569);
and UO_202 (O_202,N_29214,N_29875);
nand UO_203 (O_203,N_29459,N_29112);
and UO_204 (O_204,N_29458,N_29288);
nand UO_205 (O_205,N_29480,N_29203);
nand UO_206 (O_206,N_29279,N_29763);
or UO_207 (O_207,N_29535,N_29461);
or UO_208 (O_208,N_29001,N_29982);
xor UO_209 (O_209,N_29079,N_29625);
or UO_210 (O_210,N_29191,N_29251);
xnor UO_211 (O_211,N_29281,N_29560);
xnor UO_212 (O_212,N_29858,N_29731);
nand UO_213 (O_213,N_29373,N_29248);
nand UO_214 (O_214,N_29641,N_29455);
xor UO_215 (O_215,N_29876,N_29867);
nand UO_216 (O_216,N_29401,N_29706);
or UO_217 (O_217,N_29412,N_29944);
nor UO_218 (O_218,N_29042,N_29797);
or UO_219 (O_219,N_29411,N_29464);
nor UO_220 (O_220,N_29240,N_29686);
and UO_221 (O_221,N_29175,N_29400);
nor UO_222 (O_222,N_29000,N_29142);
nor UO_223 (O_223,N_29975,N_29448);
xnor UO_224 (O_224,N_29393,N_29820);
or UO_225 (O_225,N_29648,N_29378);
nor UO_226 (O_226,N_29642,N_29544);
or UO_227 (O_227,N_29181,N_29016);
xor UO_228 (O_228,N_29423,N_29218);
or UO_229 (O_229,N_29370,N_29852);
nor UO_230 (O_230,N_29986,N_29118);
xnor UO_231 (O_231,N_29276,N_29997);
or UO_232 (O_232,N_29872,N_29335);
and UO_233 (O_233,N_29418,N_29102);
or UO_234 (O_234,N_29012,N_29682);
nand UO_235 (O_235,N_29045,N_29907);
and UO_236 (O_236,N_29526,N_29347);
nor UO_237 (O_237,N_29968,N_29487);
nor UO_238 (O_238,N_29784,N_29634);
or UO_239 (O_239,N_29210,N_29683);
and UO_240 (O_240,N_29519,N_29424);
and UO_241 (O_241,N_29568,N_29597);
and UO_242 (O_242,N_29476,N_29576);
nor UO_243 (O_243,N_29097,N_29667);
or UO_244 (O_244,N_29172,N_29201);
nand UO_245 (O_245,N_29403,N_29949);
xnor UO_246 (O_246,N_29178,N_29696);
nand UO_247 (O_247,N_29900,N_29931);
nor UO_248 (O_248,N_29387,N_29196);
nor UO_249 (O_249,N_29854,N_29577);
xnor UO_250 (O_250,N_29849,N_29326);
xnor UO_251 (O_251,N_29099,N_29620);
or UO_252 (O_252,N_29722,N_29323);
and UO_253 (O_253,N_29094,N_29297);
nand UO_254 (O_254,N_29776,N_29015);
nor UO_255 (O_255,N_29285,N_29679);
and UO_256 (O_256,N_29592,N_29959);
and UO_257 (O_257,N_29995,N_29213);
and UO_258 (O_258,N_29286,N_29881);
or UO_259 (O_259,N_29889,N_29515);
or UO_260 (O_260,N_29238,N_29446);
or UO_261 (O_261,N_29209,N_29300);
and UO_262 (O_262,N_29920,N_29691);
nor UO_263 (O_263,N_29502,N_29548);
xnor UO_264 (O_264,N_29236,N_29126);
and UO_265 (O_265,N_29382,N_29110);
nand UO_266 (O_266,N_29584,N_29189);
and UO_267 (O_267,N_29467,N_29421);
and UO_268 (O_268,N_29507,N_29434);
or UO_269 (O_269,N_29303,N_29735);
xor UO_270 (O_270,N_29088,N_29869);
xor UO_271 (O_271,N_29851,N_29216);
or UO_272 (O_272,N_29713,N_29702);
and UO_273 (O_273,N_29253,N_29668);
and UO_274 (O_274,N_29573,N_29541);
nor UO_275 (O_275,N_29947,N_29331);
xor UO_276 (O_276,N_29491,N_29320);
xor UO_277 (O_277,N_29773,N_29829);
nor UO_278 (O_278,N_29389,N_29553);
and UO_279 (O_279,N_29902,N_29984);
xor UO_280 (O_280,N_29146,N_29107);
nand UO_281 (O_281,N_29538,N_29844);
xor UO_282 (O_282,N_29719,N_29167);
and UO_283 (O_283,N_29605,N_29427);
xnor UO_284 (O_284,N_29879,N_29469);
or UO_285 (O_285,N_29334,N_29224);
xor UO_286 (O_286,N_29426,N_29206);
xnor UO_287 (O_287,N_29980,N_29235);
nand UO_288 (O_288,N_29863,N_29414);
or UO_289 (O_289,N_29589,N_29994);
xor UO_290 (O_290,N_29835,N_29258);
and UO_291 (O_291,N_29772,N_29145);
and UO_292 (O_292,N_29148,N_29559);
and UO_293 (O_293,N_29952,N_29022);
and UO_294 (O_294,N_29760,N_29744);
nor UO_295 (O_295,N_29375,N_29897);
nor UO_296 (O_296,N_29836,N_29381);
nand UO_297 (O_297,N_29068,N_29352);
and UO_298 (O_298,N_29033,N_29080);
xnor UO_299 (O_299,N_29048,N_29439);
nand UO_300 (O_300,N_29687,N_29321);
nand UO_301 (O_301,N_29254,N_29302);
xor UO_302 (O_302,N_29814,N_29774);
xnor UO_303 (O_303,N_29018,N_29108);
nand UO_304 (O_304,N_29379,N_29028);
and UO_305 (O_305,N_29413,N_29842);
xnor UO_306 (O_306,N_29607,N_29154);
xnor UO_307 (O_307,N_29807,N_29204);
nand UO_308 (O_308,N_29060,N_29309);
nor UO_309 (O_309,N_29402,N_29525);
and UO_310 (O_310,N_29222,N_29977);
xor UO_311 (O_311,N_29921,N_29991);
xor UO_312 (O_312,N_29437,N_29394);
nor UO_313 (O_313,N_29860,N_29729);
nand UO_314 (O_314,N_29005,N_29761);
nand UO_315 (O_315,N_29996,N_29442);
nand UO_316 (O_316,N_29898,N_29228);
and UO_317 (O_317,N_29859,N_29533);
or UO_318 (O_318,N_29289,N_29417);
nor UO_319 (O_319,N_29485,N_29732);
xnor UO_320 (O_320,N_29801,N_29014);
or UO_321 (O_321,N_29436,N_29564);
nor UO_322 (O_322,N_29751,N_29870);
nor UO_323 (O_323,N_29027,N_29850);
and UO_324 (O_324,N_29925,N_29628);
nor UO_325 (O_325,N_29818,N_29067);
nand UO_326 (O_326,N_29940,N_29561);
or UO_327 (O_327,N_29839,N_29475);
or UO_328 (O_328,N_29728,N_29026);
xor UO_329 (O_329,N_29408,N_29399);
nor UO_330 (O_330,N_29249,N_29257);
xor UO_331 (O_331,N_29055,N_29681);
xnor UO_332 (O_332,N_29861,N_29345);
xnor UO_333 (O_333,N_29006,N_29463);
nand UO_334 (O_334,N_29932,N_29710);
and UO_335 (O_335,N_29031,N_29680);
or UO_336 (O_336,N_29009,N_29430);
nor UO_337 (O_337,N_29599,N_29450);
nand UO_338 (O_338,N_29976,N_29611);
nor UO_339 (O_339,N_29063,N_29726);
xor UO_340 (O_340,N_29610,N_29120);
nand UO_341 (O_341,N_29185,N_29416);
nor UO_342 (O_342,N_29639,N_29091);
nor UO_343 (O_343,N_29523,N_29082);
nor UO_344 (O_344,N_29404,N_29974);
or UO_345 (O_345,N_29847,N_29065);
xor UO_346 (O_346,N_29904,N_29354);
nand UO_347 (O_347,N_29374,N_29545);
nand UO_348 (O_348,N_29520,N_29333);
and UO_349 (O_349,N_29550,N_29813);
nand UO_350 (O_350,N_29089,N_29941);
nor UO_351 (O_351,N_29106,N_29590);
and UO_352 (O_352,N_29229,N_29685);
or UO_353 (O_353,N_29407,N_29518);
nor UO_354 (O_354,N_29277,N_29695);
and UO_355 (O_355,N_29585,N_29105);
nand UO_356 (O_356,N_29318,N_29336);
nand UO_357 (O_357,N_29232,N_29616);
and UO_358 (O_358,N_29808,N_29197);
or UO_359 (O_359,N_29987,N_29489);
and UO_360 (O_360,N_29961,N_29753);
and UO_361 (O_361,N_29527,N_29371);
nand UO_362 (O_362,N_29350,N_29243);
or UO_363 (O_363,N_29294,N_29939);
xnor UO_364 (O_364,N_29650,N_29824);
nor UO_365 (O_365,N_29202,N_29833);
nand UO_366 (O_366,N_29565,N_29062);
xor UO_367 (O_367,N_29139,N_29084);
nand UO_368 (O_368,N_29946,N_29054);
and UO_369 (O_369,N_29322,N_29182);
xor UO_370 (O_370,N_29466,N_29617);
nor UO_371 (O_371,N_29140,N_29372);
nand UO_372 (O_372,N_29308,N_29822);
xnor UO_373 (O_373,N_29521,N_29896);
and UO_374 (O_374,N_29831,N_29840);
nor UO_375 (O_375,N_29622,N_29051);
or UO_376 (O_376,N_29330,N_29873);
and UO_377 (O_377,N_29764,N_29815);
nand UO_378 (O_378,N_29432,N_29002);
xnor UO_379 (O_379,N_29662,N_29004);
and UO_380 (O_380,N_29073,N_29386);
nor UO_381 (O_381,N_29445,N_29090);
nand UO_382 (O_382,N_29928,N_29179);
nor UO_383 (O_383,N_29539,N_29342);
and UO_384 (O_384,N_29786,N_29298);
nor UO_385 (O_385,N_29633,N_29778);
nand UO_386 (O_386,N_29494,N_29365);
and UO_387 (O_387,N_29056,N_29916);
nor UO_388 (O_388,N_29384,N_29391);
and UO_389 (O_389,N_29800,N_29711);
or UO_390 (O_390,N_29708,N_29160);
or UO_391 (O_391,N_29658,N_29066);
or UO_392 (O_392,N_29910,N_29791);
nor UO_393 (O_393,N_29555,N_29396);
xor UO_394 (O_394,N_29890,N_29884);
nor UO_395 (O_395,N_29811,N_29649);
or UO_396 (O_396,N_29098,N_29093);
xor UO_397 (O_397,N_29259,N_29187);
and UO_398 (O_398,N_29540,N_29183);
xor UO_399 (O_399,N_29443,N_29324);
nand UO_400 (O_400,N_29862,N_29828);
nor UO_401 (O_401,N_29409,N_29496);
and UO_402 (O_402,N_29913,N_29972);
and UO_403 (O_403,N_29039,N_29798);
nand UO_404 (O_404,N_29096,N_29013);
xnor UO_405 (O_405,N_29803,N_29837);
nand UO_406 (O_406,N_29036,N_29125);
nor UO_407 (O_407,N_29355,N_29747);
and UO_408 (O_408,N_29758,N_29688);
nand UO_409 (O_409,N_29124,N_29733);
nand UO_410 (O_410,N_29603,N_29425);
and UO_411 (O_411,N_29727,N_29168);
or UO_412 (O_412,N_29263,N_29547);
or UO_413 (O_413,N_29796,N_29343);
nor UO_414 (O_414,N_29512,N_29762);
nand UO_415 (O_415,N_29644,N_29052);
xnor UO_416 (O_416,N_29086,N_29954);
nand UO_417 (O_417,N_29356,N_29819);
nor UO_418 (O_418,N_29767,N_29647);
nor UO_419 (O_419,N_29832,N_29575);
or UO_420 (O_420,N_29981,N_29227);
nor UO_421 (O_421,N_29245,N_29868);
and UO_422 (O_422,N_29989,N_29693);
nor UO_423 (O_423,N_29582,N_29101);
and UO_424 (O_424,N_29626,N_29826);
nand UO_425 (O_425,N_29675,N_29736);
or UO_426 (O_426,N_29998,N_29656);
xor UO_427 (O_427,N_29883,N_29194);
nand UO_428 (O_428,N_29349,N_29008);
xor UO_429 (O_429,N_29856,N_29217);
and UO_430 (O_430,N_29878,N_29632);
nand UO_431 (O_431,N_29273,N_29935);
nor UO_432 (O_432,N_29223,N_29233);
nor UO_433 (O_433,N_29282,N_29549);
nand UO_434 (O_434,N_29287,N_29122);
and UO_435 (O_435,N_29563,N_29211);
and UO_436 (O_436,N_29985,N_29003);
nor UO_437 (O_437,N_29019,N_29593);
nor UO_438 (O_438,N_29546,N_29664);
xnor UO_439 (O_439,N_29781,N_29810);
xnor UO_440 (O_440,N_29035,N_29823);
xor UO_441 (O_441,N_29516,N_29509);
nor UO_442 (O_442,N_29169,N_29806);
nand UO_443 (O_443,N_29433,N_29957);
xor UO_444 (O_444,N_29730,N_29141);
or UO_445 (O_445,N_29363,N_29587);
nor UO_446 (O_446,N_29029,N_29864);
or UO_447 (O_447,N_29635,N_29193);
nand UO_448 (O_448,N_29583,N_29247);
or UO_449 (O_449,N_29136,N_29291);
xor UO_450 (O_450,N_29369,N_29542);
or UO_451 (O_451,N_29993,N_29310);
nand UO_452 (O_452,N_29543,N_29058);
xor UO_453 (O_453,N_29780,N_29670);
and UO_454 (O_454,N_29383,N_29700);
or UO_455 (O_455,N_29478,N_29495);
nand UO_456 (O_456,N_29697,N_29958);
xor UO_457 (O_457,N_29312,N_29115);
or UO_458 (O_458,N_29221,N_29877);
nor UO_459 (O_459,N_29845,N_29514);
nor UO_460 (O_460,N_29376,N_29348);
nor UO_461 (O_461,N_29151,N_29195);
nor UO_462 (O_462,N_29830,N_29078);
nor UO_463 (O_463,N_29465,N_29380);
nor UO_464 (O_464,N_29319,N_29721);
nand UO_465 (O_465,N_29083,N_29933);
or UO_466 (O_466,N_29505,N_29295);
nand UO_467 (O_467,N_29135,N_29121);
or UO_468 (O_468,N_29341,N_29908);
or UO_469 (O_469,N_29990,N_29011);
or UO_470 (O_470,N_29103,N_29452);
nor UO_471 (O_471,N_29244,N_29766);
nand UO_472 (O_472,N_29482,N_29397);
nand UO_473 (O_473,N_29200,N_29315);
and UO_474 (O_474,N_29473,N_29219);
nand UO_475 (O_475,N_29556,N_29061);
nand UO_476 (O_476,N_29072,N_29570);
nand UO_477 (O_477,N_29077,N_29261);
and UO_478 (O_478,N_29795,N_29149);
nor UO_479 (O_479,N_29723,N_29271);
or UO_480 (O_480,N_29296,N_29768);
and UO_481 (O_481,N_29361,N_29963);
nand UO_482 (O_482,N_29924,N_29351);
and UO_483 (O_483,N_29186,N_29499);
nand UO_484 (O_484,N_29230,N_29745);
and UO_485 (O_485,N_29627,N_29714);
and UO_486 (O_486,N_29043,N_29843);
xor UO_487 (O_487,N_29262,N_29770);
nand UO_488 (O_488,N_29483,N_29684);
nor UO_489 (O_489,N_29275,N_29757);
or UO_490 (O_490,N_29225,N_29161);
nor UO_491 (O_491,N_29207,N_29929);
or UO_492 (O_492,N_29955,N_29821);
nand UO_493 (O_493,N_29552,N_29805);
nand UO_494 (O_494,N_29783,N_29449);
nor UO_495 (O_495,N_29891,N_29915);
or UO_496 (O_496,N_29612,N_29069);
nand UO_497 (O_497,N_29562,N_29645);
nand UO_498 (O_498,N_29789,N_29049);
xor UO_499 (O_499,N_29057,N_29156);
xnor UO_500 (O_500,N_29667,N_29310);
nand UO_501 (O_501,N_29699,N_29655);
or UO_502 (O_502,N_29461,N_29121);
or UO_503 (O_503,N_29619,N_29623);
nor UO_504 (O_504,N_29083,N_29343);
nand UO_505 (O_505,N_29026,N_29134);
nor UO_506 (O_506,N_29894,N_29202);
or UO_507 (O_507,N_29255,N_29525);
nand UO_508 (O_508,N_29066,N_29188);
nor UO_509 (O_509,N_29514,N_29804);
and UO_510 (O_510,N_29306,N_29036);
nand UO_511 (O_511,N_29865,N_29975);
xnor UO_512 (O_512,N_29881,N_29484);
nand UO_513 (O_513,N_29981,N_29095);
and UO_514 (O_514,N_29576,N_29046);
xor UO_515 (O_515,N_29839,N_29169);
nor UO_516 (O_516,N_29879,N_29453);
and UO_517 (O_517,N_29621,N_29473);
nor UO_518 (O_518,N_29433,N_29707);
or UO_519 (O_519,N_29280,N_29742);
nand UO_520 (O_520,N_29709,N_29089);
xor UO_521 (O_521,N_29758,N_29750);
nor UO_522 (O_522,N_29013,N_29681);
and UO_523 (O_523,N_29427,N_29131);
xor UO_524 (O_524,N_29121,N_29955);
xor UO_525 (O_525,N_29845,N_29008);
or UO_526 (O_526,N_29917,N_29757);
and UO_527 (O_527,N_29379,N_29309);
xnor UO_528 (O_528,N_29458,N_29086);
nor UO_529 (O_529,N_29820,N_29744);
nor UO_530 (O_530,N_29287,N_29170);
and UO_531 (O_531,N_29567,N_29265);
or UO_532 (O_532,N_29056,N_29151);
nor UO_533 (O_533,N_29873,N_29985);
xnor UO_534 (O_534,N_29665,N_29925);
or UO_535 (O_535,N_29888,N_29238);
and UO_536 (O_536,N_29923,N_29045);
nor UO_537 (O_537,N_29984,N_29607);
xor UO_538 (O_538,N_29878,N_29578);
xnor UO_539 (O_539,N_29780,N_29660);
xor UO_540 (O_540,N_29458,N_29720);
and UO_541 (O_541,N_29166,N_29858);
nand UO_542 (O_542,N_29049,N_29513);
xnor UO_543 (O_543,N_29866,N_29684);
nor UO_544 (O_544,N_29434,N_29611);
or UO_545 (O_545,N_29388,N_29498);
nand UO_546 (O_546,N_29299,N_29392);
xnor UO_547 (O_547,N_29253,N_29256);
nor UO_548 (O_548,N_29441,N_29013);
xor UO_549 (O_549,N_29595,N_29674);
and UO_550 (O_550,N_29253,N_29645);
xor UO_551 (O_551,N_29913,N_29197);
nor UO_552 (O_552,N_29844,N_29960);
xnor UO_553 (O_553,N_29796,N_29762);
or UO_554 (O_554,N_29027,N_29491);
nor UO_555 (O_555,N_29566,N_29509);
and UO_556 (O_556,N_29083,N_29650);
nor UO_557 (O_557,N_29875,N_29586);
nand UO_558 (O_558,N_29979,N_29209);
nand UO_559 (O_559,N_29612,N_29811);
and UO_560 (O_560,N_29646,N_29180);
and UO_561 (O_561,N_29929,N_29118);
nand UO_562 (O_562,N_29811,N_29404);
and UO_563 (O_563,N_29718,N_29189);
or UO_564 (O_564,N_29623,N_29471);
nor UO_565 (O_565,N_29119,N_29825);
and UO_566 (O_566,N_29044,N_29724);
or UO_567 (O_567,N_29481,N_29405);
nor UO_568 (O_568,N_29892,N_29858);
nand UO_569 (O_569,N_29398,N_29551);
or UO_570 (O_570,N_29289,N_29437);
or UO_571 (O_571,N_29318,N_29377);
and UO_572 (O_572,N_29656,N_29018);
and UO_573 (O_573,N_29932,N_29985);
or UO_574 (O_574,N_29190,N_29644);
or UO_575 (O_575,N_29012,N_29171);
nor UO_576 (O_576,N_29208,N_29597);
nor UO_577 (O_577,N_29445,N_29764);
or UO_578 (O_578,N_29563,N_29352);
nor UO_579 (O_579,N_29698,N_29552);
nand UO_580 (O_580,N_29106,N_29414);
nor UO_581 (O_581,N_29354,N_29297);
and UO_582 (O_582,N_29914,N_29929);
nor UO_583 (O_583,N_29201,N_29462);
xnor UO_584 (O_584,N_29258,N_29314);
nand UO_585 (O_585,N_29390,N_29931);
nand UO_586 (O_586,N_29335,N_29420);
xnor UO_587 (O_587,N_29518,N_29553);
xor UO_588 (O_588,N_29043,N_29841);
nand UO_589 (O_589,N_29683,N_29365);
nor UO_590 (O_590,N_29150,N_29468);
nor UO_591 (O_591,N_29366,N_29815);
or UO_592 (O_592,N_29738,N_29725);
and UO_593 (O_593,N_29571,N_29492);
nand UO_594 (O_594,N_29776,N_29423);
nand UO_595 (O_595,N_29767,N_29617);
and UO_596 (O_596,N_29500,N_29059);
and UO_597 (O_597,N_29142,N_29248);
or UO_598 (O_598,N_29395,N_29768);
and UO_599 (O_599,N_29974,N_29386);
and UO_600 (O_600,N_29877,N_29520);
or UO_601 (O_601,N_29153,N_29923);
nand UO_602 (O_602,N_29738,N_29656);
and UO_603 (O_603,N_29578,N_29169);
nor UO_604 (O_604,N_29568,N_29920);
xor UO_605 (O_605,N_29435,N_29197);
xor UO_606 (O_606,N_29572,N_29924);
xnor UO_607 (O_607,N_29578,N_29050);
nand UO_608 (O_608,N_29957,N_29094);
xnor UO_609 (O_609,N_29357,N_29792);
and UO_610 (O_610,N_29177,N_29534);
and UO_611 (O_611,N_29968,N_29408);
nand UO_612 (O_612,N_29893,N_29721);
xnor UO_613 (O_613,N_29176,N_29047);
nand UO_614 (O_614,N_29372,N_29476);
nand UO_615 (O_615,N_29080,N_29274);
or UO_616 (O_616,N_29063,N_29222);
or UO_617 (O_617,N_29198,N_29822);
nand UO_618 (O_618,N_29386,N_29533);
nand UO_619 (O_619,N_29552,N_29048);
and UO_620 (O_620,N_29417,N_29890);
nor UO_621 (O_621,N_29210,N_29733);
and UO_622 (O_622,N_29982,N_29444);
xnor UO_623 (O_623,N_29081,N_29679);
nand UO_624 (O_624,N_29911,N_29275);
nor UO_625 (O_625,N_29263,N_29129);
or UO_626 (O_626,N_29742,N_29595);
xor UO_627 (O_627,N_29904,N_29327);
nor UO_628 (O_628,N_29735,N_29577);
nand UO_629 (O_629,N_29925,N_29669);
or UO_630 (O_630,N_29414,N_29891);
xor UO_631 (O_631,N_29010,N_29719);
and UO_632 (O_632,N_29445,N_29606);
or UO_633 (O_633,N_29621,N_29919);
xor UO_634 (O_634,N_29784,N_29172);
nand UO_635 (O_635,N_29485,N_29351);
or UO_636 (O_636,N_29256,N_29456);
xnor UO_637 (O_637,N_29156,N_29335);
nor UO_638 (O_638,N_29243,N_29919);
or UO_639 (O_639,N_29698,N_29163);
and UO_640 (O_640,N_29107,N_29172);
xor UO_641 (O_641,N_29483,N_29463);
or UO_642 (O_642,N_29839,N_29147);
or UO_643 (O_643,N_29932,N_29278);
or UO_644 (O_644,N_29820,N_29707);
nand UO_645 (O_645,N_29449,N_29215);
and UO_646 (O_646,N_29234,N_29302);
nand UO_647 (O_647,N_29441,N_29784);
nor UO_648 (O_648,N_29833,N_29822);
nand UO_649 (O_649,N_29023,N_29155);
xnor UO_650 (O_650,N_29564,N_29931);
and UO_651 (O_651,N_29880,N_29968);
nand UO_652 (O_652,N_29608,N_29028);
nand UO_653 (O_653,N_29161,N_29075);
or UO_654 (O_654,N_29188,N_29532);
nand UO_655 (O_655,N_29212,N_29585);
or UO_656 (O_656,N_29144,N_29021);
nand UO_657 (O_657,N_29164,N_29592);
and UO_658 (O_658,N_29377,N_29518);
nand UO_659 (O_659,N_29630,N_29672);
nor UO_660 (O_660,N_29482,N_29393);
and UO_661 (O_661,N_29439,N_29482);
xnor UO_662 (O_662,N_29310,N_29679);
nor UO_663 (O_663,N_29568,N_29792);
nor UO_664 (O_664,N_29914,N_29562);
nand UO_665 (O_665,N_29897,N_29076);
nand UO_666 (O_666,N_29966,N_29713);
nor UO_667 (O_667,N_29251,N_29891);
nor UO_668 (O_668,N_29919,N_29566);
xnor UO_669 (O_669,N_29301,N_29500);
nand UO_670 (O_670,N_29264,N_29772);
nand UO_671 (O_671,N_29542,N_29212);
and UO_672 (O_672,N_29290,N_29214);
xnor UO_673 (O_673,N_29693,N_29237);
nor UO_674 (O_674,N_29013,N_29141);
nor UO_675 (O_675,N_29682,N_29401);
and UO_676 (O_676,N_29674,N_29447);
xnor UO_677 (O_677,N_29007,N_29442);
nor UO_678 (O_678,N_29594,N_29443);
and UO_679 (O_679,N_29598,N_29538);
nand UO_680 (O_680,N_29552,N_29321);
nor UO_681 (O_681,N_29493,N_29421);
nor UO_682 (O_682,N_29401,N_29213);
nand UO_683 (O_683,N_29751,N_29510);
xnor UO_684 (O_684,N_29817,N_29804);
or UO_685 (O_685,N_29490,N_29451);
or UO_686 (O_686,N_29235,N_29417);
and UO_687 (O_687,N_29591,N_29281);
nor UO_688 (O_688,N_29274,N_29948);
nor UO_689 (O_689,N_29818,N_29564);
or UO_690 (O_690,N_29712,N_29631);
xor UO_691 (O_691,N_29965,N_29365);
and UO_692 (O_692,N_29376,N_29335);
or UO_693 (O_693,N_29496,N_29434);
xnor UO_694 (O_694,N_29494,N_29023);
nor UO_695 (O_695,N_29140,N_29600);
nor UO_696 (O_696,N_29209,N_29727);
or UO_697 (O_697,N_29071,N_29655);
xnor UO_698 (O_698,N_29482,N_29128);
nand UO_699 (O_699,N_29507,N_29207);
or UO_700 (O_700,N_29775,N_29928);
and UO_701 (O_701,N_29928,N_29101);
or UO_702 (O_702,N_29553,N_29410);
and UO_703 (O_703,N_29838,N_29379);
xnor UO_704 (O_704,N_29971,N_29064);
or UO_705 (O_705,N_29734,N_29967);
xor UO_706 (O_706,N_29257,N_29156);
xnor UO_707 (O_707,N_29419,N_29644);
nor UO_708 (O_708,N_29448,N_29261);
or UO_709 (O_709,N_29951,N_29893);
nand UO_710 (O_710,N_29669,N_29736);
xor UO_711 (O_711,N_29178,N_29033);
nand UO_712 (O_712,N_29603,N_29556);
xnor UO_713 (O_713,N_29913,N_29449);
nor UO_714 (O_714,N_29845,N_29422);
nor UO_715 (O_715,N_29192,N_29608);
xnor UO_716 (O_716,N_29317,N_29609);
and UO_717 (O_717,N_29971,N_29065);
and UO_718 (O_718,N_29746,N_29429);
xor UO_719 (O_719,N_29389,N_29602);
and UO_720 (O_720,N_29823,N_29305);
xor UO_721 (O_721,N_29995,N_29314);
and UO_722 (O_722,N_29274,N_29693);
or UO_723 (O_723,N_29697,N_29488);
or UO_724 (O_724,N_29272,N_29397);
or UO_725 (O_725,N_29008,N_29326);
nand UO_726 (O_726,N_29066,N_29415);
xor UO_727 (O_727,N_29443,N_29531);
nor UO_728 (O_728,N_29613,N_29126);
nand UO_729 (O_729,N_29302,N_29021);
xnor UO_730 (O_730,N_29944,N_29799);
and UO_731 (O_731,N_29111,N_29813);
and UO_732 (O_732,N_29462,N_29921);
or UO_733 (O_733,N_29860,N_29455);
nand UO_734 (O_734,N_29738,N_29152);
and UO_735 (O_735,N_29443,N_29851);
or UO_736 (O_736,N_29126,N_29887);
nor UO_737 (O_737,N_29013,N_29717);
nand UO_738 (O_738,N_29770,N_29872);
or UO_739 (O_739,N_29408,N_29896);
xnor UO_740 (O_740,N_29796,N_29918);
or UO_741 (O_741,N_29335,N_29452);
nand UO_742 (O_742,N_29263,N_29503);
xnor UO_743 (O_743,N_29659,N_29156);
nand UO_744 (O_744,N_29466,N_29369);
nand UO_745 (O_745,N_29473,N_29392);
nor UO_746 (O_746,N_29917,N_29510);
nor UO_747 (O_747,N_29643,N_29773);
or UO_748 (O_748,N_29467,N_29618);
nand UO_749 (O_749,N_29599,N_29911);
nand UO_750 (O_750,N_29676,N_29634);
nand UO_751 (O_751,N_29628,N_29759);
or UO_752 (O_752,N_29896,N_29915);
or UO_753 (O_753,N_29280,N_29054);
xor UO_754 (O_754,N_29580,N_29492);
xor UO_755 (O_755,N_29727,N_29719);
nand UO_756 (O_756,N_29266,N_29610);
nand UO_757 (O_757,N_29211,N_29610);
or UO_758 (O_758,N_29751,N_29931);
and UO_759 (O_759,N_29211,N_29261);
nor UO_760 (O_760,N_29698,N_29429);
and UO_761 (O_761,N_29979,N_29110);
or UO_762 (O_762,N_29399,N_29486);
or UO_763 (O_763,N_29047,N_29698);
nor UO_764 (O_764,N_29874,N_29895);
or UO_765 (O_765,N_29452,N_29627);
or UO_766 (O_766,N_29195,N_29541);
nand UO_767 (O_767,N_29823,N_29179);
or UO_768 (O_768,N_29851,N_29714);
or UO_769 (O_769,N_29380,N_29647);
nor UO_770 (O_770,N_29530,N_29997);
or UO_771 (O_771,N_29032,N_29922);
and UO_772 (O_772,N_29870,N_29375);
nor UO_773 (O_773,N_29691,N_29102);
and UO_774 (O_774,N_29343,N_29389);
nand UO_775 (O_775,N_29449,N_29097);
or UO_776 (O_776,N_29202,N_29085);
and UO_777 (O_777,N_29658,N_29821);
and UO_778 (O_778,N_29014,N_29562);
nand UO_779 (O_779,N_29866,N_29328);
nor UO_780 (O_780,N_29384,N_29236);
xor UO_781 (O_781,N_29890,N_29943);
nand UO_782 (O_782,N_29439,N_29135);
or UO_783 (O_783,N_29301,N_29693);
and UO_784 (O_784,N_29042,N_29166);
and UO_785 (O_785,N_29915,N_29232);
or UO_786 (O_786,N_29968,N_29969);
xnor UO_787 (O_787,N_29280,N_29269);
nor UO_788 (O_788,N_29679,N_29690);
and UO_789 (O_789,N_29536,N_29152);
nand UO_790 (O_790,N_29020,N_29110);
nor UO_791 (O_791,N_29742,N_29869);
xor UO_792 (O_792,N_29245,N_29395);
xor UO_793 (O_793,N_29954,N_29707);
nand UO_794 (O_794,N_29804,N_29837);
and UO_795 (O_795,N_29622,N_29068);
and UO_796 (O_796,N_29385,N_29214);
xnor UO_797 (O_797,N_29559,N_29145);
nor UO_798 (O_798,N_29199,N_29264);
or UO_799 (O_799,N_29774,N_29732);
or UO_800 (O_800,N_29737,N_29206);
xnor UO_801 (O_801,N_29228,N_29611);
and UO_802 (O_802,N_29004,N_29892);
xnor UO_803 (O_803,N_29117,N_29649);
and UO_804 (O_804,N_29571,N_29220);
nor UO_805 (O_805,N_29551,N_29270);
or UO_806 (O_806,N_29747,N_29347);
or UO_807 (O_807,N_29832,N_29909);
nand UO_808 (O_808,N_29924,N_29127);
or UO_809 (O_809,N_29393,N_29564);
nand UO_810 (O_810,N_29138,N_29687);
nor UO_811 (O_811,N_29609,N_29124);
nor UO_812 (O_812,N_29540,N_29495);
nand UO_813 (O_813,N_29489,N_29857);
nor UO_814 (O_814,N_29645,N_29718);
or UO_815 (O_815,N_29422,N_29072);
and UO_816 (O_816,N_29396,N_29648);
xor UO_817 (O_817,N_29169,N_29454);
nand UO_818 (O_818,N_29553,N_29104);
nand UO_819 (O_819,N_29327,N_29131);
nand UO_820 (O_820,N_29265,N_29394);
or UO_821 (O_821,N_29547,N_29947);
or UO_822 (O_822,N_29177,N_29366);
nor UO_823 (O_823,N_29198,N_29799);
or UO_824 (O_824,N_29210,N_29198);
and UO_825 (O_825,N_29139,N_29133);
nor UO_826 (O_826,N_29071,N_29838);
or UO_827 (O_827,N_29200,N_29330);
nor UO_828 (O_828,N_29806,N_29819);
nor UO_829 (O_829,N_29179,N_29927);
or UO_830 (O_830,N_29783,N_29604);
xnor UO_831 (O_831,N_29069,N_29456);
nor UO_832 (O_832,N_29691,N_29088);
or UO_833 (O_833,N_29958,N_29097);
xor UO_834 (O_834,N_29875,N_29947);
or UO_835 (O_835,N_29060,N_29305);
or UO_836 (O_836,N_29573,N_29640);
nor UO_837 (O_837,N_29736,N_29188);
xnor UO_838 (O_838,N_29683,N_29068);
nor UO_839 (O_839,N_29560,N_29194);
and UO_840 (O_840,N_29305,N_29692);
nand UO_841 (O_841,N_29177,N_29943);
nand UO_842 (O_842,N_29303,N_29515);
xnor UO_843 (O_843,N_29680,N_29114);
xor UO_844 (O_844,N_29872,N_29165);
nand UO_845 (O_845,N_29219,N_29265);
and UO_846 (O_846,N_29940,N_29457);
nand UO_847 (O_847,N_29903,N_29482);
nor UO_848 (O_848,N_29229,N_29059);
or UO_849 (O_849,N_29829,N_29936);
or UO_850 (O_850,N_29699,N_29547);
xnor UO_851 (O_851,N_29023,N_29026);
nand UO_852 (O_852,N_29798,N_29925);
xor UO_853 (O_853,N_29249,N_29127);
xnor UO_854 (O_854,N_29235,N_29900);
nand UO_855 (O_855,N_29236,N_29481);
nand UO_856 (O_856,N_29076,N_29662);
and UO_857 (O_857,N_29013,N_29196);
nor UO_858 (O_858,N_29796,N_29416);
nand UO_859 (O_859,N_29855,N_29337);
nand UO_860 (O_860,N_29450,N_29553);
nand UO_861 (O_861,N_29768,N_29439);
xnor UO_862 (O_862,N_29620,N_29777);
nand UO_863 (O_863,N_29212,N_29316);
or UO_864 (O_864,N_29811,N_29824);
nor UO_865 (O_865,N_29528,N_29359);
nand UO_866 (O_866,N_29448,N_29548);
and UO_867 (O_867,N_29659,N_29635);
or UO_868 (O_868,N_29804,N_29526);
and UO_869 (O_869,N_29026,N_29115);
xnor UO_870 (O_870,N_29716,N_29967);
nand UO_871 (O_871,N_29312,N_29042);
xnor UO_872 (O_872,N_29857,N_29065);
or UO_873 (O_873,N_29258,N_29243);
xnor UO_874 (O_874,N_29328,N_29789);
nor UO_875 (O_875,N_29478,N_29025);
or UO_876 (O_876,N_29490,N_29831);
nor UO_877 (O_877,N_29994,N_29777);
nand UO_878 (O_878,N_29216,N_29594);
and UO_879 (O_879,N_29919,N_29870);
xnor UO_880 (O_880,N_29299,N_29930);
xor UO_881 (O_881,N_29033,N_29938);
or UO_882 (O_882,N_29972,N_29769);
nand UO_883 (O_883,N_29827,N_29152);
xor UO_884 (O_884,N_29541,N_29275);
nor UO_885 (O_885,N_29314,N_29979);
nand UO_886 (O_886,N_29094,N_29039);
nor UO_887 (O_887,N_29325,N_29630);
nor UO_888 (O_888,N_29075,N_29987);
nor UO_889 (O_889,N_29702,N_29054);
nor UO_890 (O_890,N_29032,N_29682);
nor UO_891 (O_891,N_29886,N_29706);
xor UO_892 (O_892,N_29937,N_29058);
nand UO_893 (O_893,N_29885,N_29924);
nor UO_894 (O_894,N_29728,N_29304);
and UO_895 (O_895,N_29603,N_29386);
nand UO_896 (O_896,N_29246,N_29510);
and UO_897 (O_897,N_29853,N_29249);
or UO_898 (O_898,N_29496,N_29707);
xor UO_899 (O_899,N_29697,N_29386);
or UO_900 (O_900,N_29796,N_29177);
or UO_901 (O_901,N_29627,N_29844);
and UO_902 (O_902,N_29404,N_29296);
xnor UO_903 (O_903,N_29389,N_29908);
and UO_904 (O_904,N_29624,N_29564);
nor UO_905 (O_905,N_29756,N_29785);
nand UO_906 (O_906,N_29803,N_29659);
nor UO_907 (O_907,N_29459,N_29381);
or UO_908 (O_908,N_29609,N_29497);
nor UO_909 (O_909,N_29062,N_29860);
xnor UO_910 (O_910,N_29960,N_29143);
nor UO_911 (O_911,N_29922,N_29892);
and UO_912 (O_912,N_29009,N_29290);
nor UO_913 (O_913,N_29066,N_29812);
xnor UO_914 (O_914,N_29440,N_29611);
and UO_915 (O_915,N_29650,N_29827);
xnor UO_916 (O_916,N_29558,N_29592);
and UO_917 (O_917,N_29639,N_29302);
nor UO_918 (O_918,N_29526,N_29834);
nor UO_919 (O_919,N_29128,N_29607);
and UO_920 (O_920,N_29140,N_29113);
or UO_921 (O_921,N_29544,N_29359);
nand UO_922 (O_922,N_29173,N_29547);
xnor UO_923 (O_923,N_29869,N_29820);
xnor UO_924 (O_924,N_29496,N_29508);
xnor UO_925 (O_925,N_29329,N_29099);
xor UO_926 (O_926,N_29067,N_29628);
nand UO_927 (O_927,N_29806,N_29884);
nand UO_928 (O_928,N_29085,N_29809);
or UO_929 (O_929,N_29085,N_29214);
nor UO_930 (O_930,N_29240,N_29103);
xnor UO_931 (O_931,N_29048,N_29170);
nor UO_932 (O_932,N_29418,N_29864);
nand UO_933 (O_933,N_29593,N_29342);
nor UO_934 (O_934,N_29550,N_29635);
xor UO_935 (O_935,N_29408,N_29087);
and UO_936 (O_936,N_29010,N_29307);
or UO_937 (O_937,N_29815,N_29238);
nor UO_938 (O_938,N_29594,N_29774);
xnor UO_939 (O_939,N_29266,N_29090);
nor UO_940 (O_940,N_29602,N_29474);
or UO_941 (O_941,N_29366,N_29661);
and UO_942 (O_942,N_29483,N_29469);
xor UO_943 (O_943,N_29483,N_29991);
nand UO_944 (O_944,N_29070,N_29952);
nand UO_945 (O_945,N_29376,N_29842);
and UO_946 (O_946,N_29727,N_29312);
or UO_947 (O_947,N_29119,N_29140);
nand UO_948 (O_948,N_29824,N_29757);
and UO_949 (O_949,N_29451,N_29955);
nor UO_950 (O_950,N_29458,N_29231);
nand UO_951 (O_951,N_29512,N_29583);
nand UO_952 (O_952,N_29883,N_29308);
nand UO_953 (O_953,N_29135,N_29042);
xnor UO_954 (O_954,N_29576,N_29249);
nand UO_955 (O_955,N_29612,N_29588);
and UO_956 (O_956,N_29632,N_29125);
and UO_957 (O_957,N_29265,N_29576);
nor UO_958 (O_958,N_29096,N_29656);
xor UO_959 (O_959,N_29474,N_29303);
xnor UO_960 (O_960,N_29087,N_29244);
or UO_961 (O_961,N_29630,N_29831);
and UO_962 (O_962,N_29973,N_29877);
xor UO_963 (O_963,N_29515,N_29098);
and UO_964 (O_964,N_29701,N_29047);
nor UO_965 (O_965,N_29518,N_29508);
nor UO_966 (O_966,N_29574,N_29484);
xnor UO_967 (O_967,N_29149,N_29167);
nand UO_968 (O_968,N_29632,N_29019);
and UO_969 (O_969,N_29240,N_29983);
and UO_970 (O_970,N_29293,N_29360);
or UO_971 (O_971,N_29117,N_29360);
xor UO_972 (O_972,N_29390,N_29159);
nand UO_973 (O_973,N_29393,N_29745);
or UO_974 (O_974,N_29927,N_29895);
xnor UO_975 (O_975,N_29701,N_29330);
or UO_976 (O_976,N_29070,N_29244);
xnor UO_977 (O_977,N_29454,N_29374);
xnor UO_978 (O_978,N_29662,N_29834);
or UO_979 (O_979,N_29617,N_29224);
nor UO_980 (O_980,N_29001,N_29327);
and UO_981 (O_981,N_29486,N_29799);
or UO_982 (O_982,N_29622,N_29364);
or UO_983 (O_983,N_29499,N_29750);
and UO_984 (O_984,N_29878,N_29949);
nor UO_985 (O_985,N_29209,N_29013);
nor UO_986 (O_986,N_29312,N_29792);
or UO_987 (O_987,N_29144,N_29899);
or UO_988 (O_988,N_29212,N_29743);
nor UO_989 (O_989,N_29630,N_29447);
or UO_990 (O_990,N_29672,N_29501);
nor UO_991 (O_991,N_29951,N_29749);
xnor UO_992 (O_992,N_29020,N_29588);
nand UO_993 (O_993,N_29363,N_29129);
and UO_994 (O_994,N_29286,N_29219);
xor UO_995 (O_995,N_29665,N_29780);
nand UO_996 (O_996,N_29054,N_29841);
xor UO_997 (O_997,N_29914,N_29244);
or UO_998 (O_998,N_29532,N_29791);
or UO_999 (O_999,N_29274,N_29909);
and UO_1000 (O_1000,N_29952,N_29239);
or UO_1001 (O_1001,N_29077,N_29772);
and UO_1002 (O_1002,N_29499,N_29972);
nand UO_1003 (O_1003,N_29090,N_29695);
nand UO_1004 (O_1004,N_29816,N_29283);
nand UO_1005 (O_1005,N_29118,N_29653);
or UO_1006 (O_1006,N_29905,N_29125);
xnor UO_1007 (O_1007,N_29961,N_29052);
or UO_1008 (O_1008,N_29589,N_29218);
or UO_1009 (O_1009,N_29198,N_29577);
xnor UO_1010 (O_1010,N_29365,N_29103);
xnor UO_1011 (O_1011,N_29059,N_29586);
nand UO_1012 (O_1012,N_29593,N_29986);
nor UO_1013 (O_1013,N_29782,N_29726);
nand UO_1014 (O_1014,N_29623,N_29629);
xnor UO_1015 (O_1015,N_29828,N_29126);
nor UO_1016 (O_1016,N_29568,N_29368);
nand UO_1017 (O_1017,N_29368,N_29715);
or UO_1018 (O_1018,N_29373,N_29334);
nor UO_1019 (O_1019,N_29286,N_29444);
nand UO_1020 (O_1020,N_29157,N_29652);
and UO_1021 (O_1021,N_29997,N_29258);
xnor UO_1022 (O_1022,N_29553,N_29465);
and UO_1023 (O_1023,N_29439,N_29810);
nand UO_1024 (O_1024,N_29880,N_29113);
or UO_1025 (O_1025,N_29151,N_29978);
xnor UO_1026 (O_1026,N_29747,N_29237);
nor UO_1027 (O_1027,N_29450,N_29049);
nand UO_1028 (O_1028,N_29146,N_29998);
xor UO_1029 (O_1029,N_29422,N_29278);
or UO_1030 (O_1030,N_29579,N_29436);
nor UO_1031 (O_1031,N_29131,N_29203);
or UO_1032 (O_1032,N_29272,N_29977);
or UO_1033 (O_1033,N_29243,N_29776);
or UO_1034 (O_1034,N_29954,N_29321);
and UO_1035 (O_1035,N_29936,N_29078);
nor UO_1036 (O_1036,N_29472,N_29440);
or UO_1037 (O_1037,N_29232,N_29535);
nor UO_1038 (O_1038,N_29420,N_29529);
nand UO_1039 (O_1039,N_29701,N_29262);
and UO_1040 (O_1040,N_29736,N_29630);
nor UO_1041 (O_1041,N_29636,N_29110);
nor UO_1042 (O_1042,N_29362,N_29192);
nor UO_1043 (O_1043,N_29249,N_29758);
or UO_1044 (O_1044,N_29449,N_29858);
and UO_1045 (O_1045,N_29820,N_29774);
and UO_1046 (O_1046,N_29707,N_29974);
or UO_1047 (O_1047,N_29266,N_29821);
xor UO_1048 (O_1048,N_29951,N_29950);
nor UO_1049 (O_1049,N_29331,N_29612);
xor UO_1050 (O_1050,N_29058,N_29406);
xnor UO_1051 (O_1051,N_29451,N_29570);
nor UO_1052 (O_1052,N_29953,N_29931);
or UO_1053 (O_1053,N_29941,N_29942);
nand UO_1054 (O_1054,N_29919,N_29175);
nand UO_1055 (O_1055,N_29222,N_29082);
nor UO_1056 (O_1056,N_29630,N_29384);
nand UO_1057 (O_1057,N_29056,N_29937);
nor UO_1058 (O_1058,N_29598,N_29129);
and UO_1059 (O_1059,N_29849,N_29462);
nor UO_1060 (O_1060,N_29128,N_29775);
or UO_1061 (O_1061,N_29790,N_29050);
and UO_1062 (O_1062,N_29754,N_29420);
or UO_1063 (O_1063,N_29379,N_29186);
nand UO_1064 (O_1064,N_29361,N_29736);
nor UO_1065 (O_1065,N_29700,N_29611);
xnor UO_1066 (O_1066,N_29296,N_29195);
and UO_1067 (O_1067,N_29920,N_29041);
nor UO_1068 (O_1068,N_29030,N_29166);
xnor UO_1069 (O_1069,N_29816,N_29507);
xor UO_1070 (O_1070,N_29602,N_29700);
xor UO_1071 (O_1071,N_29994,N_29492);
xor UO_1072 (O_1072,N_29537,N_29621);
nor UO_1073 (O_1073,N_29775,N_29224);
or UO_1074 (O_1074,N_29678,N_29956);
nor UO_1075 (O_1075,N_29491,N_29102);
and UO_1076 (O_1076,N_29252,N_29041);
or UO_1077 (O_1077,N_29751,N_29825);
and UO_1078 (O_1078,N_29159,N_29086);
or UO_1079 (O_1079,N_29573,N_29278);
or UO_1080 (O_1080,N_29891,N_29083);
or UO_1081 (O_1081,N_29390,N_29789);
and UO_1082 (O_1082,N_29605,N_29398);
and UO_1083 (O_1083,N_29363,N_29463);
and UO_1084 (O_1084,N_29016,N_29948);
xnor UO_1085 (O_1085,N_29911,N_29828);
or UO_1086 (O_1086,N_29467,N_29430);
nand UO_1087 (O_1087,N_29841,N_29603);
xnor UO_1088 (O_1088,N_29505,N_29026);
xor UO_1089 (O_1089,N_29046,N_29939);
xor UO_1090 (O_1090,N_29758,N_29401);
xor UO_1091 (O_1091,N_29263,N_29348);
nor UO_1092 (O_1092,N_29277,N_29428);
and UO_1093 (O_1093,N_29720,N_29812);
and UO_1094 (O_1094,N_29349,N_29204);
or UO_1095 (O_1095,N_29695,N_29189);
nor UO_1096 (O_1096,N_29225,N_29066);
or UO_1097 (O_1097,N_29897,N_29548);
nor UO_1098 (O_1098,N_29354,N_29407);
or UO_1099 (O_1099,N_29068,N_29463);
xnor UO_1100 (O_1100,N_29375,N_29869);
and UO_1101 (O_1101,N_29239,N_29956);
or UO_1102 (O_1102,N_29954,N_29261);
nand UO_1103 (O_1103,N_29775,N_29057);
nor UO_1104 (O_1104,N_29516,N_29425);
and UO_1105 (O_1105,N_29568,N_29855);
or UO_1106 (O_1106,N_29989,N_29648);
nand UO_1107 (O_1107,N_29720,N_29123);
nand UO_1108 (O_1108,N_29287,N_29899);
and UO_1109 (O_1109,N_29518,N_29612);
nor UO_1110 (O_1110,N_29757,N_29788);
nand UO_1111 (O_1111,N_29113,N_29251);
nand UO_1112 (O_1112,N_29765,N_29333);
xnor UO_1113 (O_1113,N_29010,N_29713);
xor UO_1114 (O_1114,N_29771,N_29139);
nor UO_1115 (O_1115,N_29246,N_29317);
nor UO_1116 (O_1116,N_29718,N_29942);
and UO_1117 (O_1117,N_29602,N_29043);
nor UO_1118 (O_1118,N_29559,N_29634);
nor UO_1119 (O_1119,N_29773,N_29726);
nand UO_1120 (O_1120,N_29325,N_29754);
or UO_1121 (O_1121,N_29128,N_29933);
or UO_1122 (O_1122,N_29043,N_29629);
and UO_1123 (O_1123,N_29212,N_29409);
and UO_1124 (O_1124,N_29288,N_29379);
or UO_1125 (O_1125,N_29319,N_29918);
nand UO_1126 (O_1126,N_29857,N_29441);
nand UO_1127 (O_1127,N_29992,N_29957);
nand UO_1128 (O_1128,N_29362,N_29703);
or UO_1129 (O_1129,N_29707,N_29490);
and UO_1130 (O_1130,N_29350,N_29177);
nor UO_1131 (O_1131,N_29578,N_29314);
and UO_1132 (O_1132,N_29114,N_29531);
and UO_1133 (O_1133,N_29789,N_29297);
xor UO_1134 (O_1134,N_29527,N_29422);
xnor UO_1135 (O_1135,N_29953,N_29337);
xnor UO_1136 (O_1136,N_29649,N_29082);
or UO_1137 (O_1137,N_29257,N_29962);
nand UO_1138 (O_1138,N_29844,N_29127);
nand UO_1139 (O_1139,N_29607,N_29106);
and UO_1140 (O_1140,N_29725,N_29802);
or UO_1141 (O_1141,N_29444,N_29257);
nor UO_1142 (O_1142,N_29933,N_29988);
nand UO_1143 (O_1143,N_29165,N_29527);
nor UO_1144 (O_1144,N_29955,N_29718);
xor UO_1145 (O_1145,N_29827,N_29617);
xor UO_1146 (O_1146,N_29933,N_29685);
or UO_1147 (O_1147,N_29157,N_29432);
xnor UO_1148 (O_1148,N_29312,N_29297);
or UO_1149 (O_1149,N_29584,N_29466);
xor UO_1150 (O_1150,N_29913,N_29891);
xnor UO_1151 (O_1151,N_29596,N_29076);
nand UO_1152 (O_1152,N_29626,N_29538);
or UO_1153 (O_1153,N_29444,N_29203);
and UO_1154 (O_1154,N_29924,N_29423);
or UO_1155 (O_1155,N_29323,N_29600);
xor UO_1156 (O_1156,N_29766,N_29393);
nand UO_1157 (O_1157,N_29983,N_29277);
or UO_1158 (O_1158,N_29717,N_29758);
nand UO_1159 (O_1159,N_29429,N_29283);
nand UO_1160 (O_1160,N_29034,N_29550);
or UO_1161 (O_1161,N_29991,N_29760);
or UO_1162 (O_1162,N_29620,N_29809);
or UO_1163 (O_1163,N_29851,N_29625);
or UO_1164 (O_1164,N_29598,N_29126);
nor UO_1165 (O_1165,N_29777,N_29388);
and UO_1166 (O_1166,N_29588,N_29877);
nand UO_1167 (O_1167,N_29873,N_29242);
nand UO_1168 (O_1168,N_29754,N_29611);
xor UO_1169 (O_1169,N_29545,N_29568);
xnor UO_1170 (O_1170,N_29396,N_29212);
nand UO_1171 (O_1171,N_29186,N_29841);
xnor UO_1172 (O_1172,N_29694,N_29733);
xor UO_1173 (O_1173,N_29800,N_29808);
nor UO_1174 (O_1174,N_29414,N_29170);
or UO_1175 (O_1175,N_29049,N_29806);
xnor UO_1176 (O_1176,N_29959,N_29203);
nand UO_1177 (O_1177,N_29135,N_29356);
nand UO_1178 (O_1178,N_29126,N_29248);
nor UO_1179 (O_1179,N_29693,N_29905);
and UO_1180 (O_1180,N_29158,N_29773);
or UO_1181 (O_1181,N_29448,N_29909);
and UO_1182 (O_1182,N_29592,N_29774);
xor UO_1183 (O_1183,N_29273,N_29681);
xor UO_1184 (O_1184,N_29446,N_29485);
or UO_1185 (O_1185,N_29216,N_29693);
xnor UO_1186 (O_1186,N_29857,N_29817);
and UO_1187 (O_1187,N_29579,N_29524);
or UO_1188 (O_1188,N_29728,N_29766);
or UO_1189 (O_1189,N_29213,N_29612);
nand UO_1190 (O_1190,N_29340,N_29734);
or UO_1191 (O_1191,N_29332,N_29702);
xnor UO_1192 (O_1192,N_29104,N_29759);
and UO_1193 (O_1193,N_29970,N_29773);
and UO_1194 (O_1194,N_29717,N_29918);
or UO_1195 (O_1195,N_29728,N_29396);
and UO_1196 (O_1196,N_29570,N_29054);
or UO_1197 (O_1197,N_29918,N_29819);
or UO_1198 (O_1198,N_29669,N_29228);
nor UO_1199 (O_1199,N_29382,N_29084);
and UO_1200 (O_1200,N_29133,N_29188);
nand UO_1201 (O_1201,N_29031,N_29292);
nor UO_1202 (O_1202,N_29276,N_29245);
nor UO_1203 (O_1203,N_29626,N_29288);
and UO_1204 (O_1204,N_29817,N_29343);
nor UO_1205 (O_1205,N_29374,N_29674);
or UO_1206 (O_1206,N_29302,N_29709);
and UO_1207 (O_1207,N_29102,N_29583);
and UO_1208 (O_1208,N_29496,N_29428);
and UO_1209 (O_1209,N_29075,N_29825);
and UO_1210 (O_1210,N_29239,N_29334);
or UO_1211 (O_1211,N_29324,N_29901);
nor UO_1212 (O_1212,N_29631,N_29639);
and UO_1213 (O_1213,N_29680,N_29033);
or UO_1214 (O_1214,N_29577,N_29449);
nand UO_1215 (O_1215,N_29354,N_29479);
xor UO_1216 (O_1216,N_29461,N_29148);
and UO_1217 (O_1217,N_29056,N_29789);
nand UO_1218 (O_1218,N_29714,N_29854);
xnor UO_1219 (O_1219,N_29842,N_29999);
or UO_1220 (O_1220,N_29806,N_29001);
nand UO_1221 (O_1221,N_29740,N_29984);
or UO_1222 (O_1222,N_29423,N_29191);
or UO_1223 (O_1223,N_29748,N_29186);
nand UO_1224 (O_1224,N_29964,N_29124);
nor UO_1225 (O_1225,N_29981,N_29928);
or UO_1226 (O_1226,N_29054,N_29150);
and UO_1227 (O_1227,N_29774,N_29276);
and UO_1228 (O_1228,N_29083,N_29698);
nand UO_1229 (O_1229,N_29051,N_29706);
or UO_1230 (O_1230,N_29070,N_29519);
xor UO_1231 (O_1231,N_29354,N_29384);
nand UO_1232 (O_1232,N_29061,N_29670);
and UO_1233 (O_1233,N_29358,N_29940);
or UO_1234 (O_1234,N_29149,N_29684);
or UO_1235 (O_1235,N_29666,N_29568);
xor UO_1236 (O_1236,N_29058,N_29304);
nand UO_1237 (O_1237,N_29386,N_29208);
xnor UO_1238 (O_1238,N_29412,N_29100);
and UO_1239 (O_1239,N_29693,N_29595);
and UO_1240 (O_1240,N_29773,N_29217);
xnor UO_1241 (O_1241,N_29582,N_29623);
and UO_1242 (O_1242,N_29627,N_29116);
and UO_1243 (O_1243,N_29909,N_29802);
and UO_1244 (O_1244,N_29759,N_29314);
nor UO_1245 (O_1245,N_29354,N_29018);
and UO_1246 (O_1246,N_29161,N_29088);
or UO_1247 (O_1247,N_29119,N_29625);
nor UO_1248 (O_1248,N_29839,N_29794);
and UO_1249 (O_1249,N_29495,N_29324);
and UO_1250 (O_1250,N_29128,N_29265);
nand UO_1251 (O_1251,N_29758,N_29510);
or UO_1252 (O_1252,N_29765,N_29707);
xnor UO_1253 (O_1253,N_29978,N_29469);
nor UO_1254 (O_1254,N_29467,N_29402);
xnor UO_1255 (O_1255,N_29676,N_29651);
and UO_1256 (O_1256,N_29786,N_29694);
nand UO_1257 (O_1257,N_29600,N_29907);
nor UO_1258 (O_1258,N_29245,N_29278);
xnor UO_1259 (O_1259,N_29570,N_29062);
nor UO_1260 (O_1260,N_29126,N_29869);
or UO_1261 (O_1261,N_29574,N_29224);
nand UO_1262 (O_1262,N_29830,N_29100);
or UO_1263 (O_1263,N_29616,N_29231);
nor UO_1264 (O_1264,N_29854,N_29403);
xor UO_1265 (O_1265,N_29195,N_29558);
nor UO_1266 (O_1266,N_29242,N_29865);
or UO_1267 (O_1267,N_29740,N_29750);
xnor UO_1268 (O_1268,N_29557,N_29638);
nand UO_1269 (O_1269,N_29463,N_29102);
xor UO_1270 (O_1270,N_29909,N_29107);
nand UO_1271 (O_1271,N_29681,N_29064);
xor UO_1272 (O_1272,N_29051,N_29018);
nor UO_1273 (O_1273,N_29421,N_29928);
or UO_1274 (O_1274,N_29738,N_29300);
or UO_1275 (O_1275,N_29025,N_29482);
nor UO_1276 (O_1276,N_29629,N_29162);
xnor UO_1277 (O_1277,N_29428,N_29785);
or UO_1278 (O_1278,N_29615,N_29180);
xnor UO_1279 (O_1279,N_29355,N_29634);
nand UO_1280 (O_1280,N_29830,N_29712);
nand UO_1281 (O_1281,N_29018,N_29774);
and UO_1282 (O_1282,N_29690,N_29073);
or UO_1283 (O_1283,N_29623,N_29720);
and UO_1284 (O_1284,N_29954,N_29356);
xnor UO_1285 (O_1285,N_29463,N_29857);
nand UO_1286 (O_1286,N_29201,N_29027);
and UO_1287 (O_1287,N_29802,N_29453);
xnor UO_1288 (O_1288,N_29192,N_29799);
or UO_1289 (O_1289,N_29906,N_29444);
nor UO_1290 (O_1290,N_29045,N_29879);
and UO_1291 (O_1291,N_29205,N_29054);
nand UO_1292 (O_1292,N_29237,N_29185);
or UO_1293 (O_1293,N_29561,N_29093);
xnor UO_1294 (O_1294,N_29645,N_29506);
nand UO_1295 (O_1295,N_29668,N_29772);
nor UO_1296 (O_1296,N_29221,N_29983);
and UO_1297 (O_1297,N_29635,N_29223);
and UO_1298 (O_1298,N_29555,N_29447);
nor UO_1299 (O_1299,N_29940,N_29337);
nand UO_1300 (O_1300,N_29900,N_29985);
and UO_1301 (O_1301,N_29919,N_29110);
and UO_1302 (O_1302,N_29155,N_29638);
nand UO_1303 (O_1303,N_29233,N_29842);
nand UO_1304 (O_1304,N_29295,N_29176);
and UO_1305 (O_1305,N_29596,N_29297);
nor UO_1306 (O_1306,N_29231,N_29757);
nand UO_1307 (O_1307,N_29234,N_29722);
and UO_1308 (O_1308,N_29323,N_29496);
nor UO_1309 (O_1309,N_29852,N_29184);
nand UO_1310 (O_1310,N_29445,N_29203);
xor UO_1311 (O_1311,N_29242,N_29257);
nand UO_1312 (O_1312,N_29858,N_29392);
xor UO_1313 (O_1313,N_29169,N_29262);
or UO_1314 (O_1314,N_29501,N_29480);
nor UO_1315 (O_1315,N_29489,N_29922);
and UO_1316 (O_1316,N_29665,N_29022);
and UO_1317 (O_1317,N_29292,N_29397);
or UO_1318 (O_1318,N_29808,N_29892);
or UO_1319 (O_1319,N_29351,N_29584);
nand UO_1320 (O_1320,N_29266,N_29216);
nor UO_1321 (O_1321,N_29388,N_29118);
nand UO_1322 (O_1322,N_29496,N_29730);
xnor UO_1323 (O_1323,N_29347,N_29711);
nand UO_1324 (O_1324,N_29221,N_29808);
or UO_1325 (O_1325,N_29331,N_29592);
and UO_1326 (O_1326,N_29506,N_29728);
xnor UO_1327 (O_1327,N_29728,N_29773);
nor UO_1328 (O_1328,N_29799,N_29293);
and UO_1329 (O_1329,N_29548,N_29422);
nand UO_1330 (O_1330,N_29120,N_29373);
and UO_1331 (O_1331,N_29613,N_29485);
and UO_1332 (O_1332,N_29580,N_29784);
and UO_1333 (O_1333,N_29124,N_29244);
xor UO_1334 (O_1334,N_29892,N_29369);
or UO_1335 (O_1335,N_29616,N_29101);
and UO_1336 (O_1336,N_29486,N_29209);
or UO_1337 (O_1337,N_29805,N_29913);
xnor UO_1338 (O_1338,N_29384,N_29282);
nor UO_1339 (O_1339,N_29838,N_29900);
nor UO_1340 (O_1340,N_29878,N_29466);
or UO_1341 (O_1341,N_29273,N_29699);
nand UO_1342 (O_1342,N_29720,N_29986);
nand UO_1343 (O_1343,N_29074,N_29199);
or UO_1344 (O_1344,N_29322,N_29612);
nor UO_1345 (O_1345,N_29362,N_29509);
xnor UO_1346 (O_1346,N_29067,N_29463);
nand UO_1347 (O_1347,N_29129,N_29460);
xnor UO_1348 (O_1348,N_29940,N_29737);
nand UO_1349 (O_1349,N_29889,N_29555);
or UO_1350 (O_1350,N_29572,N_29321);
nand UO_1351 (O_1351,N_29106,N_29485);
and UO_1352 (O_1352,N_29487,N_29560);
nor UO_1353 (O_1353,N_29717,N_29350);
xor UO_1354 (O_1354,N_29129,N_29185);
nor UO_1355 (O_1355,N_29897,N_29137);
and UO_1356 (O_1356,N_29402,N_29633);
or UO_1357 (O_1357,N_29674,N_29804);
nor UO_1358 (O_1358,N_29594,N_29174);
nor UO_1359 (O_1359,N_29150,N_29380);
nor UO_1360 (O_1360,N_29414,N_29885);
or UO_1361 (O_1361,N_29907,N_29552);
nand UO_1362 (O_1362,N_29495,N_29319);
or UO_1363 (O_1363,N_29638,N_29992);
nand UO_1364 (O_1364,N_29256,N_29153);
nor UO_1365 (O_1365,N_29506,N_29289);
nor UO_1366 (O_1366,N_29146,N_29206);
xnor UO_1367 (O_1367,N_29088,N_29269);
xnor UO_1368 (O_1368,N_29974,N_29647);
nand UO_1369 (O_1369,N_29061,N_29609);
and UO_1370 (O_1370,N_29970,N_29866);
nand UO_1371 (O_1371,N_29094,N_29449);
nor UO_1372 (O_1372,N_29880,N_29598);
nor UO_1373 (O_1373,N_29601,N_29168);
or UO_1374 (O_1374,N_29389,N_29665);
xnor UO_1375 (O_1375,N_29361,N_29808);
nand UO_1376 (O_1376,N_29660,N_29704);
xor UO_1377 (O_1377,N_29854,N_29677);
nor UO_1378 (O_1378,N_29463,N_29876);
or UO_1379 (O_1379,N_29917,N_29749);
xnor UO_1380 (O_1380,N_29896,N_29120);
xnor UO_1381 (O_1381,N_29434,N_29606);
nand UO_1382 (O_1382,N_29716,N_29408);
nor UO_1383 (O_1383,N_29458,N_29269);
and UO_1384 (O_1384,N_29340,N_29975);
or UO_1385 (O_1385,N_29737,N_29002);
and UO_1386 (O_1386,N_29218,N_29005);
nor UO_1387 (O_1387,N_29686,N_29208);
xor UO_1388 (O_1388,N_29205,N_29659);
xor UO_1389 (O_1389,N_29531,N_29750);
nand UO_1390 (O_1390,N_29635,N_29883);
nand UO_1391 (O_1391,N_29162,N_29731);
and UO_1392 (O_1392,N_29522,N_29314);
xor UO_1393 (O_1393,N_29959,N_29374);
or UO_1394 (O_1394,N_29708,N_29382);
xor UO_1395 (O_1395,N_29133,N_29278);
nand UO_1396 (O_1396,N_29634,N_29373);
nand UO_1397 (O_1397,N_29651,N_29463);
nand UO_1398 (O_1398,N_29751,N_29228);
nor UO_1399 (O_1399,N_29206,N_29526);
nor UO_1400 (O_1400,N_29118,N_29009);
and UO_1401 (O_1401,N_29870,N_29061);
nand UO_1402 (O_1402,N_29627,N_29962);
xor UO_1403 (O_1403,N_29593,N_29935);
nand UO_1404 (O_1404,N_29351,N_29173);
or UO_1405 (O_1405,N_29178,N_29425);
xnor UO_1406 (O_1406,N_29352,N_29930);
nand UO_1407 (O_1407,N_29379,N_29880);
nand UO_1408 (O_1408,N_29783,N_29814);
nor UO_1409 (O_1409,N_29797,N_29722);
xor UO_1410 (O_1410,N_29028,N_29642);
and UO_1411 (O_1411,N_29064,N_29206);
nor UO_1412 (O_1412,N_29245,N_29151);
nor UO_1413 (O_1413,N_29637,N_29649);
or UO_1414 (O_1414,N_29369,N_29251);
and UO_1415 (O_1415,N_29184,N_29587);
or UO_1416 (O_1416,N_29789,N_29141);
nor UO_1417 (O_1417,N_29978,N_29630);
or UO_1418 (O_1418,N_29617,N_29159);
nand UO_1419 (O_1419,N_29171,N_29090);
xnor UO_1420 (O_1420,N_29796,N_29733);
and UO_1421 (O_1421,N_29106,N_29279);
nand UO_1422 (O_1422,N_29950,N_29947);
xnor UO_1423 (O_1423,N_29291,N_29275);
xnor UO_1424 (O_1424,N_29509,N_29422);
nor UO_1425 (O_1425,N_29375,N_29338);
nand UO_1426 (O_1426,N_29083,N_29067);
nor UO_1427 (O_1427,N_29234,N_29415);
or UO_1428 (O_1428,N_29105,N_29974);
and UO_1429 (O_1429,N_29050,N_29494);
xnor UO_1430 (O_1430,N_29737,N_29971);
or UO_1431 (O_1431,N_29521,N_29765);
nand UO_1432 (O_1432,N_29307,N_29886);
nand UO_1433 (O_1433,N_29069,N_29429);
xor UO_1434 (O_1434,N_29638,N_29815);
nor UO_1435 (O_1435,N_29784,N_29837);
or UO_1436 (O_1436,N_29123,N_29445);
or UO_1437 (O_1437,N_29198,N_29456);
and UO_1438 (O_1438,N_29440,N_29107);
nand UO_1439 (O_1439,N_29171,N_29008);
nand UO_1440 (O_1440,N_29052,N_29254);
and UO_1441 (O_1441,N_29573,N_29848);
and UO_1442 (O_1442,N_29011,N_29279);
xnor UO_1443 (O_1443,N_29678,N_29058);
xor UO_1444 (O_1444,N_29956,N_29849);
or UO_1445 (O_1445,N_29693,N_29837);
nor UO_1446 (O_1446,N_29079,N_29803);
nor UO_1447 (O_1447,N_29551,N_29155);
or UO_1448 (O_1448,N_29091,N_29426);
xnor UO_1449 (O_1449,N_29923,N_29564);
and UO_1450 (O_1450,N_29657,N_29500);
or UO_1451 (O_1451,N_29643,N_29219);
nand UO_1452 (O_1452,N_29553,N_29257);
nor UO_1453 (O_1453,N_29660,N_29493);
nand UO_1454 (O_1454,N_29417,N_29748);
xnor UO_1455 (O_1455,N_29185,N_29083);
and UO_1456 (O_1456,N_29248,N_29383);
and UO_1457 (O_1457,N_29966,N_29019);
nor UO_1458 (O_1458,N_29696,N_29195);
nor UO_1459 (O_1459,N_29823,N_29268);
and UO_1460 (O_1460,N_29777,N_29849);
or UO_1461 (O_1461,N_29266,N_29750);
xnor UO_1462 (O_1462,N_29642,N_29565);
xnor UO_1463 (O_1463,N_29527,N_29063);
nand UO_1464 (O_1464,N_29657,N_29517);
or UO_1465 (O_1465,N_29280,N_29614);
nor UO_1466 (O_1466,N_29791,N_29863);
and UO_1467 (O_1467,N_29164,N_29755);
nor UO_1468 (O_1468,N_29441,N_29492);
or UO_1469 (O_1469,N_29879,N_29150);
and UO_1470 (O_1470,N_29026,N_29223);
xor UO_1471 (O_1471,N_29097,N_29291);
nand UO_1472 (O_1472,N_29631,N_29783);
or UO_1473 (O_1473,N_29099,N_29354);
nor UO_1474 (O_1474,N_29184,N_29609);
xor UO_1475 (O_1475,N_29256,N_29487);
and UO_1476 (O_1476,N_29327,N_29054);
nor UO_1477 (O_1477,N_29552,N_29257);
or UO_1478 (O_1478,N_29048,N_29817);
nor UO_1479 (O_1479,N_29342,N_29527);
nor UO_1480 (O_1480,N_29214,N_29461);
and UO_1481 (O_1481,N_29016,N_29544);
and UO_1482 (O_1482,N_29842,N_29938);
or UO_1483 (O_1483,N_29652,N_29687);
nand UO_1484 (O_1484,N_29409,N_29485);
nand UO_1485 (O_1485,N_29726,N_29564);
nand UO_1486 (O_1486,N_29424,N_29550);
nor UO_1487 (O_1487,N_29975,N_29092);
xnor UO_1488 (O_1488,N_29540,N_29604);
nand UO_1489 (O_1489,N_29061,N_29397);
nand UO_1490 (O_1490,N_29795,N_29652);
and UO_1491 (O_1491,N_29607,N_29892);
or UO_1492 (O_1492,N_29105,N_29989);
or UO_1493 (O_1493,N_29865,N_29251);
nor UO_1494 (O_1494,N_29903,N_29972);
or UO_1495 (O_1495,N_29524,N_29831);
nor UO_1496 (O_1496,N_29730,N_29810);
and UO_1497 (O_1497,N_29875,N_29854);
xnor UO_1498 (O_1498,N_29566,N_29825);
and UO_1499 (O_1499,N_29929,N_29558);
nand UO_1500 (O_1500,N_29047,N_29890);
and UO_1501 (O_1501,N_29422,N_29194);
nand UO_1502 (O_1502,N_29527,N_29239);
xor UO_1503 (O_1503,N_29661,N_29223);
nand UO_1504 (O_1504,N_29532,N_29504);
and UO_1505 (O_1505,N_29374,N_29441);
or UO_1506 (O_1506,N_29668,N_29621);
and UO_1507 (O_1507,N_29971,N_29743);
nand UO_1508 (O_1508,N_29096,N_29721);
xnor UO_1509 (O_1509,N_29586,N_29832);
nor UO_1510 (O_1510,N_29017,N_29837);
or UO_1511 (O_1511,N_29652,N_29616);
xor UO_1512 (O_1512,N_29065,N_29591);
nand UO_1513 (O_1513,N_29343,N_29147);
or UO_1514 (O_1514,N_29326,N_29944);
and UO_1515 (O_1515,N_29923,N_29326);
nand UO_1516 (O_1516,N_29539,N_29750);
and UO_1517 (O_1517,N_29093,N_29451);
and UO_1518 (O_1518,N_29631,N_29159);
or UO_1519 (O_1519,N_29759,N_29203);
and UO_1520 (O_1520,N_29101,N_29795);
nor UO_1521 (O_1521,N_29896,N_29157);
and UO_1522 (O_1522,N_29846,N_29376);
or UO_1523 (O_1523,N_29657,N_29904);
nor UO_1524 (O_1524,N_29990,N_29241);
xor UO_1525 (O_1525,N_29581,N_29659);
or UO_1526 (O_1526,N_29316,N_29853);
and UO_1527 (O_1527,N_29798,N_29738);
nand UO_1528 (O_1528,N_29651,N_29889);
or UO_1529 (O_1529,N_29709,N_29463);
nand UO_1530 (O_1530,N_29998,N_29035);
and UO_1531 (O_1531,N_29518,N_29069);
xnor UO_1532 (O_1532,N_29624,N_29661);
xor UO_1533 (O_1533,N_29402,N_29471);
and UO_1534 (O_1534,N_29848,N_29774);
nor UO_1535 (O_1535,N_29472,N_29277);
nand UO_1536 (O_1536,N_29482,N_29800);
nand UO_1537 (O_1537,N_29777,N_29475);
nor UO_1538 (O_1538,N_29776,N_29455);
nor UO_1539 (O_1539,N_29139,N_29921);
and UO_1540 (O_1540,N_29760,N_29922);
nand UO_1541 (O_1541,N_29254,N_29221);
xnor UO_1542 (O_1542,N_29588,N_29595);
nor UO_1543 (O_1543,N_29482,N_29171);
and UO_1544 (O_1544,N_29415,N_29014);
nand UO_1545 (O_1545,N_29002,N_29109);
and UO_1546 (O_1546,N_29368,N_29192);
xnor UO_1547 (O_1547,N_29877,N_29916);
or UO_1548 (O_1548,N_29730,N_29606);
xor UO_1549 (O_1549,N_29825,N_29725);
and UO_1550 (O_1550,N_29030,N_29897);
xnor UO_1551 (O_1551,N_29266,N_29270);
nor UO_1552 (O_1552,N_29558,N_29635);
and UO_1553 (O_1553,N_29474,N_29605);
nor UO_1554 (O_1554,N_29708,N_29911);
nor UO_1555 (O_1555,N_29407,N_29695);
nor UO_1556 (O_1556,N_29420,N_29573);
nor UO_1557 (O_1557,N_29766,N_29962);
xnor UO_1558 (O_1558,N_29323,N_29024);
or UO_1559 (O_1559,N_29037,N_29470);
or UO_1560 (O_1560,N_29190,N_29328);
xor UO_1561 (O_1561,N_29333,N_29539);
or UO_1562 (O_1562,N_29352,N_29728);
and UO_1563 (O_1563,N_29258,N_29736);
nand UO_1564 (O_1564,N_29024,N_29321);
nand UO_1565 (O_1565,N_29372,N_29866);
or UO_1566 (O_1566,N_29742,N_29220);
nor UO_1567 (O_1567,N_29206,N_29723);
nor UO_1568 (O_1568,N_29081,N_29048);
or UO_1569 (O_1569,N_29423,N_29772);
and UO_1570 (O_1570,N_29096,N_29351);
xor UO_1571 (O_1571,N_29978,N_29682);
and UO_1572 (O_1572,N_29040,N_29818);
nor UO_1573 (O_1573,N_29787,N_29309);
nand UO_1574 (O_1574,N_29866,N_29986);
nand UO_1575 (O_1575,N_29868,N_29741);
and UO_1576 (O_1576,N_29995,N_29776);
xnor UO_1577 (O_1577,N_29205,N_29893);
nor UO_1578 (O_1578,N_29349,N_29611);
nand UO_1579 (O_1579,N_29931,N_29873);
or UO_1580 (O_1580,N_29168,N_29540);
nor UO_1581 (O_1581,N_29933,N_29216);
and UO_1582 (O_1582,N_29195,N_29881);
and UO_1583 (O_1583,N_29552,N_29828);
nor UO_1584 (O_1584,N_29976,N_29469);
or UO_1585 (O_1585,N_29773,N_29442);
nor UO_1586 (O_1586,N_29910,N_29505);
nand UO_1587 (O_1587,N_29916,N_29993);
xnor UO_1588 (O_1588,N_29254,N_29970);
nand UO_1589 (O_1589,N_29213,N_29309);
nor UO_1590 (O_1590,N_29438,N_29451);
xnor UO_1591 (O_1591,N_29564,N_29816);
and UO_1592 (O_1592,N_29851,N_29749);
nor UO_1593 (O_1593,N_29535,N_29974);
xnor UO_1594 (O_1594,N_29545,N_29103);
and UO_1595 (O_1595,N_29853,N_29389);
and UO_1596 (O_1596,N_29575,N_29482);
xor UO_1597 (O_1597,N_29728,N_29906);
or UO_1598 (O_1598,N_29932,N_29712);
nor UO_1599 (O_1599,N_29521,N_29839);
and UO_1600 (O_1600,N_29931,N_29295);
xor UO_1601 (O_1601,N_29437,N_29167);
or UO_1602 (O_1602,N_29112,N_29625);
nand UO_1603 (O_1603,N_29480,N_29658);
nor UO_1604 (O_1604,N_29801,N_29252);
or UO_1605 (O_1605,N_29423,N_29467);
and UO_1606 (O_1606,N_29339,N_29038);
nor UO_1607 (O_1607,N_29251,N_29087);
nor UO_1608 (O_1608,N_29746,N_29747);
or UO_1609 (O_1609,N_29685,N_29841);
xnor UO_1610 (O_1610,N_29318,N_29966);
xor UO_1611 (O_1611,N_29249,N_29753);
and UO_1612 (O_1612,N_29516,N_29589);
nand UO_1613 (O_1613,N_29686,N_29358);
and UO_1614 (O_1614,N_29766,N_29442);
and UO_1615 (O_1615,N_29067,N_29813);
and UO_1616 (O_1616,N_29100,N_29348);
nand UO_1617 (O_1617,N_29313,N_29682);
nor UO_1618 (O_1618,N_29812,N_29282);
nor UO_1619 (O_1619,N_29192,N_29136);
xnor UO_1620 (O_1620,N_29999,N_29181);
nand UO_1621 (O_1621,N_29416,N_29657);
or UO_1622 (O_1622,N_29176,N_29040);
nand UO_1623 (O_1623,N_29281,N_29754);
and UO_1624 (O_1624,N_29109,N_29093);
or UO_1625 (O_1625,N_29585,N_29115);
or UO_1626 (O_1626,N_29353,N_29165);
nor UO_1627 (O_1627,N_29799,N_29771);
nand UO_1628 (O_1628,N_29949,N_29560);
or UO_1629 (O_1629,N_29759,N_29949);
xnor UO_1630 (O_1630,N_29734,N_29401);
or UO_1631 (O_1631,N_29628,N_29119);
nand UO_1632 (O_1632,N_29563,N_29751);
nand UO_1633 (O_1633,N_29970,N_29761);
xnor UO_1634 (O_1634,N_29438,N_29520);
nand UO_1635 (O_1635,N_29959,N_29833);
nor UO_1636 (O_1636,N_29436,N_29463);
xnor UO_1637 (O_1637,N_29066,N_29811);
or UO_1638 (O_1638,N_29839,N_29883);
and UO_1639 (O_1639,N_29539,N_29940);
nand UO_1640 (O_1640,N_29459,N_29108);
nor UO_1641 (O_1641,N_29696,N_29424);
nor UO_1642 (O_1642,N_29588,N_29830);
or UO_1643 (O_1643,N_29775,N_29458);
or UO_1644 (O_1644,N_29974,N_29564);
nand UO_1645 (O_1645,N_29672,N_29527);
and UO_1646 (O_1646,N_29875,N_29284);
or UO_1647 (O_1647,N_29950,N_29182);
and UO_1648 (O_1648,N_29649,N_29469);
xnor UO_1649 (O_1649,N_29167,N_29732);
or UO_1650 (O_1650,N_29847,N_29613);
xor UO_1651 (O_1651,N_29487,N_29078);
nand UO_1652 (O_1652,N_29726,N_29235);
and UO_1653 (O_1653,N_29167,N_29970);
or UO_1654 (O_1654,N_29607,N_29788);
nor UO_1655 (O_1655,N_29275,N_29403);
nand UO_1656 (O_1656,N_29067,N_29966);
nand UO_1657 (O_1657,N_29738,N_29438);
xor UO_1658 (O_1658,N_29347,N_29653);
nor UO_1659 (O_1659,N_29762,N_29315);
nand UO_1660 (O_1660,N_29164,N_29757);
or UO_1661 (O_1661,N_29893,N_29547);
and UO_1662 (O_1662,N_29983,N_29996);
xor UO_1663 (O_1663,N_29948,N_29612);
nor UO_1664 (O_1664,N_29607,N_29418);
nand UO_1665 (O_1665,N_29803,N_29875);
xor UO_1666 (O_1666,N_29210,N_29669);
and UO_1667 (O_1667,N_29672,N_29480);
nor UO_1668 (O_1668,N_29238,N_29325);
nor UO_1669 (O_1669,N_29092,N_29883);
nand UO_1670 (O_1670,N_29187,N_29625);
and UO_1671 (O_1671,N_29687,N_29291);
nand UO_1672 (O_1672,N_29038,N_29411);
and UO_1673 (O_1673,N_29282,N_29145);
or UO_1674 (O_1674,N_29834,N_29586);
xor UO_1675 (O_1675,N_29432,N_29954);
and UO_1676 (O_1676,N_29915,N_29110);
or UO_1677 (O_1677,N_29973,N_29010);
nor UO_1678 (O_1678,N_29190,N_29544);
nor UO_1679 (O_1679,N_29718,N_29409);
xnor UO_1680 (O_1680,N_29770,N_29580);
nand UO_1681 (O_1681,N_29377,N_29380);
or UO_1682 (O_1682,N_29965,N_29483);
or UO_1683 (O_1683,N_29032,N_29265);
and UO_1684 (O_1684,N_29382,N_29805);
nand UO_1685 (O_1685,N_29562,N_29624);
and UO_1686 (O_1686,N_29750,N_29520);
nor UO_1687 (O_1687,N_29642,N_29090);
nand UO_1688 (O_1688,N_29109,N_29193);
nand UO_1689 (O_1689,N_29560,N_29514);
nand UO_1690 (O_1690,N_29500,N_29049);
or UO_1691 (O_1691,N_29465,N_29866);
nor UO_1692 (O_1692,N_29187,N_29273);
or UO_1693 (O_1693,N_29572,N_29125);
nand UO_1694 (O_1694,N_29213,N_29765);
xnor UO_1695 (O_1695,N_29387,N_29204);
nor UO_1696 (O_1696,N_29397,N_29849);
or UO_1697 (O_1697,N_29114,N_29855);
nand UO_1698 (O_1698,N_29211,N_29781);
and UO_1699 (O_1699,N_29988,N_29453);
nor UO_1700 (O_1700,N_29410,N_29375);
nor UO_1701 (O_1701,N_29518,N_29563);
nor UO_1702 (O_1702,N_29654,N_29414);
or UO_1703 (O_1703,N_29763,N_29667);
and UO_1704 (O_1704,N_29783,N_29405);
nor UO_1705 (O_1705,N_29906,N_29992);
xnor UO_1706 (O_1706,N_29244,N_29201);
xor UO_1707 (O_1707,N_29484,N_29732);
or UO_1708 (O_1708,N_29219,N_29987);
or UO_1709 (O_1709,N_29207,N_29620);
and UO_1710 (O_1710,N_29686,N_29602);
xnor UO_1711 (O_1711,N_29321,N_29970);
nand UO_1712 (O_1712,N_29507,N_29494);
nor UO_1713 (O_1713,N_29122,N_29211);
or UO_1714 (O_1714,N_29767,N_29268);
or UO_1715 (O_1715,N_29101,N_29465);
nor UO_1716 (O_1716,N_29608,N_29251);
and UO_1717 (O_1717,N_29504,N_29319);
nand UO_1718 (O_1718,N_29382,N_29671);
and UO_1719 (O_1719,N_29860,N_29961);
or UO_1720 (O_1720,N_29367,N_29884);
nand UO_1721 (O_1721,N_29912,N_29590);
or UO_1722 (O_1722,N_29365,N_29643);
xnor UO_1723 (O_1723,N_29901,N_29996);
nand UO_1724 (O_1724,N_29654,N_29727);
nand UO_1725 (O_1725,N_29755,N_29660);
and UO_1726 (O_1726,N_29358,N_29232);
xnor UO_1727 (O_1727,N_29345,N_29061);
xnor UO_1728 (O_1728,N_29200,N_29378);
and UO_1729 (O_1729,N_29160,N_29007);
or UO_1730 (O_1730,N_29330,N_29660);
or UO_1731 (O_1731,N_29137,N_29451);
and UO_1732 (O_1732,N_29191,N_29589);
nor UO_1733 (O_1733,N_29932,N_29827);
nand UO_1734 (O_1734,N_29364,N_29746);
xor UO_1735 (O_1735,N_29843,N_29006);
nand UO_1736 (O_1736,N_29139,N_29171);
or UO_1737 (O_1737,N_29455,N_29628);
nor UO_1738 (O_1738,N_29572,N_29718);
nand UO_1739 (O_1739,N_29843,N_29373);
nand UO_1740 (O_1740,N_29977,N_29481);
or UO_1741 (O_1741,N_29211,N_29254);
or UO_1742 (O_1742,N_29732,N_29727);
nor UO_1743 (O_1743,N_29655,N_29907);
or UO_1744 (O_1744,N_29159,N_29345);
nor UO_1745 (O_1745,N_29743,N_29879);
xnor UO_1746 (O_1746,N_29140,N_29172);
nand UO_1747 (O_1747,N_29133,N_29754);
xor UO_1748 (O_1748,N_29365,N_29331);
xor UO_1749 (O_1749,N_29674,N_29913);
xnor UO_1750 (O_1750,N_29326,N_29498);
nor UO_1751 (O_1751,N_29608,N_29770);
nor UO_1752 (O_1752,N_29609,N_29577);
nor UO_1753 (O_1753,N_29017,N_29141);
nand UO_1754 (O_1754,N_29659,N_29436);
nand UO_1755 (O_1755,N_29807,N_29324);
nand UO_1756 (O_1756,N_29989,N_29256);
and UO_1757 (O_1757,N_29532,N_29231);
nor UO_1758 (O_1758,N_29307,N_29343);
nor UO_1759 (O_1759,N_29123,N_29447);
and UO_1760 (O_1760,N_29788,N_29487);
nand UO_1761 (O_1761,N_29110,N_29042);
xor UO_1762 (O_1762,N_29088,N_29380);
or UO_1763 (O_1763,N_29883,N_29629);
and UO_1764 (O_1764,N_29287,N_29189);
nor UO_1765 (O_1765,N_29599,N_29043);
nand UO_1766 (O_1766,N_29157,N_29112);
nor UO_1767 (O_1767,N_29777,N_29793);
and UO_1768 (O_1768,N_29631,N_29581);
nand UO_1769 (O_1769,N_29782,N_29780);
xor UO_1770 (O_1770,N_29470,N_29440);
or UO_1771 (O_1771,N_29846,N_29176);
nand UO_1772 (O_1772,N_29051,N_29464);
or UO_1773 (O_1773,N_29952,N_29161);
xnor UO_1774 (O_1774,N_29307,N_29972);
and UO_1775 (O_1775,N_29943,N_29922);
nand UO_1776 (O_1776,N_29673,N_29363);
and UO_1777 (O_1777,N_29945,N_29911);
nand UO_1778 (O_1778,N_29218,N_29877);
xor UO_1779 (O_1779,N_29009,N_29845);
or UO_1780 (O_1780,N_29201,N_29898);
or UO_1781 (O_1781,N_29304,N_29451);
or UO_1782 (O_1782,N_29560,N_29391);
xor UO_1783 (O_1783,N_29825,N_29233);
and UO_1784 (O_1784,N_29295,N_29425);
or UO_1785 (O_1785,N_29651,N_29483);
and UO_1786 (O_1786,N_29310,N_29638);
xor UO_1787 (O_1787,N_29998,N_29880);
xor UO_1788 (O_1788,N_29386,N_29099);
nor UO_1789 (O_1789,N_29080,N_29883);
and UO_1790 (O_1790,N_29539,N_29104);
xnor UO_1791 (O_1791,N_29810,N_29543);
nand UO_1792 (O_1792,N_29608,N_29056);
nor UO_1793 (O_1793,N_29751,N_29823);
nand UO_1794 (O_1794,N_29766,N_29180);
xnor UO_1795 (O_1795,N_29549,N_29765);
and UO_1796 (O_1796,N_29604,N_29125);
nor UO_1797 (O_1797,N_29632,N_29554);
nand UO_1798 (O_1798,N_29134,N_29460);
nand UO_1799 (O_1799,N_29770,N_29791);
xor UO_1800 (O_1800,N_29993,N_29155);
and UO_1801 (O_1801,N_29072,N_29874);
and UO_1802 (O_1802,N_29458,N_29620);
nor UO_1803 (O_1803,N_29135,N_29874);
and UO_1804 (O_1804,N_29632,N_29154);
nor UO_1805 (O_1805,N_29263,N_29596);
xor UO_1806 (O_1806,N_29980,N_29377);
xnor UO_1807 (O_1807,N_29247,N_29147);
xor UO_1808 (O_1808,N_29521,N_29463);
nand UO_1809 (O_1809,N_29258,N_29750);
xor UO_1810 (O_1810,N_29551,N_29643);
nor UO_1811 (O_1811,N_29015,N_29519);
nand UO_1812 (O_1812,N_29660,N_29063);
and UO_1813 (O_1813,N_29150,N_29756);
nor UO_1814 (O_1814,N_29855,N_29011);
nor UO_1815 (O_1815,N_29920,N_29110);
nor UO_1816 (O_1816,N_29930,N_29134);
nor UO_1817 (O_1817,N_29145,N_29985);
or UO_1818 (O_1818,N_29244,N_29620);
nor UO_1819 (O_1819,N_29210,N_29407);
nand UO_1820 (O_1820,N_29212,N_29053);
nand UO_1821 (O_1821,N_29441,N_29434);
xnor UO_1822 (O_1822,N_29982,N_29967);
xnor UO_1823 (O_1823,N_29255,N_29622);
nand UO_1824 (O_1824,N_29403,N_29310);
or UO_1825 (O_1825,N_29990,N_29024);
or UO_1826 (O_1826,N_29921,N_29811);
nand UO_1827 (O_1827,N_29052,N_29498);
or UO_1828 (O_1828,N_29796,N_29596);
nand UO_1829 (O_1829,N_29216,N_29909);
nor UO_1830 (O_1830,N_29401,N_29672);
and UO_1831 (O_1831,N_29745,N_29296);
or UO_1832 (O_1832,N_29717,N_29371);
xnor UO_1833 (O_1833,N_29315,N_29463);
nor UO_1834 (O_1834,N_29559,N_29538);
and UO_1835 (O_1835,N_29134,N_29878);
nor UO_1836 (O_1836,N_29262,N_29632);
or UO_1837 (O_1837,N_29940,N_29104);
nor UO_1838 (O_1838,N_29210,N_29561);
or UO_1839 (O_1839,N_29324,N_29263);
nand UO_1840 (O_1840,N_29527,N_29770);
xor UO_1841 (O_1841,N_29224,N_29675);
xor UO_1842 (O_1842,N_29240,N_29206);
nor UO_1843 (O_1843,N_29209,N_29051);
and UO_1844 (O_1844,N_29842,N_29290);
xor UO_1845 (O_1845,N_29250,N_29662);
nand UO_1846 (O_1846,N_29242,N_29849);
and UO_1847 (O_1847,N_29422,N_29043);
nand UO_1848 (O_1848,N_29711,N_29950);
xor UO_1849 (O_1849,N_29756,N_29095);
nor UO_1850 (O_1850,N_29739,N_29903);
and UO_1851 (O_1851,N_29401,N_29053);
xnor UO_1852 (O_1852,N_29312,N_29373);
xor UO_1853 (O_1853,N_29278,N_29250);
or UO_1854 (O_1854,N_29511,N_29811);
xnor UO_1855 (O_1855,N_29989,N_29024);
or UO_1856 (O_1856,N_29497,N_29130);
xor UO_1857 (O_1857,N_29453,N_29877);
nand UO_1858 (O_1858,N_29504,N_29022);
or UO_1859 (O_1859,N_29845,N_29250);
nand UO_1860 (O_1860,N_29127,N_29610);
xor UO_1861 (O_1861,N_29095,N_29327);
xnor UO_1862 (O_1862,N_29704,N_29051);
nor UO_1863 (O_1863,N_29542,N_29377);
xnor UO_1864 (O_1864,N_29015,N_29652);
and UO_1865 (O_1865,N_29353,N_29631);
nor UO_1866 (O_1866,N_29398,N_29886);
or UO_1867 (O_1867,N_29552,N_29031);
or UO_1868 (O_1868,N_29593,N_29424);
nand UO_1869 (O_1869,N_29951,N_29550);
nand UO_1870 (O_1870,N_29867,N_29629);
and UO_1871 (O_1871,N_29671,N_29937);
xor UO_1872 (O_1872,N_29172,N_29363);
or UO_1873 (O_1873,N_29024,N_29396);
and UO_1874 (O_1874,N_29554,N_29133);
and UO_1875 (O_1875,N_29259,N_29998);
nand UO_1876 (O_1876,N_29625,N_29082);
nor UO_1877 (O_1877,N_29433,N_29630);
nand UO_1878 (O_1878,N_29792,N_29435);
nand UO_1879 (O_1879,N_29291,N_29889);
nor UO_1880 (O_1880,N_29472,N_29878);
and UO_1881 (O_1881,N_29685,N_29047);
or UO_1882 (O_1882,N_29245,N_29121);
xnor UO_1883 (O_1883,N_29552,N_29517);
or UO_1884 (O_1884,N_29038,N_29397);
xnor UO_1885 (O_1885,N_29741,N_29411);
and UO_1886 (O_1886,N_29002,N_29922);
nor UO_1887 (O_1887,N_29590,N_29980);
nor UO_1888 (O_1888,N_29006,N_29632);
or UO_1889 (O_1889,N_29172,N_29482);
or UO_1890 (O_1890,N_29997,N_29709);
nand UO_1891 (O_1891,N_29455,N_29947);
and UO_1892 (O_1892,N_29103,N_29873);
nor UO_1893 (O_1893,N_29532,N_29239);
or UO_1894 (O_1894,N_29455,N_29853);
nand UO_1895 (O_1895,N_29309,N_29433);
and UO_1896 (O_1896,N_29226,N_29195);
or UO_1897 (O_1897,N_29099,N_29169);
nor UO_1898 (O_1898,N_29158,N_29590);
nand UO_1899 (O_1899,N_29583,N_29110);
nor UO_1900 (O_1900,N_29680,N_29539);
nand UO_1901 (O_1901,N_29487,N_29043);
nand UO_1902 (O_1902,N_29942,N_29261);
nand UO_1903 (O_1903,N_29465,N_29153);
nor UO_1904 (O_1904,N_29105,N_29759);
nand UO_1905 (O_1905,N_29352,N_29250);
or UO_1906 (O_1906,N_29702,N_29368);
nand UO_1907 (O_1907,N_29078,N_29595);
nor UO_1908 (O_1908,N_29856,N_29558);
nor UO_1909 (O_1909,N_29352,N_29918);
and UO_1910 (O_1910,N_29988,N_29620);
xnor UO_1911 (O_1911,N_29743,N_29655);
xor UO_1912 (O_1912,N_29965,N_29294);
nor UO_1913 (O_1913,N_29828,N_29905);
xor UO_1914 (O_1914,N_29780,N_29838);
or UO_1915 (O_1915,N_29492,N_29086);
xnor UO_1916 (O_1916,N_29763,N_29605);
nand UO_1917 (O_1917,N_29904,N_29810);
xor UO_1918 (O_1918,N_29245,N_29640);
nor UO_1919 (O_1919,N_29532,N_29208);
xor UO_1920 (O_1920,N_29142,N_29652);
or UO_1921 (O_1921,N_29821,N_29070);
nand UO_1922 (O_1922,N_29136,N_29443);
xor UO_1923 (O_1923,N_29996,N_29786);
nor UO_1924 (O_1924,N_29499,N_29507);
or UO_1925 (O_1925,N_29790,N_29592);
or UO_1926 (O_1926,N_29389,N_29153);
nor UO_1927 (O_1927,N_29447,N_29928);
nor UO_1928 (O_1928,N_29361,N_29864);
nand UO_1929 (O_1929,N_29037,N_29469);
nand UO_1930 (O_1930,N_29877,N_29091);
nor UO_1931 (O_1931,N_29545,N_29211);
nor UO_1932 (O_1932,N_29844,N_29467);
nand UO_1933 (O_1933,N_29515,N_29481);
nand UO_1934 (O_1934,N_29145,N_29136);
or UO_1935 (O_1935,N_29885,N_29848);
nand UO_1936 (O_1936,N_29120,N_29335);
nand UO_1937 (O_1937,N_29439,N_29815);
nand UO_1938 (O_1938,N_29836,N_29524);
xor UO_1939 (O_1939,N_29080,N_29411);
nor UO_1940 (O_1940,N_29297,N_29333);
and UO_1941 (O_1941,N_29841,N_29593);
and UO_1942 (O_1942,N_29901,N_29119);
or UO_1943 (O_1943,N_29213,N_29193);
or UO_1944 (O_1944,N_29299,N_29268);
nor UO_1945 (O_1945,N_29060,N_29957);
xor UO_1946 (O_1946,N_29840,N_29346);
or UO_1947 (O_1947,N_29198,N_29288);
or UO_1948 (O_1948,N_29548,N_29828);
xnor UO_1949 (O_1949,N_29411,N_29034);
nand UO_1950 (O_1950,N_29682,N_29230);
nor UO_1951 (O_1951,N_29255,N_29441);
and UO_1952 (O_1952,N_29852,N_29083);
xor UO_1953 (O_1953,N_29199,N_29228);
xor UO_1954 (O_1954,N_29633,N_29582);
and UO_1955 (O_1955,N_29758,N_29146);
nand UO_1956 (O_1956,N_29914,N_29171);
xnor UO_1957 (O_1957,N_29753,N_29181);
xnor UO_1958 (O_1958,N_29141,N_29942);
nor UO_1959 (O_1959,N_29120,N_29359);
nor UO_1960 (O_1960,N_29231,N_29503);
nor UO_1961 (O_1961,N_29234,N_29401);
or UO_1962 (O_1962,N_29593,N_29050);
or UO_1963 (O_1963,N_29879,N_29534);
nor UO_1964 (O_1964,N_29063,N_29061);
nand UO_1965 (O_1965,N_29876,N_29759);
or UO_1966 (O_1966,N_29625,N_29285);
xor UO_1967 (O_1967,N_29941,N_29320);
nand UO_1968 (O_1968,N_29778,N_29562);
and UO_1969 (O_1969,N_29057,N_29933);
nor UO_1970 (O_1970,N_29661,N_29040);
or UO_1971 (O_1971,N_29195,N_29031);
nand UO_1972 (O_1972,N_29587,N_29888);
nand UO_1973 (O_1973,N_29164,N_29015);
xnor UO_1974 (O_1974,N_29793,N_29386);
nor UO_1975 (O_1975,N_29729,N_29899);
nand UO_1976 (O_1976,N_29098,N_29450);
nor UO_1977 (O_1977,N_29143,N_29712);
nor UO_1978 (O_1978,N_29670,N_29939);
nor UO_1979 (O_1979,N_29325,N_29820);
nor UO_1980 (O_1980,N_29168,N_29226);
and UO_1981 (O_1981,N_29419,N_29096);
xor UO_1982 (O_1982,N_29235,N_29719);
nor UO_1983 (O_1983,N_29377,N_29929);
nor UO_1984 (O_1984,N_29027,N_29858);
and UO_1985 (O_1985,N_29293,N_29594);
nand UO_1986 (O_1986,N_29248,N_29427);
nand UO_1987 (O_1987,N_29783,N_29055);
nand UO_1988 (O_1988,N_29735,N_29053);
nor UO_1989 (O_1989,N_29036,N_29772);
and UO_1990 (O_1990,N_29295,N_29716);
nand UO_1991 (O_1991,N_29566,N_29387);
nor UO_1992 (O_1992,N_29263,N_29285);
xnor UO_1993 (O_1993,N_29384,N_29531);
or UO_1994 (O_1994,N_29246,N_29910);
nand UO_1995 (O_1995,N_29443,N_29591);
nand UO_1996 (O_1996,N_29684,N_29453);
nor UO_1997 (O_1997,N_29480,N_29469);
nor UO_1998 (O_1998,N_29098,N_29130);
nand UO_1999 (O_1999,N_29276,N_29469);
xnor UO_2000 (O_2000,N_29987,N_29200);
nor UO_2001 (O_2001,N_29516,N_29752);
or UO_2002 (O_2002,N_29993,N_29261);
xor UO_2003 (O_2003,N_29897,N_29070);
and UO_2004 (O_2004,N_29842,N_29208);
nor UO_2005 (O_2005,N_29300,N_29028);
nand UO_2006 (O_2006,N_29271,N_29302);
nand UO_2007 (O_2007,N_29322,N_29007);
nor UO_2008 (O_2008,N_29588,N_29141);
and UO_2009 (O_2009,N_29855,N_29284);
nor UO_2010 (O_2010,N_29601,N_29903);
nand UO_2011 (O_2011,N_29653,N_29099);
nor UO_2012 (O_2012,N_29437,N_29422);
nor UO_2013 (O_2013,N_29655,N_29632);
xnor UO_2014 (O_2014,N_29784,N_29453);
nor UO_2015 (O_2015,N_29532,N_29672);
or UO_2016 (O_2016,N_29721,N_29495);
and UO_2017 (O_2017,N_29822,N_29075);
xor UO_2018 (O_2018,N_29882,N_29280);
and UO_2019 (O_2019,N_29235,N_29475);
xor UO_2020 (O_2020,N_29070,N_29881);
xor UO_2021 (O_2021,N_29288,N_29569);
nor UO_2022 (O_2022,N_29650,N_29008);
or UO_2023 (O_2023,N_29889,N_29280);
and UO_2024 (O_2024,N_29565,N_29026);
or UO_2025 (O_2025,N_29934,N_29296);
xnor UO_2026 (O_2026,N_29493,N_29112);
and UO_2027 (O_2027,N_29373,N_29694);
and UO_2028 (O_2028,N_29121,N_29993);
nor UO_2029 (O_2029,N_29887,N_29888);
xor UO_2030 (O_2030,N_29919,N_29965);
and UO_2031 (O_2031,N_29683,N_29067);
and UO_2032 (O_2032,N_29373,N_29960);
nor UO_2033 (O_2033,N_29499,N_29875);
nor UO_2034 (O_2034,N_29987,N_29595);
xor UO_2035 (O_2035,N_29010,N_29478);
or UO_2036 (O_2036,N_29649,N_29539);
or UO_2037 (O_2037,N_29791,N_29426);
nand UO_2038 (O_2038,N_29390,N_29707);
nor UO_2039 (O_2039,N_29958,N_29174);
nand UO_2040 (O_2040,N_29002,N_29129);
nor UO_2041 (O_2041,N_29789,N_29578);
and UO_2042 (O_2042,N_29762,N_29797);
nand UO_2043 (O_2043,N_29012,N_29711);
and UO_2044 (O_2044,N_29488,N_29473);
xor UO_2045 (O_2045,N_29173,N_29939);
xnor UO_2046 (O_2046,N_29978,N_29919);
xor UO_2047 (O_2047,N_29625,N_29799);
or UO_2048 (O_2048,N_29298,N_29437);
and UO_2049 (O_2049,N_29334,N_29644);
nand UO_2050 (O_2050,N_29485,N_29399);
or UO_2051 (O_2051,N_29086,N_29358);
nand UO_2052 (O_2052,N_29008,N_29933);
and UO_2053 (O_2053,N_29733,N_29174);
nor UO_2054 (O_2054,N_29981,N_29913);
and UO_2055 (O_2055,N_29776,N_29099);
or UO_2056 (O_2056,N_29235,N_29684);
and UO_2057 (O_2057,N_29165,N_29200);
nor UO_2058 (O_2058,N_29288,N_29835);
xor UO_2059 (O_2059,N_29606,N_29391);
nand UO_2060 (O_2060,N_29363,N_29958);
xnor UO_2061 (O_2061,N_29772,N_29636);
and UO_2062 (O_2062,N_29850,N_29611);
or UO_2063 (O_2063,N_29562,N_29537);
and UO_2064 (O_2064,N_29955,N_29128);
and UO_2065 (O_2065,N_29197,N_29490);
nor UO_2066 (O_2066,N_29353,N_29364);
and UO_2067 (O_2067,N_29611,N_29790);
nand UO_2068 (O_2068,N_29934,N_29575);
and UO_2069 (O_2069,N_29224,N_29159);
xor UO_2070 (O_2070,N_29885,N_29412);
and UO_2071 (O_2071,N_29974,N_29522);
and UO_2072 (O_2072,N_29794,N_29295);
nor UO_2073 (O_2073,N_29849,N_29268);
nand UO_2074 (O_2074,N_29725,N_29192);
nor UO_2075 (O_2075,N_29551,N_29750);
and UO_2076 (O_2076,N_29953,N_29127);
xnor UO_2077 (O_2077,N_29763,N_29728);
xnor UO_2078 (O_2078,N_29442,N_29213);
nand UO_2079 (O_2079,N_29604,N_29119);
and UO_2080 (O_2080,N_29767,N_29447);
or UO_2081 (O_2081,N_29078,N_29449);
or UO_2082 (O_2082,N_29807,N_29339);
xnor UO_2083 (O_2083,N_29031,N_29441);
and UO_2084 (O_2084,N_29208,N_29295);
nor UO_2085 (O_2085,N_29267,N_29222);
nand UO_2086 (O_2086,N_29284,N_29709);
xor UO_2087 (O_2087,N_29364,N_29577);
or UO_2088 (O_2088,N_29286,N_29379);
nand UO_2089 (O_2089,N_29156,N_29912);
xnor UO_2090 (O_2090,N_29552,N_29869);
or UO_2091 (O_2091,N_29650,N_29062);
and UO_2092 (O_2092,N_29199,N_29189);
nand UO_2093 (O_2093,N_29763,N_29212);
or UO_2094 (O_2094,N_29617,N_29702);
or UO_2095 (O_2095,N_29133,N_29623);
xnor UO_2096 (O_2096,N_29205,N_29915);
xor UO_2097 (O_2097,N_29784,N_29642);
xnor UO_2098 (O_2098,N_29969,N_29165);
nand UO_2099 (O_2099,N_29549,N_29238);
nand UO_2100 (O_2100,N_29203,N_29313);
or UO_2101 (O_2101,N_29354,N_29609);
xnor UO_2102 (O_2102,N_29422,N_29818);
and UO_2103 (O_2103,N_29513,N_29378);
and UO_2104 (O_2104,N_29258,N_29096);
nor UO_2105 (O_2105,N_29505,N_29804);
nor UO_2106 (O_2106,N_29740,N_29917);
nand UO_2107 (O_2107,N_29342,N_29208);
xnor UO_2108 (O_2108,N_29995,N_29528);
and UO_2109 (O_2109,N_29109,N_29699);
and UO_2110 (O_2110,N_29453,N_29754);
or UO_2111 (O_2111,N_29419,N_29143);
and UO_2112 (O_2112,N_29705,N_29374);
xor UO_2113 (O_2113,N_29856,N_29058);
or UO_2114 (O_2114,N_29173,N_29896);
or UO_2115 (O_2115,N_29689,N_29924);
xnor UO_2116 (O_2116,N_29005,N_29581);
xnor UO_2117 (O_2117,N_29492,N_29529);
and UO_2118 (O_2118,N_29658,N_29778);
or UO_2119 (O_2119,N_29407,N_29514);
and UO_2120 (O_2120,N_29538,N_29211);
nand UO_2121 (O_2121,N_29790,N_29055);
or UO_2122 (O_2122,N_29712,N_29418);
nor UO_2123 (O_2123,N_29691,N_29576);
xnor UO_2124 (O_2124,N_29623,N_29066);
nor UO_2125 (O_2125,N_29511,N_29673);
nor UO_2126 (O_2126,N_29885,N_29300);
nor UO_2127 (O_2127,N_29151,N_29526);
and UO_2128 (O_2128,N_29915,N_29464);
nor UO_2129 (O_2129,N_29156,N_29290);
nand UO_2130 (O_2130,N_29440,N_29328);
or UO_2131 (O_2131,N_29020,N_29858);
nand UO_2132 (O_2132,N_29711,N_29226);
nand UO_2133 (O_2133,N_29485,N_29776);
nor UO_2134 (O_2134,N_29603,N_29041);
and UO_2135 (O_2135,N_29116,N_29099);
or UO_2136 (O_2136,N_29893,N_29827);
or UO_2137 (O_2137,N_29655,N_29107);
and UO_2138 (O_2138,N_29700,N_29928);
and UO_2139 (O_2139,N_29409,N_29680);
nand UO_2140 (O_2140,N_29957,N_29065);
nor UO_2141 (O_2141,N_29753,N_29875);
nor UO_2142 (O_2142,N_29401,N_29934);
and UO_2143 (O_2143,N_29833,N_29963);
or UO_2144 (O_2144,N_29303,N_29696);
nor UO_2145 (O_2145,N_29116,N_29083);
nand UO_2146 (O_2146,N_29463,N_29752);
nor UO_2147 (O_2147,N_29034,N_29519);
and UO_2148 (O_2148,N_29006,N_29185);
and UO_2149 (O_2149,N_29574,N_29345);
nor UO_2150 (O_2150,N_29383,N_29191);
nor UO_2151 (O_2151,N_29566,N_29816);
and UO_2152 (O_2152,N_29996,N_29331);
nor UO_2153 (O_2153,N_29421,N_29810);
nand UO_2154 (O_2154,N_29357,N_29959);
nand UO_2155 (O_2155,N_29591,N_29310);
nand UO_2156 (O_2156,N_29080,N_29007);
or UO_2157 (O_2157,N_29675,N_29316);
xnor UO_2158 (O_2158,N_29641,N_29319);
xnor UO_2159 (O_2159,N_29989,N_29951);
or UO_2160 (O_2160,N_29568,N_29581);
or UO_2161 (O_2161,N_29545,N_29917);
xnor UO_2162 (O_2162,N_29015,N_29257);
and UO_2163 (O_2163,N_29708,N_29879);
nor UO_2164 (O_2164,N_29052,N_29244);
nand UO_2165 (O_2165,N_29101,N_29478);
xor UO_2166 (O_2166,N_29273,N_29560);
xor UO_2167 (O_2167,N_29522,N_29614);
and UO_2168 (O_2168,N_29863,N_29612);
and UO_2169 (O_2169,N_29092,N_29452);
and UO_2170 (O_2170,N_29115,N_29681);
or UO_2171 (O_2171,N_29898,N_29916);
xor UO_2172 (O_2172,N_29611,N_29244);
xnor UO_2173 (O_2173,N_29928,N_29980);
nor UO_2174 (O_2174,N_29276,N_29913);
xor UO_2175 (O_2175,N_29940,N_29788);
and UO_2176 (O_2176,N_29722,N_29621);
nor UO_2177 (O_2177,N_29406,N_29293);
or UO_2178 (O_2178,N_29708,N_29133);
xnor UO_2179 (O_2179,N_29353,N_29179);
and UO_2180 (O_2180,N_29653,N_29085);
nor UO_2181 (O_2181,N_29088,N_29542);
nand UO_2182 (O_2182,N_29958,N_29380);
or UO_2183 (O_2183,N_29136,N_29673);
nand UO_2184 (O_2184,N_29029,N_29642);
xor UO_2185 (O_2185,N_29844,N_29072);
and UO_2186 (O_2186,N_29219,N_29867);
or UO_2187 (O_2187,N_29051,N_29803);
nor UO_2188 (O_2188,N_29283,N_29957);
and UO_2189 (O_2189,N_29121,N_29258);
or UO_2190 (O_2190,N_29342,N_29566);
and UO_2191 (O_2191,N_29436,N_29740);
or UO_2192 (O_2192,N_29034,N_29315);
nor UO_2193 (O_2193,N_29522,N_29935);
and UO_2194 (O_2194,N_29283,N_29883);
nand UO_2195 (O_2195,N_29436,N_29332);
or UO_2196 (O_2196,N_29328,N_29314);
or UO_2197 (O_2197,N_29743,N_29570);
or UO_2198 (O_2198,N_29027,N_29387);
xnor UO_2199 (O_2199,N_29321,N_29525);
nand UO_2200 (O_2200,N_29040,N_29452);
nor UO_2201 (O_2201,N_29845,N_29523);
or UO_2202 (O_2202,N_29503,N_29245);
nand UO_2203 (O_2203,N_29597,N_29867);
or UO_2204 (O_2204,N_29332,N_29961);
xnor UO_2205 (O_2205,N_29277,N_29888);
and UO_2206 (O_2206,N_29052,N_29784);
xnor UO_2207 (O_2207,N_29042,N_29929);
and UO_2208 (O_2208,N_29195,N_29718);
nand UO_2209 (O_2209,N_29774,N_29910);
xnor UO_2210 (O_2210,N_29863,N_29644);
or UO_2211 (O_2211,N_29003,N_29963);
or UO_2212 (O_2212,N_29295,N_29702);
nor UO_2213 (O_2213,N_29710,N_29541);
xnor UO_2214 (O_2214,N_29973,N_29919);
nand UO_2215 (O_2215,N_29165,N_29990);
nand UO_2216 (O_2216,N_29356,N_29174);
nor UO_2217 (O_2217,N_29648,N_29887);
nand UO_2218 (O_2218,N_29004,N_29552);
or UO_2219 (O_2219,N_29703,N_29114);
xor UO_2220 (O_2220,N_29790,N_29782);
nor UO_2221 (O_2221,N_29635,N_29623);
xor UO_2222 (O_2222,N_29611,N_29856);
and UO_2223 (O_2223,N_29955,N_29772);
nor UO_2224 (O_2224,N_29542,N_29258);
xnor UO_2225 (O_2225,N_29658,N_29168);
nor UO_2226 (O_2226,N_29427,N_29136);
xor UO_2227 (O_2227,N_29148,N_29894);
and UO_2228 (O_2228,N_29061,N_29836);
and UO_2229 (O_2229,N_29525,N_29274);
xnor UO_2230 (O_2230,N_29851,N_29144);
or UO_2231 (O_2231,N_29000,N_29588);
and UO_2232 (O_2232,N_29427,N_29106);
or UO_2233 (O_2233,N_29404,N_29340);
nor UO_2234 (O_2234,N_29972,N_29951);
xor UO_2235 (O_2235,N_29889,N_29816);
nor UO_2236 (O_2236,N_29011,N_29471);
nor UO_2237 (O_2237,N_29581,N_29501);
nor UO_2238 (O_2238,N_29433,N_29981);
nor UO_2239 (O_2239,N_29016,N_29284);
nand UO_2240 (O_2240,N_29508,N_29627);
or UO_2241 (O_2241,N_29617,N_29454);
and UO_2242 (O_2242,N_29028,N_29714);
xor UO_2243 (O_2243,N_29328,N_29635);
xor UO_2244 (O_2244,N_29510,N_29067);
or UO_2245 (O_2245,N_29418,N_29759);
xnor UO_2246 (O_2246,N_29126,N_29650);
nor UO_2247 (O_2247,N_29976,N_29085);
nand UO_2248 (O_2248,N_29618,N_29079);
nand UO_2249 (O_2249,N_29533,N_29907);
nor UO_2250 (O_2250,N_29932,N_29145);
nor UO_2251 (O_2251,N_29111,N_29671);
and UO_2252 (O_2252,N_29652,N_29003);
xnor UO_2253 (O_2253,N_29272,N_29843);
xnor UO_2254 (O_2254,N_29177,N_29749);
and UO_2255 (O_2255,N_29481,N_29642);
nor UO_2256 (O_2256,N_29720,N_29876);
nor UO_2257 (O_2257,N_29929,N_29847);
xnor UO_2258 (O_2258,N_29210,N_29120);
and UO_2259 (O_2259,N_29656,N_29612);
or UO_2260 (O_2260,N_29008,N_29793);
and UO_2261 (O_2261,N_29668,N_29836);
or UO_2262 (O_2262,N_29560,N_29075);
and UO_2263 (O_2263,N_29896,N_29413);
xnor UO_2264 (O_2264,N_29124,N_29006);
nand UO_2265 (O_2265,N_29327,N_29323);
and UO_2266 (O_2266,N_29314,N_29030);
nand UO_2267 (O_2267,N_29067,N_29553);
xnor UO_2268 (O_2268,N_29352,N_29760);
and UO_2269 (O_2269,N_29528,N_29322);
and UO_2270 (O_2270,N_29625,N_29431);
nor UO_2271 (O_2271,N_29979,N_29669);
or UO_2272 (O_2272,N_29204,N_29301);
nor UO_2273 (O_2273,N_29287,N_29493);
xor UO_2274 (O_2274,N_29555,N_29924);
nand UO_2275 (O_2275,N_29195,N_29762);
xor UO_2276 (O_2276,N_29378,N_29801);
and UO_2277 (O_2277,N_29622,N_29754);
or UO_2278 (O_2278,N_29092,N_29447);
or UO_2279 (O_2279,N_29435,N_29829);
nand UO_2280 (O_2280,N_29994,N_29342);
or UO_2281 (O_2281,N_29589,N_29972);
nand UO_2282 (O_2282,N_29799,N_29475);
and UO_2283 (O_2283,N_29987,N_29407);
or UO_2284 (O_2284,N_29318,N_29079);
nor UO_2285 (O_2285,N_29313,N_29467);
xor UO_2286 (O_2286,N_29590,N_29695);
and UO_2287 (O_2287,N_29016,N_29686);
and UO_2288 (O_2288,N_29526,N_29108);
or UO_2289 (O_2289,N_29767,N_29498);
nor UO_2290 (O_2290,N_29949,N_29657);
xor UO_2291 (O_2291,N_29668,N_29486);
nand UO_2292 (O_2292,N_29837,N_29888);
nand UO_2293 (O_2293,N_29235,N_29107);
xor UO_2294 (O_2294,N_29238,N_29154);
nor UO_2295 (O_2295,N_29362,N_29616);
xnor UO_2296 (O_2296,N_29071,N_29387);
nand UO_2297 (O_2297,N_29868,N_29483);
nor UO_2298 (O_2298,N_29138,N_29342);
and UO_2299 (O_2299,N_29418,N_29358);
xor UO_2300 (O_2300,N_29212,N_29914);
and UO_2301 (O_2301,N_29079,N_29552);
and UO_2302 (O_2302,N_29029,N_29671);
and UO_2303 (O_2303,N_29923,N_29344);
or UO_2304 (O_2304,N_29338,N_29885);
xor UO_2305 (O_2305,N_29819,N_29893);
xnor UO_2306 (O_2306,N_29552,N_29864);
or UO_2307 (O_2307,N_29160,N_29396);
nand UO_2308 (O_2308,N_29389,N_29233);
nand UO_2309 (O_2309,N_29837,N_29770);
and UO_2310 (O_2310,N_29378,N_29073);
or UO_2311 (O_2311,N_29146,N_29578);
and UO_2312 (O_2312,N_29687,N_29893);
or UO_2313 (O_2313,N_29224,N_29542);
nor UO_2314 (O_2314,N_29305,N_29664);
nor UO_2315 (O_2315,N_29852,N_29211);
or UO_2316 (O_2316,N_29629,N_29272);
nand UO_2317 (O_2317,N_29836,N_29129);
and UO_2318 (O_2318,N_29700,N_29724);
or UO_2319 (O_2319,N_29471,N_29002);
xnor UO_2320 (O_2320,N_29613,N_29474);
nor UO_2321 (O_2321,N_29649,N_29203);
xor UO_2322 (O_2322,N_29124,N_29462);
xnor UO_2323 (O_2323,N_29967,N_29516);
and UO_2324 (O_2324,N_29873,N_29929);
and UO_2325 (O_2325,N_29163,N_29458);
nor UO_2326 (O_2326,N_29872,N_29837);
nand UO_2327 (O_2327,N_29703,N_29168);
xor UO_2328 (O_2328,N_29136,N_29573);
nand UO_2329 (O_2329,N_29949,N_29241);
nand UO_2330 (O_2330,N_29168,N_29985);
and UO_2331 (O_2331,N_29017,N_29980);
or UO_2332 (O_2332,N_29714,N_29662);
or UO_2333 (O_2333,N_29456,N_29335);
xor UO_2334 (O_2334,N_29096,N_29905);
and UO_2335 (O_2335,N_29843,N_29750);
or UO_2336 (O_2336,N_29737,N_29867);
and UO_2337 (O_2337,N_29181,N_29505);
xor UO_2338 (O_2338,N_29855,N_29457);
nand UO_2339 (O_2339,N_29759,N_29741);
or UO_2340 (O_2340,N_29064,N_29753);
nand UO_2341 (O_2341,N_29936,N_29457);
or UO_2342 (O_2342,N_29923,N_29213);
nand UO_2343 (O_2343,N_29447,N_29600);
or UO_2344 (O_2344,N_29654,N_29460);
and UO_2345 (O_2345,N_29866,N_29895);
nor UO_2346 (O_2346,N_29386,N_29104);
nand UO_2347 (O_2347,N_29540,N_29482);
xnor UO_2348 (O_2348,N_29631,N_29388);
or UO_2349 (O_2349,N_29974,N_29178);
xor UO_2350 (O_2350,N_29872,N_29788);
and UO_2351 (O_2351,N_29173,N_29805);
nand UO_2352 (O_2352,N_29893,N_29401);
or UO_2353 (O_2353,N_29732,N_29450);
xnor UO_2354 (O_2354,N_29587,N_29897);
xor UO_2355 (O_2355,N_29545,N_29936);
and UO_2356 (O_2356,N_29242,N_29816);
xor UO_2357 (O_2357,N_29879,N_29324);
nor UO_2358 (O_2358,N_29396,N_29997);
nor UO_2359 (O_2359,N_29599,N_29187);
or UO_2360 (O_2360,N_29717,N_29212);
nor UO_2361 (O_2361,N_29526,N_29767);
nor UO_2362 (O_2362,N_29567,N_29683);
nand UO_2363 (O_2363,N_29149,N_29067);
xor UO_2364 (O_2364,N_29857,N_29519);
nor UO_2365 (O_2365,N_29369,N_29221);
and UO_2366 (O_2366,N_29706,N_29936);
and UO_2367 (O_2367,N_29629,N_29039);
nand UO_2368 (O_2368,N_29404,N_29050);
or UO_2369 (O_2369,N_29431,N_29252);
or UO_2370 (O_2370,N_29932,N_29889);
nor UO_2371 (O_2371,N_29852,N_29314);
or UO_2372 (O_2372,N_29299,N_29877);
nand UO_2373 (O_2373,N_29953,N_29359);
nand UO_2374 (O_2374,N_29566,N_29917);
or UO_2375 (O_2375,N_29979,N_29372);
and UO_2376 (O_2376,N_29627,N_29771);
nor UO_2377 (O_2377,N_29394,N_29802);
or UO_2378 (O_2378,N_29213,N_29226);
xnor UO_2379 (O_2379,N_29377,N_29067);
xor UO_2380 (O_2380,N_29538,N_29045);
xor UO_2381 (O_2381,N_29716,N_29024);
or UO_2382 (O_2382,N_29197,N_29931);
nand UO_2383 (O_2383,N_29656,N_29459);
xnor UO_2384 (O_2384,N_29616,N_29098);
nand UO_2385 (O_2385,N_29934,N_29332);
or UO_2386 (O_2386,N_29119,N_29222);
and UO_2387 (O_2387,N_29411,N_29113);
or UO_2388 (O_2388,N_29878,N_29532);
and UO_2389 (O_2389,N_29718,N_29112);
nand UO_2390 (O_2390,N_29443,N_29182);
and UO_2391 (O_2391,N_29342,N_29173);
nor UO_2392 (O_2392,N_29254,N_29701);
xnor UO_2393 (O_2393,N_29143,N_29261);
and UO_2394 (O_2394,N_29739,N_29722);
xor UO_2395 (O_2395,N_29326,N_29470);
nor UO_2396 (O_2396,N_29081,N_29706);
nand UO_2397 (O_2397,N_29154,N_29046);
or UO_2398 (O_2398,N_29752,N_29066);
or UO_2399 (O_2399,N_29349,N_29364);
nor UO_2400 (O_2400,N_29603,N_29671);
and UO_2401 (O_2401,N_29035,N_29166);
and UO_2402 (O_2402,N_29959,N_29900);
or UO_2403 (O_2403,N_29376,N_29561);
nand UO_2404 (O_2404,N_29157,N_29405);
or UO_2405 (O_2405,N_29394,N_29955);
and UO_2406 (O_2406,N_29850,N_29428);
xor UO_2407 (O_2407,N_29588,N_29422);
nor UO_2408 (O_2408,N_29511,N_29152);
nor UO_2409 (O_2409,N_29656,N_29259);
and UO_2410 (O_2410,N_29229,N_29521);
or UO_2411 (O_2411,N_29845,N_29947);
and UO_2412 (O_2412,N_29202,N_29725);
nand UO_2413 (O_2413,N_29549,N_29178);
xor UO_2414 (O_2414,N_29349,N_29050);
nor UO_2415 (O_2415,N_29672,N_29219);
or UO_2416 (O_2416,N_29079,N_29068);
nor UO_2417 (O_2417,N_29555,N_29699);
nand UO_2418 (O_2418,N_29734,N_29947);
nand UO_2419 (O_2419,N_29400,N_29864);
nor UO_2420 (O_2420,N_29304,N_29017);
nand UO_2421 (O_2421,N_29726,N_29721);
nand UO_2422 (O_2422,N_29228,N_29594);
nor UO_2423 (O_2423,N_29454,N_29213);
nand UO_2424 (O_2424,N_29952,N_29129);
nor UO_2425 (O_2425,N_29470,N_29146);
xnor UO_2426 (O_2426,N_29719,N_29829);
nor UO_2427 (O_2427,N_29405,N_29823);
nand UO_2428 (O_2428,N_29048,N_29109);
or UO_2429 (O_2429,N_29267,N_29546);
and UO_2430 (O_2430,N_29704,N_29139);
and UO_2431 (O_2431,N_29753,N_29781);
or UO_2432 (O_2432,N_29710,N_29804);
nand UO_2433 (O_2433,N_29572,N_29760);
nand UO_2434 (O_2434,N_29986,N_29346);
xor UO_2435 (O_2435,N_29624,N_29051);
or UO_2436 (O_2436,N_29322,N_29098);
and UO_2437 (O_2437,N_29848,N_29345);
nor UO_2438 (O_2438,N_29274,N_29139);
nand UO_2439 (O_2439,N_29155,N_29762);
and UO_2440 (O_2440,N_29986,N_29873);
nand UO_2441 (O_2441,N_29348,N_29665);
and UO_2442 (O_2442,N_29352,N_29910);
xor UO_2443 (O_2443,N_29811,N_29285);
and UO_2444 (O_2444,N_29214,N_29546);
nand UO_2445 (O_2445,N_29424,N_29935);
xnor UO_2446 (O_2446,N_29591,N_29780);
and UO_2447 (O_2447,N_29091,N_29696);
or UO_2448 (O_2448,N_29679,N_29296);
and UO_2449 (O_2449,N_29116,N_29215);
nor UO_2450 (O_2450,N_29883,N_29403);
and UO_2451 (O_2451,N_29202,N_29548);
and UO_2452 (O_2452,N_29758,N_29947);
nor UO_2453 (O_2453,N_29241,N_29749);
xor UO_2454 (O_2454,N_29179,N_29901);
nand UO_2455 (O_2455,N_29189,N_29815);
xnor UO_2456 (O_2456,N_29332,N_29450);
and UO_2457 (O_2457,N_29807,N_29258);
or UO_2458 (O_2458,N_29779,N_29092);
xnor UO_2459 (O_2459,N_29268,N_29857);
and UO_2460 (O_2460,N_29101,N_29957);
and UO_2461 (O_2461,N_29642,N_29199);
xor UO_2462 (O_2462,N_29442,N_29892);
nor UO_2463 (O_2463,N_29535,N_29108);
or UO_2464 (O_2464,N_29561,N_29790);
xor UO_2465 (O_2465,N_29599,N_29762);
or UO_2466 (O_2466,N_29200,N_29860);
or UO_2467 (O_2467,N_29365,N_29624);
nor UO_2468 (O_2468,N_29471,N_29382);
nand UO_2469 (O_2469,N_29378,N_29031);
or UO_2470 (O_2470,N_29973,N_29712);
and UO_2471 (O_2471,N_29920,N_29890);
xnor UO_2472 (O_2472,N_29230,N_29440);
nor UO_2473 (O_2473,N_29841,N_29089);
or UO_2474 (O_2474,N_29706,N_29590);
and UO_2475 (O_2475,N_29029,N_29790);
nand UO_2476 (O_2476,N_29583,N_29301);
or UO_2477 (O_2477,N_29432,N_29750);
and UO_2478 (O_2478,N_29462,N_29850);
and UO_2479 (O_2479,N_29709,N_29698);
xnor UO_2480 (O_2480,N_29620,N_29837);
xor UO_2481 (O_2481,N_29273,N_29391);
nor UO_2482 (O_2482,N_29611,N_29819);
and UO_2483 (O_2483,N_29026,N_29967);
xor UO_2484 (O_2484,N_29992,N_29526);
nor UO_2485 (O_2485,N_29041,N_29640);
nor UO_2486 (O_2486,N_29758,N_29107);
and UO_2487 (O_2487,N_29072,N_29831);
and UO_2488 (O_2488,N_29602,N_29333);
nor UO_2489 (O_2489,N_29534,N_29084);
or UO_2490 (O_2490,N_29854,N_29477);
nand UO_2491 (O_2491,N_29201,N_29803);
and UO_2492 (O_2492,N_29262,N_29645);
and UO_2493 (O_2493,N_29748,N_29587);
nand UO_2494 (O_2494,N_29433,N_29352);
or UO_2495 (O_2495,N_29078,N_29599);
nand UO_2496 (O_2496,N_29219,N_29514);
nand UO_2497 (O_2497,N_29124,N_29151);
or UO_2498 (O_2498,N_29553,N_29236);
xnor UO_2499 (O_2499,N_29761,N_29081);
and UO_2500 (O_2500,N_29985,N_29093);
or UO_2501 (O_2501,N_29000,N_29674);
nor UO_2502 (O_2502,N_29923,N_29423);
nand UO_2503 (O_2503,N_29541,N_29693);
nor UO_2504 (O_2504,N_29095,N_29232);
or UO_2505 (O_2505,N_29967,N_29018);
xnor UO_2506 (O_2506,N_29968,N_29717);
xor UO_2507 (O_2507,N_29517,N_29293);
nand UO_2508 (O_2508,N_29466,N_29848);
or UO_2509 (O_2509,N_29154,N_29745);
or UO_2510 (O_2510,N_29186,N_29265);
or UO_2511 (O_2511,N_29712,N_29187);
nand UO_2512 (O_2512,N_29734,N_29156);
xor UO_2513 (O_2513,N_29398,N_29480);
nand UO_2514 (O_2514,N_29336,N_29605);
nand UO_2515 (O_2515,N_29234,N_29275);
xnor UO_2516 (O_2516,N_29448,N_29272);
xnor UO_2517 (O_2517,N_29723,N_29847);
or UO_2518 (O_2518,N_29137,N_29300);
and UO_2519 (O_2519,N_29701,N_29845);
nand UO_2520 (O_2520,N_29116,N_29061);
xnor UO_2521 (O_2521,N_29885,N_29851);
nand UO_2522 (O_2522,N_29435,N_29918);
xor UO_2523 (O_2523,N_29604,N_29989);
and UO_2524 (O_2524,N_29590,N_29218);
or UO_2525 (O_2525,N_29227,N_29481);
xnor UO_2526 (O_2526,N_29622,N_29443);
or UO_2527 (O_2527,N_29579,N_29607);
or UO_2528 (O_2528,N_29877,N_29327);
and UO_2529 (O_2529,N_29189,N_29779);
nand UO_2530 (O_2530,N_29805,N_29301);
xor UO_2531 (O_2531,N_29514,N_29570);
or UO_2532 (O_2532,N_29557,N_29210);
or UO_2533 (O_2533,N_29019,N_29253);
or UO_2534 (O_2534,N_29753,N_29080);
xnor UO_2535 (O_2535,N_29504,N_29879);
or UO_2536 (O_2536,N_29018,N_29733);
xor UO_2537 (O_2537,N_29529,N_29193);
nand UO_2538 (O_2538,N_29891,N_29019);
xnor UO_2539 (O_2539,N_29558,N_29078);
and UO_2540 (O_2540,N_29623,N_29896);
or UO_2541 (O_2541,N_29495,N_29016);
and UO_2542 (O_2542,N_29768,N_29566);
and UO_2543 (O_2543,N_29510,N_29342);
nor UO_2544 (O_2544,N_29118,N_29656);
nor UO_2545 (O_2545,N_29325,N_29015);
xor UO_2546 (O_2546,N_29452,N_29075);
or UO_2547 (O_2547,N_29241,N_29778);
nand UO_2548 (O_2548,N_29789,N_29300);
and UO_2549 (O_2549,N_29659,N_29145);
nor UO_2550 (O_2550,N_29726,N_29702);
and UO_2551 (O_2551,N_29817,N_29225);
xor UO_2552 (O_2552,N_29063,N_29152);
and UO_2553 (O_2553,N_29721,N_29105);
or UO_2554 (O_2554,N_29659,N_29237);
nor UO_2555 (O_2555,N_29811,N_29156);
and UO_2556 (O_2556,N_29737,N_29457);
and UO_2557 (O_2557,N_29448,N_29040);
nand UO_2558 (O_2558,N_29470,N_29786);
nor UO_2559 (O_2559,N_29812,N_29315);
xor UO_2560 (O_2560,N_29782,N_29821);
nor UO_2561 (O_2561,N_29375,N_29113);
or UO_2562 (O_2562,N_29161,N_29915);
nor UO_2563 (O_2563,N_29496,N_29958);
or UO_2564 (O_2564,N_29305,N_29285);
and UO_2565 (O_2565,N_29456,N_29683);
xnor UO_2566 (O_2566,N_29870,N_29733);
xnor UO_2567 (O_2567,N_29568,N_29984);
nand UO_2568 (O_2568,N_29810,N_29949);
and UO_2569 (O_2569,N_29348,N_29507);
nor UO_2570 (O_2570,N_29856,N_29102);
and UO_2571 (O_2571,N_29411,N_29997);
nand UO_2572 (O_2572,N_29489,N_29331);
or UO_2573 (O_2573,N_29994,N_29980);
or UO_2574 (O_2574,N_29459,N_29110);
or UO_2575 (O_2575,N_29847,N_29907);
or UO_2576 (O_2576,N_29061,N_29765);
or UO_2577 (O_2577,N_29168,N_29155);
nand UO_2578 (O_2578,N_29640,N_29199);
nand UO_2579 (O_2579,N_29535,N_29254);
nand UO_2580 (O_2580,N_29785,N_29231);
and UO_2581 (O_2581,N_29280,N_29319);
xor UO_2582 (O_2582,N_29877,N_29774);
nand UO_2583 (O_2583,N_29382,N_29328);
and UO_2584 (O_2584,N_29813,N_29481);
or UO_2585 (O_2585,N_29856,N_29890);
nor UO_2586 (O_2586,N_29084,N_29489);
xor UO_2587 (O_2587,N_29799,N_29900);
and UO_2588 (O_2588,N_29252,N_29891);
nor UO_2589 (O_2589,N_29957,N_29420);
or UO_2590 (O_2590,N_29013,N_29058);
and UO_2591 (O_2591,N_29652,N_29379);
nor UO_2592 (O_2592,N_29091,N_29176);
nand UO_2593 (O_2593,N_29378,N_29132);
or UO_2594 (O_2594,N_29098,N_29165);
xnor UO_2595 (O_2595,N_29685,N_29861);
and UO_2596 (O_2596,N_29438,N_29115);
or UO_2597 (O_2597,N_29992,N_29831);
nand UO_2598 (O_2598,N_29998,N_29534);
or UO_2599 (O_2599,N_29311,N_29001);
or UO_2600 (O_2600,N_29273,N_29428);
nor UO_2601 (O_2601,N_29641,N_29892);
or UO_2602 (O_2602,N_29403,N_29202);
nor UO_2603 (O_2603,N_29064,N_29469);
nand UO_2604 (O_2604,N_29074,N_29518);
or UO_2605 (O_2605,N_29142,N_29801);
xor UO_2606 (O_2606,N_29539,N_29650);
xor UO_2607 (O_2607,N_29981,N_29295);
and UO_2608 (O_2608,N_29825,N_29018);
nand UO_2609 (O_2609,N_29037,N_29596);
or UO_2610 (O_2610,N_29051,N_29950);
nor UO_2611 (O_2611,N_29581,N_29072);
nor UO_2612 (O_2612,N_29895,N_29753);
xor UO_2613 (O_2613,N_29640,N_29447);
and UO_2614 (O_2614,N_29449,N_29003);
or UO_2615 (O_2615,N_29766,N_29802);
and UO_2616 (O_2616,N_29736,N_29069);
nor UO_2617 (O_2617,N_29079,N_29323);
nor UO_2618 (O_2618,N_29361,N_29561);
nor UO_2619 (O_2619,N_29282,N_29525);
and UO_2620 (O_2620,N_29402,N_29914);
xnor UO_2621 (O_2621,N_29232,N_29924);
nand UO_2622 (O_2622,N_29419,N_29696);
and UO_2623 (O_2623,N_29301,N_29872);
xnor UO_2624 (O_2624,N_29926,N_29535);
xor UO_2625 (O_2625,N_29182,N_29899);
or UO_2626 (O_2626,N_29866,N_29817);
and UO_2627 (O_2627,N_29503,N_29334);
xor UO_2628 (O_2628,N_29932,N_29682);
nor UO_2629 (O_2629,N_29454,N_29755);
and UO_2630 (O_2630,N_29640,N_29951);
nor UO_2631 (O_2631,N_29169,N_29307);
xnor UO_2632 (O_2632,N_29181,N_29783);
nor UO_2633 (O_2633,N_29677,N_29349);
nand UO_2634 (O_2634,N_29941,N_29102);
nand UO_2635 (O_2635,N_29367,N_29192);
nor UO_2636 (O_2636,N_29612,N_29268);
nand UO_2637 (O_2637,N_29166,N_29890);
and UO_2638 (O_2638,N_29433,N_29078);
xor UO_2639 (O_2639,N_29513,N_29682);
nor UO_2640 (O_2640,N_29260,N_29925);
nor UO_2641 (O_2641,N_29388,N_29099);
xnor UO_2642 (O_2642,N_29264,N_29047);
and UO_2643 (O_2643,N_29108,N_29040);
or UO_2644 (O_2644,N_29003,N_29232);
and UO_2645 (O_2645,N_29872,N_29184);
and UO_2646 (O_2646,N_29146,N_29936);
and UO_2647 (O_2647,N_29487,N_29803);
nand UO_2648 (O_2648,N_29018,N_29682);
or UO_2649 (O_2649,N_29470,N_29711);
or UO_2650 (O_2650,N_29887,N_29098);
and UO_2651 (O_2651,N_29258,N_29199);
or UO_2652 (O_2652,N_29389,N_29204);
xor UO_2653 (O_2653,N_29365,N_29525);
and UO_2654 (O_2654,N_29271,N_29261);
xor UO_2655 (O_2655,N_29378,N_29428);
nand UO_2656 (O_2656,N_29995,N_29386);
nor UO_2657 (O_2657,N_29740,N_29234);
xnor UO_2658 (O_2658,N_29418,N_29210);
xnor UO_2659 (O_2659,N_29862,N_29485);
nor UO_2660 (O_2660,N_29580,N_29174);
or UO_2661 (O_2661,N_29295,N_29348);
nor UO_2662 (O_2662,N_29011,N_29035);
or UO_2663 (O_2663,N_29731,N_29777);
nor UO_2664 (O_2664,N_29775,N_29687);
and UO_2665 (O_2665,N_29240,N_29286);
xor UO_2666 (O_2666,N_29242,N_29400);
xor UO_2667 (O_2667,N_29922,N_29669);
xnor UO_2668 (O_2668,N_29786,N_29889);
xor UO_2669 (O_2669,N_29159,N_29994);
or UO_2670 (O_2670,N_29097,N_29859);
nor UO_2671 (O_2671,N_29690,N_29409);
and UO_2672 (O_2672,N_29073,N_29142);
xor UO_2673 (O_2673,N_29426,N_29776);
nor UO_2674 (O_2674,N_29687,N_29455);
nand UO_2675 (O_2675,N_29048,N_29828);
and UO_2676 (O_2676,N_29649,N_29691);
xor UO_2677 (O_2677,N_29922,N_29714);
nand UO_2678 (O_2678,N_29529,N_29489);
and UO_2679 (O_2679,N_29401,N_29687);
and UO_2680 (O_2680,N_29018,N_29770);
nand UO_2681 (O_2681,N_29801,N_29619);
nor UO_2682 (O_2682,N_29782,N_29682);
and UO_2683 (O_2683,N_29324,N_29660);
or UO_2684 (O_2684,N_29196,N_29715);
and UO_2685 (O_2685,N_29708,N_29938);
nand UO_2686 (O_2686,N_29664,N_29794);
nor UO_2687 (O_2687,N_29876,N_29287);
xor UO_2688 (O_2688,N_29902,N_29442);
and UO_2689 (O_2689,N_29305,N_29752);
and UO_2690 (O_2690,N_29126,N_29451);
nand UO_2691 (O_2691,N_29938,N_29000);
nor UO_2692 (O_2692,N_29604,N_29009);
and UO_2693 (O_2693,N_29882,N_29871);
nor UO_2694 (O_2694,N_29015,N_29176);
and UO_2695 (O_2695,N_29771,N_29034);
and UO_2696 (O_2696,N_29658,N_29960);
nor UO_2697 (O_2697,N_29774,N_29585);
and UO_2698 (O_2698,N_29251,N_29364);
or UO_2699 (O_2699,N_29489,N_29585);
or UO_2700 (O_2700,N_29931,N_29307);
nand UO_2701 (O_2701,N_29537,N_29966);
or UO_2702 (O_2702,N_29168,N_29532);
nand UO_2703 (O_2703,N_29520,N_29936);
and UO_2704 (O_2704,N_29498,N_29922);
or UO_2705 (O_2705,N_29914,N_29625);
and UO_2706 (O_2706,N_29743,N_29944);
and UO_2707 (O_2707,N_29325,N_29385);
or UO_2708 (O_2708,N_29576,N_29981);
and UO_2709 (O_2709,N_29314,N_29725);
nor UO_2710 (O_2710,N_29225,N_29553);
nor UO_2711 (O_2711,N_29079,N_29007);
and UO_2712 (O_2712,N_29525,N_29489);
nor UO_2713 (O_2713,N_29379,N_29356);
xor UO_2714 (O_2714,N_29418,N_29566);
or UO_2715 (O_2715,N_29383,N_29703);
nor UO_2716 (O_2716,N_29745,N_29928);
nand UO_2717 (O_2717,N_29496,N_29311);
or UO_2718 (O_2718,N_29278,N_29625);
xor UO_2719 (O_2719,N_29206,N_29819);
nand UO_2720 (O_2720,N_29532,N_29236);
xor UO_2721 (O_2721,N_29624,N_29541);
nand UO_2722 (O_2722,N_29585,N_29346);
nor UO_2723 (O_2723,N_29498,N_29952);
or UO_2724 (O_2724,N_29634,N_29049);
nor UO_2725 (O_2725,N_29875,N_29554);
or UO_2726 (O_2726,N_29909,N_29235);
xnor UO_2727 (O_2727,N_29804,N_29099);
nand UO_2728 (O_2728,N_29762,N_29955);
xor UO_2729 (O_2729,N_29972,N_29827);
nor UO_2730 (O_2730,N_29954,N_29094);
nor UO_2731 (O_2731,N_29459,N_29556);
nand UO_2732 (O_2732,N_29895,N_29513);
and UO_2733 (O_2733,N_29239,N_29205);
or UO_2734 (O_2734,N_29179,N_29627);
or UO_2735 (O_2735,N_29727,N_29766);
nand UO_2736 (O_2736,N_29759,N_29557);
nand UO_2737 (O_2737,N_29398,N_29958);
or UO_2738 (O_2738,N_29920,N_29775);
nand UO_2739 (O_2739,N_29420,N_29998);
xor UO_2740 (O_2740,N_29019,N_29987);
and UO_2741 (O_2741,N_29880,N_29631);
nand UO_2742 (O_2742,N_29510,N_29269);
xor UO_2743 (O_2743,N_29000,N_29956);
nor UO_2744 (O_2744,N_29874,N_29187);
nor UO_2745 (O_2745,N_29793,N_29988);
nor UO_2746 (O_2746,N_29132,N_29020);
nand UO_2747 (O_2747,N_29123,N_29614);
and UO_2748 (O_2748,N_29374,N_29608);
nand UO_2749 (O_2749,N_29741,N_29115);
xor UO_2750 (O_2750,N_29807,N_29784);
and UO_2751 (O_2751,N_29361,N_29317);
nor UO_2752 (O_2752,N_29395,N_29741);
nor UO_2753 (O_2753,N_29385,N_29144);
xor UO_2754 (O_2754,N_29254,N_29034);
nor UO_2755 (O_2755,N_29634,N_29757);
xnor UO_2756 (O_2756,N_29135,N_29831);
or UO_2757 (O_2757,N_29115,N_29390);
or UO_2758 (O_2758,N_29547,N_29890);
nor UO_2759 (O_2759,N_29259,N_29500);
xnor UO_2760 (O_2760,N_29502,N_29759);
xor UO_2761 (O_2761,N_29858,N_29887);
and UO_2762 (O_2762,N_29313,N_29835);
nor UO_2763 (O_2763,N_29717,N_29852);
and UO_2764 (O_2764,N_29403,N_29492);
nand UO_2765 (O_2765,N_29920,N_29200);
nand UO_2766 (O_2766,N_29635,N_29803);
xor UO_2767 (O_2767,N_29322,N_29937);
or UO_2768 (O_2768,N_29023,N_29455);
xor UO_2769 (O_2769,N_29625,N_29838);
nand UO_2770 (O_2770,N_29874,N_29846);
or UO_2771 (O_2771,N_29230,N_29003);
nor UO_2772 (O_2772,N_29590,N_29398);
nor UO_2773 (O_2773,N_29240,N_29987);
and UO_2774 (O_2774,N_29943,N_29543);
nand UO_2775 (O_2775,N_29109,N_29053);
or UO_2776 (O_2776,N_29155,N_29882);
nand UO_2777 (O_2777,N_29370,N_29056);
or UO_2778 (O_2778,N_29196,N_29188);
nand UO_2779 (O_2779,N_29796,N_29825);
xor UO_2780 (O_2780,N_29105,N_29363);
xor UO_2781 (O_2781,N_29971,N_29850);
nand UO_2782 (O_2782,N_29030,N_29750);
or UO_2783 (O_2783,N_29627,N_29761);
nand UO_2784 (O_2784,N_29384,N_29046);
nand UO_2785 (O_2785,N_29260,N_29305);
nand UO_2786 (O_2786,N_29048,N_29290);
nor UO_2787 (O_2787,N_29891,N_29450);
xnor UO_2788 (O_2788,N_29704,N_29735);
nand UO_2789 (O_2789,N_29217,N_29594);
nand UO_2790 (O_2790,N_29226,N_29064);
nor UO_2791 (O_2791,N_29295,N_29267);
nand UO_2792 (O_2792,N_29213,N_29949);
or UO_2793 (O_2793,N_29147,N_29092);
and UO_2794 (O_2794,N_29516,N_29298);
or UO_2795 (O_2795,N_29152,N_29930);
or UO_2796 (O_2796,N_29048,N_29467);
xnor UO_2797 (O_2797,N_29255,N_29507);
and UO_2798 (O_2798,N_29724,N_29219);
xor UO_2799 (O_2799,N_29204,N_29856);
or UO_2800 (O_2800,N_29957,N_29976);
nand UO_2801 (O_2801,N_29380,N_29706);
nor UO_2802 (O_2802,N_29921,N_29800);
nand UO_2803 (O_2803,N_29806,N_29460);
and UO_2804 (O_2804,N_29805,N_29186);
nor UO_2805 (O_2805,N_29188,N_29451);
and UO_2806 (O_2806,N_29424,N_29107);
and UO_2807 (O_2807,N_29516,N_29562);
and UO_2808 (O_2808,N_29371,N_29357);
and UO_2809 (O_2809,N_29557,N_29213);
xor UO_2810 (O_2810,N_29138,N_29932);
or UO_2811 (O_2811,N_29618,N_29366);
and UO_2812 (O_2812,N_29782,N_29125);
xor UO_2813 (O_2813,N_29459,N_29756);
or UO_2814 (O_2814,N_29919,N_29367);
nor UO_2815 (O_2815,N_29977,N_29409);
xor UO_2816 (O_2816,N_29175,N_29066);
or UO_2817 (O_2817,N_29107,N_29297);
and UO_2818 (O_2818,N_29829,N_29256);
xnor UO_2819 (O_2819,N_29372,N_29172);
or UO_2820 (O_2820,N_29677,N_29255);
xnor UO_2821 (O_2821,N_29561,N_29441);
or UO_2822 (O_2822,N_29668,N_29178);
and UO_2823 (O_2823,N_29897,N_29612);
xor UO_2824 (O_2824,N_29456,N_29237);
nand UO_2825 (O_2825,N_29069,N_29379);
or UO_2826 (O_2826,N_29625,N_29514);
nor UO_2827 (O_2827,N_29628,N_29545);
nand UO_2828 (O_2828,N_29181,N_29082);
xnor UO_2829 (O_2829,N_29456,N_29749);
nor UO_2830 (O_2830,N_29162,N_29393);
xor UO_2831 (O_2831,N_29840,N_29448);
nand UO_2832 (O_2832,N_29633,N_29089);
or UO_2833 (O_2833,N_29805,N_29849);
nand UO_2834 (O_2834,N_29774,N_29227);
xnor UO_2835 (O_2835,N_29848,N_29182);
nor UO_2836 (O_2836,N_29760,N_29817);
or UO_2837 (O_2837,N_29978,N_29571);
xnor UO_2838 (O_2838,N_29528,N_29753);
or UO_2839 (O_2839,N_29341,N_29028);
and UO_2840 (O_2840,N_29698,N_29885);
xnor UO_2841 (O_2841,N_29213,N_29520);
nor UO_2842 (O_2842,N_29211,N_29360);
or UO_2843 (O_2843,N_29620,N_29251);
or UO_2844 (O_2844,N_29472,N_29906);
nor UO_2845 (O_2845,N_29575,N_29786);
xor UO_2846 (O_2846,N_29378,N_29124);
and UO_2847 (O_2847,N_29914,N_29357);
or UO_2848 (O_2848,N_29504,N_29318);
or UO_2849 (O_2849,N_29072,N_29832);
nor UO_2850 (O_2850,N_29870,N_29309);
xnor UO_2851 (O_2851,N_29107,N_29081);
nand UO_2852 (O_2852,N_29700,N_29815);
and UO_2853 (O_2853,N_29397,N_29517);
xnor UO_2854 (O_2854,N_29474,N_29384);
or UO_2855 (O_2855,N_29815,N_29934);
and UO_2856 (O_2856,N_29944,N_29834);
and UO_2857 (O_2857,N_29971,N_29753);
nor UO_2858 (O_2858,N_29038,N_29947);
nor UO_2859 (O_2859,N_29738,N_29988);
and UO_2860 (O_2860,N_29797,N_29292);
and UO_2861 (O_2861,N_29567,N_29555);
nand UO_2862 (O_2862,N_29036,N_29680);
and UO_2863 (O_2863,N_29140,N_29199);
xor UO_2864 (O_2864,N_29917,N_29843);
nand UO_2865 (O_2865,N_29290,N_29469);
nand UO_2866 (O_2866,N_29427,N_29649);
nor UO_2867 (O_2867,N_29667,N_29197);
nand UO_2868 (O_2868,N_29030,N_29861);
and UO_2869 (O_2869,N_29595,N_29208);
and UO_2870 (O_2870,N_29202,N_29398);
and UO_2871 (O_2871,N_29648,N_29831);
or UO_2872 (O_2872,N_29054,N_29976);
nor UO_2873 (O_2873,N_29935,N_29120);
nand UO_2874 (O_2874,N_29042,N_29618);
nand UO_2875 (O_2875,N_29714,N_29242);
and UO_2876 (O_2876,N_29642,N_29994);
xor UO_2877 (O_2877,N_29917,N_29682);
nand UO_2878 (O_2878,N_29164,N_29145);
xnor UO_2879 (O_2879,N_29943,N_29732);
xnor UO_2880 (O_2880,N_29430,N_29961);
nand UO_2881 (O_2881,N_29249,N_29224);
nand UO_2882 (O_2882,N_29739,N_29392);
nand UO_2883 (O_2883,N_29805,N_29966);
or UO_2884 (O_2884,N_29726,N_29116);
nand UO_2885 (O_2885,N_29408,N_29197);
nor UO_2886 (O_2886,N_29695,N_29637);
nand UO_2887 (O_2887,N_29815,N_29798);
nor UO_2888 (O_2888,N_29012,N_29869);
nand UO_2889 (O_2889,N_29494,N_29444);
nor UO_2890 (O_2890,N_29049,N_29861);
or UO_2891 (O_2891,N_29590,N_29501);
and UO_2892 (O_2892,N_29356,N_29837);
xnor UO_2893 (O_2893,N_29138,N_29141);
nor UO_2894 (O_2894,N_29054,N_29397);
nor UO_2895 (O_2895,N_29493,N_29016);
nand UO_2896 (O_2896,N_29954,N_29916);
and UO_2897 (O_2897,N_29311,N_29080);
xnor UO_2898 (O_2898,N_29535,N_29568);
and UO_2899 (O_2899,N_29477,N_29426);
nand UO_2900 (O_2900,N_29472,N_29423);
nand UO_2901 (O_2901,N_29684,N_29302);
nand UO_2902 (O_2902,N_29045,N_29316);
nand UO_2903 (O_2903,N_29112,N_29139);
xor UO_2904 (O_2904,N_29245,N_29996);
or UO_2905 (O_2905,N_29858,N_29430);
and UO_2906 (O_2906,N_29973,N_29923);
or UO_2907 (O_2907,N_29290,N_29178);
xnor UO_2908 (O_2908,N_29285,N_29612);
xnor UO_2909 (O_2909,N_29865,N_29498);
nand UO_2910 (O_2910,N_29644,N_29798);
nor UO_2911 (O_2911,N_29934,N_29675);
nand UO_2912 (O_2912,N_29310,N_29558);
xor UO_2913 (O_2913,N_29697,N_29290);
xor UO_2914 (O_2914,N_29562,N_29971);
xnor UO_2915 (O_2915,N_29204,N_29486);
or UO_2916 (O_2916,N_29582,N_29970);
nand UO_2917 (O_2917,N_29595,N_29080);
or UO_2918 (O_2918,N_29286,N_29971);
nand UO_2919 (O_2919,N_29290,N_29333);
xor UO_2920 (O_2920,N_29349,N_29620);
xor UO_2921 (O_2921,N_29069,N_29400);
nand UO_2922 (O_2922,N_29153,N_29559);
nor UO_2923 (O_2923,N_29094,N_29798);
nor UO_2924 (O_2924,N_29553,N_29874);
nor UO_2925 (O_2925,N_29327,N_29910);
xnor UO_2926 (O_2926,N_29489,N_29387);
nor UO_2927 (O_2927,N_29270,N_29109);
xnor UO_2928 (O_2928,N_29633,N_29442);
nor UO_2929 (O_2929,N_29021,N_29186);
nor UO_2930 (O_2930,N_29685,N_29879);
and UO_2931 (O_2931,N_29381,N_29232);
or UO_2932 (O_2932,N_29363,N_29427);
or UO_2933 (O_2933,N_29658,N_29229);
nor UO_2934 (O_2934,N_29903,N_29811);
or UO_2935 (O_2935,N_29555,N_29456);
and UO_2936 (O_2936,N_29579,N_29253);
or UO_2937 (O_2937,N_29514,N_29300);
or UO_2938 (O_2938,N_29390,N_29235);
xor UO_2939 (O_2939,N_29936,N_29897);
nand UO_2940 (O_2940,N_29163,N_29703);
nand UO_2941 (O_2941,N_29154,N_29488);
nand UO_2942 (O_2942,N_29312,N_29892);
nand UO_2943 (O_2943,N_29297,N_29988);
or UO_2944 (O_2944,N_29101,N_29687);
or UO_2945 (O_2945,N_29876,N_29899);
nand UO_2946 (O_2946,N_29888,N_29149);
or UO_2947 (O_2947,N_29580,N_29248);
or UO_2948 (O_2948,N_29311,N_29584);
nor UO_2949 (O_2949,N_29056,N_29091);
nor UO_2950 (O_2950,N_29030,N_29054);
and UO_2951 (O_2951,N_29287,N_29847);
nor UO_2952 (O_2952,N_29282,N_29344);
and UO_2953 (O_2953,N_29385,N_29215);
nor UO_2954 (O_2954,N_29383,N_29990);
nand UO_2955 (O_2955,N_29878,N_29806);
nor UO_2956 (O_2956,N_29854,N_29405);
nand UO_2957 (O_2957,N_29684,N_29275);
and UO_2958 (O_2958,N_29985,N_29404);
and UO_2959 (O_2959,N_29146,N_29896);
nand UO_2960 (O_2960,N_29817,N_29950);
or UO_2961 (O_2961,N_29827,N_29012);
or UO_2962 (O_2962,N_29154,N_29719);
and UO_2963 (O_2963,N_29236,N_29202);
nand UO_2964 (O_2964,N_29397,N_29480);
or UO_2965 (O_2965,N_29391,N_29849);
and UO_2966 (O_2966,N_29641,N_29895);
and UO_2967 (O_2967,N_29521,N_29067);
nor UO_2968 (O_2968,N_29491,N_29973);
and UO_2969 (O_2969,N_29282,N_29096);
or UO_2970 (O_2970,N_29147,N_29752);
nand UO_2971 (O_2971,N_29761,N_29339);
and UO_2972 (O_2972,N_29073,N_29314);
or UO_2973 (O_2973,N_29475,N_29793);
nor UO_2974 (O_2974,N_29956,N_29092);
and UO_2975 (O_2975,N_29737,N_29045);
nor UO_2976 (O_2976,N_29561,N_29457);
nand UO_2977 (O_2977,N_29476,N_29260);
xnor UO_2978 (O_2978,N_29408,N_29317);
nor UO_2979 (O_2979,N_29471,N_29652);
and UO_2980 (O_2980,N_29151,N_29564);
and UO_2981 (O_2981,N_29261,N_29633);
and UO_2982 (O_2982,N_29113,N_29242);
nor UO_2983 (O_2983,N_29105,N_29998);
and UO_2984 (O_2984,N_29030,N_29214);
or UO_2985 (O_2985,N_29825,N_29656);
or UO_2986 (O_2986,N_29013,N_29138);
nor UO_2987 (O_2987,N_29233,N_29009);
nand UO_2988 (O_2988,N_29199,N_29002);
nor UO_2989 (O_2989,N_29107,N_29771);
nand UO_2990 (O_2990,N_29817,N_29498);
xnor UO_2991 (O_2991,N_29367,N_29846);
or UO_2992 (O_2992,N_29937,N_29869);
nor UO_2993 (O_2993,N_29164,N_29820);
nand UO_2994 (O_2994,N_29795,N_29563);
xor UO_2995 (O_2995,N_29047,N_29537);
or UO_2996 (O_2996,N_29470,N_29263);
xnor UO_2997 (O_2997,N_29376,N_29273);
or UO_2998 (O_2998,N_29662,N_29272);
or UO_2999 (O_2999,N_29574,N_29254);
and UO_3000 (O_3000,N_29283,N_29131);
nand UO_3001 (O_3001,N_29178,N_29052);
or UO_3002 (O_3002,N_29860,N_29437);
xnor UO_3003 (O_3003,N_29649,N_29037);
and UO_3004 (O_3004,N_29303,N_29633);
and UO_3005 (O_3005,N_29312,N_29542);
nor UO_3006 (O_3006,N_29050,N_29684);
or UO_3007 (O_3007,N_29102,N_29037);
nand UO_3008 (O_3008,N_29906,N_29622);
nor UO_3009 (O_3009,N_29147,N_29933);
and UO_3010 (O_3010,N_29626,N_29012);
xor UO_3011 (O_3011,N_29719,N_29534);
nor UO_3012 (O_3012,N_29954,N_29503);
xor UO_3013 (O_3013,N_29502,N_29630);
xnor UO_3014 (O_3014,N_29692,N_29815);
nor UO_3015 (O_3015,N_29734,N_29290);
xor UO_3016 (O_3016,N_29009,N_29513);
and UO_3017 (O_3017,N_29578,N_29202);
nand UO_3018 (O_3018,N_29521,N_29804);
nand UO_3019 (O_3019,N_29907,N_29278);
xor UO_3020 (O_3020,N_29788,N_29848);
nor UO_3021 (O_3021,N_29864,N_29744);
or UO_3022 (O_3022,N_29300,N_29829);
nor UO_3023 (O_3023,N_29070,N_29165);
nand UO_3024 (O_3024,N_29741,N_29749);
and UO_3025 (O_3025,N_29638,N_29300);
and UO_3026 (O_3026,N_29720,N_29247);
nand UO_3027 (O_3027,N_29996,N_29863);
nand UO_3028 (O_3028,N_29193,N_29361);
nor UO_3029 (O_3029,N_29081,N_29376);
and UO_3030 (O_3030,N_29120,N_29752);
nor UO_3031 (O_3031,N_29461,N_29366);
xnor UO_3032 (O_3032,N_29577,N_29512);
or UO_3033 (O_3033,N_29901,N_29439);
nor UO_3034 (O_3034,N_29354,N_29471);
nand UO_3035 (O_3035,N_29010,N_29147);
nand UO_3036 (O_3036,N_29059,N_29605);
nor UO_3037 (O_3037,N_29347,N_29566);
xor UO_3038 (O_3038,N_29736,N_29716);
or UO_3039 (O_3039,N_29648,N_29769);
or UO_3040 (O_3040,N_29438,N_29686);
nand UO_3041 (O_3041,N_29412,N_29190);
xor UO_3042 (O_3042,N_29421,N_29482);
nand UO_3043 (O_3043,N_29648,N_29424);
nand UO_3044 (O_3044,N_29275,N_29100);
and UO_3045 (O_3045,N_29640,N_29809);
and UO_3046 (O_3046,N_29928,N_29264);
nor UO_3047 (O_3047,N_29619,N_29368);
xnor UO_3048 (O_3048,N_29148,N_29749);
and UO_3049 (O_3049,N_29332,N_29251);
nor UO_3050 (O_3050,N_29684,N_29986);
xnor UO_3051 (O_3051,N_29960,N_29951);
nor UO_3052 (O_3052,N_29752,N_29428);
xnor UO_3053 (O_3053,N_29503,N_29781);
xor UO_3054 (O_3054,N_29311,N_29749);
nor UO_3055 (O_3055,N_29698,N_29529);
or UO_3056 (O_3056,N_29257,N_29240);
and UO_3057 (O_3057,N_29324,N_29415);
nand UO_3058 (O_3058,N_29110,N_29325);
nor UO_3059 (O_3059,N_29003,N_29812);
or UO_3060 (O_3060,N_29058,N_29371);
nand UO_3061 (O_3061,N_29129,N_29130);
and UO_3062 (O_3062,N_29631,N_29312);
xnor UO_3063 (O_3063,N_29837,N_29116);
nand UO_3064 (O_3064,N_29486,N_29988);
or UO_3065 (O_3065,N_29690,N_29415);
nor UO_3066 (O_3066,N_29238,N_29012);
or UO_3067 (O_3067,N_29737,N_29339);
and UO_3068 (O_3068,N_29296,N_29420);
and UO_3069 (O_3069,N_29041,N_29568);
or UO_3070 (O_3070,N_29598,N_29985);
nand UO_3071 (O_3071,N_29734,N_29824);
nor UO_3072 (O_3072,N_29096,N_29474);
xnor UO_3073 (O_3073,N_29185,N_29656);
nor UO_3074 (O_3074,N_29101,N_29244);
nand UO_3075 (O_3075,N_29025,N_29761);
nor UO_3076 (O_3076,N_29944,N_29454);
or UO_3077 (O_3077,N_29601,N_29472);
nor UO_3078 (O_3078,N_29784,N_29854);
nand UO_3079 (O_3079,N_29127,N_29457);
nor UO_3080 (O_3080,N_29814,N_29773);
xor UO_3081 (O_3081,N_29318,N_29009);
nor UO_3082 (O_3082,N_29106,N_29553);
or UO_3083 (O_3083,N_29175,N_29876);
and UO_3084 (O_3084,N_29703,N_29388);
nor UO_3085 (O_3085,N_29010,N_29156);
and UO_3086 (O_3086,N_29316,N_29583);
or UO_3087 (O_3087,N_29915,N_29220);
xor UO_3088 (O_3088,N_29658,N_29902);
or UO_3089 (O_3089,N_29679,N_29383);
nor UO_3090 (O_3090,N_29184,N_29634);
nor UO_3091 (O_3091,N_29196,N_29885);
xor UO_3092 (O_3092,N_29985,N_29451);
nand UO_3093 (O_3093,N_29744,N_29413);
and UO_3094 (O_3094,N_29139,N_29635);
xnor UO_3095 (O_3095,N_29253,N_29891);
nand UO_3096 (O_3096,N_29373,N_29107);
nand UO_3097 (O_3097,N_29837,N_29636);
nand UO_3098 (O_3098,N_29968,N_29774);
or UO_3099 (O_3099,N_29693,N_29552);
xnor UO_3100 (O_3100,N_29270,N_29640);
nor UO_3101 (O_3101,N_29536,N_29613);
and UO_3102 (O_3102,N_29216,N_29378);
nor UO_3103 (O_3103,N_29887,N_29590);
nand UO_3104 (O_3104,N_29803,N_29047);
or UO_3105 (O_3105,N_29854,N_29497);
or UO_3106 (O_3106,N_29660,N_29687);
and UO_3107 (O_3107,N_29618,N_29560);
nor UO_3108 (O_3108,N_29047,N_29350);
or UO_3109 (O_3109,N_29794,N_29360);
nand UO_3110 (O_3110,N_29051,N_29674);
nand UO_3111 (O_3111,N_29439,N_29044);
and UO_3112 (O_3112,N_29055,N_29962);
nor UO_3113 (O_3113,N_29213,N_29157);
xor UO_3114 (O_3114,N_29880,N_29264);
nand UO_3115 (O_3115,N_29586,N_29524);
nand UO_3116 (O_3116,N_29973,N_29280);
xnor UO_3117 (O_3117,N_29906,N_29723);
nor UO_3118 (O_3118,N_29939,N_29991);
nand UO_3119 (O_3119,N_29150,N_29247);
xor UO_3120 (O_3120,N_29658,N_29479);
and UO_3121 (O_3121,N_29940,N_29493);
or UO_3122 (O_3122,N_29746,N_29393);
nand UO_3123 (O_3123,N_29253,N_29535);
or UO_3124 (O_3124,N_29563,N_29550);
or UO_3125 (O_3125,N_29217,N_29560);
xor UO_3126 (O_3126,N_29199,N_29687);
and UO_3127 (O_3127,N_29183,N_29825);
and UO_3128 (O_3128,N_29464,N_29421);
or UO_3129 (O_3129,N_29973,N_29967);
nand UO_3130 (O_3130,N_29056,N_29724);
xor UO_3131 (O_3131,N_29067,N_29531);
xor UO_3132 (O_3132,N_29854,N_29456);
nand UO_3133 (O_3133,N_29075,N_29424);
and UO_3134 (O_3134,N_29355,N_29260);
nor UO_3135 (O_3135,N_29284,N_29177);
or UO_3136 (O_3136,N_29894,N_29499);
or UO_3137 (O_3137,N_29055,N_29820);
nor UO_3138 (O_3138,N_29753,N_29779);
and UO_3139 (O_3139,N_29166,N_29196);
xnor UO_3140 (O_3140,N_29944,N_29961);
and UO_3141 (O_3141,N_29201,N_29646);
nor UO_3142 (O_3142,N_29717,N_29083);
nor UO_3143 (O_3143,N_29069,N_29393);
or UO_3144 (O_3144,N_29496,N_29861);
nor UO_3145 (O_3145,N_29961,N_29842);
xnor UO_3146 (O_3146,N_29709,N_29768);
nand UO_3147 (O_3147,N_29767,N_29156);
or UO_3148 (O_3148,N_29229,N_29533);
nand UO_3149 (O_3149,N_29495,N_29271);
nand UO_3150 (O_3150,N_29936,N_29586);
or UO_3151 (O_3151,N_29991,N_29431);
xor UO_3152 (O_3152,N_29426,N_29306);
nand UO_3153 (O_3153,N_29212,N_29746);
nor UO_3154 (O_3154,N_29579,N_29401);
xnor UO_3155 (O_3155,N_29551,N_29718);
xor UO_3156 (O_3156,N_29841,N_29703);
nor UO_3157 (O_3157,N_29454,N_29362);
nand UO_3158 (O_3158,N_29297,N_29697);
and UO_3159 (O_3159,N_29725,N_29853);
or UO_3160 (O_3160,N_29965,N_29447);
nor UO_3161 (O_3161,N_29162,N_29206);
nor UO_3162 (O_3162,N_29782,N_29602);
nor UO_3163 (O_3163,N_29695,N_29085);
xnor UO_3164 (O_3164,N_29502,N_29666);
and UO_3165 (O_3165,N_29858,N_29026);
nand UO_3166 (O_3166,N_29078,N_29791);
nor UO_3167 (O_3167,N_29949,N_29068);
or UO_3168 (O_3168,N_29846,N_29537);
or UO_3169 (O_3169,N_29747,N_29185);
xor UO_3170 (O_3170,N_29634,N_29171);
xnor UO_3171 (O_3171,N_29133,N_29134);
and UO_3172 (O_3172,N_29611,N_29407);
xnor UO_3173 (O_3173,N_29225,N_29145);
and UO_3174 (O_3174,N_29630,N_29734);
or UO_3175 (O_3175,N_29768,N_29739);
or UO_3176 (O_3176,N_29732,N_29723);
nand UO_3177 (O_3177,N_29077,N_29748);
xnor UO_3178 (O_3178,N_29868,N_29684);
xnor UO_3179 (O_3179,N_29484,N_29864);
and UO_3180 (O_3180,N_29790,N_29991);
nand UO_3181 (O_3181,N_29892,N_29079);
and UO_3182 (O_3182,N_29009,N_29420);
or UO_3183 (O_3183,N_29802,N_29924);
and UO_3184 (O_3184,N_29188,N_29504);
and UO_3185 (O_3185,N_29687,N_29322);
and UO_3186 (O_3186,N_29298,N_29347);
nand UO_3187 (O_3187,N_29763,N_29048);
or UO_3188 (O_3188,N_29398,N_29794);
or UO_3189 (O_3189,N_29822,N_29476);
xnor UO_3190 (O_3190,N_29487,N_29111);
nor UO_3191 (O_3191,N_29952,N_29720);
nor UO_3192 (O_3192,N_29594,N_29274);
xnor UO_3193 (O_3193,N_29569,N_29428);
nand UO_3194 (O_3194,N_29727,N_29340);
or UO_3195 (O_3195,N_29350,N_29345);
nor UO_3196 (O_3196,N_29235,N_29918);
nor UO_3197 (O_3197,N_29169,N_29435);
xor UO_3198 (O_3198,N_29559,N_29483);
and UO_3199 (O_3199,N_29574,N_29102);
nand UO_3200 (O_3200,N_29917,N_29181);
nand UO_3201 (O_3201,N_29210,N_29124);
or UO_3202 (O_3202,N_29783,N_29249);
and UO_3203 (O_3203,N_29732,N_29559);
nand UO_3204 (O_3204,N_29164,N_29978);
or UO_3205 (O_3205,N_29276,N_29190);
or UO_3206 (O_3206,N_29806,N_29113);
and UO_3207 (O_3207,N_29569,N_29508);
nand UO_3208 (O_3208,N_29503,N_29918);
nand UO_3209 (O_3209,N_29636,N_29795);
or UO_3210 (O_3210,N_29816,N_29084);
xor UO_3211 (O_3211,N_29379,N_29748);
nand UO_3212 (O_3212,N_29199,N_29700);
or UO_3213 (O_3213,N_29967,N_29658);
xor UO_3214 (O_3214,N_29187,N_29200);
nor UO_3215 (O_3215,N_29106,N_29775);
and UO_3216 (O_3216,N_29486,N_29214);
nand UO_3217 (O_3217,N_29990,N_29303);
or UO_3218 (O_3218,N_29427,N_29180);
nand UO_3219 (O_3219,N_29356,N_29706);
nand UO_3220 (O_3220,N_29841,N_29554);
xor UO_3221 (O_3221,N_29557,N_29294);
or UO_3222 (O_3222,N_29102,N_29185);
or UO_3223 (O_3223,N_29811,N_29463);
xnor UO_3224 (O_3224,N_29685,N_29036);
nor UO_3225 (O_3225,N_29985,N_29547);
and UO_3226 (O_3226,N_29521,N_29502);
or UO_3227 (O_3227,N_29111,N_29962);
xnor UO_3228 (O_3228,N_29223,N_29227);
or UO_3229 (O_3229,N_29135,N_29088);
xnor UO_3230 (O_3230,N_29602,N_29786);
xor UO_3231 (O_3231,N_29973,N_29188);
and UO_3232 (O_3232,N_29538,N_29558);
xor UO_3233 (O_3233,N_29027,N_29681);
xnor UO_3234 (O_3234,N_29951,N_29796);
xor UO_3235 (O_3235,N_29700,N_29426);
or UO_3236 (O_3236,N_29064,N_29721);
or UO_3237 (O_3237,N_29655,N_29169);
or UO_3238 (O_3238,N_29955,N_29575);
and UO_3239 (O_3239,N_29411,N_29440);
xor UO_3240 (O_3240,N_29957,N_29709);
and UO_3241 (O_3241,N_29779,N_29425);
nor UO_3242 (O_3242,N_29632,N_29854);
nand UO_3243 (O_3243,N_29187,N_29558);
and UO_3244 (O_3244,N_29477,N_29175);
nand UO_3245 (O_3245,N_29456,N_29162);
or UO_3246 (O_3246,N_29669,N_29509);
nor UO_3247 (O_3247,N_29365,N_29665);
xnor UO_3248 (O_3248,N_29741,N_29327);
xnor UO_3249 (O_3249,N_29659,N_29582);
nand UO_3250 (O_3250,N_29835,N_29377);
nand UO_3251 (O_3251,N_29139,N_29432);
xor UO_3252 (O_3252,N_29707,N_29220);
nand UO_3253 (O_3253,N_29743,N_29523);
xor UO_3254 (O_3254,N_29857,N_29199);
or UO_3255 (O_3255,N_29864,N_29519);
and UO_3256 (O_3256,N_29751,N_29493);
nand UO_3257 (O_3257,N_29466,N_29622);
nor UO_3258 (O_3258,N_29945,N_29752);
and UO_3259 (O_3259,N_29303,N_29394);
and UO_3260 (O_3260,N_29406,N_29509);
nor UO_3261 (O_3261,N_29033,N_29462);
nand UO_3262 (O_3262,N_29305,N_29124);
nand UO_3263 (O_3263,N_29057,N_29998);
nand UO_3264 (O_3264,N_29735,N_29629);
nand UO_3265 (O_3265,N_29136,N_29631);
or UO_3266 (O_3266,N_29865,N_29624);
and UO_3267 (O_3267,N_29536,N_29641);
nand UO_3268 (O_3268,N_29782,N_29783);
nand UO_3269 (O_3269,N_29258,N_29713);
and UO_3270 (O_3270,N_29339,N_29950);
nor UO_3271 (O_3271,N_29365,N_29507);
or UO_3272 (O_3272,N_29688,N_29859);
and UO_3273 (O_3273,N_29207,N_29654);
or UO_3274 (O_3274,N_29494,N_29697);
xnor UO_3275 (O_3275,N_29428,N_29931);
xor UO_3276 (O_3276,N_29231,N_29873);
nor UO_3277 (O_3277,N_29711,N_29146);
nor UO_3278 (O_3278,N_29582,N_29056);
and UO_3279 (O_3279,N_29886,N_29496);
nand UO_3280 (O_3280,N_29616,N_29499);
and UO_3281 (O_3281,N_29974,N_29241);
xnor UO_3282 (O_3282,N_29541,N_29454);
or UO_3283 (O_3283,N_29823,N_29948);
nand UO_3284 (O_3284,N_29925,N_29301);
nor UO_3285 (O_3285,N_29735,N_29594);
xnor UO_3286 (O_3286,N_29799,N_29918);
and UO_3287 (O_3287,N_29283,N_29623);
nor UO_3288 (O_3288,N_29419,N_29474);
or UO_3289 (O_3289,N_29222,N_29841);
nand UO_3290 (O_3290,N_29455,N_29736);
or UO_3291 (O_3291,N_29122,N_29395);
nand UO_3292 (O_3292,N_29390,N_29679);
and UO_3293 (O_3293,N_29992,N_29037);
nor UO_3294 (O_3294,N_29885,N_29181);
and UO_3295 (O_3295,N_29709,N_29354);
or UO_3296 (O_3296,N_29182,N_29281);
and UO_3297 (O_3297,N_29917,N_29271);
nor UO_3298 (O_3298,N_29235,N_29960);
nor UO_3299 (O_3299,N_29795,N_29898);
xor UO_3300 (O_3300,N_29664,N_29960);
nand UO_3301 (O_3301,N_29545,N_29335);
nand UO_3302 (O_3302,N_29845,N_29687);
and UO_3303 (O_3303,N_29463,N_29554);
nor UO_3304 (O_3304,N_29936,N_29705);
and UO_3305 (O_3305,N_29574,N_29335);
or UO_3306 (O_3306,N_29741,N_29729);
and UO_3307 (O_3307,N_29563,N_29754);
or UO_3308 (O_3308,N_29223,N_29794);
and UO_3309 (O_3309,N_29406,N_29830);
or UO_3310 (O_3310,N_29510,N_29439);
xor UO_3311 (O_3311,N_29063,N_29038);
nand UO_3312 (O_3312,N_29485,N_29345);
xnor UO_3313 (O_3313,N_29587,N_29513);
and UO_3314 (O_3314,N_29318,N_29244);
nor UO_3315 (O_3315,N_29049,N_29117);
xor UO_3316 (O_3316,N_29562,N_29694);
nand UO_3317 (O_3317,N_29303,N_29727);
xor UO_3318 (O_3318,N_29623,N_29708);
nand UO_3319 (O_3319,N_29305,N_29136);
xnor UO_3320 (O_3320,N_29587,N_29673);
nand UO_3321 (O_3321,N_29450,N_29187);
or UO_3322 (O_3322,N_29136,N_29665);
and UO_3323 (O_3323,N_29447,N_29527);
nor UO_3324 (O_3324,N_29104,N_29996);
and UO_3325 (O_3325,N_29402,N_29426);
or UO_3326 (O_3326,N_29566,N_29167);
or UO_3327 (O_3327,N_29795,N_29299);
xor UO_3328 (O_3328,N_29032,N_29424);
nand UO_3329 (O_3329,N_29938,N_29803);
xnor UO_3330 (O_3330,N_29383,N_29470);
nand UO_3331 (O_3331,N_29130,N_29444);
and UO_3332 (O_3332,N_29822,N_29784);
xnor UO_3333 (O_3333,N_29753,N_29762);
nor UO_3334 (O_3334,N_29330,N_29113);
and UO_3335 (O_3335,N_29122,N_29379);
nand UO_3336 (O_3336,N_29926,N_29388);
nand UO_3337 (O_3337,N_29910,N_29527);
nand UO_3338 (O_3338,N_29533,N_29552);
or UO_3339 (O_3339,N_29341,N_29184);
xor UO_3340 (O_3340,N_29642,N_29354);
nor UO_3341 (O_3341,N_29213,N_29742);
nor UO_3342 (O_3342,N_29875,N_29876);
or UO_3343 (O_3343,N_29039,N_29500);
nor UO_3344 (O_3344,N_29797,N_29658);
nor UO_3345 (O_3345,N_29114,N_29576);
xor UO_3346 (O_3346,N_29470,N_29941);
xor UO_3347 (O_3347,N_29068,N_29119);
and UO_3348 (O_3348,N_29045,N_29520);
nor UO_3349 (O_3349,N_29211,N_29766);
or UO_3350 (O_3350,N_29874,N_29137);
nand UO_3351 (O_3351,N_29513,N_29054);
nand UO_3352 (O_3352,N_29163,N_29753);
nand UO_3353 (O_3353,N_29775,N_29921);
and UO_3354 (O_3354,N_29270,N_29176);
or UO_3355 (O_3355,N_29493,N_29041);
nor UO_3356 (O_3356,N_29629,N_29000);
xnor UO_3357 (O_3357,N_29275,N_29700);
xnor UO_3358 (O_3358,N_29990,N_29146);
and UO_3359 (O_3359,N_29655,N_29838);
or UO_3360 (O_3360,N_29300,N_29994);
or UO_3361 (O_3361,N_29933,N_29300);
or UO_3362 (O_3362,N_29206,N_29042);
nor UO_3363 (O_3363,N_29929,N_29741);
nor UO_3364 (O_3364,N_29212,N_29123);
xnor UO_3365 (O_3365,N_29905,N_29062);
and UO_3366 (O_3366,N_29657,N_29234);
or UO_3367 (O_3367,N_29058,N_29800);
nor UO_3368 (O_3368,N_29077,N_29281);
or UO_3369 (O_3369,N_29504,N_29664);
or UO_3370 (O_3370,N_29274,N_29256);
xor UO_3371 (O_3371,N_29813,N_29223);
or UO_3372 (O_3372,N_29749,N_29690);
and UO_3373 (O_3373,N_29708,N_29819);
nand UO_3374 (O_3374,N_29981,N_29230);
nand UO_3375 (O_3375,N_29078,N_29252);
nand UO_3376 (O_3376,N_29378,N_29679);
or UO_3377 (O_3377,N_29030,N_29596);
nor UO_3378 (O_3378,N_29571,N_29658);
or UO_3379 (O_3379,N_29444,N_29007);
xor UO_3380 (O_3380,N_29800,N_29220);
nor UO_3381 (O_3381,N_29172,N_29756);
nor UO_3382 (O_3382,N_29391,N_29901);
nor UO_3383 (O_3383,N_29774,N_29765);
nor UO_3384 (O_3384,N_29104,N_29401);
or UO_3385 (O_3385,N_29293,N_29662);
or UO_3386 (O_3386,N_29814,N_29010);
xnor UO_3387 (O_3387,N_29401,N_29639);
nor UO_3388 (O_3388,N_29582,N_29560);
or UO_3389 (O_3389,N_29896,N_29871);
nand UO_3390 (O_3390,N_29131,N_29813);
nor UO_3391 (O_3391,N_29130,N_29212);
nor UO_3392 (O_3392,N_29778,N_29012);
nor UO_3393 (O_3393,N_29701,N_29766);
nor UO_3394 (O_3394,N_29896,N_29026);
or UO_3395 (O_3395,N_29512,N_29032);
or UO_3396 (O_3396,N_29566,N_29005);
and UO_3397 (O_3397,N_29199,N_29922);
and UO_3398 (O_3398,N_29562,N_29960);
or UO_3399 (O_3399,N_29720,N_29843);
xnor UO_3400 (O_3400,N_29949,N_29294);
nor UO_3401 (O_3401,N_29417,N_29789);
and UO_3402 (O_3402,N_29167,N_29973);
nand UO_3403 (O_3403,N_29576,N_29895);
nand UO_3404 (O_3404,N_29670,N_29850);
or UO_3405 (O_3405,N_29868,N_29217);
xor UO_3406 (O_3406,N_29180,N_29008);
or UO_3407 (O_3407,N_29233,N_29570);
or UO_3408 (O_3408,N_29614,N_29003);
nor UO_3409 (O_3409,N_29770,N_29689);
nand UO_3410 (O_3410,N_29374,N_29204);
nand UO_3411 (O_3411,N_29986,N_29628);
nand UO_3412 (O_3412,N_29953,N_29402);
xnor UO_3413 (O_3413,N_29348,N_29966);
or UO_3414 (O_3414,N_29450,N_29711);
or UO_3415 (O_3415,N_29868,N_29025);
and UO_3416 (O_3416,N_29273,N_29968);
or UO_3417 (O_3417,N_29411,N_29096);
and UO_3418 (O_3418,N_29796,N_29178);
nor UO_3419 (O_3419,N_29304,N_29530);
and UO_3420 (O_3420,N_29203,N_29251);
nor UO_3421 (O_3421,N_29975,N_29123);
or UO_3422 (O_3422,N_29086,N_29329);
or UO_3423 (O_3423,N_29454,N_29751);
nand UO_3424 (O_3424,N_29389,N_29988);
xnor UO_3425 (O_3425,N_29837,N_29744);
nand UO_3426 (O_3426,N_29837,N_29721);
nor UO_3427 (O_3427,N_29913,N_29580);
or UO_3428 (O_3428,N_29721,N_29727);
nand UO_3429 (O_3429,N_29376,N_29812);
and UO_3430 (O_3430,N_29689,N_29423);
and UO_3431 (O_3431,N_29260,N_29469);
nand UO_3432 (O_3432,N_29451,N_29172);
nand UO_3433 (O_3433,N_29939,N_29002);
nand UO_3434 (O_3434,N_29595,N_29006);
and UO_3435 (O_3435,N_29934,N_29338);
nand UO_3436 (O_3436,N_29804,N_29213);
and UO_3437 (O_3437,N_29179,N_29478);
xnor UO_3438 (O_3438,N_29731,N_29431);
xnor UO_3439 (O_3439,N_29659,N_29932);
nor UO_3440 (O_3440,N_29014,N_29358);
and UO_3441 (O_3441,N_29137,N_29937);
nor UO_3442 (O_3442,N_29496,N_29480);
or UO_3443 (O_3443,N_29400,N_29712);
nand UO_3444 (O_3444,N_29622,N_29309);
xor UO_3445 (O_3445,N_29068,N_29518);
or UO_3446 (O_3446,N_29667,N_29965);
or UO_3447 (O_3447,N_29732,N_29815);
nor UO_3448 (O_3448,N_29426,N_29339);
xor UO_3449 (O_3449,N_29260,N_29082);
xnor UO_3450 (O_3450,N_29666,N_29835);
nand UO_3451 (O_3451,N_29684,N_29564);
xor UO_3452 (O_3452,N_29750,N_29162);
nand UO_3453 (O_3453,N_29470,N_29375);
nand UO_3454 (O_3454,N_29890,N_29540);
and UO_3455 (O_3455,N_29689,N_29771);
and UO_3456 (O_3456,N_29148,N_29423);
xor UO_3457 (O_3457,N_29881,N_29410);
nand UO_3458 (O_3458,N_29121,N_29833);
nor UO_3459 (O_3459,N_29548,N_29616);
or UO_3460 (O_3460,N_29098,N_29204);
or UO_3461 (O_3461,N_29244,N_29885);
and UO_3462 (O_3462,N_29687,N_29151);
nand UO_3463 (O_3463,N_29553,N_29254);
nand UO_3464 (O_3464,N_29453,N_29796);
nor UO_3465 (O_3465,N_29574,N_29141);
xor UO_3466 (O_3466,N_29141,N_29740);
nor UO_3467 (O_3467,N_29204,N_29405);
and UO_3468 (O_3468,N_29215,N_29639);
nand UO_3469 (O_3469,N_29998,N_29257);
xnor UO_3470 (O_3470,N_29647,N_29256);
and UO_3471 (O_3471,N_29710,N_29948);
or UO_3472 (O_3472,N_29516,N_29348);
xor UO_3473 (O_3473,N_29151,N_29335);
or UO_3474 (O_3474,N_29469,N_29204);
nand UO_3475 (O_3475,N_29297,N_29782);
or UO_3476 (O_3476,N_29008,N_29319);
or UO_3477 (O_3477,N_29207,N_29453);
and UO_3478 (O_3478,N_29610,N_29830);
or UO_3479 (O_3479,N_29633,N_29745);
and UO_3480 (O_3480,N_29022,N_29668);
nor UO_3481 (O_3481,N_29454,N_29034);
and UO_3482 (O_3482,N_29723,N_29509);
nand UO_3483 (O_3483,N_29257,N_29546);
and UO_3484 (O_3484,N_29325,N_29269);
nand UO_3485 (O_3485,N_29772,N_29626);
and UO_3486 (O_3486,N_29990,N_29054);
xnor UO_3487 (O_3487,N_29481,N_29392);
xnor UO_3488 (O_3488,N_29520,N_29515);
nand UO_3489 (O_3489,N_29292,N_29839);
xor UO_3490 (O_3490,N_29337,N_29420);
xor UO_3491 (O_3491,N_29957,N_29671);
nor UO_3492 (O_3492,N_29034,N_29057);
or UO_3493 (O_3493,N_29348,N_29049);
or UO_3494 (O_3494,N_29672,N_29008);
nand UO_3495 (O_3495,N_29227,N_29975);
or UO_3496 (O_3496,N_29884,N_29976);
or UO_3497 (O_3497,N_29984,N_29860);
and UO_3498 (O_3498,N_29033,N_29891);
nand UO_3499 (O_3499,N_29872,N_29085);
endmodule