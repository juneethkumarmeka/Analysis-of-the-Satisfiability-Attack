module basic_1000_10000_1500_4_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_152,In_808);
or U1 (N_1,In_549,In_560);
and U2 (N_2,In_624,In_155);
nand U3 (N_3,In_853,In_695);
and U4 (N_4,In_211,In_645);
nor U5 (N_5,In_438,In_82);
nor U6 (N_6,In_567,In_589);
or U7 (N_7,In_237,In_218);
and U8 (N_8,In_283,In_395);
nor U9 (N_9,In_970,In_71);
and U10 (N_10,In_277,In_382);
nand U11 (N_11,In_790,In_122);
nand U12 (N_12,In_904,In_553);
and U13 (N_13,In_272,In_592);
nand U14 (N_14,In_230,In_56);
nor U15 (N_15,In_255,In_956);
and U16 (N_16,In_239,In_366);
or U17 (N_17,In_169,In_207);
nand U18 (N_18,In_313,In_47);
nor U19 (N_19,In_146,In_259);
or U20 (N_20,In_17,In_727);
and U21 (N_21,In_343,In_284);
nor U22 (N_22,In_603,In_620);
or U23 (N_23,In_988,In_951);
and U24 (N_24,In_583,In_104);
and U25 (N_25,In_637,In_662);
nand U26 (N_26,In_550,In_745);
nor U27 (N_27,In_643,In_200);
nand U28 (N_28,In_209,In_714);
nor U29 (N_29,In_423,In_163);
and U30 (N_30,In_716,In_445);
nor U31 (N_31,In_717,In_947);
nand U32 (N_32,In_139,In_723);
xor U33 (N_33,In_866,In_124);
and U34 (N_34,In_764,In_945);
nor U35 (N_35,In_447,In_81);
or U36 (N_36,In_985,In_983);
xor U37 (N_37,In_276,In_667);
nor U38 (N_38,In_960,In_969);
nor U39 (N_39,In_450,In_765);
xor U40 (N_40,In_208,In_523);
or U41 (N_41,In_850,In_776);
xnor U42 (N_42,In_958,In_663);
or U43 (N_43,In_793,In_678);
and U44 (N_44,In_650,In_436);
or U45 (N_45,In_49,In_646);
nand U46 (N_46,In_556,In_883);
nand U47 (N_47,In_180,In_261);
and U48 (N_48,In_310,In_368);
xnor U49 (N_49,In_734,In_340);
nand U50 (N_50,In_720,In_761);
nor U51 (N_51,In_575,In_164);
and U52 (N_52,In_303,In_409);
nor U53 (N_53,In_400,In_529);
or U54 (N_54,In_235,In_434);
and U55 (N_55,In_309,In_151);
xnor U56 (N_56,In_360,In_747);
nor U57 (N_57,In_333,In_769);
and U58 (N_58,In_145,In_711);
nand U59 (N_59,In_666,In_741);
xnor U60 (N_60,In_240,In_348);
and U61 (N_61,In_574,In_927);
or U62 (N_62,In_779,In_617);
nor U63 (N_63,In_119,In_763);
nor U64 (N_64,In_675,In_568);
or U65 (N_65,In_472,In_886);
nor U66 (N_66,In_202,In_314);
nand U67 (N_67,In_319,In_470);
or U68 (N_68,In_127,In_700);
and U69 (N_69,In_330,In_561);
or U70 (N_70,In_888,In_521);
and U71 (N_71,In_821,In_564);
nor U72 (N_72,In_681,In_785);
or U73 (N_73,In_852,In_851);
and U74 (N_74,In_913,In_759);
or U75 (N_75,In_223,In_690);
nor U76 (N_76,In_531,In_535);
xnor U77 (N_77,In_471,In_842);
nand U78 (N_78,In_329,In_459);
nand U79 (N_79,In_994,In_915);
or U80 (N_80,In_267,In_751);
and U81 (N_81,In_347,In_772);
nand U82 (N_82,In_632,In_972);
and U83 (N_83,In_386,In_285);
xor U84 (N_84,In_385,In_599);
or U85 (N_85,In_115,In_909);
nor U86 (N_86,In_50,In_647);
nor U87 (N_87,In_376,In_993);
nand U88 (N_88,In_424,In_140);
or U89 (N_89,In_537,In_840);
and U90 (N_90,In_444,In_244);
nor U91 (N_91,In_522,In_42);
nor U92 (N_92,In_26,In_844);
nor U93 (N_93,In_510,In_220);
nor U94 (N_94,In_57,In_879);
nor U95 (N_95,In_439,In_45);
nor U96 (N_96,In_62,In_925);
nand U97 (N_97,In_755,In_88);
and U98 (N_98,In_818,In_167);
nor U99 (N_99,In_482,In_615);
nand U100 (N_100,In_105,In_388);
nor U101 (N_101,In_486,In_750);
xor U102 (N_102,In_0,In_379);
or U103 (N_103,In_500,In_190);
xnor U104 (N_104,In_106,In_23);
nor U105 (N_105,In_724,In_664);
nand U106 (N_106,In_495,In_296);
nor U107 (N_107,In_53,In_318);
and U108 (N_108,In_874,In_926);
or U109 (N_109,In_614,In_829);
nand U110 (N_110,In_843,In_804);
and U111 (N_111,In_813,In_532);
xor U112 (N_112,In_483,In_756);
or U113 (N_113,In_350,In_412);
xnor U114 (N_114,In_541,In_777);
xor U115 (N_115,In_422,In_515);
nand U116 (N_116,In_378,In_394);
nand U117 (N_117,In_460,In_30);
or U118 (N_118,In_584,In_77);
or U119 (N_119,In_875,In_217);
nand U120 (N_120,In_810,In_89);
nor U121 (N_121,In_786,In_782);
and U122 (N_122,In_100,In_501);
nor U123 (N_123,In_511,In_487);
and U124 (N_124,In_744,In_430);
or U125 (N_125,In_507,In_757);
or U126 (N_126,In_280,In_701);
nand U127 (N_127,In_526,In_22);
nor U128 (N_128,In_943,In_948);
nor U129 (N_129,In_257,In_128);
nor U130 (N_130,In_801,In_950);
and U131 (N_131,In_578,In_335);
nand U132 (N_132,In_628,In_192);
and U133 (N_133,In_939,In_626);
or U134 (N_134,In_469,In_743);
and U135 (N_135,In_232,In_655);
nand U136 (N_136,In_107,In_33);
or U137 (N_137,In_260,In_233);
or U138 (N_138,In_282,In_706);
nand U139 (N_139,In_936,In_796);
and U140 (N_140,In_389,In_393);
or U141 (N_141,In_225,In_691);
or U142 (N_142,In_456,In_18);
and U143 (N_143,In_497,In_981);
nand U144 (N_144,In_536,In_832);
nand U145 (N_145,In_867,In_35);
or U146 (N_146,In_421,In_496);
nand U147 (N_147,In_109,In_868);
nand U148 (N_148,In_344,In_451);
nand U149 (N_149,In_76,In_827);
or U150 (N_150,In_10,In_427);
or U151 (N_151,In_58,In_885);
nor U152 (N_152,In_353,In_685);
xor U153 (N_153,In_307,In_594);
nor U154 (N_154,In_798,In_40);
nor U155 (N_155,In_437,In_41);
nand U156 (N_156,In_907,In_593);
or U157 (N_157,In_227,In_823);
or U158 (N_158,In_351,In_381);
and U159 (N_159,In_485,In_363);
or U160 (N_160,In_383,In_884);
and U161 (N_161,In_836,In_954);
and U162 (N_162,In_141,In_214);
or U163 (N_163,In_229,In_248);
and U164 (N_164,In_934,In_498);
or U165 (N_165,In_730,In_815);
or U166 (N_166,In_302,In_175);
nor U167 (N_167,In_203,In_586);
and U168 (N_168,In_858,In_513);
xor U169 (N_169,In_998,In_14);
or U170 (N_170,In_838,In_228);
and U171 (N_171,In_289,In_95);
and U172 (N_172,In_660,In_238);
and U173 (N_173,In_547,In_941);
nand U174 (N_174,In_820,In_847);
and U175 (N_175,In_554,In_508);
nor U176 (N_176,In_509,In_9);
nor U177 (N_177,In_373,In_653);
nor U178 (N_178,In_197,In_295);
nand U179 (N_179,In_299,In_652);
and U180 (N_180,In_899,In_922);
nor U181 (N_181,In_93,In_384);
nand U182 (N_182,In_396,In_754);
nand U183 (N_183,In_631,In_737);
and U184 (N_184,In_43,In_429);
xor U185 (N_185,In_961,In_73);
and U186 (N_186,In_391,In_12);
or U187 (N_187,In_189,In_625);
or U188 (N_188,In_872,In_775);
nor U189 (N_189,In_463,In_387);
and U190 (N_190,In_931,In_986);
or U191 (N_191,In_708,In_725);
and U192 (N_192,In_719,In_516);
and U193 (N_193,In_489,In_742);
or U194 (N_194,In_494,In_935);
or U195 (N_195,In_921,In_640);
xnor U196 (N_196,In_11,In_317);
and U197 (N_197,In_336,In_738);
or U198 (N_198,In_890,In_69);
nor U199 (N_199,In_216,In_3);
xnor U200 (N_200,In_736,In_147);
or U201 (N_201,In_659,In_466);
xnor U202 (N_202,In_590,In_403);
nand U203 (N_203,In_413,In_349);
and U204 (N_204,In_903,In_657);
and U205 (N_205,In_540,In_817);
and U206 (N_206,In_432,In_612);
and U207 (N_207,In_362,In_99);
nor U208 (N_208,In_895,In_372);
and U209 (N_209,In_20,In_34);
or U210 (N_210,In_377,In_746);
nor U211 (N_211,In_355,In_601);
nor U212 (N_212,In_36,In_894);
xor U213 (N_213,In_91,In_656);
xnor U214 (N_214,In_420,In_1);
or U215 (N_215,In_671,In_468);
xnor U216 (N_216,In_577,In_324);
nor U217 (N_217,In_305,In_552);
or U218 (N_218,In_773,In_67);
and U219 (N_219,In_64,In_856);
or U220 (N_220,In_609,In_582);
xnor U221 (N_221,In_103,In_365);
or U222 (N_222,In_183,In_807);
nor U223 (N_223,In_722,In_406);
or U224 (N_224,In_178,In_900);
nand U225 (N_225,In_997,In_264);
and U226 (N_226,In_967,In_286);
and U227 (N_227,In_576,In_992);
and U228 (N_228,In_311,In_514);
or U229 (N_229,In_987,In_544);
nor U230 (N_230,In_416,In_811);
nor U231 (N_231,In_8,In_37);
nor U232 (N_232,In_731,In_672);
nor U233 (N_233,In_542,In_845);
or U234 (N_234,In_467,In_144);
nor U235 (N_235,In_783,In_153);
or U236 (N_236,In_132,In_749);
or U237 (N_237,In_221,In_946);
nor U238 (N_238,In_753,In_607);
nor U239 (N_239,In_517,In_157);
nor U240 (N_240,In_705,In_458);
and U241 (N_241,In_633,In_713);
nand U242 (N_242,In_364,In_125);
or U243 (N_243,In_390,In_59);
nor U244 (N_244,In_431,In_996);
nor U245 (N_245,In_787,In_559);
nand U246 (N_246,In_610,In_917);
or U247 (N_247,In_881,In_892);
or U248 (N_248,In_877,In_805);
or U249 (N_249,In_327,In_195);
nand U250 (N_250,In_54,In_579);
nor U251 (N_251,In_789,In_462);
nor U252 (N_252,In_359,In_294);
nor U253 (N_253,In_848,In_154);
nand U254 (N_254,In_627,In_619);
xor U255 (N_255,In_704,In_959);
nor U256 (N_256,In_25,In_480);
or U257 (N_257,In_279,In_506);
nor U258 (N_258,In_933,In_520);
xnor U259 (N_259,In_512,In_802);
nor U260 (N_260,In_504,In_253);
or U261 (N_261,In_715,In_331);
xnor U262 (N_262,In_369,In_611);
or U263 (N_263,In_748,In_457);
and U264 (N_264,In_962,In_712);
or U265 (N_265,In_108,In_942);
or U266 (N_266,In_545,In_938);
and U267 (N_267,In_346,In_999);
and U268 (N_268,In_557,In_762);
nand U269 (N_269,In_898,In_126);
nand U270 (N_270,In_964,In_308);
and U271 (N_271,In_910,In_179);
nand U272 (N_272,In_29,In_519);
and U273 (N_273,In_825,In_358);
nand U274 (N_274,In_803,In_839);
xnor U275 (N_275,In_121,In_380);
xor U276 (N_276,In_709,In_806);
nor U277 (N_277,In_905,In_860);
nor U278 (N_278,In_116,In_873);
and U279 (N_279,In_953,In_172);
and U280 (N_280,In_61,In_689);
nor U281 (N_281,In_158,In_301);
nor U282 (N_282,In_912,In_944);
nor U283 (N_283,In_306,In_809);
and U284 (N_284,In_957,In_326);
nor U285 (N_285,In_13,In_266);
nand U286 (N_286,In_316,In_923);
nand U287 (N_287,In_137,In_928);
xnor U288 (N_288,In_930,In_732);
nor U289 (N_289,In_995,In_916);
or U290 (N_290,In_702,In_694);
nand U291 (N_291,In_680,In_826);
nor U292 (N_292,In_84,In_674);
nor U293 (N_293,In_581,In_974);
xnor U294 (N_294,In_435,In_97);
nand U295 (N_295,In_79,In_236);
nand U296 (N_296,In_204,In_402);
nand U297 (N_297,In_919,In_19);
and U298 (N_298,In_914,In_258);
nand U299 (N_299,In_415,In_452);
and U300 (N_300,In_661,In_528);
and U301 (N_301,In_461,In_191);
nand U302 (N_302,In_142,In_975);
and U303 (N_303,In_841,In_210);
nor U304 (N_304,In_133,In_677);
or U305 (N_305,In_613,In_48);
and U306 (N_306,In_977,In_479);
nand U307 (N_307,In_555,In_268);
nand U308 (N_308,In_605,In_558);
or U309 (N_309,In_7,In_275);
or U310 (N_310,In_426,In_397);
nor U311 (N_311,In_683,In_530);
xnor U312 (N_312,In_352,In_658);
and U313 (N_313,In_597,In_863);
and U314 (N_314,In_6,In_673);
nor U315 (N_315,In_835,In_924);
or U316 (N_316,In_337,In_699);
nand U317 (N_317,In_641,In_679);
and U318 (N_318,In_265,In_138);
xnor U319 (N_319,In_794,In_102);
nor U320 (N_320,In_830,In_991);
or U321 (N_321,In_322,In_940);
nand U322 (N_322,In_184,In_134);
or U323 (N_323,In_159,In_566);
and U324 (N_324,In_323,In_224);
and U325 (N_325,In_897,In_166);
or U326 (N_326,In_46,In_870);
or U327 (N_327,In_623,In_143);
xor U328 (N_328,In_425,In_668);
or U329 (N_329,In_399,In_70);
or U330 (N_330,In_342,In_973);
and U331 (N_331,In_325,In_38);
xor U332 (N_332,In_630,In_251);
and U333 (N_333,In_182,In_474);
nor U334 (N_334,In_570,In_602);
nand U335 (N_335,In_367,In_478);
or U336 (N_336,In_493,In_173);
nand U337 (N_337,In_864,In_505);
nand U338 (N_338,In_833,In_822);
nor U339 (N_339,In_814,In_320);
nor U340 (N_340,In_252,In_168);
nor U341 (N_341,In_123,In_865);
nand U342 (N_342,In_649,In_644);
or U343 (N_343,In_792,In_538);
xnor U344 (N_344,In_414,In_697);
and U345 (N_345,In_816,In_984);
or U346 (N_346,In_354,In_51);
or U347 (N_347,In_788,In_148);
nor U348 (N_348,In_475,In_539);
nor U349 (N_349,In_441,In_85);
and U350 (N_350,In_533,In_408);
nand U351 (N_351,In_569,In_334);
and U352 (N_352,In_846,In_728);
nand U353 (N_353,In_600,In_118);
or U354 (N_354,In_932,In_407);
and U355 (N_355,In_911,In_112);
or U356 (N_356,In_418,In_87);
and U357 (N_357,In_966,In_871);
nor U358 (N_358,In_449,In_375);
nor U359 (N_359,In_55,In_618);
or U360 (N_360,In_591,In_129);
or U361 (N_361,In_370,In_758);
nor U362 (N_362,In_799,In_249);
nor U363 (N_363,In_193,In_24);
xor U364 (N_364,In_698,In_187);
or U365 (N_365,In_242,In_186);
nand U366 (N_366,In_32,In_965);
and U367 (N_367,In_206,In_404);
or U368 (N_368,In_740,In_332);
nand U369 (N_369,In_636,In_524);
nor U370 (N_370,In_819,In_733);
nor U371 (N_371,In_194,In_831);
and U372 (N_372,In_250,In_448);
or U373 (N_373,In_688,In_862);
nor U374 (N_374,In_31,In_428);
nand U375 (N_375,In_901,In_15);
nor U376 (N_376,In_80,In_442);
nand U377 (N_377,In_241,In_149);
and U378 (N_378,In_196,In_185);
and U379 (N_379,In_114,In_484);
and U380 (N_380,In_735,In_135);
and U381 (N_381,In_648,In_968);
or U382 (N_382,In_629,In_634);
nand U383 (N_383,In_726,In_784);
or U384 (N_384,In_896,In_411);
or U385 (N_385,In_767,In_491);
nor U386 (N_386,In_345,In_979);
or U387 (N_387,In_682,In_580);
nand U388 (N_388,In_488,In_571);
or U389 (N_389,In_291,In_120);
or U390 (N_390,In_243,In_551);
nand U391 (N_391,In_595,In_72);
xor U392 (N_392,In_502,In_174);
xor U393 (N_393,In_476,In_297);
or U394 (N_394,In_176,In_693);
xor U395 (N_395,In_60,In_791);
or U396 (N_396,In_780,In_608);
nand U397 (N_397,In_490,In_274);
nand U398 (N_398,In_949,In_642);
nand U399 (N_399,In_918,In_982);
nand U400 (N_400,In_28,In_440);
nor U401 (N_401,In_63,In_21);
nand U402 (N_402,In_906,In_66);
and U403 (N_403,In_392,In_638);
or U404 (N_404,In_254,In_978);
nand U405 (N_405,In_215,In_859);
nand U406 (N_406,In_181,In_684);
nand U407 (N_407,In_161,In_718);
and U408 (N_408,In_889,In_869);
xnor U409 (N_409,In_281,In_587);
nand U410 (N_410,In_341,In_247);
nor U411 (N_411,In_16,In_878);
nor U412 (N_412,In_621,In_205);
nand U413 (N_413,In_170,In_721);
and U414 (N_414,In_339,In_929);
or U415 (N_415,In_882,In_503);
nor U416 (N_416,In_278,In_293);
nand U417 (N_417,In_908,In_855);
and U418 (N_418,In_271,In_198);
xnor U419 (N_419,In_263,In_766);
nand U420 (N_420,In_477,In_357);
xnor U421 (N_421,In_96,In_920);
nand U422 (N_422,In_563,In_131);
nor U423 (N_423,In_687,In_952);
nand U424 (N_424,In_876,In_980);
xnor U425 (N_425,In_446,In_219);
nand U426 (N_426,In_92,In_857);
or U427 (N_427,In_596,In_771);
nand U428 (N_428,In_880,In_136);
nor U429 (N_429,In_703,In_269);
or U430 (N_430,In_113,In_887);
nor U431 (N_431,In_499,In_111);
xor U432 (N_432,In_246,In_616);
and U433 (N_433,In_465,In_94);
and U434 (N_434,In_562,In_543);
nor U435 (N_435,In_622,In_83);
nor U436 (N_436,In_891,In_676);
or U437 (N_437,In_824,In_963);
and U438 (N_438,In_971,In_78);
nand U439 (N_439,In_902,In_356);
nor U440 (N_440,In_739,In_234);
nor U441 (N_441,In_797,In_328);
xor U442 (N_442,In_419,In_101);
or U443 (N_443,In_226,In_565);
and U444 (N_444,In_433,In_692);
nand U445 (N_445,In_453,In_262);
or U446 (N_446,In_165,In_492);
nor U447 (N_447,In_774,In_321);
nor U448 (N_448,In_710,In_795);
and U449 (N_449,In_443,In_270);
or U450 (N_450,In_231,In_598);
or U451 (N_451,In_604,In_273);
or U452 (N_452,In_5,In_288);
nand U453 (N_453,In_162,In_473);
nand U454 (N_454,In_989,In_90);
and U455 (N_455,In_188,In_686);
nand U456 (N_456,In_781,In_525);
nor U457 (N_457,In_707,In_150);
or U458 (N_458,In_527,In_778);
and U459 (N_459,In_606,In_405);
and U460 (N_460,In_976,In_39);
nand U461 (N_461,In_752,In_548);
xor U462 (N_462,In_893,In_245);
nand U463 (N_463,In_464,In_156);
nand U464 (N_464,In_199,In_770);
and U465 (N_465,In_670,In_834);
or U466 (N_466,In_481,In_374);
nor U467 (N_467,In_417,In_201);
nand U468 (N_468,In_410,In_828);
and U469 (N_469,In_222,In_177);
nand U470 (N_470,In_256,In_2);
or U471 (N_471,In_635,In_315);
xnor U472 (N_472,In_290,In_729);
nor U473 (N_473,In_654,In_572);
or U474 (N_474,In_573,In_454);
or U475 (N_475,In_455,In_371);
nand U476 (N_476,In_849,In_955);
and U477 (N_477,In_86,In_651);
nand U478 (N_478,In_665,In_27);
xnor U479 (N_479,In_768,In_300);
and U480 (N_480,In_338,In_401);
and U481 (N_481,In_854,In_398);
nand U482 (N_482,In_361,In_130);
nand U483 (N_483,In_760,In_44);
nor U484 (N_484,In_98,In_546);
and U485 (N_485,In_160,In_534);
nor U486 (N_486,In_292,In_696);
xnor U487 (N_487,In_117,In_4);
or U488 (N_488,In_68,In_312);
nand U489 (N_489,In_65,In_585);
and U490 (N_490,In_171,In_990);
nand U491 (N_491,In_800,In_937);
nand U492 (N_492,In_52,In_837);
nand U493 (N_493,In_669,In_812);
nor U494 (N_494,In_287,In_304);
xor U495 (N_495,In_75,In_74);
nand U496 (N_496,In_639,In_588);
xor U497 (N_497,In_518,In_212);
nand U498 (N_498,In_298,In_110);
nor U499 (N_499,In_213,In_861);
and U500 (N_500,In_314,In_944);
nor U501 (N_501,In_769,In_518);
nor U502 (N_502,In_284,In_644);
xor U503 (N_503,In_754,In_663);
xor U504 (N_504,In_95,In_430);
and U505 (N_505,In_810,In_99);
nor U506 (N_506,In_388,In_104);
nand U507 (N_507,In_47,In_882);
and U508 (N_508,In_965,In_365);
nor U509 (N_509,In_205,In_276);
nor U510 (N_510,In_713,In_152);
or U511 (N_511,In_936,In_587);
or U512 (N_512,In_91,In_424);
xnor U513 (N_513,In_170,In_266);
nand U514 (N_514,In_343,In_181);
xnor U515 (N_515,In_533,In_5);
and U516 (N_516,In_216,In_249);
and U517 (N_517,In_863,In_622);
xor U518 (N_518,In_441,In_903);
nand U519 (N_519,In_208,In_151);
nor U520 (N_520,In_820,In_592);
nor U521 (N_521,In_296,In_683);
xnor U522 (N_522,In_688,In_427);
and U523 (N_523,In_312,In_34);
and U524 (N_524,In_660,In_528);
xor U525 (N_525,In_806,In_399);
xor U526 (N_526,In_550,In_548);
nand U527 (N_527,In_475,In_135);
nand U528 (N_528,In_343,In_719);
xnor U529 (N_529,In_747,In_542);
xor U530 (N_530,In_686,In_623);
nor U531 (N_531,In_148,In_536);
and U532 (N_532,In_343,In_604);
nand U533 (N_533,In_559,In_550);
nor U534 (N_534,In_962,In_620);
or U535 (N_535,In_118,In_642);
or U536 (N_536,In_367,In_497);
nor U537 (N_537,In_486,In_409);
nand U538 (N_538,In_396,In_939);
nor U539 (N_539,In_416,In_683);
and U540 (N_540,In_140,In_889);
nand U541 (N_541,In_94,In_428);
or U542 (N_542,In_615,In_926);
nor U543 (N_543,In_537,In_587);
or U544 (N_544,In_867,In_584);
nand U545 (N_545,In_661,In_374);
and U546 (N_546,In_713,In_485);
and U547 (N_547,In_934,In_891);
and U548 (N_548,In_425,In_636);
nor U549 (N_549,In_290,In_296);
and U550 (N_550,In_407,In_242);
nand U551 (N_551,In_843,In_831);
and U552 (N_552,In_801,In_538);
and U553 (N_553,In_8,In_404);
or U554 (N_554,In_773,In_989);
and U555 (N_555,In_129,In_292);
and U556 (N_556,In_680,In_958);
nand U557 (N_557,In_259,In_909);
nand U558 (N_558,In_778,In_491);
and U559 (N_559,In_635,In_694);
xnor U560 (N_560,In_916,In_466);
xnor U561 (N_561,In_527,In_65);
nor U562 (N_562,In_993,In_936);
nand U563 (N_563,In_802,In_63);
xnor U564 (N_564,In_266,In_590);
nor U565 (N_565,In_997,In_700);
nand U566 (N_566,In_849,In_523);
or U567 (N_567,In_85,In_955);
nand U568 (N_568,In_290,In_517);
nand U569 (N_569,In_396,In_656);
nand U570 (N_570,In_646,In_501);
or U571 (N_571,In_307,In_624);
nor U572 (N_572,In_446,In_764);
nand U573 (N_573,In_189,In_52);
and U574 (N_574,In_906,In_733);
and U575 (N_575,In_372,In_676);
and U576 (N_576,In_666,In_63);
and U577 (N_577,In_280,In_257);
nand U578 (N_578,In_19,In_325);
nand U579 (N_579,In_45,In_855);
nor U580 (N_580,In_543,In_942);
nor U581 (N_581,In_650,In_513);
nand U582 (N_582,In_685,In_772);
or U583 (N_583,In_159,In_98);
or U584 (N_584,In_919,In_928);
nor U585 (N_585,In_521,In_210);
and U586 (N_586,In_27,In_404);
or U587 (N_587,In_897,In_378);
nand U588 (N_588,In_460,In_631);
nand U589 (N_589,In_327,In_638);
nand U590 (N_590,In_989,In_934);
nand U591 (N_591,In_281,In_147);
and U592 (N_592,In_872,In_101);
nand U593 (N_593,In_396,In_548);
nand U594 (N_594,In_575,In_186);
nand U595 (N_595,In_711,In_760);
or U596 (N_596,In_28,In_722);
or U597 (N_597,In_524,In_541);
nand U598 (N_598,In_987,In_554);
nor U599 (N_599,In_666,In_92);
nand U600 (N_600,In_981,In_475);
nor U601 (N_601,In_657,In_315);
xor U602 (N_602,In_657,In_217);
xor U603 (N_603,In_618,In_931);
xor U604 (N_604,In_320,In_703);
nor U605 (N_605,In_819,In_664);
or U606 (N_606,In_471,In_301);
nand U607 (N_607,In_545,In_270);
and U608 (N_608,In_959,In_510);
nand U609 (N_609,In_615,In_829);
and U610 (N_610,In_301,In_455);
xnor U611 (N_611,In_924,In_72);
and U612 (N_612,In_270,In_154);
nor U613 (N_613,In_153,In_769);
and U614 (N_614,In_228,In_140);
nand U615 (N_615,In_895,In_589);
and U616 (N_616,In_705,In_998);
nor U617 (N_617,In_355,In_464);
nand U618 (N_618,In_3,In_356);
nand U619 (N_619,In_343,In_990);
nand U620 (N_620,In_523,In_351);
xnor U621 (N_621,In_185,In_182);
or U622 (N_622,In_848,In_293);
and U623 (N_623,In_638,In_192);
and U624 (N_624,In_759,In_140);
and U625 (N_625,In_294,In_344);
nor U626 (N_626,In_291,In_522);
and U627 (N_627,In_353,In_85);
nand U628 (N_628,In_576,In_677);
or U629 (N_629,In_163,In_299);
or U630 (N_630,In_635,In_669);
or U631 (N_631,In_474,In_967);
or U632 (N_632,In_92,In_671);
nand U633 (N_633,In_659,In_141);
nand U634 (N_634,In_479,In_35);
nor U635 (N_635,In_680,In_140);
or U636 (N_636,In_529,In_721);
and U637 (N_637,In_236,In_177);
xnor U638 (N_638,In_27,In_198);
nor U639 (N_639,In_253,In_36);
nand U640 (N_640,In_659,In_839);
and U641 (N_641,In_623,In_98);
and U642 (N_642,In_232,In_128);
nor U643 (N_643,In_12,In_775);
xnor U644 (N_644,In_908,In_430);
nand U645 (N_645,In_931,In_951);
or U646 (N_646,In_397,In_610);
and U647 (N_647,In_531,In_907);
nand U648 (N_648,In_763,In_36);
and U649 (N_649,In_413,In_672);
nand U650 (N_650,In_38,In_587);
and U651 (N_651,In_330,In_688);
and U652 (N_652,In_717,In_732);
or U653 (N_653,In_51,In_559);
nand U654 (N_654,In_574,In_593);
or U655 (N_655,In_717,In_692);
nor U656 (N_656,In_443,In_102);
nand U657 (N_657,In_681,In_181);
or U658 (N_658,In_291,In_633);
nor U659 (N_659,In_179,In_733);
and U660 (N_660,In_473,In_387);
and U661 (N_661,In_197,In_328);
nand U662 (N_662,In_392,In_433);
xnor U663 (N_663,In_940,In_241);
nand U664 (N_664,In_196,In_56);
or U665 (N_665,In_786,In_392);
nand U666 (N_666,In_140,In_826);
nor U667 (N_667,In_136,In_545);
or U668 (N_668,In_691,In_169);
nor U669 (N_669,In_768,In_472);
or U670 (N_670,In_119,In_463);
or U671 (N_671,In_814,In_508);
or U672 (N_672,In_475,In_561);
nor U673 (N_673,In_675,In_817);
nor U674 (N_674,In_407,In_870);
nand U675 (N_675,In_158,In_680);
nor U676 (N_676,In_14,In_963);
and U677 (N_677,In_249,In_792);
and U678 (N_678,In_899,In_32);
and U679 (N_679,In_511,In_751);
and U680 (N_680,In_867,In_612);
or U681 (N_681,In_444,In_646);
nand U682 (N_682,In_716,In_427);
and U683 (N_683,In_244,In_471);
or U684 (N_684,In_965,In_199);
or U685 (N_685,In_902,In_447);
and U686 (N_686,In_296,In_259);
nor U687 (N_687,In_4,In_174);
nor U688 (N_688,In_703,In_53);
nand U689 (N_689,In_772,In_933);
nand U690 (N_690,In_129,In_58);
nor U691 (N_691,In_592,In_340);
nand U692 (N_692,In_511,In_539);
nor U693 (N_693,In_331,In_731);
or U694 (N_694,In_560,In_41);
nand U695 (N_695,In_212,In_838);
or U696 (N_696,In_781,In_506);
or U697 (N_697,In_781,In_520);
and U698 (N_698,In_861,In_763);
or U699 (N_699,In_334,In_527);
xnor U700 (N_700,In_694,In_601);
nor U701 (N_701,In_674,In_774);
nand U702 (N_702,In_917,In_45);
and U703 (N_703,In_891,In_666);
or U704 (N_704,In_622,In_205);
nor U705 (N_705,In_15,In_221);
xor U706 (N_706,In_753,In_913);
nand U707 (N_707,In_187,In_578);
nor U708 (N_708,In_349,In_968);
nand U709 (N_709,In_534,In_149);
or U710 (N_710,In_982,In_648);
and U711 (N_711,In_257,In_802);
or U712 (N_712,In_291,In_911);
nand U713 (N_713,In_688,In_809);
or U714 (N_714,In_798,In_644);
and U715 (N_715,In_76,In_724);
and U716 (N_716,In_937,In_477);
and U717 (N_717,In_390,In_133);
nor U718 (N_718,In_443,In_917);
nor U719 (N_719,In_69,In_946);
nand U720 (N_720,In_750,In_939);
nor U721 (N_721,In_702,In_746);
xor U722 (N_722,In_195,In_286);
nor U723 (N_723,In_471,In_498);
nor U724 (N_724,In_932,In_523);
xnor U725 (N_725,In_983,In_761);
xor U726 (N_726,In_642,In_841);
and U727 (N_727,In_470,In_157);
nand U728 (N_728,In_499,In_687);
xnor U729 (N_729,In_913,In_712);
or U730 (N_730,In_389,In_903);
or U731 (N_731,In_804,In_297);
nor U732 (N_732,In_559,In_418);
nand U733 (N_733,In_954,In_122);
nor U734 (N_734,In_389,In_711);
or U735 (N_735,In_846,In_638);
and U736 (N_736,In_631,In_251);
and U737 (N_737,In_902,In_931);
nand U738 (N_738,In_705,In_590);
nand U739 (N_739,In_820,In_185);
or U740 (N_740,In_651,In_805);
or U741 (N_741,In_450,In_758);
nand U742 (N_742,In_553,In_141);
xnor U743 (N_743,In_245,In_754);
nand U744 (N_744,In_592,In_12);
nand U745 (N_745,In_955,In_995);
nor U746 (N_746,In_808,In_127);
and U747 (N_747,In_784,In_246);
and U748 (N_748,In_566,In_404);
or U749 (N_749,In_229,In_571);
or U750 (N_750,In_524,In_672);
nand U751 (N_751,In_814,In_475);
and U752 (N_752,In_684,In_441);
and U753 (N_753,In_828,In_499);
or U754 (N_754,In_600,In_105);
or U755 (N_755,In_712,In_106);
nor U756 (N_756,In_155,In_773);
and U757 (N_757,In_346,In_690);
and U758 (N_758,In_916,In_967);
nor U759 (N_759,In_668,In_624);
nor U760 (N_760,In_864,In_509);
and U761 (N_761,In_911,In_661);
and U762 (N_762,In_485,In_408);
nand U763 (N_763,In_660,In_880);
and U764 (N_764,In_195,In_585);
and U765 (N_765,In_14,In_709);
nand U766 (N_766,In_227,In_143);
or U767 (N_767,In_371,In_436);
and U768 (N_768,In_737,In_209);
and U769 (N_769,In_504,In_584);
or U770 (N_770,In_147,In_472);
and U771 (N_771,In_346,In_936);
or U772 (N_772,In_726,In_832);
and U773 (N_773,In_341,In_498);
nor U774 (N_774,In_693,In_595);
and U775 (N_775,In_317,In_60);
nand U776 (N_776,In_233,In_766);
nor U777 (N_777,In_667,In_369);
or U778 (N_778,In_184,In_302);
and U779 (N_779,In_777,In_333);
nor U780 (N_780,In_772,In_140);
nor U781 (N_781,In_179,In_191);
xor U782 (N_782,In_923,In_669);
and U783 (N_783,In_777,In_661);
and U784 (N_784,In_383,In_83);
or U785 (N_785,In_423,In_818);
nor U786 (N_786,In_195,In_840);
nand U787 (N_787,In_156,In_36);
xnor U788 (N_788,In_689,In_921);
nand U789 (N_789,In_74,In_36);
xnor U790 (N_790,In_248,In_893);
nand U791 (N_791,In_501,In_840);
nor U792 (N_792,In_653,In_44);
or U793 (N_793,In_663,In_735);
nor U794 (N_794,In_931,In_689);
or U795 (N_795,In_374,In_918);
and U796 (N_796,In_253,In_663);
or U797 (N_797,In_197,In_511);
nand U798 (N_798,In_446,In_531);
and U799 (N_799,In_161,In_421);
nand U800 (N_800,In_108,In_662);
nand U801 (N_801,In_309,In_654);
xnor U802 (N_802,In_220,In_642);
and U803 (N_803,In_954,In_770);
or U804 (N_804,In_261,In_681);
nor U805 (N_805,In_58,In_534);
and U806 (N_806,In_413,In_216);
and U807 (N_807,In_938,In_86);
and U808 (N_808,In_210,In_803);
or U809 (N_809,In_133,In_34);
nor U810 (N_810,In_886,In_595);
nor U811 (N_811,In_621,In_158);
or U812 (N_812,In_505,In_224);
nand U813 (N_813,In_481,In_695);
or U814 (N_814,In_291,In_5);
xnor U815 (N_815,In_833,In_780);
and U816 (N_816,In_635,In_659);
xnor U817 (N_817,In_582,In_528);
nand U818 (N_818,In_204,In_821);
nand U819 (N_819,In_519,In_673);
or U820 (N_820,In_545,In_429);
nand U821 (N_821,In_778,In_384);
or U822 (N_822,In_333,In_492);
and U823 (N_823,In_86,In_235);
nand U824 (N_824,In_127,In_374);
nor U825 (N_825,In_699,In_125);
or U826 (N_826,In_840,In_491);
nand U827 (N_827,In_158,In_137);
xnor U828 (N_828,In_122,In_244);
nor U829 (N_829,In_659,In_287);
nand U830 (N_830,In_298,In_614);
nand U831 (N_831,In_71,In_148);
and U832 (N_832,In_241,In_523);
nor U833 (N_833,In_620,In_261);
nor U834 (N_834,In_879,In_560);
nor U835 (N_835,In_882,In_880);
nor U836 (N_836,In_408,In_169);
nor U837 (N_837,In_299,In_155);
nor U838 (N_838,In_416,In_212);
nor U839 (N_839,In_244,In_376);
and U840 (N_840,In_531,In_337);
nor U841 (N_841,In_100,In_372);
nand U842 (N_842,In_32,In_438);
or U843 (N_843,In_17,In_11);
and U844 (N_844,In_503,In_802);
and U845 (N_845,In_170,In_806);
xor U846 (N_846,In_808,In_364);
or U847 (N_847,In_277,In_344);
nor U848 (N_848,In_55,In_364);
or U849 (N_849,In_956,In_831);
nand U850 (N_850,In_309,In_767);
or U851 (N_851,In_132,In_704);
xor U852 (N_852,In_768,In_341);
xor U853 (N_853,In_201,In_72);
and U854 (N_854,In_240,In_15);
nand U855 (N_855,In_658,In_602);
nor U856 (N_856,In_580,In_45);
nor U857 (N_857,In_845,In_776);
nor U858 (N_858,In_155,In_77);
nand U859 (N_859,In_475,In_718);
nor U860 (N_860,In_161,In_615);
and U861 (N_861,In_790,In_714);
nor U862 (N_862,In_284,In_161);
and U863 (N_863,In_115,In_678);
nor U864 (N_864,In_371,In_300);
nor U865 (N_865,In_204,In_147);
nor U866 (N_866,In_653,In_151);
and U867 (N_867,In_437,In_104);
and U868 (N_868,In_328,In_756);
and U869 (N_869,In_999,In_657);
nand U870 (N_870,In_418,In_353);
and U871 (N_871,In_618,In_791);
and U872 (N_872,In_839,In_49);
nand U873 (N_873,In_161,In_253);
or U874 (N_874,In_945,In_3);
nand U875 (N_875,In_274,In_681);
or U876 (N_876,In_12,In_491);
or U877 (N_877,In_156,In_747);
and U878 (N_878,In_290,In_941);
and U879 (N_879,In_687,In_715);
or U880 (N_880,In_232,In_714);
or U881 (N_881,In_130,In_943);
or U882 (N_882,In_5,In_375);
nor U883 (N_883,In_56,In_446);
or U884 (N_884,In_442,In_787);
and U885 (N_885,In_599,In_211);
and U886 (N_886,In_690,In_860);
and U887 (N_887,In_25,In_529);
or U888 (N_888,In_44,In_664);
and U889 (N_889,In_10,In_525);
nor U890 (N_890,In_342,In_667);
nand U891 (N_891,In_517,In_19);
nor U892 (N_892,In_245,In_889);
xnor U893 (N_893,In_812,In_143);
and U894 (N_894,In_791,In_325);
and U895 (N_895,In_257,In_167);
nor U896 (N_896,In_573,In_928);
xor U897 (N_897,In_521,In_374);
or U898 (N_898,In_425,In_179);
and U899 (N_899,In_800,In_625);
nand U900 (N_900,In_748,In_170);
or U901 (N_901,In_960,In_158);
or U902 (N_902,In_775,In_721);
or U903 (N_903,In_24,In_705);
xor U904 (N_904,In_291,In_542);
nor U905 (N_905,In_59,In_674);
xnor U906 (N_906,In_115,In_38);
nor U907 (N_907,In_274,In_999);
nand U908 (N_908,In_854,In_138);
or U909 (N_909,In_249,In_270);
nor U910 (N_910,In_970,In_32);
or U911 (N_911,In_193,In_774);
and U912 (N_912,In_470,In_874);
xor U913 (N_913,In_692,In_814);
nand U914 (N_914,In_622,In_286);
xnor U915 (N_915,In_60,In_302);
and U916 (N_916,In_535,In_395);
and U917 (N_917,In_654,In_885);
nor U918 (N_918,In_538,In_746);
nor U919 (N_919,In_360,In_68);
and U920 (N_920,In_65,In_693);
and U921 (N_921,In_815,In_795);
nor U922 (N_922,In_531,In_663);
and U923 (N_923,In_795,In_690);
nand U924 (N_924,In_73,In_587);
nor U925 (N_925,In_612,In_747);
nor U926 (N_926,In_250,In_860);
nand U927 (N_927,In_887,In_271);
nor U928 (N_928,In_386,In_539);
nor U929 (N_929,In_735,In_650);
nor U930 (N_930,In_835,In_869);
xnor U931 (N_931,In_143,In_743);
or U932 (N_932,In_178,In_263);
or U933 (N_933,In_825,In_268);
or U934 (N_934,In_478,In_293);
and U935 (N_935,In_925,In_604);
nand U936 (N_936,In_546,In_100);
nor U937 (N_937,In_818,In_181);
nand U938 (N_938,In_620,In_933);
nor U939 (N_939,In_3,In_326);
and U940 (N_940,In_313,In_387);
xnor U941 (N_941,In_202,In_644);
nor U942 (N_942,In_64,In_333);
nor U943 (N_943,In_101,In_534);
xnor U944 (N_944,In_443,In_715);
and U945 (N_945,In_190,In_143);
nor U946 (N_946,In_49,In_0);
xnor U947 (N_947,In_218,In_80);
xor U948 (N_948,In_249,In_396);
xnor U949 (N_949,In_595,In_883);
nor U950 (N_950,In_678,In_551);
and U951 (N_951,In_177,In_291);
nor U952 (N_952,In_835,In_710);
or U953 (N_953,In_910,In_562);
or U954 (N_954,In_180,In_872);
nor U955 (N_955,In_222,In_520);
and U956 (N_956,In_576,In_605);
nor U957 (N_957,In_745,In_618);
or U958 (N_958,In_879,In_701);
and U959 (N_959,In_253,In_314);
xor U960 (N_960,In_408,In_677);
xor U961 (N_961,In_980,In_58);
nand U962 (N_962,In_260,In_986);
and U963 (N_963,In_814,In_971);
xor U964 (N_964,In_733,In_42);
nor U965 (N_965,In_911,In_489);
nor U966 (N_966,In_667,In_547);
and U967 (N_967,In_127,In_879);
or U968 (N_968,In_676,In_900);
nor U969 (N_969,In_831,In_259);
and U970 (N_970,In_27,In_721);
and U971 (N_971,In_448,In_337);
nand U972 (N_972,In_881,In_466);
nor U973 (N_973,In_587,In_814);
or U974 (N_974,In_320,In_770);
or U975 (N_975,In_726,In_546);
nor U976 (N_976,In_992,In_728);
nor U977 (N_977,In_330,In_45);
or U978 (N_978,In_239,In_387);
nor U979 (N_979,In_368,In_7);
xor U980 (N_980,In_467,In_970);
xor U981 (N_981,In_48,In_557);
nor U982 (N_982,In_930,In_873);
nor U983 (N_983,In_275,In_310);
nor U984 (N_984,In_283,In_771);
and U985 (N_985,In_69,In_510);
and U986 (N_986,In_88,In_328);
nor U987 (N_987,In_514,In_10);
or U988 (N_988,In_377,In_833);
and U989 (N_989,In_839,In_117);
and U990 (N_990,In_399,In_988);
and U991 (N_991,In_496,In_990);
nor U992 (N_992,In_860,In_193);
and U993 (N_993,In_74,In_890);
nand U994 (N_994,In_52,In_858);
nand U995 (N_995,In_705,In_350);
xor U996 (N_996,In_74,In_340);
nand U997 (N_997,In_835,In_518);
nor U998 (N_998,In_682,In_302);
nor U999 (N_999,In_926,In_995);
or U1000 (N_1000,In_776,In_535);
nand U1001 (N_1001,In_10,In_595);
nand U1002 (N_1002,In_256,In_458);
and U1003 (N_1003,In_816,In_193);
nand U1004 (N_1004,In_994,In_891);
xor U1005 (N_1005,In_61,In_640);
nand U1006 (N_1006,In_856,In_723);
or U1007 (N_1007,In_227,In_857);
and U1008 (N_1008,In_28,In_973);
and U1009 (N_1009,In_113,In_574);
or U1010 (N_1010,In_640,In_116);
nand U1011 (N_1011,In_679,In_617);
or U1012 (N_1012,In_719,In_208);
and U1013 (N_1013,In_757,In_148);
nor U1014 (N_1014,In_882,In_112);
nor U1015 (N_1015,In_557,In_546);
nand U1016 (N_1016,In_616,In_99);
and U1017 (N_1017,In_936,In_150);
nor U1018 (N_1018,In_553,In_801);
or U1019 (N_1019,In_10,In_25);
nand U1020 (N_1020,In_498,In_811);
nand U1021 (N_1021,In_508,In_238);
nor U1022 (N_1022,In_849,In_929);
nand U1023 (N_1023,In_736,In_425);
nor U1024 (N_1024,In_10,In_486);
or U1025 (N_1025,In_680,In_345);
or U1026 (N_1026,In_170,In_662);
or U1027 (N_1027,In_803,In_79);
nor U1028 (N_1028,In_30,In_615);
nand U1029 (N_1029,In_815,In_423);
and U1030 (N_1030,In_518,In_614);
and U1031 (N_1031,In_817,In_419);
nand U1032 (N_1032,In_381,In_912);
and U1033 (N_1033,In_208,In_549);
nor U1034 (N_1034,In_392,In_653);
nand U1035 (N_1035,In_921,In_869);
and U1036 (N_1036,In_981,In_638);
and U1037 (N_1037,In_687,In_105);
nor U1038 (N_1038,In_77,In_430);
nand U1039 (N_1039,In_143,In_560);
and U1040 (N_1040,In_871,In_626);
or U1041 (N_1041,In_483,In_339);
nand U1042 (N_1042,In_636,In_942);
or U1043 (N_1043,In_185,In_892);
nand U1044 (N_1044,In_779,In_160);
nand U1045 (N_1045,In_600,In_95);
nor U1046 (N_1046,In_350,In_871);
xnor U1047 (N_1047,In_65,In_222);
and U1048 (N_1048,In_737,In_712);
nor U1049 (N_1049,In_549,In_598);
nand U1050 (N_1050,In_890,In_736);
xnor U1051 (N_1051,In_160,In_203);
nand U1052 (N_1052,In_341,In_774);
nor U1053 (N_1053,In_134,In_407);
or U1054 (N_1054,In_291,In_482);
and U1055 (N_1055,In_304,In_347);
nand U1056 (N_1056,In_577,In_706);
or U1057 (N_1057,In_69,In_479);
nor U1058 (N_1058,In_840,In_219);
nand U1059 (N_1059,In_977,In_653);
and U1060 (N_1060,In_768,In_455);
nand U1061 (N_1061,In_890,In_40);
and U1062 (N_1062,In_210,In_354);
nor U1063 (N_1063,In_488,In_994);
nand U1064 (N_1064,In_144,In_575);
nand U1065 (N_1065,In_574,In_227);
and U1066 (N_1066,In_89,In_724);
nand U1067 (N_1067,In_578,In_597);
and U1068 (N_1068,In_306,In_206);
nor U1069 (N_1069,In_766,In_72);
nor U1070 (N_1070,In_318,In_996);
nand U1071 (N_1071,In_524,In_332);
nand U1072 (N_1072,In_818,In_93);
and U1073 (N_1073,In_906,In_727);
or U1074 (N_1074,In_736,In_910);
nand U1075 (N_1075,In_437,In_352);
nand U1076 (N_1076,In_211,In_614);
xor U1077 (N_1077,In_462,In_295);
or U1078 (N_1078,In_57,In_832);
nor U1079 (N_1079,In_466,In_379);
or U1080 (N_1080,In_769,In_415);
nand U1081 (N_1081,In_237,In_850);
and U1082 (N_1082,In_729,In_806);
nand U1083 (N_1083,In_733,In_167);
nand U1084 (N_1084,In_546,In_140);
and U1085 (N_1085,In_785,In_93);
and U1086 (N_1086,In_418,In_688);
xor U1087 (N_1087,In_887,In_35);
nand U1088 (N_1088,In_693,In_561);
nor U1089 (N_1089,In_20,In_599);
nand U1090 (N_1090,In_144,In_836);
nand U1091 (N_1091,In_560,In_57);
xor U1092 (N_1092,In_424,In_843);
or U1093 (N_1093,In_420,In_425);
and U1094 (N_1094,In_331,In_6);
nor U1095 (N_1095,In_26,In_480);
or U1096 (N_1096,In_481,In_293);
and U1097 (N_1097,In_514,In_549);
nand U1098 (N_1098,In_460,In_293);
and U1099 (N_1099,In_314,In_470);
and U1100 (N_1100,In_29,In_763);
nand U1101 (N_1101,In_508,In_648);
nor U1102 (N_1102,In_738,In_96);
nand U1103 (N_1103,In_77,In_494);
or U1104 (N_1104,In_362,In_743);
and U1105 (N_1105,In_365,In_261);
nor U1106 (N_1106,In_807,In_981);
xnor U1107 (N_1107,In_170,In_911);
nand U1108 (N_1108,In_389,In_989);
or U1109 (N_1109,In_934,In_255);
or U1110 (N_1110,In_38,In_76);
nand U1111 (N_1111,In_850,In_349);
nor U1112 (N_1112,In_882,In_468);
and U1113 (N_1113,In_86,In_738);
nand U1114 (N_1114,In_819,In_817);
nand U1115 (N_1115,In_635,In_711);
and U1116 (N_1116,In_348,In_799);
xnor U1117 (N_1117,In_885,In_465);
nor U1118 (N_1118,In_213,In_696);
and U1119 (N_1119,In_658,In_500);
nor U1120 (N_1120,In_688,In_675);
or U1121 (N_1121,In_407,In_919);
or U1122 (N_1122,In_261,In_18);
or U1123 (N_1123,In_409,In_790);
nor U1124 (N_1124,In_173,In_197);
and U1125 (N_1125,In_885,In_578);
nor U1126 (N_1126,In_725,In_90);
nor U1127 (N_1127,In_640,In_714);
and U1128 (N_1128,In_610,In_287);
nor U1129 (N_1129,In_878,In_877);
and U1130 (N_1130,In_335,In_240);
xnor U1131 (N_1131,In_794,In_7);
nor U1132 (N_1132,In_417,In_353);
and U1133 (N_1133,In_532,In_498);
nand U1134 (N_1134,In_608,In_527);
nand U1135 (N_1135,In_213,In_632);
or U1136 (N_1136,In_765,In_593);
xor U1137 (N_1137,In_333,In_790);
or U1138 (N_1138,In_895,In_933);
nor U1139 (N_1139,In_362,In_924);
nor U1140 (N_1140,In_68,In_791);
or U1141 (N_1141,In_789,In_895);
nor U1142 (N_1142,In_657,In_990);
and U1143 (N_1143,In_206,In_776);
nand U1144 (N_1144,In_125,In_293);
or U1145 (N_1145,In_515,In_993);
or U1146 (N_1146,In_793,In_377);
nand U1147 (N_1147,In_172,In_169);
or U1148 (N_1148,In_996,In_523);
or U1149 (N_1149,In_885,In_683);
nor U1150 (N_1150,In_961,In_254);
or U1151 (N_1151,In_705,In_834);
nor U1152 (N_1152,In_116,In_219);
or U1153 (N_1153,In_422,In_900);
xnor U1154 (N_1154,In_29,In_851);
nand U1155 (N_1155,In_267,In_838);
and U1156 (N_1156,In_598,In_213);
and U1157 (N_1157,In_472,In_506);
nor U1158 (N_1158,In_582,In_891);
and U1159 (N_1159,In_799,In_735);
nand U1160 (N_1160,In_488,In_210);
xnor U1161 (N_1161,In_834,In_833);
nand U1162 (N_1162,In_689,In_540);
or U1163 (N_1163,In_885,In_875);
and U1164 (N_1164,In_592,In_932);
and U1165 (N_1165,In_957,In_40);
nand U1166 (N_1166,In_265,In_743);
or U1167 (N_1167,In_900,In_404);
or U1168 (N_1168,In_992,In_211);
and U1169 (N_1169,In_62,In_188);
and U1170 (N_1170,In_392,In_49);
and U1171 (N_1171,In_281,In_297);
or U1172 (N_1172,In_818,In_576);
nand U1173 (N_1173,In_854,In_941);
or U1174 (N_1174,In_666,In_294);
nor U1175 (N_1175,In_124,In_293);
nand U1176 (N_1176,In_382,In_508);
or U1177 (N_1177,In_917,In_200);
and U1178 (N_1178,In_125,In_558);
nand U1179 (N_1179,In_10,In_287);
nand U1180 (N_1180,In_358,In_308);
and U1181 (N_1181,In_139,In_1);
nor U1182 (N_1182,In_198,In_203);
nand U1183 (N_1183,In_271,In_977);
nand U1184 (N_1184,In_592,In_845);
or U1185 (N_1185,In_657,In_639);
nor U1186 (N_1186,In_221,In_244);
nor U1187 (N_1187,In_692,In_720);
or U1188 (N_1188,In_141,In_598);
or U1189 (N_1189,In_412,In_201);
and U1190 (N_1190,In_173,In_90);
or U1191 (N_1191,In_398,In_458);
xnor U1192 (N_1192,In_352,In_764);
xnor U1193 (N_1193,In_171,In_272);
and U1194 (N_1194,In_983,In_284);
nand U1195 (N_1195,In_777,In_706);
and U1196 (N_1196,In_267,In_826);
or U1197 (N_1197,In_872,In_559);
or U1198 (N_1198,In_728,In_715);
xor U1199 (N_1199,In_87,In_831);
and U1200 (N_1200,In_581,In_460);
or U1201 (N_1201,In_24,In_627);
or U1202 (N_1202,In_89,In_517);
nor U1203 (N_1203,In_258,In_193);
or U1204 (N_1204,In_913,In_740);
and U1205 (N_1205,In_666,In_237);
or U1206 (N_1206,In_868,In_995);
and U1207 (N_1207,In_329,In_226);
nand U1208 (N_1208,In_99,In_583);
nor U1209 (N_1209,In_486,In_952);
and U1210 (N_1210,In_499,In_803);
or U1211 (N_1211,In_968,In_433);
nor U1212 (N_1212,In_497,In_967);
nor U1213 (N_1213,In_465,In_305);
nand U1214 (N_1214,In_884,In_554);
nand U1215 (N_1215,In_62,In_932);
nor U1216 (N_1216,In_286,In_563);
or U1217 (N_1217,In_79,In_853);
xnor U1218 (N_1218,In_911,In_873);
or U1219 (N_1219,In_638,In_111);
xnor U1220 (N_1220,In_884,In_276);
xnor U1221 (N_1221,In_684,In_861);
and U1222 (N_1222,In_23,In_350);
and U1223 (N_1223,In_49,In_205);
nand U1224 (N_1224,In_168,In_32);
and U1225 (N_1225,In_984,In_409);
xor U1226 (N_1226,In_185,In_386);
or U1227 (N_1227,In_881,In_397);
nand U1228 (N_1228,In_723,In_720);
nor U1229 (N_1229,In_889,In_520);
and U1230 (N_1230,In_646,In_433);
and U1231 (N_1231,In_195,In_344);
and U1232 (N_1232,In_640,In_946);
or U1233 (N_1233,In_354,In_611);
and U1234 (N_1234,In_747,In_494);
and U1235 (N_1235,In_714,In_187);
and U1236 (N_1236,In_362,In_583);
nor U1237 (N_1237,In_955,In_776);
xnor U1238 (N_1238,In_989,In_102);
and U1239 (N_1239,In_792,In_967);
xnor U1240 (N_1240,In_270,In_317);
nand U1241 (N_1241,In_456,In_665);
and U1242 (N_1242,In_739,In_218);
and U1243 (N_1243,In_562,In_205);
or U1244 (N_1244,In_508,In_943);
nor U1245 (N_1245,In_562,In_210);
and U1246 (N_1246,In_983,In_739);
or U1247 (N_1247,In_497,In_248);
and U1248 (N_1248,In_338,In_804);
nor U1249 (N_1249,In_663,In_242);
nor U1250 (N_1250,In_147,In_877);
nor U1251 (N_1251,In_568,In_310);
or U1252 (N_1252,In_776,In_209);
xor U1253 (N_1253,In_873,In_70);
or U1254 (N_1254,In_594,In_295);
and U1255 (N_1255,In_104,In_952);
nor U1256 (N_1256,In_852,In_58);
and U1257 (N_1257,In_57,In_195);
nand U1258 (N_1258,In_876,In_762);
or U1259 (N_1259,In_225,In_886);
nor U1260 (N_1260,In_781,In_657);
xor U1261 (N_1261,In_316,In_143);
and U1262 (N_1262,In_524,In_366);
or U1263 (N_1263,In_280,In_343);
xor U1264 (N_1264,In_584,In_254);
nor U1265 (N_1265,In_114,In_169);
nand U1266 (N_1266,In_155,In_611);
or U1267 (N_1267,In_529,In_333);
xnor U1268 (N_1268,In_401,In_472);
and U1269 (N_1269,In_768,In_18);
nand U1270 (N_1270,In_601,In_15);
nor U1271 (N_1271,In_626,In_479);
or U1272 (N_1272,In_502,In_145);
nand U1273 (N_1273,In_536,In_422);
nand U1274 (N_1274,In_109,In_430);
and U1275 (N_1275,In_1,In_16);
xor U1276 (N_1276,In_338,In_501);
nand U1277 (N_1277,In_69,In_368);
nor U1278 (N_1278,In_656,In_154);
and U1279 (N_1279,In_731,In_972);
nand U1280 (N_1280,In_991,In_555);
nand U1281 (N_1281,In_470,In_184);
xor U1282 (N_1282,In_208,In_20);
nor U1283 (N_1283,In_431,In_291);
nor U1284 (N_1284,In_109,In_389);
or U1285 (N_1285,In_927,In_367);
nor U1286 (N_1286,In_296,In_563);
or U1287 (N_1287,In_57,In_495);
nand U1288 (N_1288,In_818,In_68);
nand U1289 (N_1289,In_371,In_64);
nor U1290 (N_1290,In_86,In_66);
nand U1291 (N_1291,In_23,In_659);
nor U1292 (N_1292,In_342,In_157);
xnor U1293 (N_1293,In_876,In_341);
and U1294 (N_1294,In_436,In_481);
or U1295 (N_1295,In_669,In_233);
and U1296 (N_1296,In_431,In_427);
or U1297 (N_1297,In_673,In_232);
nor U1298 (N_1298,In_370,In_126);
xnor U1299 (N_1299,In_376,In_309);
nor U1300 (N_1300,In_739,In_433);
nand U1301 (N_1301,In_162,In_437);
xor U1302 (N_1302,In_852,In_938);
or U1303 (N_1303,In_440,In_932);
or U1304 (N_1304,In_257,In_251);
and U1305 (N_1305,In_46,In_82);
nand U1306 (N_1306,In_584,In_862);
xor U1307 (N_1307,In_59,In_931);
nand U1308 (N_1308,In_353,In_465);
nor U1309 (N_1309,In_713,In_838);
and U1310 (N_1310,In_241,In_485);
or U1311 (N_1311,In_216,In_37);
nor U1312 (N_1312,In_359,In_431);
or U1313 (N_1313,In_114,In_670);
or U1314 (N_1314,In_174,In_827);
nand U1315 (N_1315,In_671,In_366);
nor U1316 (N_1316,In_793,In_522);
and U1317 (N_1317,In_388,In_747);
nand U1318 (N_1318,In_177,In_422);
xnor U1319 (N_1319,In_68,In_59);
nand U1320 (N_1320,In_145,In_373);
or U1321 (N_1321,In_657,In_318);
and U1322 (N_1322,In_140,In_883);
nand U1323 (N_1323,In_746,In_547);
xnor U1324 (N_1324,In_32,In_734);
nand U1325 (N_1325,In_684,In_969);
nor U1326 (N_1326,In_333,In_100);
nand U1327 (N_1327,In_6,In_534);
or U1328 (N_1328,In_304,In_828);
or U1329 (N_1329,In_628,In_979);
and U1330 (N_1330,In_318,In_839);
or U1331 (N_1331,In_483,In_301);
or U1332 (N_1332,In_867,In_677);
and U1333 (N_1333,In_263,In_817);
nand U1334 (N_1334,In_691,In_531);
and U1335 (N_1335,In_550,In_851);
nor U1336 (N_1336,In_499,In_32);
nor U1337 (N_1337,In_660,In_947);
nand U1338 (N_1338,In_212,In_731);
nand U1339 (N_1339,In_85,In_722);
or U1340 (N_1340,In_906,In_798);
nand U1341 (N_1341,In_673,In_382);
and U1342 (N_1342,In_779,In_598);
and U1343 (N_1343,In_781,In_530);
nor U1344 (N_1344,In_999,In_605);
nand U1345 (N_1345,In_800,In_155);
nand U1346 (N_1346,In_266,In_757);
nand U1347 (N_1347,In_376,In_213);
or U1348 (N_1348,In_461,In_552);
and U1349 (N_1349,In_126,In_418);
and U1350 (N_1350,In_50,In_681);
nor U1351 (N_1351,In_722,In_327);
nor U1352 (N_1352,In_906,In_606);
or U1353 (N_1353,In_741,In_119);
and U1354 (N_1354,In_833,In_492);
and U1355 (N_1355,In_0,In_3);
nor U1356 (N_1356,In_545,In_457);
and U1357 (N_1357,In_859,In_736);
or U1358 (N_1358,In_284,In_30);
and U1359 (N_1359,In_229,In_550);
nor U1360 (N_1360,In_362,In_150);
nand U1361 (N_1361,In_683,In_526);
or U1362 (N_1362,In_472,In_898);
nor U1363 (N_1363,In_863,In_208);
nor U1364 (N_1364,In_998,In_36);
or U1365 (N_1365,In_858,In_295);
or U1366 (N_1366,In_840,In_31);
and U1367 (N_1367,In_816,In_465);
and U1368 (N_1368,In_489,In_766);
nor U1369 (N_1369,In_508,In_691);
xor U1370 (N_1370,In_310,In_928);
and U1371 (N_1371,In_421,In_414);
nor U1372 (N_1372,In_910,In_686);
and U1373 (N_1373,In_200,In_726);
nor U1374 (N_1374,In_801,In_972);
nor U1375 (N_1375,In_159,In_286);
and U1376 (N_1376,In_675,In_451);
nand U1377 (N_1377,In_400,In_507);
nand U1378 (N_1378,In_337,In_387);
nand U1379 (N_1379,In_322,In_181);
or U1380 (N_1380,In_289,In_878);
and U1381 (N_1381,In_78,In_308);
nor U1382 (N_1382,In_674,In_565);
and U1383 (N_1383,In_595,In_536);
and U1384 (N_1384,In_128,In_871);
and U1385 (N_1385,In_919,In_337);
nand U1386 (N_1386,In_37,In_128);
and U1387 (N_1387,In_93,In_217);
and U1388 (N_1388,In_362,In_972);
and U1389 (N_1389,In_413,In_877);
xnor U1390 (N_1390,In_119,In_539);
nor U1391 (N_1391,In_874,In_292);
and U1392 (N_1392,In_727,In_504);
nand U1393 (N_1393,In_826,In_599);
nor U1394 (N_1394,In_312,In_174);
or U1395 (N_1395,In_288,In_194);
nand U1396 (N_1396,In_96,In_918);
xor U1397 (N_1397,In_286,In_81);
xnor U1398 (N_1398,In_865,In_634);
nand U1399 (N_1399,In_233,In_213);
and U1400 (N_1400,In_680,In_538);
xnor U1401 (N_1401,In_189,In_223);
xnor U1402 (N_1402,In_247,In_846);
nand U1403 (N_1403,In_384,In_55);
and U1404 (N_1404,In_398,In_673);
or U1405 (N_1405,In_665,In_369);
nor U1406 (N_1406,In_996,In_449);
or U1407 (N_1407,In_529,In_101);
or U1408 (N_1408,In_983,In_637);
nand U1409 (N_1409,In_182,In_266);
nor U1410 (N_1410,In_857,In_155);
nand U1411 (N_1411,In_8,In_380);
or U1412 (N_1412,In_271,In_680);
nor U1413 (N_1413,In_990,In_677);
and U1414 (N_1414,In_458,In_28);
and U1415 (N_1415,In_911,In_120);
nand U1416 (N_1416,In_959,In_110);
or U1417 (N_1417,In_502,In_3);
and U1418 (N_1418,In_22,In_104);
and U1419 (N_1419,In_188,In_209);
or U1420 (N_1420,In_972,In_368);
or U1421 (N_1421,In_179,In_692);
and U1422 (N_1422,In_815,In_261);
nor U1423 (N_1423,In_962,In_30);
nor U1424 (N_1424,In_495,In_114);
nor U1425 (N_1425,In_87,In_429);
nor U1426 (N_1426,In_896,In_63);
nor U1427 (N_1427,In_803,In_810);
nand U1428 (N_1428,In_209,In_688);
and U1429 (N_1429,In_823,In_159);
nor U1430 (N_1430,In_2,In_184);
xnor U1431 (N_1431,In_704,In_9);
nor U1432 (N_1432,In_729,In_585);
nand U1433 (N_1433,In_467,In_735);
nand U1434 (N_1434,In_30,In_926);
or U1435 (N_1435,In_717,In_875);
nand U1436 (N_1436,In_927,In_391);
and U1437 (N_1437,In_770,In_747);
nor U1438 (N_1438,In_270,In_146);
xor U1439 (N_1439,In_580,In_574);
nor U1440 (N_1440,In_537,In_585);
or U1441 (N_1441,In_196,In_740);
or U1442 (N_1442,In_481,In_514);
nand U1443 (N_1443,In_402,In_940);
or U1444 (N_1444,In_416,In_607);
nor U1445 (N_1445,In_703,In_468);
xnor U1446 (N_1446,In_140,In_66);
xnor U1447 (N_1447,In_177,In_475);
and U1448 (N_1448,In_193,In_319);
and U1449 (N_1449,In_522,In_338);
nor U1450 (N_1450,In_842,In_214);
nand U1451 (N_1451,In_251,In_336);
nor U1452 (N_1452,In_848,In_244);
and U1453 (N_1453,In_501,In_27);
nor U1454 (N_1454,In_628,In_744);
nand U1455 (N_1455,In_986,In_332);
nor U1456 (N_1456,In_584,In_210);
or U1457 (N_1457,In_194,In_236);
nor U1458 (N_1458,In_636,In_235);
or U1459 (N_1459,In_30,In_16);
or U1460 (N_1460,In_358,In_491);
or U1461 (N_1461,In_763,In_665);
or U1462 (N_1462,In_859,In_616);
and U1463 (N_1463,In_134,In_950);
and U1464 (N_1464,In_681,In_244);
or U1465 (N_1465,In_538,In_182);
and U1466 (N_1466,In_492,In_209);
or U1467 (N_1467,In_792,In_63);
xor U1468 (N_1468,In_404,In_491);
and U1469 (N_1469,In_342,In_406);
nor U1470 (N_1470,In_584,In_880);
and U1471 (N_1471,In_31,In_906);
nand U1472 (N_1472,In_621,In_566);
or U1473 (N_1473,In_299,In_377);
and U1474 (N_1474,In_700,In_29);
or U1475 (N_1475,In_730,In_509);
and U1476 (N_1476,In_140,In_538);
nand U1477 (N_1477,In_547,In_840);
nor U1478 (N_1478,In_523,In_278);
nor U1479 (N_1479,In_284,In_437);
or U1480 (N_1480,In_782,In_171);
or U1481 (N_1481,In_411,In_762);
or U1482 (N_1482,In_62,In_377);
or U1483 (N_1483,In_380,In_31);
and U1484 (N_1484,In_613,In_824);
nand U1485 (N_1485,In_445,In_577);
nor U1486 (N_1486,In_303,In_98);
and U1487 (N_1487,In_209,In_591);
and U1488 (N_1488,In_946,In_327);
or U1489 (N_1489,In_627,In_311);
xor U1490 (N_1490,In_385,In_505);
nor U1491 (N_1491,In_259,In_167);
nand U1492 (N_1492,In_422,In_27);
xor U1493 (N_1493,In_689,In_752);
or U1494 (N_1494,In_867,In_840);
nor U1495 (N_1495,In_345,In_577);
nor U1496 (N_1496,In_140,In_365);
nor U1497 (N_1497,In_961,In_536);
xnor U1498 (N_1498,In_70,In_148);
and U1499 (N_1499,In_201,In_738);
nor U1500 (N_1500,In_765,In_557);
nor U1501 (N_1501,In_840,In_276);
and U1502 (N_1502,In_973,In_296);
nor U1503 (N_1503,In_511,In_661);
nor U1504 (N_1504,In_138,In_24);
and U1505 (N_1505,In_861,In_993);
nor U1506 (N_1506,In_894,In_305);
and U1507 (N_1507,In_474,In_386);
nand U1508 (N_1508,In_948,In_149);
nor U1509 (N_1509,In_58,In_471);
or U1510 (N_1510,In_232,In_352);
nor U1511 (N_1511,In_124,In_851);
nor U1512 (N_1512,In_323,In_199);
nand U1513 (N_1513,In_204,In_330);
or U1514 (N_1514,In_285,In_727);
and U1515 (N_1515,In_338,In_274);
and U1516 (N_1516,In_878,In_784);
xor U1517 (N_1517,In_581,In_142);
nand U1518 (N_1518,In_32,In_181);
xnor U1519 (N_1519,In_478,In_369);
or U1520 (N_1520,In_850,In_350);
nand U1521 (N_1521,In_59,In_29);
and U1522 (N_1522,In_419,In_773);
nand U1523 (N_1523,In_461,In_900);
nor U1524 (N_1524,In_98,In_619);
nor U1525 (N_1525,In_725,In_435);
and U1526 (N_1526,In_273,In_164);
nand U1527 (N_1527,In_221,In_455);
xor U1528 (N_1528,In_115,In_375);
xor U1529 (N_1529,In_462,In_360);
and U1530 (N_1530,In_677,In_81);
or U1531 (N_1531,In_325,In_146);
or U1532 (N_1532,In_75,In_533);
and U1533 (N_1533,In_733,In_803);
or U1534 (N_1534,In_206,In_431);
or U1535 (N_1535,In_513,In_659);
and U1536 (N_1536,In_304,In_134);
and U1537 (N_1537,In_615,In_638);
nor U1538 (N_1538,In_369,In_68);
or U1539 (N_1539,In_866,In_763);
and U1540 (N_1540,In_89,In_38);
and U1541 (N_1541,In_382,In_649);
xnor U1542 (N_1542,In_438,In_221);
xnor U1543 (N_1543,In_383,In_300);
or U1544 (N_1544,In_198,In_669);
nor U1545 (N_1545,In_879,In_743);
nand U1546 (N_1546,In_664,In_400);
nand U1547 (N_1547,In_907,In_919);
or U1548 (N_1548,In_415,In_11);
or U1549 (N_1549,In_96,In_962);
or U1550 (N_1550,In_556,In_597);
nor U1551 (N_1551,In_879,In_100);
nor U1552 (N_1552,In_51,In_53);
and U1553 (N_1553,In_762,In_875);
nand U1554 (N_1554,In_395,In_812);
nor U1555 (N_1555,In_581,In_628);
and U1556 (N_1556,In_645,In_789);
or U1557 (N_1557,In_44,In_805);
and U1558 (N_1558,In_971,In_904);
nand U1559 (N_1559,In_514,In_576);
or U1560 (N_1560,In_698,In_983);
nand U1561 (N_1561,In_749,In_22);
and U1562 (N_1562,In_727,In_667);
nand U1563 (N_1563,In_476,In_731);
xnor U1564 (N_1564,In_751,In_600);
and U1565 (N_1565,In_675,In_867);
nand U1566 (N_1566,In_732,In_421);
and U1567 (N_1567,In_937,In_23);
nand U1568 (N_1568,In_10,In_896);
nor U1569 (N_1569,In_879,In_550);
nand U1570 (N_1570,In_207,In_982);
nor U1571 (N_1571,In_263,In_905);
nand U1572 (N_1572,In_239,In_910);
nand U1573 (N_1573,In_920,In_370);
nor U1574 (N_1574,In_655,In_291);
or U1575 (N_1575,In_598,In_275);
nand U1576 (N_1576,In_808,In_859);
nor U1577 (N_1577,In_7,In_948);
xnor U1578 (N_1578,In_534,In_775);
or U1579 (N_1579,In_827,In_602);
nand U1580 (N_1580,In_415,In_896);
nor U1581 (N_1581,In_963,In_775);
nand U1582 (N_1582,In_537,In_176);
and U1583 (N_1583,In_679,In_912);
xor U1584 (N_1584,In_988,In_319);
xnor U1585 (N_1585,In_745,In_684);
nor U1586 (N_1586,In_728,In_984);
and U1587 (N_1587,In_257,In_218);
and U1588 (N_1588,In_839,In_233);
or U1589 (N_1589,In_989,In_353);
nand U1590 (N_1590,In_369,In_438);
or U1591 (N_1591,In_297,In_0);
nor U1592 (N_1592,In_368,In_103);
nor U1593 (N_1593,In_127,In_446);
nor U1594 (N_1594,In_987,In_185);
and U1595 (N_1595,In_629,In_2);
or U1596 (N_1596,In_950,In_755);
and U1597 (N_1597,In_989,In_616);
and U1598 (N_1598,In_829,In_605);
or U1599 (N_1599,In_483,In_961);
and U1600 (N_1600,In_639,In_600);
nand U1601 (N_1601,In_390,In_443);
or U1602 (N_1602,In_566,In_364);
or U1603 (N_1603,In_727,In_919);
nand U1604 (N_1604,In_999,In_90);
or U1605 (N_1605,In_997,In_441);
nand U1606 (N_1606,In_988,In_861);
nand U1607 (N_1607,In_791,In_733);
nor U1608 (N_1608,In_628,In_741);
nand U1609 (N_1609,In_707,In_818);
xor U1610 (N_1610,In_886,In_884);
nor U1611 (N_1611,In_847,In_275);
nor U1612 (N_1612,In_567,In_878);
or U1613 (N_1613,In_285,In_632);
nand U1614 (N_1614,In_384,In_170);
xor U1615 (N_1615,In_538,In_889);
or U1616 (N_1616,In_514,In_51);
or U1617 (N_1617,In_6,In_472);
or U1618 (N_1618,In_826,In_387);
xor U1619 (N_1619,In_197,In_658);
and U1620 (N_1620,In_889,In_391);
nand U1621 (N_1621,In_280,In_115);
and U1622 (N_1622,In_879,In_742);
nor U1623 (N_1623,In_397,In_774);
and U1624 (N_1624,In_420,In_736);
or U1625 (N_1625,In_283,In_897);
xor U1626 (N_1626,In_878,In_72);
or U1627 (N_1627,In_58,In_989);
or U1628 (N_1628,In_855,In_971);
nand U1629 (N_1629,In_29,In_67);
and U1630 (N_1630,In_28,In_282);
nand U1631 (N_1631,In_900,In_785);
and U1632 (N_1632,In_115,In_608);
nor U1633 (N_1633,In_107,In_937);
nor U1634 (N_1634,In_311,In_505);
and U1635 (N_1635,In_302,In_542);
xor U1636 (N_1636,In_857,In_60);
nor U1637 (N_1637,In_317,In_567);
and U1638 (N_1638,In_39,In_486);
nand U1639 (N_1639,In_880,In_860);
nand U1640 (N_1640,In_794,In_655);
nor U1641 (N_1641,In_409,In_981);
xnor U1642 (N_1642,In_320,In_949);
and U1643 (N_1643,In_734,In_423);
or U1644 (N_1644,In_68,In_625);
nor U1645 (N_1645,In_402,In_250);
nor U1646 (N_1646,In_753,In_77);
and U1647 (N_1647,In_428,In_225);
or U1648 (N_1648,In_966,In_345);
nor U1649 (N_1649,In_756,In_425);
nand U1650 (N_1650,In_202,In_470);
and U1651 (N_1651,In_852,In_523);
xnor U1652 (N_1652,In_406,In_373);
nand U1653 (N_1653,In_687,In_140);
or U1654 (N_1654,In_329,In_985);
nor U1655 (N_1655,In_165,In_214);
or U1656 (N_1656,In_291,In_513);
and U1657 (N_1657,In_777,In_671);
and U1658 (N_1658,In_146,In_299);
or U1659 (N_1659,In_141,In_72);
xor U1660 (N_1660,In_791,In_310);
or U1661 (N_1661,In_994,In_104);
and U1662 (N_1662,In_801,In_323);
nand U1663 (N_1663,In_232,In_810);
or U1664 (N_1664,In_649,In_697);
or U1665 (N_1665,In_891,In_62);
and U1666 (N_1666,In_868,In_935);
and U1667 (N_1667,In_84,In_8);
nor U1668 (N_1668,In_840,In_925);
nor U1669 (N_1669,In_601,In_185);
nand U1670 (N_1670,In_520,In_802);
nand U1671 (N_1671,In_614,In_360);
and U1672 (N_1672,In_116,In_544);
nor U1673 (N_1673,In_555,In_81);
and U1674 (N_1674,In_375,In_708);
or U1675 (N_1675,In_198,In_622);
nand U1676 (N_1676,In_979,In_25);
and U1677 (N_1677,In_318,In_412);
xnor U1678 (N_1678,In_948,In_116);
and U1679 (N_1679,In_641,In_488);
nand U1680 (N_1680,In_474,In_488);
or U1681 (N_1681,In_495,In_938);
and U1682 (N_1682,In_846,In_42);
and U1683 (N_1683,In_320,In_636);
nor U1684 (N_1684,In_262,In_263);
and U1685 (N_1685,In_830,In_441);
nor U1686 (N_1686,In_175,In_354);
or U1687 (N_1687,In_229,In_685);
and U1688 (N_1688,In_619,In_301);
nor U1689 (N_1689,In_26,In_704);
and U1690 (N_1690,In_502,In_390);
nor U1691 (N_1691,In_783,In_290);
and U1692 (N_1692,In_19,In_149);
nor U1693 (N_1693,In_661,In_37);
xnor U1694 (N_1694,In_382,In_31);
nor U1695 (N_1695,In_126,In_974);
nand U1696 (N_1696,In_910,In_220);
nand U1697 (N_1697,In_412,In_472);
and U1698 (N_1698,In_690,In_940);
nor U1699 (N_1699,In_191,In_395);
nor U1700 (N_1700,In_628,In_577);
or U1701 (N_1701,In_961,In_151);
nand U1702 (N_1702,In_758,In_430);
nor U1703 (N_1703,In_674,In_283);
nor U1704 (N_1704,In_752,In_415);
nand U1705 (N_1705,In_300,In_644);
xnor U1706 (N_1706,In_182,In_312);
nor U1707 (N_1707,In_442,In_343);
or U1708 (N_1708,In_244,In_650);
xor U1709 (N_1709,In_430,In_363);
and U1710 (N_1710,In_270,In_815);
or U1711 (N_1711,In_47,In_387);
nor U1712 (N_1712,In_770,In_883);
xor U1713 (N_1713,In_442,In_593);
nand U1714 (N_1714,In_630,In_379);
nor U1715 (N_1715,In_476,In_688);
xor U1716 (N_1716,In_899,In_293);
or U1717 (N_1717,In_174,In_890);
nand U1718 (N_1718,In_759,In_645);
xnor U1719 (N_1719,In_44,In_526);
nand U1720 (N_1720,In_811,In_878);
and U1721 (N_1721,In_214,In_726);
xnor U1722 (N_1722,In_951,In_801);
and U1723 (N_1723,In_705,In_420);
or U1724 (N_1724,In_46,In_292);
nor U1725 (N_1725,In_123,In_238);
or U1726 (N_1726,In_741,In_321);
nor U1727 (N_1727,In_962,In_713);
nand U1728 (N_1728,In_559,In_624);
or U1729 (N_1729,In_443,In_545);
and U1730 (N_1730,In_610,In_577);
nor U1731 (N_1731,In_33,In_314);
or U1732 (N_1732,In_878,In_164);
nand U1733 (N_1733,In_385,In_127);
nand U1734 (N_1734,In_581,In_802);
nand U1735 (N_1735,In_944,In_543);
xor U1736 (N_1736,In_726,In_206);
nor U1737 (N_1737,In_333,In_269);
nand U1738 (N_1738,In_602,In_906);
and U1739 (N_1739,In_976,In_337);
nor U1740 (N_1740,In_573,In_112);
nand U1741 (N_1741,In_678,In_372);
xor U1742 (N_1742,In_233,In_253);
nand U1743 (N_1743,In_122,In_305);
xor U1744 (N_1744,In_150,In_662);
xor U1745 (N_1745,In_593,In_42);
or U1746 (N_1746,In_600,In_670);
nand U1747 (N_1747,In_703,In_92);
nand U1748 (N_1748,In_727,In_202);
or U1749 (N_1749,In_698,In_158);
and U1750 (N_1750,In_763,In_703);
and U1751 (N_1751,In_404,In_754);
or U1752 (N_1752,In_741,In_980);
nand U1753 (N_1753,In_17,In_27);
and U1754 (N_1754,In_786,In_464);
nand U1755 (N_1755,In_585,In_41);
or U1756 (N_1756,In_218,In_867);
nor U1757 (N_1757,In_243,In_774);
nor U1758 (N_1758,In_257,In_425);
nand U1759 (N_1759,In_144,In_323);
or U1760 (N_1760,In_765,In_346);
nor U1761 (N_1761,In_383,In_136);
or U1762 (N_1762,In_673,In_473);
nand U1763 (N_1763,In_396,In_250);
nand U1764 (N_1764,In_39,In_194);
nand U1765 (N_1765,In_171,In_683);
nor U1766 (N_1766,In_155,In_960);
nor U1767 (N_1767,In_594,In_382);
or U1768 (N_1768,In_870,In_318);
nand U1769 (N_1769,In_371,In_661);
or U1770 (N_1770,In_882,In_729);
and U1771 (N_1771,In_188,In_869);
nand U1772 (N_1772,In_443,In_392);
nor U1773 (N_1773,In_394,In_350);
and U1774 (N_1774,In_19,In_332);
nor U1775 (N_1775,In_185,In_913);
nor U1776 (N_1776,In_706,In_636);
and U1777 (N_1777,In_218,In_55);
xnor U1778 (N_1778,In_775,In_92);
nor U1779 (N_1779,In_350,In_714);
nor U1780 (N_1780,In_918,In_270);
and U1781 (N_1781,In_852,In_524);
nand U1782 (N_1782,In_222,In_838);
nor U1783 (N_1783,In_212,In_954);
or U1784 (N_1784,In_5,In_778);
nand U1785 (N_1785,In_671,In_634);
or U1786 (N_1786,In_439,In_900);
or U1787 (N_1787,In_573,In_455);
and U1788 (N_1788,In_468,In_868);
nand U1789 (N_1789,In_477,In_21);
and U1790 (N_1790,In_198,In_438);
and U1791 (N_1791,In_566,In_692);
and U1792 (N_1792,In_10,In_588);
and U1793 (N_1793,In_866,In_558);
nor U1794 (N_1794,In_573,In_535);
nor U1795 (N_1795,In_621,In_492);
and U1796 (N_1796,In_754,In_588);
xnor U1797 (N_1797,In_190,In_547);
nand U1798 (N_1798,In_386,In_534);
nand U1799 (N_1799,In_549,In_706);
and U1800 (N_1800,In_562,In_843);
nor U1801 (N_1801,In_996,In_582);
nand U1802 (N_1802,In_733,In_756);
or U1803 (N_1803,In_649,In_89);
nor U1804 (N_1804,In_161,In_764);
xnor U1805 (N_1805,In_457,In_423);
and U1806 (N_1806,In_665,In_566);
and U1807 (N_1807,In_578,In_500);
nor U1808 (N_1808,In_264,In_531);
or U1809 (N_1809,In_903,In_826);
nor U1810 (N_1810,In_741,In_671);
and U1811 (N_1811,In_568,In_3);
nor U1812 (N_1812,In_161,In_334);
and U1813 (N_1813,In_81,In_228);
nand U1814 (N_1814,In_25,In_934);
and U1815 (N_1815,In_693,In_238);
nand U1816 (N_1816,In_197,In_1);
nand U1817 (N_1817,In_35,In_861);
nand U1818 (N_1818,In_347,In_723);
nand U1819 (N_1819,In_790,In_391);
and U1820 (N_1820,In_729,In_362);
and U1821 (N_1821,In_489,In_806);
or U1822 (N_1822,In_620,In_637);
nand U1823 (N_1823,In_838,In_310);
and U1824 (N_1824,In_310,In_823);
nand U1825 (N_1825,In_89,In_416);
or U1826 (N_1826,In_112,In_676);
nand U1827 (N_1827,In_969,In_976);
and U1828 (N_1828,In_436,In_243);
nand U1829 (N_1829,In_438,In_342);
nand U1830 (N_1830,In_722,In_477);
and U1831 (N_1831,In_88,In_962);
or U1832 (N_1832,In_400,In_457);
or U1833 (N_1833,In_19,In_177);
nand U1834 (N_1834,In_188,In_384);
nand U1835 (N_1835,In_860,In_570);
and U1836 (N_1836,In_286,In_423);
and U1837 (N_1837,In_316,In_37);
or U1838 (N_1838,In_935,In_642);
xor U1839 (N_1839,In_293,In_291);
and U1840 (N_1840,In_270,In_796);
nand U1841 (N_1841,In_583,In_969);
and U1842 (N_1842,In_437,In_429);
nor U1843 (N_1843,In_372,In_852);
and U1844 (N_1844,In_718,In_237);
or U1845 (N_1845,In_510,In_769);
nand U1846 (N_1846,In_743,In_788);
xor U1847 (N_1847,In_928,In_802);
or U1848 (N_1848,In_565,In_88);
xnor U1849 (N_1849,In_472,In_681);
or U1850 (N_1850,In_466,In_658);
and U1851 (N_1851,In_533,In_921);
and U1852 (N_1852,In_808,In_826);
or U1853 (N_1853,In_242,In_180);
xnor U1854 (N_1854,In_531,In_93);
nor U1855 (N_1855,In_933,In_785);
or U1856 (N_1856,In_687,In_19);
and U1857 (N_1857,In_229,In_60);
xor U1858 (N_1858,In_11,In_456);
nand U1859 (N_1859,In_453,In_288);
or U1860 (N_1860,In_787,In_492);
and U1861 (N_1861,In_329,In_603);
or U1862 (N_1862,In_260,In_943);
nor U1863 (N_1863,In_570,In_152);
and U1864 (N_1864,In_564,In_110);
nand U1865 (N_1865,In_340,In_820);
and U1866 (N_1866,In_771,In_286);
xor U1867 (N_1867,In_198,In_373);
and U1868 (N_1868,In_754,In_681);
or U1869 (N_1869,In_35,In_712);
xor U1870 (N_1870,In_679,In_326);
nand U1871 (N_1871,In_740,In_448);
nand U1872 (N_1872,In_809,In_51);
nand U1873 (N_1873,In_530,In_339);
and U1874 (N_1874,In_10,In_502);
nor U1875 (N_1875,In_46,In_128);
or U1876 (N_1876,In_685,In_67);
xnor U1877 (N_1877,In_229,In_297);
or U1878 (N_1878,In_592,In_486);
nor U1879 (N_1879,In_483,In_895);
xnor U1880 (N_1880,In_473,In_800);
nor U1881 (N_1881,In_716,In_793);
or U1882 (N_1882,In_54,In_313);
or U1883 (N_1883,In_103,In_180);
or U1884 (N_1884,In_380,In_697);
and U1885 (N_1885,In_67,In_937);
or U1886 (N_1886,In_199,In_873);
xor U1887 (N_1887,In_114,In_122);
or U1888 (N_1888,In_559,In_660);
nor U1889 (N_1889,In_450,In_563);
or U1890 (N_1890,In_367,In_627);
or U1891 (N_1891,In_924,In_705);
and U1892 (N_1892,In_520,In_544);
nor U1893 (N_1893,In_562,In_599);
nor U1894 (N_1894,In_706,In_623);
xnor U1895 (N_1895,In_742,In_133);
or U1896 (N_1896,In_334,In_272);
nand U1897 (N_1897,In_884,In_447);
nand U1898 (N_1898,In_835,In_426);
or U1899 (N_1899,In_504,In_184);
nor U1900 (N_1900,In_244,In_604);
and U1901 (N_1901,In_7,In_158);
nor U1902 (N_1902,In_570,In_783);
nor U1903 (N_1903,In_8,In_51);
nand U1904 (N_1904,In_640,In_78);
nand U1905 (N_1905,In_459,In_974);
nand U1906 (N_1906,In_815,In_834);
nand U1907 (N_1907,In_444,In_832);
nand U1908 (N_1908,In_723,In_587);
nand U1909 (N_1909,In_356,In_191);
and U1910 (N_1910,In_367,In_9);
nand U1911 (N_1911,In_449,In_583);
nand U1912 (N_1912,In_612,In_708);
xor U1913 (N_1913,In_695,In_630);
or U1914 (N_1914,In_689,In_120);
nand U1915 (N_1915,In_610,In_661);
nor U1916 (N_1916,In_320,In_111);
nand U1917 (N_1917,In_795,In_577);
nand U1918 (N_1918,In_324,In_915);
nand U1919 (N_1919,In_703,In_132);
nand U1920 (N_1920,In_952,In_803);
or U1921 (N_1921,In_309,In_186);
nand U1922 (N_1922,In_750,In_319);
nor U1923 (N_1923,In_539,In_719);
nand U1924 (N_1924,In_578,In_765);
nand U1925 (N_1925,In_46,In_997);
and U1926 (N_1926,In_20,In_201);
and U1927 (N_1927,In_405,In_748);
or U1928 (N_1928,In_107,In_314);
and U1929 (N_1929,In_919,In_125);
nor U1930 (N_1930,In_714,In_83);
nor U1931 (N_1931,In_512,In_457);
nand U1932 (N_1932,In_852,In_392);
nand U1933 (N_1933,In_619,In_794);
or U1934 (N_1934,In_534,In_249);
nand U1935 (N_1935,In_92,In_171);
or U1936 (N_1936,In_557,In_662);
nor U1937 (N_1937,In_46,In_624);
nor U1938 (N_1938,In_767,In_603);
and U1939 (N_1939,In_745,In_384);
nand U1940 (N_1940,In_245,In_948);
and U1941 (N_1941,In_981,In_261);
and U1942 (N_1942,In_428,In_515);
xor U1943 (N_1943,In_20,In_409);
nand U1944 (N_1944,In_332,In_770);
and U1945 (N_1945,In_374,In_672);
nand U1946 (N_1946,In_563,In_140);
and U1947 (N_1947,In_629,In_83);
or U1948 (N_1948,In_653,In_758);
nor U1949 (N_1949,In_748,In_369);
and U1950 (N_1950,In_982,In_226);
or U1951 (N_1951,In_658,In_992);
and U1952 (N_1952,In_606,In_697);
and U1953 (N_1953,In_426,In_101);
nand U1954 (N_1954,In_412,In_20);
nor U1955 (N_1955,In_588,In_259);
nand U1956 (N_1956,In_368,In_435);
and U1957 (N_1957,In_815,In_81);
xnor U1958 (N_1958,In_154,In_35);
and U1959 (N_1959,In_671,In_345);
xnor U1960 (N_1960,In_864,In_581);
xnor U1961 (N_1961,In_754,In_715);
and U1962 (N_1962,In_743,In_970);
nand U1963 (N_1963,In_543,In_224);
nor U1964 (N_1964,In_377,In_756);
nor U1965 (N_1965,In_610,In_350);
nand U1966 (N_1966,In_957,In_766);
xnor U1967 (N_1967,In_48,In_831);
and U1968 (N_1968,In_557,In_434);
xnor U1969 (N_1969,In_989,In_64);
nor U1970 (N_1970,In_485,In_504);
nand U1971 (N_1971,In_191,In_948);
nor U1972 (N_1972,In_485,In_639);
nor U1973 (N_1973,In_156,In_336);
nor U1974 (N_1974,In_897,In_388);
nor U1975 (N_1975,In_520,In_662);
nor U1976 (N_1976,In_993,In_582);
nand U1977 (N_1977,In_744,In_532);
and U1978 (N_1978,In_1,In_163);
nand U1979 (N_1979,In_379,In_625);
nand U1980 (N_1980,In_350,In_22);
xor U1981 (N_1981,In_417,In_249);
and U1982 (N_1982,In_702,In_124);
or U1983 (N_1983,In_401,In_807);
and U1984 (N_1984,In_765,In_364);
nand U1985 (N_1985,In_881,In_785);
or U1986 (N_1986,In_861,In_867);
nand U1987 (N_1987,In_946,In_839);
or U1988 (N_1988,In_915,In_152);
nand U1989 (N_1989,In_677,In_794);
nand U1990 (N_1990,In_545,In_701);
or U1991 (N_1991,In_128,In_199);
nand U1992 (N_1992,In_842,In_213);
xor U1993 (N_1993,In_238,In_295);
and U1994 (N_1994,In_925,In_585);
or U1995 (N_1995,In_382,In_513);
nand U1996 (N_1996,In_77,In_844);
nand U1997 (N_1997,In_499,In_38);
nand U1998 (N_1998,In_368,In_399);
nand U1999 (N_1999,In_327,In_753);
or U2000 (N_2000,In_992,In_715);
nand U2001 (N_2001,In_931,In_569);
or U2002 (N_2002,In_310,In_692);
nor U2003 (N_2003,In_676,In_851);
nand U2004 (N_2004,In_271,In_566);
nand U2005 (N_2005,In_604,In_323);
and U2006 (N_2006,In_652,In_430);
nor U2007 (N_2007,In_159,In_655);
or U2008 (N_2008,In_410,In_557);
nand U2009 (N_2009,In_796,In_97);
and U2010 (N_2010,In_117,In_887);
nor U2011 (N_2011,In_734,In_773);
xnor U2012 (N_2012,In_813,In_125);
xor U2013 (N_2013,In_343,In_38);
nand U2014 (N_2014,In_150,In_61);
nor U2015 (N_2015,In_468,In_173);
xor U2016 (N_2016,In_180,In_788);
nand U2017 (N_2017,In_413,In_555);
nand U2018 (N_2018,In_378,In_484);
nand U2019 (N_2019,In_285,In_806);
nor U2020 (N_2020,In_779,In_618);
or U2021 (N_2021,In_346,In_725);
nor U2022 (N_2022,In_867,In_287);
and U2023 (N_2023,In_562,In_866);
nor U2024 (N_2024,In_480,In_374);
nor U2025 (N_2025,In_535,In_156);
nor U2026 (N_2026,In_250,In_568);
and U2027 (N_2027,In_42,In_871);
and U2028 (N_2028,In_342,In_594);
nand U2029 (N_2029,In_157,In_533);
nand U2030 (N_2030,In_640,In_347);
and U2031 (N_2031,In_899,In_93);
and U2032 (N_2032,In_315,In_961);
and U2033 (N_2033,In_519,In_351);
nand U2034 (N_2034,In_288,In_176);
and U2035 (N_2035,In_783,In_879);
nor U2036 (N_2036,In_807,In_746);
nor U2037 (N_2037,In_566,In_562);
and U2038 (N_2038,In_836,In_172);
and U2039 (N_2039,In_717,In_562);
xnor U2040 (N_2040,In_708,In_596);
and U2041 (N_2041,In_778,In_149);
and U2042 (N_2042,In_179,In_417);
or U2043 (N_2043,In_611,In_207);
nor U2044 (N_2044,In_945,In_899);
nor U2045 (N_2045,In_115,In_49);
or U2046 (N_2046,In_82,In_515);
or U2047 (N_2047,In_837,In_142);
nor U2048 (N_2048,In_163,In_973);
or U2049 (N_2049,In_437,In_678);
and U2050 (N_2050,In_90,In_784);
or U2051 (N_2051,In_497,In_0);
nor U2052 (N_2052,In_993,In_770);
and U2053 (N_2053,In_353,In_70);
or U2054 (N_2054,In_447,In_868);
or U2055 (N_2055,In_654,In_93);
or U2056 (N_2056,In_39,In_622);
or U2057 (N_2057,In_919,In_448);
or U2058 (N_2058,In_270,In_622);
xor U2059 (N_2059,In_639,In_84);
nor U2060 (N_2060,In_921,In_393);
and U2061 (N_2061,In_600,In_987);
nor U2062 (N_2062,In_660,In_11);
or U2063 (N_2063,In_987,In_591);
xor U2064 (N_2064,In_533,In_285);
or U2065 (N_2065,In_777,In_56);
nor U2066 (N_2066,In_59,In_221);
nand U2067 (N_2067,In_632,In_919);
nand U2068 (N_2068,In_475,In_117);
and U2069 (N_2069,In_382,In_411);
and U2070 (N_2070,In_856,In_62);
nand U2071 (N_2071,In_799,In_749);
nand U2072 (N_2072,In_214,In_838);
or U2073 (N_2073,In_429,In_229);
or U2074 (N_2074,In_272,In_153);
nand U2075 (N_2075,In_147,In_766);
nand U2076 (N_2076,In_295,In_514);
nor U2077 (N_2077,In_80,In_400);
nand U2078 (N_2078,In_644,In_635);
and U2079 (N_2079,In_166,In_58);
or U2080 (N_2080,In_911,In_283);
nor U2081 (N_2081,In_223,In_410);
nand U2082 (N_2082,In_713,In_666);
or U2083 (N_2083,In_501,In_220);
nand U2084 (N_2084,In_797,In_560);
xor U2085 (N_2085,In_651,In_661);
nand U2086 (N_2086,In_486,In_200);
and U2087 (N_2087,In_541,In_410);
nand U2088 (N_2088,In_274,In_945);
nand U2089 (N_2089,In_916,In_516);
or U2090 (N_2090,In_927,In_153);
and U2091 (N_2091,In_296,In_883);
and U2092 (N_2092,In_495,In_648);
or U2093 (N_2093,In_311,In_292);
nand U2094 (N_2094,In_583,In_654);
and U2095 (N_2095,In_417,In_734);
and U2096 (N_2096,In_954,In_868);
nor U2097 (N_2097,In_891,In_932);
and U2098 (N_2098,In_659,In_160);
nand U2099 (N_2099,In_303,In_45);
nand U2100 (N_2100,In_902,In_572);
nand U2101 (N_2101,In_358,In_403);
or U2102 (N_2102,In_162,In_184);
and U2103 (N_2103,In_997,In_688);
nand U2104 (N_2104,In_806,In_178);
xnor U2105 (N_2105,In_764,In_464);
nor U2106 (N_2106,In_144,In_284);
or U2107 (N_2107,In_465,In_581);
nor U2108 (N_2108,In_574,In_777);
and U2109 (N_2109,In_118,In_502);
nand U2110 (N_2110,In_162,In_577);
or U2111 (N_2111,In_131,In_577);
or U2112 (N_2112,In_784,In_852);
nand U2113 (N_2113,In_837,In_959);
nor U2114 (N_2114,In_979,In_372);
and U2115 (N_2115,In_142,In_619);
xor U2116 (N_2116,In_989,In_968);
and U2117 (N_2117,In_906,In_779);
or U2118 (N_2118,In_896,In_367);
or U2119 (N_2119,In_141,In_429);
nand U2120 (N_2120,In_450,In_956);
nand U2121 (N_2121,In_579,In_41);
nand U2122 (N_2122,In_717,In_449);
or U2123 (N_2123,In_760,In_887);
and U2124 (N_2124,In_859,In_59);
and U2125 (N_2125,In_947,In_935);
nand U2126 (N_2126,In_834,In_544);
nor U2127 (N_2127,In_907,In_886);
or U2128 (N_2128,In_256,In_401);
or U2129 (N_2129,In_226,In_678);
nor U2130 (N_2130,In_749,In_970);
nor U2131 (N_2131,In_714,In_392);
or U2132 (N_2132,In_246,In_353);
or U2133 (N_2133,In_429,In_666);
xnor U2134 (N_2134,In_304,In_782);
nor U2135 (N_2135,In_807,In_978);
nand U2136 (N_2136,In_822,In_715);
nor U2137 (N_2137,In_137,In_889);
nor U2138 (N_2138,In_913,In_369);
xor U2139 (N_2139,In_284,In_520);
nor U2140 (N_2140,In_571,In_946);
nor U2141 (N_2141,In_99,In_973);
or U2142 (N_2142,In_319,In_386);
xor U2143 (N_2143,In_641,In_389);
or U2144 (N_2144,In_313,In_409);
nor U2145 (N_2145,In_347,In_424);
nor U2146 (N_2146,In_232,In_783);
nor U2147 (N_2147,In_849,In_93);
or U2148 (N_2148,In_773,In_604);
nand U2149 (N_2149,In_130,In_720);
nand U2150 (N_2150,In_726,In_585);
nand U2151 (N_2151,In_496,In_511);
and U2152 (N_2152,In_536,In_242);
and U2153 (N_2153,In_980,In_240);
nor U2154 (N_2154,In_856,In_836);
nand U2155 (N_2155,In_849,In_596);
nand U2156 (N_2156,In_383,In_895);
nand U2157 (N_2157,In_783,In_697);
or U2158 (N_2158,In_275,In_905);
or U2159 (N_2159,In_232,In_6);
xor U2160 (N_2160,In_889,In_735);
nand U2161 (N_2161,In_835,In_672);
and U2162 (N_2162,In_265,In_930);
or U2163 (N_2163,In_353,In_500);
or U2164 (N_2164,In_628,In_689);
and U2165 (N_2165,In_709,In_386);
nor U2166 (N_2166,In_545,In_789);
and U2167 (N_2167,In_716,In_310);
xor U2168 (N_2168,In_138,In_197);
or U2169 (N_2169,In_358,In_21);
nor U2170 (N_2170,In_390,In_474);
nor U2171 (N_2171,In_275,In_581);
nand U2172 (N_2172,In_119,In_441);
nand U2173 (N_2173,In_603,In_33);
xnor U2174 (N_2174,In_257,In_326);
nand U2175 (N_2175,In_814,In_584);
nor U2176 (N_2176,In_908,In_944);
or U2177 (N_2177,In_522,In_615);
nand U2178 (N_2178,In_127,In_205);
nor U2179 (N_2179,In_76,In_915);
and U2180 (N_2180,In_866,In_102);
nor U2181 (N_2181,In_510,In_593);
nand U2182 (N_2182,In_550,In_672);
nor U2183 (N_2183,In_929,In_41);
nor U2184 (N_2184,In_350,In_543);
nor U2185 (N_2185,In_982,In_105);
nand U2186 (N_2186,In_849,In_721);
nand U2187 (N_2187,In_812,In_683);
or U2188 (N_2188,In_724,In_615);
or U2189 (N_2189,In_123,In_591);
xor U2190 (N_2190,In_739,In_934);
nand U2191 (N_2191,In_331,In_940);
and U2192 (N_2192,In_515,In_192);
nand U2193 (N_2193,In_153,In_207);
and U2194 (N_2194,In_433,In_240);
nand U2195 (N_2195,In_711,In_840);
and U2196 (N_2196,In_761,In_909);
and U2197 (N_2197,In_916,In_45);
nand U2198 (N_2198,In_115,In_920);
or U2199 (N_2199,In_932,In_376);
or U2200 (N_2200,In_600,In_208);
or U2201 (N_2201,In_940,In_748);
xnor U2202 (N_2202,In_707,In_859);
and U2203 (N_2203,In_407,In_100);
nand U2204 (N_2204,In_987,In_610);
or U2205 (N_2205,In_517,In_953);
nand U2206 (N_2206,In_685,In_362);
nand U2207 (N_2207,In_627,In_564);
and U2208 (N_2208,In_487,In_921);
or U2209 (N_2209,In_479,In_197);
nor U2210 (N_2210,In_595,In_373);
or U2211 (N_2211,In_458,In_708);
nor U2212 (N_2212,In_469,In_520);
nand U2213 (N_2213,In_508,In_62);
nor U2214 (N_2214,In_659,In_86);
nand U2215 (N_2215,In_231,In_793);
xnor U2216 (N_2216,In_455,In_766);
nor U2217 (N_2217,In_901,In_695);
and U2218 (N_2218,In_822,In_995);
or U2219 (N_2219,In_933,In_155);
nor U2220 (N_2220,In_749,In_111);
nand U2221 (N_2221,In_223,In_781);
and U2222 (N_2222,In_208,In_194);
or U2223 (N_2223,In_894,In_666);
and U2224 (N_2224,In_406,In_424);
or U2225 (N_2225,In_324,In_681);
or U2226 (N_2226,In_285,In_791);
or U2227 (N_2227,In_356,In_296);
nor U2228 (N_2228,In_639,In_815);
nand U2229 (N_2229,In_906,In_209);
and U2230 (N_2230,In_854,In_596);
nand U2231 (N_2231,In_693,In_761);
nand U2232 (N_2232,In_479,In_643);
nand U2233 (N_2233,In_900,In_823);
or U2234 (N_2234,In_952,In_959);
nor U2235 (N_2235,In_189,In_276);
or U2236 (N_2236,In_74,In_98);
or U2237 (N_2237,In_955,In_647);
nor U2238 (N_2238,In_313,In_658);
and U2239 (N_2239,In_565,In_897);
nand U2240 (N_2240,In_115,In_894);
nor U2241 (N_2241,In_124,In_867);
nor U2242 (N_2242,In_944,In_701);
nand U2243 (N_2243,In_807,In_98);
nor U2244 (N_2244,In_135,In_228);
nand U2245 (N_2245,In_686,In_325);
or U2246 (N_2246,In_801,In_0);
or U2247 (N_2247,In_457,In_866);
or U2248 (N_2248,In_239,In_958);
nor U2249 (N_2249,In_277,In_672);
nand U2250 (N_2250,In_8,In_665);
and U2251 (N_2251,In_94,In_616);
and U2252 (N_2252,In_394,In_420);
and U2253 (N_2253,In_883,In_809);
nand U2254 (N_2254,In_320,In_730);
nand U2255 (N_2255,In_95,In_191);
xor U2256 (N_2256,In_924,In_58);
and U2257 (N_2257,In_216,In_414);
or U2258 (N_2258,In_554,In_134);
nor U2259 (N_2259,In_250,In_427);
or U2260 (N_2260,In_506,In_487);
nand U2261 (N_2261,In_487,In_924);
and U2262 (N_2262,In_313,In_173);
nor U2263 (N_2263,In_607,In_96);
and U2264 (N_2264,In_487,In_864);
or U2265 (N_2265,In_710,In_65);
and U2266 (N_2266,In_37,In_775);
nand U2267 (N_2267,In_494,In_461);
nand U2268 (N_2268,In_401,In_899);
or U2269 (N_2269,In_845,In_978);
nor U2270 (N_2270,In_405,In_478);
nor U2271 (N_2271,In_908,In_180);
nand U2272 (N_2272,In_681,In_172);
or U2273 (N_2273,In_991,In_38);
nand U2274 (N_2274,In_753,In_157);
nand U2275 (N_2275,In_843,In_901);
nand U2276 (N_2276,In_272,In_429);
and U2277 (N_2277,In_82,In_69);
nor U2278 (N_2278,In_15,In_965);
xnor U2279 (N_2279,In_929,In_806);
or U2280 (N_2280,In_280,In_360);
nand U2281 (N_2281,In_12,In_652);
nand U2282 (N_2282,In_988,In_736);
or U2283 (N_2283,In_416,In_650);
nor U2284 (N_2284,In_476,In_478);
nor U2285 (N_2285,In_251,In_515);
nand U2286 (N_2286,In_856,In_114);
nand U2287 (N_2287,In_416,In_646);
and U2288 (N_2288,In_928,In_988);
and U2289 (N_2289,In_452,In_525);
nand U2290 (N_2290,In_296,In_947);
xnor U2291 (N_2291,In_962,In_520);
nor U2292 (N_2292,In_457,In_951);
or U2293 (N_2293,In_752,In_283);
or U2294 (N_2294,In_501,In_852);
nor U2295 (N_2295,In_737,In_580);
nand U2296 (N_2296,In_665,In_37);
or U2297 (N_2297,In_93,In_62);
and U2298 (N_2298,In_519,In_750);
nor U2299 (N_2299,In_590,In_8);
nand U2300 (N_2300,In_46,In_536);
and U2301 (N_2301,In_707,In_485);
nand U2302 (N_2302,In_50,In_948);
nor U2303 (N_2303,In_627,In_582);
nor U2304 (N_2304,In_583,In_385);
and U2305 (N_2305,In_583,In_544);
nand U2306 (N_2306,In_887,In_111);
nand U2307 (N_2307,In_534,In_788);
nor U2308 (N_2308,In_773,In_408);
xor U2309 (N_2309,In_763,In_112);
and U2310 (N_2310,In_268,In_850);
nor U2311 (N_2311,In_808,In_568);
nor U2312 (N_2312,In_786,In_14);
nor U2313 (N_2313,In_434,In_231);
nor U2314 (N_2314,In_190,In_838);
nor U2315 (N_2315,In_779,In_636);
xor U2316 (N_2316,In_127,In_567);
or U2317 (N_2317,In_454,In_581);
or U2318 (N_2318,In_274,In_619);
nand U2319 (N_2319,In_175,In_438);
nor U2320 (N_2320,In_854,In_922);
or U2321 (N_2321,In_852,In_485);
or U2322 (N_2322,In_705,In_658);
nor U2323 (N_2323,In_234,In_905);
nor U2324 (N_2324,In_865,In_189);
nand U2325 (N_2325,In_975,In_313);
nor U2326 (N_2326,In_471,In_510);
nand U2327 (N_2327,In_150,In_460);
and U2328 (N_2328,In_471,In_525);
nand U2329 (N_2329,In_494,In_746);
and U2330 (N_2330,In_193,In_997);
and U2331 (N_2331,In_623,In_294);
or U2332 (N_2332,In_481,In_219);
xnor U2333 (N_2333,In_517,In_231);
or U2334 (N_2334,In_992,In_788);
nand U2335 (N_2335,In_195,In_51);
or U2336 (N_2336,In_355,In_78);
xnor U2337 (N_2337,In_107,In_497);
and U2338 (N_2338,In_52,In_544);
or U2339 (N_2339,In_110,In_605);
nor U2340 (N_2340,In_493,In_29);
and U2341 (N_2341,In_883,In_125);
or U2342 (N_2342,In_544,In_212);
and U2343 (N_2343,In_326,In_723);
or U2344 (N_2344,In_808,In_671);
nor U2345 (N_2345,In_653,In_177);
nand U2346 (N_2346,In_282,In_852);
nor U2347 (N_2347,In_395,In_418);
or U2348 (N_2348,In_662,In_456);
nor U2349 (N_2349,In_461,In_916);
xor U2350 (N_2350,In_209,In_992);
nor U2351 (N_2351,In_618,In_587);
nor U2352 (N_2352,In_36,In_214);
nor U2353 (N_2353,In_592,In_474);
or U2354 (N_2354,In_673,In_551);
and U2355 (N_2355,In_994,In_757);
nor U2356 (N_2356,In_482,In_604);
nor U2357 (N_2357,In_201,In_527);
or U2358 (N_2358,In_790,In_555);
nand U2359 (N_2359,In_832,In_723);
or U2360 (N_2360,In_95,In_858);
nor U2361 (N_2361,In_559,In_415);
nand U2362 (N_2362,In_893,In_627);
and U2363 (N_2363,In_414,In_597);
and U2364 (N_2364,In_454,In_771);
xnor U2365 (N_2365,In_333,In_701);
or U2366 (N_2366,In_399,In_9);
and U2367 (N_2367,In_223,In_569);
nand U2368 (N_2368,In_677,In_474);
nor U2369 (N_2369,In_18,In_661);
nor U2370 (N_2370,In_826,In_437);
nor U2371 (N_2371,In_22,In_832);
or U2372 (N_2372,In_390,In_809);
nand U2373 (N_2373,In_520,In_892);
and U2374 (N_2374,In_239,In_188);
and U2375 (N_2375,In_25,In_994);
nand U2376 (N_2376,In_319,In_37);
or U2377 (N_2377,In_917,In_844);
nor U2378 (N_2378,In_416,In_545);
and U2379 (N_2379,In_877,In_626);
nand U2380 (N_2380,In_386,In_209);
nand U2381 (N_2381,In_316,In_718);
nor U2382 (N_2382,In_928,In_244);
nand U2383 (N_2383,In_497,In_806);
or U2384 (N_2384,In_685,In_786);
and U2385 (N_2385,In_631,In_573);
or U2386 (N_2386,In_469,In_712);
nor U2387 (N_2387,In_545,In_106);
and U2388 (N_2388,In_38,In_926);
nand U2389 (N_2389,In_113,In_379);
nand U2390 (N_2390,In_898,In_666);
nor U2391 (N_2391,In_685,In_523);
nand U2392 (N_2392,In_735,In_994);
or U2393 (N_2393,In_7,In_45);
nor U2394 (N_2394,In_673,In_982);
xnor U2395 (N_2395,In_188,In_268);
or U2396 (N_2396,In_520,In_796);
and U2397 (N_2397,In_144,In_173);
and U2398 (N_2398,In_35,In_583);
nor U2399 (N_2399,In_211,In_10);
or U2400 (N_2400,In_260,In_904);
nor U2401 (N_2401,In_739,In_989);
and U2402 (N_2402,In_102,In_682);
nand U2403 (N_2403,In_633,In_573);
nor U2404 (N_2404,In_208,In_216);
nand U2405 (N_2405,In_853,In_928);
or U2406 (N_2406,In_314,In_573);
and U2407 (N_2407,In_236,In_705);
nor U2408 (N_2408,In_831,In_11);
nand U2409 (N_2409,In_546,In_685);
or U2410 (N_2410,In_51,In_531);
or U2411 (N_2411,In_51,In_395);
nand U2412 (N_2412,In_296,In_383);
or U2413 (N_2413,In_834,In_158);
nor U2414 (N_2414,In_835,In_851);
nand U2415 (N_2415,In_262,In_853);
or U2416 (N_2416,In_832,In_25);
nand U2417 (N_2417,In_192,In_760);
nor U2418 (N_2418,In_878,In_281);
nor U2419 (N_2419,In_692,In_603);
and U2420 (N_2420,In_934,In_464);
or U2421 (N_2421,In_125,In_239);
and U2422 (N_2422,In_343,In_861);
nor U2423 (N_2423,In_288,In_803);
or U2424 (N_2424,In_449,In_284);
and U2425 (N_2425,In_72,In_759);
nand U2426 (N_2426,In_453,In_475);
xor U2427 (N_2427,In_515,In_831);
or U2428 (N_2428,In_358,In_674);
or U2429 (N_2429,In_646,In_995);
or U2430 (N_2430,In_952,In_964);
nand U2431 (N_2431,In_554,In_104);
and U2432 (N_2432,In_207,In_709);
nor U2433 (N_2433,In_917,In_298);
or U2434 (N_2434,In_291,In_731);
and U2435 (N_2435,In_623,In_197);
or U2436 (N_2436,In_458,In_197);
xnor U2437 (N_2437,In_931,In_549);
or U2438 (N_2438,In_414,In_749);
and U2439 (N_2439,In_158,In_325);
or U2440 (N_2440,In_619,In_926);
and U2441 (N_2441,In_712,In_114);
or U2442 (N_2442,In_463,In_28);
nor U2443 (N_2443,In_652,In_145);
or U2444 (N_2444,In_272,In_584);
nand U2445 (N_2445,In_640,In_654);
and U2446 (N_2446,In_278,In_767);
nand U2447 (N_2447,In_937,In_485);
and U2448 (N_2448,In_432,In_615);
and U2449 (N_2449,In_190,In_822);
nor U2450 (N_2450,In_181,In_12);
or U2451 (N_2451,In_389,In_638);
and U2452 (N_2452,In_380,In_658);
xor U2453 (N_2453,In_103,In_111);
nand U2454 (N_2454,In_855,In_836);
or U2455 (N_2455,In_695,In_278);
nand U2456 (N_2456,In_56,In_661);
nand U2457 (N_2457,In_549,In_709);
and U2458 (N_2458,In_780,In_157);
nor U2459 (N_2459,In_526,In_855);
or U2460 (N_2460,In_111,In_811);
nand U2461 (N_2461,In_992,In_174);
and U2462 (N_2462,In_194,In_855);
nand U2463 (N_2463,In_659,In_871);
or U2464 (N_2464,In_883,In_80);
or U2465 (N_2465,In_552,In_12);
nor U2466 (N_2466,In_918,In_286);
xor U2467 (N_2467,In_206,In_602);
or U2468 (N_2468,In_917,In_396);
nor U2469 (N_2469,In_359,In_724);
and U2470 (N_2470,In_253,In_507);
nor U2471 (N_2471,In_503,In_923);
or U2472 (N_2472,In_786,In_344);
and U2473 (N_2473,In_582,In_560);
nor U2474 (N_2474,In_261,In_986);
and U2475 (N_2475,In_530,In_793);
or U2476 (N_2476,In_74,In_879);
nor U2477 (N_2477,In_286,In_469);
and U2478 (N_2478,In_809,In_872);
or U2479 (N_2479,In_983,In_130);
or U2480 (N_2480,In_15,In_491);
nand U2481 (N_2481,In_987,In_616);
nand U2482 (N_2482,In_77,In_426);
nand U2483 (N_2483,In_894,In_137);
xnor U2484 (N_2484,In_225,In_423);
and U2485 (N_2485,In_897,In_369);
or U2486 (N_2486,In_232,In_525);
nor U2487 (N_2487,In_256,In_337);
or U2488 (N_2488,In_156,In_34);
or U2489 (N_2489,In_952,In_791);
nand U2490 (N_2490,In_641,In_433);
nand U2491 (N_2491,In_997,In_875);
and U2492 (N_2492,In_911,In_711);
and U2493 (N_2493,In_367,In_708);
or U2494 (N_2494,In_540,In_522);
nor U2495 (N_2495,In_554,In_299);
nor U2496 (N_2496,In_416,In_353);
or U2497 (N_2497,In_794,In_25);
nand U2498 (N_2498,In_740,In_687);
and U2499 (N_2499,In_766,In_31);
nor U2500 (N_2500,N_1949,N_2256);
or U2501 (N_2501,N_953,N_802);
nand U2502 (N_2502,N_2371,N_942);
nand U2503 (N_2503,N_371,N_2293);
and U2504 (N_2504,N_558,N_407);
nand U2505 (N_2505,N_335,N_270);
nor U2506 (N_2506,N_232,N_79);
and U2507 (N_2507,N_1803,N_2282);
or U2508 (N_2508,N_1778,N_2115);
and U2509 (N_2509,N_1311,N_2117);
nand U2510 (N_2510,N_1369,N_2474);
nor U2511 (N_2511,N_295,N_2082);
nor U2512 (N_2512,N_2167,N_561);
xnor U2513 (N_2513,N_639,N_793);
xor U2514 (N_2514,N_1876,N_1859);
nand U2515 (N_2515,N_1097,N_965);
and U2516 (N_2516,N_952,N_279);
and U2517 (N_2517,N_488,N_476);
xor U2518 (N_2518,N_1122,N_1764);
and U2519 (N_2519,N_2468,N_258);
and U2520 (N_2520,N_1210,N_10);
and U2521 (N_2521,N_582,N_85);
or U2522 (N_2522,N_1760,N_2477);
nor U2523 (N_2523,N_2011,N_818);
and U2524 (N_2524,N_119,N_897);
and U2525 (N_2525,N_706,N_579);
nand U2526 (N_2526,N_1249,N_1468);
nand U2527 (N_2527,N_2187,N_1491);
or U2528 (N_2528,N_1966,N_1553);
nor U2529 (N_2529,N_57,N_181);
and U2530 (N_2530,N_66,N_2423);
nor U2531 (N_2531,N_846,N_349);
and U2532 (N_2532,N_1813,N_2027);
nor U2533 (N_2533,N_1717,N_1639);
and U2534 (N_2534,N_1610,N_633);
nand U2535 (N_2535,N_1893,N_1686);
and U2536 (N_2536,N_1772,N_282);
nor U2537 (N_2537,N_2179,N_1008);
and U2538 (N_2538,N_2220,N_506);
nand U2539 (N_2539,N_525,N_1405);
nand U2540 (N_2540,N_1502,N_679);
and U2541 (N_2541,N_1573,N_675);
and U2542 (N_2542,N_1946,N_1499);
or U2543 (N_2543,N_2302,N_1461);
xnor U2544 (N_2544,N_1349,N_2358);
nand U2545 (N_2545,N_2057,N_1913);
nand U2546 (N_2546,N_821,N_625);
nand U2547 (N_2547,N_2460,N_912);
nand U2548 (N_2548,N_1022,N_858);
or U2549 (N_2549,N_2253,N_1234);
or U2550 (N_2550,N_2376,N_1364);
or U2551 (N_2551,N_1714,N_2014);
or U2552 (N_2552,N_510,N_1908);
nand U2553 (N_2553,N_2486,N_636);
nor U2554 (N_2554,N_1986,N_573);
nand U2555 (N_2555,N_1058,N_2160);
nand U2556 (N_2556,N_273,N_137);
or U2557 (N_2557,N_1339,N_712);
and U2558 (N_2558,N_1888,N_2444);
or U2559 (N_2559,N_2055,N_1947);
and U2560 (N_2560,N_1821,N_139);
and U2561 (N_2561,N_452,N_1872);
nor U2562 (N_2562,N_2459,N_1514);
and U2563 (N_2563,N_1165,N_167);
xor U2564 (N_2564,N_728,N_2191);
and U2565 (N_2565,N_461,N_146);
or U2566 (N_2566,N_347,N_1029);
and U2567 (N_2567,N_894,N_1288);
or U2568 (N_2568,N_2306,N_977);
nor U2569 (N_2569,N_2307,N_8);
xor U2570 (N_2570,N_1451,N_1623);
nand U2571 (N_2571,N_751,N_812);
xnor U2572 (N_2572,N_606,N_4);
xor U2573 (N_2573,N_1089,N_958);
and U2574 (N_2574,N_740,N_1634);
or U2575 (N_2575,N_1270,N_2465);
and U2576 (N_2576,N_2332,N_686);
nor U2577 (N_2577,N_1408,N_2135);
and U2578 (N_2578,N_1696,N_1635);
or U2579 (N_2579,N_2397,N_83);
or U2580 (N_2580,N_830,N_1512);
nand U2581 (N_2581,N_1702,N_1419);
or U2582 (N_2582,N_121,N_1409);
nand U2583 (N_2583,N_1593,N_409);
nand U2584 (N_2584,N_304,N_2096);
nand U2585 (N_2585,N_1214,N_1528);
nor U2586 (N_2586,N_1895,N_2217);
or U2587 (N_2587,N_1738,N_2363);
nor U2588 (N_2588,N_382,N_641);
and U2589 (N_2589,N_2399,N_2364);
nand U2590 (N_2590,N_93,N_966);
nor U2591 (N_2591,N_1312,N_1550);
and U2592 (N_2592,N_1358,N_107);
nand U2593 (N_2593,N_1281,N_1681);
or U2594 (N_2594,N_101,N_1636);
nand U2595 (N_2595,N_1782,N_237);
or U2596 (N_2596,N_1551,N_2124);
nor U2597 (N_2597,N_867,N_1077);
nor U2598 (N_2598,N_1651,N_140);
or U2599 (N_2599,N_2294,N_1683);
nor U2600 (N_2600,N_870,N_350);
or U2601 (N_2601,N_22,N_2069);
and U2602 (N_2602,N_1658,N_1154);
nand U2603 (N_2603,N_2456,N_976);
xor U2604 (N_2604,N_1325,N_815);
or U2605 (N_2605,N_1797,N_2114);
or U2606 (N_2606,N_1044,N_1384);
nor U2607 (N_2607,N_2433,N_1924);
nand U2608 (N_2608,N_1383,N_1773);
nand U2609 (N_2609,N_1804,N_441);
nor U2610 (N_2610,N_881,N_127);
nor U2611 (N_2611,N_1024,N_212);
and U2612 (N_2612,N_2046,N_950);
or U2613 (N_2613,N_2085,N_796);
or U2614 (N_2614,N_272,N_138);
or U2615 (N_2615,N_330,N_245);
and U2616 (N_2616,N_709,N_1692);
or U2617 (N_2617,N_1045,N_2080);
xor U2618 (N_2618,N_731,N_2031);
nor U2619 (N_2619,N_789,N_1678);
xor U2620 (N_2620,N_1544,N_188);
nand U2621 (N_2621,N_1386,N_1535);
or U2622 (N_2622,N_586,N_2266);
nand U2623 (N_2623,N_1646,N_192);
and U2624 (N_2624,N_785,N_1227);
nand U2625 (N_2625,N_182,N_1126);
or U2626 (N_2626,N_1439,N_762);
nand U2627 (N_2627,N_1716,N_2149);
nor U2628 (N_2628,N_1516,N_610);
nand U2629 (N_2629,N_780,N_2021);
or U2630 (N_2630,N_1991,N_2182);
or U2631 (N_2631,N_230,N_1508);
and U2632 (N_2632,N_961,N_948);
and U2633 (N_2633,N_2146,N_1236);
xor U2634 (N_2634,N_2095,N_1866);
nand U2635 (N_2635,N_2431,N_309);
and U2636 (N_2636,N_2164,N_2204);
nand U2637 (N_2637,N_102,N_1267);
nand U2638 (N_2638,N_930,N_971);
xor U2639 (N_2639,N_2303,N_2476);
and U2640 (N_2640,N_1243,N_1769);
nor U2641 (N_2641,N_185,N_2375);
and U2642 (N_2642,N_2367,N_296);
nor U2643 (N_2643,N_1590,N_2339);
nor U2644 (N_2644,N_118,N_1560);
xor U2645 (N_2645,N_1273,N_2480);
nand U2646 (N_2646,N_2079,N_1103);
nor U2647 (N_2647,N_1335,N_1819);
and U2648 (N_2648,N_536,N_2059);
nand U2649 (N_2649,N_2242,N_1563);
nand U2650 (N_2650,N_1722,N_219);
nand U2651 (N_2651,N_2331,N_1320);
and U2652 (N_2652,N_1370,N_2207);
nor U2653 (N_2653,N_1071,N_373);
nand U2654 (N_2654,N_736,N_577);
nor U2655 (N_2655,N_1116,N_2357);
and U2656 (N_2656,N_1942,N_1179);
xnor U2657 (N_2657,N_2216,N_1496);
and U2658 (N_2658,N_1928,N_1290);
xor U2659 (N_2659,N_1219,N_2226);
and U2660 (N_2660,N_1840,N_2304);
nand U2661 (N_2661,N_2071,N_143);
xnor U2662 (N_2662,N_1836,N_741);
and U2663 (N_2663,N_984,N_594);
nor U2664 (N_2664,N_1121,N_1604);
nor U2665 (N_2665,N_2052,N_2466);
nor U2666 (N_2666,N_2349,N_1470);
and U2667 (N_2667,N_2263,N_1822);
or U2668 (N_2668,N_38,N_1372);
and U2669 (N_2669,N_822,N_1130);
or U2670 (N_2670,N_1120,N_1504);
xor U2671 (N_2671,N_1157,N_387);
xor U2672 (N_2672,N_206,N_1817);
nand U2673 (N_2673,N_2168,N_1920);
and U2674 (N_2674,N_277,N_571);
nor U2675 (N_2675,N_1968,N_2118);
xnor U2676 (N_2676,N_754,N_547);
or U2677 (N_2677,N_1333,N_1601);
or U2678 (N_2678,N_2255,N_149);
nand U2679 (N_2679,N_554,N_1135);
and U2680 (N_2680,N_1025,N_678);
and U2681 (N_2681,N_2018,N_1088);
and U2682 (N_2682,N_756,N_1919);
nand U2683 (N_2683,N_276,N_1707);
or U2684 (N_2684,N_1595,N_1423);
or U2685 (N_2685,N_2065,N_1753);
nand U2686 (N_2686,N_864,N_2239);
and U2687 (N_2687,N_2224,N_1648);
nor U2688 (N_2688,N_2316,N_2297);
nor U2689 (N_2689,N_49,N_1360);
nand U2690 (N_2690,N_1858,N_2140);
nor U2691 (N_2691,N_1177,N_1425);
or U2692 (N_2692,N_1072,N_1448);
nand U2693 (N_2693,N_1955,N_833);
and U2694 (N_2694,N_2479,N_377);
and U2695 (N_2695,N_1084,N_483);
and U2696 (N_2696,N_1253,N_1390);
and U2697 (N_2697,N_205,N_429);
nor U2698 (N_2698,N_1277,N_1505);
nand U2699 (N_2699,N_60,N_1418);
nor U2700 (N_2700,N_2251,N_1501);
nand U2701 (N_2701,N_346,N_964);
nand U2702 (N_2702,N_1155,N_2133);
nand U2703 (N_2703,N_943,N_220);
nand U2704 (N_2704,N_2038,N_196);
nand U2705 (N_2705,N_1559,N_2436);
or U2706 (N_2706,N_400,N_597);
and U2707 (N_2707,N_2310,N_462);
and U2708 (N_2708,N_334,N_1049);
or U2709 (N_2709,N_502,N_2449);
nand U2710 (N_2710,N_1123,N_1540);
and U2711 (N_2711,N_2193,N_1818);
and U2712 (N_2712,N_1279,N_567);
and U2713 (N_2713,N_1256,N_1331);
or U2714 (N_2714,N_988,N_869);
and U2715 (N_2715,N_499,N_289);
nor U2716 (N_2716,N_1034,N_1060);
and U2717 (N_2717,N_29,N_2268);
nand U2718 (N_2718,N_1857,N_3);
or U2719 (N_2719,N_2377,N_2211);
nor U2720 (N_2720,N_2231,N_260);
xor U2721 (N_2721,N_353,N_148);
nand U2722 (N_2722,N_1790,N_743);
and U2723 (N_2723,N_231,N_1322);
xor U2724 (N_2724,N_836,N_2284);
nor U2725 (N_2725,N_1851,N_100);
and U2726 (N_2726,N_1464,N_1999);
and U2727 (N_2727,N_458,N_543);
nor U2728 (N_2728,N_1201,N_253);
xor U2729 (N_2729,N_877,N_227);
nor U2730 (N_2730,N_255,N_635);
or U2731 (N_2731,N_2396,N_379);
nand U2732 (N_2732,N_120,N_325);
and U2733 (N_2733,N_2298,N_2170);
nand U2734 (N_2734,N_959,N_1276);
nand U2735 (N_2735,N_1712,N_1189);
or U2736 (N_2736,N_1095,N_1028);
nor U2737 (N_2737,N_294,N_1957);
xnor U2738 (N_2738,N_1411,N_696);
nor U2739 (N_2739,N_1997,N_655);
nand U2740 (N_2740,N_2188,N_1641);
xor U2741 (N_2741,N_2393,N_292);
nand U2742 (N_2742,N_742,N_1996);
xnor U2743 (N_2743,N_2219,N_713);
nand U2744 (N_2744,N_565,N_332);
nor U2745 (N_2745,N_1188,N_381);
and U2746 (N_2746,N_16,N_1691);
xnor U2747 (N_2747,N_753,N_218);
nor U2748 (N_2748,N_595,N_1624);
or U2749 (N_2749,N_1291,N_1713);
or U2750 (N_2750,N_2347,N_1037);
xor U2751 (N_2751,N_1298,N_97);
or U2752 (N_2752,N_694,N_1463);
xnor U2753 (N_2753,N_2192,N_122);
xor U2754 (N_2754,N_374,N_1264);
nor U2755 (N_2755,N_1534,N_2309);
or U2756 (N_2756,N_361,N_1096);
and U2757 (N_2757,N_71,N_460);
nor U2758 (N_2758,N_1373,N_541);
or U2759 (N_2759,N_1495,N_1266);
or U2760 (N_2760,N_911,N_962);
nor U2761 (N_2761,N_1376,N_1964);
and U2762 (N_2762,N_421,N_1345);
nor U2763 (N_2763,N_578,N_1557);
or U2764 (N_2764,N_1558,N_774);
xnor U2765 (N_2765,N_1018,N_566);
or U2766 (N_2766,N_689,N_1825);
xor U2767 (N_2767,N_1410,N_1937);
nor U2768 (N_2768,N_1257,N_446);
nand U2769 (N_2769,N_714,N_1216);
nor U2770 (N_2770,N_1746,N_2173);
and U2771 (N_2771,N_2186,N_498);
or U2772 (N_2772,N_2333,N_352);
nor U2773 (N_2773,N_490,N_2241);
and U2774 (N_2774,N_1200,N_267);
or U2775 (N_2775,N_1533,N_1588);
or U2776 (N_2776,N_19,N_1389);
and U2777 (N_2777,N_1391,N_2439);
nor U2778 (N_2778,N_454,N_74);
nand U2779 (N_2779,N_1417,N_1568);
xor U2780 (N_2780,N_393,N_1810);
and U2781 (N_2781,N_23,N_365);
xnor U2782 (N_2782,N_1260,N_87);
nor U2783 (N_2783,N_986,N_702);
nand U2784 (N_2784,N_35,N_1854);
nor U2785 (N_2785,N_505,N_366);
nor U2786 (N_2786,N_624,N_312);
or U2787 (N_2787,N_301,N_851);
or U2788 (N_2788,N_602,N_481);
nor U2789 (N_2789,N_1066,N_399);
and U2790 (N_2790,N_797,N_674);
and U2791 (N_2791,N_1205,N_985);
or U2792 (N_2792,N_1903,N_1412);
nand U2793 (N_2793,N_2485,N_482);
and U2794 (N_2794,N_176,N_1371);
or U2795 (N_2795,N_197,N_521);
nand U2796 (N_2796,N_103,N_1787);
or U2797 (N_2797,N_1892,N_1101);
nand U2798 (N_2798,N_782,N_2395);
xor U2799 (N_2799,N_1190,N_1548);
nor U2800 (N_2800,N_1742,N_336);
and U2801 (N_2801,N_348,N_2350);
nand U2802 (N_2802,N_2155,N_1067);
xor U2803 (N_2803,N_557,N_2249);
and U2804 (N_2804,N_1992,N_1546);
and U2805 (N_2805,N_88,N_601);
and U2806 (N_2806,N_1013,N_1382);
and U2807 (N_2807,N_947,N_1351);
or U2808 (N_2808,N_1299,N_2390);
xnor U2809 (N_2809,N_144,N_2199);
and U2810 (N_2810,N_204,N_1415);
nor U2811 (N_2811,N_738,N_1631);
xor U2812 (N_2812,N_2153,N_522);
nor U2813 (N_2813,N_175,N_1283);
or U2814 (N_2814,N_1282,N_1757);
and U2815 (N_2815,N_2441,N_2006);
and U2816 (N_2816,N_297,N_2003);
xor U2817 (N_2817,N_1628,N_2097);
nor U2818 (N_2818,N_2092,N_263);
or U2819 (N_2819,N_1380,N_1758);
xor U2820 (N_2820,N_2156,N_437);
nand U2821 (N_2821,N_456,N_632);
and U2822 (N_2822,N_2081,N_248);
or U2823 (N_2823,N_1365,N_974);
xor U2824 (N_2824,N_1687,N_2391);
and U2825 (N_2825,N_657,N_173);
or U2826 (N_2826,N_1827,N_1110);
and U2827 (N_2827,N_1134,N_1161);
nor U2828 (N_2828,N_750,N_584);
or U2829 (N_2829,N_1951,N_2105);
nor U2830 (N_2830,N_1950,N_2119);
xnor U2831 (N_2831,N_1662,N_1600);
nand U2832 (N_2832,N_615,N_715);
or U2833 (N_2833,N_1860,N_302);
nand U2834 (N_2834,N_1846,N_1186);
nand U2835 (N_2835,N_2404,N_810);
and U2836 (N_2836,N_198,N_544);
and U2837 (N_2837,N_1584,N_613);
nand U2838 (N_2838,N_708,N_2301);
nand U2839 (N_2839,N_1536,N_600);
or U2840 (N_2840,N_2120,N_767);
or U2841 (N_2841,N_76,N_2416);
nand U2842 (N_2842,N_1618,N_1286);
and U2843 (N_2843,N_1296,N_1021);
nor U2844 (N_2844,N_654,N_72);
nand U2845 (N_2845,N_2317,N_420);
nor U2846 (N_2846,N_653,N_2469);
and U2847 (N_2847,N_628,N_2190);
nor U2848 (N_2848,N_287,N_1209);
or U2849 (N_2849,N_359,N_519);
or U2850 (N_2850,N_2341,N_1245);
nand U2851 (N_2851,N_464,N_2374);
or U2852 (N_2852,N_1674,N_1147);
nand U2853 (N_2853,N_2305,N_2398);
or U2854 (N_2854,N_468,N_1010);
xor U2855 (N_2855,N_939,N_993);
or U2856 (N_2856,N_1578,N_1863);
nand U2857 (N_2857,N_44,N_882);
and U2858 (N_2858,N_752,N_1106);
nand U2859 (N_2859,N_2337,N_707);
nand U2860 (N_2860,N_683,N_323);
xnor U2861 (N_2861,N_735,N_164);
nand U2862 (N_2862,N_795,N_1901);
nand U2863 (N_2863,N_765,N_115);
nor U2864 (N_2864,N_2176,N_2159);
and U2865 (N_2865,N_2023,N_2194);
and U2866 (N_2866,N_885,N_1941);
nand U2867 (N_2867,N_887,N_1706);
nor U2868 (N_2868,N_1800,N_2045);
nor U2869 (N_2869,N_1459,N_643);
nand U2870 (N_2870,N_2148,N_2288);
nand U2871 (N_2871,N_792,N_2030);
nor U2872 (N_2872,N_1726,N_2024);
or U2873 (N_2873,N_883,N_1500);
xnor U2874 (N_2874,N_2126,N_1052);
and U2875 (N_2875,N_906,N_1180);
nor U2876 (N_2876,N_2329,N_430);
nor U2877 (N_2877,N_801,N_2265);
and U2878 (N_2878,N_1137,N_328);
or U2879 (N_2879,N_1416,N_94);
nand U2880 (N_2880,N_945,N_2311);
and U2881 (N_2881,N_1934,N_1329);
nand U2882 (N_2882,N_288,N_426);
and U2883 (N_2883,N_2324,N_2162);
nor U2884 (N_2884,N_886,N_2382);
or U2885 (N_2885,N_2200,N_1644);
nand U2886 (N_2886,N_1393,N_2);
xor U2887 (N_2887,N_484,N_477);
nor U2888 (N_2888,N_1323,N_11);
nand U2889 (N_2889,N_262,N_311);
xor U2890 (N_2890,N_229,N_850);
and U2891 (N_2891,N_473,N_1663);
and U2892 (N_2892,N_788,N_860);
and U2893 (N_2893,N_54,N_711);
and U2894 (N_2894,N_1269,N_1444);
nor U2895 (N_2895,N_1945,N_1927);
and U2896 (N_2896,N_1395,N_2353);
nor U2897 (N_2897,N_507,N_759);
nand U2898 (N_2898,N_1594,N_55);
or U2899 (N_2899,N_1603,N_249);
and U2900 (N_2900,N_2223,N_254);
and U2901 (N_2901,N_2270,N_202);
nand U2902 (N_2902,N_1397,N_1420);
or U2903 (N_2903,N_1642,N_2325);
nand U2904 (N_2904,N_1626,N_1915);
nand U2905 (N_2905,N_256,N_1394);
nor U2906 (N_2906,N_2323,N_1206);
xor U2907 (N_2907,N_1645,N_1525);
nor U2908 (N_2908,N_1781,N_1454);
xor U2909 (N_2909,N_1509,N_1820);
nand U2910 (N_2910,N_2336,N_1515);
nand U2911 (N_2911,N_1304,N_2108);
nor U2912 (N_2912,N_1324,N_369);
xnor U2913 (N_2913,N_2209,N_618);
nor U2914 (N_2914,N_730,N_284);
nor U2915 (N_2915,N_1151,N_1602);
or U2916 (N_2916,N_994,N_898);
xnor U2917 (N_2917,N_1208,N_1359);
xnor U2918 (N_2918,N_533,N_917);
and U2919 (N_2919,N_300,N_1105);
and U2920 (N_2920,N_2446,N_1486);
xnor U2921 (N_2921,N_1056,N_1975);
nand U2922 (N_2922,N_1099,N_1798);
or U2923 (N_2923,N_1343,N_2257);
and U2924 (N_2924,N_2442,N_677);
or U2925 (N_2925,N_1970,N_2036);
or U2926 (N_2926,N_1102,N_1313);
nand U2927 (N_2927,N_1649,N_757);
or U2928 (N_2928,N_2484,N_1144);
or U2929 (N_2929,N_1792,N_408);
nor U2930 (N_2930,N_2315,N_1739);
or U2931 (N_2931,N_370,N_2401);
nor U2932 (N_2932,N_946,N_1995);
and U2933 (N_2933,N_2411,N_384);
nand U2934 (N_2934,N_24,N_1353);
xor U2935 (N_2935,N_2487,N_1724);
nor U2936 (N_2936,N_41,N_1829);
xnor U2937 (N_2937,N_367,N_2061);
or U2938 (N_2938,N_1910,N_2440);
xor U2939 (N_2939,N_775,N_790);
or U2940 (N_2940,N_890,N_2145);
nor U2941 (N_2941,N_438,N_2229);
or U2942 (N_2942,N_1719,N_852);
or U2943 (N_2943,N_1062,N_1736);
or U2944 (N_2944,N_2383,N_56);
xnor U2945 (N_2945,N_469,N_150);
or U2946 (N_2946,N_1421,N_899);
nor U2947 (N_2947,N_1047,N_1319);
nand U2948 (N_2948,N_171,N_1875);
nand U2949 (N_2949,N_1033,N_2058);
nand U2950 (N_2950,N_997,N_2247);
nor U2951 (N_2951,N_59,N_0);
or U2952 (N_2952,N_1543,N_2131);
or U2953 (N_2953,N_1556,N_726);
and U2954 (N_2954,N_159,N_394);
xnor U2955 (N_2955,N_1520,N_1671);
nor U2956 (N_2956,N_82,N_1115);
nand U2957 (N_2957,N_1148,N_1612);
or U2958 (N_2958,N_1576,N_1577);
or U2959 (N_2959,N_1063,N_563);
and U2960 (N_2960,N_1952,N_2472);
nor U2961 (N_2961,N_1805,N_1087);
nand U2962 (N_2962,N_2129,N_2280);
and U2963 (N_2963,N_1332,N_1861);
xor U2964 (N_2964,N_827,N_1567);
or U2965 (N_2965,N_638,N_940);
nor U2966 (N_2966,N_857,N_2429);
nand U2967 (N_2967,N_424,N_327);
or U2968 (N_2968,N_2434,N_2165);
nand U2969 (N_2969,N_1251,N_2041);
or U2970 (N_2970,N_2286,N_1480);
or U2971 (N_2971,N_1677,N_1657);
nand U2972 (N_2972,N_329,N_1869);
or U2973 (N_2973,N_1633,N_918);
nor U2974 (N_2974,N_2053,N_1166);
nand U2975 (N_2975,N_794,N_1262);
nor U2976 (N_2976,N_1441,N_748);
nor U2977 (N_2977,N_1561,N_524);
and U2978 (N_2978,N_2330,N_1494);
or U2979 (N_2979,N_1898,N_937);
nand U2980 (N_2980,N_1228,N_1669);
nand U2981 (N_2981,N_259,N_320);
and U2982 (N_2982,N_194,N_1090);
or U2983 (N_2983,N_695,N_2451);
or U2984 (N_2984,N_1842,N_2013);
nor U2985 (N_2985,N_433,N_1011);
or U2986 (N_2986,N_1850,N_298);
or U2987 (N_2987,N_1235,N_2491);
or U2988 (N_2988,N_904,N_703);
or U2989 (N_2989,N_1962,N_1990);
or U2990 (N_2990,N_658,N_839);
and U2991 (N_2991,N_644,N_69);
or U2992 (N_2992,N_855,N_271);
nand U2993 (N_2993,N_184,N_2010);
and U2994 (N_2994,N_1751,N_58);
nand U2995 (N_2995,N_2327,N_135);
and U2996 (N_2996,N_444,N_1140);
and U2997 (N_2997,N_2067,N_1057);
nand U2998 (N_2998,N_1318,N_819);
xnor U2999 (N_2999,N_2461,N_876);
or U3000 (N_3000,N_1430,N_411);
nor U3001 (N_3001,N_500,N_64);
nor U3002 (N_3002,N_1539,N_250);
nor U3003 (N_3003,N_2152,N_2314);
and U3004 (N_3004,N_1806,N_308);
or U3005 (N_3005,N_729,N_758);
nand U3006 (N_3006,N_1885,N_2389);
nand U3007 (N_3007,N_2379,N_65);
nor U3008 (N_3008,N_1972,N_113);
and U3009 (N_3009,N_992,N_496);
nand U3010 (N_3010,N_280,N_1443);
xor U3011 (N_3011,N_1704,N_1607);
or U3012 (N_3012,N_1967,N_1104);
nor U3013 (N_3013,N_515,N_1579);
nand U3014 (N_3014,N_1993,N_147);
or U3015 (N_3015,N_395,N_666);
nor U3016 (N_3016,N_647,N_2195);
nor U3017 (N_3017,N_239,N_1985);
nand U3018 (N_3018,N_2415,N_1882);
and U3019 (N_3019,N_1672,N_222);
or U3020 (N_3020,N_1939,N_693);
nand U3021 (N_3021,N_436,N_124);
nand U3022 (N_3022,N_1776,N_1197);
or U3023 (N_3023,N_1173,N_2218);
or U3024 (N_3024,N_1268,N_1868);
nand U3025 (N_3025,N_1149,N_2005);
nand U3026 (N_3026,N_1799,N_1562);
nor U3027 (N_3027,N_1081,N_682);
nor U3028 (N_3028,N_616,N_2320);
nand U3029 (N_3029,N_1462,N_1936);
or U3030 (N_3030,N_537,N_1093);
or U3031 (N_3031,N_591,N_1215);
xnor U3032 (N_3032,N_1472,N_106);
or U3033 (N_3033,N_786,N_866);
or U3034 (N_3034,N_199,N_2002);
nand U3035 (N_3035,N_2161,N_1959);
nand U3036 (N_3036,N_2272,N_576);
nand U3037 (N_3037,N_1795,N_234);
and U3038 (N_3038,N_1807,N_1517);
nor U3039 (N_3039,N_501,N_133);
and U3040 (N_3040,N_1466,N_1682);
nand U3041 (N_3041,N_1473,N_1656);
or U3042 (N_3042,N_474,N_623);
and U3043 (N_3043,N_2134,N_1930);
or U3044 (N_3044,N_2483,N_648);
nand U3045 (N_3045,N_1295,N_1478);
nand U3046 (N_3046,N_1867,N_2369);
and U3047 (N_3047,N_92,N_2368);
nor U3048 (N_3048,N_1853,N_1668);
nor U3049 (N_3049,N_995,N_281);
or U3050 (N_3050,N_1727,N_667);
and U3051 (N_3051,N_183,N_2107);
and U3052 (N_3052,N_955,N_2443);
nor U3053 (N_3053,N_634,N_1597);
nor U3054 (N_3054,N_2009,N_2174);
nor U3055 (N_3055,N_47,N_1401);
nand U3056 (N_3056,N_2457,N_2025);
nor U3057 (N_3057,N_2360,N_180);
nor U3058 (N_3058,N_1225,N_1447);
nand U3059 (N_3059,N_931,N_831);
and U3060 (N_3060,N_450,N_1879);
nand U3061 (N_3061,N_2130,N_1944);
nand U3062 (N_3062,N_529,N_2295);
and U3063 (N_3063,N_2427,N_1921);
or U3064 (N_3064,N_1613,N_2233);
and U3065 (N_3065,N_1326,N_2151);
nand U3066 (N_3066,N_2322,N_2111);
nor U3067 (N_3067,N_1172,N_2277);
and U3068 (N_3068,N_585,N_1321);
and U3069 (N_3069,N_1844,N_687);
or U3070 (N_3070,N_2414,N_1552);
or U3071 (N_3071,N_2158,N_210);
nand U3072 (N_3072,N_1356,N_157);
or U3073 (N_3073,N_62,N_1660);
xor U3074 (N_3074,N_1469,N_1434);
or U3075 (N_3075,N_2403,N_1278);
or U3076 (N_3076,N_1199,N_1455);
nand U3077 (N_3077,N_514,N_1566);
and U3078 (N_3078,N_900,N_2210);
nand U3079 (N_3079,N_745,N_228);
and U3080 (N_3080,N_321,N_152);
or U3081 (N_3081,N_1183,N_261);
nand U3082 (N_3082,N_1767,N_1114);
xor U3083 (N_3083,N_451,N_98);
xnor U3084 (N_3084,N_1377,N_1485);
nand U3085 (N_3085,N_1922,N_2432);
and U3086 (N_3086,N_1752,N_165);
or U3087 (N_3087,N_142,N_2127);
and U3088 (N_3088,N_1185,N_987);
xnor U3089 (N_3089,N_246,N_1178);
nand U3090 (N_3090,N_1788,N_1303);
or U3091 (N_3091,N_1531,N_861);
nor U3092 (N_3092,N_1541,N_1965);
and U3093 (N_3093,N_854,N_1877);
and U3094 (N_3094,N_247,N_2387);
and U3095 (N_3095,N_1629,N_863);
and U3096 (N_3096,N_1715,N_2267);
nor U3097 (N_3097,N_642,N_999);
nand U3098 (N_3098,N_1241,N_1524);
and U3099 (N_3099,N_516,N_1575);
or U3100 (N_3100,N_375,N_604);
nor U3101 (N_3101,N_1847,N_1248);
or U3102 (N_3102,N_1399,N_823);
nand U3103 (N_3103,N_391,N_1652);
or U3104 (N_3104,N_935,N_1522);
nand U3105 (N_3105,N_672,N_1182);
or U3106 (N_3106,N_739,N_208);
nor U3107 (N_3107,N_2008,N_1221);
or U3108 (N_3108,N_2100,N_914);
xnor U3109 (N_3109,N_1865,N_1438);
or U3110 (N_3110,N_572,N_1368);
nor U3111 (N_3111,N_665,N_829);
or U3112 (N_3112,N_189,N_1721);
and U3113 (N_3113,N_523,N_303);
xor U3114 (N_3114,N_2437,N_1055);
and U3115 (N_3115,N_1744,N_938);
or U3116 (N_3116,N_1620,N_1310);
or U3117 (N_3117,N_1271,N_661);
nand U3118 (N_3118,N_1342,N_1073);
nand U3119 (N_3119,N_1042,N_535);
nand U3120 (N_3120,N_2462,N_2467);
nand U3121 (N_3121,N_1887,N_1431);
nand U3122 (N_3122,N_1453,N_128);
nand U3123 (N_3123,N_727,N_2222);
or U3124 (N_3124,N_2410,N_214);
xor U3125 (N_3125,N_1133,N_916);
nor U3126 (N_3126,N_1786,N_1796);
or U3127 (N_3127,N_2227,N_1163);
and U3128 (N_3128,N_1314,N_1589);
nor U3129 (N_3129,N_1129,N_1619);
nand U3130 (N_3130,N_2422,N_2089);
xor U3131 (N_3131,N_1694,N_2043);
or U3132 (N_3132,N_936,N_1159);
nand U3133 (N_3133,N_1481,N_487);
nand U3134 (N_3134,N_1213,N_2064);
or U3135 (N_3135,N_1374,N_1246);
and U3136 (N_3136,N_129,N_800);
nand U3137 (N_3137,N_1925,N_1327);
and U3138 (N_3138,N_778,N_626);
or U3139 (N_3139,N_791,N_2421);
and U3140 (N_3140,N_1723,N_2048);
nand U3141 (N_3141,N_372,N_105);
or U3142 (N_3142,N_2000,N_2094);
or U3143 (N_3143,N_2348,N_1740);
and U3144 (N_3144,N_2208,N_2197);
xnor U3145 (N_3145,N_46,N_310);
xnor U3146 (N_3146,N_1605,N_2488);
and U3147 (N_3147,N_2426,N_1139);
xor U3148 (N_3148,N_1476,N_104);
xor U3149 (N_3149,N_455,N_2121);
nand U3150 (N_3150,N_223,N_680);
nor U3151 (N_3151,N_1006,N_1301);
or U3152 (N_3152,N_1239,N_466);
xor U3153 (N_3153,N_1280,N_629);
and U3154 (N_3154,N_2245,N_575);
and U3155 (N_3155,N_344,N_1414);
and U3156 (N_3156,N_186,N_1880);
nand U3157 (N_3157,N_1814,N_2250);
xor U3158 (N_3158,N_1244,N_673);
and U3159 (N_3159,N_1890,N_542);
or U3160 (N_3160,N_834,N_2478);
nor U3161 (N_3161,N_1307,N_2034);
or U3162 (N_3162,N_1363,N_607);
or U3163 (N_3163,N_1031,N_2300);
and U3164 (N_3164,N_832,N_1987);
or U3165 (N_3165,N_211,N_427);
xnor U3166 (N_3166,N_1069,N_2066);
nand U3167 (N_3167,N_954,N_744);
and U3168 (N_3168,N_2319,N_1168);
nor U3169 (N_3169,N_583,N_405);
xnor U3170 (N_3170,N_389,N_603);
and U3171 (N_3171,N_590,N_1608);
and U3172 (N_3172,N_435,N_2101);
nor U3173 (N_3173,N_449,N_843);
or U3174 (N_3174,N_1585,N_1145);
nand U3175 (N_3175,N_1923,N_2345);
nand U3176 (N_3176,N_1160,N_1259);
or U3177 (N_3177,N_1053,N_1554);
nor U3178 (N_3178,N_2290,N_1697);
or U3179 (N_3179,N_494,N_2262);
nand U3180 (N_3180,N_1432,N_1467);
nand U3181 (N_3181,N_766,N_177);
or U3182 (N_3182,N_773,N_1730);
nand U3183 (N_3183,N_2489,N_760);
nor U3184 (N_3184,N_1000,N_316);
nand U3185 (N_3185,N_805,N_560);
nand U3186 (N_3186,N_688,N_1708);
or U3187 (N_3187,N_1980,N_1076);
nand U3188 (N_3188,N_879,N_403);
nand U3189 (N_3189,N_1916,N_532);
and U3190 (N_3190,N_2335,N_1917);
nor U3191 (N_3191,N_95,N_1938);
nand U3192 (N_3192,N_1435,N_1125);
nand U3193 (N_3193,N_1622,N_895);
nand U3194 (N_3194,N_1222,N_216);
xnor U3195 (N_3195,N_978,N_996);
or U3196 (N_3196,N_608,N_1855);
and U3197 (N_3197,N_213,N_1445);
and U3198 (N_3198,N_7,N_207);
or U3199 (N_3199,N_1014,N_528);
nor U3200 (N_3200,N_238,N_2084);
and U3201 (N_3201,N_875,N_2498);
and U3202 (N_3202,N_720,N_546);
nor U3203 (N_3203,N_2125,N_919);
or U3204 (N_3204,N_1136,N_1763);
and U3205 (N_3205,N_2106,N_2384);
and U3206 (N_3206,N_1316,N_2296);
and U3207 (N_3207,N_1775,N_650);
and U3208 (N_3208,N_1429,N_1263);
or U3209 (N_3209,N_901,N_1240);
nor U3210 (N_3210,N_1926,N_949);
xnor U3211 (N_3211,N_2385,N_2196);
and U3212 (N_3212,N_1741,N_360);
and U3213 (N_3213,N_423,N_564);
nor U3214 (N_3214,N_2054,N_385);
nand U3215 (N_3215,N_283,N_574);
or U3216 (N_3216,N_1287,N_2198);
xor U3217 (N_3217,N_2016,N_691);
or U3218 (N_3218,N_1785,N_2378);
or U3219 (N_3219,N_457,N_274);
and U3220 (N_3220,N_587,N_1091);
nor U3221 (N_3221,N_1074,N_2037);
and U3222 (N_3222,N_1529,N_1085);
and U3223 (N_3223,N_431,N_1344);
and U3224 (N_3224,N_1212,N_1848);
nand U3225 (N_3225,N_718,N_878);
nor U3226 (N_3226,N_1718,N_676);
or U3227 (N_3227,N_1511,N_934);
and U3228 (N_3228,N_1737,N_2139);
nand U3229 (N_3229,N_1020,N_520);
or U3230 (N_3230,N_1357,N_2112);
nor U3231 (N_3231,N_2033,N_620);
nor U3232 (N_3232,N_2490,N_1315);
nand U3233 (N_3233,N_358,N_290);
xor U3234 (N_3234,N_299,N_2340);
or U3235 (N_3235,N_783,N_1498);
nor U3236 (N_3236,N_873,N_209);
and U3237 (N_3237,N_2494,N_2235);
or U3238 (N_3238,N_1150,N_1547);
or U3239 (N_3239,N_538,N_160);
nor U3240 (N_3240,N_1611,N_925);
and U3241 (N_3241,N_923,N_432);
nor U3242 (N_3242,N_2497,N_1218);
or U3243 (N_3243,N_1,N_2470);
and U3244 (N_3244,N_1041,N_2022);
nand U3245 (N_3245,N_251,N_397);
or U3246 (N_3246,N_2362,N_472);
and U3247 (N_3247,N_1079,N_1233);
or U3248 (N_3248,N_1774,N_1156);
or U3249 (N_3249,N_2234,N_660);
and U3250 (N_3250,N_1873,N_637);
and U3251 (N_3251,N_1852,N_2318);
or U3252 (N_3252,N_179,N_2452);
nand U3253 (N_3253,N_2438,N_1978);
and U3254 (N_3254,N_1061,N_1667);
and U3255 (N_3255,N_326,N_2419);
or U3256 (N_3256,N_2264,N_1143);
nor U3257 (N_3257,N_401,N_2418);
nand U3258 (N_3258,N_2028,N_701);
xor U3259 (N_3259,N_2007,N_443);
and U3260 (N_3260,N_1523,N_699);
and U3261 (N_3261,N_224,N_592);
nor U3262 (N_3262,N_2275,N_1725);
or U3263 (N_3263,N_1490,N_1900);
or U3264 (N_3264,N_1699,N_252);
and U3265 (N_3265,N_1907,N_86);
or U3266 (N_3266,N_1302,N_2380);
nand U3267 (N_3267,N_380,N_1038);
or U3268 (N_3268,N_1754,N_1684);
and U3269 (N_3269,N_178,N_725);
xnor U3270 (N_3270,N_508,N_145);
nand U3271 (N_3271,N_631,N_1293);
and U3272 (N_3272,N_605,N_2086);
nor U3273 (N_3273,N_1791,N_1902);
nand U3274 (N_3274,N_844,N_2287);
or U3275 (N_3275,N_428,N_2074);
nor U3276 (N_3276,N_1487,N_787);
nand U3277 (N_3277,N_151,N_2400);
and U3278 (N_3278,N_698,N_413);
nor U3279 (N_3279,N_2271,N_1832);
and U3280 (N_3280,N_1929,N_217);
nor U3281 (N_3281,N_2409,N_840);
or U3282 (N_3282,N_2450,N_2103);
nor U3283 (N_3283,N_18,N_485);
nand U3284 (N_3284,N_1175,N_315);
xnor U3285 (N_3285,N_73,N_504);
nor U3286 (N_3286,N_2189,N_1442);
or U3287 (N_3287,N_1630,N_1100);
nand U3288 (N_3288,N_1030,N_2424);
and U3289 (N_3289,N_2458,N_842);
or U3290 (N_3290,N_1317,N_1527);
and U3291 (N_3291,N_1731,N_2281);
and U3292 (N_3292,N_659,N_617);
and U3293 (N_3293,N_1015,N_2313);
and U3294 (N_3294,N_2202,N_168);
xor U3295 (N_3295,N_1007,N_1747);
nor U3296 (N_3296,N_770,N_2068);
nor U3297 (N_3297,N_1346,N_871);
or U3298 (N_3298,N_1695,N_1347);
and U3299 (N_3299,N_1164,N_920);
xnor U3300 (N_3300,N_2040,N_2001);
nand U3301 (N_3301,N_410,N_599);
or U3302 (N_3302,N_396,N_1894);
or U3303 (N_3303,N_1881,N_1194);
or U3304 (N_3304,N_1545,N_1255);
or U3305 (N_3305,N_513,N_811);
or U3306 (N_3306,N_90,N_779);
and U3307 (N_3307,N_1456,N_51);
nand U3308 (N_3308,N_2206,N_1387);
nand U3309 (N_3309,N_969,N_33);
or U3310 (N_3310,N_1988,N_266);
nor U3311 (N_3311,N_67,N_1340);
or U3312 (N_3312,N_1083,N_1911);
xnor U3313 (N_3313,N_453,N_717);
and U3314 (N_3314,N_816,N_1606);
and U3315 (N_3315,N_1366,N_2060);
nor U3316 (N_3316,N_1174,N_1184);
nand U3317 (N_3317,N_1392,N_1693);
and U3318 (N_3318,N_1689,N_956);
and U3319 (N_3319,N_1771,N_2289);
nor U3320 (N_3320,N_497,N_2276);
and U3321 (N_3321,N_749,N_80);
and U3322 (N_3322,N_1292,N_865);
and U3323 (N_3323,N_1113,N_2445);
or U3324 (N_3324,N_467,N_1661);
xor U3325 (N_3325,N_1768,N_1407);
nand U3326 (N_3326,N_2019,N_1617);
or U3327 (N_3327,N_1207,N_1142);
or U3328 (N_3328,N_1032,N_1046);
nor U3329 (N_3329,N_378,N_927);
or U3330 (N_3330,N_671,N_161);
or U3331 (N_3331,N_1109,N_611);
or U3332 (N_3332,N_1632,N_1958);
or U3333 (N_3333,N_1705,N_1587);
nand U3334 (N_3334,N_1948,N_2248);
nor U3335 (N_3335,N_2312,N_2413);
nand U3336 (N_3336,N_2128,N_700);
or U3337 (N_3337,N_1258,N_2388);
nand U3338 (N_3338,N_318,N_305);
and U3339 (N_3339,N_418,N_1665);
or U3340 (N_3340,N_243,N_1569);
nor U3341 (N_3341,N_61,N_1874);
and U3342 (N_3342,N_190,N_1638);
or U3343 (N_3343,N_434,N_1841);
nor U3344 (N_3344,N_1979,N_2252);
or U3345 (N_3345,N_363,N_1537);
nor U3346 (N_3346,N_2428,N_354);
xor U3347 (N_3347,N_1223,N_448);
and U3348 (N_3348,N_1023,N_1749);
nor U3349 (N_3349,N_941,N_527);
or U3350 (N_3350,N_627,N_1275);
and U3351 (N_3351,N_2230,N_37);
and U3352 (N_3352,N_1914,N_853);
and U3353 (N_3353,N_1756,N_2029);
or U3354 (N_3354,N_1809,N_89);
and U3355 (N_3355,N_1982,N_1337);
and U3356 (N_3356,N_817,N_1479);
or U3357 (N_3357,N_828,N_1870);
and U3358 (N_3358,N_1743,N_235);
nor U3359 (N_3359,N_1935,N_1035);
nor U3360 (N_3360,N_2123,N_1506);
or U3361 (N_3361,N_589,N_1127);
and U3362 (N_3362,N_1477,N_1974);
or U3363 (N_3363,N_1654,N_75);
nor U3364 (N_3364,N_130,N_2328);
and U3365 (N_3365,N_286,N_970);
xor U3366 (N_3366,N_1780,N_1489);
nor U3367 (N_3367,N_849,N_1350);
xnor U3368 (N_3368,N_341,N_1849);
and U3369 (N_3369,N_1450,N_1354);
nand U3370 (N_3370,N_30,N_503);
and U3371 (N_3371,N_1131,N_908);
nor U3372 (N_3372,N_517,N_2180);
nand U3373 (N_3373,N_1808,N_1224);
nor U3374 (N_3374,N_1878,N_1564);
nor U3375 (N_3375,N_685,N_1572);
or U3376 (N_3376,N_2326,N_1176);
and U3377 (N_3377,N_1750,N_2232);
nand U3378 (N_3378,N_201,N_1729);
nand U3379 (N_3379,N_2406,N_2254);
nand U3380 (N_3380,N_540,N_841);
xnor U3381 (N_3381,N_968,N_2473);
and U3382 (N_3382,N_357,N_1082);
and U3383 (N_3383,N_722,N_803);
nor U3384 (N_3384,N_1679,N_1794);
nand U3385 (N_3385,N_848,N_53);
and U3386 (N_3386,N_116,N_2015);
and U3387 (N_3387,N_265,N_2407);
nand U3388 (N_3388,N_2279,N_131);
nand U3389 (N_3389,N_1250,N_215);
nor U3390 (N_3390,N_798,N_1274);
nor U3391 (N_3391,N_1532,N_2394);
nor U3392 (N_3392,N_307,N_910);
and U3393 (N_3393,N_1766,N_1027);
nand U3394 (N_3394,N_1124,N_390);
xor U3395 (N_3395,N_1284,N_1308);
nor U3396 (N_3396,N_559,N_772);
nand U3397 (N_3397,N_915,N_203);
and U3398 (N_3398,N_109,N_612);
nor U3399 (N_3399,N_593,N_376);
or U3400 (N_3400,N_981,N_2463);
or U3401 (N_3401,N_2482,N_913);
nand U3402 (N_3402,N_1977,N_1513);
nand U3403 (N_3403,N_534,N_2291);
and U3404 (N_3404,N_1761,N_721);
nor U3405 (N_3405,N_475,N_2408);
nand U3406 (N_3406,N_903,N_1493);
nor U3407 (N_3407,N_569,N_1098);
nor U3408 (N_3408,N_856,N_2070);
or U3409 (N_3409,N_2344,N_1092);
and U3410 (N_3410,N_1181,N_670);
xor U3411 (N_3411,N_1375,N_1217);
and U3412 (N_3412,N_48,N_1904);
nand U3413 (N_3413,N_1801,N_732);
nand U3414 (N_3414,N_581,N_1720);
or U3415 (N_3415,N_692,N_1586);
or U3416 (N_3416,N_1864,N_1666);
and U3417 (N_3417,N_21,N_478);
nand U3418 (N_3418,N_2361,N_2144);
and U3419 (N_3419,N_907,N_153);
nor U3420 (N_3420,N_1265,N_2237);
and U3421 (N_3421,N_1003,N_580);
and U3422 (N_3422,N_929,N_425);
nor U3423 (N_3423,N_406,N_1242);
or U3424 (N_3424,N_1192,N_1670);
nor U3425 (N_3425,N_902,N_1475);
or U3426 (N_3426,N_2273,N_1709);
and U3427 (N_3427,N_39,N_645);
nor U3428 (N_3428,N_1581,N_862);
xnor U3429 (N_3429,N_163,N_2078);
xnor U3430 (N_3430,N_1026,N_690);
nand U3431 (N_3431,N_233,N_442);
xnor U3432 (N_3432,N_1465,N_1457);
and U3433 (N_3433,N_1896,N_2228);
nand U3434 (N_3434,N_268,N_471);
nand U3435 (N_3435,N_1048,N_957);
and U3436 (N_3436,N_402,N_1379);
or U3437 (N_3437,N_1680,N_1823);
nand U3438 (N_3438,N_291,N_2354);
and U3439 (N_3439,N_697,N_1141);
and U3440 (N_3440,N_975,N_1676);
nor U3441 (N_3441,N_562,N_2177);
nor U3442 (N_3442,N_2214,N_114);
nand U3443 (N_3443,N_221,N_1956);
nor U3444 (N_3444,N_1783,N_1690);
xnor U3445 (N_3445,N_621,N_1019);
nor U3446 (N_3446,N_1427,N_2020);
nor U3447 (N_3447,N_1381,N_1843);
and U3448 (N_3448,N_1897,N_1883);
nor U3449 (N_3449,N_14,N_2076);
or U3450 (N_3450,N_1297,N_1779);
or U3451 (N_3451,N_825,N_1309);
nor U3452 (N_3452,N_392,N_2343);
xor U3453 (N_3453,N_1838,N_1784);
nor U3454 (N_3454,N_275,N_1002);
nor U3455 (N_3455,N_1300,N_2285);
nor U3456 (N_3456,N_136,N_555);
nor U3457 (N_3457,N_166,N_1659);
or U3458 (N_3458,N_619,N_1005);
nor U3459 (N_3459,N_383,N_470);
or U3460 (N_3460,N_1596,N_1146);
nand U3461 (N_3461,N_1336,N_664);
nor U3462 (N_3462,N_763,N_77);
nand U3463 (N_3463,N_1247,N_880);
nor U3464 (N_3464,N_761,N_1001);
and U3465 (N_3465,N_1111,N_1793);
nor U3466 (N_3466,N_2430,N_2475);
nand U3467 (N_3467,N_84,N_440);
nor U3468 (N_3468,N_896,N_1650);
or U3469 (N_3469,N_663,N_1458);
or U3470 (N_3470,N_651,N_1711);
nor U3471 (N_3471,N_42,N_872);
or U3472 (N_3472,N_493,N_1503);
nor U3473 (N_3473,N_1701,N_776);
nor U3474 (N_3474,N_1167,N_652);
nand U3475 (N_3475,N_884,N_2372);
nor U3476 (N_3476,N_2481,N_1152);
and U3477 (N_3477,N_1640,N_172);
nor U3478 (N_3478,N_1191,N_734);
nand U3479 (N_3479,N_1837,N_1811);
nand U3480 (N_3480,N_921,N_1009);
or U3481 (N_3481,N_1086,N_1460);
or U3482 (N_3482,N_570,N_1862);
or U3483 (N_3483,N_1070,N_2499);
nand U3484 (N_3484,N_1542,N_2246);
or U3485 (N_3485,N_2213,N_70);
or U3486 (N_3486,N_447,N_2104);
and U3487 (N_3487,N_2093,N_1673);
nor U3488 (N_3488,N_1204,N_1334);
nand U3489 (N_3489,N_1983,N_2417);
and U3490 (N_3490,N_1507,N_905);
or U3491 (N_3491,N_2035,N_1436);
or U3492 (N_3492,N_847,N_972);
nor U3493 (N_3493,N_1969,N_716);
and U3494 (N_3494,N_552,N_1452);
and U3495 (N_3495,N_1230,N_43);
nand U3496 (N_3496,N_1403,N_746);
nand U3497 (N_3497,N_656,N_134);
and U3498 (N_3498,N_1138,N_889);
nand U3499 (N_3499,N_2163,N_2175);
or U3500 (N_3500,N_459,N_1510);
nand U3501 (N_3501,N_25,N_1254);
or U3502 (N_3502,N_1549,N_1285);
and U3503 (N_3503,N_1961,N_465);
nor U3504 (N_3504,N_1426,N_386);
nor U3505 (N_3505,N_781,N_1078);
nor U3506 (N_3506,N_339,N_814);
or U3507 (N_3507,N_596,N_1616);
nor U3508 (N_3508,N_944,N_2032);
or U3509 (N_3509,N_355,N_1976);
and U3510 (N_3510,N_1953,N_351);
or U3511 (N_3511,N_241,N_342);
nand U3512 (N_3512,N_1835,N_989);
nor U3513 (N_3513,N_1973,N_1580);
or U3514 (N_3514,N_486,N_1203);
nor U3515 (N_3515,N_244,N_1521);
nand U3516 (N_3516,N_807,N_2225);
nor U3517 (N_3517,N_2044,N_1710);
or U3518 (N_3518,N_2185,N_195);
xor U3519 (N_3519,N_2269,N_1252);
nand U3520 (N_3520,N_2171,N_1918);
nor U3521 (N_3521,N_1828,N_518);
nor U3522 (N_3522,N_2308,N_1653);
or U3523 (N_3523,N_1833,N_1449);
nand U3524 (N_3524,N_2454,N_2143);
and U3525 (N_3525,N_804,N_419);
and U3526 (N_3526,N_1396,N_512);
nand U3527 (N_3527,N_2299,N_1385);
nor U3528 (N_3528,N_492,N_1943);
and U3529 (N_3529,N_837,N_112);
nor U3530 (N_3530,N_2017,N_156);
and U3531 (N_3531,N_737,N_2136);
or U3532 (N_3532,N_1538,N_191);
nand U3533 (N_3533,N_1981,N_640);
nand U3534 (N_3534,N_2221,N_2455);
nand U3535 (N_3535,N_2138,N_622);
and U3536 (N_3536,N_2091,N_824);
xor U3537 (N_3537,N_416,N_1826);
nor U3538 (N_3538,N_556,N_2205);
nand U3539 (N_3539,N_31,N_1348);
nand U3540 (N_3540,N_550,N_1211);
nand U3541 (N_3541,N_1871,N_1051);
or U3542 (N_3542,N_1064,N_422);
xor U3543 (N_3543,N_630,N_2258);
nand U3544 (N_3544,N_568,N_20);
xor U3545 (N_3545,N_2236,N_799);
and U3546 (N_3546,N_2338,N_2172);
and U3547 (N_3547,N_1884,N_123);
or U3548 (N_3548,N_2088,N_1400);
or U3549 (N_3549,N_724,N_1759);
nor U3550 (N_3550,N_2405,N_764);
or U3551 (N_3551,N_2169,N_1599);
and U3552 (N_3552,N_548,N_2072);
or U3553 (N_3553,N_649,N_356);
or U3554 (N_3554,N_526,N_1162);
nor U3555 (N_3555,N_2392,N_257);
or U3556 (N_3556,N_768,N_1198);
xor U3557 (N_3557,N_32,N_1158);
nor U3558 (N_3558,N_1889,N_2063);
or U3559 (N_3559,N_990,N_1931);
nor U3560 (N_3560,N_1355,N_845);
and U3561 (N_3561,N_1906,N_1107);
nand U3562 (N_3562,N_187,N_553);
nand U3563 (N_3563,N_1187,N_960);
and U3564 (N_3564,N_1446,N_1075);
and U3565 (N_3565,N_2259,N_1591);
or U3566 (N_3566,N_398,N_1582);
or U3567 (N_3567,N_982,N_1153);
and U3568 (N_3568,N_1132,N_2049);
nor U3569 (N_3569,N_1994,N_2260);
and U3570 (N_3570,N_1570,N_1940);
nor U3571 (N_3571,N_1261,N_1068);
and U3572 (N_3572,N_646,N_1195);
or U3573 (N_3573,N_826,N_417);
nor U3574 (N_3574,N_2141,N_909);
nor U3575 (N_3575,N_52,N_2087);
or U3576 (N_3576,N_240,N_2244);
nand U3577 (N_3577,N_2386,N_1675);
xnor U3578 (N_3578,N_1755,N_317);
or U3579 (N_3579,N_922,N_2099);
or U3580 (N_3580,N_963,N_2004);
or U3581 (N_3581,N_1655,N_893);
and U3582 (N_3582,N_1080,N_2132);
nor U3583 (N_3583,N_445,N_1238);
xnor U3584 (N_3584,N_1119,N_1647);
nor U3585 (N_3585,N_169,N_242);
and U3586 (N_3586,N_2109,N_1816);
or U3587 (N_3587,N_813,N_769);
nand U3588 (N_3588,N_1592,N_1615);
nand U3589 (N_3589,N_1220,N_1627);
or U3590 (N_3590,N_723,N_1700);
nor U3591 (N_3591,N_681,N_154);
nor U3592 (N_3592,N_874,N_1202);
nand U3593 (N_3593,N_609,N_933);
xnor U3594 (N_3594,N_2448,N_2026);
or U3595 (N_3595,N_489,N_108);
nand U3596 (N_3596,N_99,N_1932);
or U3597 (N_3597,N_809,N_888);
nor U3598 (N_3598,N_162,N_2073);
nor U3599 (N_3599,N_117,N_1574);
nor U3600 (N_3600,N_806,N_1643);
nor U3601 (N_3601,N_1306,N_2238);
or U3602 (N_3602,N_980,N_2110);
or U3603 (N_3603,N_226,N_719);
nand U3604 (N_3604,N_530,N_2464);
and U3605 (N_3605,N_1289,N_155);
and U3606 (N_3606,N_322,N_662);
nand U3607 (N_3607,N_2142,N_1413);
and U3608 (N_3608,N_891,N_1971);
and U3609 (N_3609,N_859,N_2359);
and U3610 (N_3610,N_364,N_771);
nand U3611 (N_3611,N_2292,N_2184);
nand U3612 (N_3612,N_2471,N_1583);
xor U3613 (N_3613,N_2122,N_479);
xnor U3614 (N_3614,N_1565,N_2365);
and U3615 (N_3615,N_1765,N_306);
nor U3616 (N_3616,N_495,N_1621);
nand U3617 (N_3617,N_1770,N_2342);
or U3618 (N_3618,N_285,N_1398);
and U3619 (N_3619,N_808,N_2240);
or U3620 (N_3620,N_1341,N_2283);
nor U3621 (N_3621,N_324,N_1231);
nor U3622 (N_3622,N_200,N_1909);
or U3623 (N_3623,N_1526,N_125);
and U3624 (N_3624,N_1732,N_1040);
nand U3625 (N_3625,N_2012,N_2381);
nor U3626 (N_3626,N_1406,N_2373);
and U3627 (N_3627,N_2261,N_293);
nor U3628 (N_3628,N_1933,N_2495);
and U3629 (N_3629,N_998,N_983);
or U3630 (N_3630,N_2278,N_1428);
xor U3631 (N_3631,N_2056,N_539);
nand U3632 (N_3632,N_132,N_2051);
nand U3633 (N_3633,N_1519,N_193);
or U3634 (N_3634,N_141,N_2453);
xor U3635 (N_3635,N_1571,N_225);
nor U3636 (N_3636,N_924,N_509);
or U3637 (N_3637,N_1899,N_2447);
and U3638 (N_3638,N_340,N_2166);
nor U3639 (N_3639,N_710,N_511);
nor U3640 (N_3640,N_733,N_1748);
nor U3641 (N_3641,N_50,N_705);
nand U3642 (N_3642,N_1471,N_2137);
nor U3643 (N_3643,N_2157,N_1171);
nor U3644 (N_3644,N_174,N_1017);
nor U3645 (N_3645,N_2334,N_236);
nand U3646 (N_3646,N_838,N_1330);
nor U3647 (N_3647,N_2203,N_1039);
or U3648 (N_3648,N_549,N_1845);
xnor U3649 (N_3649,N_2047,N_551);
and U3650 (N_3650,N_1812,N_1815);
nor U3651 (N_3651,N_1762,N_1839);
and U3652 (N_3652,N_1960,N_1294);
or U3653 (N_3653,N_1094,N_1170);
or U3654 (N_3654,N_598,N_951);
and U3655 (N_3655,N_1734,N_1488);
nand U3656 (N_3656,N_2042,N_1054);
or U3657 (N_3657,N_2492,N_1474);
and U3658 (N_3658,N_1745,N_2150);
nand U3659 (N_3659,N_439,N_1352);
nor U3660 (N_3660,N_1664,N_1118);
nand U3661 (N_3661,N_333,N_2147);
nor U3662 (N_3662,N_2435,N_668);
and U3663 (N_3663,N_126,N_6);
nand U3664 (N_3664,N_1912,N_1685);
and U3665 (N_3665,N_1378,N_13);
nand U3666 (N_3666,N_1328,N_1728);
nand U3667 (N_3667,N_588,N_1886);
and U3668 (N_3668,N_1989,N_1703);
or U3669 (N_3669,N_1050,N_1043);
nor U3670 (N_3670,N_1016,N_1117);
nor U3671 (N_3671,N_1614,N_1361);
nor U3672 (N_3672,N_28,N_2352);
nor U3673 (N_3673,N_1834,N_1422);
and U3674 (N_3674,N_1012,N_1905);
nor U3675 (N_3675,N_1433,N_1492);
nor U3676 (N_3676,N_1169,N_2183);
or U3677 (N_3677,N_777,N_1733);
nand U3678 (N_3678,N_1482,N_2039);
and U3679 (N_3679,N_1229,N_2113);
nand U3680 (N_3680,N_2412,N_1530);
and U3681 (N_3681,N_343,N_2212);
nor U3682 (N_3682,N_110,N_1226);
nand U3683 (N_3683,N_926,N_1232);
or U3684 (N_3684,N_1036,N_784);
nor U3685 (N_3685,N_34,N_331);
and U3686 (N_3686,N_26,N_1108);
or U3687 (N_3687,N_2181,N_1404);
or U3688 (N_3688,N_2370,N_2493);
and U3689 (N_3689,N_1598,N_1112);
or U3690 (N_3690,N_1998,N_2201);
nand U3691 (N_3691,N_1518,N_1891);
nand U3692 (N_3692,N_1272,N_1388);
xnor U3693 (N_3693,N_973,N_337);
or U3694 (N_3694,N_2356,N_1984);
and U3695 (N_3695,N_2366,N_1831);
and U3696 (N_3696,N_2346,N_368);
and U3697 (N_3697,N_1424,N_2083);
or U3698 (N_3698,N_2090,N_111);
nand U3699 (N_3699,N_2243,N_319);
and U3700 (N_3700,N_2062,N_313);
and U3701 (N_3701,N_480,N_2154);
and U3702 (N_3702,N_1698,N_81);
and U3703 (N_3703,N_40,N_967);
or U3704 (N_3704,N_1735,N_2274);
nand U3705 (N_3705,N_1237,N_868);
xor U3706 (N_3706,N_1484,N_78);
nand U3707 (N_3707,N_1777,N_414);
nand U3708 (N_3708,N_2321,N_892);
nand U3709 (N_3709,N_2351,N_932);
or U3710 (N_3710,N_1128,N_1625);
and U3711 (N_3711,N_2050,N_2402);
xnor U3712 (N_3712,N_2215,N_1362);
xnor U3713 (N_3713,N_2425,N_1856);
nand U3714 (N_3714,N_91,N_491);
nand U3715 (N_3715,N_704,N_991);
and U3716 (N_3716,N_314,N_1440);
xnor U3717 (N_3717,N_264,N_545);
nand U3718 (N_3718,N_63,N_755);
and U3719 (N_3719,N_531,N_388);
xor U3720 (N_3720,N_269,N_2178);
and U3721 (N_3721,N_463,N_2496);
nand U3722 (N_3722,N_820,N_2075);
nor U3723 (N_3723,N_170,N_68);
and U3724 (N_3724,N_1637,N_1963);
nand U3725 (N_3725,N_1483,N_15);
nand U3726 (N_3726,N_2077,N_1305);
nand U3727 (N_3727,N_5,N_2116);
and U3728 (N_3728,N_1059,N_2098);
nor U3729 (N_3729,N_2102,N_1609);
or U3730 (N_3730,N_1954,N_684);
or U3731 (N_3731,N_747,N_1402);
nor U3732 (N_3732,N_362,N_338);
nand U3733 (N_3733,N_1802,N_1193);
and U3734 (N_3734,N_2355,N_45);
nand U3735 (N_3735,N_1367,N_1004);
nand U3736 (N_3736,N_12,N_669);
or U3737 (N_3737,N_2420,N_1497);
or U3738 (N_3738,N_1065,N_96);
or U3739 (N_3739,N_1338,N_412);
nand U3740 (N_3740,N_415,N_835);
nor U3741 (N_3741,N_1824,N_404);
nor U3742 (N_3742,N_928,N_27);
nand U3743 (N_3743,N_345,N_1555);
and U3744 (N_3744,N_1789,N_36);
and U3745 (N_3745,N_17,N_1196);
or U3746 (N_3746,N_158,N_979);
and U3747 (N_3747,N_614,N_1830);
or U3748 (N_3748,N_9,N_1437);
or U3749 (N_3749,N_278,N_1688);
xnor U3750 (N_3750,N_951,N_1218);
or U3751 (N_3751,N_1533,N_845);
nand U3752 (N_3752,N_1911,N_1009);
nand U3753 (N_3753,N_1021,N_2327);
and U3754 (N_3754,N_353,N_1644);
and U3755 (N_3755,N_2492,N_503);
nor U3756 (N_3756,N_1627,N_2450);
nor U3757 (N_3757,N_688,N_1091);
xor U3758 (N_3758,N_1450,N_2116);
xor U3759 (N_3759,N_1831,N_761);
nand U3760 (N_3760,N_1246,N_2086);
xor U3761 (N_3761,N_62,N_607);
or U3762 (N_3762,N_2331,N_775);
nor U3763 (N_3763,N_686,N_139);
nand U3764 (N_3764,N_991,N_514);
or U3765 (N_3765,N_2408,N_1864);
and U3766 (N_3766,N_2467,N_1771);
and U3767 (N_3767,N_662,N_1934);
nor U3768 (N_3768,N_2422,N_2072);
and U3769 (N_3769,N_100,N_999);
nor U3770 (N_3770,N_729,N_2129);
or U3771 (N_3771,N_2258,N_614);
nor U3772 (N_3772,N_99,N_1867);
or U3773 (N_3773,N_1418,N_1208);
and U3774 (N_3774,N_100,N_1202);
or U3775 (N_3775,N_1862,N_2219);
nor U3776 (N_3776,N_1675,N_769);
and U3777 (N_3777,N_1224,N_1774);
nor U3778 (N_3778,N_1008,N_526);
nand U3779 (N_3779,N_188,N_1350);
and U3780 (N_3780,N_2384,N_1573);
nor U3781 (N_3781,N_2426,N_690);
nand U3782 (N_3782,N_393,N_2348);
xor U3783 (N_3783,N_1948,N_464);
or U3784 (N_3784,N_1659,N_1109);
and U3785 (N_3785,N_1675,N_885);
nand U3786 (N_3786,N_340,N_1420);
xnor U3787 (N_3787,N_1976,N_1393);
nor U3788 (N_3788,N_1995,N_2295);
or U3789 (N_3789,N_1252,N_138);
nor U3790 (N_3790,N_228,N_1360);
nand U3791 (N_3791,N_6,N_367);
nor U3792 (N_3792,N_421,N_1914);
or U3793 (N_3793,N_917,N_524);
nand U3794 (N_3794,N_1159,N_2140);
or U3795 (N_3795,N_1217,N_123);
nor U3796 (N_3796,N_1148,N_117);
nand U3797 (N_3797,N_995,N_1001);
nor U3798 (N_3798,N_2188,N_1519);
nor U3799 (N_3799,N_1225,N_2120);
or U3800 (N_3800,N_1337,N_1209);
or U3801 (N_3801,N_410,N_1544);
and U3802 (N_3802,N_1765,N_1488);
or U3803 (N_3803,N_2442,N_529);
or U3804 (N_3804,N_2122,N_2088);
nand U3805 (N_3805,N_1346,N_2453);
nor U3806 (N_3806,N_1837,N_1433);
nor U3807 (N_3807,N_2358,N_144);
xor U3808 (N_3808,N_2272,N_1566);
or U3809 (N_3809,N_7,N_1854);
or U3810 (N_3810,N_782,N_956);
or U3811 (N_3811,N_212,N_2448);
and U3812 (N_3812,N_1786,N_24);
and U3813 (N_3813,N_237,N_2480);
and U3814 (N_3814,N_1566,N_269);
or U3815 (N_3815,N_2086,N_801);
and U3816 (N_3816,N_595,N_1194);
or U3817 (N_3817,N_948,N_2324);
and U3818 (N_3818,N_622,N_2404);
nand U3819 (N_3819,N_1712,N_1729);
or U3820 (N_3820,N_2264,N_867);
xnor U3821 (N_3821,N_1672,N_2258);
and U3822 (N_3822,N_1922,N_1115);
xnor U3823 (N_3823,N_2149,N_1213);
and U3824 (N_3824,N_2291,N_498);
or U3825 (N_3825,N_2216,N_812);
and U3826 (N_3826,N_697,N_1340);
nand U3827 (N_3827,N_1153,N_1606);
nand U3828 (N_3828,N_840,N_6);
nand U3829 (N_3829,N_874,N_392);
nor U3830 (N_3830,N_673,N_946);
or U3831 (N_3831,N_1186,N_2403);
nor U3832 (N_3832,N_1086,N_605);
and U3833 (N_3833,N_486,N_2290);
or U3834 (N_3834,N_1639,N_1943);
xnor U3835 (N_3835,N_450,N_1385);
and U3836 (N_3836,N_1987,N_1971);
and U3837 (N_3837,N_717,N_1512);
or U3838 (N_3838,N_1366,N_1909);
nand U3839 (N_3839,N_1855,N_2415);
and U3840 (N_3840,N_382,N_1575);
nand U3841 (N_3841,N_1214,N_1758);
nand U3842 (N_3842,N_2024,N_2299);
or U3843 (N_3843,N_2052,N_396);
nor U3844 (N_3844,N_1393,N_2156);
xor U3845 (N_3845,N_453,N_1714);
and U3846 (N_3846,N_863,N_618);
or U3847 (N_3847,N_616,N_1812);
or U3848 (N_3848,N_1773,N_1226);
or U3849 (N_3849,N_1602,N_622);
or U3850 (N_3850,N_2168,N_1574);
nor U3851 (N_3851,N_1330,N_718);
or U3852 (N_3852,N_2115,N_1143);
xnor U3853 (N_3853,N_494,N_918);
and U3854 (N_3854,N_267,N_1116);
or U3855 (N_3855,N_2268,N_687);
nand U3856 (N_3856,N_1654,N_166);
and U3857 (N_3857,N_839,N_2073);
or U3858 (N_3858,N_1482,N_530);
nor U3859 (N_3859,N_346,N_1288);
nor U3860 (N_3860,N_1518,N_2294);
nand U3861 (N_3861,N_264,N_2396);
nand U3862 (N_3862,N_2389,N_1402);
xnor U3863 (N_3863,N_1677,N_659);
and U3864 (N_3864,N_2066,N_1753);
nand U3865 (N_3865,N_1780,N_1061);
or U3866 (N_3866,N_140,N_1153);
and U3867 (N_3867,N_182,N_63);
nand U3868 (N_3868,N_2352,N_1327);
or U3869 (N_3869,N_1052,N_952);
or U3870 (N_3870,N_1,N_1403);
nor U3871 (N_3871,N_906,N_1357);
xnor U3872 (N_3872,N_2340,N_2175);
nand U3873 (N_3873,N_1240,N_2429);
nor U3874 (N_3874,N_24,N_1487);
or U3875 (N_3875,N_2191,N_1009);
and U3876 (N_3876,N_471,N_1445);
or U3877 (N_3877,N_1683,N_1883);
nor U3878 (N_3878,N_206,N_1566);
and U3879 (N_3879,N_491,N_1603);
and U3880 (N_3880,N_1451,N_735);
nand U3881 (N_3881,N_1852,N_873);
nand U3882 (N_3882,N_1629,N_1906);
nand U3883 (N_3883,N_1644,N_1268);
or U3884 (N_3884,N_1718,N_703);
or U3885 (N_3885,N_79,N_455);
and U3886 (N_3886,N_380,N_1333);
nor U3887 (N_3887,N_2419,N_1910);
and U3888 (N_3888,N_1560,N_216);
xnor U3889 (N_3889,N_938,N_803);
nand U3890 (N_3890,N_2418,N_278);
and U3891 (N_3891,N_1488,N_207);
or U3892 (N_3892,N_2080,N_2197);
nor U3893 (N_3893,N_2025,N_782);
or U3894 (N_3894,N_949,N_1279);
nor U3895 (N_3895,N_1568,N_2087);
nor U3896 (N_3896,N_2142,N_1618);
nor U3897 (N_3897,N_720,N_1788);
or U3898 (N_3898,N_1506,N_44);
or U3899 (N_3899,N_13,N_2345);
or U3900 (N_3900,N_1862,N_790);
nand U3901 (N_3901,N_291,N_1348);
or U3902 (N_3902,N_387,N_2262);
and U3903 (N_3903,N_1832,N_1396);
and U3904 (N_3904,N_2081,N_1455);
nand U3905 (N_3905,N_2103,N_1427);
xor U3906 (N_3906,N_1894,N_1446);
or U3907 (N_3907,N_1769,N_882);
and U3908 (N_3908,N_1735,N_472);
or U3909 (N_3909,N_79,N_1040);
nand U3910 (N_3910,N_2367,N_1232);
or U3911 (N_3911,N_2244,N_71);
nor U3912 (N_3912,N_1795,N_915);
xnor U3913 (N_3913,N_0,N_1070);
or U3914 (N_3914,N_1825,N_1246);
nor U3915 (N_3915,N_1469,N_1851);
nor U3916 (N_3916,N_1843,N_1489);
nor U3917 (N_3917,N_164,N_2258);
and U3918 (N_3918,N_2052,N_1631);
nor U3919 (N_3919,N_1764,N_1085);
nor U3920 (N_3920,N_311,N_1106);
nor U3921 (N_3921,N_2494,N_1524);
nand U3922 (N_3922,N_380,N_1783);
and U3923 (N_3923,N_2044,N_1831);
and U3924 (N_3924,N_2079,N_330);
or U3925 (N_3925,N_1400,N_2376);
nand U3926 (N_3926,N_65,N_1299);
and U3927 (N_3927,N_774,N_722);
nand U3928 (N_3928,N_2015,N_1260);
nor U3929 (N_3929,N_869,N_877);
or U3930 (N_3930,N_1375,N_1756);
or U3931 (N_3931,N_421,N_1754);
or U3932 (N_3932,N_117,N_2241);
nand U3933 (N_3933,N_2280,N_1044);
or U3934 (N_3934,N_850,N_2395);
or U3935 (N_3935,N_1249,N_1648);
nand U3936 (N_3936,N_2466,N_589);
nor U3937 (N_3937,N_1922,N_2067);
and U3938 (N_3938,N_289,N_2031);
or U3939 (N_3939,N_586,N_331);
xor U3940 (N_3940,N_401,N_793);
nor U3941 (N_3941,N_197,N_1310);
nand U3942 (N_3942,N_1993,N_253);
nor U3943 (N_3943,N_1508,N_1768);
nor U3944 (N_3944,N_1901,N_492);
nand U3945 (N_3945,N_1955,N_1819);
or U3946 (N_3946,N_1326,N_1559);
nand U3947 (N_3947,N_805,N_413);
nor U3948 (N_3948,N_424,N_1448);
xnor U3949 (N_3949,N_1010,N_555);
and U3950 (N_3950,N_837,N_15);
nor U3951 (N_3951,N_1559,N_1993);
nor U3952 (N_3952,N_935,N_2084);
or U3953 (N_3953,N_2488,N_1273);
or U3954 (N_3954,N_203,N_1878);
nand U3955 (N_3955,N_1676,N_1355);
or U3956 (N_3956,N_2019,N_1216);
nand U3957 (N_3957,N_620,N_1859);
xor U3958 (N_3958,N_1791,N_2043);
nor U3959 (N_3959,N_1256,N_477);
or U3960 (N_3960,N_2197,N_1407);
nor U3961 (N_3961,N_605,N_1213);
xnor U3962 (N_3962,N_595,N_1546);
nor U3963 (N_3963,N_232,N_2032);
or U3964 (N_3964,N_872,N_2214);
or U3965 (N_3965,N_1562,N_2022);
xnor U3966 (N_3966,N_1249,N_605);
or U3967 (N_3967,N_724,N_796);
or U3968 (N_3968,N_1108,N_803);
or U3969 (N_3969,N_1722,N_145);
or U3970 (N_3970,N_1248,N_1256);
xor U3971 (N_3971,N_670,N_2344);
nor U3972 (N_3972,N_1739,N_254);
or U3973 (N_3973,N_30,N_2371);
nand U3974 (N_3974,N_2272,N_503);
nor U3975 (N_3975,N_2425,N_523);
or U3976 (N_3976,N_1477,N_1710);
or U3977 (N_3977,N_1700,N_197);
and U3978 (N_3978,N_130,N_367);
nand U3979 (N_3979,N_1077,N_820);
or U3980 (N_3980,N_996,N_1832);
or U3981 (N_3981,N_336,N_1914);
nand U3982 (N_3982,N_173,N_2207);
and U3983 (N_3983,N_1292,N_634);
or U3984 (N_3984,N_449,N_1);
or U3985 (N_3985,N_1759,N_1250);
or U3986 (N_3986,N_1101,N_342);
nor U3987 (N_3987,N_685,N_1602);
nand U3988 (N_3988,N_2238,N_2189);
or U3989 (N_3989,N_2153,N_762);
nand U3990 (N_3990,N_559,N_1804);
and U3991 (N_3991,N_523,N_1608);
nor U3992 (N_3992,N_988,N_776);
nor U3993 (N_3993,N_1318,N_134);
nor U3994 (N_3994,N_2407,N_1684);
or U3995 (N_3995,N_1055,N_911);
xnor U3996 (N_3996,N_550,N_1111);
and U3997 (N_3997,N_318,N_1331);
nand U3998 (N_3998,N_2189,N_582);
and U3999 (N_3999,N_2074,N_959);
xor U4000 (N_4000,N_1668,N_806);
nand U4001 (N_4001,N_1921,N_2286);
xnor U4002 (N_4002,N_2288,N_351);
nand U4003 (N_4003,N_1892,N_1028);
or U4004 (N_4004,N_1353,N_1044);
nand U4005 (N_4005,N_471,N_1840);
nand U4006 (N_4006,N_2101,N_164);
nand U4007 (N_4007,N_1642,N_2177);
or U4008 (N_4008,N_264,N_109);
and U4009 (N_4009,N_1435,N_1647);
nand U4010 (N_4010,N_1220,N_1246);
nand U4011 (N_4011,N_2273,N_421);
and U4012 (N_4012,N_961,N_1667);
nor U4013 (N_4013,N_2311,N_2301);
nor U4014 (N_4014,N_1911,N_2265);
nor U4015 (N_4015,N_314,N_250);
nand U4016 (N_4016,N_2137,N_1574);
or U4017 (N_4017,N_2096,N_2306);
or U4018 (N_4018,N_1118,N_2267);
nor U4019 (N_4019,N_1952,N_2165);
nand U4020 (N_4020,N_2391,N_1106);
and U4021 (N_4021,N_169,N_1102);
nor U4022 (N_4022,N_2270,N_1182);
or U4023 (N_4023,N_871,N_185);
and U4024 (N_4024,N_724,N_1388);
and U4025 (N_4025,N_993,N_1306);
nand U4026 (N_4026,N_221,N_1187);
nor U4027 (N_4027,N_2422,N_398);
or U4028 (N_4028,N_1890,N_1952);
and U4029 (N_4029,N_144,N_758);
or U4030 (N_4030,N_2282,N_1296);
and U4031 (N_4031,N_650,N_434);
nand U4032 (N_4032,N_2431,N_629);
or U4033 (N_4033,N_949,N_1605);
nand U4034 (N_4034,N_477,N_436);
or U4035 (N_4035,N_642,N_939);
nor U4036 (N_4036,N_976,N_286);
or U4037 (N_4037,N_217,N_1089);
nand U4038 (N_4038,N_516,N_1661);
nor U4039 (N_4039,N_685,N_1130);
and U4040 (N_4040,N_1297,N_2169);
nand U4041 (N_4041,N_1795,N_1197);
nand U4042 (N_4042,N_2092,N_252);
xor U4043 (N_4043,N_356,N_29);
or U4044 (N_4044,N_1038,N_37);
and U4045 (N_4045,N_2483,N_1765);
xnor U4046 (N_4046,N_2285,N_2093);
nor U4047 (N_4047,N_829,N_2011);
and U4048 (N_4048,N_1478,N_2083);
or U4049 (N_4049,N_708,N_1233);
nand U4050 (N_4050,N_1164,N_667);
nor U4051 (N_4051,N_2352,N_1798);
and U4052 (N_4052,N_1254,N_390);
and U4053 (N_4053,N_1683,N_715);
nor U4054 (N_4054,N_2396,N_42);
nand U4055 (N_4055,N_1240,N_215);
and U4056 (N_4056,N_1055,N_1206);
or U4057 (N_4057,N_1755,N_414);
xor U4058 (N_4058,N_1353,N_722);
xnor U4059 (N_4059,N_2446,N_1737);
nand U4060 (N_4060,N_809,N_1742);
or U4061 (N_4061,N_1925,N_65);
and U4062 (N_4062,N_33,N_2234);
or U4063 (N_4063,N_2220,N_443);
or U4064 (N_4064,N_1881,N_1289);
nand U4065 (N_4065,N_2447,N_1205);
or U4066 (N_4066,N_2054,N_123);
or U4067 (N_4067,N_1133,N_2143);
and U4068 (N_4068,N_501,N_1853);
and U4069 (N_4069,N_1689,N_666);
nor U4070 (N_4070,N_1963,N_2483);
and U4071 (N_4071,N_1787,N_1632);
and U4072 (N_4072,N_2419,N_597);
nand U4073 (N_4073,N_490,N_8);
nand U4074 (N_4074,N_787,N_1985);
and U4075 (N_4075,N_919,N_2140);
and U4076 (N_4076,N_1607,N_813);
nand U4077 (N_4077,N_1439,N_2018);
or U4078 (N_4078,N_26,N_2470);
nand U4079 (N_4079,N_835,N_1836);
nor U4080 (N_4080,N_1368,N_1214);
nor U4081 (N_4081,N_267,N_509);
xor U4082 (N_4082,N_56,N_251);
nand U4083 (N_4083,N_1062,N_2326);
nand U4084 (N_4084,N_63,N_1887);
or U4085 (N_4085,N_1046,N_1295);
nor U4086 (N_4086,N_1285,N_1198);
nand U4087 (N_4087,N_2280,N_742);
or U4088 (N_4088,N_1707,N_582);
nand U4089 (N_4089,N_1555,N_2497);
and U4090 (N_4090,N_2080,N_1692);
and U4091 (N_4091,N_442,N_424);
and U4092 (N_4092,N_1390,N_1686);
nand U4093 (N_4093,N_2012,N_2079);
nand U4094 (N_4094,N_1383,N_370);
or U4095 (N_4095,N_526,N_1171);
and U4096 (N_4096,N_2184,N_2400);
nor U4097 (N_4097,N_912,N_1754);
and U4098 (N_4098,N_2376,N_2042);
nor U4099 (N_4099,N_884,N_95);
xor U4100 (N_4100,N_531,N_329);
and U4101 (N_4101,N_2449,N_1404);
or U4102 (N_4102,N_1027,N_670);
or U4103 (N_4103,N_1452,N_66);
xnor U4104 (N_4104,N_553,N_1434);
and U4105 (N_4105,N_1860,N_481);
or U4106 (N_4106,N_2166,N_1144);
nand U4107 (N_4107,N_46,N_1495);
nor U4108 (N_4108,N_606,N_1825);
or U4109 (N_4109,N_1821,N_2114);
and U4110 (N_4110,N_253,N_1303);
nand U4111 (N_4111,N_1026,N_305);
and U4112 (N_4112,N_1667,N_718);
and U4113 (N_4113,N_1399,N_94);
nand U4114 (N_4114,N_1265,N_655);
nand U4115 (N_4115,N_1669,N_1749);
and U4116 (N_4116,N_2409,N_73);
nor U4117 (N_4117,N_94,N_963);
nand U4118 (N_4118,N_2202,N_1455);
nand U4119 (N_4119,N_1950,N_1033);
nand U4120 (N_4120,N_2283,N_1737);
or U4121 (N_4121,N_1546,N_30);
or U4122 (N_4122,N_1746,N_2312);
and U4123 (N_4123,N_1782,N_426);
nor U4124 (N_4124,N_1526,N_1053);
nor U4125 (N_4125,N_776,N_2194);
xnor U4126 (N_4126,N_705,N_1270);
or U4127 (N_4127,N_875,N_82);
and U4128 (N_4128,N_1761,N_1493);
nand U4129 (N_4129,N_929,N_262);
and U4130 (N_4130,N_2434,N_56);
nand U4131 (N_4131,N_1918,N_1123);
nor U4132 (N_4132,N_156,N_1025);
and U4133 (N_4133,N_1817,N_1314);
xor U4134 (N_4134,N_2270,N_1868);
xor U4135 (N_4135,N_275,N_2203);
xor U4136 (N_4136,N_496,N_787);
xor U4137 (N_4137,N_153,N_701);
nand U4138 (N_4138,N_187,N_1987);
or U4139 (N_4139,N_2328,N_1527);
nor U4140 (N_4140,N_214,N_229);
nor U4141 (N_4141,N_109,N_2126);
or U4142 (N_4142,N_2044,N_152);
nor U4143 (N_4143,N_578,N_656);
nand U4144 (N_4144,N_927,N_978);
nor U4145 (N_4145,N_12,N_41);
nand U4146 (N_4146,N_806,N_1117);
and U4147 (N_4147,N_2124,N_1112);
nand U4148 (N_4148,N_1716,N_1290);
or U4149 (N_4149,N_422,N_24);
and U4150 (N_4150,N_1708,N_1288);
xnor U4151 (N_4151,N_860,N_1419);
nand U4152 (N_4152,N_142,N_137);
and U4153 (N_4153,N_1797,N_1700);
nand U4154 (N_4154,N_1138,N_1654);
or U4155 (N_4155,N_207,N_1850);
nand U4156 (N_4156,N_1338,N_1381);
nand U4157 (N_4157,N_7,N_152);
or U4158 (N_4158,N_737,N_2236);
and U4159 (N_4159,N_987,N_1792);
xor U4160 (N_4160,N_1709,N_1998);
or U4161 (N_4161,N_830,N_1213);
nand U4162 (N_4162,N_2206,N_776);
nor U4163 (N_4163,N_1777,N_1415);
nand U4164 (N_4164,N_815,N_1903);
and U4165 (N_4165,N_480,N_2030);
and U4166 (N_4166,N_42,N_2060);
or U4167 (N_4167,N_826,N_2120);
and U4168 (N_4168,N_924,N_2173);
nand U4169 (N_4169,N_729,N_59);
nand U4170 (N_4170,N_1422,N_1785);
or U4171 (N_4171,N_2395,N_161);
nor U4172 (N_4172,N_874,N_1952);
nor U4173 (N_4173,N_2240,N_2403);
or U4174 (N_4174,N_889,N_2344);
xnor U4175 (N_4175,N_1929,N_312);
or U4176 (N_4176,N_356,N_2237);
and U4177 (N_4177,N_2408,N_704);
or U4178 (N_4178,N_2471,N_1620);
xnor U4179 (N_4179,N_1667,N_2039);
or U4180 (N_4180,N_2186,N_2459);
or U4181 (N_4181,N_1160,N_578);
nand U4182 (N_4182,N_1832,N_2372);
and U4183 (N_4183,N_2117,N_1909);
nand U4184 (N_4184,N_1912,N_101);
or U4185 (N_4185,N_1990,N_1412);
nand U4186 (N_4186,N_2205,N_717);
nand U4187 (N_4187,N_844,N_271);
and U4188 (N_4188,N_546,N_351);
nand U4189 (N_4189,N_2071,N_262);
and U4190 (N_4190,N_1951,N_725);
or U4191 (N_4191,N_144,N_2379);
nor U4192 (N_4192,N_751,N_1039);
and U4193 (N_4193,N_1224,N_527);
and U4194 (N_4194,N_395,N_834);
xnor U4195 (N_4195,N_1986,N_2438);
and U4196 (N_4196,N_257,N_219);
nand U4197 (N_4197,N_712,N_166);
or U4198 (N_4198,N_1941,N_1349);
or U4199 (N_4199,N_882,N_2416);
nor U4200 (N_4200,N_1587,N_1678);
xnor U4201 (N_4201,N_2392,N_2407);
nand U4202 (N_4202,N_78,N_1048);
or U4203 (N_4203,N_628,N_145);
nand U4204 (N_4204,N_790,N_595);
or U4205 (N_4205,N_360,N_1666);
or U4206 (N_4206,N_2268,N_2129);
and U4207 (N_4207,N_866,N_2358);
nor U4208 (N_4208,N_2200,N_7);
nand U4209 (N_4209,N_823,N_2294);
and U4210 (N_4210,N_982,N_642);
and U4211 (N_4211,N_932,N_1895);
nor U4212 (N_4212,N_2183,N_1385);
nor U4213 (N_4213,N_1418,N_1459);
nor U4214 (N_4214,N_2132,N_587);
xor U4215 (N_4215,N_170,N_262);
and U4216 (N_4216,N_538,N_445);
nand U4217 (N_4217,N_2307,N_1579);
or U4218 (N_4218,N_1677,N_1569);
nor U4219 (N_4219,N_2483,N_105);
nor U4220 (N_4220,N_1450,N_2367);
nor U4221 (N_4221,N_911,N_1868);
and U4222 (N_4222,N_1463,N_807);
nor U4223 (N_4223,N_393,N_2255);
or U4224 (N_4224,N_1120,N_768);
nor U4225 (N_4225,N_644,N_345);
and U4226 (N_4226,N_1640,N_2426);
xor U4227 (N_4227,N_1180,N_1210);
nand U4228 (N_4228,N_1783,N_2043);
and U4229 (N_4229,N_887,N_2338);
xnor U4230 (N_4230,N_1822,N_1018);
nand U4231 (N_4231,N_1604,N_2122);
nand U4232 (N_4232,N_1102,N_2454);
nor U4233 (N_4233,N_1278,N_848);
nor U4234 (N_4234,N_700,N_25);
and U4235 (N_4235,N_1426,N_757);
or U4236 (N_4236,N_852,N_487);
nand U4237 (N_4237,N_2391,N_680);
nor U4238 (N_4238,N_1796,N_354);
and U4239 (N_4239,N_359,N_1217);
nor U4240 (N_4240,N_2111,N_1427);
and U4241 (N_4241,N_1158,N_1235);
or U4242 (N_4242,N_1595,N_2331);
and U4243 (N_4243,N_2122,N_1751);
or U4244 (N_4244,N_905,N_1521);
nand U4245 (N_4245,N_184,N_288);
or U4246 (N_4246,N_996,N_2428);
nand U4247 (N_4247,N_2140,N_405);
and U4248 (N_4248,N_1331,N_1040);
and U4249 (N_4249,N_2365,N_974);
nor U4250 (N_4250,N_1642,N_1748);
or U4251 (N_4251,N_1078,N_802);
nand U4252 (N_4252,N_1735,N_1719);
and U4253 (N_4253,N_1869,N_2156);
or U4254 (N_4254,N_51,N_924);
nor U4255 (N_4255,N_911,N_628);
nand U4256 (N_4256,N_1704,N_221);
or U4257 (N_4257,N_1079,N_1977);
and U4258 (N_4258,N_695,N_291);
nand U4259 (N_4259,N_1156,N_1243);
or U4260 (N_4260,N_157,N_1000);
and U4261 (N_4261,N_90,N_2057);
nand U4262 (N_4262,N_789,N_967);
nand U4263 (N_4263,N_276,N_2450);
nor U4264 (N_4264,N_1749,N_1614);
nor U4265 (N_4265,N_2395,N_2281);
nor U4266 (N_4266,N_346,N_1903);
nand U4267 (N_4267,N_2304,N_1847);
nand U4268 (N_4268,N_219,N_1206);
and U4269 (N_4269,N_112,N_651);
nor U4270 (N_4270,N_2103,N_1523);
or U4271 (N_4271,N_364,N_880);
and U4272 (N_4272,N_683,N_1327);
and U4273 (N_4273,N_461,N_1078);
or U4274 (N_4274,N_232,N_329);
nand U4275 (N_4275,N_1085,N_2455);
nand U4276 (N_4276,N_1916,N_379);
and U4277 (N_4277,N_1666,N_801);
or U4278 (N_4278,N_577,N_2374);
nand U4279 (N_4279,N_937,N_899);
or U4280 (N_4280,N_1116,N_1740);
nor U4281 (N_4281,N_1253,N_223);
nand U4282 (N_4282,N_728,N_1586);
and U4283 (N_4283,N_2342,N_1273);
xnor U4284 (N_4284,N_2308,N_1025);
or U4285 (N_4285,N_1185,N_2060);
or U4286 (N_4286,N_204,N_174);
xnor U4287 (N_4287,N_1088,N_1422);
nor U4288 (N_4288,N_750,N_2227);
xor U4289 (N_4289,N_1261,N_967);
nor U4290 (N_4290,N_1214,N_228);
nand U4291 (N_4291,N_251,N_2271);
nand U4292 (N_4292,N_2242,N_2055);
xnor U4293 (N_4293,N_2190,N_1580);
nor U4294 (N_4294,N_576,N_2274);
or U4295 (N_4295,N_537,N_1251);
or U4296 (N_4296,N_1700,N_2203);
or U4297 (N_4297,N_1190,N_2473);
nor U4298 (N_4298,N_2403,N_1959);
nor U4299 (N_4299,N_2162,N_2212);
nor U4300 (N_4300,N_347,N_27);
nor U4301 (N_4301,N_392,N_1348);
nor U4302 (N_4302,N_1529,N_2128);
or U4303 (N_4303,N_2493,N_1440);
nor U4304 (N_4304,N_17,N_2042);
nor U4305 (N_4305,N_2269,N_251);
nand U4306 (N_4306,N_1354,N_279);
or U4307 (N_4307,N_1547,N_431);
nor U4308 (N_4308,N_1807,N_1794);
and U4309 (N_4309,N_1287,N_1462);
xor U4310 (N_4310,N_318,N_814);
or U4311 (N_4311,N_1971,N_2202);
xnor U4312 (N_4312,N_726,N_1825);
or U4313 (N_4313,N_786,N_876);
nor U4314 (N_4314,N_1434,N_556);
nand U4315 (N_4315,N_1899,N_115);
nand U4316 (N_4316,N_1632,N_248);
and U4317 (N_4317,N_1633,N_2065);
and U4318 (N_4318,N_2206,N_712);
xor U4319 (N_4319,N_2056,N_668);
nand U4320 (N_4320,N_1625,N_13);
nor U4321 (N_4321,N_2356,N_1831);
nor U4322 (N_4322,N_2062,N_1349);
and U4323 (N_4323,N_1958,N_1714);
or U4324 (N_4324,N_1172,N_1923);
and U4325 (N_4325,N_1864,N_1890);
or U4326 (N_4326,N_1,N_569);
or U4327 (N_4327,N_2316,N_1685);
or U4328 (N_4328,N_681,N_1532);
or U4329 (N_4329,N_279,N_1733);
nor U4330 (N_4330,N_1735,N_2418);
and U4331 (N_4331,N_45,N_1537);
or U4332 (N_4332,N_92,N_968);
nor U4333 (N_4333,N_665,N_687);
or U4334 (N_4334,N_206,N_1459);
and U4335 (N_4335,N_15,N_50);
nand U4336 (N_4336,N_1178,N_510);
and U4337 (N_4337,N_761,N_1300);
or U4338 (N_4338,N_535,N_631);
and U4339 (N_4339,N_279,N_1737);
and U4340 (N_4340,N_1565,N_76);
nand U4341 (N_4341,N_646,N_2316);
xor U4342 (N_4342,N_1994,N_1778);
nor U4343 (N_4343,N_1758,N_2477);
and U4344 (N_4344,N_2378,N_1667);
xnor U4345 (N_4345,N_2107,N_318);
xnor U4346 (N_4346,N_1132,N_451);
nor U4347 (N_4347,N_7,N_1488);
xnor U4348 (N_4348,N_2207,N_1801);
and U4349 (N_4349,N_745,N_1683);
and U4350 (N_4350,N_1052,N_2125);
and U4351 (N_4351,N_1697,N_1904);
or U4352 (N_4352,N_1190,N_322);
or U4353 (N_4353,N_720,N_1022);
nor U4354 (N_4354,N_1022,N_946);
nor U4355 (N_4355,N_2125,N_2379);
nand U4356 (N_4356,N_666,N_1700);
nor U4357 (N_4357,N_347,N_190);
nor U4358 (N_4358,N_732,N_1802);
nand U4359 (N_4359,N_1531,N_491);
nand U4360 (N_4360,N_656,N_394);
nor U4361 (N_4361,N_1611,N_409);
nor U4362 (N_4362,N_866,N_452);
nand U4363 (N_4363,N_2208,N_1767);
and U4364 (N_4364,N_1496,N_685);
xor U4365 (N_4365,N_241,N_1298);
nor U4366 (N_4366,N_618,N_1868);
and U4367 (N_4367,N_1809,N_1549);
nor U4368 (N_4368,N_2065,N_416);
nor U4369 (N_4369,N_1490,N_665);
nor U4370 (N_4370,N_1434,N_79);
nor U4371 (N_4371,N_2236,N_610);
nand U4372 (N_4372,N_2361,N_1766);
and U4373 (N_4373,N_2466,N_1159);
nand U4374 (N_4374,N_2130,N_1174);
or U4375 (N_4375,N_2353,N_1324);
and U4376 (N_4376,N_757,N_1554);
or U4377 (N_4377,N_1647,N_1969);
and U4378 (N_4378,N_577,N_1900);
nor U4379 (N_4379,N_1828,N_1077);
xnor U4380 (N_4380,N_952,N_592);
or U4381 (N_4381,N_712,N_2132);
nand U4382 (N_4382,N_122,N_139);
or U4383 (N_4383,N_1717,N_2138);
nor U4384 (N_4384,N_2133,N_1807);
xnor U4385 (N_4385,N_2315,N_2438);
and U4386 (N_4386,N_771,N_306);
nor U4387 (N_4387,N_1169,N_9);
xnor U4388 (N_4388,N_1040,N_1265);
xnor U4389 (N_4389,N_1224,N_2093);
or U4390 (N_4390,N_88,N_972);
nor U4391 (N_4391,N_1504,N_20);
or U4392 (N_4392,N_1675,N_565);
or U4393 (N_4393,N_1402,N_1244);
xor U4394 (N_4394,N_2029,N_1293);
nand U4395 (N_4395,N_747,N_1670);
nand U4396 (N_4396,N_852,N_1198);
nand U4397 (N_4397,N_2135,N_1243);
nand U4398 (N_4398,N_437,N_2168);
or U4399 (N_4399,N_773,N_2229);
or U4400 (N_4400,N_818,N_1441);
nor U4401 (N_4401,N_2168,N_2391);
xnor U4402 (N_4402,N_1931,N_1922);
and U4403 (N_4403,N_1028,N_1927);
nand U4404 (N_4404,N_1824,N_1782);
or U4405 (N_4405,N_1567,N_1328);
or U4406 (N_4406,N_168,N_1892);
and U4407 (N_4407,N_992,N_682);
or U4408 (N_4408,N_2378,N_1839);
and U4409 (N_4409,N_168,N_1152);
and U4410 (N_4410,N_971,N_1319);
nor U4411 (N_4411,N_1795,N_2319);
nand U4412 (N_4412,N_1115,N_4);
nor U4413 (N_4413,N_617,N_460);
xor U4414 (N_4414,N_1216,N_691);
or U4415 (N_4415,N_1919,N_2285);
nand U4416 (N_4416,N_314,N_1388);
nand U4417 (N_4417,N_1873,N_2422);
or U4418 (N_4418,N_532,N_838);
nor U4419 (N_4419,N_41,N_695);
or U4420 (N_4420,N_1196,N_1920);
and U4421 (N_4421,N_721,N_1277);
nor U4422 (N_4422,N_1268,N_1513);
and U4423 (N_4423,N_1657,N_898);
xor U4424 (N_4424,N_960,N_578);
nand U4425 (N_4425,N_2159,N_1692);
or U4426 (N_4426,N_164,N_91);
nor U4427 (N_4427,N_1669,N_1885);
or U4428 (N_4428,N_1163,N_1331);
or U4429 (N_4429,N_44,N_1698);
or U4430 (N_4430,N_1126,N_2307);
or U4431 (N_4431,N_2304,N_1336);
nand U4432 (N_4432,N_16,N_713);
or U4433 (N_4433,N_1451,N_21);
or U4434 (N_4434,N_50,N_47);
nand U4435 (N_4435,N_584,N_723);
nor U4436 (N_4436,N_153,N_2435);
nor U4437 (N_4437,N_1235,N_2002);
and U4438 (N_4438,N_712,N_2295);
nand U4439 (N_4439,N_1145,N_2178);
nor U4440 (N_4440,N_1865,N_776);
nor U4441 (N_4441,N_2429,N_2187);
or U4442 (N_4442,N_1834,N_1978);
nor U4443 (N_4443,N_1061,N_1030);
or U4444 (N_4444,N_1363,N_518);
nor U4445 (N_4445,N_1673,N_1097);
nand U4446 (N_4446,N_540,N_1659);
nor U4447 (N_4447,N_897,N_2068);
nor U4448 (N_4448,N_578,N_500);
xor U4449 (N_4449,N_2344,N_608);
nor U4450 (N_4450,N_2399,N_1207);
and U4451 (N_4451,N_1077,N_710);
nand U4452 (N_4452,N_1625,N_11);
nor U4453 (N_4453,N_1641,N_1044);
nand U4454 (N_4454,N_2011,N_572);
nand U4455 (N_4455,N_927,N_855);
or U4456 (N_4456,N_2406,N_1970);
nand U4457 (N_4457,N_446,N_133);
xnor U4458 (N_4458,N_2164,N_1795);
xnor U4459 (N_4459,N_2002,N_1754);
nand U4460 (N_4460,N_773,N_578);
nor U4461 (N_4461,N_2321,N_1149);
nor U4462 (N_4462,N_827,N_1983);
nor U4463 (N_4463,N_1602,N_2384);
and U4464 (N_4464,N_1032,N_1365);
nand U4465 (N_4465,N_759,N_728);
or U4466 (N_4466,N_1017,N_61);
xor U4467 (N_4467,N_1336,N_695);
and U4468 (N_4468,N_635,N_1954);
or U4469 (N_4469,N_533,N_1768);
and U4470 (N_4470,N_1437,N_47);
or U4471 (N_4471,N_129,N_894);
or U4472 (N_4472,N_538,N_48);
nor U4473 (N_4473,N_517,N_958);
nand U4474 (N_4474,N_683,N_1562);
or U4475 (N_4475,N_524,N_1230);
xnor U4476 (N_4476,N_1928,N_1185);
nor U4477 (N_4477,N_2475,N_274);
nand U4478 (N_4478,N_568,N_1074);
nor U4479 (N_4479,N_570,N_953);
nand U4480 (N_4480,N_1553,N_994);
or U4481 (N_4481,N_263,N_224);
and U4482 (N_4482,N_1867,N_42);
nand U4483 (N_4483,N_2111,N_1982);
nor U4484 (N_4484,N_2329,N_738);
xor U4485 (N_4485,N_120,N_2064);
nand U4486 (N_4486,N_1460,N_1957);
nand U4487 (N_4487,N_1810,N_2480);
nor U4488 (N_4488,N_678,N_1298);
xor U4489 (N_4489,N_2198,N_1969);
or U4490 (N_4490,N_2013,N_1464);
nand U4491 (N_4491,N_2251,N_46);
and U4492 (N_4492,N_1027,N_1594);
nor U4493 (N_4493,N_52,N_600);
and U4494 (N_4494,N_1229,N_598);
or U4495 (N_4495,N_1696,N_835);
or U4496 (N_4496,N_766,N_1098);
or U4497 (N_4497,N_2127,N_2366);
nor U4498 (N_4498,N_348,N_2163);
or U4499 (N_4499,N_342,N_378);
nor U4500 (N_4500,N_685,N_1915);
and U4501 (N_4501,N_1971,N_1917);
and U4502 (N_4502,N_1980,N_555);
nand U4503 (N_4503,N_1645,N_1018);
nor U4504 (N_4504,N_363,N_2111);
or U4505 (N_4505,N_610,N_1926);
xnor U4506 (N_4506,N_375,N_2479);
nand U4507 (N_4507,N_261,N_326);
nand U4508 (N_4508,N_1555,N_410);
xor U4509 (N_4509,N_611,N_2278);
nor U4510 (N_4510,N_2441,N_2154);
or U4511 (N_4511,N_152,N_1553);
and U4512 (N_4512,N_241,N_938);
or U4513 (N_4513,N_2028,N_686);
xnor U4514 (N_4514,N_1104,N_867);
or U4515 (N_4515,N_2006,N_1082);
nor U4516 (N_4516,N_1274,N_632);
nand U4517 (N_4517,N_1913,N_1168);
or U4518 (N_4518,N_2231,N_1633);
xor U4519 (N_4519,N_2054,N_1615);
or U4520 (N_4520,N_2477,N_2411);
and U4521 (N_4521,N_2371,N_1373);
nor U4522 (N_4522,N_1496,N_240);
nand U4523 (N_4523,N_507,N_1150);
nand U4524 (N_4524,N_41,N_588);
nand U4525 (N_4525,N_1621,N_2140);
xnor U4526 (N_4526,N_562,N_2434);
xor U4527 (N_4527,N_650,N_527);
and U4528 (N_4528,N_78,N_1729);
nor U4529 (N_4529,N_432,N_2450);
and U4530 (N_4530,N_1000,N_2163);
or U4531 (N_4531,N_1956,N_1832);
xor U4532 (N_4532,N_235,N_714);
nor U4533 (N_4533,N_2190,N_1881);
nand U4534 (N_4534,N_1970,N_2358);
or U4535 (N_4535,N_1320,N_2229);
nor U4536 (N_4536,N_813,N_1446);
or U4537 (N_4537,N_984,N_279);
xnor U4538 (N_4538,N_1570,N_1909);
and U4539 (N_4539,N_989,N_1100);
or U4540 (N_4540,N_1282,N_746);
nor U4541 (N_4541,N_128,N_2028);
and U4542 (N_4542,N_885,N_2154);
nand U4543 (N_4543,N_1570,N_1695);
nor U4544 (N_4544,N_699,N_2075);
and U4545 (N_4545,N_561,N_1092);
and U4546 (N_4546,N_552,N_2410);
xor U4547 (N_4547,N_723,N_406);
or U4548 (N_4548,N_1826,N_614);
and U4549 (N_4549,N_324,N_2176);
and U4550 (N_4550,N_1891,N_1821);
xor U4551 (N_4551,N_452,N_965);
xnor U4552 (N_4552,N_2428,N_9);
and U4553 (N_4553,N_2351,N_1587);
nor U4554 (N_4554,N_625,N_1030);
and U4555 (N_4555,N_1650,N_141);
and U4556 (N_4556,N_1487,N_434);
or U4557 (N_4557,N_1402,N_1735);
nand U4558 (N_4558,N_1190,N_1881);
nor U4559 (N_4559,N_1776,N_1408);
nand U4560 (N_4560,N_2362,N_875);
nor U4561 (N_4561,N_2086,N_761);
nand U4562 (N_4562,N_1621,N_2451);
xor U4563 (N_4563,N_2337,N_1334);
nand U4564 (N_4564,N_904,N_690);
nor U4565 (N_4565,N_1334,N_486);
or U4566 (N_4566,N_2214,N_2454);
nand U4567 (N_4567,N_1599,N_1905);
and U4568 (N_4568,N_2246,N_1280);
or U4569 (N_4569,N_273,N_1510);
or U4570 (N_4570,N_157,N_1451);
or U4571 (N_4571,N_2147,N_171);
nor U4572 (N_4572,N_1565,N_1012);
and U4573 (N_4573,N_1654,N_79);
or U4574 (N_4574,N_1046,N_178);
nor U4575 (N_4575,N_2312,N_184);
or U4576 (N_4576,N_398,N_1129);
nor U4577 (N_4577,N_1753,N_2244);
nor U4578 (N_4578,N_1124,N_831);
and U4579 (N_4579,N_610,N_1104);
nor U4580 (N_4580,N_1646,N_2411);
or U4581 (N_4581,N_957,N_164);
nor U4582 (N_4582,N_404,N_1294);
or U4583 (N_4583,N_1576,N_1626);
nor U4584 (N_4584,N_219,N_1894);
and U4585 (N_4585,N_51,N_1454);
nand U4586 (N_4586,N_397,N_429);
or U4587 (N_4587,N_249,N_1331);
xnor U4588 (N_4588,N_1207,N_360);
nand U4589 (N_4589,N_1127,N_2403);
and U4590 (N_4590,N_2154,N_120);
or U4591 (N_4591,N_311,N_1872);
nor U4592 (N_4592,N_215,N_999);
nor U4593 (N_4593,N_1640,N_1361);
or U4594 (N_4594,N_1308,N_1439);
nand U4595 (N_4595,N_634,N_1283);
or U4596 (N_4596,N_546,N_130);
and U4597 (N_4597,N_2163,N_2063);
and U4598 (N_4598,N_1350,N_288);
nor U4599 (N_4599,N_1978,N_1832);
nor U4600 (N_4600,N_1022,N_376);
and U4601 (N_4601,N_2459,N_331);
or U4602 (N_4602,N_726,N_1272);
and U4603 (N_4603,N_2037,N_2430);
or U4604 (N_4604,N_1505,N_1073);
xor U4605 (N_4605,N_1438,N_1160);
nor U4606 (N_4606,N_1978,N_879);
nand U4607 (N_4607,N_1949,N_1476);
nand U4608 (N_4608,N_524,N_259);
and U4609 (N_4609,N_1394,N_1929);
nand U4610 (N_4610,N_1144,N_2176);
or U4611 (N_4611,N_1149,N_1345);
and U4612 (N_4612,N_1854,N_2218);
nand U4613 (N_4613,N_848,N_1243);
nand U4614 (N_4614,N_124,N_2024);
nor U4615 (N_4615,N_2241,N_1168);
nor U4616 (N_4616,N_1677,N_176);
and U4617 (N_4617,N_1392,N_1201);
and U4618 (N_4618,N_1067,N_569);
nor U4619 (N_4619,N_1906,N_500);
nor U4620 (N_4620,N_1468,N_711);
nand U4621 (N_4621,N_1211,N_326);
and U4622 (N_4622,N_811,N_1790);
nor U4623 (N_4623,N_246,N_23);
xor U4624 (N_4624,N_1511,N_1553);
nor U4625 (N_4625,N_1916,N_2131);
and U4626 (N_4626,N_2161,N_375);
nor U4627 (N_4627,N_1452,N_2003);
and U4628 (N_4628,N_743,N_2228);
or U4629 (N_4629,N_1745,N_2149);
xor U4630 (N_4630,N_867,N_169);
nor U4631 (N_4631,N_1345,N_1955);
xor U4632 (N_4632,N_2469,N_2398);
xor U4633 (N_4633,N_175,N_638);
or U4634 (N_4634,N_781,N_794);
nand U4635 (N_4635,N_834,N_1598);
nand U4636 (N_4636,N_754,N_1272);
or U4637 (N_4637,N_2290,N_1628);
nand U4638 (N_4638,N_592,N_1581);
nand U4639 (N_4639,N_792,N_916);
nor U4640 (N_4640,N_1074,N_1124);
nand U4641 (N_4641,N_68,N_838);
or U4642 (N_4642,N_279,N_2033);
nand U4643 (N_4643,N_443,N_2224);
or U4644 (N_4644,N_1850,N_1908);
nand U4645 (N_4645,N_677,N_1062);
nand U4646 (N_4646,N_780,N_1828);
or U4647 (N_4647,N_1631,N_1311);
or U4648 (N_4648,N_2082,N_464);
nor U4649 (N_4649,N_710,N_364);
nand U4650 (N_4650,N_1842,N_177);
nand U4651 (N_4651,N_1933,N_2117);
xnor U4652 (N_4652,N_2470,N_1797);
nand U4653 (N_4653,N_615,N_138);
xor U4654 (N_4654,N_2209,N_162);
nor U4655 (N_4655,N_796,N_1491);
and U4656 (N_4656,N_854,N_1148);
and U4657 (N_4657,N_2342,N_1456);
nor U4658 (N_4658,N_806,N_264);
nand U4659 (N_4659,N_809,N_1458);
nand U4660 (N_4660,N_1337,N_2258);
nor U4661 (N_4661,N_678,N_570);
nor U4662 (N_4662,N_657,N_12);
and U4663 (N_4663,N_243,N_1681);
and U4664 (N_4664,N_1952,N_2288);
nand U4665 (N_4665,N_2130,N_574);
or U4666 (N_4666,N_322,N_1850);
or U4667 (N_4667,N_640,N_473);
nand U4668 (N_4668,N_1446,N_1886);
or U4669 (N_4669,N_1153,N_2053);
nand U4670 (N_4670,N_1550,N_2447);
or U4671 (N_4671,N_2352,N_241);
xnor U4672 (N_4672,N_2298,N_962);
and U4673 (N_4673,N_992,N_1410);
and U4674 (N_4674,N_1859,N_737);
nor U4675 (N_4675,N_727,N_1468);
nand U4676 (N_4676,N_189,N_1535);
xnor U4677 (N_4677,N_906,N_619);
xnor U4678 (N_4678,N_94,N_2304);
nand U4679 (N_4679,N_192,N_273);
xor U4680 (N_4680,N_586,N_1441);
or U4681 (N_4681,N_534,N_1360);
and U4682 (N_4682,N_1314,N_310);
and U4683 (N_4683,N_2213,N_195);
xnor U4684 (N_4684,N_1172,N_1497);
nor U4685 (N_4685,N_2438,N_987);
and U4686 (N_4686,N_2243,N_35);
nand U4687 (N_4687,N_1227,N_860);
nand U4688 (N_4688,N_2456,N_706);
nor U4689 (N_4689,N_2038,N_2276);
or U4690 (N_4690,N_1363,N_2213);
nor U4691 (N_4691,N_1003,N_671);
and U4692 (N_4692,N_353,N_740);
xnor U4693 (N_4693,N_1678,N_912);
nor U4694 (N_4694,N_1138,N_675);
nand U4695 (N_4695,N_1559,N_2295);
nand U4696 (N_4696,N_789,N_1841);
and U4697 (N_4697,N_1025,N_225);
and U4698 (N_4698,N_1411,N_1736);
nor U4699 (N_4699,N_2365,N_1152);
nand U4700 (N_4700,N_119,N_927);
nor U4701 (N_4701,N_1451,N_278);
or U4702 (N_4702,N_753,N_2404);
xor U4703 (N_4703,N_774,N_1208);
nor U4704 (N_4704,N_2190,N_583);
or U4705 (N_4705,N_2493,N_338);
nand U4706 (N_4706,N_832,N_2165);
or U4707 (N_4707,N_2300,N_2039);
nor U4708 (N_4708,N_912,N_1077);
nor U4709 (N_4709,N_2325,N_2209);
or U4710 (N_4710,N_1051,N_1321);
nor U4711 (N_4711,N_1694,N_2491);
or U4712 (N_4712,N_413,N_1988);
xnor U4713 (N_4713,N_1616,N_2215);
or U4714 (N_4714,N_692,N_2451);
nand U4715 (N_4715,N_1092,N_2201);
or U4716 (N_4716,N_1270,N_873);
and U4717 (N_4717,N_1558,N_669);
and U4718 (N_4718,N_962,N_484);
or U4719 (N_4719,N_2127,N_2344);
nor U4720 (N_4720,N_2183,N_1951);
or U4721 (N_4721,N_926,N_379);
or U4722 (N_4722,N_2168,N_273);
nand U4723 (N_4723,N_1409,N_1665);
nor U4724 (N_4724,N_1261,N_628);
nor U4725 (N_4725,N_1055,N_732);
nand U4726 (N_4726,N_1807,N_90);
or U4727 (N_4727,N_946,N_2201);
or U4728 (N_4728,N_1037,N_1867);
nand U4729 (N_4729,N_2404,N_1541);
and U4730 (N_4730,N_992,N_489);
nand U4731 (N_4731,N_563,N_240);
or U4732 (N_4732,N_701,N_60);
or U4733 (N_4733,N_1696,N_1481);
or U4734 (N_4734,N_542,N_869);
and U4735 (N_4735,N_2290,N_1825);
or U4736 (N_4736,N_135,N_2181);
nor U4737 (N_4737,N_1282,N_597);
nor U4738 (N_4738,N_1773,N_1426);
and U4739 (N_4739,N_2192,N_1947);
or U4740 (N_4740,N_2187,N_1030);
nor U4741 (N_4741,N_1696,N_2397);
or U4742 (N_4742,N_579,N_1682);
and U4743 (N_4743,N_1079,N_1537);
or U4744 (N_4744,N_1436,N_1131);
xnor U4745 (N_4745,N_2159,N_1892);
or U4746 (N_4746,N_1709,N_872);
or U4747 (N_4747,N_1994,N_447);
nor U4748 (N_4748,N_1971,N_1265);
nor U4749 (N_4749,N_820,N_1129);
nor U4750 (N_4750,N_2305,N_1297);
nand U4751 (N_4751,N_672,N_1684);
and U4752 (N_4752,N_1162,N_1203);
and U4753 (N_4753,N_709,N_1567);
nor U4754 (N_4754,N_1286,N_939);
nand U4755 (N_4755,N_745,N_481);
nor U4756 (N_4756,N_54,N_319);
xor U4757 (N_4757,N_243,N_782);
xnor U4758 (N_4758,N_1166,N_1134);
and U4759 (N_4759,N_2375,N_1161);
and U4760 (N_4760,N_2161,N_70);
or U4761 (N_4761,N_182,N_1662);
and U4762 (N_4762,N_908,N_1467);
nand U4763 (N_4763,N_1539,N_614);
nand U4764 (N_4764,N_356,N_163);
nor U4765 (N_4765,N_430,N_1874);
and U4766 (N_4766,N_563,N_1937);
and U4767 (N_4767,N_2204,N_937);
nor U4768 (N_4768,N_2338,N_1506);
nor U4769 (N_4769,N_1723,N_1788);
nand U4770 (N_4770,N_691,N_887);
nand U4771 (N_4771,N_1827,N_669);
and U4772 (N_4772,N_725,N_1893);
nor U4773 (N_4773,N_994,N_858);
nor U4774 (N_4774,N_1735,N_142);
nor U4775 (N_4775,N_1380,N_23);
nor U4776 (N_4776,N_1869,N_1127);
nor U4777 (N_4777,N_2266,N_1377);
nor U4778 (N_4778,N_1017,N_2484);
nand U4779 (N_4779,N_1316,N_1903);
or U4780 (N_4780,N_1602,N_1822);
nor U4781 (N_4781,N_849,N_1409);
and U4782 (N_4782,N_504,N_261);
and U4783 (N_4783,N_1973,N_1263);
nand U4784 (N_4784,N_484,N_1605);
and U4785 (N_4785,N_1986,N_82);
and U4786 (N_4786,N_679,N_1552);
xor U4787 (N_4787,N_821,N_2042);
xor U4788 (N_4788,N_1414,N_1571);
and U4789 (N_4789,N_2329,N_308);
and U4790 (N_4790,N_2133,N_2059);
and U4791 (N_4791,N_1574,N_1875);
and U4792 (N_4792,N_391,N_888);
or U4793 (N_4793,N_83,N_2211);
xnor U4794 (N_4794,N_619,N_309);
xnor U4795 (N_4795,N_2395,N_2074);
or U4796 (N_4796,N_2381,N_36);
and U4797 (N_4797,N_1377,N_2112);
and U4798 (N_4798,N_273,N_657);
nor U4799 (N_4799,N_1366,N_1510);
nor U4800 (N_4800,N_9,N_20);
nor U4801 (N_4801,N_1645,N_964);
nand U4802 (N_4802,N_1531,N_2360);
nor U4803 (N_4803,N_1738,N_873);
or U4804 (N_4804,N_315,N_2306);
and U4805 (N_4805,N_698,N_532);
and U4806 (N_4806,N_2377,N_1108);
or U4807 (N_4807,N_1632,N_2265);
and U4808 (N_4808,N_1389,N_1023);
or U4809 (N_4809,N_2174,N_1708);
nor U4810 (N_4810,N_395,N_1829);
and U4811 (N_4811,N_391,N_207);
and U4812 (N_4812,N_433,N_1303);
nor U4813 (N_4813,N_1712,N_1764);
nor U4814 (N_4814,N_2387,N_684);
nand U4815 (N_4815,N_1553,N_2482);
nor U4816 (N_4816,N_379,N_1621);
or U4817 (N_4817,N_2263,N_114);
or U4818 (N_4818,N_299,N_475);
or U4819 (N_4819,N_2105,N_1089);
and U4820 (N_4820,N_451,N_453);
or U4821 (N_4821,N_583,N_1297);
nor U4822 (N_4822,N_302,N_131);
or U4823 (N_4823,N_295,N_2025);
and U4824 (N_4824,N_634,N_993);
nand U4825 (N_4825,N_1032,N_1217);
xnor U4826 (N_4826,N_310,N_264);
nand U4827 (N_4827,N_2472,N_941);
nor U4828 (N_4828,N_426,N_478);
nand U4829 (N_4829,N_2310,N_86);
nand U4830 (N_4830,N_962,N_5);
or U4831 (N_4831,N_1596,N_1653);
nand U4832 (N_4832,N_915,N_2213);
nand U4833 (N_4833,N_2210,N_1689);
nor U4834 (N_4834,N_1426,N_1174);
and U4835 (N_4835,N_1273,N_1477);
or U4836 (N_4836,N_5,N_2219);
or U4837 (N_4837,N_32,N_1165);
nand U4838 (N_4838,N_1263,N_257);
nor U4839 (N_4839,N_128,N_972);
or U4840 (N_4840,N_1981,N_423);
nand U4841 (N_4841,N_2168,N_481);
nand U4842 (N_4842,N_1150,N_2197);
nand U4843 (N_4843,N_1454,N_2280);
xnor U4844 (N_4844,N_1966,N_298);
nand U4845 (N_4845,N_1077,N_428);
and U4846 (N_4846,N_2477,N_953);
or U4847 (N_4847,N_110,N_1442);
or U4848 (N_4848,N_555,N_1851);
nor U4849 (N_4849,N_467,N_893);
or U4850 (N_4850,N_1634,N_2446);
and U4851 (N_4851,N_666,N_1013);
nand U4852 (N_4852,N_1872,N_822);
nand U4853 (N_4853,N_1156,N_404);
or U4854 (N_4854,N_2099,N_89);
or U4855 (N_4855,N_1287,N_483);
or U4856 (N_4856,N_1534,N_60);
and U4857 (N_4857,N_1714,N_2349);
nand U4858 (N_4858,N_1629,N_885);
nand U4859 (N_4859,N_1148,N_2281);
nand U4860 (N_4860,N_1582,N_2350);
or U4861 (N_4861,N_742,N_700);
and U4862 (N_4862,N_2200,N_322);
nor U4863 (N_4863,N_244,N_65);
or U4864 (N_4864,N_1925,N_2181);
or U4865 (N_4865,N_1669,N_445);
nand U4866 (N_4866,N_1306,N_1448);
nand U4867 (N_4867,N_1168,N_899);
or U4868 (N_4868,N_32,N_1404);
or U4869 (N_4869,N_389,N_987);
or U4870 (N_4870,N_2152,N_1704);
nor U4871 (N_4871,N_625,N_2341);
and U4872 (N_4872,N_536,N_1397);
and U4873 (N_4873,N_788,N_475);
xor U4874 (N_4874,N_406,N_2482);
or U4875 (N_4875,N_874,N_2189);
nor U4876 (N_4876,N_1743,N_481);
nand U4877 (N_4877,N_676,N_1802);
or U4878 (N_4878,N_1062,N_1231);
nor U4879 (N_4879,N_2000,N_2324);
nor U4880 (N_4880,N_604,N_1535);
nor U4881 (N_4881,N_510,N_2070);
and U4882 (N_4882,N_9,N_2258);
nor U4883 (N_4883,N_1578,N_2077);
nor U4884 (N_4884,N_412,N_339);
or U4885 (N_4885,N_368,N_1974);
nand U4886 (N_4886,N_1820,N_493);
and U4887 (N_4887,N_2232,N_395);
nand U4888 (N_4888,N_1740,N_1429);
nand U4889 (N_4889,N_1927,N_2307);
nor U4890 (N_4890,N_2252,N_898);
or U4891 (N_4891,N_1900,N_1018);
and U4892 (N_4892,N_406,N_1098);
nand U4893 (N_4893,N_930,N_388);
nand U4894 (N_4894,N_2498,N_1792);
nand U4895 (N_4895,N_2220,N_2138);
or U4896 (N_4896,N_612,N_1883);
and U4897 (N_4897,N_180,N_1219);
nand U4898 (N_4898,N_1563,N_1607);
and U4899 (N_4899,N_1719,N_333);
nand U4900 (N_4900,N_528,N_497);
nand U4901 (N_4901,N_1058,N_974);
and U4902 (N_4902,N_495,N_2384);
nand U4903 (N_4903,N_535,N_1731);
and U4904 (N_4904,N_802,N_1436);
or U4905 (N_4905,N_1554,N_1633);
or U4906 (N_4906,N_1171,N_746);
and U4907 (N_4907,N_267,N_927);
and U4908 (N_4908,N_98,N_1455);
or U4909 (N_4909,N_108,N_1949);
and U4910 (N_4910,N_2078,N_1456);
nor U4911 (N_4911,N_1110,N_953);
xnor U4912 (N_4912,N_683,N_199);
nor U4913 (N_4913,N_4,N_44);
and U4914 (N_4914,N_1843,N_269);
xnor U4915 (N_4915,N_341,N_199);
and U4916 (N_4916,N_1473,N_448);
or U4917 (N_4917,N_1670,N_541);
nor U4918 (N_4918,N_1165,N_1213);
or U4919 (N_4919,N_195,N_1993);
nand U4920 (N_4920,N_2031,N_116);
and U4921 (N_4921,N_2132,N_1842);
or U4922 (N_4922,N_977,N_351);
nand U4923 (N_4923,N_1296,N_1448);
nor U4924 (N_4924,N_591,N_2363);
nor U4925 (N_4925,N_455,N_2434);
and U4926 (N_4926,N_2139,N_197);
and U4927 (N_4927,N_1190,N_1370);
and U4928 (N_4928,N_98,N_1329);
xnor U4929 (N_4929,N_2225,N_1357);
nand U4930 (N_4930,N_1201,N_2388);
or U4931 (N_4931,N_1817,N_989);
or U4932 (N_4932,N_810,N_1969);
nor U4933 (N_4933,N_2152,N_299);
and U4934 (N_4934,N_1646,N_114);
nor U4935 (N_4935,N_217,N_880);
nand U4936 (N_4936,N_203,N_1076);
and U4937 (N_4937,N_1012,N_2063);
nor U4938 (N_4938,N_893,N_1068);
or U4939 (N_4939,N_1240,N_662);
or U4940 (N_4940,N_600,N_1190);
nand U4941 (N_4941,N_813,N_2042);
or U4942 (N_4942,N_1791,N_1235);
nand U4943 (N_4943,N_746,N_2067);
nand U4944 (N_4944,N_1420,N_2002);
nor U4945 (N_4945,N_1100,N_274);
and U4946 (N_4946,N_1929,N_2313);
or U4947 (N_4947,N_2178,N_1892);
nor U4948 (N_4948,N_1308,N_679);
nor U4949 (N_4949,N_802,N_590);
nor U4950 (N_4950,N_2333,N_2476);
nand U4951 (N_4951,N_1641,N_1322);
and U4952 (N_4952,N_1769,N_1358);
and U4953 (N_4953,N_2210,N_1119);
nand U4954 (N_4954,N_659,N_1120);
nand U4955 (N_4955,N_374,N_874);
nand U4956 (N_4956,N_1164,N_806);
and U4957 (N_4957,N_368,N_1316);
nand U4958 (N_4958,N_1718,N_2322);
nor U4959 (N_4959,N_2028,N_934);
or U4960 (N_4960,N_484,N_350);
nand U4961 (N_4961,N_569,N_931);
xor U4962 (N_4962,N_2293,N_322);
and U4963 (N_4963,N_2336,N_155);
and U4964 (N_4964,N_120,N_512);
or U4965 (N_4965,N_86,N_2233);
or U4966 (N_4966,N_2072,N_2461);
or U4967 (N_4967,N_1151,N_323);
or U4968 (N_4968,N_874,N_2393);
nor U4969 (N_4969,N_1216,N_885);
nor U4970 (N_4970,N_2397,N_2145);
or U4971 (N_4971,N_1248,N_2217);
nand U4972 (N_4972,N_649,N_39);
or U4973 (N_4973,N_1723,N_1061);
xnor U4974 (N_4974,N_2168,N_2021);
or U4975 (N_4975,N_1023,N_825);
xnor U4976 (N_4976,N_2203,N_573);
xnor U4977 (N_4977,N_1468,N_1042);
nand U4978 (N_4978,N_587,N_580);
nor U4979 (N_4979,N_503,N_1510);
nor U4980 (N_4980,N_555,N_509);
or U4981 (N_4981,N_2263,N_2064);
and U4982 (N_4982,N_1878,N_1475);
nand U4983 (N_4983,N_1278,N_1688);
nand U4984 (N_4984,N_1074,N_2388);
or U4985 (N_4985,N_2196,N_339);
or U4986 (N_4986,N_89,N_1739);
nor U4987 (N_4987,N_1088,N_201);
and U4988 (N_4988,N_1233,N_693);
or U4989 (N_4989,N_1105,N_1489);
or U4990 (N_4990,N_184,N_2137);
nor U4991 (N_4991,N_878,N_2448);
or U4992 (N_4992,N_2154,N_371);
nand U4993 (N_4993,N_633,N_2116);
nand U4994 (N_4994,N_1471,N_549);
and U4995 (N_4995,N_1484,N_1481);
xor U4996 (N_4996,N_2286,N_2076);
nand U4997 (N_4997,N_406,N_412);
nand U4998 (N_4998,N_1850,N_1813);
nor U4999 (N_4999,N_465,N_1034);
or U5000 (N_5000,N_3847,N_2543);
or U5001 (N_5001,N_3501,N_3185);
or U5002 (N_5002,N_2666,N_4837);
or U5003 (N_5003,N_4139,N_4951);
xor U5004 (N_5004,N_4011,N_3591);
or U5005 (N_5005,N_4599,N_4493);
or U5006 (N_5006,N_3587,N_3671);
nor U5007 (N_5007,N_4087,N_3356);
xor U5008 (N_5008,N_2871,N_2664);
nor U5009 (N_5009,N_4534,N_3167);
nand U5010 (N_5010,N_2514,N_3786);
nor U5011 (N_5011,N_4147,N_4044);
and U5012 (N_5012,N_3498,N_3808);
or U5013 (N_5013,N_3239,N_3720);
nor U5014 (N_5014,N_4145,N_3870);
nor U5015 (N_5015,N_4926,N_3863);
nand U5016 (N_5016,N_2857,N_3445);
nor U5017 (N_5017,N_3419,N_4201);
or U5018 (N_5018,N_3363,N_4971);
nand U5019 (N_5019,N_4385,N_4670);
and U5020 (N_5020,N_2650,N_4866);
and U5021 (N_5021,N_4227,N_3288);
xor U5022 (N_5022,N_2604,N_4880);
or U5023 (N_5023,N_4252,N_2715);
nand U5024 (N_5024,N_4047,N_4914);
nor U5025 (N_5025,N_4715,N_3007);
nand U5026 (N_5026,N_2959,N_3281);
or U5027 (N_5027,N_4787,N_3509);
nor U5028 (N_5028,N_3451,N_4104);
and U5029 (N_5029,N_2960,N_4682);
nand U5030 (N_5030,N_4939,N_3276);
and U5031 (N_5031,N_4825,N_2649);
or U5032 (N_5032,N_3506,N_2709);
nand U5033 (N_5033,N_4707,N_4000);
and U5034 (N_5034,N_4968,N_3214);
nand U5035 (N_5035,N_3161,N_4983);
or U5036 (N_5036,N_2587,N_4383);
or U5037 (N_5037,N_2785,N_3066);
and U5038 (N_5038,N_2767,N_3841);
nor U5039 (N_5039,N_4105,N_3289);
nand U5040 (N_5040,N_3751,N_3822);
and U5041 (N_5041,N_4676,N_3758);
or U5042 (N_5042,N_4026,N_4325);
xnor U5043 (N_5043,N_4486,N_4538);
and U5044 (N_5044,N_3658,N_4588);
nand U5045 (N_5045,N_2733,N_3343);
or U5046 (N_5046,N_3206,N_3595);
nor U5047 (N_5047,N_3471,N_4204);
and U5048 (N_5048,N_4378,N_4346);
nor U5049 (N_5049,N_3086,N_3393);
and U5050 (N_5050,N_3902,N_3547);
xor U5051 (N_5051,N_4432,N_3176);
or U5052 (N_5052,N_4527,N_4459);
nor U5053 (N_5053,N_3186,N_4580);
xor U5054 (N_5054,N_2591,N_4053);
and U5055 (N_5055,N_4901,N_3050);
and U5056 (N_5056,N_3064,N_2723);
nor U5057 (N_5057,N_4125,N_4547);
or U5058 (N_5058,N_2845,N_4436);
nor U5059 (N_5059,N_3551,N_4194);
nand U5060 (N_5060,N_4393,N_3963);
or U5061 (N_5061,N_2523,N_3302);
or U5062 (N_5062,N_4350,N_3712);
nand U5063 (N_5063,N_4250,N_3602);
and U5064 (N_5064,N_2758,N_2789);
nand U5065 (N_5065,N_2773,N_2938);
nor U5066 (N_5066,N_4180,N_3006);
and U5067 (N_5067,N_3588,N_2838);
and U5068 (N_5068,N_4769,N_3436);
nand U5069 (N_5069,N_2945,N_4363);
and U5070 (N_5070,N_3949,N_4730);
nand U5071 (N_5071,N_3901,N_4045);
nand U5072 (N_5072,N_3518,N_4594);
and U5073 (N_5073,N_4311,N_4868);
and U5074 (N_5074,N_4111,N_2634);
or U5075 (N_5075,N_2505,N_4131);
and U5076 (N_5076,N_4460,N_4115);
nand U5077 (N_5077,N_3828,N_3269);
nor U5078 (N_5078,N_3839,N_3705);
nor U5079 (N_5079,N_2575,N_4160);
nor U5080 (N_5080,N_2796,N_2512);
or U5081 (N_5081,N_3931,N_4055);
nor U5082 (N_5082,N_4503,N_3265);
nor U5083 (N_5083,N_4631,N_2724);
nor U5084 (N_5084,N_3494,N_3654);
or U5085 (N_5085,N_4351,N_4326);
xnor U5086 (N_5086,N_2783,N_2521);
nand U5087 (N_5087,N_4354,N_4470);
nor U5088 (N_5088,N_2896,N_4638);
and U5089 (N_5089,N_4724,N_4620);
nor U5090 (N_5090,N_4415,N_2995);
nand U5091 (N_5091,N_4543,N_4618);
and U5092 (N_5092,N_2574,N_4709);
and U5093 (N_5093,N_3369,N_4211);
nor U5094 (N_5094,N_3775,N_3562);
xnor U5095 (N_5095,N_3051,N_3908);
or U5096 (N_5096,N_4826,N_2772);
and U5097 (N_5097,N_2595,N_2668);
nor U5098 (N_5098,N_4226,N_4069);
and U5099 (N_5099,N_3253,N_3296);
and U5100 (N_5100,N_3953,N_3584);
nor U5101 (N_5101,N_3076,N_4161);
nand U5102 (N_5102,N_3464,N_3627);
or U5103 (N_5103,N_3838,N_4058);
and U5104 (N_5104,N_3913,N_3017);
nand U5105 (N_5105,N_3427,N_4895);
and U5106 (N_5106,N_3090,N_3935);
nor U5107 (N_5107,N_3041,N_3643);
and U5108 (N_5108,N_4124,N_4627);
and U5109 (N_5109,N_3065,N_4873);
nor U5110 (N_5110,N_3300,N_3301);
nand U5111 (N_5111,N_3692,N_2606);
nand U5112 (N_5112,N_3976,N_2775);
nor U5113 (N_5113,N_4758,N_4722);
nand U5114 (N_5114,N_3385,N_4217);
nor U5115 (N_5115,N_2781,N_2866);
nor U5116 (N_5116,N_4947,N_4529);
nand U5117 (N_5117,N_3796,N_3073);
and U5118 (N_5118,N_4146,N_4187);
and U5119 (N_5119,N_4987,N_4285);
or U5120 (N_5120,N_4289,N_4213);
nor U5121 (N_5121,N_2588,N_3392);
nand U5122 (N_5122,N_3774,N_3619);
xnor U5123 (N_5123,N_3394,N_2531);
nand U5124 (N_5124,N_3229,N_3083);
and U5125 (N_5125,N_3336,N_3697);
xnor U5126 (N_5126,N_4483,N_4535);
and U5127 (N_5127,N_4335,N_3155);
xor U5128 (N_5128,N_3499,N_3406);
and U5129 (N_5129,N_4672,N_3816);
nor U5130 (N_5130,N_3618,N_2947);
nor U5131 (N_5131,N_3687,N_3340);
xor U5132 (N_5132,N_4280,N_4640);
nor U5133 (N_5133,N_4659,N_4804);
nor U5134 (N_5134,N_2951,N_2788);
or U5135 (N_5135,N_4108,N_3440);
xnor U5136 (N_5136,N_3384,N_4872);
nor U5137 (N_5137,N_4027,N_3803);
nor U5138 (N_5138,N_3271,N_3635);
or U5139 (N_5139,N_2860,N_2834);
and U5140 (N_5140,N_2608,N_4466);
or U5141 (N_5141,N_3761,N_3467);
nand U5142 (N_5142,N_3212,N_3215);
xnor U5143 (N_5143,N_3119,N_3868);
or U5144 (N_5144,N_3071,N_4691);
or U5145 (N_5145,N_2906,N_4428);
nand U5146 (N_5146,N_4288,N_3107);
nor U5147 (N_5147,N_4963,N_3850);
nand U5148 (N_5148,N_4009,N_4566);
or U5149 (N_5149,N_3579,N_2892);
nand U5150 (N_5150,N_2807,N_2889);
nor U5151 (N_5151,N_3171,N_4173);
nand U5152 (N_5152,N_3951,N_4510);
and U5153 (N_5153,N_2822,N_4404);
nand U5154 (N_5154,N_3067,N_3299);
nor U5155 (N_5155,N_4059,N_4673);
nand U5156 (N_5156,N_4696,N_3137);
nor U5157 (N_5157,N_4944,N_4708);
xnor U5158 (N_5158,N_3959,N_3650);
nand U5159 (N_5159,N_3059,N_4266);
nand U5160 (N_5160,N_3663,N_2662);
nor U5161 (N_5161,N_4929,N_3515);
nand U5162 (N_5162,N_3237,N_3315);
nand U5163 (N_5163,N_3946,N_4295);
or U5164 (N_5164,N_3743,N_3057);
and U5165 (N_5165,N_2862,N_2979);
or U5166 (N_5166,N_4746,N_3887);
and U5167 (N_5167,N_2755,N_3603);
nor U5168 (N_5168,N_4384,N_3084);
and U5169 (N_5169,N_4300,N_2519);
xor U5170 (N_5170,N_4005,N_4754);
nor U5171 (N_5171,N_2984,N_4525);
or U5172 (N_5172,N_3319,N_3564);
or U5173 (N_5173,N_3801,N_4581);
or U5174 (N_5174,N_2509,N_3968);
nand U5175 (N_5175,N_4887,N_3347);
or U5176 (N_5176,N_2676,N_4706);
nand U5177 (N_5177,N_4560,N_4001);
or U5178 (N_5178,N_3069,N_4829);
xnor U5179 (N_5179,N_3166,N_4875);
or U5180 (N_5180,N_2501,N_3583);
and U5181 (N_5181,N_2770,N_4847);
xnor U5182 (N_5182,N_3903,N_4487);
nand U5183 (N_5183,N_3972,N_3091);
or U5184 (N_5184,N_2729,N_3306);
xnor U5185 (N_5185,N_4541,N_4070);
nand U5186 (N_5186,N_4228,N_3311);
and U5187 (N_5187,N_2544,N_3827);
or U5188 (N_5188,N_3272,N_3268);
or U5189 (N_5189,N_4723,N_4597);
nand U5190 (N_5190,N_2516,N_3372);
nand U5191 (N_5191,N_4156,N_4478);
xor U5192 (N_5192,N_3832,N_2555);
nor U5193 (N_5193,N_3365,N_3157);
nor U5194 (N_5194,N_2560,N_3438);
nand U5195 (N_5195,N_3975,N_3893);
nand U5196 (N_5196,N_2637,N_3552);
nand U5197 (N_5197,N_4342,N_3566);
nor U5198 (N_5198,N_3505,N_3492);
or U5199 (N_5199,N_3804,N_4553);
xor U5200 (N_5200,N_4773,N_3273);
xnor U5201 (N_5201,N_3628,N_4406);
and U5202 (N_5202,N_3548,N_4817);
or U5203 (N_5203,N_3560,N_4743);
xnor U5204 (N_5204,N_4562,N_3230);
nand U5205 (N_5205,N_2554,N_4761);
or U5206 (N_5206,N_4141,N_2759);
nor U5207 (N_5207,N_3495,N_4686);
or U5208 (N_5208,N_4776,N_3715);
nor U5209 (N_5209,N_4035,N_3355);
nor U5210 (N_5210,N_2869,N_4034);
or U5211 (N_5211,N_2811,N_3741);
and U5212 (N_5212,N_3207,N_3383);
or U5213 (N_5213,N_4348,N_2943);
nand U5214 (N_5214,N_2875,N_2748);
nand U5215 (N_5215,N_2687,N_3811);
and U5216 (N_5216,N_4996,N_2966);
nor U5217 (N_5217,N_2846,N_4593);
and U5218 (N_5218,N_3632,N_4972);
or U5219 (N_5219,N_3459,N_4559);
nor U5220 (N_5220,N_3189,N_4570);
nor U5221 (N_5221,N_2702,N_4595);
nor U5222 (N_5222,N_3213,N_4511);
nor U5223 (N_5223,N_3681,N_4123);
nor U5224 (N_5224,N_2779,N_4729);
and U5225 (N_5225,N_4297,N_3134);
nand U5226 (N_5226,N_4995,N_2734);
nor U5227 (N_5227,N_3797,N_4279);
nand U5228 (N_5228,N_2526,N_4809);
and U5229 (N_5229,N_3001,N_3318);
nor U5230 (N_5230,N_3694,N_4813);
nand U5231 (N_5231,N_3631,N_2593);
nand U5232 (N_5232,N_3196,N_2562);
and U5233 (N_5233,N_4109,N_2534);
or U5234 (N_5234,N_3104,N_4172);
nor U5235 (N_5235,N_3942,N_4544);
nand U5236 (N_5236,N_2944,N_4867);
or U5237 (N_5237,N_4048,N_4750);
and U5238 (N_5238,N_3918,N_2753);
xor U5239 (N_5239,N_3139,N_3449);
and U5240 (N_5240,N_3922,N_4438);
or U5241 (N_5241,N_3826,N_4355);
nor U5242 (N_5242,N_3993,N_4003);
and U5243 (N_5243,N_3981,N_3937);
and U5244 (N_5244,N_4231,N_4292);
nor U5245 (N_5245,N_3063,N_3800);
or U5246 (N_5246,N_2571,N_3753);
nand U5247 (N_5247,N_4666,N_2828);
or U5248 (N_5248,N_3991,N_3553);
nor U5249 (N_5249,N_3188,N_3874);
nor U5250 (N_5250,N_4653,N_4451);
nor U5251 (N_5251,N_4100,N_4306);
or U5252 (N_5252,N_2747,N_2712);
nor U5253 (N_5253,N_3228,N_4361);
nor U5254 (N_5254,N_4241,N_3485);
nor U5255 (N_5255,N_4775,N_3648);
xor U5256 (N_5256,N_3244,N_2617);
nor U5257 (N_5257,N_2527,N_3367);
nor U5258 (N_5258,N_3864,N_2970);
or U5259 (N_5259,N_4032,N_3245);
nor U5260 (N_5260,N_2583,N_3928);
nor U5261 (N_5261,N_2814,N_2589);
and U5262 (N_5262,N_3790,N_3487);
or U5263 (N_5263,N_3201,N_4596);
xnor U5264 (N_5264,N_3008,N_2752);
nor U5265 (N_5265,N_3373,N_4814);
nand U5266 (N_5266,N_3018,N_3033);
nand U5267 (N_5267,N_3056,N_4853);
or U5268 (N_5268,N_2953,N_3594);
or U5269 (N_5269,N_4565,N_4705);
xnor U5270 (N_5270,N_2518,N_4993);
nand U5271 (N_5271,N_2809,N_3014);
xor U5272 (N_5272,N_4029,N_3368);
nor U5273 (N_5273,N_4396,N_4677);
nand U5274 (N_5274,N_3439,N_4907);
or U5275 (N_5275,N_3223,N_3558);
or U5276 (N_5276,N_4688,N_3128);
or U5277 (N_5277,N_4422,N_2533);
and U5278 (N_5278,N_4891,N_4423);
and U5279 (N_5279,N_3251,N_3909);
or U5280 (N_5280,N_3752,N_2539);
nand U5281 (N_5281,N_4121,N_4084);
nor U5282 (N_5282,N_4749,N_4976);
and U5283 (N_5283,N_3667,N_3535);
xor U5284 (N_5284,N_3873,N_3813);
nand U5285 (N_5285,N_3335,N_4685);
nor U5286 (N_5286,N_4421,N_4196);
nand U5287 (N_5287,N_4756,N_4790);
and U5288 (N_5288,N_4894,N_4992);
nand U5289 (N_5289,N_3825,N_4695);
nor U5290 (N_5290,N_4382,N_4941);
or U5291 (N_5291,N_3749,N_4540);
or U5292 (N_5292,N_4293,N_3433);
nor U5293 (N_5293,N_3794,N_4073);
and U5294 (N_5294,N_4892,N_2751);
or U5295 (N_5295,N_4469,N_4800);
xnor U5296 (N_5296,N_3995,N_3576);
nand U5297 (N_5297,N_4392,N_4785);
and U5298 (N_5298,N_4357,N_3361);
or U5299 (N_5299,N_3224,N_4925);
and U5300 (N_5300,N_3397,N_4924);
or U5301 (N_5301,N_3103,N_3755);
nor U5302 (N_5302,N_3747,N_3293);
and U5303 (N_5303,N_3160,N_4259);
and U5304 (N_5304,N_3719,N_4683);
or U5305 (N_5305,N_4626,N_4513);
nor U5306 (N_5306,N_4919,N_2806);
nand U5307 (N_5307,N_4747,N_4616);
nand U5308 (N_5308,N_3162,N_4964);
nand U5309 (N_5309,N_3112,N_2618);
or U5310 (N_5310,N_3305,N_3403);
or U5311 (N_5311,N_3641,N_4917);
or U5312 (N_5312,N_4054,N_3982);
or U5313 (N_5313,N_4352,N_2663);
and U5314 (N_5314,N_3012,N_3136);
or U5315 (N_5315,N_3899,N_2909);
nor U5316 (N_5316,N_4879,N_2754);
nand U5317 (N_5317,N_2642,N_3570);
xor U5318 (N_5318,N_4978,N_4835);
nand U5319 (N_5319,N_3470,N_4797);
xnor U5320 (N_5320,N_3364,N_3525);
or U5321 (N_5321,N_3225,N_3733);
or U5322 (N_5322,N_4248,N_2961);
or U5323 (N_5323,N_3173,N_3082);
nor U5324 (N_5324,N_3197,N_3200);
and U5325 (N_5325,N_3074,N_2898);
or U5326 (N_5326,N_3195,N_2999);
xor U5327 (N_5327,N_4766,N_2631);
or U5328 (N_5328,N_3483,N_3170);
or U5329 (N_5329,N_3731,N_3737);
nand U5330 (N_5330,N_2852,N_3938);
nand U5331 (N_5331,N_4943,N_2873);
nand U5332 (N_5332,N_4229,N_3612);
nand U5333 (N_5333,N_2992,N_3691);
nand U5334 (N_5334,N_4374,N_4886);
nand U5335 (N_5335,N_2675,N_4237);
and U5336 (N_5336,N_2937,N_3652);
nand U5337 (N_5337,N_4025,N_2812);
or U5338 (N_5338,N_4358,N_4186);
nand U5339 (N_5339,N_4712,N_4262);
xnor U5340 (N_5340,N_4302,N_3855);
nand U5341 (N_5341,N_2952,N_2877);
nor U5342 (N_5342,N_3567,N_3290);
nand U5343 (N_5343,N_4198,N_3629);
nor U5344 (N_5344,N_3117,N_3405);
xor U5345 (N_5345,N_2647,N_3198);
and U5346 (N_5346,N_4270,N_2780);
and U5347 (N_5347,N_4772,N_3545);
or U5348 (N_5348,N_3930,N_4613);
nand U5349 (N_5349,N_2703,N_4657);
or U5350 (N_5350,N_4450,N_2586);
nor U5351 (N_5351,N_3590,N_4757);
nor U5352 (N_5352,N_4786,N_3354);
nand U5353 (N_5353,N_3099,N_4341);
or U5354 (N_5354,N_2965,N_4607);
nand U5355 (N_5355,N_4251,N_2594);
and U5356 (N_5356,N_3651,N_2762);
nand U5357 (N_5357,N_3280,N_2671);
nor U5358 (N_5358,N_2599,N_4744);
or U5359 (N_5359,N_4619,N_3413);
and U5360 (N_5360,N_3573,N_3118);
nor U5361 (N_5361,N_4665,N_4737);
or U5362 (N_5362,N_4497,N_4689);
xnor U5363 (N_5363,N_3709,N_2602);
and U5364 (N_5364,N_4654,N_4359);
and U5365 (N_5365,N_2918,N_2613);
and U5366 (N_5366,N_4449,N_3925);
nor U5367 (N_5367,N_4651,N_4871);
or U5368 (N_5368,N_4549,N_3061);
or U5369 (N_5369,N_3482,N_3002);
nand U5370 (N_5370,N_3582,N_4182);
or U5371 (N_5371,N_3138,N_3912);
nor U5372 (N_5372,N_4479,N_3236);
nand U5373 (N_5373,N_2769,N_3689);
and U5374 (N_5374,N_3757,N_4608);
and U5375 (N_5375,N_4782,N_3154);
nand U5376 (N_5376,N_3662,N_4253);
nor U5377 (N_5377,N_3530,N_3539);
nand U5378 (N_5378,N_3060,N_4759);
nand U5379 (N_5379,N_2749,N_2743);
nor U5380 (N_5380,N_2645,N_3295);
nand U5381 (N_5381,N_3914,N_3115);
or U5382 (N_5382,N_4751,N_3606);
or U5383 (N_5383,N_4883,N_3123);
nor U5384 (N_5384,N_3325,N_3219);
nor U5385 (N_5385,N_3852,N_4795);
and U5386 (N_5386,N_4148,N_4504);
nand U5387 (N_5387,N_4079,N_3164);
nand U5388 (N_5388,N_3054,N_3202);
or U5389 (N_5389,N_4681,N_3423);
or U5390 (N_5390,N_3572,N_2745);
nor U5391 (N_5391,N_3789,N_3399);
nand U5392 (N_5392,N_2651,N_4441);
or U5393 (N_5393,N_4063,N_3145);
nor U5394 (N_5394,N_3542,N_4010);
nand U5395 (N_5395,N_4485,N_4434);
or U5396 (N_5396,N_3969,N_3298);
nand U5397 (N_5397,N_3638,N_4379);
and U5398 (N_5398,N_2736,N_2946);
nor U5399 (N_5399,N_3520,N_3221);
nor U5400 (N_5400,N_4836,N_4905);
nor U5401 (N_5401,N_2682,N_4071);
and U5402 (N_5402,N_3131,N_2927);
nand U5403 (N_5403,N_2967,N_3819);
and U5404 (N_5404,N_3983,N_4684);
xnor U5405 (N_5405,N_2503,N_4427);
nor U5406 (N_5406,N_3127,N_2901);
or U5407 (N_5407,N_2528,N_4575);
or U5408 (N_5408,N_3835,N_4090);
nor U5409 (N_5409,N_3777,N_4212);
and U5410 (N_5410,N_3916,N_4448);
or U5411 (N_5411,N_3994,N_2830);
nor U5412 (N_5412,N_4224,N_3058);
nor U5413 (N_5413,N_4395,N_3313);
or U5414 (N_5414,N_4661,N_3932);
nand U5415 (N_5415,N_4360,N_3146);
or U5416 (N_5416,N_3611,N_3622);
and U5417 (N_5417,N_3782,N_2737);
or U5418 (N_5418,N_3661,N_4630);
and U5419 (N_5419,N_2919,N_4416);
or U5420 (N_5420,N_3317,N_3872);
and U5421 (N_5421,N_4419,N_4309);
nor U5422 (N_5422,N_4037,N_3585);
or U5423 (N_5423,N_2530,N_4642);
and U5424 (N_5424,N_3607,N_4014);
and U5425 (N_5425,N_2686,N_3701);
nand U5426 (N_5426,N_2854,N_2988);
nor U5427 (N_5427,N_3260,N_3675);
nand U5428 (N_5428,N_2654,N_4962);
nand U5429 (N_5429,N_4126,N_2700);
and U5430 (N_5430,N_2764,N_4694);
nand U5431 (N_5431,N_3665,N_4845);
nor U5432 (N_5432,N_4304,N_3400);
nand U5433 (N_5433,N_4337,N_2532);
nand U5434 (N_5434,N_3025,N_3831);
or U5435 (N_5435,N_3389,N_3806);
and U5436 (N_5436,N_2685,N_3209);
or U5437 (N_5437,N_3177,N_4663);
or U5438 (N_5438,N_2794,N_2547);
and U5439 (N_5439,N_4430,N_2815);
nor U5440 (N_5440,N_4265,N_2688);
nor U5441 (N_5441,N_3324,N_3407);
nor U5442 (N_5442,N_4999,N_3532);
nor U5443 (N_5443,N_3586,N_3783);
nor U5444 (N_5444,N_4457,N_3881);
nand U5445 (N_5445,N_4465,N_4937);
nand U5446 (N_5446,N_2884,N_4366);
nand U5447 (N_5447,N_4509,N_3358);
or U5448 (N_5448,N_3149,N_4220);
nor U5449 (N_5449,N_3754,N_3756);
nor U5450 (N_5450,N_2673,N_3234);
nand U5451 (N_5451,N_2707,N_2930);
and U5452 (N_5452,N_4846,N_3070);
xor U5453 (N_5453,N_3517,N_2585);
and U5454 (N_5454,N_4664,N_3500);
or U5455 (N_5455,N_4656,N_4247);
or U5456 (N_5456,N_3860,N_4328);
or U5457 (N_5457,N_3792,N_2697);
or U5458 (N_5458,N_4343,N_4961);
or U5459 (N_5459,N_4958,N_2908);
or U5460 (N_5460,N_4710,N_3217);
nor U5461 (N_5461,N_4208,N_3152);
and U5462 (N_5462,N_2925,N_4046);
xnor U5463 (N_5463,N_3646,N_2706);
nor U5464 (N_5464,N_3488,N_2566);
nor U5465 (N_5465,N_2972,N_3574);
nand U5466 (N_5466,N_3078,N_4455);
and U5467 (N_5467,N_3763,N_4946);
nor U5468 (N_5468,N_4557,N_2643);
or U5469 (N_5469,N_2922,N_3966);
nor U5470 (N_5470,N_4051,N_2831);
nor U5471 (N_5471,N_4942,N_2541);
and U5472 (N_5472,N_4704,N_4974);
or U5473 (N_5473,N_2558,N_3528);
nand U5474 (N_5474,N_4519,N_3254);
nor U5475 (N_5475,N_4163,N_4521);
or U5476 (N_5476,N_3921,N_2810);
and U5477 (N_5477,N_3088,N_2782);
and U5478 (N_5478,N_3259,N_2717);
and U5479 (N_5479,N_2552,N_2893);
nand U5480 (N_5480,N_3843,N_3817);
or U5481 (N_5481,N_3604,N_3140);
or U5482 (N_5482,N_2716,N_3767);
nand U5483 (N_5483,N_2926,N_3917);
or U5484 (N_5484,N_2982,N_4823);
nand U5485 (N_5485,N_2941,N_2843);
nand U5486 (N_5486,N_3571,N_3247);
nor U5487 (N_5487,N_3342,N_3894);
or U5488 (N_5488,N_4878,N_4874);
nand U5489 (N_5489,N_2610,N_4870);
nand U5490 (N_5490,N_4796,N_3546);
or U5491 (N_5491,N_4429,N_2517);
or U5492 (N_5492,N_4098,N_4331);
or U5493 (N_5493,N_2590,N_4721);
or U5494 (N_5494,N_4036,N_3204);
and U5495 (N_5495,N_2568,N_3022);
nor U5496 (N_5496,N_2962,N_4426);
xnor U5497 (N_5497,N_4556,N_3954);
xnor U5498 (N_5498,N_4505,N_2768);
nor U5499 (N_5499,N_4784,N_3746);
and U5500 (N_5500,N_3890,N_2600);
and U5501 (N_5501,N_4008,N_3442);
nor U5502 (N_5502,N_3821,N_4542);
xnor U5503 (N_5503,N_4548,N_3113);
or U5504 (N_5504,N_4893,N_4902);
nand U5505 (N_5505,N_3793,N_4377);
and U5506 (N_5506,N_2730,N_4023);
and U5507 (N_5507,N_3906,N_3609);
or U5508 (N_5508,N_2894,N_4339);
or U5509 (N_5509,N_2868,N_4731);
nor U5510 (N_5510,N_4533,N_3729);
and U5511 (N_5511,N_4243,N_2548);
and U5512 (N_5512,N_4407,N_3538);
nor U5513 (N_5513,N_2787,N_4305);
and U5514 (N_5514,N_3941,N_3267);
nand U5515 (N_5515,N_2994,N_3504);
and U5516 (N_5516,N_2955,N_4985);
xnor U5517 (N_5517,N_4365,N_2524);
or U5518 (N_5518,N_3307,N_3610);
or U5519 (N_5519,N_3460,N_4906);
nand U5520 (N_5520,N_4516,N_4904);
xnor U5521 (N_5521,N_3208,N_4110);
xnor U5522 (N_5522,N_2832,N_3926);
or U5523 (N_5523,N_4839,N_4477);
and U5524 (N_5524,N_4072,N_2958);
or U5525 (N_5525,N_3434,N_4822);
or U5526 (N_5526,N_4601,N_3333);
xnor U5527 (N_5527,N_3316,N_4499);
xnor U5528 (N_5528,N_2626,N_4550);
or U5529 (N_5529,N_2720,N_2880);
and U5530 (N_5530,N_2542,N_4162);
and U5531 (N_5531,N_3258,N_2813);
and U5532 (N_5532,N_3042,N_4118);
nor U5533 (N_5533,N_4316,N_3910);
nor U5534 (N_5534,N_2861,N_4203);
or U5535 (N_5535,N_2538,N_2818);
nand U5536 (N_5536,N_4498,N_4889);
xnor U5537 (N_5537,N_2656,N_3190);
xnor U5538 (N_5538,N_4913,N_4492);
nand U5539 (N_5539,N_4838,N_4698);
nand U5540 (N_5540,N_3559,N_4202);
and U5541 (N_5541,N_4372,N_3948);
and U5542 (N_5542,N_4320,N_3220);
and U5543 (N_5543,N_3980,N_3334);
nand U5544 (N_5544,N_3072,N_3444);
and U5545 (N_5545,N_3100,N_4514);
nor U5546 (N_5546,N_3685,N_2933);
nor U5547 (N_5547,N_3462,N_3766);
nand U5548 (N_5548,N_4390,N_3010);
or U5549 (N_5549,N_3352,N_3321);
nand U5550 (N_5550,N_4604,N_3329);
nor U5551 (N_5551,N_3845,N_2742);
nor U5552 (N_5552,N_2850,N_2990);
nor U5553 (N_5553,N_2974,N_4291);
nor U5554 (N_5554,N_3762,N_3446);
nand U5555 (N_5555,N_3391,N_4727);
nand U5556 (N_5556,N_3376,N_4020);
and U5557 (N_5557,N_3799,N_3896);
and U5558 (N_5558,N_3669,N_4068);
or U5559 (N_5559,N_2652,N_2678);
nor U5560 (N_5560,N_4649,N_4957);
or U5561 (N_5561,N_4473,N_3366);
nand U5562 (N_5562,N_3659,N_3029);
nor U5563 (N_5563,N_4512,N_3895);
or U5564 (N_5564,N_3911,N_3344);
nor U5565 (N_5565,N_3348,N_4984);
or U5566 (N_5566,N_2867,N_4235);
or U5567 (N_5567,N_3718,N_4674);
or U5568 (N_5568,N_3156,N_4127);
nand U5569 (N_5569,N_2540,N_4197);
and U5570 (N_5570,N_3653,N_4274);
and U5571 (N_5571,N_3772,N_4474);
nand U5572 (N_5572,N_2551,N_3600);
nand U5573 (N_5573,N_3802,N_4007);
nand U5574 (N_5574,N_2739,N_4155);
and U5575 (N_5575,N_3401,N_4107);
nand U5576 (N_5576,N_4129,N_2612);
or U5577 (N_5577,N_3011,N_2816);
nor U5578 (N_5578,N_3274,N_3235);
or U5579 (N_5579,N_2506,N_4960);
nand U5580 (N_5580,N_4517,N_2969);
or U5581 (N_5581,N_2525,N_4792);
xnor U5582 (N_5582,N_4832,N_4307);
or U5583 (N_5583,N_4269,N_2607);
or U5584 (N_5584,N_3292,N_2580);
and U5585 (N_5585,N_3277,N_3454);
xnor U5586 (N_5586,N_2504,N_2907);
and U5587 (N_5587,N_4840,N_4471);
and U5588 (N_5588,N_3780,N_4959);
or U5589 (N_5589,N_3770,N_3867);
xnor U5590 (N_5590,N_3469,N_3851);
or U5591 (N_5591,N_3698,N_3266);
or U5592 (N_5592,N_4934,N_4452);
or U5593 (N_5593,N_2765,N_3047);
or U5594 (N_5594,N_3519,N_4169);
nor U5595 (N_5595,N_2954,N_2971);
nand U5596 (N_5596,N_3032,N_4066);
and U5597 (N_5597,N_2680,N_2732);
or U5598 (N_5598,N_4523,N_3544);
or U5599 (N_5599,N_4848,N_4828);
xor U5600 (N_5600,N_4060,N_4799);
nand U5601 (N_5601,N_4568,N_4388);
nor U5602 (N_5602,N_3668,N_4501);
xnor U5603 (N_5603,N_3168,N_3818);
xnor U5604 (N_5604,N_4668,N_3973);
and U5605 (N_5605,N_3889,N_4149);
nand U5606 (N_5606,N_4494,N_4998);
and U5607 (N_5607,N_3456,N_2856);
xnor U5608 (N_5608,N_3891,N_4461);
xnor U5609 (N_5609,N_3479,N_4635);
nand U5610 (N_5610,N_3048,N_4719);
or U5611 (N_5611,N_3106,N_3481);
xor U5612 (N_5612,N_3785,N_3357);
xnor U5613 (N_5613,N_4778,N_3093);
nand U5614 (N_5614,N_4134,N_2620);
nand U5615 (N_5615,N_4445,N_3143);
and U5616 (N_5616,N_3349,N_4603);
or U5617 (N_5617,N_3095,N_2929);
nand U5618 (N_5618,N_4258,N_3523);
and U5619 (N_5619,N_4765,N_4935);
nor U5620 (N_5620,N_3634,N_3879);
xnor U5621 (N_5621,N_2557,N_4592);
nor U5622 (N_5622,N_4590,N_3987);
and U5623 (N_5623,N_2728,N_2916);
or U5624 (N_5624,N_2840,N_3526);
nand U5625 (N_5625,N_3374,N_4271);
nand U5626 (N_5626,N_4779,N_4210);
nor U5627 (N_5627,N_3416,N_4815);
nor U5628 (N_5628,N_4353,N_2690);
or U5629 (N_5629,N_4818,N_4082);
nor U5630 (N_5630,N_4555,N_3323);
nand U5631 (N_5631,N_2644,N_3779);
and U5632 (N_5632,N_4798,N_4387);
and U5633 (N_5633,N_4482,N_3278);
or U5634 (N_5634,N_3110,N_4621);
or U5635 (N_5635,N_4057,N_3647);
nor U5636 (N_5636,N_4854,N_4536);
nor U5637 (N_5637,N_4859,N_4515);
or U5638 (N_5638,N_2885,N_4281);
and U5639 (N_5639,N_4344,N_4639);
xnor U5640 (N_5640,N_3933,N_3960);
or U5641 (N_5641,N_3837,N_2819);
nand U5642 (N_5642,N_3700,N_2903);
nor U5643 (N_5643,N_3417,N_3997);
nand U5644 (N_5644,N_3534,N_3568);
or U5645 (N_5645,N_4327,N_4329);
nor U5646 (N_5646,N_2872,N_3861);
nor U5647 (N_5647,N_4193,N_2790);
nand U5648 (N_5648,N_3053,N_3569);
xnor U5649 (N_5649,N_2956,N_4373);
nor U5650 (N_5650,N_4791,N_3764);
nor U5651 (N_5651,N_2839,N_4140);
or U5652 (N_5652,N_4178,N_4244);
or U5653 (N_5653,N_3513,N_2855);
or U5654 (N_5654,N_4089,N_3129);
nand U5655 (N_5655,N_3153,N_4600);
or U5656 (N_5656,N_3836,N_3727);
xnor U5657 (N_5657,N_4317,N_2546);
nor U5658 (N_5658,N_4425,N_2598);
nand U5659 (N_5659,N_4572,N_2750);
or U5660 (N_5660,N_4065,N_4417);
or U5661 (N_5661,N_3452,N_4238);
and U5662 (N_5662,N_3771,N_4380);
and U5663 (N_5663,N_3502,N_4692);
or U5664 (N_5664,N_2837,N_3408);
xor U5665 (N_5665,N_4966,N_4234);
and U5666 (N_5666,N_2741,N_3723);
or U5667 (N_5667,N_4184,N_4012);
nand U5668 (N_5668,N_4074,N_4770);
nand U5669 (N_5669,N_4701,N_3592);
nor U5670 (N_5670,N_2520,N_3508);
nor U5671 (N_5671,N_4783,N_4805);
nand U5672 (N_5672,N_2576,N_4154);
nand U5673 (N_5673,N_4700,N_4464);
or U5674 (N_5674,N_4323,N_4816);
nor U5675 (N_5675,N_3387,N_4881);
nor U5676 (N_5676,N_3003,N_2567);
or U5677 (N_5677,N_4591,N_3684);
and U5678 (N_5678,N_2510,N_2823);
or U5679 (N_5679,N_3805,N_4830);
nand U5680 (N_5680,N_4130,N_3285);
nor U5681 (N_5681,N_2628,N_4539);
and U5682 (N_5682,N_3561,N_3122);
xor U5683 (N_5683,N_4083,N_3089);
xnor U5684 (N_5684,N_4117,N_4199);
nand U5685 (N_5685,N_3927,N_3605);
and U5686 (N_5686,N_3484,N_4368);
nand U5687 (N_5687,N_2923,N_4043);
xor U5688 (N_5688,N_2978,N_2963);
nor U5689 (N_5689,N_2719,N_4056);
xor U5690 (N_5690,N_4143,N_4039);
or U5691 (N_5691,N_2853,N_3175);
and U5692 (N_5692,N_4741,N_2572);
nand U5693 (N_5693,N_3614,N_2507);
nor U5694 (N_5694,N_3283,N_4850);
or U5695 (N_5695,N_3322,N_4855);
nand U5696 (N_5696,N_3536,N_3016);
nor U5697 (N_5697,N_2756,N_4246);
nand U5698 (N_5698,N_3680,N_3414);
or U5699 (N_5699,N_3578,N_3810);
nand U5700 (N_5700,N_3615,N_3232);
and U5701 (N_5701,N_4577,N_2973);
and U5702 (N_5702,N_4970,N_2985);
or U5703 (N_5703,N_3013,N_4249);
nand U5704 (N_5704,N_4582,N_3765);
and U5705 (N_5705,N_4114,N_2777);
nand U5706 (N_5706,N_4132,N_4456);
nand U5707 (N_5707,N_3026,N_3341);
nand U5708 (N_5708,N_3141,N_3351);
nor U5709 (N_5709,N_3130,N_4345);
or U5710 (N_5710,N_2792,N_3345);
and U5711 (N_5711,N_4006,N_3249);
nor U5712 (N_5712,N_4738,N_3453);
nand U5713 (N_5713,N_4400,N_2914);
and U5714 (N_5714,N_4702,N_2699);
or U5715 (N_5715,N_3241,N_4435);
or U5716 (N_5716,N_3092,N_2910);
or U5717 (N_5717,N_4444,N_3672);
xnor U5718 (N_5718,N_2681,N_4586);
xor U5719 (N_5719,N_4192,N_4697);
and U5720 (N_5720,N_2592,N_3732);
or U5721 (N_5721,N_3279,N_4732);
nand U5722 (N_5722,N_3540,N_2847);
xor U5723 (N_5723,N_2627,N_3144);
nand U5724 (N_5724,N_4567,N_4257);
nand U5725 (N_5725,N_3286,N_2817);
and U5726 (N_5726,N_4762,N_3039);
nand U5727 (N_5727,N_3098,N_2603);
nand U5728 (N_5728,N_2611,N_3420);
nand U5729 (N_5729,N_4067,N_4965);
or U5730 (N_5730,N_3989,N_4909);
or U5731 (N_5731,N_4877,N_4050);
nand U5732 (N_5732,N_4038,N_3725);
or U5733 (N_5733,N_3121,N_4506);
nand U5734 (N_5734,N_4119,N_2932);
and U5735 (N_5735,N_3477,N_2820);
and U5736 (N_5736,N_3330,N_4956);
and U5737 (N_5737,N_4641,N_3320);
xnor U5738 (N_5738,N_3900,N_2989);
and U5739 (N_5739,N_3380,N_2549);
or U5740 (N_5740,N_3437,N_2888);
nor U5741 (N_5741,N_4205,N_4347);
nor U5742 (N_5742,N_4578,N_3965);
and U5743 (N_5743,N_4233,N_4820);
and U5744 (N_5744,N_2508,N_3848);
nor U5745 (N_5745,N_4076,N_2581);
nand U5746 (N_5746,N_3589,N_4078);
nor U5747 (N_5747,N_4605,N_4864);
nor U5748 (N_5748,N_4954,N_2537);
nand U5749 (N_5749,N_4322,N_3049);
nor U5750 (N_5750,N_3180,N_3111);
or U5751 (N_5751,N_3956,N_2874);
xor U5752 (N_5752,N_3402,N_3284);
nor U5753 (N_5753,N_2711,N_3183);
and U5754 (N_5754,N_3978,N_4189);
and U5755 (N_5755,N_4411,N_4748);
or U5756 (N_5756,N_3915,N_2609);
or U5757 (N_5757,N_2949,N_4106);
xnor U5758 (N_5758,N_3620,N_2596);
nor U5759 (N_5759,N_2529,N_4860);
and U5760 (N_5760,N_2698,N_4440);
or U5761 (N_5761,N_3310,N_4819);
xor U5762 (N_5762,N_4190,N_4015);
or U5763 (N_5763,N_4255,N_4648);
nor U5764 (N_5764,N_2760,N_3529);
nor U5765 (N_5765,N_3448,N_4589);
nand U5766 (N_5766,N_3472,N_3639);
nand U5767 (N_5767,N_3187,N_4221);
xor U5768 (N_5768,N_4116,N_4940);
and U5769 (N_5769,N_4980,N_4138);
and U5770 (N_5770,N_4174,N_2597);
or U5771 (N_5771,N_4164,N_3699);
and U5772 (N_5772,N_4097,N_3812);
nor U5773 (N_5773,N_4953,N_3939);
or U5774 (N_5774,N_3326,N_4170);
nand U5775 (N_5775,N_3934,N_4583);
or U5776 (N_5776,N_3522,N_2913);
and U5777 (N_5777,N_3625,N_4997);
nor U5778 (N_5778,N_4254,N_3759);
or U5779 (N_5779,N_4077,N_2891);
and U5780 (N_5780,N_3248,N_4101);
nand U5781 (N_5781,N_4447,N_2900);
or U5782 (N_5782,N_2624,N_3182);
or U5783 (N_5783,N_3346,N_4200);
and U5784 (N_5784,N_4086,N_4475);
xor U5785 (N_5785,N_2605,N_4061);
or U5786 (N_5786,N_4080,N_3984);
nor U5787 (N_5787,N_3036,N_2793);
or U5788 (N_5788,N_4398,N_2653);
and U5789 (N_5789,N_3556,N_4679);
nor U5790 (N_5790,N_3443,N_3728);
or U5791 (N_5791,N_3854,N_4973);
and U5792 (N_5792,N_4481,N_3516);
nand U5793 (N_5793,N_3194,N_3450);
nor U5794 (N_5794,N_4468,N_3637);
nand U5795 (N_5795,N_3418,N_3490);
xor U5796 (N_5796,N_3776,N_3491);
or U5797 (N_5797,N_4214,N_3781);
and U5798 (N_5798,N_3308,N_2563);
or U5799 (N_5799,N_4643,N_4041);
or U5800 (N_5800,N_3216,N_3824);
xor U5801 (N_5801,N_3998,N_4381);
and U5802 (N_5802,N_4617,N_4781);
xnor U5803 (N_5803,N_3608,N_4564);
nand U5804 (N_5804,N_4720,N_3875);
nor U5805 (N_5805,N_2667,N_4718);
xor U5806 (N_5806,N_3596,N_3884);
nor U5807 (N_5807,N_4780,N_3422);
nand U5808 (N_5808,N_2646,N_4611);
xor U5809 (N_5809,N_3205,N_3846);
and U5810 (N_5810,N_3958,N_4882);
nand U5811 (N_5811,N_3359,N_3486);
or U5812 (N_5812,N_3426,N_2935);
and U5813 (N_5813,N_2648,N_2658);
nand U5814 (N_5814,N_2964,N_4443);
and U5815 (N_5815,N_4209,N_4897);
and U5816 (N_5816,N_4167,N_3097);
and U5817 (N_5817,N_3882,N_3222);
and U5818 (N_5818,N_3878,N_3303);
nand U5819 (N_5819,N_3945,N_2774);
or U5820 (N_5820,N_3382,N_2936);
nand U5821 (N_5821,N_2713,N_4662);
nor U5822 (N_5822,N_3711,N_3642);
nand U5823 (N_5823,N_2826,N_3503);
nand U5824 (N_5824,N_4166,N_3199);
and U5825 (N_5825,N_4725,N_3888);
nand U5826 (N_5826,N_3673,N_3261);
nor U5827 (N_5827,N_3395,N_3907);
or U5828 (N_5828,N_2740,N_3593);
and U5829 (N_5829,N_3974,N_4095);
nor U5830 (N_5830,N_2500,N_2615);
and U5831 (N_5831,N_3676,N_2535);
or U5832 (N_5832,N_2661,N_4558);
xor U5833 (N_5833,N_3943,N_4264);
nor U5834 (N_5834,N_3327,N_2569);
nor U5835 (N_5835,N_4176,N_4310);
nand U5836 (N_5836,N_3105,N_4526);
or U5837 (N_5837,N_3114,N_4803);
xnor U5838 (N_5838,N_4502,N_3031);
xnor U5839 (N_5839,N_4898,N_3521);
xor U5840 (N_5840,N_4584,N_3866);
and U5841 (N_5841,N_2696,N_4812);
or U5842 (N_5842,N_3554,N_4981);
or U5843 (N_5843,N_4389,N_2977);
and U5844 (N_5844,N_3601,N_4975);
xnor U5845 (N_5845,N_2691,N_4371);
nor U5846 (N_5846,N_2983,N_4370);
xor U5847 (N_5847,N_2915,N_3717);
nand U5848 (N_5848,N_3985,N_4763);
or U5849 (N_5849,N_4401,N_4742);
and U5850 (N_5850,N_4120,N_3151);
xnor U5851 (N_5851,N_3543,N_4977);
and U5852 (N_5852,N_3964,N_4842);
xnor U5853 (N_5853,N_3905,N_4391);
or U5854 (N_5854,N_2791,N_3613);
nor U5855 (N_5855,N_3563,N_2948);
nor U5856 (N_5856,N_3304,N_4017);
nor U5857 (N_5857,N_4185,N_3079);
and U5858 (N_5858,N_4319,N_3377);
nor U5859 (N_5859,N_4488,N_4408);
nand U5860 (N_5860,N_3688,N_3398);
nor U5861 (N_5861,N_3255,N_4669);
or U5862 (N_5862,N_4496,N_4938);
or U5863 (N_5863,N_3227,N_3883);
xor U5864 (N_5864,N_2996,N_4680);
nand U5865 (N_5865,N_3390,N_3429);
nor U5866 (N_5866,N_3877,N_4561);
and U5867 (N_5867,N_4982,N_2550);
or U5868 (N_5868,N_4927,N_4490);
or U5869 (N_5869,N_3465,N_3706);
and U5870 (N_5870,N_3555,N_2939);
and U5871 (N_5871,N_2912,N_3081);
and U5872 (N_5872,N_4225,N_2895);
xnor U5873 (N_5873,N_4092,N_3169);
xor U5874 (N_5874,N_3557,N_4936);
or U5875 (N_5875,N_3655,N_4177);
and U5876 (N_5876,N_4755,N_2616);
nand U5877 (N_5877,N_3683,N_4952);
nand U5878 (N_5878,N_4933,N_2731);
and U5879 (N_5879,N_4122,N_2899);
and U5880 (N_5880,N_2625,N_3125);
nor U5881 (N_5881,N_4402,N_3435);
or U5882 (N_5882,N_4386,N_4075);
xor U5883 (N_5883,N_4979,N_3080);
or U5884 (N_5884,N_4171,N_3971);
and U5885 (N_5885,N_3421,N_4717);
nor U5886 (N_5886,N_4113,N_2798);
and U5887 (N_5887,N_2640,N_3496);
nor U5888 (N_5888,N_4612,N_3695);
nand U5889 (N_5889,N_4049,N_3193);
or U5890 (N_5890,N_3174,N_2735);
xnor U5891 (N_5891,N_4863,N_2766);
or U5892 (N_5892,N_4085,N_4990);
or U5893 (N_5893,N_3052,N_4865);
and U5894 (N_5894,N_3739,N_4739);
nand U5895 (N_5895,N_2897,N_4801);
nor U5896 (N_5896,N_3455,N_3869);
and U5897 (N_5897,N_3623,N_3537);
nor U5898 (N_5898,N_2689,N_4491);
nor U5899 (N_5899,N_3507,N_4298);
and U5900 (N_5900,N_4633,N_3858);
or U5901 (N_5901,N_4040,N_4849);
and U5902 (N_5902,N_3876,N_3988);
and U5903 (N_5903,N_4852,N_4336);
xor U5904 (N_5904,N_4645,N_3704);
and U5905 (N_5905,N_4303,N_3674);
or U5906 (N_5906,N_4467,N_2674);
nor U5907 (N_5907,N_4753,N_4520);
nand U5908 (N_5908,N_2695,N_4195);
or U5909 (N_5909,N_2621,N_4667);
and U5910 (N_5910,N_2887,N_2511);
and U5911 (N_5911,N_3740,N_3430);
or U5912 (N_5912,N_4287,N_4312);
and U5913 (N_5913,N_3203,N_3809);
xnor U5914 (N_5914,N_4165,N_3386);
nand U5915 (N_5915,N_4318,N_4437);
nor U5916 (N_5916,N_3024,N_2950);
nor U5917 (N_5917,N_2848,N_4267);
and U5918 (N_5918,N_3807,N_3885);
and U5919 (N_5919,N_4168,N_3378);
nand U5920 (N_5920,N_4207,N_4531);
nand U5921 (N_5921,N_3970,N_3035);
nor U5922 (N_5922,N_4239,N_2863);
nor U5923 (N_5923,N_4042,N_3246);
and U5924 (N_5924,N_4576,N_2836);
or U5925 (N_5925,N_4308,N_4841);
nor U5926 (N_5926,N_3742,N_4019);
or U5927 (N_5927,N_4183,N_4230);
or U5928 (N_5928,N_3524,N_3085);
nand U5929 (N_5929,N_3859,N_4690);
xor U5930 (N_5930,N_3497,N_3120);
nand U5931 (N_5931,N_3730,N_4236);
or U5932 (N_5932,N_3238,N_4314);
and U5933 (N_5933,N_2940,N_4918);
xnor U5934 (N_5934,N_3833,N_4102);
nor U5935 (N_5935,N_2801,N_4136);
nand U5936 (N_5936,N_4703,N_4884);
or U5937 (N_5937,N_3784,N_4137);
and U5938 (N_5938,N_2694,N_3474);
nand U5939 (N_5939,N_2976,N_3849);
nor U5940 (N_5940,N_4340,N_3150);
nor U5941 (N_5941,N_4955,N_4856);
and U5942 (N_5942,N_3892,N_3871);
and U5943 (N_5943,N_4024,N_3898);
nand U5944 (N_5944,N_4245,N_3424);
and U5945 (N_5945,N_3360,N_4885);
and U5946 (N_5946,N_4736,N_3431);
nor U5947 (N_5947,N_4945,N_4862);
or U5948 (N_5948,N_4489,N_4409);
nor U5949 (N_5949,N_2659,N_3999);
nor U5950 (N_5950,N_4623,N_4321);
xor U5951 (N_5951,N_4858,N_4296);
xor U5952 (N_5952,N_4376,N_3493);
xor U5953 (N_5953,N_3463,N_2998);
or U5954 (N_5954,N_3677,N_3077);
nand U5955 (N_5955,N_3787,N_4811);
nand U5956 (N_5956,N_4206,N_4290);
nand U5957 (N_5957,N_4313,N_3332);
and U5958 (N_5958,N_4833,N_4500);
xor U5959 (N_5959,N_2570,N_3231);
nor U5960 (N_5960,N_4151,N_4424);
nand U5961 (N_5961,N_4598,N_3457);
or U5962 (N_5962,N_4734,N_3184);
and U5963 (N_5963,N_4637,N_3015);
nand U5964 (N_5964,N_3788,N_2630);
nand U5965 (N_5965,N_2757,N_3447);
or U5966 (N_5966,N_3598,N_4334);
or U5967 (N_5967,N_3768,N_4433);
nand U5968 (N_5968,N_3844,N_2835);
or U5969 (N_5969,N_2619,N_4278);
and U5970 (N_5970,N_3565,N_4324);
or U5971 (N_5971,N_4112,N_3696);
nor U5972 (N_5972,N_3314,N_3339);
xnor U5973 (N_5973,N_3702,N_4735);
and U5974 (N_5974,N_2821,N_2928);
or U5975 (N_5975,N_3957,N_4678);
or U5976 (N_5976,N_2882,N_2683);
xnor U5977 (N_5977,N_2679,N_3853);
nand U5978 (N_5978,N_4714,N_2931);
xnor U5979 (N_5979,N_3726,N_3055);
nor U5980 (N_5980,N_2744,N_4652);
nand U5981 (N_5981,N_4282,N_2573);
nor U5982 (N_5982,N_2997,N_2799);
xor U5983 (N_5983,N_3461,N_4931);
or U5984 (N_5984,N_3147,N_4462);
and U5985 (N_5985,N_3986,N_3678);
and U5986 (N_5986,N_4277,N_4454);
nand U5987 (N_5987,N_3735,N_3769);
nor U5988 (N_5988,N_3599,N_3626);
or U5989 (N_5989,N_4476,N_3045);
nand U5990 (N_5990,N_2726,N_3815);
nand U5991 (N_5991,N_3473,N_4713);
and U5992 (N_5992,N_3331,N_3270);
nand U5993 (N_5993,N_3475,N_4299);
xor U5994 (N_5994,N_3178,N_4463);
and U5995 (N_5995,N_2556,N_4367);
xor U5996 (N_5996,N_4632,N_4646);
or U5997 (N_5997,N_3670,N_4418);
or U5998 (N_5998,N_4571,N_4275);
or U5999 (N_5999,N_4921,N_3028);
and U6000 (N_6000,N_4333,N_2993);
nor U6001 (N_6001,N_4222,N_3722);
xnor U6002 (N_6002,N_4031,N_4446);
or U6003 (N_6003,N_2842,N_4876);
xnor U6004 (N_6004,N_3527,N_3621);
and U6005 (N_6005,N_3371,N_4888);
xnor U6006 (N_6006,N_3961,N_4774);
nand U6007 (N_6007,N_4369,N_4610);
or U6008 (N_6008,N_4912,N_2924);
or U6009 (N_6009,N_3037,N_4232);
and U6010 (N_6010,N_4764,N_3291);
or U6011 (N_6011,N_4453,N_4219);
and U6012 (N_6012,N_4923,N_4128);
or U6013 (N_6013,N_3511,N_4771);
or U6014 (N_6014,N_3649,N_3886);
nor U6015 (N_6015,N_4349,N_4625);
nor U6016 (N_6016,N_2561,N_2771);
or U6017 (N_6017,N_3075,N_3004);
or U6018 (N_6018,N_4330,N_3312);
nor U6019 (N_6019,N_4530,N_3624);
nand U6020 (N_6020,N_4508,N_3458);
nand U6021 (N_6021,N_4930,N_3736);
and U6022 (N_6022,N_4064,N_3682);
xor U6023 (N_6023,N_3550,N_3880);
or U6024 (N_6024,N_3857,N_2865);
nand U6025 (N_6025,N_3233,N_4338);
and U6026 (N_6026,N_4021,N_2725);
nand U6027 (N_6027,N_4153,N_4789);
or U6028 (N_6028,N_2864,N_4986);
or U6029 (N_6029,N_4301,N_2641);
or U6030 (N_6030,N_4991,N_2665);
and U6031 (N_6031,N_4135,N_4223);
and U6032 (N_6032,N_3773,N_4412);
nand U6033 (N_6033,N_2657,N_4806);
nor U6034 (N_6034,N_4760,N_4159);
xnor U6035 (N_6035,N_4405,N_4403);
and U6036 (N_6036,N_2727,N_3109);
and U6037 (N_6037,N_3630,N_3409);
and U6038 (N_6038,N_3967,N_3226);
nand U6039 (N_6039,N_3798,N_4216);
or U6040 (N_6040,N_2975,N_3411);
and U6041 (N_6041,N_4994,N_3165);
nand U6042 (N_6042,N_4294,N_3686);
nand U6043 (N_6043,N_4948,N_3666);
and U6044 (N_6044,N_4394,N_3415);
nor U6045 (N_6045,N_3023,N_4091);
and U6046 (N_6046,N_3159,N_4157);
nand U6047 (N_6047,N_3842,N_3116);
and U6048 (N_6048,N_2565,N_4910);
or U6049 (N_6049,N_3132,N_3791);
or U6050 (N_6050,N_3297,N_3660);
and U6051 (N_6051,N_4016,N_4609);
or U6052 (N_6052,N_2701,N_3750);
nand U6053 (N_6053,N_4495,N_3287);
nand U6054 (N_6054,N_4094,N_2881);
and U6055 (N_6055,N_3309,N_3990);
xnor U6056 (N_6056,N_4093,N_3616);
and U6057 (N_6057,N_4675,N_3703);
and U6058 (N_6058,N_4602,N_3952);
nand U6059 (N_6059,N_2804,N_3124);
nor U6060 (N_6060,N_4622,N_4484);
xnor U6061 (N_6061,N_3710,N_4728);
nor U6062 (N_6062,N_3929,N_4733);
nand U6063 (N_6063,N_3936,N_3412);
xnor U6064 (N_6064,N_3034,N_3919);
and U6065 (N_6065,N_3388,N_2553);
xnor U6066 (N_6066,N_2824,N_4507);
or U6067 (N_6067,N_3977,N_3478);
nor U6068 (N_6068,N_3257,N_2632);
or U6069 (N_6069,N_2623,N_2601);
xor U6070 (N_6070,N_3549,N_2851);
nand U6071 (N_6071,N_4726,N_4606);
nand U6072 (N_6072,N_3714,N_2670);
and U6073 (N_6073,N_4218,N_3158);
nand U6074 (N_6074,N_2633,N_2692);
nor U6075 (N_6075,N_3068,N_3019);
nor U6076 (N_6076,N_3679,N_4315);
nor U6077 (N_6077,N_3940,N_2677);
nor U6078 (N_6078,N_4844,N_2515);
xnor U6079 (N_6079,N_2584,N_4869);
nand U6080 (N_6080,N_2921,N_3046);
nor U6081 (N_6081,N_3531,N_4810);
nand U6082 (N_6082,N_4950,N_3996);
or U6083 (N_6083,N_4191,N_3375);
nand U6084 (N_6084,N_3541,N_2803);
xnor U6085 (N_6085,N_4013,N_3533);
nand U6086 (N_6086,N_4587,N_4524);
nor U6087 (N_6087,N_2917,N_2672);
nand U6088 (N_6088,N_2905,N_3381);
nor U6089 (N_6089,N_3191,N_2513);
or U6090 (N_6090,N_3262,N_2638);
or U6091 (N_6091,N_4843,N_2635);
or U6092 (N_6092,N_2827,N_3829);
or U6093 (N_6093,N_4579,N_3512);
or U6094 (N_6094,N_4033,N_2986);
or U6095 (N_6095,N_3181,N_2957);
xnor U6096 (N_6096,N_3337,N_2761);
and U6097 (N_6097,N_3126,N_2614);
nor U6098 (N_6098,N_3108,N_3211);
or U6099 (N_6099,N_2684,N_4375);
and U6100 (N_6100,N_4857,N_3142);
and U6101 (N_6101,N_4081,N_4546);
or U6102 (N_6102,N_4949,N_3924);
nor U6103 (N_6103,N_3707,N_2991);
nand U6104 (N_6104,N_3830,N_4660);
or U6105 (N_6105,N_4807,N_3466);
or U6106 (N_6106,N_3721,N_4967);
nor U6107 (N_6107,N_4284,N_4777);
nand U6108 (N_6108,N_3432,N_4522);
nor U6109 (N_6109,N_4152,N_3745);
or U6110 (N_6110,N_2545,N_2902);
nand U6111 (N_6111,N_3947,N_3428);
and U6112 (N_6112,N_4242,N_4922);
nor U6113 (N_6113,N_2784,N_3575);
or U6114 (N_6114,N_3148,N_4552);
nand U6115 (N_6115,N_4793,N_4687);
or U6116 (N_6116,N_2776,N_3404);
nand U6117 (N_6117,N_3617,N_2981);
nor U6118 (N_6118,N_2829,N_2870);
nor U6119 (N_6119,N_4831,N_3693);
and U6120 (N_6120,N_4920,N_3396);
or U6121 (N_6121,N_3510,N_2980);
or U6122 (N_6122,N_4788,N_3087);
nor U6123 (N_6123,N_4903,N_4142);
and U6124 (N_6124,N_4808,N_2536);
nor U6125 (N_6125,N_4911,N_2786);
or U6126 (N_6126,N_3823,N_4362);
or U6127 (N_6127,N_4821,N_4256);
nand U6128 (N_6128,N_2559,N_4215);
nand U6129 (N_6129,N_3920,N_4397);
nor U6130 (N_6130,N_3179,N_3865);
or U6131 (N_6131,N_3904,N_4002);
or U6132 (N_6132,N_3476,N_4150);
or U6133 (N_6133,N_2886,N_4551);
nor U6134 (N_6134,N_3441,N_4573);
and U6135 (N_6135,N_2795,N_4022);
nor U6136 (N_6136,N_4276,N_3005);
nor U6137 (N_6137,N_4563,N_3657);
or U6138 (N_6138,N_3734,N_2904);
nand U6139 (N_6139,N_4263,N_3040);
nand U6140 (N_6140,N_2714,N_2987);
xnor U6141 (N_6141,N_2629,N_4969);
nand U6142 (N_6142,N_4268,N_2578);
xnor U6143 (N_6143,N_4480,N_4752);
or U6144 (N_6144,N_3468,N_2746);
xnor U6145 (N_6145,N_3328,N_2522);
nor U6146 (N_6146,N_4915,N_4636);
nand U6147 (N_6147,N_4899,N_4834);
nor U6148 (N_6148,N_4399,N_3379);
or U6149 (N_6149,N_2797,N_4518);
nand U6150 (N_6150,N_3243,N_3713);
nor U6151 (N_6151,N_3172,N_3096);
nand U6152 (N_6152,N_3102,N_3640);
nor U6153 (N_6153,N_2858,N_4414);
nand U6154 (N_6154,N_4261,N_3030);
nor U6155 (N_6155,N_4671,N_4413);
nor U6156 (N_6156,N_3636,N_4144);
and U6157 (N_6157,N_3820,N_2763);
or U6158 (N_6158,N_2805,N_4932);
nand U6159 (N_6159,N_3708,N_3644);
and U6160 (N_6160,N_4004,N_2968);
and U6161 (N_6161,N_4624,N_3294);
or U6162 (N_6162,N_3256,N_2883);
or U6163 (N_6163,N_4545,N_2655);
or U6164 (N_6164,N_4628,N_4644);
xnor U6165 (N_6165,N_4028,N_4794);
nor U6166 (N_6166,N_4716,N_4181);
nand U6167 (N_6167,N_3577,N_3094);
xnor U6168 (N_6168,N_4420,N_4537);
or U6169 (N_6169,N_4099,N_3580);
nor U6170 (N_6170,N_3778,N_2564);
and U6171 (N_6171,N_4030,N_3009);
or U6172 (N_6172,N_2833,N_2849);
and U6173 (N_6173,N_4740,N_2942);
or U6174 (N_6174,N_3748,N_3263);
or U6175 (N_6175,N_2738,N_3021);
nand U6176 (N_6176,N_3044,N_3101);
and U6177 (N_6177,N_4802,N_3514);
or U6178 (N_6178,N_2693,N_3362);
and U6179 (N_6179,N_2859,N_4364);
or U6180 (N_6180,N_3135,N_2722);
and U6181 (N_6181,N_3962,N_3923);
and U6182 (N_6182,N_4018,N_4629);
nor U6183 (N_6183,N_4890,N_2920);
and U6184 (N_6184,N_3350,N_3043);
or U6185 (N_6185,N_3218,N_2577);
nor U6186 (N_6186,N_4188,N_4693);
nor U6187 (N_6187,N_4585,N_4332);
nor U6188 (N_6188,N_4647,N_4528);
and U6189 (N_6189,N_3656,N_3664);
or U6190 (N_6190,N_3489,N_3370);
and U6191 (N_6191,N_2911,N_4442);
or U6192 (N_6192,N_3163,N_4896);
nor U6193 (N_6193,N_2708,N_2841);
xnor U6194 (N_6194,N_4900,N_3242);
and U6195 (N_6195,N_3210,N_4989);
or U6196 (N_6196,N_4096,N_3250);
nor U6197 (N_6197,N_2890,N_4088);
and U6198 (N_6198,N_4655,N_3275);
nand U6199 (N_6199,N_3252,N_2876);
nand U6200 (N_6200,N_4356,N_4988);
nor U6201 (N_6201,N_3192,N_4286);
nor U6202 (N_6202,N_3020,N_3133);
or U6203 (N_6203,N_2778,N_4615);
nor U6204 (N_6204,N_4634,N_2825);
and U6205 (N_6205,N_3795,N_3264);
or U6206 (N_6206,N_4179,N_4431);
and U6207 (N_6207,N_3856,N_3744);
nand U6208 (N_6208,N_2669,N_3955);
and U6209 (N_6209,N_2844,N_2879);
or U6210 (N_6210,N_3038,N_3425);
or U6211 (N_6211,N_3760,N_3410);
nor U6212 (N_6212,N_3353,N_3897);
and U6213 (N_6213,N_4472,N_3338);
or U6214 (N_6214,N_3738,N_3979);
nand U6215 (N_6215,N_4614,N_4745);
nor U6216 (N_6216,N_4916,N_4283);
nand U6217 (N_6217,N_3992,N_4658);
or U6218 (N_6218,N_4103,N_3716);
and U6219 (N_6219,N_4052,N_4574);
or U6220 (N_6220,N_3062,N_4928);
nand U6221 (N_6221,N_4851,N_4175);
or U6222 (N_6222,N_4699,N_4062);
nand U6223 (N_6223,N_2582,N_4272);
and U6224 (N_6224,N_2622,N_4569);
nor U6225 (N_6225,N_4650,N_4458);
nand U6226 (N_6226,N_2721,N_4768);
nor U6227 (N_6227,N_2704,N_2660);
and U6228 (N_6228,N_3633,N_4273);
and U6229 (N_6229,N_4554,N_4824);
nand U6230 (N_6230,N_4260,N_3645);
and U6231 (N_6231,N_3944,N_3834);
and U6232 (N_6232,N_4133,N_3282);
or U6233 (N_6233,N_2934,N_2639);
or U6234 (N_6234,N_3724,N_3814);
xor U6235 (N_6235,N_3597,N_4439);
and U6236 (N_6236,N_4410,N_4908);
nand U6237 (N_6237,N_2800,N_3581);
and U6238 (N_6238,N_3027,N_2579);
and U6239 (N_6239,N_4827,N_3690);
and U6240 (N_6240,N_3240,N_3480);
nor U6241 (N_6241,N_3862,N_4532);
and U6242 (N_6242,N_4711,N_2878);
nor U6243 (N_6243,N_2705,N_4158);
and U6244 (N_6244,N_2636,N_2710);
nor U6245 (N_6245,N_2802,N_4861);
and U6246 (N_6246,N_2808,N_4240);
or U6247 (N_6247,N_2718,N_3000);
or U6248 (N_6248,N_3950,N_3840);
and U6249 (N_6249,N_4767,N_2502);
nor U6250 (N_6250,N_4482,N_3513);
nand U6251 (N_6251,N_3686,N_3223);
and U6252 (N_6252,N_4074,N_2906);
or U6253 (N_6253,N_4161,N_2641);
xor U6254 (N_6254,N_4228,N_4899);
or U6255 (N_6255,N_3793,N_2881);
or U6256 (N_6256,N_3417,N_2578);
or U6257 (N_6257,N_4481,N_4364);
and U6258 (N_6258,N_3963,N_3354);
xnor U6259 (N_6259,N_3163,N_3496);
xor U6260 (N_6260,N_2962,N_3832);
nor U6261 (N_6261,N_3408,N_3067);
or U6262 (N_6262,N_3963,N_2695);
nor U6263 (N_6263,N_2840,N_4558);
and U6264 (N_6264,N_3689,N_4835);
and U6265 (N_6265,N_2972,N_3614);
nor U6266 (N_6266,N_2891,N_4340);
and U6267 (N_6267,N_3037,N_3272);
nand U6268 (N_6268,N_3687,N_3175);
and U6269 (N_6269,N_4904,N_3742);
nor U6270 (N_6270,N_3502,N_4342);
xor U6271 (N_6271,N_3340,N_2709);
or U6272 (N_6272,N_2943,N_4432);
or U6273 (N_6273,N_4989,N_3385);
xor U6274 (N_6274,N_3390,N_4763);
nor U6275 (N_6275,N_4556,N_2644);
or U6276 (N_6276,N_2895,N_4245);
and U6277 (N_6277,N_3228,N_3898);
or U6278 (N_6278,N_3205,N_3617);
nor U6279 (N_6279,N_4502,N_4818);
and U6280 (N_6280,N_3664,N_4577);
nor U6281 (N_6281,N_2846,N_3058);
nand U6282 (N_6282,N_3752,N_3953);
xor U6283 (N_6283,N_4675,N_4699);
nor U6284 (N_6284,N_4315,N_4691);
or U6285 (N_6285,N_3375,N_4823);
nor U6286 (N_6286,N_2956,N_3212);
and U6287 (N_6287,N_4403,N_3677);
and U6288 (N_6288,N_4317,N_3044);
nor U6289 (N_6289,N_3914,N_2700);
and U6290 (N_6290,N_3966,N_3523);
or U6291 (N_6291,N_3358,N_3305);
and U6292 (N_6292,N_4784,N_4197);
and U6293 (N_6293,N_3374,N_4651);
nand U6294 (N_6294,N_3462,N_4454);
nand U6295 (N_6295,N_2728,N_3157);
xor U6296 (N_6296,N_4403,N_4633);
or U6297 (N_6297,N_3852,N_3524);
or U6298 (N_6298,N_4691,N_4283);
or U6299 (N_6299,N_3769,N_3441);
xnor U6300 (N_6300,N_3378,N_2730);
nand U6301 (N_6301,N_3859,N_2679);
or U6302 (N_6302,N_4235,N_2572);
nand U6303 (N_6303,N_3988,N_3168);
nand U6304 (N_6304,N_4982,N_3660);
and U6305 (N_6305,N_4588,N_2514);
or U6306 (N_6306,N_4801,N_3036);
nor U6307 (N_6307,N_3961,N_4698);
nand U6308 (N_6308,N_3950,N_4653);
nand U6309 (N_6309,N_2866,N_4272);
or U6310 (N_6310,N_4334,N_4462);
and U6311 (N_6311,N_3804,N_4756);
nand U6312 (N_6312,N_3272,N_4017);
or U6313 (N_6313,N_4835,N_3011);
and U6314 (N_6314,N_3570,N_3635);
or U6315 (N_6315,N_3817,N_3069);
or U6316 (N_6316,N_4245,N_3219);
or U6317 (N_6317,N_4568,N_3869);
and U6318 (N_6318,N_3434,N_3549);
and U6319 (N_6319,N_4624,N_2596);
nor U6320 (N_6320,N_4409,N_3642);
or U6321 (N_6321,N_3373,N_3859);
nand U6322 (N_6322,N_3971,N_4387);
and U6323 (N_6323,N_2907,N_4023);
nand U6324 (N_6324,N_4192,N_4226);
or U6325 (N_6325,N_4874,N_3626);
nor U6326 (N_6326,N_2950,N_4712);
or U6327 (N_6327,N_4281,N_3671);
or U6328 (N_6328,N_4044,N_3606);
or U6329 (N_6329,N_3115,N_3578);
or U6330 (N_6330,N_4010,N_4234);
nor U6331 (N_6331,N_4927,N_3105);
nand U6332 (N_6332,N_2699,N_3110);
nand U6333 (N_6333,N_3933,N_4824);
or U6334 (N_6334,N_2989,N_3868);
or U6335 (N_6335,N_4863,N_4788);
nor U6336 (N_6336,N_4057,N_3938);
xor U6337 (N_6337,N_2942,N_4996);
nand U6338 (N_6338,N_4738,N_3095);
and U6339 (N_6339,N_3677,N_2812);
or U6340 (N_6340,N_3538,N_2756);
nor U6341 (N_6341,N_4863,N_2904);
or U6342 (N_6342,N_4792,N_3995);
and U6343 (N_6343,N_4207,N_4422);
nand U6344 (N_6344,N_4447,N_4760);
or U6345 (N_6345,N_2613,N_2700);
or U6346 (N_6346,N_4759,N_3268);
xor U6347 (N_6347,N_2575,N_2973);
and U6348 (N_6348,N_3848,N_4612);
nand U6349 (N_6349,N_4267,N_4340);
and U6350 (N_6350,N_4662,N_3119);
xor U6351 (N_6351,N_4690,N_4738);
nand U6352 (N_6352,N_3773,N_2584);
and U6353 (N_6353,N_4066,N_2677);
nor U6354 (N_6354,N_4774,N_3652);
nor U6355 (N_6355,N_4515,N_4957);
nand U6356 (N_6356,N_4605,N_4121);
and U6357 (N_6357,N_3569,N_2915);
nand U6358 (N_6358,N_4314,N_2587);
nor U6359 (N_6359,N_2721,N_2885);
and U6360 (N_6360,N_4227,N_2505);
and U6361 (N_6361,N_3348,N_4914);
nand U6362 (N_6362,N_3346,N_4226);
and U6363 (N_6363,N_4431,N_4358);
and U6364 (N_6364,N_2825,N_4066);
and U6365 (N_6365,N_4004,N_3822);
or U6366 (N_6366,N_2527,N_4265);
xor U6367 (N_6367,N_2871,N_4573);
nor U6368 (N_6368,N_3197,N_4833);
nand U6369 (N_6369,N_3165,N_4234);
or U6370 (N_6370,N_3796,N_4485);
nand U6371 (N_6371,N_4084,N_2616);
xor U6372 (N_6372,N_4091,N_3155);
nand U6373 (N_6373,N_2924,N_4987);
nand U6374 (N_6374,N_4074,N_2787);
and U6375 (N_6375,N_4009,N_4117);
and U6376 (N_6376,N_3385,N_3482);
nand U6377 (N_6377,N_4711,N_4623);
nor U6378 (N_6378,N_2896,N_4475);
xor U6379 (N_6379,N_4596,N_3688);
or U6380 (N_6380,N_2756,N_4031);
and U6381 (N_6381,N_3766,N_4041);
and U6382 (N_6382,N_4888,N_4481);
nor U6383 (N_6383,N_3724,N_2792);
or U6384 (N_6384,N_4329,N_4074);
and U6385 (N_6385,N_4077,N_3274);
or U6386 (N_6386,N_2970,N_3402);
or U6387 (N_6387,N_2534,N_4326);
nor U6388 (N_6388,N_4877,N_3462);
or U6389 (N_6389,N_3751,N_3896);
and U6390 (N_6390,N_2869,N_4298);
or U6391 (N_6391,N_4651,N_2528);
nor U6392 (N_6392,N_4467,N_3710);
nor U6393 (N_6393,N_4267,N_4302);
nand U6394 (N_6394,N_2553,N_3579);
nand U6395 (N_6395,N_3440,N_4397);
nand U6396 (N_6396,N_3806,N_3213);
or U6397 (N_6397,N_4396,N_4774);
nor U6398 (N_6398,N_4389,N_4083);
nor U6399 (N_6399,N_4890,N_2855);
nand U6400 (N_6400,N_4837,N_4126);
nor U6401 (N_6401,N_4835,N_4701);
or U6402 (N_6402,N_2790,N_3262);
xnor U6403 (N_6403,N_3716,N_4439);
nand U6404 (N_6404,N_4894,N_3694);
xnor U6405 (N_6405,N_3930,N_2618);
and U6406 (N_6406,N_4597,N_4623);
and U6407 (N_6407,N_4384,N_3465);
nor U6408 (N_6408,N_4452,N_3878);
xnor U6409 (N_6409,N_4206,N_3934);
nand U6410 (N_6410,N_3136,N_4595);
nor U6411 (N_6411,N_3934,N_4002);
or U6412 (N_6412,N_4712,N_3977);
or U6413 (N_6413,N_2802,N_3396);
and U6414 (N_6414,N_4660,N_3434);
nand U6415 (N_6415,N_3802,N_4743);
nor U6416 (N_6416,N_4929,N_4634);
and U6417 (N_6417,N_4100,N_4650);
or U6418 (N_6418,N_4479,N_4694);
xor U6419 (N_6419,N_3998,N_4214);
or U6420 (N_6420,N_3463,N_2727);
and U6421 (N_6421,N_3670,N_3890);
or U6422 (N_6422,N_3248,N_4745);
or U6423 (N_6423,N_2560,N_3024);
xnor U6424 (N_6424,N_3993,N_4887);
nand U6425 (N_6425,N_3443,N_3556);
and U6426 (N_6426,N_2630,N_4540);
nor U6427 (N_6427,N_4403,N_2610);
and U6428 (N_6428,N_4719,N_4478);
nand U6429 (N_6429,N_2748,N_2611);
nor U6430 (N_6430,N_4525,N_4917);
or U6431 (N_6431,N_4746,N_3625);
or U6432 (N_6432,N_4217,N_3602);
or U6433 (N_6433,N_3057,N_4317);
nor U6434 (N_6434,N_3086,N_2928);
nor U6435 (N_6435,N_2921,N_4456);
nor U6436 (N_6436,N_4124,N_2853);
or U6437 (N_6437,N_4786,N_4020);
nor U6438 (N_6438,N_4877,N_3771);
nand U6439 (N_6439,N_2904,N_3792);
or U6440 (N_6440,N_4030,N_3776);
or U6441 (N_6441,N_3758,N_3301);
or U6442 (N_6442,N_2613,N_2546);
nand U6443 (N_6443,N_3738,N_4798);
and U6444 (N_6444,N_3201,N_4233);
nand U6445 (N_6445,N_3602,N_4963);
or U6446 (N_6446,N_3217,N_3918);
nand U6447 (N_6447,N_4519,N_3665);
or U6448 (N_6448,N_3548,N_4426);
nand U6449 (N_6449,N_3761,N_3763);
and U6450 (N_6450,N_2603,N_4751);
or U6451 (N_6451,N_3433,N_4750);
nor U6452 (N_6452,N_4364,N_4788);
and U6453 (N_6453,N_4575,N_2934);
or U6454 (N_6454,N_4942,N_2960);
nor U6455 (N_6455,N_4302,N_2837);
or U6456 (N_6456,N_2713,N_3014);
or U6457 (N_6457,N_3542,N_2676);
nand U6458 (N_6458,N_4096,N_3252);
and U6459 (N_6459,N_3647,N_4988);
nand U6460 (N_6460,N_3477,N_4044);
nand U6461 (N_6461,N_4109,N_3812);
and U6462 (N_6462,N_3141,N_2507);
nand U6463 (N_6463,N_3576,N_4787);
xor U6464 (N_6464,N_2732,N_3221);
nor U6465 (N_6465,N_2633,N_3865);
nand U6466 (N_6466,N_2948,N_2521);
xor U6467 (N_6467,N_2660,N_2591);
nand U6468 (N_6468,N_3023,N_4113);
nor U6469 (N_6469,N_4145,N_4342);
nor U6470 (N_6470,N_3887,N_4695);
nand U6471 (N_6471,N_3316,N_3659);
or U6472 (N_6472,N_4427,N_4056);
nand U6473 (N_6473,N_3720,N_3187);
and U6474 (N_6474,N_3794,N_3944);
nand U6475 (N_6475,N_3390,N_2989);
nor U6476 (N_6476,N_3379,N_3258);
nand U6477 (N_6477,N_4366,N_3116);
nor U6478 (N_6478,N_4840,N_2594);
or U6479 (N_6479,N_4839,N_4545);
and U6480 (N_6480,N_3288,N_2759);
nand U6481 (N_6481,N_4157,N_4634);
and U6482 (N_6482,N_3001,N_4594);
and U6483 (N_6483,N_4676,N_3573);
nor U6484 (N_6484,N_3296,N_3500);
nand U6485 (N_6485,N_3263,N_3704);
nor U6486 (N_6486,N_4125,N_3565);
nor U6487 (N_6487,N_4613,N_3746);
nor U6488 (N_6488,N_2603,N_4163);
and U6489 (N_6489,N_4298,N_4605);
nor U6490 (N_6490,N_3783,N_4085);
nor U6491 (N_6491,N_2563,N_3497);
nor U6492 (N_6492,N_3028,N_3943);
or U6493 (N_6493,N_4036,N_4322);
and U6494 (N_6494,N_4022,N_3882);
nand U6495 (N_6495,N_2665,N_2500);
and U6496 (N_6496,N_4683,N_3641);
and U6497 (N_6497,N_4276,N_2727);
or U6498 (N_6498,N_3756,N_3519);
nor U6499 (N_6499,N_4612,N_4046);
or U6500 (N_6500,N_3795,N_3583);
nor U6501 (N_6501,N_2554,N_2989);
xnor U6502 (N_6502,N_4808,N_3629);
nor U6503 (N_6503,N_2838,N_2684);
or U6504 (N_6504,N_2940,N_4566);
or U6505 (N_6505,N_2795,N_3699);
and U6506 (N_6506,N_3327,N_2824);
and U6507 (N_6507,N_3320,N_4162);
or U6508 (N_6508,N_4680,N_4120);
and U6509 (N_6509,N_3320,N_2812);
nor U6510 (N_6510,N_3555,N_3963);
and U6511 (N_6511,N_3140,N_2540);
nor U6512 (N_6512,N_3275,N_4993);
or U6513 (N_6513,N_4300,N_4092);
nor U6514 (N_6514,N_4344,N_2655);
and U6515 (N_6515,N_3845,N_4278);
nand U6516 (N_6516,N_4684,N_2929);
or U6517 (N_6517,N_2771,N_4420);
and U6518 (N_6518,N_3391,N_4153);
nand U6519 (N_6519,N_3398,N_4841);
and U6520 (N_6520,N_3678,N_4923);
nand U6521 (N_6521,N_4646,N_4591);
or U6522 (N_6522,N_3254,N_3821);
and U6523 (N_6523,N_2705,N_2549);
xor U6524 (N_6524,N_4898,N_4800);
and U6525 (N_6525,N_2940,N_4415);
and U6526 (N_6526,N_3035,N_2689);
nor U6527 (N_6527,N_3988,N_3050);
or U6528 (N_6528,N_2904,N_2777);
nor U6529 (N_6529,N_3342,N_3398);
and U6530 (N_6530,N_3316,N_2639);
nor U6531 (N_6531,N_4609,N_3168);
xor U6532 (N_6532,N_4131,N_4511);
nor U6533 (N_6533,N_4091,N_2928);
nor U6534 (N_6534,N_3568,N_4810);
or U6535 (N_6535,N_4299,N_3333);
nor U6536 (N_6536,N_3064,N_4819);
nand U6537 (N_6537,N_3713,N_3278);
or U6538 (N_6538,N_2676,N_3024);
nand U6539 (N_6539,N_2608,N_3009);
nor U6540 (N_6540,N_2580,N_3828);
nor U6541 (N_6541,N_3939,N_3080);
and U6542 (N_6542,N_2539,N_4905);
or U6543 (N_6543,N_4827,N_4289);
nor U6544 (N_6544,N_2684,N_2987);
nand U6545 (N_6545,N_3812,N_4180);
or U6546 (N_6546,N_2509,N_2776);
and U6547 (N_6547,N_4976,N_4110);
nor U6548 (N_6548,N_4302,N_2754);
or U6549 (N_6549,N_2533,N_4440);
and U6550 (N_6550,N_4816,N_3922);
nand U6551 (N_6551,N_3799,N_4422);
nor U6552 (N_6552,N_2964,N_4924);
or U6553 (N_6553,N_4129,N_3682);
nand U6554 (N_6554,N_3448,N_3547);
nor U6555 (N_6555,N_3931,N_3762);
nor U6556 (N_6556,N_4844,N_3254);
nand U6557 (N_6557,N_2547,N_3931);
and U6558 (N_6558,N_2963,N_4457);
nand U6559 (N_6559,N_2808,N_2846);
or U6560 (N_6560,N_2975,N_4721);
nor U6561 (N_6561,N_4721,N_2776);
nor U6562 (N_6562,N_3245,N_2508);
nand U6563 (N_6563,N_2958,N_4693);
or U6564 (N_6564,N_4374,N_4549);
or U6565 (N_6565,N_3578,N_3095);
and U6566 (N_6566,N_3017,N_4096);
nor U6567 (N_6567,N_3696,N_4111);
or U6568 (N_6568,N_4576,N_2791);
or U6569 (N_6569,N_4772,N_3746);
nand U6570 (N_6570,N_3657,N_4481);
or U6571 (N_6571,N_4003,N_3302);
or U6572 (N_6572,N_3118,N_4345);
nand U6573 (N_6573,N_2520,N_3016);
or U6574 (N_6574,N_2953,N_3390);
or U6575 (N_6575,N_4939,N_3878);
or U6576 (N_6576,N_2896,N_3529);
nor U6577 (N_6577,N_2939,N_2657);
nor U6578 (N_6578,N_3340,N_2514);
xnor U6579 (N_6579,N_2751,N_4414);
nand U6580 (N_6580,N_2508,N_4551);
nand U6581 (N_6581,N_2947,N_3921);
and U6582 (N_6582,N_2987,N_4753);
nor U6583 (N_6583,N_3937,N_3900);
nor U6584 (N_6584,N_4551,N_4000);
and U6585 (N_6585,N_3606,N_4415);
nor U6586 (N_6586,N_4210,N_4445);
nand U6587 (N_6587,N_4456,N_4696);
and U6588 (N_6588,N_3859,N_3830);
and U6589 (N_6589,N_2722,N_2661);
nor U6590 (N_6590,N_4653,N_3267);
or U6591 (N_6591,N_3623,N_4148);
and U6592 (N_6592,N_2888,N_4703);
nand U6593 (N_6593,N_3649,N_3327);
or U6594 (N_6594,N_3719,N_4161);
and U6595 (N_6595,N_4529,N_4447);
and U6596 (N_6596,N_4571,N_4858);
nand U6597 (N_6597,N_3811,N_3949);
nor U6598 (N_6598,N_4320,N_3286);
and U6599 (N_6599,N_4184,N_3945);
nor U6600 (N_6600,N_4108,N_4198);
nand U6601 (N_6601,N_4546,N_4545);
or U6602 (N_6602,N_4597,N_4493);
or U6603 (N_6603,N_2937,N_2990);
or U6604 (N_6604,N_3247,N_2683);
xnor U6605 (N_6605,N_2838,N_4075);
and U6606 (N_6606,N_3881,N_4827);
xor U6607 (N_6607,N_3436,N_2677);
nor U6608 (N_6608,N_4626,N_4076);
xnor U6609 (N_6609,N_4346,N_3208);
or U6610 (N_6610,N_3087,N_3878);
nand U6611 (N_6611,N_3295,N_3690);
or U6612 (N_6612,N_2937,N_3506);
or U6613 (N_6613,N_2792,N_3783);
and U6614 (N_6614,N_3808,N_2676);
and U6615 (N_6615,N_3073,N_4925);
or U6616 (N_6616,N_2901,N_4146);
nor U6617 (N_6617,N_4595,N_3165);
xnor U6618 (N_6618,N_4866,N_3713);
nor U6619 (N_6619,N_3833,N_3782);
xnor U6620 (N_6620,N_2571,N_3755);
nor U6621 (N_6621,N_2733,N_2698);
nor U6622 (N_6622,N_2681,N_2850);
and U6623 (N_6623,N_4739,N_3221);
nor U6624 (N_6624,N_3987,N_3035);
and U6625 (N_6625,N_2579,N_3209);
xnor U6626 (N_6626,N_3085,N_3897);
nor U6627 (N_6627,N_4427,N_3337);
nand U6628 (N_6628,N_3838,N_4482);
or U6629 (N_6629,N_2656,N_4798);
xnor U6630 (N_6630,N_4865,N_4426);
and U6631 (N_6631,N_2799,N_2594);
or U6632 (N_6632,N_2587,N_3169);
and U6633 (N_6633,N_2825,N_3904);
and U6634 (N_6634,N_3126,N_4137);
nor U6635 (N_6635,N_3921,N_4185);
nor U6636 (N_6636,N_3936,N_3147);
and U6637 (N_6637,N_2627,N_3060);
xor U6638 (N_6638,N_3992,N_2756);
and U6639 (N_6639,N_4899,N_3289);
nor U6640 (N_6640,N_3466,N_4023);
nand U6641 (N_6641,N_3511,N_2795);
and U6642 (N_6642,N_4467,N_4160);
nand U6643 (N_6643,N_4144,N_4368);
and U6644 (N_6644,N_4019,N_2726);
nor U6645 (N_6645,N_4568,N_3364);
xnor U6646 (N_6646,N_4163,N_3468);
and U6647 (N_6647,N_2907,N_3062);
nand U6648 (N_6648,N_3406,N_4236);
nor U6649 (N_6649,N_3669,N_3330);
or U6650 (N_6650,N_3010,N_4140);
or U6651 (N_6651,N_4255,N_4061);
nor U6652 (N_6652,N_4350,N_3678);
nor U6653 (N_6653,N_2841,N_3001);
xor U6654 (N_6654,N_3478,N_4838);
nor U6655 (N_6655,N_2686,N_4309);
nor U6656 (N_6656,N_3506,N_3863);
nor U6657 (N_6657,N_3108,N_3096);
nor U6658 (N_6658,N_2643,N_3699);
and U6659 (N_6659,N_3173,N_2710);
nor U6660 (N_6660,N_4951,N_4691);
and U6661 (N_6661,N_4186,N_4172);
nor U6662 (N_6662,N_4717,N_4199);
nor U6663 (N_6663,N_2591,N_4196);
nand U6664 (N_6664,N_4340,N_4301);
nor U6665 (N_6665,N_4717,N_4027);
and U6666 (N_6666,N_4798,N_4300);
nand U6667 (N_6667,N_4107,N_3609);
and U6668 (N_6668,N_3342,N_3141);
and U6669 (N_6669,N_3788,N_3869);
and U6670 (N_6670,N_4883,N_4506);
or U6671 (N_6671,N_2755,N_4578);
and U6672 (N_6672,N_2611,N_4691);
and U6673 (N_6673,N_2949,N_3799);
and U6674 (N_6674,N_4480,N_3744);
and U6675 (N_6675,N_2972,N_2910);
nor U6676 (N_6676,N_2742,N_3755);
nor U6677 (N_6677,N_3578,N_4745);
or U6678 (N_6678,N_4735,N_4114);
nor U6679 (N_6679,N_4388,N_4681);
xor U6680 (N_6680,N_3044,N_3321);
or U6681 (N_6681,N_2678,N_3839);
xor U6682 (N_6682,N_4363,N_2909);
nor U6683 (N_6683,N_3080,N_3246);
xor U6684 (N_6684,N_4907,N_2715);
nor U6685 (N_6685,N_4768,N_3978);
xnor U6686 (N_6686,N_4366,N_3886);
xor U6687 (N_6687,N_4468,N_3417);
xor U6688 (N_6688,N_3581,N_4975);
nor U6689 (N_6689,N_2964,N_4775);
xnor U6690 (N_6690,N_4738,N_4579);
nor U6691 (N_6691,N_2807,N_4773);
or U6692 (N_6692,N_2613,N_4582);
nand U6693 (N_6693,N_2735,N_3021);
nand U6694 (N_6694,N_3811,N_2735);
nand U6695 (N_6695,N_4945,N_3883);
nand U6696 (N_6696,N_4413,N_3412);
nor U6697 (N_6697,N_4851,N_2900);
nor U6698 (N_6698,N_4537,N_2630);
or U6699 (N_6699,N_2635,N_2801);
nor U6700 (N_6700,N_2904,N_3882);
nor U6701 (N_6701,N_4936,N_4989);
nand U6702 (N_6702,N_3054,N_4111);
nand U6703 (N_6703,N_4121,N_4541);
xnor U6704 (N_6704,N_4131,N_2889);
nor U6705 (N_6705,N_3645,N_3588);
xnor U6706 (N_6706,N_3471,N_4062);
and U6707 (N_6707,N_4764,N_4421);
nor U6708 (N_6708,N_3776,N_3060);
nand U6709 (N_6709,N_4843,N_4093);
or U6710 (N_6710,N_4846,N_4466);
or U6711 (N_6711,N_3594,N_3742);
nand U6712 (N_6712,N_4683,N_3395);
nand U6713 (N_6713,N_3797,N_4378);
or U6714 (N_6714,N_2933,N_4485);
nor U6715 (N_6715,N_4805,N_3765);
and U6716 (N_6716,N_3231,N_2974);
nor U6717 (N_6717,N_2873,N_3657);
or U6718 (N_6718,N_3551,N_3729);
nand U6719 (N_6719,N_2726,N_4403);
or U6720 (N_6720,N_4050,N_3793);
and U6721 (N_6721,N_3956,N_3321);
nand U6722 (N_6722,N_3717,N_3402);
and U6723 (N_6723,N_2751,N_3348);
or U6724 (N_6724,N_3649,N_4992);
nand U6725 (N_6725,N_3911,N_3038);
and U6726 (N_6726,N_4623,N_4947);
xnor U6727 (N_6727,N_2723,N_3795);
nor U6728 (N_6728,N_4591,N_3678);
and U6729 (N_6729,N_3304,N_4484);
nand U6730 (N_6730,N_2578,N_4233);
nor U6731 (N_6731,N_3229,N_2828);
xnor U6732 (N_6732,N_4589,N_4634);
and U6733 (N_6733,N_4153,N_4046);
xnor U6734 (N_6734,N_3246,N_2683);
nor U6735 (N_6735,N_2663,N_4015);
and U6736 (N_6736,N_3241,N_4499);
or U6737 (N_6737,N_4538,N_3078);
xnor U6738 (N_6738,N_3111,N_3714);
and U6739 (N_6739,N_3751,N_3615);
nor U6740 (N_6740,N_3049,N_3087);
and U6741 (N_6741,N_2604,N_4328);
and U6742 (N_6742,N_3508,N_4061);
nand U6743 (N_6743,N_4773,N_3508);
xor U6744 (N_6744,N_3037,N_2794);
or U6745 (N_6745,N_3973,N_2567);
nand U6746 (N_6746,N_4201,N_3193);
and U6747 (N_6747,N_4344,N_4545);
nand U6748 (N_6748,N_3821,N_3433);
nor U6749 (N_6749,N_4153,N_2921);
nand U6750 (N_6750,N_2889,N_3287);
nor U6751 (N_6751,N_3286,N_3360);
and U6752 (N_6752,N_4257,N_3592);
and U6753 (N_6753,N_3590,N_3869);
nand U6754 (N_6754,N_4701,N_3085);
and U6755 (N_6755,N_2842,N_3732);
nor U6756 (N_6756,N_3449,N_4772);
nand U6757 (N_6757,N_3092,N_3094);
nand U6758 (N_6758,N_3230,N_2626);
nand U6759 (N_6759,N_3160,N_2574);
nor U6760 (N_6760,N_3479,N_3629);
nand U6761 (N_6761,N_4279,N_3356);
and U6762 (N_6762,N_4989,N_3817);
and U6763 (N_6763,N_3961,N_2585);
xor U6764 (N_6764,N_3347,N_4427);
xor U6765 (N_6765,N_3694,N_2813);
nor U6766 (N_6766,N_3467,N_3756);
and U6767 (N_6767,N_3979,N_4264);
nor U6768 (N_6768,N_2810,N_2849);
or U6769 (N_6769,N_3616,N_3458);
or U6770 (N_6770,N_3390,N_3996);
nor U6771 (N_6771,N_3660,N_2541);
or U6772 (N_6772,N_3983,N_2947);
or U6773 (N_6773,N_3397,N_3707);
nand U6774 (N_6774,N_3711,N_4285);
nor U6775 (N_6775,N_3080,N_4038);
and U6776 (N_6776,N_4015,N_3957);
nor U6777 (N_6777,N_3140,N_3872);
xnor U6778 (N_6778,N_4001,N_4850);
nand U6779 (N_6779,N_3697,N_4709);
nor U6780 (N_6780,N_3692,N_3073);
nor U6781 (N_6781,N_4699,N_2777);
nand U6782 (N_6782,N_2727,N_3545);
nand U6783 (N_6783,N_2867,N_4475);
nor U6784 (N_6784,N_3328,N_3835);
or U6785 (N_6785,N_3661,N_3421);
nand U6786 (N_6786,N_3926,N_3570);
nor U6787 (N_6787,N_4703,N_4622);
nor U6788 (N_6788,N_2561,N_3709);
or U6789 (N_6789,N_2957,N_4235);
nand U6790 (N_6790,N_3114,N_3981);
nor U6791 (N_6791,N_3365,N_4488);
nor U6792 (N_6792,N_4633,N_4194);
or U6793 (N_6793,N_4804,N_3567);
nand U6794 (N_6794,N_3707,N_3515);
nand U6795 (N_6795,N_3278,N_4441);
and U6796 (N_6796,N_3750,N_3751);
and U6797 (N_6797,N_4429,N_4353);
or U6798 (N_6798,N_2850,N_3307);
nor U6799 (N_6799,N_3899,N_4391);
nor U6800 (N_6800,N_2963,N_3323);
and U6801 (N_6801,N_3177,N_4414);
and U6802 (N_6802,N_4761,N_3512);
or U6803 (N_6803,N_3809,N_3313);
xor U6804 (N_6804,N_2898,N_4576);
nand U6805 (N_6805,N_4454,N_4896);
nor U6806 (N_6806,N_4400,N_4064);
nand U6807 (N_6807,N_4224,N_3906);
xnor U6808 (N_6808,N_4393,N_4936);
and U6809 (N_6809,N_3109,N_4088);
or U6810 (N_6810,N_3999,N_4293);
nand U6811 (N_6811,N_2885,N_3794);
nand U6812 (N_6812,N_3214,N_2742);
nor U6813 (N_6813,N_3929,N_4262);
or U6814 (N_6814,N_4321,N_2822);
nand U6815 (N_6815,N_3894,N_2536);
and U6816 (N_6816,N_3244,N_4146);
and U6817 (N_6817,N_3156,N_2962);
nand U6818 (N_6818,N_3307,N_2940);
nand U6819 (N_6819,N_3868,N_3638);
nand U6820 (N_6820,N_4833,N_4023);
nor U6821 (N_6821,N_3533,N_3440);
or U6822 (N_6822,N_3097,N_2505);
nor U6823 (N_6823,N_3490,N_2893);
or U6824 (N_6824,N_3159,N_3003);
nand U6825 (N_6825,N_2524,N_2875);
nor U6826 (N_6826,N_4598,N_4875);
or U6827 (N_6827,N_3165,N_4657);
nor U6828 (N_6828,N_2851,N_4120);
nand U6829 (N_6829,N_4385,N_2740);
and U6830 (N_6830,N_4156,N_3374);
and U6831 (N_6831,N_3039,N_4051);
nor U6832 (N_6832,N_4826,N_3387);
nand U6833 (N_6833,N_3245,N_4324);
nand U6834 (N_6834,N_3761,N_4819);
nor U6835 (N_6835,N_3836,N_2581);
nor U6836 (N_6836,N_4877,N_4455);
nor U6837 (N_6837,N_3830,N_4030);
or U6838 (N_6838,N_4377,N_4382);
nand U6839 (N_6839,N_3101,N_4868);
xnor U6840 (N_6840,N_3510,N_3190);
xnor U6841 (N_6841,N_2963,N_4610);
nand U6842 (N_6842,N_4195,N_4260);
and U6843 (N_6843,N_4778,N_3779);
nand U6844 (N_6844,N_4303,N_4474);
or U6845 (N_6845,N_3820,N_3581);
nand U6846 (N_6846,N_3016,N_4046);
nor U6847 (N_6847,N_3050,N_2820);
xor U6848 (N_6848,N_4600,N_4188);
and U6849 (N_6849,N_4514,N_4213);
or U6850 (N_6850,N_2874,N_3607);
or U6851 (N_6851,N_4946,N_2691);
nand U6852 (N_6852,N_3042,N_2901);
or U6853 (N_6853,N_4742,N_4661);
nand U6854 (N_6854,N_4353,N_3347);
and U6855 (N_6855,N_2738,N_3173);
xnor U6856 (N_6856,N_4943,N_3084);
nand U6857 (N_6857,N_4227,N_4320);
nor U6858 (N_6858,N_2743,N_3710);
and U6859 (N_6859,N_4525,N_3434);
and U6860 (N_6860,N_3387,N_4198);
or U6861 (N_6861,N_4480,N_2721);
xnor U6862 (N_6862,N_4318,N_4116);
nor U6863 (N_6863,N_3990,N_4085);
and U6864 (N_6864,N_2505,N_3547);
nand U6865 (N_6865,N_3500,N_4200);
xnor U6866 (N_6866,N_4797,N_4943);
nand U6867 (N_6867,N_3536,N_4658);
or U6868 (N_6868,N_3988,N_4473);
nand U6869 (N_6869,N_2504,N_3579);
nand U6870 (N_6870,N_4638,N_2518);
or U6871 (N_6871,N_3940,N_3603);
or U6872 (N_6872,N_4224,N_4968);
and U6873 (N_6873,N_3687,N_2970);
and U6874 (N_6874,N_4695,N_3518);
nand U6875 (N_6875,N_2677,N_4379);
nand U6876 (N_6876,N_4902,N_3026);
nor U6877 (N_6877,N_2622,N_3397);
xor U6878 (N_6878,N_2720,N_3614);
nand U6879 (N_6879,N_4313,N_3062);
nor U6880 (N_6880,N_3886,N_4191);
nand U6881 (N_6881,N_2712,N_3000);
nand U6882 (N_6882,N_3886,N_3085);
xor U6883 (N_6883,N_2814,N_4762);
or U6884 (N_6884,N_3405,N_4384);
xnor U6885 (N_6885,N_4188,N_4149);
or U6886 (N_6886,N_3009,N_3848);
nand U6887 (N_6887,N_4810,N_4797);
or U6888 (N_6888,N_4562,N_4406);
and U6889 (N_6889,N_3427,N_4777);
or U6890 (N_6890,N_3978,N_2732);
or U6891 (N_6891,N_3520,N_3667);
nor U6892 (N_6892,N_4664,N_4315);
nand U6893 (N_6893,N_3962,N_2533);
nand U6894 (N_6894,N_4985,N_4805);
or U6895 (N_6895,N_2969,N_3570);
nand U6896 (N_6896,N_3645,N_3025);
xor U6897 (N_6897,N_2514,N_3451);
nor U6898 (N_6898,N_4146,N_3297);
or U6899 (N_6899,N_4978,N_4400);
nor U6900 (N_6900,N_4389,N_3166);
and U6901 (N_6901,N_4086,N_3855);
nand U6902 (N_6902,N_2837,N_2908);
nor U6903 (N_6903,N_3232,N_4077);
nor U6904 (N_6904,N_4082,N_3947);
or U6905 (N_6905,N_4073,N_3076);
nand U6906 (N_6906,N_4518,N_4024);
nor U6907 (N_6907,N_2663,N_3311);
xnor U6908 (N_6908,N_3377,N_3110);
and U6909 (N_6909,N_2634,N_4012);
and U6910 (N_6910,N_4879,N_4390);
nor U6911 (N_6911,N_4926,N_3172);
or U6912 (N_6912,N_3827,N_4881);
and U6913 (N_6913,N_2557,N_4122);
nand U6914 (N_6914,N_4731,N_3720);
xor U6915 (N_6915,N_2699,N_2683);
xor U6916 (N_6916,N_3142,N_3381);
or U6917 (N_6917,N_2597,N_3949);
or U6918 (N_6918,N_3315,N_3602);
nand U6919 (N_6919,N_4297,N_4639);
and U6920 (N_6920,N_4764,N_2932);
nand U6921 (N_6921,N_3010,N_2757);
and U6922 (N_6922,N_4960,N_4105);
nor U6923 (N_6923,N_4505,N_4512);
and U6924 (N_6924,N_4665,N_4365);
or U6925 (N_6925,N_4358,N_4043);
or U6926 (N_6926,N_2931,N_4252);
and U6927 (N_6927,N_2749,N_3310);
and U6928 (N_6928,N_3161,N_3425);
nor U6929 (N_6929,N_3290,N_3801);
nor U6930 (N_6930,N_4688,N_2866);
and U6931 (N_6931,N_3902,N_3247);
nor U6932 (N_6932,N_4001,N_2702);
nand U6933 (N_6933,N_4410,N_3287);
nor U6934 (N_6934,N_2896,N_3062);
or U6935 (N_6935,N_4679,N_3206);
or U6936 (N_6936,N_3476,N_4868);
xor U6937 (N_6937,N_2846,N_2961);
and U6938 (N_6938,N_4226,N_3863);
or U6939 (N_6939,N_3274,N_3892);
and U6940 (N_6940,N_4547,N_4026);
and U6941 (N_6941,N_3581,N_3517);
nand U6942 (N_6942,N_3192,N_4615);
or U6943 (N_6943,N_2720,N_3861);
and U6944 (N_6944,N_4154,N_2850);
nand U6945 (N_6945,N_4853,N_2892);
nor U6946 (N_6946,N_4407,N_3733);
nor U6947 (N_6947,N_3537,N_3629);
and U6948 (N_6948,N_4892,N_3841);
nand U6949 (N_6949,N_4834,N_2945);
and U6950 (N_6950,N_2552,N_3404);
or U6951 (N_6951,N_3279,N_3390);
or U6952 (N_6952,N_4704,N_4503);
and U6953 (N_6953,N_3194,N_4066);
or U6954 (N_6954,N_3995,N_4476);
nor U6955 (N_6955,N_3283,N_4399);
and U6956 (N_6956,N_2641,N_4775);
nand U6957 (N_6957,N_3944,N_2744);
or U6958 (N_6958,N_3637,N_3781);
or U6959 (N_6959,N_2614,N_3555);
or U6960 (N_6960,N_3526,N_2812);
nor U6961 (N_6961,N_2660,N_3403);
nand U6962 (N_6962,N_2752,N_3797);
nor U6963 (N_6963,N_4667,N_3600);
or U6964 (N_6964,N_3680,N_4967);
and U6965 (N_6965,N_3313,N_2865);
or U6966 (N_6966,N_4750,N_3448);
and U6967 (N_6967,N_4176,N_3098);
nor U6968 (N_6968,N_4552,N_2884);
nor U6969 (N_6969,N_2814,N_3196);
and U6970 (N_6970,N_2888,N_3653);
or U6971 (N_6971,N_2573,N_2658);
nor U6972 (N_6972,N_4492,N_3005);
nor U6973 (N_6973,N_4493,N_4322);
or U6974 (N_6974,N_4924,N_3320);
or U6975 (N_6975,N_4581,N_4955);
and U6976 (N_6976,N_2846,N_4346);
and U6977 (N_6977,N_4713,N_2745);
nor U6978 (N_6978,N_3395,N_3587);
nor U6979 (N_6979,N_4849,N_4456);
nor U6980 (N_6980,N_4383,N_3239);
or U6981 (N_6981,N_3283,N_3804);
nor U6982 (N_6982,N_2958,N_4470);
and U6983 (N_6983,N_4765,N_3512);
and U6984 (N_6984,N_3394,N_4474);
nand U6985 (N_6985,N_2503,N_2827);
and U6986 (N_6986,N_3138,N_3373);
nand U6987 (N_6987,N_3414,N_4448);
or U6988 (N_6988,N_4230,N_2982);
nand U6989 (N_6989,N_3410,N_4721);
or U6990 (N_6990,N_4072,N_3359);
and U6991 (N_6991,N_2983,N_4130);
nor U6992 (N_6992,N_3894,N_2911);
nor U6993 (N_6993,N_2757,N_3444);
and U6994 (N_6994,N_2689,N_4504);
nand U6995 (N_6995,N_4216,N_2864);
nand U6996 (N_6996,N_3743,N_3382);
xor U6997 (N_6997,N_2710,N_2815);
and U6998 (N_6998,N_3966,N_3463);
or U6999 (N_6999,N_2507,N_2501);
xnor U7000 (N_7000,N_2795,N_4718);
and U7001 (N_7001,N_2617,N_2849);
and U7002 (N_7002,N_3957,N_4325);
nor U7003 (N_7003,N_4651,N_4043);
and U7004 (N_7004,N_4552,N_3602);
and U7005 (N_7005,N_3350,N_2570);
nor U7006 (N_7006,N_3457,N_2512);
nor U7007 (N_7007,N_3685,N_3041);
and U7008 (N_7008,N_3223,N_3221);
and U7009 (N_7009,N_4302,N_4887);
or U7010 (N_7010,N_3594,N_3546);
xnor U7011 (N_7011,N_2810,N_4478);
or U7012 (N_7012,N_3405,N_3452);
and U7013 (N_7013,N_3397,N_3374);
nor U7014 (N_7014,N_4097,N_3764);
nand U7015 (N_7015,N_4385,N_3421);
nand U7016 (N_7016,N_4651,N_3642);
nand U7017 (N_7017,N_4937,N_4706);
and U7018 (N_7018,N_3619,N_3859);
nor U7019 (N_7019,N_2825,N_2661);
nand U7020 (N_7020,N_4256,N_4674);
or U7021 (N_7021,N_4513,N_3730);
or U7022 (N_7022,N_4714,N_2754);
and U7023 (N_7023,N_3933,N_3005);
and U7024 (N_7024,N_3338,N_4703);
nor U7025 (N_7025,N_2743,N_4418);
xor U7026 (N_7026,N_4163,N_4052);
nand U7027 (N_7027,N_4008,N_4676);
nand U7028 (N_7028,N_4956,N_3392);
nor U7029 (N_7029,N_3858,N_4819);
xnor U7030 (N_7030,N_3706,N_2559);
xor U7031 (N_7031,N_3238,N_3395);
nor U7032 (N_7032,N_4720,N_3334);
xor U7033 (N_7033,N_2968,N_4041);
or U7034 (N_7034,N_3166,N_4680);
xor U7035 (N_7035,N_2670,N_4008);
nand U7036 (N_7036,N_2596,N_3807);
nand U7037 (N_7037,N_3836,N_3667);
nand U7038 (N_7038,N_2756,N_2619);
or U7039 (N_7039,N_3908,N_4260);
nor U7040 (N_7040,N_3166,N_4097);
nor U7041 (N_7041,N_4289,N_3574);
nor U7042 (N_7042,N_2534,N_2770);
nor U7043 (N_7043,N_3731,N_4764);
or U7044 (N_7044,N_3552,N_3449);
nor U7045 (N_7045,N_2646,N_4655);
nor U7046 (N_7046,N_3605,N_4199);
nand U7047 (N_7047,N_3515,N_4262);
nor U7048 (N_7048,N_4566,N_3344);
xnor U7049 (N_7049,N_4753,N_3713);
or U7050 (N_7050,N_4720,N_2678);
nor U7051 (N_7051,N_2743,N_4571);
nor U7052 (N_7052,N_2555,N_4044);
nand U7053 (N_7053,N_4760,N_2693);
or U7054 (N_7054,N_3248,N_4664);
nand U7055 (N_7055,N_3063,N_4509);
and U7056 (N_7056,N_4007,N_2715);
nor U7057 (N_7057,N_3714,N_4122);
nand U7058 (N_7058,N_4457,N_4533);
nand U7059 (N_7059,N_2860,N_4208);
nor U7060 (N_7060,N_4259,N_3839);
or U7061 (N_7061,N_3384,N_2691);
nand U7062 (N_7062,N_4899,N_3975);
nor U7063 (N_7063,N_3186,N_3725);
nor U7064 (N_7064,N_3762,N_2768);
xnor U7065 (N_7065,N_2617,N_4829);
and U7066 (N_7066,N_3310,N_3832);
and U7067 (N_7067,N_4095,N_4295);
and U7068 (N_7068,N_4402,N_3364);
or U7069 (N_7069,N_3466,N_4863);
xor U7070 (N_7070,N_2580,N_3103);
nor U7071 (N_7071,N_4192,N_4135);
or U7072 (N_7072,N_3388,N_3485);
or U7073 (N_7073,N_2681,N_4630);
nand U7074 (N_7074,N_3565,N_4025);
nor U7075 (N_7075,N_3927,N_4907);
nor U7076 (N_7076,N_3824,N_4938);
nand U7077 (N_7077,N_4080,N_4418);
and U7078 (N_7078,N_2985,N_4098);
nand U7079 (N_7079,N_3290,N_3750);
or U7080 (N_7080,N_4021,N_4198);
xor U7081 (N_7081,N_3230,N_3578);
nor U7082 (N_7082,N_3860,N_2982);
or U7083 (N_7083,N_4004,N_4799);
and U7084 (N_7084,N_3323,N_2870);
xnor U7085 (N_7085,N_3504,N_3385);
nand U7086 (N_7086,N_4854,N_3052);
nand U7087 (N_7087,N_4106,N_3824);
nor U7088 (N_7088,N_4960,N_3512);
nor U7089 (N_7089,N_2997,N_4104);
or U7090 (N_7090,N_3295,N_3102);
nand U7091 (N_7091,N_3763,N_2829);
or U7092 (N_7092,N_4813,N_4912);
or U7093 (N_7093,N_4630,N_2941);
nor U7094 (N_7094,N_4992,N_4090);
or U7095 (N_7095,N_3452,N_4866);
xnor U7096 (N_7096,N_4418,N_4365);
and U7097 (N_7097,N_3132,N_4158);
or U7098 (N_7098,N_2765,N_4852);
or U7099 (N_7099,N_3991,N_4539);
nand U7100 (N_7100,N_4011,N_3015);
nor U7101 (N_7101,N_4589,N_2594);
or U7102 (N_7102,N_3193,N_4489);
and U7103 (N_7103,N_3799,N_4237);
xnor U7104 (N_7104,N_3421,N_3751);
and U7105 (N_7105,N_4354,N_4585);
nand U7106 (N_7106,N_3347,N_4064);
or U7107 (N_7107,N_2971,N_4909);
or U7108 (N_7108,N_3305,N_4224);
xor U7109 (N_7109,N_2600,N_3909);
nor U7110 (N_7110,N_3629,N_2860);
or U7111 (N_7111,N_2907,N_4742);
and U7112 (N_7112,N_3195,N_4465);
nand U7113 (N_7113,N_2629,N_3339);
nand U7114 (N_7114,N_2540,N_4784);
nand U7115 (N_7115,N_4723,N_3032);
or U7116 (N_7116,N_2847,N_2885);
nor U7117 (N_7117,N_4966,N_4149);
and U7118 (N_7118,N_3933,N_2803);
nor U7119 (N_7119,N_2893,N_4920);
nor U7120 (N_7120,N_2890,N_4218);
or U7121 (N_7121,N_2663,N_3626);
nor U7122 (N_7122,N_4106,N_4441);
nor U7123 (N_7123,N_4980,N_4060);
and U7124 (N_7124,N_2933,N_3056);
nand U7125 (N_7125,N_4447,N_3792);
nor U7126 (N_7126,N_3028,N_4182);
nor U7127 (N_7127,N_2790,N_3513);
or U7128 (N_7128,N_4895,N_3931);
nand U7129 (N_7129,N_4256,N_4949);
or U7130 (N_7130,N_3444,N_3714);
or U7131 (N_7131,N_4323,N_3984);
nor U7132 (N_7132,N_4297,N_4555);
or U7133 (N_7133,N_4942,N_3508);
or U7134 (N_7134,N_2526,N_4608);
nor U7135 (N_7135,N_4099,N_3645);
and U7136 (N_7136,N_3186,N_3493);
or U7137 (N_7137,N_3181,N_3108);
nand U7138 (N_7138,N_4429,N_2792);
xor U7139 (N_7139,N_3349,N_4796);
and U7140 (N_7140,N_3950,N_4949);
nand U7141 (N_7141,N_3699,N_2759);
nor U7142 (N_7142,N_3115,N_4446);
or U7143 (N_7143,N_3595,N_2515);
and U7144 (N_7144,N_2957,N_4359);
or U7145 (N_7145,N_3877,N_3620);
nor U7146 (N_7146,N_3306,N_3171);
or U7147 (N_7147,N_4270,N_2684);
or U7148 (N_7148,N_3512,N_3384);
nand U7149 (N_7149,N_4262,N_3390);
and U7150 (N_7150,N_4917,N_3375);
nor U7151 (N_7151,N_2593,N_3781);
or U7152 (N_7152,N_3545,N_3931);
and U7153 (N_7153,N_4629,N_3124);
and U7154 (N_7154,N_2928,N_4708);
and U7155 (N_7155,N_3959,N_4934);
or U7156 (N_7156,N_3247,N_3234);
nor U7157 (N_7157,N_4322,N_3672);
and U7158 (N_7158,N_4061,N_2953);
and U7159 (N_7159,N_4797,N_4913);
and U7160 (N_7160,N_4981,N_4017);
xor U7161 (N_7161,N_4856,N_4149);
nand U7162 (N_7162,N_4401,N_2825);
nand U7163 (N_7163,N_3682,N_2514);
or U7164 (N_7164,N_4739,N_3587);
nor U7165 (N_7165,N_4087,N_3880);
nor U7166 (N_7166,N_4158,N_3930);
or U7167 (N_7167,N_4234,N_4822);
or U7168 (N_7168,N_3537,N_2886);
or U7169 (N_7169,N_2878,N_3861);
and U7170 (N_7170,N_4955,N_4674);
nor U7171 (N_7171,N_3298,N_4731);
nand U7172 (N_7172,N_4906,N_3421);
or U7173 (N_7173,N_2594,N_3160);
nor U7174 (N_7174,N_4361,N_3162);
nor U7175 (N_7175,N_4929,N_4832);
nand U7176 (N_7176,N_3684,N_3022);
or U7177 (N_7177,N_4856,N_4963);
and U7178 (N_7178,N_3845,N_2749);
nand U7179 (N_7179,N_4708,N_2697);
nor U7180 (N_7180,N_4189,N_3081);
and U7181 (N_7181,N_2882,N_2591);
and U7182 (N_7182,N_4545,N_4541);
or U7183 (N_7183,N_4454,N_3701);
and U7184 (N_7184,N_4920,N_2907);
nand U7185 (N_7185,N_4244,N_2856);
and U7186 (N_7186,N_4947,N_3421);
nor U7187 (N_7187,N_4329,N_4564);
nor U7188 (N_7188,N_2641,N_4309);
and U7189 (N_7189,N_4587,N_4486);
or U7190 (N_7190,N_4216,N_2689);
or U7191 (N_7191,N_3133,N_4673);
nand U7192 (N_7192,N_2930,N_3230);
nor U7193 (N_7193,N_3263,N_3455);
nand U7194 (N_7194,N_4396,N_3555);
xnor U7195 (N_7195,N_3287,N_4497);
and U7196 (N_7196,N_3154,N_3137);
nand U7197 (N_7197,N_4336,N_3680);
nor U7198 (N_7198,N_3030,N_2777);
or U7199 (N_7199,N_3855,N_4284);
or U7200 (N_7200,N_4213,N_3939);
nor U7201 (N_7201,N_3338,N_2692);
nor U7202 (N_7202,N_3644,N_2876);
nor U7203 (N_7203,N_4441,N_4858);
and U7204 (N_7204,N_3239,N_3844);
or U7205 (N_7205,N_4481,N_3703);
nor U7206 (N_7206,N_4274,N_3695);
xor U7207 (N_7207,N_4145,N_4154);
and U7208 (N_7208,N_4865,N_2621);
nand U7209 (N_7209,N_3160,N_2570);
nand U7210 (N_7210,N_3879,N_4657);
or U7211 (N_7211,N_4844,N_4325);
nor U7212 (N_7212,N_4903,N_4335);
or U7213 (N_7213,N_4975,N_3889);
and U7214 (N_7214,N_4389,N_3781);
nand U7215 (N_7215,N_4448,N_3225);
nor U7216 (N_7216,N_3214,N_4287);
or U7217 (N_7217,N_3377,N_4647);
nor U7218 (N_7218,N_4694,N_2925);
and U7219 (N_7219,N_2898,N_3910);
and U7220 (N_7220,N_2726,N_3875);
and U7221 (N_7221,N_4298,N_3584);
xnor U7222 (N_7222,N_3197,N_4235);
or U7223 (N_7223,N_4874,N_4372);
and U7224 (N_7224,N_4108,N_4330);
nor U7225 (N_7225,N_3716,N_3277);
xor U7226 (N_7226,N_4100,N_4219);
nand U7227 (N_7227,N_3267,N_3619);
nor U7228 (N_7228,N_2696,N_3031);
or U7229 (N_7229,N_4711,N_2701);
nor U7230 (N_7230,N_3737,N_4127);
and U7231 (N_7231,N_2801,N_3351);
or U7232 (N_7232,N_2848,N_2863);
nand U7233 (N_7233,N_3929,N_3313);
nand U7234 (N_7234,N_4567,N_3550);
xnor U7235 (N_7235,N_3389,N_3614);
and U7236 (N_7236,N_2957,N_2789);
or U7237 (N_7237,N_2804,N_4363);
nand U7238 (N_7238,N_4082,N_3884);
nand U7239 (N_7239,N_4978,N_4654);
nor U7240 (N_7240,N_3541,N_3420);
xor U7241 (N_7241,N_2755,N_3404);
or U7242 (N_7242,N_4956,N_4694);
nor U7243 (N_7243,N_4737,N_2529);
nor U7244 (N_7244,N_3896,N_2893);
nand U7245 (N_7245,N_4942,N_3059);
nand U7246 (N_7246,N_3110,N_3583);
nand U7247 (N_7247,N_3152,N_3183);
xnor U7248 (N_7248,N_4895,N_3624);
nand U7249 (N_7249,N_4498,N_4018);
nor U7250 (N_7250,N_4484,N_2572);
or U7251 (N_7251,N_4798,N_4851);
nor U7252 (N_7252,N_4838,N_3906);
or U7253 (N_7253,N_4301,N_4898);
and U7254 (N_7254,N_4602,N_3454);
nor U7255 (N_7255,N_4744,N_3977);
nor U7256 (N_7256,N_3527,N_3786);
nor U7257 (N_7257,N_3729,N_2798);
nand U7258 (N_7258,N_4799,N_4223);
and U7259 (N_7259,N_3688,N_4633);
or U7260 (N_7260,N_3845,N_3201);
nand U7261 (N_7261,N_3320,N_4736);
and U7262 (N_7262,N_3150,N_2512);
and U7263 (N_7263,N_4943,N_2638);
xnor U7264 (N_7264,N_4256,N_4486);
nand U7265 (N_7265,N_3562,N_3434);
or U7266 (N_7266,N_3960,N_4976);
nand U7267 (N_7267,N_3294,N_3574);
and U7268 (N_7268,N_2556,N_2596);
nor U7269 (N_7269,N_4379,N_3499);
xor U7270 (N_7270,N_4411,N_4150);
xnor U7271 (N_7271,N_3405,N_2797);
and U7272 (N_7272,N_4128,N_4503);
or U7273 (N_7273,N_2596,N_4310);
and U7274 (N_7274,N_4263,N_2995);
or U7275 (N_7275,N_3615,N_3871);
and U7276 (N_7276,N_3884,N_4166);
and U7277 (N_7277,N_4713,N_4916);
xnor U7278 (N_7278,N_4751,N_3998);
or U7279 (N_7279,N_4146,N_2684);
and U7280 (N_7280,N_3675,N_4301);
nor U7281 (N_7281,N_4925,N_2548);
and U7282 (N_7282,N_2651,N_2673);
nor U7283 (N_7283,N_3205,N_2532);
nand U7284 (N_7284,N_3701,N_3575);
nand U7285 (N_7285,N_3687,N_3433);
nor U7286 (N_7286,N_4180,N_3576);
nand U7287 (N_7287,N_2653,N_4769);
xor U7288 (N_7288,N_3373,N_3361);
nand U7289 (N_7289,N_3017,N_4366);
nand U7290 (N_7290,N_3277,N_2797);
and U7291 (N_7291,N_4643,N_3018);
nand U7292 (N_7292,N_3523,N_4988);
nand U7293 (N_7293,N_3332,N_3253);
or U7294 (N_7294,N_4089,N_3414);
and U7295 (N_7295,N_3044,N_2605);
or U7296 (N_7296,N_3306,N_2632);
xnor U7297 (N_7297,N_4747,N_2993);
and U7298 (N_7298,N_3757,N_2710);
xor U7299 (N_7299,N_3659,N_4190);
and U7300 (N_7300,N_4835,N_2912);
and U7301 (N_7301,N_2586,N_2869);
and U7302 (N_7302,N_3893,N_3109);
nor U7303 (N_7303,N_2917,N_4460);
nand U7304 (N_7304,N_4423,N_3419);
nor U7305 (N_7305,N_4737,N_3668);
or U7306 (N_7306,N_4188,N_4984);
and U7307 (N_7307,N_3615,N_3488);
and U7308 (N_7308,N_3598,N_2665);
or U7309 (N_7309,N_3456,N_3374);
xnor U7310 (N_7310,N_4636,N_4825);
or U7311 (N_7311,N_2659,N_4887);
or U7312 (N_7312,N_2695,N_4417);
or U7313 (N_7313,N_3503,N_4497);
or U7314 (N_7314,N_4315,N_3469);
or U7315 (N_7315,N_3266,N_2678);
nor U7316 (N_7316,N_3780,N_4334);
and U7317 (N_7317,N_2787,N_2867);
and U7318 (N_7318,N_4528,N_4902);
and U7319 (N_7319,N_4681,N_4272);
or U7320 (N_7320,N_3931,N_3564);
and U7321 (N_7321,N_4978,N_3393);
or U7322 (N_7322,N_4885,N_4341);
nand U7323 (N_7323,N_4554,N_4882);
nand U7324 (N_7324,N_3932,N_2888);
nand U7325 (N_7325,N_3328,N_4879);
and U7326 (N_7326,N_2861,N_3609);
nand U7327 (N_7327,N_4994,N_4578);
nor U7328 (N_7328,N_3675,N_2992);
or U7329 (N_7329,N_3794,N_3296);
nand U7330 (N_7330,N_4021,N_3402);
xor U7331 (N_7331,N_4353,N_3478);
and U7332 (N_7332,N_2799,N_4290);
nand U7333 (N_7333,N_4076,N_4820);
nor U7334 (N_7334,N_2877,N_3323);
or U7335 (N_7335,N_4794,N_3770);
and U7336 (N_7336,N_4640,N_3714);
or U7337 (N_7337,N_2578,N_3914);
xnor U7338 (N_7338,N_4301,N_4268);
or U7339 (N_7339,N_3702,N_4914);
xnor U7340 (N_7340,N_3703,N_4719);
nor U7341 (N_7341,N_3910,N_4282);
and U7342 (N_7342,N_4409,N_3765);
nand U7343 (N_7343,N_3103,N_4996);
or U7344 (N_7344,N_2774,N_3273);
nor U7345 (N_7345,N_3247,N_2532);
nand U7346 (N_7346,N_2600,N_2737);
nand U7347 (N_7347,N_3956,N_3709);
or U7348 (N_7348,N_3301,N_4670);
or U7349 (N_7349,N_2561,N_3378);
xor U7350 (N_7350,N_4152,N_2693);
nand U7351 (N_7351,N_4946,N_3592);
nand U7352 (N_7352,N_2640,N_4215);
or U7353 (N_7353,N_4532,N_4048);
nand U7354 (N_7354,N_3642,N_3330);
or U7355 (N_7355,N_4708,N_4921);
nor U7356 (N_7356,N_2638,N_3544);
xnor U7357 (N_7357,N_2908,N_4005);
nor U7358 (N_7358,N_3484,N_4431);
and U7359 (N_7359,N_3226,N_4577);
nor U7360 (N_7360,N_4114,N_4692);
nor U7361 (N_7361,N_3051,N_3363);
or U7362 (N_7362,N_4297,N_3901);
and U7363 (N_7363,N_2578,N_3087);
and U7364 (N_7364,N_3180,N_3408);
nand U7365 (N_7365,N_4171,N_2743);
nand U7366 (N_7366,N_2591,N_3735);
xor U7367 (N_7367,N_3056,N_3752);
xnor U7368 (N_7368,N_3196,N_4314);
or U7369 (N_7369,N_3684,N_2845);
nor U7370 (N_7370,N_3668,N_3639);
nor U7371 (N_7371,N_3745,N_4546);
and U7372 (N_7372,N_2617,N_3171);
nand U7373 (N_7373,N_2656,N_4434);
or U7374 (N_7374,N_4345,N_3797);
nand U7375 (N_7375,N_3622,N_3671);
nand U7376 (N_7376,N_3012,N_4322);
nand U7377 (N_7377,N_3911,N_2978);
nor U7378 (N_7378,N_3764,N_3847);
nand U7379 (N_7379,N_2533,N_4293);
and U7380 (N_7380,N_3965,N_3228);
nand U7381 (N_7381,N_2733,N_2700);
nand U7382 (N_7382,N_3798,N_4256);
nor U7383 (N_7383,N_2852,N_3680);
or U7384 (N_7384,N_3612,N_3637);
or U7385 (N_7385,N_4778,N_3301);
or U7386 (N_7386,N_3472,N_3922);
xor U7387 (N_7387,N_2916,N_3931);
or U7388 (N_7388,N_4808,N_2589);
and U7389 (N_7389,N_3110,N_2916);
or U7390 (N_7390,N_4438,N_2781);
and U7391 (N_7391,N_2969,N_4062);
nor U7392 (N_7392,N_3128,N_3613);
nor U7393 (N_7393,N_3563,N_4578);
nand U7394 (N_7394,N_3689,N_2558);
and U7395 (N_7395,N_4565,N_2641);
or U7396 (N_7396,N_3666,N_4928);
or U7397 (N_7397,N_3126,N_4452);
nand U7398 (N_7398,N_4267,N_3435);
nor U7399 (N_7399,N_4391,N_2611);
nand U7400 (N_7400,N_4198,N_3381);
nor U7401 (N_7401,N_3189,N_4243);
and U7402 (N_7402,N_2913,N_4574);
nor U7403 (N_7403,N_4401,N_3028);
or U7404 (N_7404,N_4900,N_4297);
and U7405 (N_7405,N_4018,N_4699);
nand U7406 (N_7406,N_3077,N_3876);
or U7407 (N_7407,N_4440,N_3392);
and U7408 (N_7408,N_4786,N_4771);
or U7409 (N_7409,N_3801,N_3011);
nand U7410 (N_7410,N_3990,N_4985);
and U7411 (N_7411,N_4537,N_4092);
or U7412 (N_7412,N_4511,N_2532);
nor U7413 (N_7413,N_4645,N_4945);
nor U7414 (N_7414,N_4853,N_3141);
or U7415 (N_7415,N_2747,N_3723);
nand U7416 (N_7416,N_4649,N_3310);
or U7417 (N_7417,N_2687,N_3586);
nor U7418 (N_7418,N_3039,N_3174);
and U7419 (N_7419,N_4587,N_4924);
and U7420 (N_7420,N_2805,N_2590);
or U7421 (N_7421,N_3784,N_3915);
nor U7422 (N_7422,N_3394,N_2508);
and U7423 (N_7423,N_3041,N_3846);
nand U7424 (N_7424,N_2568,N_4836);
nand U7425 (N_7425,N_3319,N_4788);
nand U7426 (N_7426,N_4016,N_4378);
nand U7427 (N_7427,N_3747,N_4116);
and U7428 (N_7428,N_3480,N_4484);
nor U7429 (N_7429,N_4290,N_4752);
or U7430 (N_7430,N_3567,N_2853);
and U7431 (N_7431,N_3127,N_3332);
nand U7432 (N_7432,N_4538,N_2917);
nand U7433 (N_7433,N_2545,N_4746);
nand U7434 (N_7434,N_4575,N_2697);
and U7435 (N_7435,N_2631,N_3978);
nor U7436 (N_7436,N_4811,N_3479);
or U7437 (N_7437,N_4432,N_4430);
and U7438 (N_7438,N_4447,N_3247);
or U7439 (N_7439,N_3850,N_3534);
xnor U7440 (N_7440,N_3887,N_3944);
nand U7441 (N_7441,N_4523,N_4962);
or U7442 (N_7442,N_4398,N_2809);
nand U7443 (N_7443,N_4754,N_4158);
and U7444 (N_7444,N_4796,N_4987);
nor U7445 (N_7445,N_4169,N_3426);
nor U7446 (N_7446,N_4999,N_3549);
or U7447 (N_7447,N_2832,N_4732);
and U7448 (N_7448,N_3074,N_2537);
nor U7449 (N_7449,N_4769,N_4130);
nor U7450 (N_7450,N_3267,N_3349);
and U7451 (N_7451,N_4294,N_3324);
nand U7452 (N_7452,N_4569,N_4244);
and U7453 (N_7453,N_4041,N_4543);
xor U7454 (N_7454,N_4197,N_4211);
nor U7455 (N_7455,N_3185,N_3499);
or U7456 (N_7456,N_2646,N_4105);
nor U7457 (N_7457,N_2539,N_3117);
or U7458 (N_7458,N_3420,N_4531);
nand U7459 (N_7459,N_3159,N_3774);
and U7460 (N_7460,N_4483,N_3468);
nor U7461 (N_7461,N_3912,N_4109);
nor U7462 (N_7462,N_2705,N_3454);
nand U7463 (N_7463,N_4345,N_2629);
and U7464 (N_7464,N_4576,N_2531);
nor U7465 (N_7465,N_3297,N_2923);
or U7466 (N_7466,N_3851,N_3410);
nand U7467 (N_7467,N_3752,N_4719);
nor U7468 (N_7468,N_4062,N_3947);
and U7469 (N_7469,N_3616,N_2531);
nor U7470 (N_7470,N_4971,N_4546);
nand U7471 (N_7471,N_4922,N_3558);
or U7472 (N_7472,N_2694,N_3002);
nand U7473 (N_7473,N_4801,N_3402);
nand U7474 (N_7474,N_4742,N_3850);
or U7475 (N_7475,N_4198,N_4234);
and U7476 (N_7476,N_3768,N_3317);
or U7477 (N_7477,N_3176,N_2762);
nand U7478 (N_7478,N_4540,N_2827);
nor U7479 (N_7479,N_3511,N_4673);
nand U7480 (N_7480,N_3979,N_2745);
nand U7481 (N_7481,N_3880,N_4363);
nor U7482 (N_7482,N_4814,N_4308);
nor U7483 (N_7483,N_3657,N_4669);
or U7484 (N_7484,N_4958,N_3111);
nor U7485 (N_7485,N_3746,N_2966);
and U7486 (N_7486,N_2889,N_3103);
and U7487 (N_7487,N_4020,N_2604);
and U7488 (N_7488,N_4173,N_3005);
and U7489 (N_7489,N_4909,N_2584);
nor U7490 (N_7490,N_2619,N_4723);
and U7491 (N_7491,N_3566,N_4164);
nor U7492 (N_7492,N_4386,N_4155);
nor U7493 (N_7493,N_4411,N_2705);
or U7494 (N_7494,N_4621,N_3561);
xnor U7495 (N_7495,N_4359,N_4920);
or U7496 (N_7496,N_4194,N_3816);
or U7497 (N_7497,N_2802,N_3788);
and U7498 (N_7498,N_3638,N_4362);
and U7499 (N_7499,N_3580,N_3992);
nand U7500 (N_7500,N_7192,N_6698);
nand U7501 (N_7501,N_6402,N_7041);
nor U7502 (N_7502,N_6024,N_5175);
nand U7503 (N_7503,N_6890,N_6144);
and U7504 (N_7504,N_6414,N_7305);
and U7505 (N_7505,N_5480,N_7129);
and U7506 (N_7506,N_7232,N_5074);
and U7507 (N_7507,N_5772,N_7210);
nand U7508 (N_7508,N_7385,N_7440);
nand U7509 (N_7509,N_6759,N_5788);
or U7510 (N_7510,N_6128,N_6358);
nand U7511 (N_7511,N_6374,N_6828);
and U7512 (N_7512,N_6001,N_6880);
and U7513 (N_7513,N_6127,N_7081);
nand U7514 (N_7514,N_5129,N_6220);
or U7515 (N_7515,N_5849,N_7143);
and U7516 (N_7516,N_6671,N_5429);
nor U7517 (N_7517,N_5859,N_6302);
or U7518 (N_7518,N_5860,N_5867);
nor U7519 (N_7519,N_6961,N_6555);
and U7520 (N_7520,N_7278,N_6784);
xor U7521 (N_7521,N_6930,N_5560);
and U7522 (N_7522,N_6705,N_5575);
nand U7523 (N_7523,N_6049,N_5930);
and U7524 (N_7524,N_6694,N_6308);
or U7525 (N_7525,N_5080,N_7387);
xor U7526 (N_7526,N_6281,N_5692);
or U7527 (N_7527,N_5681,N_5227);
nor U7528 (N_7528,N_5231,N_5726);
or U7529 (N_7529,N_6500,N_5907);
or U7530 (N_7530,N_6467,N_7146);
nor U7531 (N_7531,N_6681,N_5220);
xor U7532 (N_7532,N_6752,N_5365);
nor U7533 (N_7533,N_5178,N_5533);
or U7534 (N_7534,N_5263,N_6431);
xor U7535 (N_7535,N_6711,N_5845);
nand U7536 (N_7536,N_5795,N_5577);
or U7537 (N_7537,N_5386,N_6917);
or U7538 (N_7538,N_6976,N_6861);
nand U7539 (N_7539,N_5761,N_5456);
or U7540 (N_7540,N_7399,N_5688);
and U7541 (N_7541,N_6549,N_5975);
xor U7542 (N_7542,N_5725,N_6359);
nand U7543 (N_7543,N_7486,N_6348);
nand U7544 (N_7544,N_5439,N_6337);
nand U7545 (N_7545,N_6137,N_5590);
nor U7546 (N_7546,N_5164,N_6903);
or U7547 (N_7547,N_6959,N_6148);
xnor U7548 (N_7548,N_6043,N_6717);
nor U7549 (N_7549,N_6026,N_5781);
and U7550 (N_7550,N_6532,N_7026);
xor U7551 (N_7551,N_5827,N_5819);
and U7552 (N_7552,N_5700,N_6092);
and U7553 (N_7553,N_5797,N_7494);
nor U7554 (N_7554,N_6588,N_6172);
and U7555 (N_7555,N_6617,N_7358);
xor U7556 (N_7556,N_7082,N_6856);
nand U7557 (N_7557,N_7227,N_5589);
nor U7558 (N_7558,N_5665,N_7222);
and U7559 (N_7559,N_5088,N_6912);
nor U7560 (N_7560,N_5019,N_5059);
nand U7561 (N_7561,N_5919,N_5655);
and U7562 (N_7562,N_5335,N_6246);
nand U7563 (N_7563,N_7018,N_6296);
nor U7564 (N_7564,N_7117,N_5448);
nor U7565 (N_7565,N_6088,N_5704);
and U7566 (N_7566,N_6622,N_5251);
nand U7567 (N_7567,N_5558,N_7005);
or U7568 (N_7568,N_5286,N_5821);
xor U7569 (N_7569,N_5553,N_6289);
and U7570 (N_7570,N_6342,N_5699);
nand U7571 (N_7571,N_6401,N_6407);
nand U7572 (N_7572,N_5464,N_6769);
and U7573 (N_7573,N_7072,N_6245);
nand U7574 (N_7574,N_6270,N_5653);
nor U7575 (N_7575,N_7073,N_6412);
nand U7576 (N_7576,N_5153,N_7107);
and U7577 (N_7577,N_7067,N_6792);
or U7578 (N_7578,N_5021,N_5817);
nand U7579 (N_7579,N_6167,N_6019);
nand U7580 (N_7580,N_5974,N_5115);
or U7581 (N_7581,N_5015,N_6802);
nand U7582 (N_7582,N_5596,N_6487);
and U7583 (N_7583,N_6803,N_7221);
nand U7584 (N_7584,N_7001,N_7231);
nor U7585 (N_7585,N_7195,N_6195);
nor U7586 (N_7586,N_5350,N_6844);
xor U7587 (N_7587,N_5205,N_5525);
or U7588 (N_7588,N_5512,N_5741);
nor U7589 (N_7589,N_7391,N_7178);
or U7590 (N_7590,N_7382,N_6193);
and U7591 (N_7591,N_7027,N_6614);
nand U7592 (N_7592,N_6371,N_6483);
nand U7593 (N_7593,N_7075,N_5082);
nor U7594 (N_7594,N_6409,N_6768);
or U7595 (N_7595,N_7393,N_5013);
nor U7596 (N_7596,N_7009,N_7176);
nor U7597 (N_7597,N_5351,N_6729);
and U7598 (N_7598,N_7314,N_6874);
and U7599 (N_7599,N_5820,N_5330);
and U7600 (N_7600,N_7159,N_6875);
nor U7601 (N_7601,N_6536,N_6251);
nand U7602 (N_7602,N_5482,N_6764);
and U7603 (N_7603,N_5275,N_6869);
or U7604 (N_7604,N_7434,N_6562);
nand U7605 (N_7605,N_6247,N_5994);
and U7606 (N_7606,N_7042,N_7337);
and U7607 (N_7607,N_5672,N_7428);
nand U7608 (N_7608,N_6336,N_5876);
nor U7609 (N_7609,N_6382,N_5454);
nor U7610 (N_7610,N_5186,N_5691);
and U7611 (N_7611,N_6130,N_6704);
xnor U7612 (N_7612,N_6369,N_5564);
or U7613 (N_7613,N_6706,N_6641);
nand U7614 (N_7614,N_5874,N_6165);
and U7615 (N_7615,N_6177,N_6899);
and U7616 (N_7616,N_5355,N_6415);
nor U7617 (N_7617,N_6811,N_5864);
or U7618 (N_7618,N_6421,N_6633);
nor U7619 (N_7619,N_6314,N_5219);
and U7620 (N_7620,N_5204,N_6993);
and U7621 (N_7621,N_6135,N_5005);
nor U7622 (N_7622,N_6827,N_7164);
or U7623 (N_7623,N_7083,N_5111);
nor U7624 (N_7624,N_6581,N_6922);
nor U7625 (N_7625,N_5910,N_6076);
nor U7626 (N_7626,N_6604,N_5522);
nor U7627 (N_7627,N_6395,N_6638);
nor U7628 (N_7628,N_7172,N_5187);
nand U7629 (N_7629,N_6994,N_5238);
nor U7630 (N_7630,N_5708,N_5904);
or U7631 (N_7631,N_5764,N_5625);
or U7632 (N_7632,N_5307,N_6339);
nor U7633 (N_7633,N_6377,N_5089);
or U7634 (N_7634,N_6373,N_6256);
and U7635 (N_7635,N_7152,N_5740);
nand U7636 (N_7636,N_5812,N_5595);
and U7637 (N_7637,N_6654,N_5176);
nand U7638 (N_7638,N_6674,N_6361);
nor U7639 (N_7639,N_6435,N_6808);
or U7640 (N_7640,N_7286,N_5034);
nand U7641 (N_7641,N_7304,N_6664);
nand U7642 (N_7642,N_6597,N_6689);
or U7643 (N_7643,N_5562,N_5780);
and U7644 (N_7644,N_5866,N_6884);
and U7645 (N_7645,N_6385,N_7071);
nor U7646 (N_7646,N_6080,N_6175);
nor U7647 (N_7647,N_5573,N_6533);
and U7648 (N_7648,N_6998,N_5640);
nand U7649 (N_7649,N_7413,N_6901);
or U7650 (N_7650,N_6790,N_5478);
or U7651 (N_7651,N_5011,N_6486);
or U7652 (N_7652,N_6754,N_7483);
nor U7653 (N_7653,N_5416,N_6058);
and U7654 (N_7654,N_5132,N_7058);
nand U7655 (N_7655,N_5824,N_7332);
or U7656 (N_7656,N_5534,N_5375);
nand U7657 (N_7657,N_6267,N_6701);
nor U7658 (N_7658,N_5254,N_6408);
or U7659 (N_7659,N_6871,N_6189);
nor U7660 (N_7660,N_5619,N_6521);
or U7661 (N_7661,N_7420,N_5169);
xor U7662 (N_7662,N_5802,N_7061);
nand U7663 (N_7663,N_5686,N_5807);
and U7664 (N_7664,N_6797,N_5731);
xor U7665 (N_7665,N_5104,N_6439);
nand U7666 (N_7666,N_5250,N_5308);
or U7667 (N_7667,N_6012,N_5184);
and U7668 (N_7668,N_5632,N_6956);
or U7669 (N_7669,N_5932,N_7468);
nor U7670 (N_7670,N_5157,N_7013);
nand U7671 (N_7671,N_6113,N_7250);
or U7672 (N_7672,N_5567,N_5607);
nor U7673 (N_7673,N_7247,N_6438);
nor U7674 (N_7674,N_6843,N_6206);
and U7675 (N_7675,N_5384,N_7321);
nor U7676 (N_7676,N_7031,N_5721);
xor U7677 (N_7677,N_5479,N_7438);
nand U7678 (N_7678,N_6918,N_5044);
nor U7679 (N_7679,N_5498,N_5126);
nor U7680 (N_7680,N_5391,N_5535);
or U7681 (N_7681,N_5912,N_6883);
or U7682 (N_7682,N_6651,N_7189);
or U7683 (N_7683,N_5077,N_5197);
or U7684 (N_7684,N_6158,N_6849);
nor U7685 (N_7685,N_6623,N_6809);
nand U7686 (N_7686,N_5278,N_5417);
or U7687 (N_7687,N_7492,N_6603);
or U7688 (N_7688,N_6326,N_6211);
nand U7689 (N_7689,N_5201,N_5159);
or U7690 (N_7690,N_5276,N_5986);
and U7691 (N_7691,N_6366,N_7331);
or U7692 (N_7692,N_5897,N_5387);
xor U7693 (N_7693,N_5646,N_6305);
or U7694 (N_7694,N_5621,N_7423);
nand U7695 (N_7695,N_5360,N_7444);
nor U7696 (N_7696,N_6821,N_5582);
or U7697 (N_7697,N_5893,N_7229);
nand U7698 (N_7698,N_6062,N_7113);
and U7699 (N_7699,N_5289,N_6071);
nor U7700 (N_7700,N_7171,N_7351);
nand U7701 (N_7701,N_5938,N_5177);
nor U7702 (N_7702,N_5639,N_6205);
and U7703 (N_7703,N_6052,N_5326);
xnor U7704 (N_7704,N_7476,N_5841);
or U7705 (N_7705,N_6464,N_5240);
or U7706 (N_7706,N_7433,N_7044);
nand U7707 (N_7707,N_6198,N_5940);
or U7708 (N_7708,N_7131,N_5946);
and U7709 (N_7709,N_6744,N_6064);
nand U7710 (N_7710,N_6571,N_5853);
or U7711 (N_7711,N_5218,N_6108);
or U7712 (N_7712,N_5285,N_6368);
nand U7713 (N_7713,N_7003,N_5331);
or U7714 (N_7714,N_7103,N_5713);
nand U7715 (N_7715,N_6653,N_5829);
or U7716 (N_7716,N_5789,N_5294);
nor U7717 (N_7717,N_5084,N_6756);
and U7718 (N_7718,N_6834,N_5787);
xnor U7719 (N_7719,N_6287,N_5142);
nand U7720 (N_7720,N_6009,N_6452);
nor U7721 (N_7721,N_7283,N_6410);
nand U7722 (N_7722,N_7353,N_7275);
or U7723 (N_7723,N_5357,N_6645);
nor U7724 (N_7724,N_5170,N_5848);
xnor U7725 (N_7725,N_7267,N_7421);
and U7726 (N_7726,N_5636,N_6320);
nand U7727 (N_7727,N_6553,N_6561);
or U7728 (N_7728,N_6788,N_5614);
nor U7729 (N_7729,N_6757,N_6657);
nor U7730 (N_7730,N_6978,N_6665);
xor U7731 (N_7731,N_5791,N_7065);
nand U7732 (N_7732,N_5673,N_6806);
or U7733 (N_7733,N_7461,N_7435);
nand U7734 (N_7734,N_7099,N_6637);
nand U7735 (N_7735,N_7274,N_5923);
xnor U7736 (N_7736,N_6776,N_7289);
nand U7737 (N_7737,N_5341,N_6225);
nand U7738 (N_7738,N_5586,N_5282);
and U7739 (N_7739,N_6789,N_6384);
and U7740 (N_7740,N_7422,N_5000);
nor U7741 (N_7741,N_6558,N_6141);
nand U7742 (N_7742,N_7108,N_5948);
xor U7743 (N_7743,N_5638,N_5099);
or U7744 (N_7744,N_6125,N_5751);
nor U7745 (N_7745,N_5046,N_6544);
nand U7746 (N_7746,N_5894,N_5947);
or U7747 (N_7747,N_5068,N_5269);
or U7748 (N_7748,N_5846,N_5580);
or U7749 (N_7749,N_6609,N_5854);
and U7750 (N_7750,N_6306,N_5112);
nand U7751 (N_7751,N_5016,N_5996);
and U7752 (N_7752,N_7115,N_6526);
nor U7753 (N_7753,N_7404,N_6568);
nor U7754 (N_7754,N_5968,N_5306);
or U7755 (N_7755,N_6892,N_6512);
xnor U7756 (N_7756,N_5650,N_5642);
nor U7757 (N_7757,N_5413,N_7038);
and U7758 (N_7758,N_5381,N_5428);
nand U7759 (N_7759,N_5838,N_6666);
nand U7760 (N_7760,N_6829,N_7153);
nand U7761 (N_7761,N_5389,N_7070);
xor U7762 (N_7762,N_7139,N_6101);
and U7763 (N_7763,N_7259,N_6819);
or U7764 (N_7764,N_6787,N_6584);
nor U7765 (N_7765,N_6037,N_5312);
nand U7766 (N_7766,N_5152,N_7484);
nor U7767 (N_7767,N_7087,N_7365);
and U7768 (N_7768,N_5143,N_6971);
xor U7769 (N_7769,N_5421,N_5096);
nand U7770 (N_7770,N_5531,N_5903);
nand U7771 (N_7771,N_6970,N_5154);
xnor U7772 (N_7772,N_7347,N_7206);
nor U7773 (N_7773,N_5235,N_6535);
or U7774 (N_7774,N_7246,N_5031);
nor U7775 (N_7775,N_6904,N_6753);
nand U7776 (N_7776,N_5784,N_5014);
nor U7777 (N_7777,N_5835,N_5051);
or U7778 (N_7778,N_5773,N_6360);
nor U7779 (N_7779,N_6157,N_5268);
or U7780 (N_7780,N_5075,N_5766);
xnor U7781 (N_7781,N_6611,N_7478);
nor U7782 (N_7782,N_6840,N_5383);
and U7783 (N_7783,N_7248,N_6825);
nand U7784 (N_7784,N_5033,N_6031);
nand U7785 (N_7785,N_5976,N_7211);
nor U7786 (N_7786,N_5258,N_6923);
and U7787 (N_7787,N_5527,N_5255);
nor U7788 (N_7788,N_5882,N_7460);
nand U7789 (N_7789,N_6404,N_7091);
nand U7790 (N_7790,N_6746,N_5585);
and U7791 (N_7791,N_6985,N_6854);
nand U7792 (N_7792,N_5737,N_6117);
nor U7793 (N_7793,N_6453,N_6065);
nand U7794 (N_7794,N_5136,N_5786);
nand U7795 (N_7795,N_6463,N_5735);
xor U7796 (N_7796,N_6488,N_5984);
or U7797 (N_7797,N_7207,N_5182);
nand U7798 (N_7798,N_6285,N_7261);
nand U7799 (N_7799,N_6362,N_6044);
and U7800 (N_7800,N_5674,N_7357);
nand U7801 (N_7801,N_6109,N_7174);
and U7802 (N_7802,N_5723,N_5362);
nor U7803 (N_7803,N_7374,N_5376);
or U7804 (N_7804,N_5851,N_7348);
nor U7805 (N_7805,N_5979,N_6477);
and U7806 (N_7806,N_5371,N_5800);
or U7807 (N_7807,N_5367,N_6028);
or U7808 (N_7808,N_6136,N_5895);
or U7809 (N_7809,N_6629,N_5314);
nor U7810 (N_7810,N_6672,N_6718);
nor U7811 (N_7811,N_6731,N_7424);
and U7812 (N_7812,N_5406,N_7403);
and U7813 (N_7813,N_6264,N_5592);
and U7814 (N_7814,N_5847,N_5191);
nand U7815 (N_7815,N_5135,N_5581);
and U7816 (N_7816,N_5506,N_5647);
or U7817 (N_7817,N_6406,N_6481);
nor U7818 (N_7818,N_6831,N_5379);
nor U7819 (N_7819,N_6086,N_6582);
nor U7820 (N_7820,N_6299,N_6707);
nor U7821 (N_7821,N_7277,N_7471);
or U7822 (N_7822,N_7355,N_6594);
nor U7823 (N_7823,N_6210,N_6250);
xor U7824 (N_7824,N_5125,N_6104);
nor U7825 (N_7825,N_5465,N_6761);
nor U7826 (N_7826,N_6986,N_6386);
or U7827 (N_7827,N_6462,N_7214);
or U7828 (N_7828,N_7238,N_7350);
xor U7829 (N_7829,N_7158,N_6868);
nand U7830 (N_7830,N_6898,N_6879);
nand U7831 (N_7831,N_5805,N_5523);
and U7832 (N_7832,N_7418,N_5792);
nand U7833 (N_7833,N_7459,N_6608);
and U7834 (N_7834,N_7055,N_5271);
or U7835 (N_7835,N_5412,N_5452);
and U7836 (N_7836,N_6094,N_5668);
and U7837 (N_7837,N_5004,N_5453);
nor U7838 (N_7838,N_5451,N_5949);
and U7839 (N_7839,N_5460,N_6590);
or U7840 (N_7840,N_7118,N_6347);
nand U7841 (N_7841,N_7485,N_5296);
or U7842 (N_7842,N_6039,N_6659);
and U7843 (N_7843,N_5680,N_7193);
nand U7844 (N_7844,N_6459,N_7161);
or U7845 (N_7845,N_5816,N_6498);
nor U7846 (N_7846,N_5888,N_6005);
nand U7847 (N_7847,N_6426,N_6566);
and U7848 (N_7848,N_6820,N_5818);
nor U7849 (N_7849,N_5980,N_5317);
or U7850 (N_7850,N_7015,N_5755);
nand U7851 (N_7851,N_5587,N_5105);
nand U7852 (N_7852,N_5635,N_7006);
and U7853 (N_7853,N_7346,N_6773);
or U7854 (N_7854,N_5257,N_7452);
and U7855 (N_7855,N_6911,N_5970);
nand U7856 (N_7856,N_5556,N_6276);
or U7857 (N_7857,N_6182,N_6714);
xnor U7858 (N_7858,N_6393,N_7062);
nand U7859 (N_7859,N_6628,N_5877);
or U7860 (N_7860,N_6798,N_5260);
nor U7861 (N_7861,N_5950,N_5880);
nand U7862 (N_7862,N_6447,N_6537);
or U7863 (N_7863,N_5608,N_5995);
or U7864 (N_7864,N_6215,N_6344);
nor U7865 (N_7865,N_6548,N_6280);
xnor U7866 (N_7866,N_6980,N_5693);
and U7867 (N_7867,N_6400,N_5858);
nand U7868 (N_7868,N_6639,N_6397);
nand U7869 (N_7869,N_5229,N_5094);
nor U7870 (N_7870,N_6579,N_6090);
xnor U7871 (N_7871,N_6363,N_5151);
nor U7872 (N_7872,N_6485,N_7345);
nand U7873 (N_7873,N_7464,N_5663);
and U7874 (N_7874,N_6927,N_6456);
or U7875 (N_7875,N_5166,N_6710);
nor U7876 (N_7876,N_7095,N_5041);
nand U7877 (N_7877,N_6838,N_5739);
and U7878 (N_7878,N_5656,N_7388);
or U7879 (N_7879,N_6387,N_6403);
nor U7880 (N_7880,N_5881,N_5863);
nor U7881 (N_7881,N_5039,N_7169);
xor U7882 (N_7882,N_5615,N_6100);
nor U7883 (N_7883,N_5572,N_6778);
or U7884 (N_7884,N_7303,N_5952);
nand U7885 (N_7885,N_6252,N_5516);
or U7886 (N_7886,N_6390,N_5422);
nand U7887 (N_7887,N_6375,N_6054);
or U7888 (N_7888,N_5079,N_5270);
nor U7889 (N_7889,N_5651,N_5511);
xnor U7890 (N_7890,N_7043,N_7446);
nand U7891 (N_7891,N_6800,N_6991);
nor U7892 (N_7892,N_7450,N_5494);
and U7893 (N_7893,N_6235,N_7023);
or U7894 (N_7894,N_6557,N_7328);
or U7895 (N_7895,N_6910,N_6942);
or U7896 (N_7896,N_6097,N_7364);
nor U7897 (N_7897,N_7296,N_7100);
nand U7898 (N_7898,N_6230,N_5137);
nor U7899 (N_7899,N_5985,N_5069);
and U7900 (N_7900,N_5469,N_5108);
nor U7901 (N_7901,N_7132,N_5850);
xnor U7902 (N_7902,N_5073,N_6528);
nor U7903 (N_7903,N_7280,N_5338);
nand U7904 (N_7904,N_6207,N_6338);
nand U7905 (N_7905,N_5554,N_6697);
and U7906 (N_7906,N_7341,N_6351);
and U7907 (N_7907,N_5687,N_6983);
and U7908 (N_7908,N_5419,N_5916);
nand U7909 (N_7909,N_5411,N_6962);
or U7910 (N_7910,N_5685,N_7122);
nor U7911 (N_7911,N_5121,N_7472);
nand U7912 (N_7912,N_7137,N_5489);
nor U7913 (N_7913,N_6936,N_6345);
and U7914 (N_7914,N_6743,N_5645);
or U7915 (N_7915,N_5915,N_5192);
and U7916 (N_7916,N_5728,N_6480);
nor U7917 (N_7917,N_6265,N_7390);
nand U7918 (N_7918,N_7299,N_6621);
or U7919 (N_7919,N_5983,N_7212);
or U7920 (N_7920,N_5618,N_7409);
or U7921 (N_7921,N_5212,N_6947);
and U7922 (N_7922,N_6661,N_5216);
xnor U7923 (N_7923,N_6479,N_5902);
nand U7924 (N_7924,N_6132,N_5203);
nor U7925 (N_7925,N_6900,N_5738);
nand U7926 (N_7926,N_5472,N_6029);
nand U7927 (N_7927,N_5281,N_6988);
nand U7928 (N_7928,N_6739,N_6124);
nand U7929 (N_7929,N_7307,N_5103);
and U7930 (N_7930,N_5359,N_6020);
nand U7931 (N_7931,N_5246,N_6679);
xnor U7932 (N_7932,N_7033,N_6855);
nand U7933 (N_7933,N_5467,N_5702);
or U7934 (N_7934,N_6888,N_6692);
and U7935 (N_7935,N_5070,N_5461);
or U7936 (N_7936,N_6428,N_7090);
nand U7937 (N_7937,N_5414,N_5502);
or U7938 (N_7938,N_6138,N_5481);
nor U7939 (N_7939,N_6059,N_5403);
and U7940 (N_7940,N_6979,N_5694);
or U7941 (N_7941,N_5868,N_5669);
nor U7942 (N_7942,N_5521,N_6253);
nor U7943 (N_7943,N_5458,N_5316);
nand U7944 (N_7944,N_6376,N_6862);
or U7945 (N_7945,N_7301,N_6217);
and U7946 (N_7946,N_7255,N_5374);
nor U7947 (N_7947,N_6448,N_5658);
and U7948 (N_7948,N_6640,N_5488);
or U7949 (N_7949,N_5487,N_5266);
or U7950 (N_7950,N_6069,N_6143);
or U7951 (N_7951,N_7149,N_6813);
nand U7952 (N_7952,N_7311,N_7088);
nand U7953 (N_7953,N_5844,N_6823);
nor U7954 (N_7954,N_6243,N_5420);
xnor U7955 (N_7955,N_7263,N_6134);
nand U7956 (N_7956,N_6902,N_6853);
and U7957 (N_7957,N_5124,N_5752);
nor U7958 (N_7958,N_6035,N_7205);
and U7959 (N_7959,N_5920,N_6105);
xnor U7960 (N_7960,N_5008,N_5783);
and U7961 (N_7961,N_5449,N_6686);
and U7962 (N_7962,N_7487,N_6047);
and U7963 (N_7963,N_6765,N_5349);
nor U7964 (N_7964,N_5892,N_6027);
and U7965 (N_7965,N_5883,N_5138);
or U7966 (N_7966,N_7086,N_6449);
nand U7967 (N_7967,N_5253,N_7019);
nand U7968 (N_7968,N_7011,N_6084);
or U7969 (N_7969,N_6506,N_7094);
or U7970 (N_7970,N_6939,N_7257);
and U7971 (N_7971,N_5295,N_5028);
xnor U7972 (N_7972,N_6214,N_7002);
or U7973 (N_7973,N_6596,N_6967);
or U7974 (N_7974,N_5392,N_6323);
nor U7975 (N_7975,N_5279,N_6471);
nor U7976 (N_7976,N_6200,N_7306);
and U7977 (N_7977,N_6122,N_6926);
nor U7978 (N_7978,N_5826,N_6437);
nand U7979 (N_7979,N_6328,N_6891);
or U7980 (N_7980,N_7226,N_5555);
nand U7981 (N_7981,N_7110,N_5243);
and U7982 (N_7982,N_5017,N_6146);
and U7983 (N_7983,N_7089,N_7431);
and U7984 (N_7984,N_6965,N_7408);
and U7985 (N_7985,N_6048,N_5675);
nand U7986 (N_7986,N_6602,N_6139);
xor U7987 (N_7987,N_6017,N_5901);
nand U7988 (N_7988,N_7217,N_5442);
or U7989 (N_7989,N_5407,N_7335);
or U7990 (N_7990,N_5963,N_5734);
nor U7991 (N_7991,N_5520,N_6233);
nand U7992 (N_7992,N_6997,N_6990);
nand U7993 (N_7993,N_7151,N_5109);
or U7994 (N_7994,N_5162,N_6524);
nand U7995 (N_7995,N_5388,N_6392);
nor U7996 (N_7996,N_7123,N_5358);
nand U7997 (N_7997,N_5654,N_6775);
or U7998 (N_7998,N_5301,N_5774);
or U7999 (N_7999,N_6591,N_7298);
or U8000 (N_8000,N_6176,N_5834);
and U8001 (N_8001,N_6068,N_6966);
or U8002 (N_8002,N_6418,N_5353);
or U8003 (N_8003,N_6896,N_6620);
and U8004 (N_8004,N_7470,N_5493);
nor U8005 (N_8005,N_6682,N_7173);
and U8006 (N_8006,N_5049,N_7441);
or U8007 (N_8007,N_5236,N_6785);
nor U8008 (N_8008,N_5973,N_5909);
nand U8009 (N_8009,N_6836,N_6041);
or U8010 (N_8010,N_6424,N_7445);
xor U8011 (N_8011,N_6209,N_5346);
and U8012 (N_8012,N_6432,N_6238);
or U8013 (N_8013,N_6042,N_5095);
nand U8014 (N_8014,N_5568,N_6630);
or U8015 (N_8015,N_5840,N_5302);
and U8016 (N_8016,N_6475,N_6070);
nor U8017 (N_8017,N_5706,N_6156);
nor U8018 (N_8018,N_5811,N_5408);
xor U8019 (N_8019,N_6199,N_6841);
nand U8020 (N_8020,N_5280,N_7479);
nor U8021 (N_8021,N_6786,N_6915);
and U8022 (N_8022,N_6131,N_5855);
nor U8023 (N_8023,N_6554,N_5382);
or U8024 (N_8024,N_5473,N_6703);
nor U8025 (N_8025,N_6212,N_6810);
and U8026 (N_8026,N_5610,N_5823);
nor U8027 (N_8027,N_7154,N_7265);
xor U8028 (N_8028,N_7096,N_6249);
nor U8029 (N_8029,N_7367,N_5398);
nor U8030 (N_8030,N_6616,N_5010);
nor U8031 (N_8031,N_6619,N_5955);
and U8032 (N_8032,N_5604,N_6675);
and U8033 (N_8033,N_5569,N_6905);
nand U8034 (N_8034,N_5274,N_6708);
nor U8035 (N_8035,N_5746,N_7354);
xor U8036 (N_8036,N_6738,N_6063);
and U8037 (N_8037,N_5232,N_6164);
nand U8038 (N_8038,N_5328,N_5156);
nand U8039 (N_8039,N_6313,N_7190);
and U8040 (N_8040,N_5050,N_5509);
nor U8041 (N_8041,N_5131,N_6218);
or U8042 (N_8042,N_6631,N_6153);
nor U8043 (N_8043,N_6564,N_5063);
nand U8044 (N_8044,N_6974,N_6067);
nor U8045 (N_8045,N_5207,N_6534);
and U8046 (N_8046,N_7180,N_7380);
and U8047 (N_8047,N_5623,N_6589);
nand U8048 (N_8048,N_6115,N_7356);
or U8049 (N_8049,N_6142,N_7064);
xnor U8050 (N_8050,N_5574,N_5933);
or U8051 (N_8051,N_7457,N_7051);
nand U8052 (N_8052,N_7454,N_6712);
and U8053 (N_8053,N_6852,N_6914);
nand U8054 (N_8054,N_5972,N_7377);
nor U8055 (N_8055,N_6388,N_5048);
xor U8056 (N_8056,N_5743,N_6670);
and U8057 (N_8057,N_6257,N_6322);
or U8058 (N_8058,N_6601,N_7035);
nand U8059 (N_8059,N_5620,N_5475);
and U8060 (N_8060,N_6678,N_6893);
nand U8061 (N_8061,N_5714,N_5961);
and U8062 (N_8062,N_5332,N_6283);
and U8063 (N_8063,N_6413,N_5223);
or U8064 (N_8064,N_6937,N_7451);
nor U8065 (N_8065,N_7053,N_6955);
and U8066 (N_8066,N_5311,N_6021);
nor U8067 (N_8067,N_6749,N_6545);
nand U8068 (N_8068,N_7135,N_5434);
or U8069 (N_8069,N_6010,N_6636);
and U8070 (N_8070,N_5689,N_7028);
nor U8071 (N_8071,N_6762,N_6443);
and U8072 (N_8072,N_5913,N_6740);
nand U8073 (N_8073,N_5093,N_6180);
nand U8074 (N_8074,N_6734,N_5796);
nand U8075 (N_8075,N_5652,N_6239);
and U8076 (N_8076,N_5168,N_5870);
or U8077 (N_8077,N_6550,N_5147);
and U8078 (N_8078,N_6179,N_7437);
nor U8079 (N_8079,N_5200,N_6719);
and U8080 (N_8080,N_5230,N_5293);
and U8081 (N_8081,N_6864,N_5340);
nand U8082 (N_8082,N_6329,N_7106);
and U8083 (N_8083,N_5744,N_7344);
nor U8084 (N_8084,N_7204,N_5173);
nand U8085 (N_8085,N_5072,N_6162);
nand U8086 (N_8086,N_6969,N_5703);
nor U8087 (N_8087,N_6953,N_6952);
xor U8088 (N_8088,N_5497,N_6040);
nand U8089 (N_8089,N_5291,N_5875);
nand U8090 (N_8090,N_6599,N_6702);
or U8091 (N_8091,N_6085,N_5036);
xor U8092 (N_8092,N_6972,N_6007);
nor U8093 (N_8093,N_5445,N_6002);
xnor U8094 (N_8094,N_5061,N_5730);
nand U8095 (N_8095,N_7223,N_7329);
xor U8096 (N_8096,N_7276,N_6807);
nand U8097 (N_8097,N_6538,N_5141);
and U8098 (N_8098,N_5202,N_6006);
or U8099 (N_8099,N_6722,N_6794);
nor U8100 (N_8100,N_6307,N_7313);
or U8101 (N_8101,N_5865,N_5160);
and U8102 (N_8102,N_6531,N_6170);
xor U8103 (N_8103,N_5579,N_5249);
xnor U8104 (N_8104,N_5884,N_6430);
xnor U8105 (N_8105,N_5519,N_5127);
nand U8106 (N_8106,N_6099,N_5116);
or U8107 (N_8107,N_6755,N_6457);
or U8108 (N_8108,N_5378,N_5529);
xor U8109 (N_8109,N_6546,N_6159);
nor U8110 (N_8110,N_5641,N_6812);
nand U8111 (N_8111,N_5552,N_6444);
nor U8112 (N_8112,N_7427,N_5999);
nand U8113 (N_8113,N_7228,N_6129);
and U8114 (N_8114,N_6520,N_5801);
nor U8115 (N_8115,N_6379,N_5622);
nor U8116 (N_8116,N_5966,N_5071);
and U8117 (N_8117,N_5158,N_6261);
or U8118 (N_8118,N_5447,N_5626);
and U8119 (N_8119,N_6502,N_6446);
nor U8120 (N_8120,N_5588,N_6325);
xor U8121 (N_8121,N_6995,N_5396);
or U8122 (N_8122,N_7037,N_5815);
nor U8123 (N_8123,N_6767,N_6881);
nand U8124 (N_8124,N_6658,N_6886);
and U8125 (N_8125,N_6022,N_6963);
and U8126 (N_8126,N_6992,N_5886);
xnor U8127 (N_8127,N_6213,N_6316);
nand U8128 (N_8128,N_6656,N_6928);
and U8129 (N_8129,N_5705,N_6349);
or U8130 (N_8130,N_5964,N_7370);
xnor U8131 (N_8131,N_7245,N_5085);
and U8132 (N_8132,N_5078,N_5532);
nor U8133 (N_8133,N_5517,N_6934);
nand U8134 (N_8134,N_6288,N_7373);
or U8135 (N_8135,N_6758,N_6751);
nor U8136 (N_8136,N_7068,N_5594);
and U8137 (N_8137,N_6867,N_6511);
nand U8138 (N_8138,N_6669,N_6833);
nor U8139 (N_8139,N_6624,N_5133);
nand U8140 (N_8140,N_7324,N_6556);
nor U8141 (N_8141,N_7249,N_6150);
nor U8142 (N_8142,N_6223,N_6793);
nand U8143 (N_8143,N_7102,N_5929);
or U8144 (N_8144,N_6495,N_6093);
or U8145 (N_8145,N_6695,N_7111);
nor U8146 (N_8146,N_5234,N_5352);
nand U8147 (N_8147,N_5025,N_7138);
nand U8148 (N_8148,N_6760,N_7239);
nand U8149 (N_8149,N_5500,N_7203);
and U8150 (N_8150,N_6747,N_7200);
nor U8151 (N_8151,N_6219,N_5290);
or U8152 (N_8152,N_7184,N_6723);
or U8153 (N_8153,N_5678,N_5758);
xor U8154 (N_8154,N_6642,N_7493);
nand U8155 (N_8155,N_7140,N_5993);
nand U8156 (N_8156,N_7079,N_6216);
nor U8157 (N_8157,N_6932,N_5637);
nand U8158 (N_8158,N_6814,N_5917);
or U8159 (N_8159,N_5287,N_5003);
nor U8160 (N_8160,N_7279,N_6957);
nor U8161 (N_8161,N_6748,N_5722);
nor U8162 (N_8162,N_7287,N_5771);
nand U8163 (N_8163,N_6297,N_6585);
or U8164 (N_8164,N_6454,N_6433);
nor U8165 (N_8165,N_5617,N_6460);
and U8166 (N_8166,N_6473,N_6075);
and U8167 (N_8167,N_5707,N_7025);
nor U8168 (N_8168,N_7260,N_6034);
nand U8169 (N_8169,N_7179,N_5657);
or U8170 (N_8170,N_7216,N_6103);
nor U8171 (N_8171,N_6763,N_6365);
and U8172 (N_8172,N_6133,N_5931);
nand U8173 (N_8173,N_5483,N_6050);
or U8174 (N_8174,N_7389,N_6291);
nand U8175 (N_8175,N_5992,N_7124);
and U8176 (N_8176,N_5262,N_6441);
nand U8177 (N_8177,N_5334,N_7490);
xor U8178 (N_8178,N_5020,N_6203);
and U8179 (N_8179,N_5941,N_5583);
nand U8180 (N_8180,N_7215,N_5206);
and U8181 (N_8181,N_5466,N_6023);
nand U8182 (N_8182,N_7098,N_5643);
nand U8183 (N_8183,N_7256,N_6237);
nand U8184 (N_8184,N_6032,N_6303);
or U8185 (N_8185,N_5491,N_6155);
nand U8186 (N_8186,N_7021,N_6184);
nor U8187 (N_8187,N_7209,N_5778);
nand U8188 (N_8188,N_5748,N_6356);
nand U8189 (N_8189,N_7213,N_6552);
and U8190 (N_8190,N_6254,N_6482);
or U8191 (N_8191,N_6476,N_6000);
nor U8192 (N_8192,N_5612,N_6004);
nor U8193 (N_8193,N_6906,N_5463);
or U8194 (N_8194,N_5769,N_5914);
nor U8195 (N_8195,N_6140,N_6352);
and U8196 (N_8196,N_5584,N_6774);
nor U8197 (N_8197,N_5027,N_5146);
nand U8198 (N_8198,N_5776,N_5601);
nor U8199 (N_8199,N_5241,N_5150);
nor U8200 (N_8200,N_7318,N_6522);
nor U8201 (N_8201,N_6173,N_6916);
and U8202 (N_8202,N_5062,N_6394);
and U8203 (N_8203,N_5321,N_5830);
nor U8204 (N_8204,N_7240,N_6655);
nand U8205 (N_8205,N_5749,N_6924);
nand U8206 (N_8206,N_5965,N_6771);
and U8207 (N_8207,N_6721,N_5043);
xnor U8208 (N_8208,N_6673,N_7077);
and U8209 (N_8209,N_6191,N_7398);
nor U8210 (N_8210,N_6355,N_5944);
nor U8211 (N_8211,N_5981,N_5924);
nor U8212 (N_8212,N_7092,N_7114);
nand U8213 (N_8213,N_6839,N_7397);
nand U8214 (N_8214,N_6713,N_7066);
nor U8215 (N_8215,N_6977,N_6635);
and U8216 (N_8216,N_7175,N_6822);
nand U8217 (N_8217,N_6647,N_5120);
nor U8218 (N_8218,N_5198,N_5283);
nor U8219 (N_8219,N_7000,N_5083);
nand U8220 (N_8220,N_5264,N_7453);
xor U8221 (N_8221,N_6341,N_7269);
and U8222 (N_8222,N_5245,N_7254);
nor U8223 (N_8223,N_5753,N_5822);
and U8224 (N_8224,N_5443,N_5717);
and U8225 (N_8225,N_6033,N_5861);
xor U8226 (N_8226,N_5742,N_7182);
and U8227 (N_8227,N_6515,N_5785);
nand U8228 (N_8228,N_5304,N_5002);
or U8229 (N_8229,N_5624,N_5444);
or U8230 (N_8230,N_5117,N_6181);
nand U8231 (N_8231,N_5609,N_6419);
or U8232 (N_8232,N_6742,N_5869);
nand U8233 (N_8233,N_7336,N_5505);
nor U8234 (N_8234,N_6882,N_5171);
or U8235 (N_8235,N_6372,N_6318);
nand U8236 (N_8236,N_5145,N_5053);
nor U8237 (N_8237,N_5323,N_6529);
and U8238 (N_8238,N_5394,N_6733);
nor U8239 (N_8239,N_7417,N_5559);
nand U8240 (N_8240,N_7155,N_5431);
xnor U8241 (N_8241,N_6688,N_6683);
nor U8242 (N_8242,N_5377,N_6805);
and U8243 (N_8243,N_7236,N_5035);
and U8244 (N_8244,N_5193,N_6948);
or U8245 (N_8245,N_7343,N_7251);
xnor U8246 (N_8246,N_7295,N_5045);
nand U8247 (N_8247,N_5066,N_7376);
and U8248 (N_8248,N_6317,N_5102);
and U8249 (N_8249,N_6417,N_6098);
nand U8250 (N_8250,N_6649,N_6866);
nor U8251 (N_8251,N_5934,N_6872);
nand U8252 (N_8252,N_6396,N_5485);
and U8253 (N_8253,N_6563,N_5300);
or U8254 (N_8254,N_6279,N_6580);
or U8255 (N_8255,N_5370,N_6527);
or U8256 (N_8256,N_5030,N_5712);
or U8257 (N_8257,N_6074,N_5055);
or U8258 (N_8258,N_5690,N_5911);
xor U8259 (N_8259,N_6737,N_7162);
and U8260 (N_8260,N_6038,N_6817);
or U8261 (N_8261,N_5404,N_7458);
or U8262 (N_8262,N_5361,N_5978);
nor U8263 (N_8263,N_7340,N_5977);
and U8264 (N_8264,N_7120,N_6848);
and U8265 (N_8265,N_7416,N_6693);
xnor U8266 (N_8266,N_5261,N_5477);
nor U8267 (N_8267,N_5715,N_5879);
and U8268 (N_8268,N_6440,N_5908);
and U8269 (N_8269,N_6434,N_7125);
or U8270 (N_8270,N_6652,N_6030);
nand U8271 (N_8271,N_6525,N_5987);
nor U8272 (N_8272,N_7291,N_5954);
xor U8273 (N_8273,N_6185,N_6465);
and U8274 (N_8274,N_5140,N_5779);
and U8275 (N_8275,N_6295,N_6147);
nand U8276 (N_8276,N_6333,N_7401);
or U8277 (N_8277,N_7379,N_5244);
and U8278 (N_8278,N_6425,N_6949);
or U8279 (N_8279,N_7187,N_5318);
and U8280 (N_8280,N_5327,N_5299);
nor U8281 (N_8281,N_6228,N_6878);
nand U8282 (N_8282,N_6015,N_5557);
nor U8283 (N_8283,N_5363,N_7167);
nand U8284 (N_8284,N_7406,N_6221);
and U8285 (N_8285,N_5199,N_6466);
xnor U8286 (N_8286,N_6540,N_6389);
and U8287 (N_8287,N_7126,N_6796);
nor U8288 (N_8288,N_5937,N_6676);
or U8289 (N_8289,N_6627,N_6102);
nor U8290 (N_8290,N_6335,N_5982);
nor U8291 (N_8291,N_7462,N_6648);
nand U8292 (N_8292,N_6196,N_5733);
nor U8293 (N_8293,N_5155,N_5969);
and U8294 (N_8294,N_6106,N_5067);
nor U8295 (N_8295,N_6981,N_5450);
and U8296 (N_8296,N_7292,N_6920);
nor U8297 (N_8297,N_6732,N_6650);
or U8298 (N_8298,N_5659,N_6999);
nor U8299 (N_8299,N_5369,N_6508);
xnor U8300 (N_8300,N_7467,N_5432);
nor U8301 (N_8301,N_6120,N_6166);
nor U8302 (N_8302,N_6091,N_5546);
nor U8303 (N_8303,N_6503,N_5056);
xnor U8304 (N_8304,N_7194,N_5179);
xnor U8305 (N_8305,N_7262,N_5189);
nor U8306 (N_8306,N_6208,N_6781);
or U8307 (N_8307,N_7225,N_5100);
or U8308 (N_8308,N_5390,N_5782);
or U8309 (N_8309,N_7273,N_6472);
nor U8310 (N_8310,N_7116,N_7439);
nor U8311 (N_8311,N_7268,N_6381);
and U8312 (N_8312,N_6859,N_5599);
nor U8313 (N_8313,N_6565,N_5081);
and U8314 (N_8314,N_7046,N_6750);
nand U8315 (N_8315,N_5697,N_6782);
nand U8316 (N_8316,N_5209,N_6575);
and U8317 (N_8317,N_6570,N_7330);
nand U8318 (N_8318,N_6057,N_6677);
nor U8319 (N_8319,N_6286,N_6436);
nand U8320 (N_8320,N_6489,N_6263);
nor U8321 (N_8321,N_7497,N_6857);
or U8322 (N_8322,N_5666,N_5898);
nor U8323 (N_8323,N_6301,N_5476);
nand U8324 (N_8324,N_6530,N_5676);
nand U8325 (N_8325,N_6931,N_6411);
nand U8326 (N_8326,N_6578,N_6229);
xor U8327 (N_8327,N_7372,N_5561);
nor U8328 (N_8328,N_5530,N_5945);
or U8329 (N_8329,N_7147,N_6583);
and U8330 (N_8330,N_7371,N_6946);
nor U8331 (N_8331,N_5167,N_5356);
and U8332 (N_8332,N_7366,N_7059);
xnor U8333 (N_8333,N_7480,N_5037);
nand U8334 (N_8334,N_6539,N_6255);
or U8335 (N_8335,N_6160,N_5899);
and U8336 (N_8336,N_5163,N_7230);
and U8337 (N_8337,N_6061,N_7375);
xor U8338 (N_8338,N_6567,N_7338);
and U8339 (N_8339,N_5648,N_6921);
nand U8340 (N_8340,N_5887,N_5309);
or U8341 (N_8341,N_7012,N_6107);
and U8342 (N_8342,N_6720,N_7201);
or U8343 (N_8343,N_7378,N_7078);
nor U8344 (N_8344,N_6493,N_5210);
nor U8345 (N_8345,N_5149,N_5727);
or U8346 (N_8346,N_6968,N_7322);
nand U8347 (N_8347,N_5393,N_6612);
nor U8348 (N_8348,N_6420,N_6735);
nor U8349 (N_8349,N_6398,N_6343);
xor U8350 (N_8350,N_7319,N_6663);
nand U8351 (N_8351,N_5225,N_5616);
and U8352 (N_8352,N_5507,N_6330);
or U8353 (N_8353,N_5926,N_5097);
nand U8354 (N_8354,N_5347,N_6877);
and U8355 (N_8355,N_6847,N_5591);
and U8356 (N_8356,N_6586,N_6518);
nand U8357 (N_8357,N_7465,N_5922);
or U8358 (N_8358,N_6236,N_5695);
nand U8359 (N_8359,N_7359,N_6818);
or U8360 (N_8360,N_6941,N_7309);
or U8361 (N_8361,N_5927,N_5878);
nor U8362 (N_8362,N_5436,N_6863);
or U8363 (N_8363,N_6304,N_6036);
and U8364 (N_8364,N_5720,N_5997);
and U8365 (N_8365,N_5188,N_7199);
nand U8366 (N_8366,N_7316,N_6560);
nor U8367 (N_8367,N_6272,N_6445);
or U8368 (N_8368,N_6492,N_7436);
nand U8369 (N_8369,N_5682,N_6592);
xnor U8370 (N_8370,N_6470,N_7191);
or U8371 (N_8371,N_6573,N_5825);
nor U8372 (N_8372,N_6699,N_7429);
or U8373 (N_8373,N_7144,N_5026);
or U8374 (N_8374,N_6095,N_5101);
nor U8375 (N_8375,N_6982,N_6851);
nand U8376 (N_8376,N_7057,N_7363);
nand U8377 (N_8377,N_7168,N_7142);
nor U8378 (N_8378,N_7333,N_6835);
nand U8379 (N_8379,N_7448,N_5042);
and U8380 (N_8380,N_5086,N_5918);
and U8381 (N_8381,N_5337,N_7016);
xor U8382 (N_8382,N_5076,N_5935);
nor U8383 (N_8383,N_5195,N_5603);
nand U8384 (N_8384,N_5925,N_5139);
nand U8385 (N_8385,N_6055,N_6242);
or U8386 (N_8386,N_7045,N_5354);
or U8387 (N_8387,N_6632,N_5563);
nand U8388 (N_8388,N_5134,N_5770);
or U8389 (N_8389,N_5988,N_6730);
and U8390 (N_8390,N_7266,N_5798);
xnor U8391 (N_8391,N_5122,N_7284);
and U8392 (N_8392,N_6954,N_7054);
or U8393 (N_8393,N_7360,N_5539);
nand U8394 (N_8394,N_5745,N_7281);
and U8395 (N_8395,N_6770,N_7177);
or U8396 (N_8396,N_6340,N_7270);
nor U8397 (N_8397,N_6378,N_6494);
nor U8398 (N_8398,N_5259,N_6079);
and U8399 (N_8399,N_7456,N_5185);
nand U8400 (N_8400,N_6727,N_5600);
or U8401 (N_8401,N_5729,N_7294);
nand U8402 (N_8402,N_5959,N_7362);
and U8403 (N_8403,N_5843,N_5891);
xor U8404 (N_8404,N_5342,N_6507);
or U8405 (N_8405,N_5329,N_6505);
xor U8406 (N_8406,N_5380,N_5344);
and U8407 (N_8407,N_7315,N_6008);
nand U8408 (N_8408,N_5183,N_7085);
and U8409 (N_8409,N_5064,N_7063);
nor U8410 (N_8410,N_6523,N_5065);
or U8411 (N_8411,N_6509,N_7425);
nand U8412 (N_8412,N_5644,N_7181);
and U8413 (N_8413,N_6996,N_5543);
and U8414 (N_8414,N_7339,N_5366);
nor U8415 (N_8415,N_5211,N_5091);
or U8416 (N_8416,N_6188,N_5526);
nand U8417 (N_8417,N_6274,N_5606);
nor U8418 (N_8418,N_7034,N_6779);
and U8419 (N_8419,N_5297,N_5711);
and U8420 (N_8420,N_5161,N_5459);
nor U8421 (N_8421,N_6815,N_6016);
nand U8422 (N_8422,N_7008,N_7121);
or U8423 (N_8423,N_5810,N_6960);
xor U8424 (N_8424,N_6543,N_6908);
or U8425 (N_8425,N_6046,N_7419);
nand U8426 (N_8426,N_5631,N_5284);
nand U8427 (N_8427,N_5990,N_5551);
nor U8428 (N_8428,N_5578,N_7400);
nor U8429 (N_8429,N_5768,N_5368);
and U8430 (N_8430,N_6478,N_6709);
and U8431 (N_8431,N_6178,N_5890);
nand U8432 (N_8432,N_7443,N_7481);
nor U8433 (N_8433,N_5438,N_6169);
nand U8434 (N_8434,N_7020,N_5277);
nor U8435 (N_8435,N_6935,N_6248);
nand U8436 (N_8436,N_6895,N_5496);
and U8437 (N_8437,N_6282,N_6187);
nand U8438 (N_8438,N_5292,N_5325);
xor U8439 (N_8439,N_5190,N_6346);
or U8440 (N_8440,N_7197,N_7396);
xor U8441 (N_8441,N_5098,N_7198);
or U8442 (N_8442,N_5305,N_5794);
xnor U8443 (N_8443,N_6940,N_5058);
nor U8444 (N_8444,N_5228,N_7290);
or U8445 (N_8445,N_6380,N_6309);
and U8446 (N_8446,N_6391,N_6060);
xor U8447 (N_8447,N_7145,N_6364);
and U8448 (N_8448,N_5710,N_5719);
nor U8449 (N_8449,N_7447,N_5597);
nand U8450 (N_8450,N_6275,N_5001);
nor U8451 (N_8451,N_7264,N_5222);
nor U8452 (N_8452,N_7157,N_6576);
and U8453 (N_8453,N_5627,N_6383);
and U8454 (N_8454,N_6950,N_6919);
xnor U8455 (N_8455,N_7032,N_7312);
or U8456 (N_8456,N_6298,N_5547);
and U8457 (N_8457,N_6837,N_5754);
and U8458 (N_8458,N_6266,N_5513);
or U8459 (N_8459,N_6011,N_5660);
and U8460 (N_8460,N_7036,N_7317);
or U8461 (N_8461,N_6232,N_6204);
and U8462 (N_8462,N_6680,N_5029);
or U8463 (N_8463,N_7488,N_5670);
nor U8464 (N_8464,N_5989,N_7234);
and U8465 (N_8465,N_5958,N_6192);
or U8466 (N_8466,N_6045,N_5399);
nor U8467 (N_8467,N_5433,N_7242);
nor U8468 (N_8468,N_5701,N_5732);
and U8469 (N_8469,N_5613,N_5446);
and U8470 (N_8470,N_7325,N_6168);
nor U8471 (N_8471,N_5397,N_5565);
and U8472 (N_8472,N_6154,N_6018);
nor U8473 (N_8473,N_5006,N_5873);
nor U8474 (N_8474,N_6577,N_6497);
and U8475 (N_8475,N_7449,N_5804);
and U8476 (N_8476,N_6271,N_5775);
nor U8477 (N_8477,N_5709,N_7049);
or U8478 (N_8478,N_5415,N_6643);
xnor U8479 (N_8479,N_6072,N_5018);
nand U8480 (N_8480,N_5090,N_7004);
nand U8481 (N_8481,N_7381,N_7300);
nand U8482 (N_8482,N_7386,N_6943);
xnor U8483 (N_8483,N_5953,N_6975);
and U8484 (N_8484,N_6224,N_7101);
or U8485 (N_8485,N_6290,N_6197);
nor U8486 (N_8486,N_5196,N_6987);
or U8487 (N_8487,N_7150,N_7410);
nand U8488 (N_8488,N_7412,N_7060);
xnor U8489 (N_8489,N_6114,N_6870);
xor U8490 (N_8490,N_7048,N_7166);
or U8491 (N_8491,N_5833,N_5032);
and U8492 (N_8492,N_6278,N_5435);
or U8493 (N_8493,N_5762,N_5951);
and U8494 (N_8494,N_5242,N_6183);
xnor U8495 (N_8495,N_5474,N_5628);
xor U8496 (N_8496,N_7342,N_6231);
xor U8497 (N_8497,N_5343,N_5942);
and U8498 (N_8498,N_6422,N_5971);
and U8499 (N_8499,N_5671,N_6826);
nand U8500 (N_8500,N_7495,N_5736);
nand U8501 (N_8501,N_6490,N_6644);
nand U8502 (N_8502,N_5806,N_5239);
nor U8503 (N_8503,N_6799,N_7498);
nor U8504 (N_8504,N_6913,N_6234);
nand U8505 (N_8505,N_6662,N_5856);
or U8506 (N_8506,N_5677,N_7165);
nand U8507 (N_8507,N_5503,N_5515);
and U8508 (N_8508,N_6367,N_5885);
and U8509 (N_8509,N_7392,N_7029);
or U8510 (N_8510,N_5106,N_5409);
nand U8511 (N_8511,N_5957,N_6569);
or U8512 (N_8512,N_7395,N_6262);
xnor U8513 (N_8513,N_5226,N_6504);
xnor U8514 (N_8514,N_5661,N_5364);
or U8515 (N_8515,N_5418,N_6726);
or U8516 (N_8516,N_6455,N_5629);
or U8517 (N_8517,N_7136,N_7369);
and U8518 (N_8518,N_7271,N_5684);
xor U8519 (N_8519,N_6056,N_7361);
nand U8520 (N_8520,N_5272,N_6310);
or U8521 (N_8521,N_5571,N_5928);
nand U8522 (N_8522,N_6646,N_5024);
and U8523 (N_8523,N_6850,N_6951);
nor U8524 (N_8524,N_5716,N_5540);
and U8525 (N_8525,N_5750,N_7186);
and U8526 (N_8526,N_5550,N_6606);
or U8527 (N_8527,N_7394,N_6783);
nand U8528 (N_8528,N_6842,N_6119);
nand U8529 (N_8529,N_6724,N_5471);
or U8530 (N_8530,N_6112,N_6083);
and U8531 (N_8531,N_7219,N_5698);
and U8532 (N_8532,N_7302,N_5960);
nor U8533 (N_8533,N_5128,N_6873);
nor U8534 (N_8534,N_6513,N_5208);
and U8535 (N_8535,N_5110,N_5267);
nand U8536 (N_8536,N_7170,N_6887);
nor U8537 (N_8537,N_5793,N_6519);
nand U8538 (N_8538,N_7109,N_5052);
nor U8539 (N_8539,N_7241,N_5256);
nor U8540 (N_8540,N_7141,N_5320);
or U8541 (N_8541,N_6725,N_7469);
or U8542 (N_8542,N_6964,N_7104);
nand U8543 (N_8543,N_5759,N_5339);
and U8544 (N_8544,N_5510,N_7134);
xor U8545 (N_8545,N_5248,N_6051);
nand U8546 (N_8546,N_5839,N_6053);
nand U8547 (N_8547,N_6450,N_6149);
and U8548 (N_8548,N_5486,N_6461);
or U8549 (N_8549,N_5499,N_6429);
or U8550 (N_8550,N_5504,N_5119);
nor U8551 (N_8551,N_6690,N_6171);
nor U8552 (N_8552,N_6324,N_5991);
and U8553 (N_8553,N_6933,N_6312);
or U8554 (N_8554,N_6269,N_5956);
nand U8555 (N_8555,N_5808,N_6989);
xnor U8556 (N_8556,N_5180,N_6087);
and U8557 (N_8557,N_5495,N_5602);
nand U8558 (N_8558,N_6830,N_5857);
nor U8559 (N_8559,N_5548,N_7244);
and U8560 (N_8560,N_7047,N_6667);
nand U8561 (N_8561,N_6163,N_5303);
nor U8562 (N_8562,N_5939,N_5538);
nor U8563 (N_8563,N_6795,N_6607);
nand U8564 (N_8564,N_5799,N_6260);
nor U8565 (N_8565,N_5872,N_7407);
xnor U8566 (N_8566,N_7074,N_5542);
or U8567 (N_8567,N_7282,N_6716);
nand U8568 (N_8568,N_6691,N_6510);
nand U8569 (N_8569,N_6174,N_5022);
nor U8570 (N_8570,N_6499,N_5194);
or U8571 (N_8571,N_5921,N_5441);
or U8572 (N_8572,N_7160,N_7156);
or U8573 (N_8573,N_5373,N_6405);
nor U8574 (N_8574,N_6089,N_5322);
or U8575 (N_8575,N_5395,N_7208);
or U8576 (N_8576,N_7288,N_5598);
or U8577 (N_8577,N_5426,N_5470);
and U8578 (N_8578,N_5468,N_5790);
nand U8579 (N_8579,N_5667,N_6073);
nor U8580 (N_8580,N_6003,N_7022);
nand U8581 (N_8581,N_5763,N_5906);
or U8582 (N_8582,N_6685,N_7323);
and U8583 (N_8583,N_5508,N_6516);
or U8584 (N_8584,N_7463,N_5570);
nand U8585 (N_8585,N_6894,N_7133);
or U8586 (N_8586,N_6259,N_6766);
xnor U8587 (N_8587,N_6780,N_6745);
and U8588 (N_8588,N_6889,N_5423);
nor U8589 (N_8589,N_6615,N_7252);
nand U8590 (N_8590,N_6593,N_6791);
or U8591 (N_8591,N_6772,N_5896);
nand U8592 (N_8592,N_5057,N_5221);
or U8593 (N_8593,N_6945,N_7127);
or U8594 (N_8594,N_6399,N_6944);
nand U8595 (N_8595,N_6984,N_7084);
or U8596 (N_8596,N_6190,N_5634);
and U8597 (N_8597,N_7235,N_7383);
or U8598 (N_8598,N_5385,N_5424);
or U8599 (N_8599,N_6123,N_5273);
xor U8600 (N_8600,N_7076,N_6907);
xnor U8601 (N_8601,N_6357,N_6268);
nor U8602 (N_8602,N_7163,N_5319);
and U8603 (N_8603,N_6013,N_7258);
nand U8604 (N_8604,N_5492,N_7327);
nand U8605 (N_8605,N_5611,N_5054);
nand U8606 (N_8606,N_7384,N_6474);
or U8607 (N_8607,N_5760,N_6077);
nand U8608 (N_8608,N_5900,N_6300);
and U8609 (N_8609,N_7196,N_5696);
nor U8610 (N_8610,N_6423,N_6334);
nand U8611 (N_8611,N_6353,N_5814);
xnor U8612 (N_8612,N_6668,N_7010);
nand U8613 (N_8613,N_7218,N_7402);
nand U8614 (N_8614,N_7334,N_6909);
nor U8615 (N_8615,N_6736,N_7056);
nand U8616 (N_8616,N_5215,N_5172);
nor U8617 (N_8617,N_7253,N_7052);
nor U8618 (N_8618,N_5544,N_6572);
or U8619 (N_8619,N_6082,N_6293);
nand U8620 (N_8620,N_6687,N_5767);
and U8621 (N_8621,N_6876,N_7499);
xnor U8622 (N_8622,N_5662,N_6152);
nand U8623 (N_8623,N_6845,N_5345);
nand U8624 (N_8624,N_7455,N_6222);
nand U8625 (N_8625,N_7349,N_5333);
nor U8626 (N_8626,N_6116,N_6126);
or U8627 (N_8627,N_5348,N_5962);
and U8628 (N_8628,N_6111,N_5047);
and U8629 (N_8629,N_5313,N_6350);
or U8630 (N_8630,N_5324,N_6605);
and U8631 (N_8631,N_5501,N_5440);
and U8632 (N_8632,N_7024,N_6728);
or U8633 (N_8633,N_5633,N_6442);
nor U8634 (N_8634,N_6610,N_5237);
or U8635 (N_8635,N_7411,N_5087);
nor U8636 (N_8636,N_7415,N_5038);
nor U8637 (N_8637,N_7320,N_7007);
xnor U8638 (N_8638,N_5664,N_7224);
or U8639 (N_8639,N_5400,N_6240);
and U8640 (N_8640,N_6741,N_6066);
nor U8641 (N_8641,N_6684,N_5777);
and U8642 (N_8642,N_5998,N_6292);
and U8643 (N_8643,N_7285,N_5490);
xor U8644 (N_8644,N_6958,N_5405);
xnor U8645 (N_8645,N_6311,N_5040);
nand U8646 (N_8646,N_7050,N_6634);
nand U8647 (N_8647,N_6542,N_7496);
nor U8648 (N_8648,N_6595,N_6081);
nor U8649 (N_8649,N_7430,N_6078);
nand U8650 (N_8650,N_7352,N_6194);
nand U8651 (N_8651,N_6118,N_5224);
xor U8652 (N_8652,N_5905,N_6468);
xor U8653 (N_8653,N_6860,N_6201);
nor U8654 (N_8654,N_6777,N_5649);
and U8655 (N_8655,N_5372,N_7105);
or U8656 (N_8656,N_6331,N_7130);
nand U8657 (N_8657,N_5524,N_7069);
and U8658 (N_8658,N_6700,N_6110);
nor U8659 (N_8659,N_7491,N_5130);
nand U8660 (N_8660,N_6925,N_6186);
nor U8661 (N_8661,N_6273,N_7475);
nor U8662 (N_8662,N_6885,N_5828);
xor U8663 (N_8663,N_6816,N_7097);
xnor U8664 (N_8664,N_7272,N_5679);
nand U8665 (N_8665,N_5536,N_5265);
nand U8666 (N_8666,N_5683,N_6096);
or U8667 (N_8667,N_6014,N_6865);
and U8668 (N_8668,N_7473,N_5009);
nor U8669 (N_8669,N_7414,N_5252);
and U8670 (N_8670,N_6626,N_5214);
nor U8671 (N_8671,N_5118,N_5092);
or U8672 (N_8672,N_7233,N_7474);
nor U8673 (N_8673,N_5410,N_6319);
nand U8674 (N_8674,N_6151,N_5967);
or U8675 (N_8675,N_7185,N_6241);
or U8676 (N_8676,N_7405,N_6541);
or U8677 (N_8677,N_5837,N_6501);
nor U8678 (N_8678,N_6321,N_5765);
nor U8679 (N_8679,N_5107,N_5174);
xnor U8680 (N_8680,N_7017,N_6613);
nand U8681 (N_8681,N_7310,N_5518);
and U8682 (N_8682,N_5060,N_5012);
or U8683 (N_8683,N_5724,N_6973);
and U8684 (N_8684,N_6469,N_5842);
nor U8685 (N_8685,N_6258,N_6484);
or U8686 (N_8686,N_6598,N_6801);
nand U8687 (N_8687,N_7482,N_7220);
and U8688 (N_8688,N_5528,N_6025);
or U8689 (N_8689,N_5549,N_7466);
nor U8690 (N_8690,N_7093,N_5148);
nand U8691 (N_8691,N_6496,N_7148);
and U8692 (N_8692,N_6244,N_5889);
nor U8693 (N_8693,N_7293,N_5437);
nand U8694 (N_8694,N_7442,N_6832);
and U8695 (N_8695,N_6370,N_7183);
nor U8696 (N_8696,N_5288,N_7326);
nor U8697 (N_8697,N_6427,N_6294);
nor U8698 (N_8698,N_6145,N_7014);
or U8699 (N_8699,N_6618,N_7243);
and U8700 (N_8700,N_5862,N_5541);
and U8701 (N_8701,N_5831,N_6696);
or U8702 (N_8702,N_7112,N_5803);
or U8703 (N_8703,N_5402,N_6846);
or U8704 (N_8704,N_5757,N_6451);
nand U8705 (N_8705,N_7297,N_5007);
nand U8706 (N_8706,N_6824,N_6121);
or U8707 (N_8707,N_6587,N_6227);
and U8708 (N_8708,N_6804,N_6929);
nand U8709 (N_8709,N_5427,N_5336);
xor U8710 (N_8710,N_5315,N_6202);
nand U8711 (N_8711,N_7128,N_5756);
nand U8712 (N_8712,N_5514,N_5852);
and U8713 (N_8713,N_5233,N_5165);
or U8714 (N_8714,N_5217,N_7477);
nand U8715 (N_8715,N_5298,N_6559);
nand U8716 (N_8716,N_5455,N_7432);
nor U8717 (N_8717,N_6574,N_5310);
and U8718 (N_8718,N_5871,N_6161);
nor U8719 (N_8719,N_6600,N_5630);
nand U8720 (N_8720,N_5114,N_5213);
nor U8721 (N_8721,N_6327,N_6315);
nor U8722 (N_8722,N_5718,N_7188);
nand U8723 (N_8723,N_7119,N_6551);
nand U8724 (N_8724,N_5813,N_5537);
nor U8725 (N_8725,N_6491,N_7489);
or U8726 (N_8726,N_6547,N_5576);
nand U8727 (N_8727,N_5144,N_7202);
nand U8728 (N_8728,N_6332,N_5113);
or U8729 (N_8729,N_5943,N_5545);
nor U8730 (N_8730,N_5457,N_6938);
or U8731 (N_8731,N_5836,N_5247);
nor U8732 (N_8732,N_7368,N_6284);
and U8733 (N_8733,N_7237,N_5123);
nand U8734 (N_8734,N_6517,N_5832);
nand U8735 (N_8735,N_5593,N_6277);
or U8736 (N_8736,N_6514,N_6660);
and U8737 (N_8737,N_6897,N_6354);
xnor U8738 (N_8738,N_7040,N_5484);
or U8739 (N_8739,N_5430,N_5566);
nor U8740 (N_8740,N_6416,N_5605);
nor U8741 (N_8741,N_7080,N_5425);
nand U8742 (N_8742,N_5023,N_5936);
or U8743 (N_8743,N_6458,N_6858);
xor U8744 (N_8744,N_5809,N_7426);
nand U8745 (N_8745,N_7039,N_7308);
and U8746 (N_8746,N_6625,N_5401);
nor U8747 (N_8747,N_7030,N_5747);
nand U8748 (N_8748,N_5462,N_6226);
and U8749 (N_8749,N_5181,N_6715);
nand U8750 (N_8750,N_5771,N_6536);
or U8751 (N_8751,N_5260,N_5353);
or U8752 (N_8752,N_5440,N_6623);
and U8753 (N_8753,N_6317,N_6003);
nor U8754 (N_8754,N_5969,N_6805);
nor U8755 (N_8755,N_7023,N_5957);
or U8756 (N_8756,N_6979,N_6351);
or U8757 (N_8757,N_6118,N_5965);
and U8758 (N_8758,N_5163,N_7255);
and U8759 (N_8759,N_5151,N_5455);
or U8760 (N_8760,N_7433,N_6836);
and U8761 (N_8761,N_5914,N_5633);
and U8762 (N_8762,N_6526,N_5420);
and U8763 (N_8763,N_5794,N_6545);
xor U8764 (N_8764,N_7113,N_5999);
nand U8765 (N_8765,N_6452,N_6503);
and U8766 (N_8766,N_6426,N_6220);
and U8767 (N_8767,N_7212,N_6256);
nor U8768 (N_8768,N_5402,N_5708);
nand U8769 (N_8769,N_5149,N_5345);
nor U8770 (N_8770,N_6503,N_7370);
and U8771 (N_8771,N_6942,N_5480);
nand U8772 (N_8772,N_5942,N_6999);
and U8773 (N_8773,N_6979,N_5135);
nand U8774 (N_8774,N_7106,N_6606);
and U8775 (N_8775,N_6846,N_7188);
and U8776 (N_8776,N_6448,N_5284);
xnor U8777 (N_8777,N_7062,N_6491);
or U8778 (N_8778,N_6036,N_5633);
xor U8779 (N_8779,N_5398,N_7128);
nor U8780 (N_8780,N_5336,N_6805);
nor U8781 (N_8781,N_5424,N_5526);
nand U8782 (N_8782,N_5673,N_6945);
or U8783 (N_8783,N_5437,N_6762);
nor U8784 (N_8784,N_5252,N_5501);
xor U8785 (N_8785,N_5883,N_6392);
xnor U8786 (N_8786,N_6612,N_5459);
nor U8787 (N_8787,N_6473,N_6552);
nor U8788 (N_8788,N_5211,N_6168);
and U8789 (N_8789,N_5427,N_6951);
and U8790 (N_8790,N_6687,N_7071);
nand U8791 (N_8791,N_6628,N_7079);
nand U8792 (N_8792,N_5076,N_5757);
nand U8793 (N_8793,N_5970,N_5496);
nor U8794 (N_8794,N_7217,N_6987);
or U8795 (N_8795,N_5209,N_5257);
nor U8796 (N_8796,N_7269,N_5242);
or U8797 (N_8797,N_7314,N_5227);
nand U8798 (N_8798,N_5391,N_6389);
nor U8799 (N_8799,N_5974,N_6548);
nor U8800 (N_8800,N_5765,N_6394);
or U8801 (N_8801,N_6157,N_5991);
nor U8802 (N_8802,N_6105,N_5657);
nor U8803 (N_8803,N_7345,N_5354);
nand U8804 (N_8804,N_6457,N_5643);
nor U8805 (N_8805,N_5120,N_5569);
xor U8806 (N_8806,N_6365,N_7493);
nand U8807 (N_8807,N_5200,N_7495);
nand U8808 (N_8808,N_6403,N_6140);
or U8809 (N_8809,N_5418,N_6741);
xnor U8810 (N_8810,N_6860,N_7228);
nor U8811 (N_8811,N_6614,N_6335);
nor U8812 (N_8812,N_5594,N_6700);
nand U8813 (N_8813,N_6212,N_6064);
or U8814 (N_8814,N_6328,N_5590);
nand U8815 (N_8815,N_5216,N_7220);
or U8816 (N_8816,N_5424,N_5134);
and U8817 (N_8817,N_7419,N_5031);
or U8818 (N_8818,N_5480,N_7308);
xor U8819 (N_8819,N_7128,N_6001);
or U8820 (N_8820,N_5975,N_5100);
or U8821 (N_8821,N_7281,N_6999);
or U8822 (N_8822,N_6496,N_6813);
or U8823 (N_8823,N_6560,N_7317);
nand U8824 (N_8824,N_7293,N_5917);
nor U8825 (N_8825,N_6624,N_5605);
nor U8826 (N_8826,N_5970,N_6630);
nand U8827 (N_8827,N_7012,N_5901);
nor U8828 (N_8828,N_6979,N_6492);
and U8829 (N_8829,N_7026,N_6159);
or U8830 (N_8830,N_5631,N_5501);
and U8831 (N_8831,N_6883,N_7059);
xnor U8832 (N_8832,N_5606,N_5583);
nand U8833 (N_8833,N_7430,N_7159);
nand U8834 (N_8834,N_7040,N_5305);
xnor U8835 (N_8835,N_6340,N_5718);
and U8836 (N_8836,N_5656,N_7029);
nor U8837 (N_8837,N_6881,N_7100);
nor U8838 (N_8838,N_6787,N_6277);
and U8839 (N_8839,N_5146,N_6862);
and U8840 (N_8840,N_5710,N_7168);
nor U8841 (N_8841,N_5778,N_6864);
xnor U8842 (N_8842,N_7392,N_6901);
nor U8843 (N_8843,N_6886,N_5450);
or U8844 (N_8844,N_6338,N_5109);
xnor U8845 (N_8845,N_5196,N_5594);
nor U8846 (N_8846,N_5240,N_7434);
and U8847 (N_8847,N_6219,N_5681);
nand U8848 (N_8848,N_5234,N_7169);
nor U8849 (N_8849,N_6579,N_6217);
nor U8850 (N_8850,N_6762,N_6283);
nor U8851 (N_8851,N_5468,N_5625);
and U8852 (N_8852,N_6598,N_6094);
and U8853 (N_8853,N_6086,N_5263);
or U8854 (N_8854,N_6916,N_7095);
and U8855 (N_8855,N_7487,N_7096);
xnor U8856 (N_8856,N_7483,N_5940);
and U8857 (N_8857,N_6747,N_6279);
and U8858 (N_8858,N_7418,N_6641);
nand U8859 (N_8859,N_5456,N_7055);
and U8860 (N_8860,N_7369,N_6092);
nor U8861 (N_8861,N_7004,N_6064);
nor U8862 (N_8862,N_5609,N_7463);
nand U8863 (N_8863,N_6057,N_7220);
nor U8864 (N_8864,N_6695,N_6130);
nor U8865 (N_8865,N_5158,N_7312);
nand U8866 (N_8866,N_5100,N_7085);
and U8867 (N_8867,N_5394,N_6332);
nor U8868 (N_8868,N_6232,N_5707);
nor U8869 (N_8869,N_6294,N_5067);
or U8870 (N_8870,N_5609,N_6523);
or U8871 (N_8871,N_7294,N_6085);
nor U8872 (N_8872,N_7321,N_6953);
and U8873 (N_8873,N_5007,N_5266);
or U8874 (N_8874,N_6738,N_6171);
nand U8875 (N_8875,N_6653,N_6763);
xor U8876 (N_8876,N_6377,N_7112);
or U8877 (N_8877,N_6549,N_6709);
and U8878 (N_8878,N_7196,N_6420);
and U8879 (N_8879,N_5774,N_6141);
nand U8880 (N_8880,N_5832,N_6776);
xor U8881 (N_8881,N_6341,N_5421);
or U8882 (N_8882,N_7388,N_7132);
nand U8883 (N_8883,N_7488,N_6192);
or U8884 (N_8884,N_7440,N_7039);
and U8885 (N_8885,N_7364,N_6814);
or U8886 (N_8886,N_6454,N_6088);
nand U8887 (N_8887,N_7119,N_6085);
nand U8888 (N_8888,N_5922,N_6260);
nor U8889 (N_8889,N_6337,N_6159);
or U8890 (N_8890,N_5522,N_7324);
nor U8891 (N_8891,N_5535,N_7300);
and U8892 (N_8892,N_5166,N_6897);
and U8893 (N_8893,N_6513,N_5191);
and U8894 (N_8894,N_7117,N_6826);
and U8895 (N_8895,N_7046,N_5716);
nand U8896 (N_8896,N_6814,N_7415);
xnor U8897 (N_8897,N_7479,N_6533);
or U8898 (N_8898,N_5320,N_7001);
and U8899 (N_8899,N_5031,N_5931);
or U8900 (N_8900,N_5546,N_6092);
xnor U8901 (N_8901,N_6711,N_5033);
nor U8902 (N_8902,N_5816,N_5181);
nor U8903 (N_8903,N_5811,N_7288);
nor U8904 (N_8904,N_5723,N_7022);
or U8905 (N_8905,N_5765,N_7297);
or U8906 (N_8906,N_5243,N_7401);
or U8907 (N_8907,N_5224,N_5147);
or U8908 (N_8908,N_5135,N_7003);
and U8909 (N_8909,N_7054,N_7457);
or U8910 (N_8910,N_6937,N_5083);
nand U8911 (N_8911,N_5591,N_7351);
xor U8912 (N_8912,N_6645,N_7288);
or U8913 (N_8913,N_5755,N_6263);
xnor U8914 (N_8914,N_6256,N_6704);
and U8915 (N_8915,N_7359,N_7104);
and U8916 (N_8916,N_7457,N_5782);
nand U8917 (N_8917,N_5338,N_5433);
nand U8918 (N_8918,N_7318,N_6867);
or U8919 (N_8919,N_7454,N_6508);
or U8920 (N_8920,N_5440,N_5003);
nor U8921 (N_8921,N_5793,N_6245);
nand U8922 (N_8922,N_5866,N_6221);
nor U8923 (N_8923,N_5959,N_6094);
nor U8924 (N_8924,N_5987,N_6966);
nor U8925 (N_8925,N_6642,N_7145);
xnor U8926 (N_8926,N_6684,N_5923);
xnor U8927 (N_8927,N_6049,N_6822);
nand U8928 (N_8928,N_5698,N_5672);
xnor U8929 (N_8929,N_5178,N_7238);
and U8930 (N_8930,N_5974,N_5285);
nand U8931 (N_8931,N_6812,N_5778);
nand U8932 (N_8932,N_5885,N_6489);
or U8933 (N_8933,N_7020,N_5090);
xor U8934 (N_8934,N_5115,N_7406);
xor U8935 (N_8935,N_5039,N_6480);
xnor U8936 (N_8936,N_7193,N_5778);
nand U8937 (N_8937,N_6555,N_7390);
nand U8938 (N_8938,N_5219,N_5150);
and U8939 (N_8939,N_5753,N_7235);
or U8940 (N_8940,N_5502,N_5271);
nor U8941 (N_8941,N_6899,N_5539);
nand U8942 (N_8942,N_7325,N_5177);
and U8943 (N_8943,N_5178,N_5465);
nand U8944 (N_8944,N_7371,N_7022);
nor U8945 (N_8945,N_5781,N_6382);
nand U8946 (N_8946,N_5912,N_6980);
or U8947 (N_8947,N_5973,N_5523);
nand U8948 (N_8948,N_6347,N_5241);
nor U8949 (N_8949,N_6294,N_5819);
or U8950 (N_8950,N_7288,N_5648);
or U8951 (N_8951,N_6217,N_7328);
nand U8952 (N_8952,N_6420,N_5088);
nor U8953 (N_8953,N_5706,N_7325);
nor U8954 (N_8954,N_5604,N_7429);
or U8955 (N_8955,N_5320,N_5846);
nor U8956 (N_8956,N_7217,N_6684);
nor U8957 (N_8957,N_6812,N_6124);
or U8958 (N_8958,N_6642,N_5171);
and U8959 (N_8959,N_6289,N_7169);
and U8960 (N_8960,N_7167,N_6231);
or U8961 (N_8961,N_5387,N_6005);
nor U8962 (N_8962,N_5555,N_6390);
or U8963 (N_8963,N_5816,N_6240);
nor U8964 (N_8964,N_6830,N_6267);
and U8965 (N_8965,N_5394,N_5199);
or U8966 (N_8966,N_6182,N_6014);
nand U8967 (N_8967,N_7449,N_6404);
nor U8968 (N_8968,N_6908,N_5037);
nand U8969 (N_8969,N_7419,N_6760);
or U8970 (N_8970,N_5103,N_6871);
or U8971 (N_8971,N_5188,N_7379);
nand U8972 (N_8972,N_5632,N_5148);
and U8973 (N_8973,N_6663,N_7493);
and U8974 (N_8974,N_7402,N_6064);
and U8975 (N_8975,N_5780,N_5373);
nor U8976 (N_8976,N_6377,N_7201);
nor U8977 (N_8977,N_5840,N_5757);
nor U8978 (N_8978,N_5283,N_7360);
and U8979 (N_8979,N_6733,N_7405);
nor U8980 (N_8980,N_6988,N_6945);
nor U8981 (N_8981,N_7498,N_6955);
and U8982 (N_8982,N_5026,N_6795);
nand U8983 (N_8983,N_5510,N_7267);
nand U8984 (N_8984,N_6045,N_6586);
nor U8985 (N_8985,N_6772,N_7092);
nor U8986 (N_8986,N_5670,N_6954);
and U8987 (N_8987,N_6458,N_7227);
nor U8988 (N_8988,N_7427,N_6685);
and U8989 (N_8989,N_7222,N_6523);
or U8990 (N_8990,N_6192,N_5032);
and U8991 (N_8991,N_6076,N_5436);
or U8992 (N_8992,N_5047,N_7176);
and U8993 (N_8993,N_6438,N_5322);
or U8994 (N_8994,N_5461,N_6538);
and U8995 (N_8995,N_6837,N_5146);
nand U8996 (N_8996,N_5976,N_5837);
xnor U8997 (N_8997,N_7217,N_7221);
xnor U8998 (N_8998,N_6486,N_5780);
or U8999 (N_8999,N_5795,N_5305);
nand U9000 (N_9000,N_6018,N_5553);
nand U9001 (N_9001,N_7113,N_6117);
xor U9002 (N_9002,N_5740,N_6959);
or U9003 (N_9003,N_6381,N_6071);
nor U9004 (N_9004,N_5608,N_5877);
nor U9005 (N_9005,N_7109,N_7128);
or U9006 (N_9006,N_6735,N_7306);
nor U9007 (N_9007,N_6197,N_5103);
or U9008 (N_9008,N_7203,N_7422);
xnor U9009 (N_9009,N_5805,N_6566);
and U9010 (N_9010,N_6895,N_7294);
nor U9011 (N_9011,N_5160,N_6888);
xnor U9012 (N_9012,N_7219,N_5819);
or U9013 (N_9013,N_7168,N_5764);
nor U9014 (N_9014,N_7086,N_5583);
and U9015 (N_9015,N_6049,N_5077);
or U9016 (N_9016,N_6609,N_5189);
nor U9017 (N_9017,N_5013,N_6265);
nor U9018 (N_9018,N_5198,N_6187);
and U9019 (N_9019,N_7233,N_6971);
and U9020 (N_9020,N_6473,N_6067);
nand U9021 (N_9021,N_7375,N_6837);
or U9022 (N_9022,N_6785,N_6019);
and U9023 (N_9023,N_6922,N_5977);
nand U9024 (N_9024,N_6962,N_5952);
nand U9025 (N_9025,N_6555,N_5798);
or U9026 (N_9026,N_7109,N_6048);
xor U9027 (N_9027,N_5698,N_5563);
or U9028 (N_9028,N_7056,N_5521);
nor U9029 (N_9029,N_6827,N_5570);
nand U9030 (N_9030,N_5425,N_7064);
nor U9031 (N_9031,N_5260,N_5110);
nor U9032 (N_9032,N_6659,N_7486);
nor U9033 (N_9033,N_6683,N_6396);
nand U9034 (N_9034,N_6317,N_7169);
nand U9035 (N_9035,N_7224,N_7321);
nor U9036 (N_9036,N_7344,N_5699);
and U9037 (N_9037,N_7329,N_5834);
or U9038 (N_9038,N_6048,N_5491);
nand U9039 (N_9039,N_5067,N_5398);
and U9040 (N_9040,N_7458,N_5623);
nor U9041 (N_9041,N_6383,N_5128);
nand U9042 (N_9042,N_6815,N_5754);
xnor U9043 (N_9043,N_6349,N_6119);
xor U9044 (N_9044,N_5098,N_6847);
xnor U9045 (N_9045,N_6549,N_5029);
and U9046 (N_9046,N_5719,N_5861);
nand U9047 (N_9047,N_5294,N_5041);
nand U9048 (N_9048,N_7215,N_5210);
nor U9049 (N_9049,N_7416,N_6839);
nor U9050 (N_9050,N_7208,N_5426);
nor U9051 (N_9051,N_5942,N_6437);
nand U9052 (N_9052,N_5290,N_6445);
nand U9053 (N_9053,N_5554,N_5697);
or U9054 (N_9054,N_6816,N_6476);
or U9055 (N_9055,N_6243,N_6174);
xor U9056 (N_9056,N_7114,N_7054);
nand U9057 (N_9057,N_5696,N_6024);
nand U9058 (N_9058,N_5781,N_6548);
and U9059 (N_9059,N_5165,N_5700);
nand U9060 (N_9060,N_6433,N_6988);
or U9061 (N_9061,N_6948,N_5213);
and U9062 (N_9062,N_5460,N_6041);
nor U9063 (N_9063,N_6097,N_5767);
or U9064 (N_9064,N_7136,N_6708);
nor U9065 (N_9065,N_5727,N_5458);
xnor U9066 (N_9066,N_6262,N_5377);
xor U9067 (N_9067,N_5619,N_5735);
and U9068 (N_9068,N_6487,N_5997);
or U9069 (N_9069,N_5679,N_6242);
or U9070 (N_9070,N_5812,N_5151);
or U9071 (N_9071,N_6791,N_6656);
nor U9072 (N_9072,N_5291,N_5476);
nand U9073 (N_9073,N_7163,N_5842);
nor U9074 (N_9074,N_5692,N_5657);
nor U9075 (N_9075,N_6590,N_7150);
nand U9076 (N_9076,N_5534,N_6424);
and U9077 (N_9077,N_5912,N_5139);
nand U9078 (N_9078,N_5017,N_7239);
nand U9079 (N_9079,N_5317,N_7347);
or U9080 (N_9080,N_5200,N_6213);
and U9081 (N_9081,N_5656,N_5756);
and U9082 (N_9082,N_6294,N_5968);
nand U9083 (N_9083,N_7122,N_6086);
nor U9084 (N_9084,N_5845,N_7210);
or U9085 (N_9085,N_5973,N_5314);
and U9086 (N_9086,N_7016,N_5669);
and U9087 (N_9087,N_6204,N_7482);
nor U9088 (N_9088,N_6281,N_7350);
or U9089 (N_9089,N_5624,N_7460);
nand U9090 (N_9090,N_6210,N_5336);
nor U9091 (N_9091,N_5327,N_5293);
or U9092 (N_9092,N_5099,N_5695);
nor U9093 (N_9093,N_5128,N_6929);
nor U9094 (N_9094,N_7067,N_5994);
nor U9095 (N_9095,N_6490,N_6201);
nand U9096 (N_9096,N_5074,N_7252);
or U9097 (N_9097,N_6924,N_5173);
xor U9098 (N_9098,N_6729,N_6831);
nand U9099 (N_9099,N_5647,N_5631);
nand U9100 (N_9100,N_7058,N_6252);
nand U9101 (N_9101,N_6641,N_6732);
or U9102 (N_9102,N_6571,N_6647);
and U9103 (N_9103,N_7356,N_6201);
nand U9104 (N_9104,N_5506,N_5288);
or U9105 (N_9105,N_6836,N_7361);
and U9106 (N_9106,N_7321,N_6159);
xor U9107 (N_9107,N_5107,N_6620);
or U9108 (N_9108,N_5029,N_6847);
and U9109 (N_9109,N_6099,N_7084);
nor U9110 (N_9110,N_7273,N_7076);
and U9111 (N_9111,N_6381,N_5304);
and U9112 (N_9112,N_6160,N_5722);
or U9113 (N_9113,N_5405,N_5557);
or U9114 (N_9114,N_5516,N_6177);
nor U9115 (N_9115,N_5091,N_5804);
and U9116 (N_9116,N_7480,N_5330);
nand U9117 (N_9117,N_7207,N_6328);
nand U9118 (N_9118,N_6028,N_7130);
nand U9119 (N_9119,N_6333,N_5202);
nand U9120 (N_9120,N_7206,N_7144);
and U9121 (N_9121,N_5999,N_6509);
nand U9122 (N_9122,N_7460,N_6017);
or U9123 (N_9123,N_5009,N_6170);
nand U9124 (N_9124,N_6310,N_6985);
and U9125 (N_9125,N_7227,N_5249);
or U9126 (N_9126,N_7188,N_6014);
nor U9127 (N_9127,N_5235,N_5443);
or U9128 (N_9128,N_5242,N_5403);
and U9129 (N_9129,N_5790,N_7400);
nand U9130 (N_9130,N_7372,N_6043);
nand U9131 (N_9131,N_5147,N_5530);
nand U9132 (N_9132,N_6652,N_6689);
or U9133 (N_9133,N_6549,N_6988);
nand U9134 (N_9134,N_6354,N_5140);
nand U9135 (N_9135,N_6095,N_6164);
and U9136 (N_9136,N_6760,N_7210);
nor U9137 (N_9137,N_6508,N_7253);
or U9138 (N_9138,N_7328,N_6178);
nand U9139 (N_9139,N_5514,N_6334);
nor U9140 (N_9140,N_5182,N_5646);
or U9141 (N_9141,N_5089,N_5616);
or U9142 (N_9142,N_5450,N_5757);
and U9143 (N_9143,N_5963,N_6976);
nor U9144 (N_9144,N_6995,N_6930);
nor U9145 (N_9145,N_5757,N_6134);
nor U9146 (N_9146,N_7438,N_6965);
nand U9147 (N_9147,N_7124,N_5644);
nor U9148 (N_9148,N_5575,N_5110);
nor U9149 (N_9149,N_5333,N_6003);
xor U9150 (N_9150,N_5071,N_6473);
and U9151 (N_9151,N_5971,N_6739);
nor U9152 (N_9152,N_6245,N_5016);
or U9153 (N_9153,N_5430,N_5434);
and U9154 (N_9154,N_5113,N_6872);
xnor U9155 (N_9155,N_6412,N_6305);
nor U9156 (N_9156,N_5459,N_6583);
nand U9157 (N_9157,N_6265,N_5249);
nor U9158 (N_9158,N_6078,N_6884);
nand U9159 (N_9159,N_5047,N_7180);
and U9160 (N_9160,N_6126,N_7165);
nor U9161 (N_9161,N_5557,N_6284);
nor U9162 (N_9162,N_6004,N_6565);
and U9163 (N_9163,N_5181,N_5787);
nor U9164 (N_9164,N_7425,N_6825);
and U9165 (N_9165,N_6215,N_6433);
nor U9166 (N_9166,N_5103,N_5542);
nor U9167 (N_9167,N_7492,N_5949);
nor U9168 (N_9168,N_7268,N_6976);
or U9169 (N_9169,N_6309,N_7363);
nor U9170 (N_9170,N_5440,N_6042);
nor U9171 (N_9171,N_6704,N_7010);
or U9172 (N_9172,N_6096,N_5826);
and U9173 (N_9173,N_6791,N_5441);
and U9174 (N_9174,N_5435,N_5765);
and U9175 (N_9175,N_6323,N_6267);
and U9176 (N_9176,N_6118,N_7041);
nand U9177 (N_9177,N_6528,N_5144);
or U9178 (N_9178,N_6620,N_6996);
nand U9179 (N_9179,N_7090,N_5745);
or U9180 (N_9180,N_6898,N_5602);
nand U9181 (N_9181,N_6805,N_6518);
nand U9182 (N_9182,N_5627,N_5599);
nor U9183 (N_9183,N_7498,N_5910);
nand U9184 (N_9184,N_7418,N_6247);
nor U9185 (N_9185,N_6131,N_6159);
nor U9186 (N_9186,N_6511,N_6187);
nand U9187 (N_9187,N_6295,N_6224);
xnor U9188 (N_9188,N_6024,N_7389);
nand U9189 (N_9189,N_5578,N_7232);
or U9190 (N_9190,N_7000,N_5611);
nand U9191 (N_9191,N_5569,N_6662);
or U9192 (N_9192,N_5290,N_5142);
or U9193 (N_9193,N_5445,N_5240);
and U9194 (N_9194,N_6656,N_6835);
nand U9195 (N_9195,N_7138,N_5031);
and U9196 (N_9196,N_6502,N_5279);
and U9197 (N_9197,N_5134,N_6027);
or U9198 (N_9198,N_5147,N_6188);
nand U9199 (N_9199,N_6600,N_6809);
xor U9200 (N_9200,N_5288,N_5247);
nand U9201 (N_9201,N_6356,N_6418);
nand U9202 (N_9202,N_5843,N_5698);
or U9203 (N_9203,N_6773,N_6906);
xor U9204 (N_9204,N_5230,N_5713);
and U9205 (N_9205,N_6113,N_6963);
xnor U9206 (N_9206,N_5111,N_6496);
nand U9207 (N_9207,N_5123,N_6264);
or U9208 (N_9208,N_7123,N_6307);
or U9209 (N_9209,N_6498,N_5994);
nand U9210 (N_9210,N_7199,N_6756);
nor U9211 (N_9211,N_5193,N_7267);
xor U9212 (N_9212,N_7209,N_6697);
and U9213 (N_9213,N_5487,N_6818);
nand U9214 (N_9214,N_6406,N_6135);
nor U9215 (N_9215,N_6392,N_6607);
nand U9216 (N_9216,N_5627,N_5788);
and U9217 (N_9217,N_6803,N_5971);
or U9218 (N_9218,N_6103,N_5446);
and U9219 (N_9219,N_7178,N_6777);
nor U9220 (N_9220,N_5187,N_6240);
xnor U9221 (N_9221,N_6214,N_5470);
nor U9222 (N_9222,N_5219,N_5547);
and U9223 (N_9223,N_5144,N_5145);
nor U9224 (N_9224,N_6713,N_6513);
or U9225 (N_9225,N_7099,N_6114);
nor U9226 (N_9226,N_5491,N_5092);
xnor U9227 (N_9227,N_5206,N_5980);
or U9228 (N_9228,N_6471,N_5772);
and U9229 (N_9229,N_6822,N_6219);
nor U9230 (N_9230,N_7484,N_6316);
and U9231 (N_9231,N_5092,N_5157);
or U9232 (N_9232,N_6060,N_5664);
xnor U9233 (N_9233,N_5464,N_5395);
nor U9234 (N_9234,N_7337,N_7226);
nand U9235 (N_9235,N_5184,N_6504);
nand U9236 (N_9236,N_6225,N_5338);
xnor U9237 (N_9237,N_5126,N_5452);
or U9238 (N_9238,N_5349,N_5453);
nor U9239 (N_9239,N_5730,N_6808);
nor U9240 (N_9240,N_5034,N_7430);
xnor U9241 (N_9241,N_5020,N_5497);
and U9242 (N_9242,N_6059,N_6873);
or U9243 (N_9243,N_6979,N_6163);
or U9244 (N_9244,N_5705,N_5847);
nor U9245 (N_9245,N_6687,N_5064);
nand U9246 (N_9246,N_7226,N_5436);
and U9247 (N_9247,N_5140,N_5194);
or U9248 (N_9248,N_6211,N_5367);
nor U9249 (N_9249,N_6717,N_6169);
nand U9250 (N_9250,N_5537,N_6713);
or U9251 (N_9251,N_6201,N_7199);
nand U9252 (N_9252,N_5011,N_5009);
xor U9253 (N_9253,N_6332,N_6937);
nand U9254 (N_9254,N_7494,N_6127);
nor U9255 (N_9255,N_6814,N_6362);
nand U9256 (N_9256,N_6991,N_6493);
xor U9257 (N_9257,N_5716,N_6443);
xor U9258 (N_9258,N_6911,N_5330);
nor U9259 (N_9259,N_6451,N_5382);
nand U9260 (N_9260,N_7037,N_6135);
nor U9261 (N_9261,N_6414,N_6371);
xnor U9262 (N_9262,N_6505,N_7135);
nor U9263 (N_9263,N_7161,N_6487);
xnor U9264 (N_9264,N_6248,N_6307);
or U9265 (N_9265,N_7486,N_5196);
nor U9266 (N_9266,N_6887,N_5790);
nor U9267 (N_9267,N_7248,N_6782);
nand U9268 (N_9268,N_7163,N_7046);
or U9269 (N_9269,N_6628,N_5586);
nor U9270 (N_9270,N_5209,N_7284);
or U9271 (N_9271,N_5492,N_6305);
or U9272 (N_9272,N_6602,N_5669);
or U9273 (N_9273,N_5138,N_6735);
or U9274 (N_9274,N_6437,N_5368);
or U9275 (N_9275,N_7232,N_6672);
nand U9276 (N_9276,N_5241,N_6679);
nor U9277 (N_9277,N_5541,N_5783);
nor U9278 (N_9278,N_6598,N_5745);
and U9279 (N_9279,N_5566,N_5735);
xnor U9280 (N_9280,N_7165,N_6381);
nor U9281 (N_9281,N_5727,N_6742);
and U9282 (N_9282,N_5752,N_6373);
and U9283 (N_9283,N_5608,N_5807);
nand U9284 (N_9284,N_6835,N_5234);
nand U9285 (N_9285,N_7306,N_6554);
or U9286 (N_9286,N_6880,N_5983);
nor U9287 (N_9287,N_6998,N_5036);
nand U9288 (N_9288,N_5620,N_6860);
or U9289 (N_9289,N_6220,N_5280);
xnor U9290 (N_9290,N_7366,N_5332);
and U9291 (N_9291,N_6832,N_5667);
nor U9292 (N_9292,N_5031,N_7133);
nand U9293 (N_9293,N_5719,N_5587);
xor U9294 (N_9294,N_5933,N_7151);
xnor U9295 (N_9295,N_6093,N_6836);
nor U9296 (N_9296,N_6865,N_5986);
nand U9297 (N_9297,N_6322,N_6533);
and U9298 (N_9298,N_5528,N_5905);
nor U9299 (N_9299,N_5463,N_6120);
xnor U9300 (N_9300,N_6402,N_6561);
nor U9301 (N_9301,N_5285,N_5429);
nor U9302 (N_9302,N_6274,N_5788);
nand U9303 (N_9303,N_5829,N_6419);
nand U9304 (N_9304,N_6057,N_5023);
xor U9305 (N_9305,N_5658,N_5260);
nor U9306 (N_9306,N_5051,N_6909);
or U9307 (N_9307,N_6044,N_6589);
and U9308 (N_9308,N_7183,N_5711);
and U9309 (N_9309,N_6860,N_7185);
nor U9310 (N_9310,N_5863,N_6741);
nor U9311 (N_9311,N_6685,N_6030);
or U9312 (N_9312,N_5715,N_6089);
or U9313 (N_9313,N_6869,N_5724);
or U9314 (N_9314,N_6100,N_7239);
nand U9315 (N_9315,N_6853,N_7167);
nand U9316 (N_9316,N_5323,N_6544);
or U9317 (N_9317,N_5733,N_6989);
and U9318 (N_9318,N_5597,N_5294);
xnor U9319 (N_9319,N_5425,N_6869);
and U9320 (N_9320,N_5886,N_5765);
nor U9321 (N_9321,N_5648,N_5013);
and U9322 (N_9322,N_6613,N_5809);
nor U9323 (N_9323,N_5908,N_5827);
or U9324 (N_9324,N_5264,N_7182);
or U9325 (N_9325,N_6307,N_6431);
nor U9326 (N_9326,N_5914,N_6193);
xor U9327 (N_9327,N_5544,N_5115);
or U9328 (N_9328,N_6898,N_7219);
or U9329 (N_9329,N_5600,N_5038);
xor U9330 (N_9330,N_5577,N_6397);
or U9331 (N_9331,N_5019,N_5135);
and U9332 (N_9332,N_7232,N_6976);
and U9333 (N_9333,N_7002,N_6041);
nand U9334 (N_9334,N_6152,N_6930);
nand U9335 (N_9335,N_6167,N_7227);
and U9336 (N_9336,N_6309,N_7330);
or U9337 (N_9337,N_5431,N_5365);
and U9338 (N_9338,N_6711,N_5391);
nand U9339 (N_9339,N_7140,N_6785);
nand U9340 (N_9340,N_6277,N_6770);
or U9341 (N_9341,N_5886,N_6891);
and U9342 (N_9342,N_7392,N_6150);
nor U9343 (N_9343,N_6597,N_6806);
xnor U9344 (N_9344,N_5869,N_6661);
or U9345 (N_9345,N_6115,N_5867);
xnor U9346 (N_9346,N_6607,N_6126);
or U9347 (N_9347,N_5517,N_5973);
or U9348 (N_9348,N_6003,N_5337);
or U9349 (N_9349,N_5572,N_5277);
nand U9350 (N_9350,N_6107,N_5774);
and U9351 (N_9351,N_6590,N_5471);
and U9352 (N_9352,N_7070,N_7428);
nand U9353 (N_9353,N_6813,N_5187);
and U9354 (N_9354,N_5979,N_7195);
and U9355 (N_9355,N_6833,N_5659);
nor U9356 (N_9356,N_7164,N_5803);
nand U9357 (N_9357,N_6918,N_6797);
nand U9358 (N_9358,N_6046,N_6796);
nand U9359 (N_9359,N_6234,N_6996);
nand U9360 (N_9360,N_5599,N_6450);
or U9361 (N_9361,N_6876,N_5471);
and U9362 (N_9362,N_5030,N_5260);
nand U9363 (N_9363,N_7010,N_5407);
xor U9364 (N_9364,N_7395,N_5865);
and U9365 (N_9365,N_5953,N_5362);
and U9366 (N_9366,N_5171,N_6864);
xor U9367 (N_9367,N_6717,N_6843);
and U9368 (N_9368,N_5009,N_7296);
or U9369 (N_9369,N_6359,N_6039);
nor U9370 (N_9370,N_5099,N_5711);
or U9371 (N_9371,N_7474,N_5649);
or U9372 (N_9372,N_6154,N_5337);
xnor U9373 (N_9373,N_5852,N_7434);
and U9374 (N_9374,N_6679,N_5670);
or U9375 (N_9375,N_6526,N_5547);
or U9376 (N_9376,N_6005,N_5827);
and U9377 (N_9377,N_7245,N_6607);
nand U9378 (N_9378,N_5074,N_5176);
or U9379 (N_9379,N_7409,N_5713);
nand U9380 (N_9380,N_6404,N_5211);
nand U9381 (N_9381,N_7230,N_7156);
nand U9382 (N_9382,N_6028,N_5386);
nor U9383 (N_9383,N_5788,N_6884);
nand U9384 (N_9384,N_6589,N_5686);
xnor U9385 (N_9385,N_5634,N_6375);
nor U9386 (N_9386,N_7071,N_7334);
and U9387 (N_9387,N_5400,N_5083);
or U9388 (N_9388,N_5473,N_7064);
nand U9389 (N_9389,N_5734,N_6788);
or U9390 (N_9390,N_5330,N_5883);
xnor U9391 (N_9391,N_6047,N_5034);
and U9392 (N_9392,N_5867,N_6527);
and U9393 (N_9393,N_5850,N_6828);
nand U9394 (N_9394,N_5514,N_7455);
and U9395 (N_9395,N_6927,N_6152);
or U9396 (N_9396,N_6204,N_7237);
nand U9397 (N_9397,N_5439,N_5745);
and U9398 (N_9398,N_5750,N_6475);
nor U9399 (N_9399,N_5451,N_6667);
and U9400 (N_9400,N_5036,N_5137);
nand U9401 (N_9401,N_5533,N_5940);
nand U9402 (N_9402,N_5782,N_7028);
and U9403 (N_9403,N_7411,N_5475);
or U9404 (N_9404,N_5587,N_6352);
nand U9405 (N_9405,N_7311,N_6361);
nand U9406 (N_9406,N_6792,N_5664);
nand U9407 (N_9407,N_6727,N_5286);
nand U9408 (N_9408,N_5775,N_5052);
or U9409 (N_9409,N_5398,N_7043);
and U9410 (N_9410,N_6474,N_5159);
nor U9411 (N_9411,N_6113,N_6502);
xnor U9412 (N_9412,N_6277,N_5080);
xnor U9413 (N_9413,N_5565,N_7142);
and U9414 (N_9414,N_5152,N_5956);
or U9415 (N_9415,N_7436,N_7236);
nand U9416 (N_9416,N_7448,N_5448);
nand U9417 (N_9417,N_6267,N_6101);
and U9418 (N_9418,N_7278,N_6879);
and U9419 (N_9419,N_5778,N_7194);
and U9420 (N_9420,N_7122,N_7477);
or U9421 (N_9421,N_6784,N_7261);
and U9422 (N_9422,N_5618,N_6220);
or U9423 (N_9423,N_7412,N_6095);
nand U9424 (N_9424,N_5054,N_6949);
nor U9425 (N_9425,N_7032,N_5952);
nand U9426 (N_9426,N_5634,N_6438);
and U9427 (N_9427,N_5776,N_5644);
nand U9428 (N_9428,N_5140,N_6546);
and U9429 (N_9429,N_6411,N_7385);
or U9430 (N_9430,N_6062,N_5536);
nor U9431 (N_9431,N_5351,N_6390);
or U9432 (N_9432,N_7250,N_6928);
xnor U9433 (N_9433,N_5504,N_6750);
nor U9434 (N_9434,N_6018,N_6119);
xor U9435 (N_9435,N_5815,N_7330);
xor U9436 (N_9436,N_5997,N_7236);
xnor U9437 (N_9437,N_6411,N_6217);
and U9438 (N_9438,N_7040,N_6490);
and U9439 (N_9439,N_6029,N_7474);
or U9440 (N_9440,N_6175,N_7245);
nor U9441 (N_9441,N_5038,N_6883);
nand U9442 (N_9442,N_5353,N_6410);
and U9443 (N_9443,N_5658,N_6088);
nor U9444 (N_9444,N_5800,N_6895);
and U9445 (N_9445,N_6096,N_5546);
nand U9446 (N_9446,N_7373,N_6449);
xnor U9447 (N_9447,N_6079,N_5556);
nand U9448 (N_9448,N_5355,N_7319);
nand U9449 (N_9449,N_6804,N_6316);
and U9450 (N_9450,N_5928,N_6740);
and U9451 (N_9451,N_5376,N_7347);
nor U9452 (N_9452,N_5785,N_5829);
nand U9453 (N_9453,N_6079,N_6462);
and U9454 (N_9454,N_5559,N_5699);
and U9455 (N_9455,N_6847,N_5916);
nand U9456 (N_9456,N_6221,N_5128);
nor U9457 (N_9457,N_5362,N_7028);
xnor U9458 (N_9458,N_5190,N_6243);
nand U9459 (N_9459,N_6567,N_7481);
and U9460 (N_9460,N_6989,N_5913);
nand U9461 (N_9461,N_5501,N_5430);
and U9462 (N_9462,N_7166,N_6131);
or U9463 (N_9463,N_5234,N_7347);
and U9464 (N_9464,N_5996,N_6227);
xor U9465 (N_9465,N_5378,N_6731);
and U9466 (N_9466,N_5202,N_6446);
and U9467 (N_9467,N_6270,N_6594);
or U9468 (N_9468,N_7271,N_6734);
and U9469 (N_9469,N_5083,N_6710);
nor U9470 (N_9470,N_6721,N_5760);
nor U9471 (N_9471,N_6211,N_7148);
nor U9472 (N_9472,N_5001,N_5608);
or U9473 (N_9473,N_6824,N_5653);
and U9474 (N_9474,N_6699,N_5298);
or U9475 (N_9475,N_7049,N_7489);
and U9476 (N_9476,N_5606,N_7368);
nand U9477 (N_9477,N_7048,N_5231);
nor U9478 (N_9478,N_5343,N_5954);
or U9479 (N_9479,N_6144,N_6636);
nand U9480 (N_9480,N_5255,N_6386);
and U9481 (N_9481,N_7200,N_7226);
nand U9482 (N_9482,N_6975,N_6594);
and U9483 (N_9483,N_5570,N_6820);
and U9484 (N_9484,N_5602,N_7348);
nor U9485 (N_9485,N_6979,N_6615);
nor U9486 (N_9486,N_5290,N_6003);
or U9487 (N_9487,N_6579,N_5811);
and U9488 (N_9488,N_7116,N_6492);
xnor U9489 (N_9489,N_7141,N_5842);
nor U9490 (N_9490,N_6049,N_6607);
and U9491 (N_9491,N_6035,N_6932);
nand U9492 (N_9492,N_6408,N_5154);
nor U9493 (N_9493,N_5268,N_6230);
and U9494 (N_9494,N_7253,N_5284);
xnor U9495 (N_9495,N_6125,N_6391);
nand U9496 (N_9496,N_5819,N_5980);
nand U9497 (N_9497,N_5470,N_5556);
nand U9498 (N_9498,N_7233,N_7080);
and U9499 (N_9499,N_7143,N_6603);
nor U9500 (N_9500,N_5967,N_6546);
nand U9501 (N_9501,N_6773,N_5644);
or U9502 (N_9502,N_5614,N_7196);
nor U9503 (N_9503,N_5624,N_5256);
or U9504 (N_9504,N_6103,N_6962);
or U9505 (N_9505,N_5723,N_6713);
or U9506 (N_9506,N_5578,N_7023);
xor U9507 (N_9507,N_5385,N_5140);
nand U9508 (N_9508,N_5141,N_5831);
nor U9509 (N_9509,N_6094,N_5526);
xnor U9510 (N_9510,N_7169,N_5563);
or U9511 (N_9511,N_5664,N_5965);
or U9512 (N_9512,N_6750,N_7157);
nor U9513 (N_9513,N_6266,N_6158);
nand U9514 (N_9514,N_6917,N_6400);
or U9515 (N_9515,N_6613,N_5752);
nand U9516 (N_9516,N_6982,N_5548);
nor U9517 (N_9517,N_7452,N_6212);
xor U9518 (N_9518,N_6034,N_7170);
or U9519 (N_9519,N_5180,N_5031);
or U9520 (N_9520,N_6147,N_5064);
and U9521 (N_9521,N_6666,N_6814);
nand U9522 (N_9522,N_6505,N_5315);
nand U9523 (N_9523,N_7490,N_6464);
or U9524 (N_9524,N_5091,N_7376);
or U9525 (N_9525,N_6052,N_6106);
and U9526 (N_9526,N_5503,N_5905);
xor U9527 (N_9527,N_6835,N_5376);
xor U9528 (N_9528,N_6856,N_7019);
nand U9529 (N_9529,N_6945,N_5046);
and U9530 (N_9530,N_5144,N_5025);
and U9531 (N_9531,N_7219,N_6518);
or U9532 (N_9532,N_6034,N_5150);
or U9533 (N_9533,N_5087,N_7046);
or U9534 (N_9534,N_5945,N_6355);
or U9535 (N_9535,N_7293,N_5466);
and U9536 (N_9536,N_6383,N_6349);
xnor U9537 (N_9537,N_6986,N_6493);
xor U9538 (N_9538,N_6650,N_6453);
or U9539 (N_9539,N_5446,N_7371);
nor U9540 (N_9540,N_5467,N_7357);
nor U9541 (N_9541,N_5723,N_6583);
nand U9542 (N_9542,N_6118,N_5556);
nor U9543 (N_9543,N_5037,N_5466);
nand U9544 (N_9544,N_5857,N_7046);
nand U9545 (N_9545,N_6301,N_5539);
and U9546 (N_9546,N_6003,N_5394);
and U9547 (N_9547,N_5793,N_5826);
nand U9548 (N_9548,N_5718,N_6551);
or U9549 (N_9549,N_7190,N_6735);
nand U9550 (N_9550,N_6700,N_7049);
nand U9551 (N_9551,N_5681,N_6929);
and U9552 (N_9552,N_6392,N_6263);
and U9553 (N_9553,N_5986,N_6898);
or U9554 (N_9554,N_7342,N_6499);
or U9555 (N_9555,N_7328,N_5116);
and U9556 (N_9556,N_5604,N_5226);
and U9557 (N_9557,N_7196,N_7080);
or U9558 (N_9558,N_5850,N_6041);
nand U9559 (N_9559,N_6757,N_5300);
nor U9560 (N_9560,N_6470,N_5729);
nor U9561 (N_9561,N_5127,N_6461);
or U9562 (N_9562,N_6082,N_5146);
nor U9563 (N_9563,N_5132,N_5364);
nand U9564 (N_9564,N_7211,N_5060);
xnor U9565 (N_9565,N_6419,N_7287);
and U9566 (N_9566,N_6854,N_5845);
or U9567 (N_9567,N_5205,N_6144);
or U9568 (N_9568,N_7175,N_7220);
nand U9569 (N_9569,N_5478,N_6868);
nand U9570 (N_9570,N_6398,N_5213);
nand U9571 (N_9571,N_5538,N_5115);
xnor U9572 (N_9572,N_7305,N_5071);
nand U9573 (N_9573,N_7417,N_7096);
nor U9574 (N_9574,N_5673,N_6548);
nand U9575 (N_9575,N_5153,N_5042);
nand U9576 (N_9576,N_6438,N_6745);
nand U9577 (N_9577,N_6106,N_7188);
and U9578 (N_9578,N_5020,N_5850);
or U9579 (N_9579,N_5649,N_5326);
and U9580 (N_9580,N_6419,N_6652);
nor U9581 (N_9581,N_7072,N_6516);
and U9582 (N_9582,N_7376,N_5515);
xnor U9583 (N_9583,N_6390,N_7103);
or U9584 (N_9584,N_5358,N_6712);
and U9585 (N_9585,N_5798,N_5548);
and U9586 (N_9586,N_7035,N_6474);
and U9587 (N_9587,N_7293,N_5742);
or U9588 (N_9588,N_5525,N_6509);
nand U9589 (N_9589,N_7434,N_6349);
nand U9590 (N_9590,N_5388,N_6874);
and U9591 (N_9591,N_6740,N_6272);
nand U9592 (N_9592,N_5638,N_6082);
xor U9593 (N_9593,N_6870,N_6830);
or U9594 (N_9594,N_5219,N_5173);
and U9595 (N_9595,N_5284,N_5909);
nand U9596 (N_9596,N_6484,N_5566);
xnor U9597 (N_9597,N_6600,N_6356);
nand U9598 (N_9598,N_6444,N_7247);
nand U9599 (N_9599,N_6237,N_6049);
or U9600 (N_9600,N_5333,N_6353);
xnor U9601 (N_9601,N_6060,N_5931);
and U9602 (N_9602,N_5294,N_7483);
nand U9603 (N_9603,N_6575,N_6968);
nor U9604 (N_9604,N_5374,N_5418);
or U9605 (N_9605,N_5632,N_5478);
xor U9606 (N_9606,N_6606,N_6062);
nand U9607 (N_9607,N_5278,N_6535);
nor U9608 (N_9608,N_5601,N_6900);
and U9609 (N_9609,N_7182,N_5982);
and U9610 (N_9610,N_6104,N_5443);
nand U9611 (N_9611,N_7166,N_6244);
or U9612 (N_9612,N_7280,N_6875);
or U9613 (N_9613,N_5891,N_6871);
nand U9614 (N_9614,N_6140,N_5936);
and U9615 (N_9615,N_5206,N_6599);
nor U9616 (N_9616,N_6775,N_5978);
nor U9617 (N_9617,N_6934,N_6746);
nor U9618 (N_9618,N_7117,N_6126);
or U9619 (N_9619,N_7319,N_5302);
nor U9620 (N_9620,N_5295,N_7328);
and U9621 (N_9621,N_6420,N_6708);
nand U9622 (N_9622,N_6114,N_7060);
nand U9623 (N_9623,N_7209,N_7117);
and U9624 (N_9624,N_5489,N_6256);
nand U9625 (N_9625,N_5955,N_6599);
xor U9626 (N_9626,N_5582,N_6508);
nor U9627 (N_9627,N_6791,N_6980);
xor U9628 (N_9628,N_7227,N_7376);
and U9629 (N_9629,N_6061,N_6079);
nor U9630 (N_9630,N_5746,N_5486);
nand U9631 (N_9631,N_7362,N_5106);
or U9632 (N_9632,N_6877,N_6217);
nor U9633 (N_9633,N_6328,N_7118);
nand U9634 (N_9634,N_7437,N_5873);
and U9635 (N_9635,N_6308,N_7211);
nand U9636 (N_9636,N_6054,N_7352);
xnor U9637 (N_9637,N_7213,N_6526);
nor U9638 (N_9638,N_5657,N_6540);
nand U9639 (N_9639,N_6427,N_6178);
and U9640 (N_9640,N_6164,N_7044);
and U9641 (N_9641,N_5319,N_6658);
nand U9642 (N_9642,N_6444,N_7112);
nor U9643 (N_9643,N_6950,N_6570);
and U9644 (N_9644,N_5934,N_6672);
or U9645 (N_9645,N_6485,N_6633);
and U9646 (N_9646,N_5724,N_6040);
or U9647 (N_9647,N_6225,N_6260);
and U9648 (N_9648,N_5836,N_5510);
nor U9649 (N_9649,N_5441,N_6758);
nand U9650 (N_9650,N_6792,N_6136);
and U9651 (N_9651,N_5071,N_7175);
nor U9652 (N_9652,N_7369,N_7101);
or U9653 (N_9653,N_6643,N_5015);
and U9654 (N_9654,N_6014,N_6077);
nand U9655 (N_9655,N_6394,N_7414);
and U9656 (N_9656,N_6027,N_5843);
or U9657 (N_9657,N_7078,N_5758);
nor U9658 (N_9658,N_5422,N_5200);
or U9659 (N_9659,N_6006,N_5330);
nor U9660 (N_9660,N_7105,N_7308);
or U9661 (N_9661,N_6822,N_6858);
nand U9662 (N_9662,N_5956,N_6130);
nor U9663 (N_9663,N_5397,N_6902);
xnor U9664 (N_9664,N_6697,N_5054);
nor U9665 (N_9665,N_6121,N_6893);
or U9666 (N_9666,N_5928,N_7176);
and U9667 (N_9667,N_5528,N_7094);
or U9668 (N_9668,N_5403,N_7397);
or U9669 (N_9669,N_7283,N_6237);
or U9670 (N_9670,N_6719,N_7058);
nor U9671 (N_9671,N_5073,N_7399);
xnor U9672 (N_9672,N_7261,N_6415);
or U9673 (N_9673,N_7165,N_7140);
nor U9674 (N_9674,N_6295,N_5214);
nand U9675 (N_9675,N_7087,N_5392);
nor U9676 (N_9676,N_7164,N_6792);
nand U9677 (N_9677,N_6110,N_6354);
and U9678 (N_9678,N_5650,N_6531);
nor U9679 (N_9679,N_5568,N_5481);
or U9680 (N_9680,N_6219,N_5566);
and U9681 (N_9681,N_5350,N_6870);
or U9682 (N_9682,N_7261,N_7400);
and U9683 (N_9683,N_5800,N_6465);
and U9684 (N_9684,N_6314,N_5308);
or U9685 (N_9685,N_5997,N_5742);
nor U9686 (N_9686,N_6914,N_6637);
xor U9687 (N_9687,N_6184,N_5446);
nor U9688 (N_9688,N_7339,N_6998);
and U9689 (N_9689,N_6776,N_5959);
nand U9690 (N_9690,N_6406,N_7105);
nor U9691 (N_9691,N_5735,N_7220);
nand U9692 (N_9692,N_5924,N_6540);
or U9693 (N_9693,N_7265,N_7453);
nand U9694 (N_9694,N_7368,N_5021);
and U9695 (N_9695,N_5000,N_7446);
or U9696 (N_9696,N_5250,N_6577);
or U9697 (N_9697,N_6538,N_6483);
nor U9698 (N_9698,N_6991,N_5870);
nor U9699 (N_9699,N_6943,N_6392);
nor U9700 (N_9700,N_7307,N_5259);
and U9701 (N_9701,N_5430,N_6878);
nand U9702 (N_9702,N_6014,N_5243);
nand U9703 (N_9703,N_6998,N_6677);
nor U9704 (N_9704,N_5820,N_6046);
and U9705 (N_9705,N_5757,N_5900);
or U9706 (N_9706,N_5796,N_7489);
nand U9707 (N_9707,N_6860,N_7091);
nor U9708 (N_9708,N_6460,N_5160);
nor U9709 (N_9709,N_6304,N_6044);
xor U9710 (N_9710,N_5746,N_6889);
and U9711 (N_9711,N_7041,N_7033);
nand U9712 (N_9712,N_5641,N_7050);
nor U9713 (N_9713,N_6642,N_5406);
or U9714 (N_9714,N_5832,N_5082);
and U9715 (N_9715,N_5740,N_6186);
xnor U9716 (N_9716,N_7134,N_7130);
nand U9717 (N_9717,N_5176,N_5033);
xor U9718 (N_9718,N_6989,N_6178);
nor U9719 (N_9719,N_6541,N_6778);
nor U9720 (N_9720,N_7314,N_6800);
and U9721 (N_9721,N_7406,N_7409);
nand U9722 (N_9722,N_6232,N_7305);
nor U9723 (N_9723,N_6825,N_5933);
xnor U9724 (N_9724,N_5951,N_5569);
and U9725 (N_9725,N_6827,N_5563);
and U9726 (N_9726,N_5235,N_6320);
nand U9727 (N_9727,N_5380,N_5248);
nand U9728 (N_9728,N_6580,N_5781);
or U9729 (N_9729,N_5776,N_7093);
nor U9730 (N_9730,N_6695,N_5094);
or U9731 (N_9731,N_5794,N_5743);
and U9732 (N_9732,N_6909,N_5472);
and U9733 (N_9733,N_5867,N_6657);
or U9734 (N_9734,N_7192,N_5803);
or U9735 (N_9735,N_6895,N_6179);
and U9736 (N_9736,N_6003,N_6848);
nand U9737 (N_9737,N_6233,N_5467);
nand U9738 (N_9738,N_5143,N_6531);
xor U9739 (N_9739,N_6026,N_6532);
or U9740 (N_9740,N_5807,N_6802);
nand U9741 (N_9741,N_5439,N_7090);
nand U9742 (N_9742,N_5224,N_5578);
or U9743 (N_9743,N_5471,N_7122);
nor U9744 (N_9744,N_5695,N_7147);
and U9745 (N_9745,N_7409,N_6923);
nand U9746 (N_9746,N_6272,N_5121);
and U9747 (N_9747,N_6574,N_6015);
nor U9748 (N_9748,N_5464,N_5943);
and U9749 (N_9749,N_5335,N_6895);
xor U9750 (N_9750,N_6442,N_5868);
nand U9751 (N_9751,N_5472,N_5857);
nor U9752 (N_9752,N_6404,N_6229);
or U9753 (N_9753,N_6994,N_6290);
nand U9754 (N_9754,N_5918,N_6315);
xnor U9755 (N_9755,N_5043,N_6386);
or U9756 (N_9756,N_5824,N_6449);
xnor U9757 (N_9757,N_5424,N_6635);
or U9758 (N_9758,N_7069,N_6137);
or U9759 (N_9759,N_7207,N_6427);
and U9760 (N_9760,N_5631,N_6033);
nand U9761 (N_9761,N_7331,N_5685);
and U9762 (N_9762,N_6327,N_5055);
nor U9763 (N_9763,N_5894,N_5008);
or U9764 (N_9764,N_5270,N_7096);
nand U9765 (N_9765,N_5913,N_6709);
xor U9766 (N_9766,N_6510,N_7346);
nor U9767 (N_9767,N_6239,N_5919);
and U9768 (N_9768,N_5233,N_5028);
or U9769 (N_9769,N_6731,N_7119);
and U9770 (N_9770,N_5635,N_5049);
or U9771 (N_9771,N_5819,N_7283);
or U9772 (N_9772,N_6590,N_5428);
nand U9773 (N_9773,N_5919,N_6337);
nand U9774 (N_9774,N_5975,N_6124);
nor U9775 (N_9775,N_7218,N_6811);
nor U9776 (N_9776,N_6012,N_5893);
nand U9777 (N_9777,N_6220,N_5075);
or U9778 (N_9778,N_5417,N_6881);
and U9779 (N_9779,N_6176,N_5429);
nand U9780 (N_9780,N_6732,N_6096);
nor U9781 (N_9781,N_6117,N_5562);
xnor U9782 (N_9782,N_5750,N_5103);
and U9783 (N_9783,N_6821,N_6601);
and U9784 (N_9784,N_6332,N_5994);
and U9785 (N_9785,N_6076,N_6211);
or U9786 (N_9786,N_7296,N_7413);
and U9787 (N_9787,N_6915,N_7428);
nand U9788 (N_9788,N_6569,N_5286);
or U9789 (N_9789,N_5116,N_6770);
or U9790 (N_9790,N_7177,N_6059);
and U9791 (N_9791,N_6902,N_7493);
and U9792 (N_9792,N_6845,N_7362);
and U9793 (N_9793,N_6150,N_6325);
nand U9794 (N_9794,N_7171,N_7215);
or U9795 (N_9795,N_6380,N_6133);
nor U9796 (N_9796,N_6992,N_6069);
and U9797 (N_9797,N_6586,N_6649);
and U9798 (N_9798,N_6548,N_5236);
nand U9799 (N_9799,N_6471,N_6300);
and U9800 (N_9800,N_5573,N_6783);
nand U9801 (N_9801,N_7104,N_5489);
or U9802 (N_9802,N_7089,N_5417);
or U9803 (N_9803,N_6295,N_5941);
xor U9804 (N_9804,N_6125,N_5610);
or U9805 (N_9805,N_5200,N_5938);
nand U9806 (N_9806,N_6667,N_6462);
nand U9807 (N_9807,N_6300,N_6873);
nor U9808 (N_9808,N_7228,N_5246);
nor U9809 (N_9809,N_5029,N_5943);
nor U9810 (N_9810,N_6627,N_5163);
or U9811 (N_9811,N_6545,N_5626);
and U9812 (N_9812,N_7127,N_7021);
xnor U9813 (N_9813,N_5127,N_5648);
or U9814 (N_9814,N_7454,N_5065);
nor U9815 (N_9815,N_7280,N_5022);
xor U9816 (N_9816,N_6402,N_5881);
and U9817 (N_9817,N_5741,N_7042);
and U9818 (N_9818,N_5785,N_5989);
nor U9819 (N_9819,N_7320,N_5306);
and U9820 (N_9820,N_6779,N_6281);
or U9821 (N_9821,N_6255,N_5721);
or U9822 (N_9822,N_5917,N_7281);
and U9823 (N_9823,N_5032,N_7012);
nand U9824 (N_9824,N_6241,N_6587);
or U9825 (N_9825,N_6742,N_7134);
nand U9826 (N_9826,N_5736,N_5311);
nand U9827 (N_9827,N_5552,N_5578);
or U9828 (N_9828,N_5457,N_6023);
nand U9829 (N_9829,N_5061,N_5472);
or U9830 (N_9830,N_5146,N_5996);
or U9831 (N_9831,N_6417,N_7049);
nor U9832 (N_9832,N_5957,N_5687);
nor U9833 (N_9833,N_7272,N_5057);
nor U9834 (N_9834,N_5934,N_5491);
nor U9835 (N_9835,N_6061,N_7216);
xor U9836 (N_9836,N_5230,N_5665);
nor U9837 (N_9837,N_5123,N_6916);
nor U9838 (N_9838,N_6069,N_6477);
or U9839 (N_9839,N_7008,N_5697);
nor U9840 (N_9840,N_7041,N_6785);
or U9841 (N_9841,N_6494,N_6203);
or U9842 (N_9842,N_5889,N_5068);
nand U9843 (N_9843,N_5672,N_5610);
nor U9844 (N_9844,N_6134,N_6004);
or U9845 (N_9845,N_5583,N_7092);
nand U9846 (N_9846,N_6102,N_7443);
nand U9847 (N_9847,N_6796,N_6742);
or U9848 (N_9848,N_6303,N_5201);
and U9849 (N_9849,N_5159,N_6483);
nor U9850 (N_9850,N_5203,N_6330);
nand U9851 (N_9851,N_6647,N_6873);
and U9852 (N_9852,N_5479,N_6012);
nand U9853 (N_9853,N_6026,N_5438);
and U9854 (N_9854,N_5544,N_5403);
nor U9855 (N_9855,N_7067,N_7095);
nor U9856 (N_9856,N_5428,N_5393);
or U9857 (N_9857,N_6485,N_5331);
nand U9858 (N_9858,N_7058,N_5322);
or U9859 (N_9859,N_5172,N_6278);
nor U9860 (N_9860,N_6719,N_7043);
nand U9861 (N_9861,N_6754,N_6304);
or U9862 (N_9862,N_7353,N_5553);
nor U9863 (N_9863,N_7345,N_7462);
or U9864 (N_9864,N_5729,N_7438);
nor U9865 (N_9865,N_6099,N_5248);
or U9866 (N_9866,N_5758,N_6094);
nand U9867 (N_9867,N_5176,N_6680);
and U9868 (N_9868,N_7151,N_7226);
or U9869 (N_9869,N_6000,N_5903);
nand U9870 (N_9870,N_5332,N_7161);
or U9871 (N_9871,N_6759,N_5209);
and U9872 (N_9872,N_6996,N_5379);
and U9873 (N_9873,N_6204,N_5397);
and U9874 (N_9874,N_6252,N_5320);
nand U9875 (N_9875,N_6918,N_6240);
xor U9876 (N_9876,N_5089,N_5628);
nand U9877 (N_9877,N_6273,N_7063);
xnor U9878 (N_9878,N_7211,N_7365);
nor U9879 (N_9879,N_6072,N_7332);
xor U9880 (N_9880,N_5266,N_5538);
nand U9881 (N_9881,N_5438,N_7256);
and U9882 (N_9882,N_5332,N_6582);
nand U9883 (N_9883,N_5595,N_7408);
or U9884 (N_9884,N_6991,N_5562);
nand U9885 (N_9885,N_5865,N_5276);
and U9886 (N_9886,N_7232,N_5198);
nand U9887 (N_9887,N_7323,N_6759);
or U9888 (N_9888,N_7216,N_7384);
and U9889 (N_9889,N_6558,N_5651);
nor U9890 (N_9890,N_5785,N_6544);
nand U9891 (N_9891,N_5402,N_5931);
and U9892 (N_9892,N_5294,N_6288);
and U9893 (N_9893,N_5780,N_6375);
xnor U9894 (N_9894,N_7168,N_6784);
and U9895 (N_9895,N_6700,N_5968);
nand U9896 (N_9896,N_5933,N_6336);
nor U9897 (N_9897,N_5246,N_7048);
nand U9898 (N_9898,N_5112,N_6953);
and U9899 (N_9899,N_5000,N_6020);
and U9900 (N_9900,N_7134,N_6775);
or U9901 (N_9901,N_5711,N_5907);
xor U9902 (N_9902,N_5184,N_5821);
nand U9903 (N_9903,N_5909,N_5066);
nand U9904 (N_9904,N_6815,N_5136);
and U9905 (N_9905,N_7448,N_5525);
nand U9906 (N_9906,N_6908,N_5687);
nor U9907 (N_9907,N_6299,N_6700);
nand U9908 (N_9908,N_6967,N_5335);
and U9909 (N_9909,N_5490,N_6057);
nor U9910 (N_9910,N_5284,N_7026);
and U9911 (N_9911,N_6119,N_6521);
or U9912 (N_9912,N_5638,N_5410);
nand U9913 (N_9913,N_7397,N_5357);
or U9914 (N_9914,N_6969,N_6588);
or U9915 (N_9915,N_5391,N_6667);
or U9916 (N_9916,N_6187,N_5723);
or U9917 (N_9917,N_5170,N_5628);
and U9918 (N_9918,N_6741,N_5946);
or U9919 (N_9919,N_6237,N_6885);
or U9920 (N_9920,N_7176,N_5400);
or U9921 (N_9921,N_5854,N_6149);
nor U9922 (N_9922,N_7438,N_5456);
nor U9923 (N_9923,N_7188,N_6981);
or U9924 (N_9924,N_5632,N_5875);
nand U9925 (N_9925,N_6566,N_7204);
nor U9926 (N_9926,N_6756,N_5285);
and U9927 (N_9927,N_6073,N_6020);
and U9928 (N_9928,N_7105,N_5154);
nand U9929 (N_9929,N_5067,N_5542);
nor U9930 (N_9930,N_6505,N_5347);
or U9931 (N_9931,N_6389,N_7337);
nor U9932 (N_9932,N_7305,N_6312);
nor U9933 (N_9933,N_5969,N_5997);
or U9934 (N_9934,N_6028,N_7053);
xor U9935 (N_9935,N_6656,N_6981);
nand U9936 (N_9936,N_5559,N_6767);
and U9937 (N_9937,N_5310,N_5682);
xnor U9938 (N_9938,N_6200,N_5997);
nor U9939 (N_9939,N_6122,N_5310);
or U9940 (N_9940,N_6298,N_6114);
and U9941 (N_9941,N_6749,N_6550);
xor U9942 (N_9942,N_6508,N_6934);
nand U9943 (N_9943,N_5400,N_5118);
nand U9944 (N_9944,N_6175,N_5417);
or U9945 (N_9945,N_6493,N_5960);
nand U9946 (N_9946,N_5892,N_6865);
nand U9947 (N_9947,N_5445,N_5747);
nor U9948 (N_9948,N_5915,N_6710);
nand U9949 (N_9949,N_6057,N_6279);
nor U9950 (N_9950,N_6268,N_5963);
and U9951 (N_9951,N_6496,N_5164);
nand U9952 (N_9952,N_5202,N_6956);
nand U9953 (N_9953,N_6130,N_6625);
or U9954 (N_9954,N_6761,N_5670);
and U9955 (N_9955,N_5344,N_6474);
nor U9956 (N_9956,N_5183,N_6227);
xnor U9957 (N_9957,N_7114,N_5319);
or U9958 (N_9958,N_5211,N_6765);
nor U9959 (N_9959,N_6783,N_6798);
nand U9960 (N_9960,N_7161,N_7311);
and U9961 (N_9961,N_5275,N_7040);
nand U9962 (N_9962,N_7253,N_5466);
xnor U9963 (N_9963,N_7493,N_6436);
nand U9964 (N_9964,N_5799,N_6917);
xor U9965 (N_9965,N_6258,N_6015);
nor U9966 (N_9966,N_6976,N_5558);
nand U9967 (N_9967,N_5476,N_6449);
or U9968 (N_9968,N_6277,N_7491);
nor U9969 (N_9969,N_5946,N_6715);
or U9970 (N_9970,N_6278,N_6717);
xor U9971 (N_9971,N_5137,N_7415);
nor U9972 (N_9972,N_6726,N_6190);
and U9973 (N_9973,N_6503,N_7301);
and U9974 (N_9974,N_6495,N_5944);
nor U9975 (N_9975,N_7323,N_5553);
and U9976 (N_9976,N_6974,N_6810);
and U9977 (N_9977,N_7444,N_7210);
nand U9978 (N_9978,N_5927,N_5712);
nand U9979 (N_9979,N_6898,N_7330);
and U9980 (N_9980,N_5856,N_5768);
and U9981 (N_9981,N_5394,N_6103);
nand U9982 (N_9982,N_5510,N_6302);
and U9983 (N_9983,N_6674,N_5574);
and U9984 (N_9984,N_5253,N_5265);
nor U9985 (N_9985,N_5829,N_5901);
nor U9986 (N_9986,N_5082,N_7450);
nor U9987 (N_9987,N_5320,N_6572);
xor U9988 (N_9988,N_5612,N_6039);
or U9989 (N_9989,N_6148,N_7261);
and U9990 (N_9990,N_7274,N_5013);
or U9991 (N_9991,N_6619,N_5858);
nor U9992 (N_9992,N_6270,N_7322);
nor U9993 (N_9993,N_6334,N_5271);
nor U9994 (N_9994,N_6615,N_6535);
and U9995 (N_9995,N_7337,N_6931);
nand U9996 (N_9996,N_5717,N_5704);
nor U9997 (N_9997,N_6857,N_5198);
and U9998 (N_9998,N_5714,N_7394);
nand U9999 (N_9999,N_7213,N_6381);
nand UO_0 (O_0,N_9046,N_8368);
nand UO_1 (O_1,N_9167,N_9237);
xor UO_2 (O_2,N_9309,N_9854);
xnor UO_3 (O_3,N_9956,N_9009);
nand UO_4 (O_4,N_8228,N_8920);
nand UO_5 (O_5,N_7987,N_8247);
nand UO_6 (O_6,N_7834,N_7807);
or UO_7 (O_7,N_9640,N_8703);
nand UO_8 (O_8,N_7598,N_9491);
or UO_9 (O_9,N_8925,N_8435);
or UO_10 (O_10,N_7515,N_8497);
nor UO_11 (O_11,N_9344,N_8307);
and UO_12 (O_12,N_7625,N_7956);
or UO_13 (O_13,N_8187,N_8130);
or UO_14 (O_14,N_8238,N_7603);
or UO_15 (O_15,N_9884,N_8677);
nor UO_16 (O_16,N_8655,N_7907);
or UO_17 (O_17,N_8980,N_9204);
nand UO_18 (O_18,N_9539,N_9739);
nand UO_19 (O_19,N_8005,N_8107);
nor UO_20 (O_20,N_9688,N_7870);
nor UO_21 (O_21,N_9432,N_9462);
nand UO_22 (O_22,N_8200,N_9814);
nand UO_23 (O_23,N_8310,N_9496);
nor UO_24 (O_24,N_8627,N_7716);
and UO_25 (O_25,N_8382,N_8082);
xor UO_26 (O_26,N_8018,N_7861);
and UO_27 (O_27,N_9725,N_9799);
nor UO_28 (O_28,N_9468,N_8838);
and UO_29 (O_29,N_8999,N_8882);
nor UO_30 (O_30,N_8557,N_8386);
nand UO_31 (O_31,N_9599,N_9114);
and UO_32 (O_32,N_9765,N_8278);
or UO_33 (O_33,N_8768,N_7761);
nand UO_34 (O_34,N_9016,N_7812);
nor UO_35 (O_35,N_8051,N_9969);
or UO_36 (O_36,N_7689,N_9377);
or UO_37 (O_37,N_8198,N_9062);
or UO_38 (O_38,N_9078,N_8601);
nor UO_39 (O_39,N_8282,N_7756);
xor UO_40 (O_40,N_7882,N_9647);
nand UO_41 (O_41,N_8816,N_9895);
and UO_42 (O_42,N_8496,N_7811);
and UO_43 (O_43,N_7579,N_7558);
nand UO_44 (O_44,N_8068,N_9897);
and UO_45 (O_45,N_8837,N_7702);
or UO_46 (O_46,N_7650,N_8258);
and UO_47 (O_47,N_8296,N_7878);
or UO_48 (O_48,N_9194,N_9545);
nand UO_49 (O_49,N_7779,N_8734);
nor UO_50 (O_50,N_7648,N_9913);
nor UO_51 (O_51,N_9181,N_9811);
or UO_52 (O_52,N_9446,N_8193);
xor UO_53 (O_53,N_9626,N_9853);
or UO_54 (O_54,N_9148,N_8305);
nor UO_55 (O_55,N_9451,N_8745);
or UO_56 (O_56,N_8050,N_7610);
nor UO_57 (O_57,N_8169,N_8602);
and UO_58 (O_58,N_8913,N_9521);
nand UO_59 (O_59,N_9748,N_8861);
or UO_60 (O_60,N_8342,N_8625);
or UO_61 (O_61,N_9924,N_9296);
or UO_62 (O_62,N_8621,N_7729);
nand UO_63 (O_63,N_8775,N_7540);
nor UO_64 (O_64,N_9749,N_8929);
xor UO_65 (O_65,N_8670,N_7970);
xnor UO_66 (O_66,N_7887,N_8979);
nor UO_67 (O_67,N_7923,N_9794);
nor UO_68 (O_68,N_9634,N_7918);
xor UO_69 (O_69,N_8385,N_7897);
and UO_70 (O_70,N_8460,N_8680);
nor UO_71 (O_71,N_7928,N_7661);
and UO_72 (O_72,N_8922,N_7613);
xor UO_73 (O_73,N_9721,N_8585);
xor UO_74 (O_74,N_9240,N_9285);
nor UO_75 (O_75,N_9017,N_7857);
and UO_76 (O_76,N_8847,N_9820);
or UO_77 (O_77,N_7662,N_8065);
and UO_78 (O_78,N_7571,N_7708);
and UO_79 (O_79,N_7858,N_7775);
xor UO_80 (O_80,N_7960,N_7977);
xnor UO_81 (O_81,N_7596,N_9067);
nor UO_82 (O_82,N_9973,N_9308);
or UO_83 (O_83,N_8459,N_9633);
nor UO_84 (O_84,N_9024,N_9733);
or UO_85 (O_85,N_8309,N_9396);
and UO_86 (O_86,N_7803,N_9759);
or UO_87 (O_87,N_9697,N_7595);
and UO_88 (O_88,N_8067,N_7880);
nand UO_89 (O_89,N_9326,N_9176);
and UO_90 (O_90,N_9949,N_8622);
or UO_91 (O_91,N_8807,N_8889);
nor UO_92 (O_92,N_9511,N_8188);
and UO_93 (O_93,N_8249,N_7532);
nor UO_94 (O_94,N_8448,N_9710);
or UO_95 (O_95,N_9034,N_9779);
and UO_96 (O_96,N_8289,N_8600);
and UO_97 (O_97,N_7594,N_9767);
nand UO_98 (O_98,N_8336,N_9330);
or UO_99 (O_99,N_9110,N_9631);
nor UO_100 (O_100,N_8832,N_8070);
and UO_101 (O_101,N_8572,N_8300);
xor UO_102 (O_102,N_7521,N_8467);
or UO_103 (O_103,N_9586,N_9984);
nor UO_104 (O_104,N_9112,N_9757);
nor UO_105 (O_105,N_9337,N_8081);
or UO_106 (O_106,N_7704,N_7673);
or UO_107 (O_107,N_7863,N_8683);
nand UO_108 (O_108,N_7743,N_8692);
nand UO_109 (O_109,N_9249,N_8842);
nand UO_110 (O_110,N_8858,N_7640);
nor UO_111 (O_111,N_9116,N_7758);
nor UO_112 (O_112,N_9758,N_9977);
nand UO_113 (O_113,N_7505,N_8091);
nand UO_114 (O_114,N_8161,N_8634);
nand UO_115 (O_115,N_9089,N_7942);
nor UO_116 (O_116,N_7721,N_9628);
nor UO_117 (O_117,N_8660,N_7591);
xnor UO_118 (O_118,N_8127,N_8209);
nor UO_119 (O_119,N_9000,N_7762);
nor UO_120 (O_120,N_9132,N_8511);
nor UO_121 (O_121,N_8916,N_8063);
nor UO_122 (O_122,N_9598,N_8001);
or UO_123 (O_123,N_9549,N_8079);
and UO_124 (O_124,N_8821,N_9904);
xor UO_125 (O_125,N_8756,N_9095);
and UO_126 (O_126,N_9713,N_7760);
and UO_127 (O_127,N_9778,N_9121);
and UO_128 (O_128,N_8545,N_8790);
nor UO_129 (O_129,N_8784,N_7685);
or UO_130 (O_130,N_9026,N_8774);
or UO_131 (O_131,N_8515,N_8725);
nand UO_132 (O_132,N_8495,N_8077);
and UO_133 (O_133,N_8513,N_8984);
nor UO_134 (O_134,N_7632,N_8960);
nand UO_135 (O_135,N_8281,N_8851);
nor UO_136 (O_136,N_9192,N_9944);
nand UO_137 (O_137,N_8854,N_8696);
nor UO_138 (O_138,N_9010,N_9130);
or UO_139 (O_139,N_9646,N_8071);
nand UO_140 (O_140,N_9102,N_8895);
nor UO_141 (O_141,N_9290,N_9146);
or UO_142 (O_142,N_9054,N_9145);
xor UO_143 (O_143,N_7774,N_9013);
nor UO_144 (O_144,N_8152,N_8679);
xnor UO_145 (O_145,N_9063,N_8226);
xnor UO_146 (O_146,N_8326,N_9193);
nand UO_147 (O_147,N_8346,N_8918);
and UO_148 (O_148,N_9244,N_7581);
or UO_149 (O_149,N_9178,N_7826);
or UO_150 (O_150,N_8678,N_9839);
nand UO_151 (O_151,N_8706,N_8803);
nor UO_152 (O_152,N_7612,N_7836);
nor UO_153 (O_153,N_8163,N_8903);
nand UO_154 (O_154,N_8186,N_9412);
and UO_155 (O_155,N_8479,N_8273);
nor UO_156 (O_156,N_9907,N_8165);
and UO_157 (O_157,N_9686,N_8761);
or UO_158 (O_158,N_7525,N_8554);
and UO_159 (O_159,N_8594,N_8325);
xnor UO_160 (O_160,N_7664,N_9528);
xnor UO_161 (O_161,N_8840,N_8164);
nor UO_162 (O_162,N_7962,N_8137);
nand UO_163 (O_163,N_7895,N_7845);
or UO_164 (O_164,N_8045,N_8713);
nor UO_165 (O_165,N_8826,N_7999);
nor UO_166 (O_166,N_8134,N_9608);
and UO_167 (O_167,N_9906,N_9845);
and UO_168 (O_168,N_9045,N_8741);
and UO_169 (O_169,N_7993,N_9606);
nor UO_170 (O_170,N_9952,N_9732);
nand UO_171 (O_171,N_9578,N_9123);
or UO_172 (O_172,N_9039,N_7922);
and UO_173 (O_173,N_7900,N_9982);
nand UO_174 (O_174,N_8264,N_9097);
or UO_175 (O_175,N_8409,N_7949);
and UO_176 (O_176,N_7957,N_8522);
nand UO_177 (O_177,N_9008,N_8879);
and UO_178 (O_178,N_9235,N_8181);
or UO_179 (O_179,N_9753,N_9573);
and UO_180 (O_180,N_7682,N_9090);
nand UO_181 (O_181,N_9442,N_7551);
nand UO_182 (O_182,N_7838,N_7941);
or UO_183 (O_183,N_9464,N_8619);
nand UO_184 (O_184,N_7599,N_8915);
and UO_185 (O_185,N_8824,N_9630);
nor UO_186 (O_186,N_9107,N_7780);
nor UO_187 (O_187,N_8773,N_9415);
and UO_188 (O_188,N_8484,N_8794);
nor UO_189 (O_189,N_8883,N_9898);
and UO_190 (O_190,N_8370,N_9447);
nand UO_191 (O_191,N_7932,N_8593);
or UO_192 (O_192,N_7731,N_8415);
and UO_193 (O_193,N_9041,N_9659);
nor UO_194 (O_194,N_9080,N_9541);
and UO_195 (O_195,N_9159,N_9623);
or UO_196 (O_196,N_9014,N_8738);
or UO_197 (O_197,N_8724,N_9938);
and UO_198 (O_198,N_7770,N_7933);
nand UO_199 (O_199,N_9066,N_8770);
or UO_200 (O_200,N_8235,N_9282);
nor UO_201 (O_201,N_9975,N_9570);
nor UO_202 (O_202,N_9142,N_9558);
nor UO_203 (O_203,N_8700,N_7914);
xnor UO_204 (O_204,N_8175,N_8269);
xnor UO_205 (O_205,N_7924,N_8553);
nor UO_206 (O_206,N_8406,N_8290);
nor UO_207 (O_207,N_8482,N_9133);
nor UO_208 (O_208,N_8072,N_7734);
xor UO_209 (O_209,N_8203,N_8168);
and UO_210 (O_210,N_8252,N_8897);
xnor UO_211 (O_211,N_9744,N_9380);
nor UO_212 (O_212,N_9997,N_9324);
or UO_213 (O_213,N_8248,N_8791);
or UO_214 (O_214,N_8280,N_8646);
nor UO_215 (O_215,N_8514,N_8982);
and UO_216 (O_216,N_8781,N_8214);
nor UO_217 (O_217,N_8195,N_8872);
xnor UO_218 (O_218,N_8739,N_8061);
or UO_219 (O_219,N_8940,N_9652);
xor UO_220 (O_220,N_9136,N_8580);
or UO_221 (O_221,N_7853,N_9156);
and UO_222 (O_222,N_9163,N_9583);
nor UO_223 (O_223,N_8444,N_7755);
nand UO_224 (O_224,N_8934,N_9632);
or UO_225 (O_225,N_9661,N_9715);
xnor UO_226 (O_226,N_8292,N_9060);
xnor UO_227 (O_227,N_8230,N_9465);
xnor UO_228 (O_228,N_8836,N_8016);
xnor UO_229 (O_229,N_9591,N_9636);
and UO_230 (O_230,N_9188,N_9401);
and UO_231 (O_231,N_9349,N_8046);
xor UO_232 (O_232,N_9049,N_9774);
nand UO_233 (O_233,N_9362,N_9702);
or UO_234 (O_234,N_9942,N_8588);
or UO_235 (O_235,N_8464,N_9727);
nand UO_236 (O_236,N_8870,N_8294);
nand UO_237 (O_237,N_8701,N_8087);
nor UO_238 (O_238,N_9453,N_9796);
nor UO_239 (O_239,N_9791,N_8517);
and UO_240 (O_240,N_9911,N_8413);
nor UO_241 (O_241,N_9352,N_7510);
nor UO_242 (O_242,N_9197,N_8062);
nand UO_243 (O_243,N_8592,N_8390);
nor UO_244 (O_244,N_9689,N_8088);
or UO_245 (O_245,N_9088,N_7604);
nand UO_246 (O_246,N_9140,N_8989);
or UO_247 (O_247,N_8287,N_8229);
nor UO_248 (O_248,N_9119,N_8623);
xor UO_249 (O_249,N_7693,N_8610);
or UO_250 (O_250,N_8695,N_8277);
xnor UO_251 (O_251,N_8035,N_7503);
nand UO_252 (O_252,N_8472,N_9797);
and UO_253 (O_253,N_8505,N_8025);
nand UO_254 (O_254,N_7618,N_7726);
nor UO_255 (O_255,N_7806,N_9775);
nor UO_256 (O_256,N_8587,N_7808);
xor UO_257 (O_257,N_8526,N_9162);
nand UO_258 (O_258,N_8059,N_8441);
and UO_259 (O_259,N_8667,N_7943);
nor UO_260 (O_260,N_9871,N_8105);
nand UO_261 (O_261,N_7679,N_9786);
nor UO_262 (O_262,N_8657,N_8122);
xor UO_263 (O_263,N_9720,N_9667);
nor UO_264 (O_264,N_8691,N_8629);
and UO_265 (O_265,N_8097,N_8952);
xnor UO_266 (O_266,N_9113,N_8179);
or UO_267 (O_267,N_8301,N_8260);
nand UO_268 (O_268,N_7874,N_9238);
nand UO_269 (O_269,N_8375,N_9379);
nand UO_270 (O_270,N_8788,N_9695);
nand UO_271 (O_271,N_9478,N_9083);
or UO_272 (O_272,N_8106,N_9025);
xnor UO_273 (O_273,N_7725,N_9649);
nor UO_274 (O_274,N_9663,N_7630);
or UO_275 (O_275,N_8686,N_9654);
xnor UO_276 (O_276,N_8008,N_8777);
nand UO_277 (O_277,N_8893,N_8757);
nor UO_278 (O_278,N_9172,N_9691);
or UO_279 (O_279,N_8101,N_7569);
and UO_280 (O_280,N_9553,N_8210);
nor UO_281 (O_281,N_9407,N_9115);
and UO_282 (O_282,N_8891,N_8769);
nor UO_283 (O_283,N_7651,N_8672);
nand UO_284 (O_284,N_9760,N_7837);
or UO_285 (O_285,N_9445,N_8446);
nand UO_286 (O_286,N_8886,N_8199);
nor UO_287 (O_287,N_8957,N_8437);
and UO_288 (O_288,N_9681,N_9053);
and UO_289 (O_289,N_8272,N_8457);
nor UO_290 (O_290,N_8365,N_8829);
nor UO_291 (O_291,N_9889,N_8284);
or UO_292 (O_292,N_9494,N_7717);
nand UO_293 (O_293,N_7930,N_9392);
nor UO_294 (O_294,N_9502,N_7681);
and UO_295 (O_295,N_8846,N_8397);
nor UO_296 (O_296,N_8033,N_7627);
or UO_297 (O_297,N_7549,N_9376);
xnor UO_298 (O_298,N_9310,N_9917);
and UO_299 (O_299,N_8149,N_9746);
and UO_300 (O_300,N_9941,N_8715);
and UO_301 (O_301,N_8407,N_9712);
or UO_302 (O_302,N_8494,N_7582);
nor UO_303 (O_303,N_9269,N_9461);
nor UO_304 (O_304,N_9229,N_7733);
xnor UO_305 (O_305,N_9666,N_7656);
xor UO_306 (O_306,N_8483,N_9831);
or UO_307 (O_307,N_9523,N_7903);
nor UO_308 (O_308,N_8919,N_8845);
nand UO_309 (O_309,N_8392,N_7840);
nand UO_310 (O_310,N_8898,N_8324);
nand UO_311 (O_311,N_8996,N_8881);
nor UO_312 (O_312,N_8500,N_8933);
nor UO_313 (O_313,N_8647,N_7884);
nand UO_314 (O_314,N_8378,N_7931);
nand UO_315 (O_315,N_8136,N_8755);
nor UO_316 (O_316,N_8477,N_9160);
xor UO_317 (O_317,N_9274,N_8147);
nand UO_318 (O_318,N_7963,N_9260);
or UO_319 (O_319,N_8314,N_8866);
and UO_320 (O_320,N_9498,N_8640);
nand UO_321 (O_321,N_9111,N_9363);
nor UO_322 (O_322,N_9481,N_9910);
and UO_323 (O_323,N_9564,N_9679);
nand UO_324 (O_324,N_8040,N_8731);
nand UO_325 (O_325,N_8772,N_8352);
xnor UO_326 (O_326,N_9307,N_8116);
nand UO_327 (O_327,N_9169,N_9439);
xor UO_328 (O_328,N_8562,N_9124);
or UO_329 (O_329,N_8053,N_7677);
nor UO_330 (O_330,N_8556,N_9387);
nand UO_331 (O_331,N_9236,N_7773);
nand UO_332 (O_332,N_7537,N_8519);
nor UO_333 (O_333,N_9700,N_9708);
or UO_334 (O_334,N_9391,N_9751);
and UO_335 (O_335,N_8128,N_7747);
or UO_336 (O_336,N_7516,N_8567);
nand UO_337 (O_337,N_9306,N_8251);
and UO_338 (O_338,N_9655,N_8434);
nand UO_339 (O_339,N_7652,N_9203);
or UO_340 (O_340,N_8732,N_8429);
xnor UO_341 (O_341,N_7683,N_8455);
nand UO_342 (O_342,N_8084,N_7601);
nor UO_343 (O_343,N_7655,N_9769);
and UO_344 (O_344,N_9635,N_8148);
nor UO_345 (O_345,N_8218,N_9345);
nand UO_346 (O_346,N_9986,N_8591);
or UO_347 (O_347,N_9218,N_7902);
nand UO_348 (O_348,N_8958,N_8792);
and UO_349 (O_349,N_7753,N_8445);
or UO_350 (O_350,N_8298,N_9288);
or UO_351 (O_351,N_9311,N_9604);
nand UO_352 (O_352,N_8574,N_9280);
xnor UO_353 (O_353,N_8937,N_8906);
or UO_354 (O_354,N_8261,N_8151);
nor UO_355 (O_355,N_7752,N_7908);
nand UO_356 (O_356,N_8674,N_9825);
nor UO_357 (O_357,N_9386,N_9576);
xor UO_358 (O_358,N_9817,N_7890);
and UO_359 (O_359,N_8205,N_9701);
and UO_360 (O_360,N_7621,N_8085);
nand UO_361 (O_361,N_9058,N_8395);
or UO_362 (O_362,N_7722,N_9619);
or UO_363 (O_363,N_8236,N_7978);
nor UO_364 (O_364,N_7827,N_9291);
xnor UO_365 (O_365,N_8146,N_7705);
or UO_366 (O_366,N_7919,N_8120);
nand UO_367 (O_367,N_7881,N_8825);
and UO_368 (O_368,N_8361,N_8034);
and UO_369 (O_369,N_7665,N_8800);
and UO_370 (O_370,N_8394,N_8564);
and UO_371 (O_371,N_9543,N_9151);
xor UO_372 (O_372,N_9228,N_8759);
nor UO_373 (O_373,N_8869,N_8389);
nand UO_374 (O_374,N_9965,N_9990);
nand UO_375 (O_375,N_8143,N_8740);
and UO_376 (O_376,N_9348,N_9245);
or UO_377 (O_377,N_7719,N_7622);
xnor UO_378 (O_378,N_9873,N_8321);
nand UO_379 (O_379,N_7940,N_9546);
or UO_380 (O_380,N_8381,N_9189);
nand UO_381 (O_381,N_9876,N_8664);
xor UO_382 (O_382,N_8002,N_8341);
or UO_383 (O_383,N_9484,N_9092);
nand UO_384 (O_384,N_8797,N_8643);
nand UO_385 (O_385,N_8243,N_8650);
nand UO_386 (O_386,N_9927,N_8004);
and UO_387 (O_387,N_9674,N_7698);
nand UO_388 (O_388,N_8661,N_7684);
and UO_389 (O_389,N_8440,N_9448);
nand UO_390 (O_390,N_8166,N_9785);
nor UO_391 (O_391,N_8132,N_7851);
nand UO_392 (O_392,N_8470,N_7706);
and UO_393 (O_393,N_8049,N_8899);
nand UO_394 (O_394,N_8583,N_9637);
nor UO_395 (O_395,N_9807,N_9668);
nor UO_396 (O_396,N_8665,N_9756);
xnor UO_397 (O_397,N_9077,N_8539);
nand UO_398 (O_398,N_7565,N_8931);
or UO_399 (O_399,N_8177,N_9592);
nand UO_400 (O_400,N_8430,N_9430);
and UO_401 (O_401,N_8417,N_8206);
xor UO_402 (O_402,N_7634,N_9566);
and UO_403 (O_403,N_7842,N_9995);
xor UO_404 (O_404,N_7678,N_9048);
or UO_405 (O_405,N_7846,N_8543);
nand UO_406 (O_406,N_9317,N_8981);
nand UO_407 (O_407,N_7660,N_8877);
and UO_408 (O_408,N_9648,N_9118);
xnor UO_409 (O_409,N_7785,N_7546);
nor UO_410 (O_410,N_8080,N_7983);
or UO_411 (O_411,N_7860,N_8157);
and UO_412 (O_412,N_9257,N_9273);
xor UO_413 (O_413,N_7669,N_9641);
and UO_414 (O_414,N_7750,N_9959);
nand UO_415 (O_415,N_9165,N_9125);
nor UO_416 (O_416,N_8758,N_8786);
or UO_417 (O_417,N_9342,N_8349);
and UO_418 (O_418,N_8345,N_9772);
nor UO_419 (O_419,N_7562,N_7805);
or UO_420 (O_420,N_9370,N_8827);
nand UO_421 (O_421,N_9364,N_9542);
nor UO_422 (O_422,N_8485,N_7982);
and UO_423 (O_423,N_8656,N_9792);
and UO_424 (O_424,N_9431,N_8379);
nand UO_425 (O_425,N_7985,N_7776);
and UO_426 (O_426,N_8427,N_8953);
and UO_427 (O_427,N_8598,N_8374);
or UO_428 (O_428,N_9886,N_8491);
nand UO_429 (O_429,N_8182,N_8632);
or UO_430 (O_430,N_9699,N_9375);
and UO_431 (O_431,N_7644,N_9537);
nand UO_432 (O_432,N_9517,N_9402);
or UO_433 (O_433,N_8548,N_7732);
nand UO_434 (O_434,N_8635,N_8612);
and UO_435 (O_435,N_8951,N_8167);
and UO_436 (O_436,N_7671,N_8862);
nand UO_437 (O_437,N_8527,N_9787);
nand UO_438 (O_438,N_9321,N_8549);
or UO_439 (O_439,N_8276,N_8596);
or UO_440 (O_440,N_9253,N_8852);
nand UO_441 (O_441,N_9444,N_9126);
nor UO_442 (O_442,N_8456,N_9656);
nor UO_443 (O_443,N_9467,N_8425);
nand UO_444 (O_444,N_8924,N_7892);
nand UO_445 (O_445,N_8969,N_8371);
or UO_446 (O_446,N_9736,N_9955);
and UO_447 (O_447,N_8254,N_9161);
nor UO_448 (O_448,N_9371,N_9294);
or UO_449 (O_449,N_8244,N_8697);
or UO_450 (O_450,N_9105,N_8092);
and UO_451 (O_451,N_8089,N_7935);
or UO_452 (O_452,N_7680,N_8098);
and UO_453 (O_453,N_8654,N_7637);
nand UO_454 (O_454,N_8323,N_8422);
and UO_455 (O_455,N_8523,N_9551);
nand UO_456 (O_456,N_8416,N_8954);
nor UO_457 (O_457,N_9851,N_8799);
or UO_458 (O_458,N_8037,N_9243);
and UO_459 (O_459,N_9532,N_9056);
and UO_460 (O_460,N_9002,N_9104);
and UO_461 (O_461,N_8871,N_9190);
or UO_462 (O_462,N_8110,N_8138);
nor UO_463 (O_463,N_9471,N_8998);
or UO_464 (O_464,N_8923,N_8652);
nand UO_465 (O_465,N_9263,N_9057);
or UO_466 (O_466,N_8579,N_7988);
or UO_467 (O_467,N_9622,N_9507);
or UO_468 (O_468,N_9771,N_9798);
nor UO_469 (O_469,N_7763,N_8538);
nand UO_470 (O_470,N_8212,N_7920);
nor UO_471 (O_471,N_8356,N_8577);
and UO_472 (O_472,N_8613,N_8744);
and UO_473 (O_473,N_8584,N_7607);
or UO_474 (O_474,N_8443,N_7667);
or UO_475 (O_475,N_8279,N_9200);
nor UO_476 (O_476,N_9241,N_9144);
nand UO_477 (O_477,N_8461,N_9770);
nor UO_478 (O_478,N_9030,N_9331);
or UO_479 (O_479,N_9084,N_9452);
or UO_480 (O_480,N_8291,N_8508);
nor UO_481 (O_481,N_7556,N_9497);
nand UO_482 (O_482,N_9847,N_8819);
nor UO_483 (O_483,N_9234,N_9281);
and UO_484 (O_484,N_7620,N_8322);
and UO_485 (O_485,N_9212,N_9168);
xnor UO_486 (O_486,N_8458,N_8340);
and UO_487 (O_487,N_7936,N_7605);
xor UO_488 (O_488,N_9037,N_8178);
and UO_489 (O_489,N_9410,N_8853);
and UO_490 (O_490,N_8946,N_8867);
and UO_491 (O_491,N_9676,N_8333);
nor UO_492 (O_492,N_9741,N_9185);
and UO_493 (O_493,N_8265,N_9888);
and UO_494 (O_494,N_8609,N_8830);
and UO_495 (O_495,N_9781,N_9355);
nor UO_496 (O_496,N_8075,N_9143);
or UO_497 (O_497,N_9696,N_7700);
or UO_498 (O_498,N_9411,N_8242);
or UO_499 (O_499,N_9488,N_9252);
xnor UO_500 (O_500,N_9091,N_8078);
xor UO_501 (O_501,N_9743,N_8058);
nor UO_502 (O_502,N_9519,N_7991);
nand UO_503 (O_503,N_9400,N_9035);
nand UO_504 (O_504,N_9584,N_9662);
nand UO_505 (O_505,N_9283,N_8771);
or UO_506 (O_506,N_9441,N_8114);
xor UO_507 (O_507,N_7759,N_8997);
or UO_508 (O_508,N_8473,N_9428);
or UO_509 (O_509,N_8928,N_9485);
nand UO_510 (O_510,N_7735,N_8331);
or UO_511 (O_511,N_9079,N_7976);
and UO_512 (O_512,N_8751,N_8710);
or UO_513 (O_513,N_8589,N_9878);
and UO_514 (O_514,N_8544,N_9803);
nor UO_515 (O_515,N_9808,N_7699);
nor UO_516 (O_516,N_8471,N_9023);
nand UO_517 (O_517,N_8343,N_7668);
nand UO_518 (O_518,N_8673,N_8512);
and UO_519 (O_519,N_9624,N_7666);
nor UO_520 (O_520,N_8848,N_8676);
nor UO_521 (O_521,N_9617,N_9303);
nand UO_522 (O_522,N_8396,N_8558);
nand UO_523 (O_523,N_8225,N_9675);
or UO_524 (O_524,N_7786,N_8237);
or UO_525 (O_525,N_8570,N_9475);
nor UO_526 (O_526,N_9065,N_9219);
nor UO_527 (O_527,N_9800,N_7889);
and UO_528 (O_528,N_9101,N_9343);
or UO_529 (O_529,N_9227,N_8224);
nand UO_530 (O_530,N_8766,N_9215);
or UO_531 (O_531,N_8955,N_7707);
and UO_532 (O_532,N_9231,N_9184);
and UO_533 (O_533,N_8787,N_9199);
or UO_534 (O_534,N_9540,N_7995);
nor UO_535 (O_535,N_9265,N_9134);
and UO_536 (O_536,N_8384,N_8438);
nand UO_537 (O_537,N_7535,N_7524);
or UO_538 (O_538,N_9585,N_7772);
nor UO_539 (O_539,N_8536,N_9479);
nor UO_540 (O_540,N_9258,N_7990);
nor UO_541 (O_541,N_7911,N_9536);
nand UO_542 (O_542,N_9301,N_8022);
or UO_543 (O_543,N_8108,N_8090);
and UO_544 (O_544,N_8297,N_9305);
or UO_545 (O_545,N_8469,N_8476);
nand UO_546 (O_546,N_8581,N_7996);
xor UO_547 (O_547,N_8874,N_7738);
nor UO_548 (O_548,N_8763,N_7597);
nand UO_549 (O_549,N_8685,N_8723);
nand UO_550 (O_550,N_9226,N_8509);
or UO_551 (O_551,N_9106,N_8991);
nor UO_552 (O_552,N_8191,N_8863);
nor UO_553 (O_553,N_8246,N_7574);
or UO_554 (O_554,N_9382,N_9826);
and UO_555 (O_555,N_8754,N_7934);
nand UO_556 (O_556,N_8023,N_9603);
nor UO_557 (O_557,N_9147,N_8817);
xnor UO_558 (O_558,N_8466,N_8319);
nand UO_559 (O_559,N_9403,N_7619);
and UO_560 (O_560,N_9454,N_9153);
and UO_561 (O_561,N_9434,N_8782);
nand UO_562 (O_562,N_7832,N_9071);
nor UO_563 (O_563,N_9544,N_9120);
or UO_564 (O_564,N_9864,N_9529);
nor UO_565 (O_565,N_7550,N_9690);
nand UO_566 (O_566,N_9810,N_9332);
nor UO_567 (O_567,N_9027,N_8971);
xnor UO_568 (O_568,N_8006,N_8890);
or UO_569 (O_569,N_9416,N_8052);
or UO_570 (O_570,N_8488,N_8943);
or UO_571 (O_571,N_8611,N_9866);
nor UO_572 (O_572,N_9266,N_7833);
and UO_573 (O_573,N_9435,N_9210);
or UO_574 (O_574,N_9354,N_9616);
or UO_575 (O_575,N_9117,N_7968);
nor UO_576 (O_576,N_9038,N_9706);
xor UO_577 (O_577,N_9378,N_8947);
xor UO_578 (O_578,N_9032,N_9154);
or UO_579 (O_579,N_8335,N_8347);
and UO_580 (O_580,N_8135,N_7636);
and UO_581 (O_581,N_8912,N_9295);
nand UO_582 (O_582,N_8303,N_7998);
nor UO_583 (O_583,N_9472,N_7568);
nor UO_584 (O_584,N_9830,N_9320);
and UO_585 (O_585,N_8144,N_9367);
or UO_586 (O_586,N_9893,N_8293);
or UO_587 (O_587,N_9683,N_9992);
and UO_588 (O_588,N_8233,N_7536);
nand UO_589 (O_589,N_8798,N_8312);
nor UO_590 (O_590,N_9985,N_9885);
nor UO_591 (O_591,N_9064,N_9398);
or UO_592 (O_592,N_7560,N_8639);
nor UO_593 (O_593,N_7590,N_8994);
and UO_594 (O_594,N_9870,N_7647);
nand UO_595 (O_595,N_8709,N_8043);
nand UO_596 (O_596,N_8820,N_9006);
nor UO_597 (O_597,N_8516,N_8631);
nand UO_598 (O_598,N_8704,N_8808);
and UO_599 (O_599,N_9590,N_9863);
or UO_600 (O_600,N_8930,N_9891);
or UO_601 (O_601,N_7641,N_8501);
and UO_602 (O_602,N_9011,N_8121);
or UO_603 (O_603,N_7514,N_7946);
xnor UO_604 (O_604,N_7791,N_9874);
or UO_605 (O_605,N_8537,N_9928);
and UO_606 (O_606,N_9859,N_8180);
xor UO_607 (O_607,N_9846,N_8487);
or UO_608 (O_608,N_8941,N_8117);
or UO_609 (O_609,N_9728,N_9552);
or UO_610 (O_610,N_8486,N_8690);
nand UO_611 (O_611,N_8131,N_9705);
nand UO_612 (O_612,N_9882,N_9642);
nor UO_613 (O_613,N_9408,N_9276);
and UO_614 (O_614,N_9561,N_9493);
and UO_615 (O_615,N_9429,N_9339);
nor UO_616 (O_616,N_8542,N_9503);
and UO_617 (O_617,N_9230,N_8119);
or UO_618 (O_618,N_8216,N_8945);
nor UO_619 (O_619,N_8990,N_8054);
nand UO_620 (O_620,N_9328,N_9868);
and UO_621 (O_621,N_7718,N_8547);
nand UO_622 (O_622,N_7703,N_7517);
and UO_623 (O_623,N_8350,N_8129);
or UO_624 (O_624,N_9206,N_9042);
nand UO_625 (O_625,N_8125,N_9179);
and UO_626 (O_626,N_7530,N_9374);
or UO_627 (O_627,N_9180,N_9588);
and UO_628 (O_628,N_7809,N_9987);
or UO_629 (O_629,N_9195,N_8843);
nor UO_630 (O_630,N_9335,N_8630);
nand UO_631 (O_631,N_8133,N_7973);
nor UO_632 (O_632,N_8172,N_7847);
nand UO_633 (O_633,N_8267,N_9963);
and UO_634 (O_634,N_8113,N_8066);
xor UO_635 (O_635,N_8103,N_8100);
nand UO_636 (O_636,N_9530,N_8648);
nor UO_637 (O_637,N_8211,N_9737);
nor UO_638 (O_638,N_8628,N_9722);
nand UO_639 (O_639,N_7764,N_9605);
nand UO_640 (O_640,N_9248,N_8256);
nand UO_641 (O_641,N_7865,N_7898);
or UO_642 (O_642,N_9670,N_9596);
nand UO_643 (O_643,N_9141,N_9182);
and UO_644 (O_644,N_7697,N_9848);
nor UO_645 (O_645,N_7580,N_8568);
or UO_646 (O_646,N_8565,N_9233);
xor UO_647 (O_647,N_8737,N_8624);
and UO_648 (O_648,N_9840,N_9004);
or UO_649 (O_649,N_8644,N_9922);
and UO_650 (O_650,N_8401,N_7927);
nand UO_651 (O_651,N_7944,N_9538);
and UO_652 (O_652,N_8687,N_9424);
and UO_653 (O_653,N_9455,N_9970);
nand UO_654 (O_654,N_8606,N_9698);
nor UO_655 (O_655,N_7511,N_9993);
or UO_656 (O_656,N_8047,N_9157);
nor UO_657 (O_657,N_8804,N_8714);
nand UO_658 (O_658,N_8746,N_9187);
nand UO_659 (O_659,N_8927,N_9805);
nand UO_660 (O_660,N_7715,N_9998);
nand UO_661 (O_661,N_7787,N_8115);
nor UO_662 (O_662,N_9466,N_7686);
and UO_663 (O_663,N_8860,N_9427);
or UO_664 (O_664,N_9012,N_9625);
nor UO_665 (O_665,N_9437,N_9593);
or UO_666 (O_666,N_9287,N_7921);
nor UO_667 (O_667,N_7531,N_8231);
and UO_668 (O_668,N_8659,N_9395);
nand UO_669 (O_669,N_8617,N_9262);
nand UO_670 (O_670,N_9806,N_8405);
xor UO_671 (O_671,N_7642,N_9338);
nand UO_672 (O_672,N_8976,N_9094);
or UO_673 (O_673,N_8400,N_8949);
nand UO_674 (O_674,N_8533,N_7984);
and UO_675 (O_675,N_8170,N_7835);
nor UO_676 (O_676,N_8096,N_7573);
xnor UO_677 (O_677,N_9535,N_7994);
or UO_678 (O_678,N_9967,N_8073);
nor UO_679 (O_679,N_8330,N_8124);
and UO_680 (O_680,N_7810,N_8876);
and UO_681 (O_681,N_9047,N_8914);
and UO_682 (O_682,N_9394,N_9043);
nand UO_683 (O_683,N_9589,N_7819);
nor UO_684 (O_684,N_9620,N_8174);
nor UO_685 (O_685,N_9372,N_7696);
xor UO_686 (O_686,N_8317,N_9718);
or UO_687 (O_687,N_7793,N_9098);
and UO_688 (O_688,N_8720,N_9368);
or UO_689 (O_689,N_8234,N_9818);
nand UO_690 (O_690,N_7958,N_9061);
nand UO_691 (O_691,N_7894,N_8353);
or UO_692 (O_692,N_8828,N_8304);
and UO_693 (O_693,N_8318,N_8268);
or UO_694 (O_694,N_9137,N_7986);
xor UO_695 (O_695,N_9334,N_9857);
nand UO_696 (O_696,N_8344,N_7901);
or UO_697 (O_697,N_8966,N_9242);
or UO_698 (O_698,N_9389,N_7623);
nand UO_699 (O_699,N_9912,N_8550);
and UO_700 (O_700,N_7638,N_8048);
xor UO_701 (O_701,N_9835,N_9671);
nor UO_702 (O_702,N_7831,N_9919);
or UO_703 (O_703,N_9764,N_8451);
nor UO_704 (O_704,N_8474,N_8559);
or UO_705 (O_705,N_8419,N_8616);
nor UO_706 (O_706,N_9515,N_7553);
nor UO_707 (O_707,N_7746,N_9714);
nor UO_708 (O_708,N_9677,N_9469);
nor UO_709 (O_709,N_8041,N_7742);
or UO_710 (O_710,N_8926,N_8299);
nand UO_711 (O_711,N_7563,N_7820);
xnor UO_712 (O_712,N_9068,N_9350);
nand UO_713 (O_713,N_9336,N_7979);
and UO_714 (O_714,N_9999,N_8126);
or UO_715 (O_715,N_9881,N_7768);
nor UO_716 (O_716,N_8393,N_8032);
nor UO_717 (O_717,N_8590,N_9657);
xor UO_718 (O_718,N_8698,N_9149);
nand UO_719 (O_719,N_8521,N_8995);
nand UO_720 (O_720,N_8420,N_8283);
nand UO_721 (O_721,N_7893,N_9173);
or UO_722 (O_722,N_8109,N_9802);
nor UO_723 (O_723,N_9202,N_7804);
or UO_724 (O_724,N_9255,N_8607);
nor UO_725 (O_725,N_9356,N_9555);
nand UO_726 (O_726,N_9417,N_7714);
or UO_727 (O_727,N_9152,N_8726);
nor UO_728 (O_728,N_7692,N_7615);
nand UO_729 (O_729,N_8074,N_8262);
and UO_730 (O_730,N_8493,N_7769);
nor UO_731 (O_731,N_9828,N_8532);
nand UO_732 (O_732,N_7789,N_7614);
nor UO_733 (O_733,N_9135,N_9833);
or UO_734 (O_734,N_9516,N_7788);
nor UO_735 (O_735,N_9658,N_9482);
and UO_736 (O_736,N_7867,N_7676);
nor UO_737 (O_737,N_9302,N_8604);
xnor UO_738 (O_738,N_9421,N_8868);
nand UO_739 (O_739,N_8973,N_9595);
nor UO_740 (O_740,N_9005,N_8963);
xor UO_741 (O_741,N_9093,N_9843);
and UO_742 (O_742,N_9790,N_9877);
or UO_743 (O_743,N_7839,N_9852);
nor UO_744 (O_744,N_8749,N_8056);
nor UO_745 (O_745,N_8197,N_7578);
and UO_746 (O_746,N_9456,N_7744);
or UO_747 (O_747,N_9347,N_7790);
nor UO_748 (O_748,N_7910,N_9246);
nor UO_749 (O_749,N_8575,N_9357);
or UO_750 (O_750,N_9001,N_8159);
or UO_751 (O_751,N_7929,N_9164);
nor UO_752 (O_752,N_7502,N_8295);
or UO_753 (O_753,N_9315,N_9100);
and UO_754 (O_754,N_9687,N_9645);
nand UO_755 (O_755,N_9196,N_9692);
and UO_756 (O_756,N_9867,N_8615);
and UO_757 (O_757,N_9947,N_8736);
nand UO_758 (O_758,N_7518,N_8932);
nand UO_759 (O_759,N_9651,N_8675);
and UO_760 (O_760,N_9353,N_8887);
or UO_761 (O_761,N_9858,N_8257);
nand UO_762 (O_762,N_8986,N_8140);
or UO_763 (O_763,N_9707,N_9286);
nand UO_764 (O_764,N_7745,N_9360);
or UO_765 (O_765,N_8366,N_9518);
nand UO_766 (O_766,N_9968,N_9709);
and UO_767 (O_767,N_7657,N_7883);
nand UO_768 (O_768,N_9860,N_7512);
and UO_769 (O_769,N_9669,N_7869);
or UO_770 (O_770,N_8069,N_9900);
or UO_771 (O_771,N_9127,N_8727);
nor UO_772 (O_772,N_8102,N_7965);
or UO_773 (O_773,N_9693,N_9438);
and UO_774 (O_774,N_8910,N_9129);
nand UO_775 (O_775,N_7913,N_9214);
nand UO_776 (O_776,N_7586,N_9894);
nor UO_777 (O_777,N_7937,N_8796);
xnor UO_778 (O_778,N_8901,N_8253);
nand UO_779 (O_779,N_8145,N_7777);
nor UO_780 (O_780,N_8728,N_9250);
and UO_781 (O_781,N_9905,N_8633);
and UO_782 (O_782,N_7792,N_9443);
nor UO_783 (O_783,N_9612,N_8850);
or UO_784 (O_784,N_8357,N_9932);
nand UO_785 (O_785,N_7794,N_9365);
nand UO_786 (O_786,N_9397,N_9665);
nor UO_787 (O_787,N_8414,N_8339);
xnor UO_788 (O_788,N_8201,N_7872);
or UO_789 (O_789,N_7961,N_8014);
or UO_790 (O_790,N_9929,N_7967);
and UO_791 (O_791,N_9954,N_7856);
or UO_792 (O_792,N_9404,N_9293);
xnor UO_793 (O_793,N_7815,N_7841);
or UO_794 (O_794,N_9903,N_9329);
nand UO_795 (O_795,N_7691,N_7823);
or UO_796 (O_796,N_9976,N_7658);
xor UO_797 (O_797,N_7824,N_7712);
or UO_798 (O_798,N_8988,N_8373);
or UO_799 (O_799,N_9572,N_8535);
nand UO_800 (O_800,N_8669,N_9856);
nand UO_801 (O_801,N_8007,N_8421);
nand UO_802 (O_802,N_9823,N_9450);
nor UO_803 (O_803,N_7947,N_8985);
or UO_804 (O_804,N_9405,N_7741);
nand UO_805 (O_805,N_7783,N_8377);
nor UO_806 (O_806,N_8974,N_7765);
nand UO_807 (O_807,N_8719,N_9128);
and UO_808 (O_808,N_9279,N_8241);
nand UO_809 (O_809,N_8546,N_8403);
or UO_810 (O_810,N_9015,N_8436);
nand UO_811 (O_811,N_9390,N_9074);
nand UO_812 (O_812,N_8399,N_7611);
nand UO_813 (O_813,N_9819,N_9961);
nand UO_814 (O_814,N_9936,N_8942);
xor UO_815 (O_815,N_7862,N_9524);
and UO_816 (O_816,N_8332,N_9815);
and UO_817 (O_817,N_7945,N_9300);
nor UO_818 (O_818,N_8908,N_8561);
nor UO_819 (O_819,N_9525,N_7570);
nand UO_820 (O_820,N_9081,N_9476);
xor UO_821 (O_821,N_8450,N_8510);
nor UO_822 (O_822,N_9514,N_9069);
nand UO_823 (O_823,N_9926,N_7544);
nand UO_824 (O_824,N_9232,N_8364);
or UO_825 (O_825,N_8428,N_9554);
nor UO_826 (O_826,N_8315,N_8823);
or UO_827 (O_827,N_9916,N_9816);
and UO_828 (O_828,N_9251,N_9527);
and UO_829 (O_829,N_8878,N_7916);
nand UO_830 (O_830,N_9580,N_8747);
and UO_831 (O_831,N_8266,N_7749);
nor UO_832 (O_832,N_9486,N_9103);
and UO_833 (O_833,N_8391,N_8935);
and UO_834 (O_834,N_8944,N_8620);
or UO_835 (O_835,N_8215,N_7915);
nand UO_836 (O_836,N_8964,N_8030);
nand UO_837 (O_837,N_9723,N_8563);
xor UO_838 (O_838,N_7844,N_8432);
nand UO_839 (O_839,N_9506,N_9562);
or UO_840 (O_840,N_9981,N_9865);
and UO_841 (O_841,N_8972,N_7906);
or UO_842 (O_842,N_7548,N_8095);
nor UO_843 (O_843,N_8658,N_7784);
and UO_844 (O_844,N_7821,N_8835);
or UO_845 (O_845,N_8813,N_8875);
or UO_846 (O_846,N_9166,N_7674);
nand UO_847 (O_847,N_9740,N_9072);
xor UO_848 (O_848,N_9931,N_9318);
or UO_849 (O_849,N_9406,N_8682);
xnor UO_850 (O_850,N_9509,N_9474);
nand UO_851 (O_851,N_7711,N_9684);
or UO_852 (O_852,N_8921,N_7800);
nor UO_853 (O_853,N_8693,N_8359);
xnor UO_854 (O_854,N_9278,N_9879);
and UO_855 (O_855,N_9019,N_8112);
and UO_856 (O_856,N_8688,N_8967);
nand UO_857 (O_857,N_7767,N_9734);
xor UO_858 (O_858,N_9569,N_9615);
or UO_859 (O_859,N_8153,N_7796);
or UO_860 (O_860,N_7520,N_9358);
nor UO_861 (O_861,N_8171,N_9614);
nor UO_862 (O_862,N_8009,N_9208);
xor UO_863 (O_863,N_8489,N_9974);
nor UO_864 (O_864,N_9018,N_9319);
xor UO_865 (O_865,N_8531,N_8019);
nor UO_866 (O_866,N_9534,N_9567);
nor UO_867 (O_867,N_9388,N_9508);
nand UO_868 (O_868,N_9385,N_7740);
or UO_869 (O_869,N_9703,N_9201);
nor UO_870 (O_870,N_7675,N_8900);
nor UO_871 (O_871,N_9076,N_7814);
or UO_872 (O_872,N_9694,N_7859);
nand UO_873 (O_873,N_9007,N_7891);
or UO_874 (O_874,N_8184,N_8123);
nor UO_875 (O_875,N_8111,N_8810);
nor UO_876 (O_876,N_9571,N_7951);
xor UO_877 (O_877,N_7538,N_9915);
nand UO_878 (O_878,N_8961,N_9827);
and UO_879 (O_879,N_7583,N_7500);
nand UO_880 (O_880,N_8662,N_8597);
or UO_881 (O_881,N_8762,N_7925);
xor UO_882 (O_882,N_9457,N_7825);
nor UO_883 (O_883,N_9685,N_8173);
nand UO_884 (O_884,N_7513,N_7875);
or UO_885 (O_885,N_9754,N_9109);
nor UO_886 (O_886,N_8442,N_7876);
nand UO_887 (O_887,N_8528,N_7948);
nor UO_888 (O_888,N_9075,N_9383);
nor UO_889 (O_889,N_7723,N_7670);
or UO_890 (O_890,N_9980,N_8223);
xnor UO_891 (O_891,N_7545,N_7828);
or UO_892 (O_892,N_9460,N_7829);
and UO_893 (O_893,N_7672,N_9836);
nor UO_894 (O_894,N_8599,N_8039);
or UO_895 (O_895,N_9678,N_7969);
nand UO_896 (O_896,N_9735,N_9221);
or UO_897 (O_897,N_9177,N_8831);
nor UO_898 (O_898,N_8185,N_7585);
nor UO_899 (O_899,N_9755,N_8959);
xnor UO_900 (O_900,N_8742,N_9579);
and UO_901 (O_901,N_8141,N_7751);
nor UO_902 (O_902,N_8042,N_8888);
xor UO_903 (O_903,N_8518,N_9021);
nor UO_904 (O_904,N_9499,N_8681);
or UO_905 (O_905,N_8334,N_8320);
nor UO_906 (O_906,N_8398,N_8003);
or UO_907 (O_907,N_8506,N_9838);
or UO_908 (O_908,N_9943,N_8540);
and UO_909 (O_909,N_8752,N_7871);
and UO_910 (O_910,N_8668,N_7509);
nor UO_911 (O_911,N_9051,N_9316);
nor UO_912 (O_912,N_9964,N_8316);
and UO_913 (O_913,N_8993,N_8263);
nand UO_914 (O_914,N_8699,N_9487);
or UO_915 (O_915,N_8271,N_8194);
nand UO_916 (O_916,N_9855,N_8055);
or UO_917 (O_917,N_9568,N_8760);
and UO_918 (O_918,N_8689,N_8894);
or UO_919 (O_919,N_8424,N_7798);
nand UO_920 (O_920,N_7541,N_9896);
nand UO_921 (O_921,N_7566,N_8478);
or UO_922 (O_922,N_9577,N_9582);
or UO_923 (O_923,N_8873,N_7849);
nand UO_924 (O_924,N_9272,N_9175);
xor UO_925 (O_925,N_8970,N_8499);
and UO_926 (O_926,N_9639,N_8498);
nor UO_927 (O_927,N_7631,N_8637);
or UO_928 (O_928,N_8809,N_8064);
nand UO_929 (O_929,N_8388,N_8475);
nor UO_930 (O_930,N_8351,N_8902);
nand UO_931 (O_931,N_9224,N_9556);
or UO_932 (O_932,N_8504,N_9271);
or UO_933 (O_933,N_8767,N_7964);
nor UO_934 (O_934,N_9784,N_7972);
nor UO_935 (O_935,N_9731,N_9322);
or UO_936 (O_936,N_9346,N_7576);
or UO_937 (O_937,N_8426,N_8507);
or UO_938 (O_938,N_9073,N_8892);
nand UO_939 (O_939,N_8560,N_7564);
and UO_940 (O_940,N_9433,N_7757);
nor UO_941 (O_941,N_9629,N_9565);
nor UO_942 (O_942,N_8849,N_7724);
or UO_943 (O_943,N_8387,N_9822);
or UO_944 (O_944,N_8239,N_7848);
nor UO_945 (O_945,N_9492,N_8844);
or UO_946 (O_946,N_8362,N_8530);
nand UO_947 (O_947,N_8452,N_8938);
and UO_948 (O_948,N_7778,N_8595);
nor UO_949 (O_949,N_7506,N_8576);
nor UO_950 (O_950,N_7617,N_9500);
or UO_951 (O_951,N_7593,N_7912);
and UO_952 (O_952,N_9277,N_8412);
nor UO_953 (O_953,N_8551,N_8404);
or UO_954 (O_954,N_9660,N_8636);
xor UO_955 (O_955,N_7852,N_9934);
nand UO_956 (O_956,N_8250,N_8571);
or UO_957 (O_957,N_9510,N_9373);
nor UO_958 (O_958,N_9801,N_9131);
nand UO_959 (O_959,N_7864,N_8118);
and UO_960 (O_960,N_9574,N_8222);
or UO_961 (O_961,N_8057,N_9384);
nor UO_962 (O_962,N_8453,N_9325);
nor UO_963 (O_963,N_8208,N_8801);
or UO_964 (O_964,N_7552,N_9183);
and UO_965 (O_965,N_8376,N_7600);
and UO_966 (O_966,N_8439,N_8806);
or UO_967 (O_967,N_8275,N_8402);
or UO_968 (O_968,N_7730,N_7539);
nor UO_969 (O_969,N_9717,N_7602);
and UO_970 (O_970,N_8534,N_7926);
and UO_971 (O_971,N_9824,N_9520);
nand UO_972 (O_972,N_8626,N_8603);
nand UO_973 (O_973,N_8864,N_7589);
xor UO_974 (O_974,N_8987,N_8904);
nand UO_975 (O_975,N_8983,N_9887);
nand UO_976 (O_976,N_7575,N_9220);
xor UO_977 (O_977,N_9420,N_8270);
xor UO_978 (O_978,N_9664,N_9908);
or UO_979 (O_979,N_8765,N_7559);
nand UO_980 (O_980,N_8423,N_8805);
nand UO_981 (O_981,N_7592,N_9899);
nand UO_982 (O_982,N_7639,N_9031);
nand UO_983 (O_983,N_7954,N_7754);
nor UO_984 (O_984,N_8814,N_9270);
and UO_985 (O_985,N_9440,N_8711);
nor UO_986 (O_986,N_9419,N_7748);
nand UO_987 (O_987,N_9747,N_7501);
nor UO_988 (O_988,N_9463,N_9361);
nor UO_989 (O_989,N_9186,N_8645);
nor UO_990 (O_990,N_9198,N_9930);
or UO_991 (O_991,N_8812,N_9426);
nand UO_992 (O_992,N_9399,N_9314);
nand UO_993 (O_993,N_8093,N_9490);
and UO_994 (O_994,N_7989,N_7905);
nor UO_995 (O_995,N_9036,N_9087);
or UO_996 (O_996,N_8492,N_8160);
nor UO_997 (O_997,N_9945,N_8083);
xor UO_998 (O_998,N_9070,N_8729);
nand UO_999 (O_999,N_9436,N_7830);
nand UO_1000 (O_1000,N_9773,N_8142);
xnor UO_1001 (O_1001,N_8031,N_7817);
nand UO_1002 (O_1002,N_8044,N_8750);
nor UO_1003 (O_1003,N_9653,N_9366);
or UO_1004 (O_1004,N_9842,N_9957);
and UO_1005 (O_1005,N_8183,N_9480);
xnor UO_1006 (O_1006,N_7523,N_8360);
nand UO_1007 (O_1007,N_9875,N_9108);
and UO_1008 (O_1008,N_8641,N_8541);
xor UO_1009 (O_1009,N_8060,N_8705);
xnor UO_1010 (O_1010,N_8369,N_7507);
or UO_1011 (O_1011,N_9526,N_9547);
and UO_1012 (O_1012,N_9312,N_8716);
or UO_1013 (O_1013,N_9033,N_8529);
or UO_1014 (O_1014,N_9972,N_9607);
nor UO_1015 (O_1015,N_9872,N_9505);
and UO_1016 (O_1016,N_9594,N_9359);
and UO_1017 (O_1017,N_8748,N_9531);
xor UO_1018 (O_1018,N_9247,N_8372);
nand UO_1019 (O_1019,N_7542,N_8431);
nor UO_1020 (O_1020,N_9044,N_9022);
nor UO_1021 (O_1021,N_8789,N_8605);
or UO_1022 (O_1022,N_9745,N_8329);
or UO_1023 (O_1023,N_7646,N_9761);
nor UO_1024 (O_1024,N_7997,N_9909);
nand UO_1025 (O_1025,N_9750,N_8753);
nand UO_1026 (O_1026,N_8013,N_7688);
nand UO_1027 (O_1027,N_9978,N_9489);
and UO_1028 (O_1028,N_9730,N_9638);
and UO_1029 (O_1029,N_9951,N_9829);
and UO_1030 (O_1030,N_9050,N_9340);
xor UO_1031 (O_1031,N_7873,N_8020);
nor UO_1032 (O_1032,N_8480,N_8783);
xor UO_1033 (O_1033,N_9883,N_8992);
or UO_1034 (O_1034,N_7739,N_7766);
and UO_1035 (O_1035,N_9946,N_8712);
nand UO_1036 (O_1036,N_8348,N_9849);
or UO_1037 (O_1037,N_9766,N_8722);
nand UO_1038 (O_1038,N_7687,N_7917);
nand UO_1039 (O_1039,N_9804,N_7799);
nand UO_1040 (O_1040,N_9841,N_8354);
nand UO_1041 (O_1041,N_9205,N_7909);
or UO_1042 (O_1042,N_9850,N_8259);
nand UO_1043 (O_1043,N_8555,N_8217);
nand UO_1044 (O_1044,N_9522,N_9059);
xor UO_1045 (O_1045,N_8730,N_8306);
and UO_1046 (O_1046,N_8196,N_8255);
nand UO_1047 (O_1047,N_9207,N_9834);
nor UO_1048 (O_1048,N_8094,N_9213);
or UO_1049 (O_1049,N_9304,N_7522);
and UO_1050 (O_1050,N_9892,N_7533);
nor UO_1051 (O_1051,N_8839,N_8880);
or UO_1052 (O_1052,N_8337,N_8015);
xor UO_1053 (O_1053,N_8447,N_8856);
nor UO_1054 (O_1054,N_8502,N_9028);
nor UO_1055 (O_1055,N_7955,N_7885);
nand UO_1056 (O_1056,N_9122,N_9298);
or UO_1057 (O_1057,N_8965,N_9869);
nor UO_1058 (O_1058,N_7782,N_9793);
nand UO_1059 (O_1059,N_9933,N_8733);
or UO_1060 (O_1060,N_9991,N_8618);
nand UO_1061 (O_1061,N_9563,N_9560);
and UO_1062 (O_1062,N_8962,N_8653);
nor UO_1063 (O_1063,N_8302,N_9425);
nor UO_1064 (O_1064,N_8651,N_9971);
and UO_1065 (O_1065,N_8029,N_8614);
and UO_1066 (O_1066,N_7802,N_8717);
xnor UO_1067 (O_1067,N_8036,N_7843);
or UO_1068 (O_1068,N_7818,N_8156);
and UO_1069 (O_1069,N_7797,N_7567);
nand UO_1070 (O_1070,N_7816,N_8694);
and UO_1071 (O_1071,N_7801,N_9052);
or UO_1072 (O_1072,N_9948,N_9618);
nor UO_1073 (O_1073,N_8367,N_8917);
and UO_1074 (O_1074,N_8977,N_9672);
nor UO_1075 (O_1075,N_7854,N_8939);
xnor UO_1076 (O_1076,N_8795,N_9621);
nor UO_1077 (O_1077,N_8380,N_8189);
and UO_1078 (O_1078,N_9597,N_9763);
nor UO_1079 (O_1079,N_9020,N_7737);
xor UO_1080 (O_1080,N_8780,N_8684);
nand UO_1081 (O_1081,N_9611,N_7727);
and UO_1082 (O_1082,N_8285,N_7561);
or UO_1083 (O_1083,N_9704,N_9966);
nand UO_1084 (O_1084,N_9292,N_9960);
and UO_1085 (O_1085,N_9752,N_9254);
and UO_1086 (O_1086,N_7975,N_9953);
or UO_1087 (O_1087,N_8956,N_9155);
nand UO_1088 (O_1088,N_7822,N_9901);
and UO_1089 (O_1089,N_7939,N_8433);
and UO_1090 (O_1090,N_9483,N_8818);
nor UO_1091 (O_1091,N_7584,N_9459);
or UO_1092 (O_1092,N_9495,N_7877);
and UO_1093 (O_1093,N_7879,N_9962);
and UO_1094 (O_1094,N_8707,N_8274);
nand UO_1095 (O_1095,N_8465,N_9610);
and UO_1096 (O_1096,N_7577,N_9085);
or UO_1097 (O_1097,N_9267,N_9581);
nand UO_1098 (O_1098,N_8011,N_9171);
nand UO_1099 (O_1099,N_9158,N_8718);
nand UO_1100 (O_1100,N_8582,N_8884);
nand UO_1101 (O_1101,N_7629,N_7555);
or UO_1102 (O_1102,N_8139,N_9925);
and UO_1103 (O_1103,N_9575,N_9513);
nor UO_1104 (O_1104,N_8663,N_8288);
and UO_1105 (O_1105,N_7526,N_9724);
xor UO_1106 (O_1106,N_9225,N_8764);
nor UO_1107 (O_1107,N_9548,N_9351);
or UO_1108 (O_1108,N_7952,N_7606);
or UO_1109 (O_1109,N_7645,N_9789);
nand UO_1110 (O_1110,N_7527,N_9920);
and UO_1111 (O_1111,N_9550,N_8232);
nor UO_1112 (O_1112,N_8909,N_9040);
xor UO_1113 (O_1113,N_9477,N_8905);
nor UO_1114 (O_1114,N_9414,N_8463);
nand UO_1115 (O_1115,N_8202,N_8468);
nor UO_1116 (O_1116,N_9673,N_9812);
nand UO_1117 (O_1117,N_8950,N_8192);
nor UO_1118 (O_1118,N_7701,N_8776);
xnor UO_1119 (O_1119,N_9809,N_9381);
nand UO_1120 (O_1120,N_9191,N_9211);
or UO_1121 (O_1121,N_8176,N_8815);
or UO_1122 (O_1122,N_8104,N_9644);
nand UO_1123 (O_1123,N_7609,N_8811);
or UO_1124 (O_1124,N_8642,N_7850);
and UO_1125 (O_1125,N_8778,N_7572);
xor UO_1126 (O_1126,N_7966,N_7649);
and UO_1127 (O_1127,N_8162,N_7713);
and UO_1128 (O_1128,N_8076,N_7950);
or UO_1129 (O_1129,N_7519,N_7971);
or UO_1130 (O_1130,N_9261,N_9983);
and UO_1131 (O_1131,N_8671,N_8907);
nor UO_1132 (O_1132,N_7626,N_8702);
xor UO_1133 (O_1133,N_8219,N_7781);
xor UO_1134 (O_1134,N_9217,N_7959);
nor UO_1135 (O_1135,N_8190,N_9082);
nand UO_1136 (O_1136,N_8896,N_8418);
nor UO_1137 (O_1137,N_9174,N_9937);
or UO_1138 (O_1138,N_7635,N_8857);
xnor UO_1139 (O_1139,N_9473,N_7653);
or UO_1140 (O_1140,N_7643,N_8245);
nor UO_1141 (O_1141,N_8503,N_7709);
nor UO_1142 (O_1142,N_8012,N_8462);
nand UO_1143 (O_1143,N_9559,N_9413);
nor UO_1144 (O_1144,N_9029,N_9780);
nor UO_1145 (O_1145,N_9921,N_8569);
nor UO_1146 (O_1146,N_8411,N_9918);
or UO_1147 (O_1147,N_9284,N_8743);
nand UO_1148 (O_1148,N_9832,N_8338);
or UO_1149 (O_1149,N_9458,N_9880);
nor UO_1150 (O_1150,N_7981,N_7504);
and UO_1151 (O_1151,N_8026,N_9783);
nor UO_1152 (O_1152,N_8975,N_9259);
nand UO_1153 (O_1153,N_9989,N_9449);
or UO_1154 (O_1154,N_8978,N_9512);
nor UO_1155 (O_1155,N_7904,N_8566);
and UO_1156 (O_1156,N_8158,N_8525);
nand UO_1157 (O_1157,N_9776,N_9777);
or UO_1158 (O_1158,N_7771,N_9643);
or UO_1159 (O_1159,N_9150,N_9844);
or UO_1160 (O_1160,N_8028,N_9003);
or UO_1161 (O_1161,N_8220,N_7543);
or UO_1162 (O_1162,N_9609,N_7554);
xnor UO_1163 (O_1163,N_9979,N_7628);
or UO_1164 (O_1164,N_8865,N_7855);
nor UO_1165 (O_1165,N_8793,N_9861);
or UO_1166 (O_1166,N_7663,N_9768);
or UO_1167 (O_1167,N_7588,N_7659);
and UO_1168 (O_1168,N_8552,N_9627);
or UO_1169 (O_1169,N_8021,N_9557);
or UO_1170 (O_1170,N_9222,N_7720);
nor UO_1171 (O_1171,N_7624,N_7529);
xnor UO_1172 (O_1172,N_9837,N_7608);
nor UO_1173 (O_1173,N_9423,N_8449);
and UO_1174 (O_1174,N_9762,N_8150);
nor UO_1175 (O_1175,N_9223,N_8524);
nor UO_1176 (O_1176,N_9821,N_9940);
or UO_1177 (O_1177,N_9216,N_8227);
or UO_1178 (O_1178,N_9958,N_8936);
or UO_1179 (O_1179,N_9600,N_9323);
nand UO_1180 (O_1180,N_8649,N_7547);
and UO_1181 (O_1181,N_8154,N_9470);
or UO_1182 (O_1182,N_9729,N_7938);
nor UO_1183 (O_1183,N_8204,N_8666);
nor UO_1184 (O_1184,N_8355,N_7690);
and UO_1185 (O_1185,N_7868,N_7813);
or UO_1186 (O_1186,N_8885,N_7616);
and UO_1187 (O_1187,N_9788,N_9418);
xor UO_1188 (O_1188,N_9782,N_8155);
or UO_1189 (O_1189,N_9988,N_8520);
xor UO_1190 (O_1190,N_8721,N_8735);
or UO_1191 (O_1191,N_7888,N_8968);
or UO_1192 (O_1192,N_7795,N_9409);
nor UO_1193 (O_1193,N_8490,N_9716);
or UO_1194 (O_1194,N_9682,N_9726);
nand UO_1195 (O_1195,N_9422,N_9256);
or UO_1196 (O_1196,N_8833,N_9533);
or UO_1197 (O_1197,N_7896,N_8578);
nand UO_1198 (O_1198,N_7886,N_8099);
or UO_1199 (O_1199,N_9923,N_8311);
nor UO_1200 (O_1200,N_9299,N_7953);
and UO_1201 (O_1201,N_9275,N_9341);
nand UO_1202 (O_1202,N_8027,N_8221);
nor UO_1203 (O_1203,N_7633,N_9086);
nor UO_1204 (O_1204,N_7736,N_7710);
nor UO_1205 (O_1205,N_9738,N_9996);
and UO_1206 (O_1206,N_8383,N_9264);
nand UO_1207 (O_1207,N_9369,N_8038);
or UO_1208 (O_1208,N_8859,N_7899);
nor UO_1209 (O_1209,N_9602,N_7654);
nand UO_1210 (O_1210,N_9613,N_8841);
nand UO_1211 (O_1211,N_9711,N_8573);
nor UO_1212 (O_1212,N_9055,N_9504);
and UO_1213 (O_1213,N_8328,N_9239);
nor UO_1214 (O_1214,N_9680,N_9297);
or UO_1215 (O_1215,N_8240,N_8286);
xnor UO_1216 (O_1216,N_7980,N_9650);
nand UO_1217 (O_1217,N_8213,N_8327);
nand UO_1218 (O_1218,N_7695,N_7587);
nor UO_1219 (O_1219,N_8024,N_9138);
or UO_1220 (O_1220,N_7974,N_8363);
or UO_1221 (O_1221,N_9393,N_9813);
nor UO_1222 (O_1222,N_8638,N_9890);
nand UO_1223 (O_1223,N_8207,N_9501);
or UO_1224 (O_1224,N_9209,N_8802);
xnor UO_1225 (O_1225,N_9719,N_7866);
nor UO_1226 (O_1226,N_8410,N_9902);
nand UO_1227 (O_1227,N_9327,N_9587);
nor UO_1228 (O_1228,N_8481,N_9935);
and UO_1229 (O_1229,N_8000,N_8308);
nand UO_1230 (O_1230,N_9914,N_9099);
nor UO_1231 (O_1231,N_8834,N_8086);
xnor UO_1232 (O_1232,N_7534,N_8586);
and UO_1233 (O_1233,N_9333,N_9139);
xnor UO_1234 (O_1234,N_8313,N_8454);
nand UO_1235 (O_1235,N_8948,N_9795);
or UO_1236 (O_1236,N_8779,N_9950);
nand UO_1237 (O_1237,N_8822,N_8408);
xnor UO_1238 (O_1238,N_7728,N_7508);
nor UO_1239 (O_1239,N_7528,N_8855);
and UO_1240 (O_1240,N_9862,N_9742);
nand UO_1241 (O_1241,N_8911,N_8017);
or UO_1242 (O_1242,N_8010,N_8358);
nor UO_1243 (O_1243,N_7992,N_9601);
xnor UO_1244 (O_1244,N_8608,N_9096);
or UO_1245 (O_1245,N_8785,N_9268);
or UO_1246 (O_1246,N_9994,N_7694);
or UO_1247 (O_1247,N_9313,N_8708);
nor UO_1248 (O_1248,N_9170,N_9939);
and UO_1249 (O_1249,N_7557,N_9289);
nand UO_1250 (O_1250,N_8140,N_8019);
or UO_1251 (O_1251,N_8016,N_8738);
xor UO_1252 (O_1252,N_7757,N_7651);
or UO_1253 (O_1253,N_7990,N_8591);
nor UO_1254 (O_1254,N_9068,N_8594);
or UO_1255 (O_1255,N_9993,N_9229);
nor UO_1256 (O_1256,N_9769,N_7553);
or UO_1257 (O_1257,N_8509,N_9524);
nor UO_1258 (O_1258,N_8348,N_9153);
and UO_1259 (O_1259,N_9886,N_8458);
nand UO_1260 (O_1260,N_9803,N_9482);
nand UO_1261 (O_1261,N_8700,N_9525);
nand UO_1262 (O_1262,N_9859,N_8900);
or UO_1263 (O_1263,N_8082,N_7654);
or UO_1264 (O_1264,N_7691,N_8076);
or UO_1265 (O_1265,N_8781,N_7694);
xnor UO_1266 (O_1266,N_8874,N_9708);
and UO_1267 (O_1267,N_8628,N_9807);
nand UO_1268 (O_1268,N_8138,N_9037);
nor UO_1269 (O_1269,N_8810,N_8650);
nor UO_1270 (O_1270,N_9594,N_8136);
nand UO_1271 (O_1271,N_9013,N_8030);
or UO_1272 (O_1272,N_7790,N_8076);
and UO_1273 (O_1273,N_8668,N_8380);
nor UO_1274 (O_1274,N_9190,N_7928);
nor UO_1275 (O_1275,N_7655,N_9937);
nor UO_1276 (O_1276,N_9548,N_8062);
and UO_1277 (O_1277,N_8734,N_9581);
xor UO_1278 (O_1278,N_9150,N_9935);
nor UO_1279 (O_1279,N_7573,N_9804);
nand UO_1280 (O_1280,N_8905,N_8514);
or UO_1281 (O_1281,N_8207,N_7832);
and UO_1282 (O_1282,N_9346,N_9506);
nand UO_1283 (O_1283,N_7548,N_8558);
nor UO_1284 (O_1284,N_7630,N_9677);
and UO_1285 (O_1285,N_9451,N_8270);
nand UO_1286 (O_1286,N_8545,N_9628);
or UO_1287 (O_1287,N_9766,N_8553);
or UO_1288 (O_1288,N_9138,N_9016);
nand UO_1289 (O_1289,N_8368,N_7595);
nand UO_1290 (O_1290,N_7847,N_8422);
nand UO_1291 (O_1291,N_8224,N_8943);
and UO_1292 (O_1292,N_7563,N_9849);
and UO_1293 (O_1293,N_8740,N_9494);
or UO_1294 (O_1294,N_9300,N_8289);
or UO_1295 (O_1295,N_7611,N_8419);
xnor UO_1296 (O_1296,N_7889,N_7891);
nand UO_1297 (O_1297,N_9217,N_7508);
or UO_1298 (O_1298,N_9987,N_8344);
and UO_1299 (O_1299,N_8848,N_9829);
and UO_1300 (O_1300,N_9260,N_7657);
and UO_1301 (O_1301,N_9283,N_8165);
xnor UO_1302 (O_1302,N_8026,N_8989);
and UO_1303 (O_1303,N_8959,N_9387);
and UO_1304 (O_1304,N_9118,N_8676);
or UO_1305 (O_1305,N_8267,N_7702);
nand UO_1306 (O_1306,N_8080,N_9883);
or UO_1307 (O_1307,N_8317,N_7758);
nor UO_1308 (O_1308,N_7783,N_8502);
or UO_1309 (O_1309,N_8531,N_9963);
and UO_1310 (O_1310,N_9347,N_9014);
nand UO_1311 (O_1311,N_7816,N_8596);
nor UO_1312 (O_1312,N_7813,N_8793);
or UO_1313 (O_1313,N_9817,N_9897);
or UO_1314 (O_1314,N_8304,N_9956);
and UO_1315 (O_1315,N_9690,N_8111);
nand UO_1316 (O_1316,N_9172,N_9330);
nand UO_1317 (O_1317,N_8524,N_7766);
nand UO_1318 (O_1318,N_7667,N_7814);
or UO_1319 (O_1319,N_7753,N_9563);
nor UO_1320 (O_1320,N_9591,N_9902);
or UO_1321 (O_1321,N_9249,N_9837);
or UO_1322 (O_1322,N_8480,N_8089);
nand UO_1323 (O_1323,N_8469,N_9738);
nand UO_1324 (O_1324,N_7841,N_9742);
nand UO_1325 (O_1325,N_9121,N_7622);
nor UO_1326 (O_1326,N_8034,N_9108);
and UO_1327 (O_1327,N_9780,N_9960);
nand UO_1328 (O_1328,N_7670,N_9010);
nor UO_1329 (O_1329,N_9503,N_7859);
xnor UO_1330 (O_1330,N_7632,N_8446);
nand UO_1331 (O_1331,N_8531,N_8377);
nand UO_1332 (O_1332,N_7843,N_8428);
nand UO_1333 (O_1333,N_8508,N_8315);
and UO_1334 (O_1334,N_9635,N_7515);
nor UO_1335 (O_1335,N_9078,N_7774);
or UO_1336 (O_1336,N_9683,N_8586);
xnor UO_1337 (O_1337,N_7672,N_8012);
nor UO_1338 (O_1338,N_9325,N_7942);
and UO_1339 (O_1339,N_9752,N_9232);
nor UO_1340 (O_1340,N_8161,N_8754);
xnor UO_1341 (O_1341,N_9664,N_8418);
and UO_1342 (O_1342,N_8317,N_9463);
nor UO_1343 (O_1343,N_8911,N_8982);
nand UO_1344 (O_1344,N_9948,N_8808);
and UO_1345 (O_1345,N_8501,N_8591);
and UO_1346 (O_1346,N_8928,N_8117);
and UO_1347 (O_1347,N_9074,N_9204);
nor UO_1348 (O_1348,N_8054,N_7777);
xnor UO_1349 (O_1349,N_9512,N_8014);
or UO_1350 (O_1350,N_8779,N_9883);
or UO_1351 (O_1351,N_9026,N_7711);
or UO_1352 (O_1352,N_9332,N_9743);
nor UO_1353 (O_1353,N_8239,N_9747);
nand UO_1354 (O_1354,N_9332,N_9150);
or UO_1355 (O_1355,N_7627,N_8504);
and UO_1356 (O_1356,N_7772,N_9893);
nor UO_1357 (O_1357,N_9208,N_9939);
nand UO_1358 (O_1358,N_9363,N_7705);
nor UO_1359 (O_1359,N_9718,N_7806);
nor UO_1360 (O_1360,N_9054,N_9592);
or UO_1361 (O_1361,N_9639,N_8452);
and UO_1362 (O_1362,N_8909,N_8517);
and UO_1363 (O_1363,N_8814,N_9407);
or UO_1364 (O_1364,N_8292,N_8121);
nor UO_1365 (O_1365,N_8989,N_7706);
nor UO_1366 (O_1366,N_8802,N_9712);
and UO_1367 (O_1367,N_8073,N_9817);
nor UO_1368 (O_1368,N_9823,N_9134);
nand UO_1369 (O_1369,N_7598,N_9939);
or UO_1370 (O_1370,N_8357,N_8945);
nor UO_1371 (O_1371,N_8584,N_7606);
nor UO_1372 (O_1372,N_9293,N_9184);
or UO_1373 (O_1373,N_9037,N_9343);
and UO_1374 (O_1374,N_8019,N_7687);
nand UO_1375 (O_1375,N_8631,N_8117);
nand UO_1376 (O_1376,N_8797,N_9841);
nor UO_1377 (O_1377,N_8495,N_8382);
xor UO_1378 (O_1378,N_9119,N_8325);
nand UO_1379 (O_1379,N_8008,N_9116);
nand UO_1380 (O_1380,N_8747,N_9845);
and UO_1381 (O_1381,N_7757,N_9296);
xnor UO_1382 (O_1382,N_7865,N_9672);
or UO_1383 (O_1383,N_8231,N_9700);
nor UO_1384 (O_1384,N_8669,N_8148);
nand UO_1385 (O_1385,N_9249,N_9303);
and UO_1386 (O_1386,N_8645,N_7649);
and UO_1387 (O_1387,N_8584,N_8340);
nor UO_1388 (O_1388,N_9780,N_9472);
or UO_1389 (O_1389,N_8176,N_9772);
or UO_1390 (O_1390,N_8050,N_7702);
and UO_1391 (O_1391,N_8058,N_9186);
nor UO_1392 (O_1392,N_8084,N_8331);
and UO_1393 (O_1393,N_8858,N_7621);
or UO_1394 (O_1394,N_8539,N_8936);
or UO_1395 (O_1395,N_9349,N_8621);
nor UO_1396 (O_1396,N_9104,N_7655);
and UO_1397 (O_1397,N_8985,N_7869);
nand UO_1398 (O_1398,N_9326,N_9858);
nand UO_1399 (O_1399,N_9846,N_7862);
xor UO_1400 (O_1400,N_9797,N_8704);
nand UO_1401 (O_1401,N_8170,N_9146);
and UO_1402 (O_1402,N_8091,N_7826);
nor UO_1403 (O_1403,N_9109,N_8678);
nor UO_1404 (O_1404,N_9153,N_7666);
nand UO_1405 (O_1405,N_8077,N_9411);
nor UO_1406 (O_1406,N_7614,N_7670);
and UO_1407 (O_1407,N_9875,N_7526);
and UO_1408 (O_1408,N_7565,N_9218);
nand UO_1409 (O_1409,N_9503,N_7613);
nor UO_1410 (O_1410,N_9445,N_9645);
or UO_1411 (O_1411,N_7861,N_9348);
or UO_1412 (O_1412,N_8131,N_9144);
or UO_1413 (O_1413,N_8434,N_8781);
or UO_1414 (O_1414,N_8224,N_8915);
and UO_1415 (O_1415,N_9348,N_8912);
nand UO_1416 (O_1416,N_9772,N_9744);
or UO_1417 (O_1417,N_9166,N_9151);
or UO_1418 (O_1418,N_8617,N_7807);
and UO_1419 (O_1419,N_8839,N_9873);
nor UO_1420 (O_1420,N_9571,N_8951);
nor UO_1421 (O_1421,N_9822,N_9334);
and UO_1422 (O_1422,N_9893,N_9889);
and UO_1423 (O_1423,N_9994,N_8814);
and UO_1424 (O_1424,N_9879,N_9268);
and UO_1425 (O_1425,N_8033,N_9710);
or UO_1426 (O_1426,N_8445,N_7862);
and UO_1427 (O_1427,N_8497,N_8245);
xnor UO_1428 (O_1428,N_9300,N_9373);
and UO_1429 (O_1429,N_8889,N_8514);
nor UO_1430 (O_1430,N_8144,N_7930);
and UO_1431 (O_1431,N_9126,N_7601);
and UO_1432 (O_1432,N_7878,N_7525);
or UO_1433 (O_1433,N_9749,N_8327);
xnor UO_1434 (O_1434,N_8557,N_8907);
and UO_1435 (O_1435,N_8950,N_9287);
nor UO_1436 (O_1436,N_7870,N_9590);
nor UO_1437 (O_1437,N_9545,N_8707);
nand UO_1438 (O_1438,N_9369,N_8371);
and UO_1439 (O_1439,N_8501,N_7875);
or UO_1440 (O_1440,N_8674,N_7658);
nor UO_1441 (O_1441,N_9787,N_9580);
nand UO_1442 (O_1442,N_9565,N_7813);
nor UO_1443 (O_1443,N_9490,N_9299);
and UO_1444 (O_1444,N_9151,N_8108);
and UO_1445 (O_1445,N_9234,N_8429);
and UO_1446 (O_1446,N_9726,N_7846);
nand UO_1447 (O_1447,N_7695,N_8921);
nor UO_1448 (O_1448,N_8111,N_7606);
nand UO_1449 (O_1449,N_9894,N_7802);
and UO_1450 (O_1450,N_8461,N_7611);
xor UO_1451 (O_1451,N_9094,N_9160);
or UO_1452 (O_1452,N_8935,N_9714);
or UO_1453 (O_1453,N_8359,N_9821);
nor UO_1454 (O_1454,N_8526,N_9130);
or UO_1455 (O_1455,N_8605,N_9647);
nand UO_1456 (O_1456,N_9115,N_9692);
nand UO_1457 (O_1457,N_9543,N_8057);
and UO_1458 (O_1458,N_9245,N_9472);
and UO_1459 (O_1459,N_9681,N_8693);
and UO_1460 (O_1460,N_9164,N_9073);
or UO_1461 (O_1461,N_8599,N_9075);
nand UO_1462 (O_1462,N_9366,N_8848);
and UO_1463 (O_1463,N_8494,N_7778);
or UO_1464 (O_1464,N_9874,N_8919);
and UO_1465 (O_1465,N_8669,N_8618);
and UO_1466 (O_1466,N_9745,N_8864);
or UO_1467 (O_1467,N_8132,N_8086);
and UO_1468 (O_1468,N_9579,N_8009);
and UO_1469 (O_1469,N_9529,N_8675);
xnor UO_1470 (O_1470,N_8380,N_8677);
or UO_1471 (O_1471,N_9431,N_7698);
nand UO_1472 (O_1472,N_9530,N_8514);
nand UO_1473 (O_1473,N_8934,N_9894);
and UO_1474 (O_1474,N_8294,N_9902);
or UO_1475 (O_1475,N_8996,N_8662);
nor UO_1476 (O_1476,N_8575,N_8748);
nand UO_1477 (O_1477,N_9762,N_9965);
nand UO_1478 (O_1478,N_9531,N_7565);
nor UO_1479 (O_1479,N_8354,N_9565);
nand UO_1480 (O_1480,N_9331,N_9877);
nand UO_1481 (O_1481,N_8934,N_9214);
nand UO_1482 (O_1482,N_7863,N_9454);
and UO_1483 (O_1483,N_9688,N_8244);
nor UO_1484 (O_1484,N_8594,N_8704);
nor UO_1485 (O_1485,N_9172,N_9740);
nand UO_1486 (O_1486,N_9136,N_8586);
nand UO_1487 (O_1487,N_9828,N_8208);
nand UO_1488 (O_1488,N_8306,N_8708);
and UO_1489 (O_1489,N_8280,N_8072);
or UO_1490 (O_1490,N_9420,N_9148);
and UO_1491 (O_1491,N_8243,N_7883);
and UO_1492 (O_1492,N_8071,N_9196);
xor UO_1493 (O_1493,N_8418,N_7686);
and UO_1494 (O_1494,N_8091,N_7757);
and UO_1495 (O_1495,N_7610,N_8523);
nor UO_1496 (O_1496,N_8939,N_8042);
nor UO_1497 (O_1497,N_9063,N_9064);
nand UO_1498 (O_1498,N_8349,N_8365);
or UO_1499 (O_1499,N_8110,N_9979);
endmodule