module basic_750_5000_1000_5_levels_2xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_116,In_515);
or U1 (N_1,In_675,In_34);
nand U2 (N_2,In_432,In_740);
or U3 (N_3,In_228,In_651);
and U4 (N_4,In_659,In_478);
nand U5 (N_5,In_63,In_237);
or U6 (N_6,In_701,In_229);
nand U7 (N_7,In_136,In_508);
nand U8 (N_8,In_102,In_207);
nor U9 (N_9,In_350,In_367);
nand U10 (N_10,In_224,In_572);
xor U11 (N_11,In_667,In_6);
nand U12 (N_12,In_21,In_568);
nor U13 (N_13,In_528,In_5);
and U14 (N_14,In_520,In_108);
or U15 (N_15,In_337,In_374);
nor U16 (N_16,In_373,In_676);
nor U17 (N_17,In_595,In_735);
or U18 (N_18,In_468,In_385);
nand U19 (N_19,In_444,In_454);
nor U20 (N_20,In_541,In_684);
nand U21 (N_21,In_55,In_377);
nor U22 (N_22,In_637,In_742);
xnor U23 (N_23,In_280,In_214);
and U24 (N_24,In_582,In_142);
nor U25 (N_25,In_268,In_279);
nor U26 (N_26,In_608,In_602);
or U27 (N_27,In_480,In_186);
nand U28 (N_28,In_141,In_704);
and U29 (N_29,In_145,In_386);
nor U30 (N_30,In_714,In_3);
nor U31 (N_31,In_680,In_408);
nor U32 (N_32,In_524,In_8);
and U33 (N_33,In_278,In_571);
nand U34 (N_34,In_435,In_297);
nor U35 (N_35,In_178,In_345);
nor U36 (N_36,In_19,In_401);
nand U37 (N_37,In_149,In_144);
nand U38 (N_38,In_275,In_548);
xnor U39 (N_39,In_677,In_573);
and U40 (N_40,In_222,In_593);
nand U41 (N_41,In_198,In_106);
and U42 (N_42,In_591,In_715);
nand U43 (N_43,In_502,In_316);
or U44 (N_44,In_39,In_580);
or U45 (N_45,In_65,In_673);
or U46 (N_46,In_68,In_653);
or U47 (N_47,In_14,In_15);
nor U48 (N_48,In_99,In_664);
or U49 (N_49,In_220,In_366);
nor U50 (N_50,In_105,In_457);
nor U51 (N_51,In_398,In_351);
xor U52 (N_52,In_327,In_193);
or U53 (N_53,In_630,In_289);
or U54 (N_54,In_211,In_588);
nor U55 (N_55,In_121,In_94);
nor U56 (N_56,In_409,In_447);
and U57 (N_57,In_293,In_183);
nor U58 (N_58,In_309,In_339);
nor U59 (N_59,In_600,In_727);
nand U60 (N_60,In_335,In_217);
nor U61 (N_61,In_197,In_78);
or U62 (N_62,In_380,In_270);
nor U63 (N_63,In_657,In_534);
nand U64 (N_64,In_259,In_705);
or U65 (N_65,In_132,In_394);
nand U66 (N_66,In_721,In_28);
nand U67 (N_67,In_257,In_473);
nand U68 (N_68,In_51,In_395);
or U69 (N_69,In_208,In_305);
nand U70 (N_70,In_470,In_564);
and U71 (N_71,In_689,In_284);
and U72 (N_72,In_707,In_134);
xor U73 (N_73,In_681,In_428);
nor U74 (N_74,In_66,In_11);
nor U75 (N_75,In_513,In_256);
nor U76 (N_76,In_190,In_294);
or U77 (N_77,In_277,In_430);
or U78 (N_78,In_272,In_492);
or U79 (N_79,In_718,In_85);
nor U80 (N_80,In_589,In_267);
and U81 (N_81,In_47,In_494);
nand U82 (N_82,In_682,In_612);
nor U83 (N_83,In_605,In_364);
or U84 (N_84,In_556,In_150);
nand U85 (N_85,In_522,In_459);
nor U86 (N_86,In_362,In_387);
or U87 (N_87,In_590,In_112);
and U88 (N_88,In_20,In_341);
or U89 (N_89,In_52,In_665);
xnor U90 (N_90,In_477,In_89);
nor U91 (N_91,In_746,In_639);
and U92 (N_92,In_210,In_722);
and U93 (N_93,In_739,In_525);
and U94 (N_94,In_647,In_700);
nor U95 (N_95,In_179,In_248);
nand U96 (N_96,In_486,In_361);
and U97 (N_97,In_180,In_295);
nand U98 (N_98,In_536,In_420);
and U99 (N_99,In_230,In_202);
nor U100 (N_100,In_584,In_679);
and U101 (N_101,In_282,In_687);
nand U102 (N_102,In_251,In_227);
nand U103 (N_103,In_97,In_188);
and U104 (N_104,In_54,In_712);
and U105 (N_105,In_660,In_720);
nand U106 (N_106,In_200,In_406);
nand U107 (N_107,In_195,In_96);
nand U108 (N_108,In_192,In_326);
nand U109 (N_109,In_342,In_732);
nand U110 (N_110,In_271,In_532);
nand U111 (N_111,In_196,In_292);
nor U112 (N_112,In_130,In_242);
nor U113 (N_113,In_57,In_38);
and U114 (N_114,In_509,In_472);
nand U115 (N_115,In_446,In_218);
and U116 (N_116,In_453,In_691);
nor U117 (N_117,In_285,In_507);
and U118 (N_118,In_317,In_163);
nand U119 (N_119,In_370,In_244);
nor U120 (N_120,In_191,In_467);
nor U121 (N_121,In_88,In_427);
and U122 (N_122,In_516,In_576);
nor U123 (N_123,In_434,In_119);
or U124 (N_124,In_255,In_231);
and U125 (N_125,In_62,In_656);
nand U126 (N_126,In_79,In_421);
nor U127 (N_127,In_542,In_422);
nor U128 (N_128,In_458,In_128);
or U129 (N_129,In_412,In_450);
nand U130 (N_130,In_349,In_497);
nor U131 (N_131,In_484,In_378);
nor U132 (N_132,In_610,In_734);
and U133 (N_133,In_308,In_464);
or U134 (N_134,In_537,In_719);
and U135 (N_135,In_561,In_565);
xnor U136 (N_136,In_250,In_118);
nor U137 (N_137,In_40,In_109);
and U138 (N_138,In_431,In_76);
nor U139 (N_139,In_694,In_418);
or U140 (N_140,In_114,In_306);
nand U141 (N_141,In_540,In_627);
nor U142 (N_142,In_369,In_417);
nor U143 (N_143,In_262,In_498);
nor U144 (N_144,In_747,In_577);
and U145 (N_145,In_736,In_30);
nand U146 (N_146,In_535,In_510);
nand U147 (N_147,In_304,In_307);
nor U148 (N_148,In_569,In_411);
xor U149 (N_149,In_357,In_60);
xor U150 (N_150,In_617,In_276);
nor U151 (N_151,In_45,In_445);
and U152 (N_152,In_64,In_405);
nor U153 (N_153,In_120,In_153);
or U154 (N_154,In_597,In_113);
and U155 (N_155,In_393,In_201);
nor U156 (N_156,In_671,In_413);
nor U157 (N_157,In_103,In_329);
and U158 (N_158,In_32,In_353);
nand U159 (N_159,In_154,In_33);
or U160 (N_160,In_549,In_529);
and U161 (N_161,In_13,In_171);
and U162 (N_162,In_343,In_92);
nand U163 (N_163,In_669,In_182);
nand U164 (N_164,In_650,In_493);
and U165 (N_165,In_274,In_703);
and U166 (N_166,In_465,In_615);
and U167 (N_167,In_300,In_433);
nand U168 (N_168,In_618,In_189);
or U169 (N_169,In_425,In_455);
and U170 (N_170,In_80,In_501);
or U171 (N_171,In_235,In_688);
xor U172 (N_172,In_567,In_558);
or U173 (N_173,In_607,In_115);
nor U174 (N_174,In_46,In_161);
and U175 (N_175,In_315,In_84);
and U176 (N_176,In_562,In_58);
nand U177 (N_177,In_426,In_613);
or U178 (N_178,In_359,In_392);
xor U179 (N_179,In_402,In_325);
or U180 (N_180,In_290,In_646);
nand U181 (N_181,In_332,In_737);
nand U182 (N_182,In_489,In_539);
and U183 (N_183,In_107,In_616);
and U184 (N_184,In_1,In_466);
nand U185 (N_185,In_555,In_205);
nor U186 (N_186,In_634,In_35);
nand U187 (N_187,In_368,In_546);
and U188 (N_188,In_389,In_519);
nand U189 (N_189,In_530,In_17);
nor U190 (N_190,In_10,In_240);
or U191 (N_191,In_436,In_59);
or U192 (N_192,In_443,In_155);
and U193 (N_193,In_490,In_2);
and U194 (N_194,In_626,In_581);
or U195 (N_195,In_574,In_625);
nor U196 (N_196,In_238,In_655);
and U197 (N_197,In_728,In_12);
nand U198 (N_198,In_662,In_496);
or U199 (N_199,In_129,In_273);
nand U200 (N_200,In_181,In_49);
nor U201 (N_201,In_518,In_169);
nand U202 (N_202,In_358,In_233);
or U203 (N_203,In_643,In_586);
and U204 (N_204,In_438,In_648);
or U205 (N_205,In_745,In_414);
nand U206 (N_206,In_461,In_288);
or U207 (N_207,In_397,In_396);
nor U208 (N_208,In_726,In_744);
nor U209 (N_209,In_437,In_139);
or U210 (N_210,In_566,In_642);
and U211 (N_211,In_286,In_223);
nand U212 (N_212,In_738,In_729);
nor U213 (N_213,In_544,In_24);
or U214 (N_214,In_449,In_506);
or U215 (N_215,In_692,In_283);
nand U216 (N_216,In_624,In_246);
or U217 (N_217,In_649,In_553);
or U218 (N_218,In_174,In_483);
nand U219 (N_219,In_717,In_658);
nand U220 (N_220,In_298,In_254);
nor U221 (N_221,In_514,In_162);
or U222 (N_222,In_448,In_331);
and U223 (N_223,In_206,In_375);
and U224 (N_224,In_72,In_44);
and U225 (N_225,In_697,In_313);
or U226 (N_226,In_451,In_603);
nor U227 (N_227,In_749,In_98);
nand U228 (N_228,In_311,In_41);
nor U229 (N_229,In_654,In_69);
nand U230 (N_230,In_531,In_234);
or U231 (N_231,In_123,In_0);
nand U232 (N_232,In_177,In_140);
or U233 (N_233,In_708,In_7);
nand U234 (N_234,In_243,In_560);
nor U235 (N_235,In_124,In_594);
and U236 (N_236,In_239,In_138);
or U237 (N_237,In_638,In_158);
nand U238 (N_238,In_400,In_71);
or U239 (N_239,In_706,In_301);
and U240 (N_240,In_670,In_61);
and U241 (N_241,In_173,In_87);
nor U242 (N_242,In_199,In_503);
nand U243 (N_243,In_668,In_724);
or U244 (N_244,In_381,In_632);
nand U245 (N_245,In_748,In_81);
or U246 (N_246,In_609,In_159);
nor U247 (N_247,In_347,In_22);
and U248 (N_248,In_252,In_212);
nor U249 (N_249,In_156,In_312);
or U250 (N_250,In_379,In_133);
nand U251 (N_251,In_194,In_187);
xor U252 (N_252,In_499,In_82);
or U253 (N_253,In_557,In_716);
nor U254 (N_254,In_695,In_570);
and U255 (N_255,In_334,In_419);
nand U256 (N_256,In_631,In_559);
nor U257 (N_257,In_391,In_296);
nor U258 (N_258,In_723,In_117);
or U259 (N_259,In_629,In_338);
or U260 (N_260,In_340,In_587);
nor U261 (N_261,In_151,In_476);
nor U262 (N_262,In_265,In_482);
and U263 (N_263,In_487,In_403);
nor U264 (N_264,In_314,In_456);
nor U265 (N_265,In_672,In_176);
or U266 (N_266,In_622,In_384);
nor U267 (N_267,In_441,In_491);
nand U268 (N_268,In_31,In_215);
nand U269 (N_269,In_640,In_416);
or U270 (N_270,In_690,In_382);
and U271 (N_271,In_26,In_376);
or U272 (N_272,In_731,In_336);
nand U273 (N_273,In_526,In_462);
nor U274 (N_274,In_371,In_563);
and U275 (N_275,In_299,In_172);
nor U276 (N_276,In_77,In_505);
nand U277 (N_277,In_481,In_203);
nor U278 (N_278,In_42,In_4);
nor U279 (N_279,In_75,In_209);
or U280 (N_280,In_148,In_641);
nor U281 (N_281,In_137,In_152);
nor U282 (N_282,In_628,In_365);
xor U283 (N_283,In_175,In_710);
nand U284 (N_284,In_439,In_696);
nor U285 (N_285,In_527,In_551);
and U286 (N_286,In_48,In_111);
or U287 (N_287,In_166,In_330);
or U288 (N_288,In_598,In_266);
or U289 (N_289,In_23,In_56);
nand U290 (N_290,In_533,In_249);
nand U291 (N_291,In_644,In_488);
and U292 (N_292,In_43,In_698);
nand U293 (N_293,In_523,In_545);
nor U294 (N_294,In_471,In_683);
or U295 (N_295,In_310,In_575);
or U296 (N_296,In_550,In_404);
nand U297 (N_297,In_50,In_424);
nand U298 (N_298,In_604,In_101);
and U299 (N_299,In_320,In_185);
nor U300 (N_300,In_463,In_543);
nand U301 (N_301,In_596,In_583);
nor U302 (N_302,In_410,In_674);
nand U303 (N_303,In_360,In_167);
and U304 (N_304,In_538,In_164);
nand U305 (N_305,In_291,In_143);
nor U306 (N_306,In_552,In_500);
or U307 (N_307,In_29,In_429);
nor U308 (N_308,In_678,In_614);
nor U309 (N_309,In_474,In_216);
nand U310 (N_310,In_355,In_620);
nand U311 (N_311,In_611,In_170);
nand U312 (N_312,In_319,In_460);
and U313 (N_313,In_372,In_127);
or U314 (N_314,In_323,In_36);
xor U315 (N_315,In_475,In_599);
nor U316 (N_316,In_352,In_247);
and U317 (N_317,In_328,In_585);
or U318 (N_318,In_16,In_741);
or U319 (N_319,In_93,In_383);
and U320 (N_320,In_390,In_90);
nor U321 (N_321,In_236,In_303);
nand U322 (N_322,In_226,In_713);
nand U323 (N_323,In_184,In_318);
and U324 (N_324,In_53,In_100);
nor U325 (N_325,In_86,In_407);
or U326 (N_326,In_709,In_733);
or U327 (N_327,In_363,In_452);
nand U328 (N_328,In_693,In_725);
nand U329 (N_329,In_423,In_122);
nor U330 (N_330,In_521,In_324);
or U331 (N_331,In_495,In_666);
nand U332 (N_332,In_601,In_225);
and U333 (N_333,In_440,In_287);
or U334 (N_334,In_346,In_554);
nand U335 (N_335,In_579,In_606);
or U336 (N_336,In_442,In_415);
or U337 (N_337,In_469,In_110);
nor U338 (N_338,In_74,In_104);
and U339 (N_339,In_241,In_135);
and U340 (N_340,In_633,In_623);
nand U341 (N_341,In_348,In_232);
or U342 (N_342,In_302,In_9);
or U343 (N_343,In_27,In_204);
nand U344 (N_344,In_711,In_125);
or U345 (N_345,In_73,In_333);
or U346 (N_346,In_621,In_663);
or U347 (N_347,In_258,In_322);
nor U348 (N_348,In_504,In_264);
and U349 (N_349,In_479,In_321);
nand U350 (N_350,In_95,In_685);
or U351 (N_351,In_147,In_126);
or U352 (N_352,In_356,In_743);
nor U353 (N_353,In_399,In_619);
and U354 (N_354,In_91,In_592);
nand U355 (N_355,In_260,In_636);
and U356 (N_356,In_635,In_686);
nand U357 (N_357,In_37,In_165);
and U358 (N_358,In_221,In_511);
nand U359 (N_359,In_146,In_485);
nand U360 (N_360,In_344,In_730);
nand U361 (N_361,In_67,In_168);
and U362 (N_362,In_645,In_652);
and U363 (N_363,In_25,In_269);
or U364 (N_364,In_699,In_219);
nand U365 (N_365,In_547,In_245);
and U366 (N_366,In_70,In_388);
nor U367 (N_367,In_261,In_83);
and U368 (N_368,In_578,In_263);
or U369 (N_369,In_18,In_157);
nor U370 (N_370,In_702,In_253);
nand U371 (N_371,In_517,In_213);
nand U372 (N_372,In_354,In_281);
or U373 (N_373,In_160,In_131);
and U374 (N_374,In_512,In_661);
and U375 (N_375,In_386,In_508);
or U376 (N_376,In_583,In_409);
nor U377 (N_377,In_360,In_213);
and U378 (N_378,In_107,In_233);
or U379 (N_379,In_497,In_453);
nand U380 (N_380,In_158,In_462);
nand U381 (N_381,In_673,In_227);
or U382 (N_382,In_407,In_74);
nor U383 (N_383,In_498,In_696);
and U384 (N_384,In_466,In_355);
xnor U385 (N_385,In_179,In_611);
or U386 (N_386,In_546,In_63);
and U387 (N_387,In_115,In_404);
nand U388 (N_388,In_114,In_633);
and U389 (N_389,In_288,In_534);
nor U390 (N_390,In_663,In_300);
nand U391 (N_391,In_135,In_454);
xor U392 (N_392,In_734,In_484);
nand U393 (N_393,In_238,In_143);
nand U394 (N_394,In_469,In_318);
and U395 (N_395,In_686,In_665);
nor U396 (N_396,In_567,In_323);
or U397 (N_397,In_188,In_516);
or U398 (N_398,In_11,In_329);
nor U399 (N_399,In_341,In_185);
and U400 (N_400,In_277,In_383);
nand U401 (N_401,In_165,In_374);
or U402 (N_402,In_625,In_109);
nand U403 (N_403,In_481,In_618);
and U404 (N_404,In_57,In_459);
nor U405 (N_405,In_191,In_309);
nand U406 (N_406,In_310,In_405);
and U407 (N_407,In_627,In_14);
nand U408 (N_408,In_439,In_588);
nor U409 (N_409,In_257,In_290);
nor U410 (N_410,In_409,In_510);
nand U411 (N_411,In_599,In_33);
nor U412 (N_412,In_209,In_628);
nor U413 (N_413,In_699,In_321);
and U414 (N_414,In_277,In_147);
and U415 (N_415,In_633,In_430);
nor U416 (N_416,In_566,In_749);
and U417 (N_417,In_467,In_126);
or U418 (N_418,In_41,In_335);
or U419 (N_419,In_397,In_474);
nand U420 (N_420,In_141,In_577);
nor U421 (N_421,In_13,In_75);
nand U422 (N_422,In_563,In_288);
nor U423 (N_423,In_419,In_445);
nand U424 (N_424,In_20,In_158);
or U425 (N_425,In_480,In_483);
nor U426 (N_426,In_275,In_206);
nor U427 (N_427,In_666,In_581);
xor U428 (N_428,In_429,In_57);
nor U429 (N_429,In_287,In_386);
xor U430 (N_430,In_521,In_441);
or U431 (N_431,In_732,In_596);
nand U432 (N_432,In_182,In_32);
and U433 (N_433,In_299,In_225);
or U434 (N_434,In_661,In_421);
or U435 (N_435,In_102,In_273);
and U436 (N_436,In_362,In_439);
xnor U437 (N_437,In_367,In_706);
nor U438 (N_438,In_216,In_714);
nor U439 (N_439,In_132,In_242);
and U440 (N_440,In_49,In_338);
and U441 (N_441,In_608,In_176);
or U442 (N_442,In_481,In_556);
nor U443 (N_443,In_157,In_420);
nand U444 (N_444,In_734,In_723);
and U445 (N_445,In_657,In_283);
nand U446 (N_446,In_217,In_583);
and U447 (N_447,In_511,In_167);
nand U448 (N_448,In_553,In_334);
and U449 (N_449,In_167,In_327);
nor U450 (N_450,In_242,In_568);
or U451 (N_451,In_713,In_32);
nor U452 (N_452,In_713,In_112);
nand U453 (N_453,In_280,In_133);
or U454 (N_454,In_185,In_572);
and U455 (N_455,In_118,In_386);
or U456 (N_456,In_184,In_183);
and U457 (N_457,In_384,In_279);
xnor U458 (N_458,In_693,In_426);
and U459 (N_459,In_212,In_238);
and U460 (N_460,In_714,In_368);
nor U461 (N_461,In_11,In_472);
or U462 (N_462,In_229,In_7);
nand U463 (N_463,In_594,In_426);
nand U464 (N_464,In_489,In_5);
and U465 (N_465,In_33,In_292);
nor U466 (N_466,In_726,In_570);
and U467 (N_467,In_292,In_217);
nand U468 (N_468,In_387,In_635);
nor U469 (N_469,In_338,In_726);
nor U470 (N_470,In_31,In_319);
nor U471 (N_471,In_749,In_643);
or U472 (N_472,In_238,In_522);
nand U473 (N_473,In_415,In_115);
or U474 (N_474,In_511,In_626);
nand U475 (N_475,In_420,In_451);
or U476 (N_476,In_424,In_201);
nor U477 (N_477,In_116,In_490);
and U478 (N_478,In_42,In_330);
or U479 (N_479,In_545,In_167);
nor U480 (N_480,In_686,In_599);
nand U481 (N_481,In_295,In_445);
nor U482 (N_482,In_526,In_3);
or U483 (N_483,In_85,In_483);
nor U484 (N_484,In_418,In_126);
and U485 (N_485,In_427,In_650);
nor U486 (N_486,In_382,In_417);
and U487 (N_487,In_337,In_694);
and U488 (N_488,In_355,In_618);
nand U489 (N_489,In_614,In_441);
or U490 (N_490,In_354,In_276);
nand U491 (N_491,In_252,In_418);
xor U492 (N_492,In_216,In_612);
nor U493 (N_493,In_481,In_448);
nor U494 (N_494,In_657,In_417);
or U495 (N_495,In_83,In_189);
and U496 (N_496,In_18,In_514);
and U497 (N_497,In_587,In_671);
nor U498 (N_498,In_368,In_260);
nor U499 (N_499,In_311,In_156);
nand U500 (N_500,In_235,In_207);
or U501 (N_501,In_232,In_431);
and U502 (N_502,In_479,In_711);
nor U503 (N_503,In_445,In_183);
nand U504 (N_504,In_597,In_680);
and U505 (N_505,In_389,In_473);
or U506 (N_506,In_24,In_135);
or U507 (N_507,In_251,In_446);
or U508 (N_508,In_179,In_263);
or U509 (N_509,In_350,In_569);
or U510 (N_510,In_615,In_121);
and U511 (N_511,In_354,In_696);
nor U512 (N_512,In_510,In_517);
and U513 (N_513,In_563,In_20);
nand U514 (N_514,In_309,In_184);
nor U515 (N_515,In_531,In_461);
or U516 (N_516,In_148,In_125);
or U517 (N_517,In_305,In_231);
nor U518 (N_518,In_479,In_554);
nand U519 (N_519,In_708,In_212);
nand U520 (N_520,In_67,In_657);
and U521 (N_521,In_390,In_666);
and U522 (N_522,In_416,In_323);
and U523 (N_523,In_698,In_412);
nand U524 (N_524,In_418,In_542);
nand U525 (N_525,In_418,In_688);
nand U526 (N_526,In_415,In_637);
or U527 (N_527,In_721,In_361);
nand U528 (N_528,In_493,In_568);
nor U529 (N_529,In_518,In_468);
nor U530 (N_530,In_44,In_540);
or U531 (N_531,In_603,In_718);
or U532 (N_532,In_701,In_231);
nor U533 (N_533,In_287,In_555);
and U534 (N_534,In_72,In_365);
or U535 (N_535,In_502,In_618);
nor U536 (N_536,In_58,In_534);
nand U537 (N_537,In_250,In_653);
nor U538 (N_538,In_525,In_472);
and U539 (N_539,In_746,In_748);
or U540 (N_540,In_35,In_123);
xnor U541 (N_541,In_591,In_204);
nor U542 (N_542,In_17,In_322);
nor U543 (N_543,In_365,In_542);
and U544 (N_544,In_601,In_616);
nand U545 (N_545,In_129,In_188);
or U546 (N_546,In_50,In_630);
nand U547 (N_547,In_440,In_618);
nand U548 (N_548,In_301,In_684);
nand U549 (N_549,In_254,In_102);
nand U550 (N_550,In_497,In_455);
xor U551 (N_551,In_721,In_427);
xor U552 (N_552,In_54,In_637);
and U553 (N_553,In_568,In_267);
nand U554 (N_554,In_42,In_333);
nor U555 (N_555,In_147,In_67);
nor U556 (N_556,In_416,In_101);
nand U557 (N_557,In_324,In_229);
nand U558 (N_558,In_442,In_693);
nand U559 (N_559,In_31,In_576);
nor U560 (N_560,In_164,In_606);
or U561 (N_561,In_169,In_570);
or U562 (N_562,In_388,In_72);
or U563 (N_563,In_681,In_492);
nor U564 (N_564,In_11,In_479);
or U565 (N_565,In_109,In_741);
and U566 (N_566,In_704,In_444);
nor U567 (N_567,In_583,In_711);
and U568 (N_568,In_406,In_701);
nor U569 (N_569,In_21,In_610);
nand U570 (N_570,In_639,In_452);
nand U571 (N_571,In_716,In_71);
xnor U572 (N_572,In_736,In_252);
or U573 (N_573,In_408,In_715);
or U574 (N_574,In_71,In_299);
nor U575 (N_575,In_624,In_292);
or U576 (N_576,In_471,In_566);
or U577 (N_577,In_16,In_205);
and U578 (N_578,In_660,In_308);
or U579 (N_579,In_498,In_40);
nor U580 (N_580,In_670,In_117);
nor U581 (N_581,In_460,In_163);
and U582 (N_582,In_138,In_574);
nand U583 (N_583,In_67,In_539);
and U584 (N_584,In_17,In_263);
nand U585 (N_585,In_538,In_269);
and U586 (N_586,In_92,In_596);
or U587 (N_587,In_688,In_469);
nand U588 (N_588,In_28,In_511);
or U589 (N_589,In_56,In_680);
and U590 (N_590,In_554,In_695);
nand U591 (N_591,In_458,In_699);
nand U592 (N_592,In_427,In_475);
and U593 (N_593,In_646,In_444);
and U594 (N_594,In_89,In_698);
nor U595 (N_595,In_513,In_209);
nand U596 (N_596,In_41,In_568);
and U597 (N_597,In_231,In_222);
and U598 (N_598,In_524,In_138);
nand U599 (N_599,In_400,In_136);
and U600 (N_600,In_300,In_16);
nor U601 (N_601,In_84,In_747);
nor U602 (N_602,In_278,In_518);
or U603 (N_603,In_384,In_377);
or U604 (N_604,In_590,In_182);
nand U605 (N_605,In_83,In_195);
and U606 (N_606,In_182,In_316);
xor U607 (N_607,In_427,In_737);
nand U608 (N_608,In_659,In_503);
nor U609 (N_609,In_422,In_231);
nand U610 (N_610,In_480,In_524);
nor U611 (N_611,In_422,In_289);
nor U612 (N_612,In_656,In_640);
and U613 (N_613,In_558,In_605);
xnor U614 (N_614,In_649,In_745);
nand U615 (N_615,In_375,In_347);
nor U616 (N_616,In_575,In_177);
nand U617 (N_617,In_613,In_427);
nor U618 (N_618,In_289,In_570);
nand U619 (N_619,In_453,In_43);
nand U620 (N_620,In_483,In_146);
and U621 (N_621,In_714,In_167);
nand U622 (N_622,In_432,In_116);
or U623 (N_623,In_582,In_647);
and U624 (N_624,In_157,In_620);
or U625 (N_625,In_560,In_500);
nor U626 (N_626,In_416,In_143);
nand U627 (N_627,In_578,In_17);
and U628 (N_628,In_56,In_705);
nand U629 (N_629,In_237,In_310);
nor U630 (N_630,In_321,In_654);
nand U631 (N_631,In_199,In_276);
xnor U632 (N_632,In_201,In_561);
and U633 (N_633,In_309,In_134);
or U634 (N_634,In_383,In_22);
and U635 (N_635,In_484,In_18);
nand U636 (N_636,In_436,In_722);
and U637 (N_637,In_700,In_191);
nand U638 (N_638,In_665,In_469);
or U639 (N_639,In_656,In_401);
nor U640 (N_640,In_251,In_176);
nand U641 (N_641,In_567,In_534);
or U642 (N_642,In_45,In_370);
or U643 (N_643,In_741,In_614);
nand U644 (N_644,In_56,In_217);
and U645 (N_645,In_609,In_723);
and U646 (N_646,In_703,In_153);
and U647 (N_647,In_36,In_457);
nand U648 (N_648,In_220,In_170);
and U649 (N_649,In_535,In_346);
xor U650 (N_650,In_349,In_550);
nand U651 (N_651,In_672,In_318);
nor U652 (N_652,In_603,In_622);
or U653 (N_653,In_468,In_489);
nor U654 (N_654,In_255,In_317);
and U655 (N_655,In_660,In_344);
nand U656 (N_656,In_397,In_383);
nor U657 (N_657,In_242,In_450);
nand U658 (N_658,In_476,In_434);
nand U659 (N_659,In_621,In_438);
and U660 (N_660,In_533,In_564);
nand U661 (N_661,In_264,In_223);
nor U662 (N_662,In_164,In_110);
xnor U663 (N_663,In_714,In_267);
and U664 (N_664,In_414,In_202);
nor U665 (N_665,In_95,In_466);
and U666 (N_666,In_305,In_562);
and U667 (N_667,In_104,In_18);
nand U668 (N_668,In_77,In_668);
and U669 (N_669,In_377,In_357);
nand U670 (N_670,In_282,In_122);
nor U671 (N_671,In_740,In_464);
nor U672 (N_672,In_284,In_25);
and U673 (N_673,In_173,In_665);
nand U674 (N_674,In_580,In_366);
or U675 (N_675,In_73,In_707);
or U676 (N_676,In_538,In_169);
or U677 (N_677,In_9,In_555);
nand U678 (N_678,In_337,In_28);
nor U679 (N_679,In_499,In_483);
or U680 (N_680,In_102,In_368);
and U681 (N_681,In_451,In_219);
and U682 (N_682,In_704,In_710);
or U683 (N_683,In_288,In_539);
nor U684 (N_684,In_31,In_129);
and U685 (N_685,In_446,In_587);
nand U686 (N_686,In_184,In_23);
nand U687 (N_687,In_331,In_447);
and U688 (N_688,In_532,In_429);
nand U689 (N_689,In_137,In_572);
nand U690 (N_690,In_348,In_504);
or U691 (N_691,In_159,In_405);
nand U692 (N_692,In_304,In_325);
nor U693 (N_693,In_480,In_601);
nor U694 (N_694,In_376,In_539);
and U695 (N_695,In_351,In_509);
or U696 (N_696,In_437,In_34);
and U697 (N_697,In_731,In_558);
xnor U698 (N_698,In_413,In_281);
and U699 (N_699,In_517,In_329);
and U700 (N_700,In_230,In_204);
nor U701 (N_701,In_695,In_265);
and U702 (N_702,In_212,In_363);
or U703 (N_703,In_711,In_171);
nor U704 (N_704,In_501,In_500);
xnor U705 (N_705,In_138,In_718);
nand U706 (N_706,In_472,In_228);
nand U707 (N_707,In_467,In_344);
nor U708 (N_708,In_660,In_459);
nor U709 (N_709,In_745,In_278);
and U710 (N_710,In_694,In_220);
or U711 (N_711,In_291,In_729);
and U712 (N_712,In_227,In_88);
nand U713 (N_713,In_635,In_507);
or U714 (N_714,In_575,In_55);
or U715 (N_715,In_4,In_287);
or U716 (N_716,In_346,In_186);
nand U717 (N_717,In_395,In_705);
nor U718 (N_718,In_343,In_142);
nand U719 (N_719,In_476,In_737);
nor U720 (N_720,In_7,In_666);
nor U721 (N_721,In_69,In_304);
or U722 (N_722,In_261,In_607);
nand U723 (N_723,In_328,In_276);
or U724 (N_724,In_111,In_2);
xor U725 (N_725,In_661,In_518);
and U726 (N_726,In_393,In_264);
nor U727 (N_727,In_5,In_720);
nor U728 (N_728,In_499,In_263);
or U729 (N_729,In_617,In_365);
or U730 (N_730,In_565,In_28);
and U731 (N_731,In_256,In_45);
or U732 (N_732,In_178,In_387);
nand U733 (N_733,In_328,In_633);
nor U734 (N_734,In_458,In_679);
nand U735 (N_735,In_586,In_557);
nor U736 (N_736,In_322,In_182);
and U737 (N_737,In_570,In_468);
nand U738 (N_738,In_709,In_643);
or U739 (N_739,In_311,In_592);
nor U740 (N_740,In_572,In_324);
or U741 (N_741,In_655,In_511);
nor U742 (N_742,In_393,In_555);
nand U743 (N_743,In_730,In_127);
nand U744 (N_744,In_107,In_573);
nor U745 (N_745,In_255,In_351);
nor U746 (N_746,In_626,In_125);
or U747 (N_747,In_335,In_145);
nor U748 (N_748,In_57,In_725);
or U749 (N_749,In_391,In_339);
nor U750 (N_750,In_716,In_270);
or U751 (N_751,In_696,In_670);
and U752 (N_752,In_130,In_55);
nor U753 (N_753,In_637,In_126);
and U754 (N_754,In_283,In_480);
nand U755 (N_755,In_37,In_195);
nand U756 (N_756,In_101,In_611);
nand U757 (N_757,In_694,In_639);
or U758 (N_758,In_576,In_727);
nor U759 (N_759,In_435,In_205);
nand U760 (N_760,In_175,In_662);
nand U761 (N_761,In_70,In_197);
nand U762 (N_762,In_511,In_126);
nor U763 (N_763,In_501,In_452);
nand U764 (N_764,In_729,In_243);
nand U765 (N_765,In_390,In_278);
and U766 (N_766,In_528,In_178);
or U767 (N_767,In_106,In_585);
nand U768 (N_768,In_96,In_704);
nor U769 (N_769,In_383,In_310);
or U770 (N_770,In_128,In_89);
nor U771 (N_771,In_141,In_156);
or U772 (N_772,In_223,In_631);
nor U773 (N_773,In_76,In_234);
or U774 (N_774,In_414,In_87);
nand U775 (N_775,In_265,In_253);
or U776 (N_776,In_547,In_584);
nor U777 (N_777,In_530,In_570);
or U778 (N_778,In_17,In_501);
nand U779 (N_779,In_5,In_373);
and U780 (N_780,In_1,In_486);
nor U781 (N_781,In_283,In_727);
nand U782 (N_782,In_18,In_203);
nor U783 (N_783,In_332,In_562);
nor U784 (N_784,In_119,In_343);
nand U785 (N_785,In_575,In_632);
nand U786 (N_786,In_131,In_96);
and U787 (N_787,In_433,In_227);
or U788 (N_788,In_721,In_157);
or U789 (N_789,In_167,In_465);
or U790 (N_790,In_201,In_258);
nor U791 (N_791,In_638,In_614);
or U792 (N_792,In_677,In_334);
and U793 (N_793,In_23,In_472);
nand U794 (N_794,In_419,In_173);
and U795 (N_795,In_95,In_364);
or U796 (N_796,In_199,In_140);
nor U797 (N_797,In_429,In_175);
nand U798 (N_798,In_116,In_616);
nand U799 (N_799,In_438,In_29);
nor U800 (N_800,In_628,In_394);
nand U801 (N_801,In_730,In_238);
or U802 (N_802,In_602,In_252);
and U803 (N_803,In_247,In_37);
nor U804 (N_804,In_380,In_319);
or U805 (N_805,In_415,In_673);
and U806 (N_806,In_92,In_522);
nor U807 (N_807,In_160,In_107);
nand U808 (N_808,In_170,In_594);
or U809 (N_809,In_78,In_710);
and U810 (N_810,In_302,In_474);
and U811 (N_811,In_102,In_360);
nor U812 (N_812,In_741,In_434);
or U813 (N_813,In_490,In_241);
nor U814 (N_814,In_529,In_14);
or U815 (N_815,In_411,In_377);
nand U816 (N_816,In_76,In_251);
and U817 (N_817,In_338,In_749);
nand U818 (N_818,In_533,In_5);
and U819 (N_819,In_304,In_649);
or U820 (N_820,In_623,In_710);
nor U821 (N_821,In_537,In_594);
and U822 (N_822,In_159,In_615);
and U823 (N_823,In_109,In_364);
or U824 (N_824,In_696,In_6);
nor U825 (N_825,In_238,In_211);
or U826 (N_826,In_239,In_314);
nand U827 (N_827,In_305,In_408);
and U828 (N_828,In_706,In_203);
nor U829 (N_829,In_743,In_212);
nand U830 (N_830,In_577,In_726);
or U831 (N_831,In_467,In_327);
nand U832 (N_832,In_741,In_245);
nor U833 (N_833,In_716,In_691);
nand U834 (N_834,In_446,In_508);
or U835 (N_835,In_677,In_628);
or U836 (N_836,In_203,In_480);
nand U837 (N_837,In_598,In_391);
and U838 (N_838,In_318,In_65);
nand U839 (N_839,In_601,In_286);
or U840 (N_840,In_246,In_550);
nor U841 (N_841,In_598,In_625);
or U842 (N_842,In_252,In_748);
or U843 (N_843,In_303,In_108);
nand U844 (N_844,In_552,In_112);
nor U845 (N_845,In_397,In_376);
or U846 (N_846,In_344,In_722);
and U847 (N_847,In_199,In_518);
and U848 (N_848,In_368,In_261);
nand U849 (N_849,In_260,In_608);
nor U850 (N_850,In_674,In_622);
and U851 (N_851,In_41,In_42);
or U852 (N_852,In_488,In_196);
nor U853 (N_853,In_626,In_585);
nand U854 (N_854,In_338,In_689);
nand U855 (N_855,In_618,In_356);
nor U856 (N_856,In_54,In_49);
and U857 (N_857,In_303,In_575);
nand U858 (N_858,In_504,In_689);
or U859 (N_859,In_140,In_190);
and U860 (N_860,In_409,In_675);
nand U861 (N_861,In_313,In_661);
nand U862 (N_862,In_575,In_374);
and U863 (N_863,In_191,In_80);
or U864 (N_864,In_679,In_734);
nand U865 (N_865,In_614,In_658);
nor U866 (N_866,In_206,In_418);
nand U867 (N_867,In_49,In_27);
xor U868 (N_868,In_588,In_108);
and U869 (N_869,In_700,In_394);
nand U870 (N_870,In_174,In_527);
nand U871 (N_871,In_396,In_266);
nand U872 (N_872,In_434,In_331);
or U873 (N_873,In_131,In_91);
or U874 (N_874,In_331,In_581);
nor U875 (N_875,In_630,In_420);
and U876 (N_876,In_506,In_655);
or U877 (N_877,In_271,In_190);
nor U878 (N_878,In_281,In_112);
nand U879 (N_879,In_237,In_158);
nand U880 (N_880,In_577,In_479);
nand U881 (N_881,In_334,In_465);
nor U882 (N_882,In_320,In_249);
nand U883 (N_883,In_225,In_140);
and U884 (N_884,In_74,In_220);
or U885 (N_885,In_590,In_617);
or U886 (N_886,In_608,In_23);
nor U887 (N_887,In_209,In_288);
and U888 (N_888,In_268,In_482);
or U889 (N_889,In_341,In_177);
nand U890 (N_890,In_156,In_298);
and U891 (N_891,In_720,In_505);
or U892 (N_892,In_207,In_731);
or U893 (N_893,In_267,In_712);
or U894 (N_894,In_71,In_186);
nor U895 (N_895,In_648,In_163);
or U896 (N_896,In_431,In_662);
nand U897 (N_897,In_313,In_1);
nor U898 (N_898,In_12,In_455);
and U899 (N_899,In_440,In_535);
nor U900 (N_900,In_111,In_276);
or U901 (N_901,In_99,In_583);
or U902 (N_902,In_489,In_82);
nand U903 (N_903,In_119,In_456);
nand U904 (N_904,In_501,In_697);
nand U905 (N_905,In_157,In_40);
nor U906 (N_906,In_600,In_298);
nand U907 (N_907,In_338,In_575);
and U908 (N_908,In_108,In_225);
nand U909 (N_909,In_202,In_596);
nor U910 (N_910,In_688,In_449);
and U911 (N_911,In_257,In_269);
nor U912 (N_912,In_730,In_557);
nor U913 (N_913,In_388,In_653);
or U914 (N_914,In_436,In_255);
or U915 (N_915,In_464,In_459);
nand U916 (N_916,In_353,In_742);
or U917 (N_917,In_73,In_153);
nor U918 (N_918,In_37,In_681);
and U919 (N_919,In_323,In_63);
and U920 (N_920,In_211,In_153);
nand U921 (N_921,In_649,In_684);
and U922 (N_922,In_218,In_257);
or U923 (N_923,In_226,In_185);
or U924 (N_924,In_446,In_197);
nand U925 (N_925,In_366,In_715);
nor U926 (N_926,In_372,In_354);
or U927 (N_927,In_396,In_683);
and U928 (N_928,In_211,In_186);
nand U929 (N_929,In_647,In_369);
nor U930 (N_930,In_343,In_661);
nand U931 (N_931,In_94,In_740);
nor U932 (N_932,In_471,In_346);
or U933 (N_933,In_70,In_698);
and U934 (N_934,In_650,In_656);
or U935 (N_935,In_1,In_44);
nor U936 (N_936,In_256,In_378);
xor U937 (N_937,In_595,In_424);
xor U938 (N_938,In_93,In_526);
and U939 (N_939,In_25,In_54);
or U940 (N_940,In_623,In_462);
nor U941 (N_941,In_338,In_676);
or U942 (N_942,In_654,In_659);
and U943 (N_943,In_641,In_576);
nand U944 (N_944,In_16,In_303);
nand U945 (N_945,In_439,In_393);
nand U946 (N_946,In_92,In_36);
nand U947 (N_947,In_471,In_281);
nor U948 (N_948,In_272,In_236);
or U949 (N_949,In_110,In_325);
nor U950 (N_950,In_427,In_167);
or U951 (N_951,In_477,In_589);
nor U952 (N_952,In_587,In_385);
or U953 (N_953,In_515,In_436);
and U954 (N_954,In_392,In_266);
nand U955 (N_955,In_619,In_262);
nor U956 (N_956,In_316,In_135);
nand U957 (N_957,In_356,In_122);
nor U958 (N_958,In_578,In_236);
nor U959 (N_959,In_548,In_608);
or U960 (N_960,In_531,In_104);
and U961 (N_961,In_729,In_639);
nor U962 (N_962,In_381,In_372);
nor U963 (N_963,In_153,In_181);
or U964 (N_964,In_157,In_531);
nand U965 (N_965,In_263,In_290);
and U966 (N_966,In_748,In_733);
nor U967 (N_967,In_700,In_149);
or U968 (N_968,In_581,In_265);
or U969 (N_969,In_82,In_376);
nand U970 (N_970,In_147,In_667);
or U971 (N_971,In_599,In_239);
nor U972 (N_972,In_638,In_136);
nand U973 (N_973,In_86,In_230);
nor U974 (N_974,In_691,In_575);
nand U975 (N_975,In_509,In_663);
or U976 (N_976,In_26,In_666);
or U977 (N_977,In_316,In_69);
nor U978 (N_978,In_147,In_390);
or U979 (N_979,In_283,In_537);
nor U980 (N_980,In_526,In_276);
or U981 (N_981,In_377,In_609);
or U982 (N_982,In_198,In_313);
nand U983 (N_983,In_668,In_577);
nor U984 (N_984,In_173,In_558);
or U985 (N_985,In_320,In_317);
or U986 (N_986,In_508,In_695);
and U987 (N_987,In_611,In_154);
and U988 (N_988,In_450,In_67);
or U989 (N_989,In_124,In_276);
and U990 (N_990,In_223,In_306);
or U991 (N_991,In_642,In_353);
nor U992 (N_992,In_739,In_434);
nand U993 (N_993,In_350,In_466);
and U994 (N_994,In_442,In_650);
nor U995 (N_995,In_40,In_73);
and U996 (N_996,In_523,In_727);
nor U997 (N_997,In_325,In_252);
or U998 (N_998,In_229,In_331);
nand U999 (N_999,In_89,In_446);
or U1000 (N_1000,N_379,N_589);
and U1001 (N_1001,N_359,N_302);
nand U1002 (N_1002,N_852,N_684);
or U1003 (N_1003,N_101,N_474);
nand U1004 (N_1004,N_710,N_886);
or U1005 (N_1005,N_885,N_707);
nor U1006 (N_1006,N_268,N_425);
nand U1007 (N_1007,N_234,N_844);
and U1008 (N_1008,N_447,N_14);
nor U1009 (N_1009,N_526,N_549);
and U1010 (N_1010,N_221,N_520);
nor U1011 (N_1011,N_409,N_832);
nor U1012 (N_1012,N_255,N_453);
and U1013 (N_1013,N_470,N_790);
nor U1014 (N_1014,N_561,N_626);
or U1015 (N_1015,N_439,N_793);
nand U1016 (N_1016,N_963,N_328);
and U1017 (N_1017,N_401,N_207);
or U1018 (N_1018,N_388,N_93);
nor U1019 (N_1019,N_87,N_729);
or U1020 (N_1020,N_116,N_45);
nand U1021 (N_1021,N_427,N_484);
nor U1022 (N_1022,N_785,N_650);
nand U1023 (N_1023,N_727,N_947);
and U1024 (N_1024,N_381,N_259);
or U1025 (N_1025,N_17,N_52);
and U1026 (N_1026,N_975,N_62);
and U1027 (N_1027,N_716,N_12);
nand U1028 (N_1028,N_536,N_332);
nor U1029 (N_1029,N_461,N_382);
or U1030 (N_1030,N_989,N_666);
nand U1031 (N_1031,N_696,N_336);
and U1032 (N_1032,N_361,N_638);
and U1033 (N_1033,N_321,N_516);
and U1034 (N_1034,N_225,N_751);
nand U1035 (N_1035,N_866,N_556);
nor U1036 (N_1036,N_421,N_30);
nand U1037 (N_1037,N_352,N_827);
nor U1038 (N_1038,N_106,N_835);
nor U1039 (N_1039,N_393,N_412);
nand U1040 (N_1040,N_506,N_616);
nand U1041 (N_1041,N_326,N_528);
nor U1042 (N_1042,N_812,N_871);
and U1043 (N_1043,N_56,N_998);
nand U1044 (N_1044,N_182,N_749);
nor U1045 (N_1045,N_910,N_685);
xnor U1046 (N_1046,N_933,N_77);
nor U1047 (N_1047,N_23,N_983);
nand U1048 (N_1048,N_800,N_246);
nand U1049 (N_1049,N_94,N_612);
nor U1050 (N_1050,N_637,N_568);
and U1051 (N_1051,N_538,N_132);
or U1052 (N_1052,N_976,N_671);
and U1053 (N_1053,N_378,N_633);
nor U1054 (N_1054,N_203,N_406);
nor U1055 (N_1055,N_599,N_490);
nand U1056 (N_1056,N_54,N_266);
nand U1057 (N_1057,N_262,N_86);
nand U1058 (N_1058,N_149,N_475);
and U1059 (N_1059,N_172,N_651);
and U1060 (N_1060,N_597,N_419);
or U1061 (N_1061,N_28,N_402);
nand U1062 (N_1062,N_801,N_937);
nor U1063 (N_1063,N_631,N_31);
nand U1064 (N_1064,N_254,N_394);
nand U1065 (N_1065,N_621,N_480);
nor U1066 (N_1066,N_542,N_60);
or U1067 (N_1067,N_263,N_219);
or U1068 (N_1068,N_691,N_605);
or U1069 (N_1069,N_237,N_3);
nor U1070 (N_1070,N_601,N_936);
nand U1071 (N_1071,N_628,N_166);
nor U1072 (N_1072,N_236,N_297);
nand U1073 (N_1073,N_810,N_532);
or U1074 (N_1074,N_25,N_856);
nand U1075 (N_1075,N_945,N_814);
xor U1076 (N_1076,N_743,N_33);
or U1077 (N_1077,N_99,N_986);
nand U1078 (N_1078,N_985,N_949);
xor U1079 (N_1079,N_652,N_501);
or U1080 (N_1080,N_428,N_803);
or U1081 (N_1081,N_569,N_586);
or U1082 (N_1082,N_741,N_134);
or U1083 (N_1083,N_774,N_72);
xor U1084 (N_1084,N_643,N_126);
nor U1085 (N_1085,N_698,N_279);
xor U1086 (N_1086,N_967,N_261);
nor U1087 (N_1087,N_251,N_113);
nor U1088 (N_1088,N_360,N_574);
nor U1089 (N_1089,N_169,N_160);
nand U1090 (N_1090,N_725,N_471);
or U1091 (N_1091,N_662,N_981);
nor U1092 (N_1092,N_747,N_179);
nor U1093 (N_1093,N_213,N_68);
and U1094 (N_1094,N_485,N_746);
or U1095 (N_1095,N_449,N_327);
and U1096 (N_1096,N_63,N_809);
or U1097 (N_1097,N_728,N_611);
or U1098 (N_1098,N_176,N_206);
and U1099 (N_1099,N_397,N_457);
nand U1100 (N_1100,N_629,N_431);
nor U1101 (N_1101,N_383,N_996);
nand U1102 (N_1102,N_994,N_585);
nor U1103 (N_1103,N_833,N_226);
nand U1104 (N_1104,N_385,N_539);
nor U1105 (N_1105,N_953,N_318);
and U1106 (N_1106,N_465,N_733);
and U1107 (N_1107,N_788,N_119);
xor U1108 (N_1108,N_120,N_962);
nor U1109 (N_1109,N_831,N_80);
and U1110 (N_1110,N_548,N_567);
and U1111 (N_1111,N_175,N_735);
nand U1112 (N_1112,N_534,N_613);
nand U1113 (N_1113,N_342,N_928);
nor U1114 (N_1114,N_39,N_181);
or U1115 (N_1115,N_913,N_271);
and U1116 (N_1116,N_712,N_952);
and U1117 (N_1117,N_584,N_906);
or U1118 (N_1118,N_9,N_35);
and U1119 (N_1119,N_111,N_514);
and U1120 (N_1120,N_604,N_647);
and U1121 (N_1121,N_300,N_414);
nand U1122 (N_1122,N_600,N_103);
nor U1123 (N_1123,N_137,N_369);
xnor U1124 (N_1124,N_267,N_156);
and U1125 (N_1125,N_893,N_990);
nor U1126 (N_1126,N_993,N_592);
xor U1127 (N_1127,N_890,N_42);
or U1128 (N_1128,N_367,N_349);
or U1129 (N_1129,N_552,N_508);
and U1130 (N_1130,N_139,N_523);
xor U1131 (N_1131,N_750,N_531);
xnor U1132 (N_1132,N_96,N_673);
nand U1133 (N_1133,N_109,N_620);
xnor U1134 (N_1134,N_242,N_277);
nor U1135 (N_1135,N_956,N_432);
nand U1136 (N_1136,N_21,N_55);
nor U1137 (N_1137,N_791,N_298);
and U1138 (N_1138,N_766,N_338);
or U1139 (N_1139,N_129,N_737);
and U1140 (N_1140,N_69,N_853);
and U1141 (N_1141,N_191,N_104);
nor U1142 (N_1142,N_16,N_407);
nor U1143 (N_1143,N_672,N_732);
nand U1144 (N_1144,N_877,N_609);
nor U1145 (N_1145,N_171,N_183);
or U1146 (N_1146,N_982,N_164);
or U1147 (N_1147,N_205,N_595);
and U1148 (N_1148,N_596,N_83);
and U1149 (N_1149,N_836,N_905);
and U1150 (N_1150,N_173,N_920);
nand U1151 (N_1151,N_224,N_822);
nand U1152 (N_1152,N_829,N_7);
and U1153 (N_1153,N_430,N_49);
or U1154 (N_1154,N_257,N_1);
nand U1155 (N_1155,N_415,N_416);
or U1156 (N_1156,N_358,N_854);
nor U1157 (N_1157,N_697,N_617);
or U1158 (N_1158,N_591,N_838);
or U1159 (N_1159,N_452,N_376);
and U1160 (N_1160,N_346,N_524);
nor U1161 (N_1161,N_888,N_840);
nor U1162 (N_1162,N_107,N_942);
and U1163 (N_1163,N_680,N_67);
nor U1164 (N_1164,N_272,N_722);
xor U1165 (N_1165,N_797,N_497);
nand U1166 (N_1166,N_5,N_876);
nand U1167 (N_1167,N_201,N_50);
nand U1168 (N_1168,N_934,N_783);
nand U1169 (N_1169,N_250,N_24);
or U1170 (N_1170,N_65,N_899);
nor U1171 (N_1171,N_75,N_105);
nor U1172 (N_1172,N_765,N_153);
or U1173 (N_1173,N_71,N_159);
or U1174 (N_1174,N_841,N_287);
nor U1175 (N_1175,N_868,N_274);
or U1176 (N_1176,N_6,N_456);
or U1177 (N_1177,N_941,N_217);
or U1178 (N_1178,N_755,N_721);
nand U1179 (N_1179,N_329,N_355);
or U1180 (N_1180,N_79,N_794);
nand U1181 (N_1181,N_420,N_608);
nor U1182 (N_1182,N_187,N_694);
nor U1183 (N_1183,N_734,N_450);
or U1184 (N_1184,N_486,N_921);
xor U1185 (N_1185,N_463,N_593);
and U1186 (N_1186,N_97,N_563);
or U1187 (N_1187,N_404,N_752);
xnor U1188 (N_1188,N_730,N_701);
or U1189 (N_1189,N_276,N_639);
nand U1190 (N_1190,N_214,N_818);
nand U1191 (N_1191,N_331,N_657);
and U1192 (N_1192,N_310,N_339);
or U1193 (N_1193,N_770,N_896);
or U1194 (N_1194,N_908,N_659);
and U1195 (N_1195,N_987,N_317);
or U1196 (N_1196,N_163,N_925);
nand U1197 (N_1197,N_140,N_984);
or U1198 (N_1198,N_964,N_566);
or U1199 (N_1199,N_411,N_708);
or U1200 (N_1200,N_195,N_862);
nand U1201 (N_1201,N_780,N_229);
nand U1202 (N_1202,N_714,N_564);
and U1203 (N_1203,N_726,N_133);
and U1204 (N_1204,N_804,N_819);
or U1205 (N_1205,N_807,N_477);
nor U1206 (N_1206,N_142,N_131);
or U1207 (N_1207,N_627,N_748);
nand U1208 (N_1208,N_951,N_285);
or U1209 (N_1209,N_437,N_648);
and U1210 (N_1210,N_162,N_618);
nor U1211 (N_1211,N_158,N_110);
nand U1212 (N_1212,N_578,N_700);
nor U1213 (N_1213,N_861,N_966);
nor U1214 (N_1214,N_972,N_959);
and U1215 (N_1215,N_577,N_570);
nand U1216 (N_1216,N_434,N_192);
nand U1217 (N_1217,N_399,N_66);
nand U1218 (N_1218,N_209,N_417);
nor U1219 (N_1219,N_881,N_114);
nand U1220 (N_1220,N_51,N_47);
nor U1221 (N_1221,N_322,N_573);
and U1222 (N_1222,N_311,N_223);
nand U1223 (N_1223,N_375,N_978);
or U1224 (N_1224,N_273,N_924);
nor U1225 (N_1225,N_773,N_34);
or U1226 (N_1226,N_681,N_828);
or U1227 (N_1227,N_436,N_806);
and U1228 (N_1228,N_923,N_0);
and U1229 (N_1229,N_674,N_527);
nor U1230 (N_1230,N_560,N_736);
nand U1231 (N_1231,N_454,N_602);
or U1232 (N_1232,N_761,N_281);
and U1233 (N_1233,N_979,N_851);
or U1234 (N_1234,N_521,N_845);
and U1235 (N_1235,N_22,N_745);
nor U1236 (N_1236,N_805,N_943);
or U1237 (N_1237,N_699,N_997);
and U1238 (N_1238,N_940,N_446);
nand U1239 (N_1239,N_880,N_948);
nor U1240 (N_1240,N_911,N_505);
nand U1241 (N_1241,N_709,N_320);
nor U1242 (N_1242,N_233,N_717);
nand U1243 (N_1243,N_879,N_429);
or U1244 (N_1244,N_922,N_194);
nor U1245 (N_1245,N_445,N_912);
nor U1246 (N_1246,N_384,N_558);
nor U1247 (N_1247,N_715,N_782);
or U1248 (N_1248,N_144,N_847);
or U1249 (N_1249,N_571,N_572);
and U1250 (N_1250,N_410,N_798);
and U1251 (N_1251,N_4,N_61);
or U1252 (N_1252,N_646,N_330);
nand U1253 (N_1253,N_395,N_290);
xnor U1254 (N_1254,N_193,N_84);
or U1255 (N_1255,N_253,N_889);
or U1256 (N_1256,N_15,N_227);
or U1257 (N_1257,N_530,N_664);
and U1258 (N_1258,N_869,N_232);
xor U1259 (N_1259,N_291,N_704);
and U1260 (N_1260,N_817,N_796);
nand U1261 (N_1261,N_895,N_240);
nand U1262 (N_1262,N_100,N_799);
or U1263 (N_1263,N_825,N_325);
nor U1264 (N_1264,N_580,N_513);
and U1265 (N_1265,N_692,N_878);
nor U1266 (N_1266,N_370,N_282);
and U1267 (N_1267,N_316,N_754);
nand U1268 (N_1268,N_517,N_81);
xnor U1269 (N_1269,N_509,N_151);
and U1270 (N_1270,N_992,N_772);
and U1271 (N_1271,N_269,N_781);
nor U1272 (N_1272,N_478,N_843);
and U1273 (N_1273,N_495,N_642);
or U1274 (N_1274,N_91,N_37);
xor U1275 (N_1275,N_625,N_653);
nand U1276 (N_1276,N_396,N_256);
and U1277 (N_1277,N_260,N_245);
xor U1278 (N_1278,N_135,N_705);
nand U1279 (N_1279,N_897,N_408);
and U1280 (N_1280,N_703,N_645);
and U1281 (N_1281,N_422,N_813);
nand U1282 (N_1282,N_622,N_220);
nor U1283 (N_1283,N_903,N_289);
nor U1284 (N_1284,N_826,N_916);
or U1285 (N_1285,N_343,N_278);
or U1286 (N_1286,N_353,N_669);
or U1287 (N_1287,N_230,N_152);
nor U1288 (N_1288,N_44,N_711);
and U1289 (N_1289,N_479,N_795);
nand U1290 (N_1290,N_632,N_540);
and U1291 (N_1291,N_875,N_340);
nor U1292 (N_1292,N_503,N_767);
or U1293 (N_1293,N_939,N_636);
and U1294 (N_1294,N_496,N_459);
nand U1295 (N_1295,N_786,N_180);
nor U1296 (N_1296,N_720,N_130);
nor U1297 (N_1297,N_27,N_18);
nand U1298 (N_1298,N_491,N_76);
or U1299 (N_1299,N_961,N_759);
or U1300 (N_1300,N_46,N_892);
or U1301 (N_1301,N_545,N_398);
nor U1302 (N_1302,N_29,N_579);
and U1303 (N_1303,N_228,N_502);
nand U1304 (N_1304,N_466,N_583);
nor U1305 (N_1305,N_954,N_347);
or U1306 (N_1306,N_124,N_48);
nand U1307 (N_1307,N_188,N_882);
and U1308 (N_1308,N_846,N_839);
and U1309 (N_1309,N_918,N_295);
and U1310 (N_1310,N_121,N_145);
and U1311 (N_1311,N_323,N_265);
and U1312 (N_1312,N_870,N_689);
nor U1313 (N_1313,N_762,N_695);
and U1314 (N_1314,N_365,N_258);
or U1315 (N_1315,N_619,N_679);
or U1316 (N_1316,N_199,N_678);
nand U1317 (N_1317,N_90,N_498);
or U1318 (N_1318,N_630,N_624);
and U1319 (N_1319,N_958,N_309);
nor U1320 (N_1320,N_644,N_901);
xor U1321 (N_1321,N_235,N_904);
or U1322 (N_1322,N_334,N_150);
and U1323 (N_1323,N_462,N_357);
or U1324 (N_1324,N_955,N_489);
or U1325 (N_1325,N_581,N_122);
nand U1326 (N_1326,N_872,N_125);
nor U1327 (N_1327,N_19,N_594);
or U1328 (N_1328,N_894,N_143);
and U1329 (N_1329,N_675,N_59);
nand U1330 (N_1330,N_864,N_283);
and U1331 (N_1331,N_543,N_373);
or U1332 (N_1332,N_834,N_248);
and U1333 (N_1333,N_756,N_64);
and U1334 (N_1334,N_706,N_165);
and U1335 (N_1335,N_582,N_946);
nor U1336 (N_1336,N_89,N_190);
nor U1337 (N_1337,N_649,N_372);
or U1338 (N_1338,N_968,N_341);
nand U1339 (N_1339,N_102,N_557);
nor U1340 (N_1340,N_73,N_351);
or U1341 (N_1341,N_211,N_304);
nand U1342 (N_1342,N_930,N_515);
and U1343 (N_1343,N_155,N_239);
nand U1344 (N_1344,N_999,N_512);
nand U1345 (N_1345,N_400,N_88);
or U1346 (N_1346,N_682,N_189);
and U1347 (N_1347,N_403,N_518);
nand U1348 (N_1348,N_319,N_969);
nor U1349 (N_1349,N_314,N_487);
and U1350 (N_1350,N_640,N_816);
nand U1351 (N_1351,N_529,N_157);
or U1352 (N_1352,N_500,N_202);
and U1353 (N_1353,N_335,N_931);
nor U1354 (N_1354,N_354,N_123);
nor U1355 (N_1355,N_757,N_740);
or U1356 (N_1356,N_820,N_483);
nand U1357 (N_1357,N_656,N_212);
nand U1358 (N_1358,N_658,N_927);
nor U1359 (N_1359,N_654,N_635);
nor U1360 (N_1360,N_10,N_92);
nor U1361 (N_1361,N_348,N_198);
and U1362 (N_1362,N_857,N_53);
or U1363 (N_1363,N_458,N_288);
and U1364 (N_1364,N_390,N_296);
or U1365 (N_1365,N_824,N_555);
nor U1366 (N_1366,N_424,N_389);
nand U1367 (N_1367,N_222,N_115);
and U1368 (N_1368,N_914,N_719);
nand U1369 (N_1369,N_301,N_686);
and U1370 (N_1370,N_185,N_441);
and U1371 (N_1371,N_270,N_960);
and U1372 (N_1372,N_128,N_623);
or U1373 (N_1373,N_210,N_11);
nor U1374 (N_1374,N_57,N_590);
nor U1375 (N_1375,N_683,N_467);
and U1376 (N_1376,N_468,N_688);
and U1377 (N_1377,N_935,N_108);
and U1378 (N_1378,N_855,N_482);
nand U1379 (N_1379,N_74,N_333);
nand U1380 (N_1380,N_693,N_26);
nor U1381 (N_1381,N_136,N_723);
and U1382 (N_1382,N_641,N_286);
and U1383 (N_1383,N_473,N_208);
nand U1384 (N_1384,N_293,N_363);
nor U1385 (N_1385,N_535,N_161);
nor U1386 (N_1386,N_859,N_95);
nand U1387 (N_1387,N_537,N_82);
nand U1388 (N_1388,N_196,N_768);
nand U1389 (N_1389,N_760,N_830);
nor U1390 (N_1390,N_547,N_443);
nor U1391 (N_1391,N_455,N_98);
nor U1392 (N_1392,N_525,N_469);
or U1393 (N_1393,N_867,N_763);
and U1394 (N_1394,N_977,N_551);
or U1395 (N_1395,N_660,N_738);
nor U1396 (N_1396,N_544,N_744);
and U1397 (N_1397,N_823,N_676);
nand U1398 (N_1398,N_554,N_607);
nor U1399 (N_1399,N_511,N_174);
or U1400 (N_1400,N_494,N_808);
and U1401 (N_1401,N_661,N_344);
nand U1402 (N_1402,N_464,N_368);
nor U1403 (N_1403,N_907,N_350);
or U1404 (N_1404,N_873,N_909);
and U1405 (N_1405,N_932,N_41);
nor U1406 (N_1406,N_777,N_837);
nor U1407 (N_1407,N_138,N_216);
nor U1408 (N_1408,N_218,N_117);
nor U1409 (N_1409,N_448,N_186);
nor U1410 (N_1410,N_519,N_247);
nor U1411 (N_1411,N_442,N_665);
and U1412 (N_1412,N_776,N_364);
nor U1413 (N_1413,N_944,N_655);
nand U1414 (N_1414,N_610,N_435);
nor U1415 (N_1415,N_178,N_702);
nand U1416 (N_1416,N_371,N_78);
and U1417 (N_1417,N_957,N_20);
nand U1418 (N_1418,N_507,N_147);
and U1419 (N_1419,N_112,N_863);
nand U1420 (N_1420,N_778,N_440);
nor U1421 (N_1421,N_575,N_973);
nand U1422 (N_1422,N_391,N_988);
nor U1423 (N_1423,N_294,N_313);
nor U1424 (N_1424,N_898,N_874);
nor U1425 (N_1425,N_154,N_902);
nand U1426 (N_1426,N_13,N_141);
nor U1427 (N_1427,N_849,N_758);
nor U1428 (N_1428,N_292,N_677);
and U1429 (N_1429,N_127,N_85);
xor U1430 (N_1430,N_433,N_418);
nor U1431 (N_1431,N_244,N_965);
and U1432 (N_1432,N_917,N_426);
nand U1433 (N_1433,N_850,N_284);
and U1434 (N_1434,N_562,N_598);
and U1435 (N_1435,N_356,N_576);
nor U1436 (N_1436,N_553,N_241);
and U1437 (N_1437,N_2,N_634);
and U1438 (N_1438,N_231,N_405);
or U1439 (N_1439,N_811,N_40);
or U1440 (N_1440,N_784,N_883);
or U1441 (N_1441,N_713,N_148);
and U1442 (N_1442,N_614,N_887);
and U1443 (N_1443,N_249,N_374);
nand U1444 (N_1444,N_771,N_451);
nor U1445 (N_1445,N_587,N_603);
or U1446 (N_1446,N_324,N_58);
or U1447 (N_1447,N_168,N_769);
or U1448 (N_1448,N_215,N_858);
nand U1449 (N_1449,N_177,N_315);
nand U1450 (N_1450,N_891,N_306);
and U1451 (N_1451,N_238,N_789);
or U1452 (N_1452,N_667,N_308);
or U1453 (N_1453,N_481,N_444);
and U1454 (N_1454,N_307,N_510);
nand U1455 (N_1455,N_775,N_387);
nand U1456 (N_1456,N_550,N_970);
or U1457 (N_1457,N_337,N_146);
nand U1458 (N_1458,N_522,N_32);
nor U1459 (N_1459,N_460,N_541);
and U1460 (N_1460,N_848,N_303);
nor U1461 (N_1461,N_36,N_559);
and U1462 (N_1462,N_974,N_615);
xnor U1463 (N_1463,N_919,N_724);
nand U1464 (N_1464,N_70,N_565);
nor U1465 (N_1465,N_299,N_687);
or U1466 (N_1466,N_312,N_377);
nor U1467 (N_1467,N_742,N_546);
and U1468 (N_1468,N_438,N_670);
nand U1469 (N_1469,N_792,N_476);
or U1470 (N_1470,N_8,N_950);
nor U1471 (N_1471,N_764,N_197);
and U1472 (N_1472,N_860,N_413);
and U1473 (N_1473,N_588,N_366);
and U1474 (N_1474,N_787,N_252);
nand U1475 (N_1475,N_668,N_929);
nor U1476 (N_1476,N_533,N_184);
and U1477 (N_1477,N_170,N_802);
and U1478 (N_1478,N_991,N_492);
nor U1479 (N_1479,N_884,N_362);
nor U1480 (N_1480,N_243,N_690);
or U1481 (N_1481,N_493,N_423);
nand U1482 (N_1482,N_204,N_43);
nor U1483 (N_1483,N_663,N_718);
and U1484 (N_1484,N_200,N_815);
nand U1485 (N_1485,N_779,N_865);
and U1486 (N_1486,N_305,N_995);
nand U1487 (N_1487,N_275,N_938);
or U1488 (N_1488,N_900,N_926);
and U1489 (N_1489,N_345,N_264);
and U1490 (N_1490,N_38,N_118);
and U1491 (N_1491,N_280,N_606);
nor U1492 (N_1492,N_753,N_392);
nor U1493 (N_1493,N_915,N_971);
nand U1494 (N_1494,N_821,N_386);
or U1495 (N_1495,N_499,N_504);
and U1496 (N_1496,N_488,N_980);
nor U1497 (N_1497,N_380,N_167);
or U1498 (N_1498,N_739,N_472);
xor U1499 (N_1499,N_842,N_731);
nor U1500 (N_1500,N_14,N_811);
or U1501 (N_1501,N_937,N_251);
nor U1502 (N_1502,N_588,N_979);
nand U1503 (N_1503,N_773,N_644);
and U1504 (N_1504,N_58,N_159);
nand U1505 (N_1505,N_306,N_210);
nor U1506 (N_1506,N_467,N_196);
or U1507 (N_1507,N_171,N_128);
nand U1508 (N_1508,N_195,N_684);
or U1509 (N_1509,N_569,N_918);
and U1510 (N_1510,N_468,N_893);
and U1511 (N_1511,N_231,N_714);
nor U1512 (N_1512,N_611,N_13);
nand U1513 (N_1513,N_770,N_421);
or U1514 (N_1514,N_485,N_297);
nor U1515 (N_1515,N_46,N_480);
nor U1516 (N_1516,N_287,N_554);
nand U1517 (N_1517,N_672,N_536);
nand U1518 (N_1518,N_972,N_39);
nor U1519 (N_1519,N_751,N_731);
or U1520 (N_1520,N_196,N_901);
or U1521 (N_1521,N_128,N_395);
or U1522 (N_1522,N_389,N_114);
nor U1523 (N_1523,N_845,N_25);
nand U1524 (N_1524,N_174,N_2);
nor U1525 (N_1525,N_324,N_960);
and U1526 (N_1526,N_560,N_159);
and U1527 (N_1527,N_882,N_533);
nor U1528 (N_1528,N_533,N_942);
nand U1529 (N_1529,N_18,N_788);
xnor U1530 (N_1530,N_64,N_44);
nor U1531 (N_1531,N_802,N_230);
nor U1532 (N_1532,N_28,N_189);
nor U1533 (N_1533,N_923,N_640);
and U1534 (N_1534,N_328,N_85);
nand U1535 (N_1535,N_594,N_235);
and U1536 (N_1536,N_598,N_634);
or U1537 (N_1537,N_866,N_535);
nand U1538 (N_1538,N_776,N_891);
nand U1539 (N_1539,N_543,N_488);
and U1540 (N_1540,N_413,N_568);
or U1541 (N_1541,N_905,N_276);
nand U1542 (N_1542,N_976,N_94);
and U1543 (N_1543,N_150,N_482);
and U1544 (N_1544,N_964,N_176);
or U1545 (N_1545,N_302,N_64);
or U1546 (N_1546,N_2,N_146);
nand U1547 (N_1547,N_579,N_380);
nor U1548 (N_1548,N_794,N_143);
or U1549 (N_1549,N_666,N_947);
nand U1550 (N_1550,N_958,N_915);
or U1551 (N_1551,N_661,N_616);
nand U1552 (N_1552,N_897,N_220);
and U1553 (N_1553,N_423,N_487);
nor U1554 (N_1554,N_239,N_456);
nand U1555 (N_1555,N_410,N_308);
or U1556 (N_1556,N_85,N_989);
nand U1557 (N_1557,N_124,N_712);
nor U1558 (N_1558,N_88,N_117);
and U1559 (N_1559,N_987,N_984);
nor U1560 (N_1560,N_258,N_394);
or U1561 (N_1561,N_706,N_671);
nand U1562 (N_1562,N_742,N_485);
nand U1563 (N_1563,N_320,N_928);
nor U1564 (N_1564,N_267,N_528);
nand U1565 (N_1565,N_841,N_374);
or U1566 (N_1566,N_62,N_102);
and U1567 (N_1567,N_285,N_799);
or U1568 (N_1568,N_617,N_441);
or U1569 (N_1569,N_942,N_718);
nand U1570 (N_1570,N_71,N_421);
nor U1571 (N_1571,N_858,N_880);
and U1572 (N_1572,N_898,N_942);
nor U1573 (N_1573,N_61,N_905);
and U1574 (N_1574,N_490,N_332);
nor U1575 (N_1575,N_508,N_911);
nor U1576 (N_1576,N_998,N_446);
nor U1577 (N_1577,N_429,N_0);
and U1578 (N_1578,N_337,N_888);
nor U1579 (N_1579,N_762,N_972);
nand U1580 (N_1580,N_47,N_127);
or U1581 (N_1581,N_805,N_799);
nand U1582 (N_1582,N_417,N_600);
nor U1583 (N_1583,N_463,N_468);
nor U1584 (N_1584,N_19,N_426);
nand U1585 (N_1585,N_36,N_116);
or U1586 (N_1586,N_879,N_778);
or U1587 (N_1587,N_459,N_973);
nand U1588 (N_1588,N_805,N_474);
nor U1589 (N_1589,N_344,N_249);
nand U1590 (N_1590,N_963,N_493);
or U1591 (N_1591,N_711,N_81);
or U1592 (N_1592,N_623,N_56);
nand U1593 (N_1593,N_280,N_830);
nand U1594 (N_1594,N_332,N_619);
nand U1595 (N_1595,N_257,N_963);
nor U1596 (N_1596,N_998,N_292);
nand U1597 (N_1597,N_515,N_243);
or U1598 (N_1598,N_766,N_904);
and U1599 (N_1599,N_587,N_100);
nand U1600 (N_1600,N_794,N_579);
and U1601 (N_1601,N_979,N_92);
nor U1602 (N_1602,N_733,N_628);
nor U1603 (N_1603,N_68,N_648);
nand U1604 (N_1604,N_227,N_683);
xnor U1605 (N_1605,N_4,N_975);
nor U1606 (N_1606,N_231,N_461);
nand U1607 (N_1607,N_263,N_458);
nand U1608 (N_1608,N_747,N_372);
or U1609 (N_1609,N_346,N_377);
nor U1610 (N_1610,N_734,N_14);
and U1611 (N_1611,N_950,N_821);
nand U1612 (N_1612,N_114,N_166);
nand U1613 (N_1613,N_666,N_693);
nor U1614 (N_1614,N_504,N_967);
or U1615 (N_1615,N_154,N_641);
nand U1616 (N_1616,N_815,N_691);
nand U1617 (N_1617,N_858,N_66);
nand U1618 (N_1618,N_917,N_14);
and U1619 (N_1619,N_718,N_78);
nor U1620 (N_1620,N_637,N_16);
or U1621 (N_1621,N_843,N_789);
xor U1622 (N_1622,N_393,N_158);
and U1623 (N_1623,N_883,N_424);
or U1624 (N_1624,N_506,N_83);
nand U1625 (N_1625,N_136,N_363);
or U1626 (N_1626,N_514,N_81);
and U1627 (N_1627,N_452,N_601);
and U1628 (N_1628,N_93,N_244);
nor U1629 (N_1629,N_698,N_889);
nand U1630 (N_1630,N_604,N_876);
nor U1631 (N_1631,N_972,N_686);
and U1632 (N_1632,N_117,N_968);
or U1633 (N_1633,N_481,N_639);
or U1634 (N_1634,N_495,N_266);
nand U1635 (N_1635,N_619,N_73);
nor U1636 (N_1636,N_386,N_845);
nor U1637 (N_1637,N_777,N_761);
or U1638 (N_1638,N_123,N_22);
or U1639 (N_1639,N_572,N_11);
and U1640 (N_1640,N_408,N_647);
or U1641 (N_1641,N_285,N_723);
or U1642 (N_1642,N_139,N_792);
nand U1643 (N_1643,N_733,N_111);
and U1644 (N_1644,N_737,N_461);
or U1645 (N_1645,N_514,N_17);
nor U1646 (N_1646,N_225,N_839);
nor U1647 (N_1647,N_688,N_959);
nor U1648 (N_1648,N_951,N_524);
nor U1649 (N_1649,N_994,N_19);
or U1650 (N_1650,N_593,N_263);
and U1651 (N_1651,N_252,N_638);
xor U1652 (N_1652,N_461,N_61);
nand U1653 (N_1653,N_840,N_368);
nand U1654 (N_1654,N_886,N_307);
and U1655 (N_1655,N_799,N_847);
nor U1656 (N_1656,N_905,N_505);
and U1657 (N_1657,N_830,N_865);
nand U1658 (N_1658,N_109,N_992);
nor U1659 (N_1659,N_553,N_7);
nor U1660 (N_1660,N_434,N_814);
nor U1661 (N_1661,N_20,N_83);
nor U1662 (N_1662,N_180,N_212);
and U1663 (N_1663,N_593,N_615);
and U1664 (N_1664,N_697,N_544);
nand U1665 (N_1665,N_355,N_558);
nor U1666 (N_1666,N_634,N_474);
nand U1667 (N_1667,N_492,N_613);
or U1668 (N_1668,N_400,N_82);
nor U1669 (N_1669,N_419,N_128);
or U1670 (N_1670,N_927,N_702);
nand U1671 (N_1671,N_634,N_165);
or U1672 (N_1672,N_668,N_310);
nand U1673 (N_1673,N_566,N_66);
nor U1674 (N_1674,N_4,N_31);
nand U1675 (N_1675,N_235,N_668);
or U1676 (N_1676,N_105,N_186);
nor U1677 (N_1677,N_141,N_237);
xor U1678 (N_1678,N_375,N_946);
and U1679 (N_1679,N_441,N_401);
or U1680 (N_1680,N_522,N_624);
nand U1681 (N_1681,N_727,N_870);
nand U1682 (N_1682,N_67,N_485);
and U1683 (N_1683,N_771,N_186);
nand U1684 (N_1684,N_604,N_846);
nand U1685 (N_1685,N_732,N_848);
and U1686 (N_1686,N_390,N_356);
or U1687 (N_1687,N_912,N_3);
or U1688 (N_1688,N_777,N_600);
and U1689 (N_1689,N_139,N_481);
nand U1690 (N_1690,N_216,N_412);
and U1691 (N_1691,N_620,N_782);
and U1692 (N_1692,N_509,N_139);
and U1693 (N_1693,N_898,N_621);
and U1694 (N_1694,N_601,N_853);
nand U1695 (N_1695,N_452,N_704);
nor U1696 (N_1696,N_833,N_361);
and U1697 (N_1697,N_956,N_395);
nor U1698 (N_1698,N_644,N_848);
nor U1699 (N_1699,N_201,N_851);
nand U1700 (N_1700,N_455,N_656);
nor U1701 (N_1701,N_279,N_898);
nor U1702 (N_1702,N_353,N_350);
nor U1703 (N_1703,N_740,N_289);
nand U1704 (N_1704,N_457,N_232);
or U1705 (N_1705,N_482,N_674);
xor U1706 (N_1706,N_707,N_751);
or U1707 (N_1707,N_665,N_16);
nand U1708 (N_1708,N_137,N_825);
nor U1709 (N_1709,N_578,N_245);
nor U1710 (N_1710,N_396,N_92);
and U1711 (N_1711,N_996,N_280);
nand U1712 (N_1712,N_597,N_926);
or U1713 (N_1713,N_504,N_760);
and U1714 (N_1714,N_697,N_355);
and U1715 (N_1715,N_330,N_484);
nor U1716 (N_1716,N_952,N_862);
or U1717 (N_1717,N_965,N_633);
nand U1718 (N_1718,N_535,N_547);
or U1719 (N_1719,N_263,N_965);
nor U1720 (N_1720,N_561,N_242);
or U1721 (N_1721,N_306,N_481);
nor U1722 (N_1722,N_67,N_526);
and U1723 (N_1723,N_941,N_127);
and U1724 (N_1724,N_692,N_236);
nand U1725 (N_1725,N_620,N_917);
nor U1726 (N_1726,N_464,N_66);
or U1727 (N_1727,N_458,N_465);
or U1728 (N_1728,N_186,N_8);
or U1729 (N_1729,N_501,N_276);
and U1730 (N_1730,N_58,N_688);
nor U1731 (N_1731,N_824,N_558);
or U1732 (N_1732,N_685,N_543);
nand U1733 (N_1733,N_748,N_907);
or U1734 (N_1734,N_229,N_797);
and U1735 (N_1735,N_210,N_800);
nand U1736 (N_1736,N_107,N_302);
or U1737 (N_1737,N_681,N_383);
nand U1738 (N_1738,N_814,N_666);
nand U1739 (N_1739,N_46,N_441);
nor U1740 (N_1740,N_328,N_357);
or U1741 (N_1741,N_788,N_534);
nand U1742 (N_1742,N_875,N_212);
and U1743 (N_1743,N_76,N_433);
or U1744 (N_1744,N_939,N_662);
nor U1745 (N_1745,N_995,N_525);
and U1746 (N_1746,N_243,N_112);
or U1747 (N_1747,N_60,N_386);
or U1748 (N_1748,N_942,N_565);
nand U1749 (N_1749,N_819,N_60);
or U1750 (N_1750,N_198,N_405);
nand U1751 (N_1751,N_14,N_139);
nand U1752 (N_1752,N_190,N_803);
nand U1753 (N_1753,N_347,N_331);
or U1754 (N_1754,N_545,N_787);
nor U1755 (N_1755,N_462,N_464);
nor U1756 (N_1756,N_233,N_35);
or U1757 (N_1757,N_98,N_240);
and U1758 (N_1758,N_719,N_607);
nand U1759 (N_1759,N_961,N_199);
and U1760 (N_1760,N_351,N_657);
or U1761 (N_1761,N_460,N_21);
nor U1762 (N_1762,N_210,N_733);
nand U1763 (N_1763,N_3,N_772);
and U1764 (N_1764,N_2,N_194);
nand U1765 (N_1765,N_295,N_199);
or U1766 (N_1766,N_803,N_792);
or U1767 (N_1767,N_690,N_900);
or U1768 (N_1768,N_418,N_677);
nor U1769 (N_1769,N_455,N_42);
and U1770 (N_1770,N_238,N_545);
and U1771 (N_1771,N_284,N_531);
nand U1772 (N_1772,N_556,N_364);
nor U1773 (N_1773,N_116,N_224);
and U1774 (N_1774,N_280,N_430);
and U1775 (N_1775,N_389,N_835);
and U1776 (N_1776,N_546,N_319);
nor U1777 (N_1777,N_176,N_927);
or U1778 (N_1778,N_466,N_238);
nand U1779 (N_1779,N_24,N_840);
nand U1780 (N_1780,N_631,N_582);
nor U1781 (N_1781,N_229,N_416);
nor U1782 (N_1782,N_276,N_616);
or U1783 (N_1783,N_429,N_768);
nor U1784 (N_1784,N_97,N_948);
nand U1785 (N_1785,N_356,N_348);
nor U1786 (N_1786,N_655,N_446);
and U1787 (N_1787,N_462,N_124);
or U1788 (N_1788,N_669,N_12);
or U1789 (N_1789,N_348,N_779);
nor U1790 (N_1790,N_154,N_752);
nand U1791 (N_1791,N_982,N_380);
xor U1792 (N_1792,N_270,N_196);
and U1793 (N_1793,N_35,N_623);
nor U1794 (N_1794,N_718,N_386);
nor U1795 (N_1795,N_848,N_603);
or U1796 (N_1796,N_305,N_932);
nand U1797 (N_1797,N_824,N_757);
or U1798 (N_1798,N_351,N_626);
and U1799 (N_1799,N_906,N_615);
nor U1800 (N_1800,N_896,N_721);
nand U1801 (N_1801,N_230,N_917);
nand U1802 (N_1802,N_814,N_205);
nor U1803 (N_1803,N_649,N_854);
nor U1804 (N_1804,N_183,N_502);
and U1805 (N_1805,N_513,N_53);
nand U1806 (N_1806,N_330,N_535);
or U1807 (N_1807,N_31,N_767);
and U1808 (N_1808,N_238,N_509);
or U1809 (N_1809,N_484,N_265);
nand U1810 (N_1810,N_667,N_507);
nor U1811 (N_1811,N_929,N_867);
or U1812 (N_1812,N_280,N_105);
nor U1813 (N_1813,N_456,N_120);
or U1814 (N_1814,N_37,N_320);
nand U1815 (N_1815,N_644,N_898);
or U1816 (N_1816,N_397,N_311);
or U1817 (N_1817,N_508,N_897);
nand U1818 (N_1818,N_497,N_396);
and U1819 (N_1819,N_598,N_180);
nor U1820 (N_1820,N_541,N_54);
nor U1821 (N_1821,N_208,N_173);
nand U1822 (N_1822,N_954,N_901);
and U1823 (N_1823,N_206,N_208);
and U1824 (N_1824,N_802,N_982);
and U1825 (N_1825,N_439,N_953);
nand U1826 (N_1826,N_99,N_123);
and U1827 (N_1827,N_748,N_806);
xnor U1828 (N_1828,N_585,N_0);
xor U1829 (N_1829,N_540,N_69);
or U1830 (N_1830,N_916,N_891);
or U1831 (N_1831,N_82,N_946);
nand U1832 (N_1832,N_619,N_710);
xnor U1833 (N_1833,N_243,N_873);
nand U1834 (N_1834,N_921,N_406);
nand U1835 (N_1835,N_376,N_590);
or U1836 (N_1836,N_84,N_431);
nor U1837 (N_1837,N_82,N_772);
xor U1838 (N_1838,N_688,N_968);
or U1839 (N_1839,N_406,N_344);
nand U1840 (N_1840,N_524,N_382);
or U1841 (N_1841,N_241,N_977);
nor U1842 (N_1842,N_91,N_670);
or U1843 (N_1843,N_116,N_909);
and U1844 (N_1844,N_834,N_877);
nand U1845 (N_1845,N_65,N_272);
or U1846 (N_1846,N_616,N_262);
nor U1847 (N_1847,N_90,N_151);
nand U1848 (N_1848,N_311,N_137);
nand U1849 (N_1849,N_922,N_119);
nand U1850 (N_1850,N_101,N_755);
nand U1851 (N_1851,N_485,N_981);
nand U1852 (N_1852,N_394,N_447);
nand U1853 (N_1853,N_859,N_82);
nand U1854 (N_1854,N_913,N_994);
nand U1855 (N_1855,N_499,N_713);
or U1856 (N_1856,N_525,N_32);
nand U1857 (N_1857,N_145,N_771);
nand U1858 (N_1858,N_428,N_795);
and U1859 (N_1859,N_579,N_124);
nand U1860 (N_1860,N_729,N_734);
nand U1861 (N_1861,N_610,N_885);
or U1862 (N_1862,N_761,N_817);
nor U1863 (N_1863,N_103,N_483);
nand U1864 (N_1864,N_297,N_538);
nand U1865 (N_1865,N_581,N_997);
and U1866 (N_1866,N_391,N_948);
or U1867 (N_1867,N_622,N_893);
nand U1868 (N_1868,N_473,N_286);
nor U1869 (N_1869,N_548,N_943);
or U1870 (N_1870,N_967,N_928);
and U1871 (N_1871,N_221,N_774);
or U1872 (N_1872,N_473,N_298);
and U1873 (N_1873,N_325,N_350);
nand U1874 (N_1874,N_133,N_277);
or U1875 (N_1875,N_341,N_34);
or U1876 (N_1876,N_358,N_642);
nand U1877 (N_1877,N_27,N_981);
xnor U1878 (N_1878,N_64,N_462);
or U1879 (N_1879,N_222,N_376);
and U1880 (N_1880,N_651,N_601);
or U1881 (N_1881,N_44,N_829);
and U1882 (N_1882,N_53,N_349);
and U1883 (N_1883,N_468,N_91);
nor U1884 (N_1884,N_758,N_355);
and U1885 (N_1885,N_740,N_229);
and U1886 (N_1886,N_479,N_902);
nor U1887 (N_1887,N_36,N_700);
or U1888 (N_1888,N_717,N_782);
and U1889 (N_1889,N_966,N_498);
nand U1890 (N_1890,N_466,N_710);
or U1891 (N_1891,N_841,N_280);
or U1892 (N_1892,N_884,N_861);
nor U1893 (N_1893,N_442,N_987);
and U1894 (N_1894,N_743,N_907);
xor U1895 (N_1895,N_311,N_786);
and U1896 (N_1896,N_739,N_631);
xor U1897 (N_1897,N_507,N_912);
nand U1898 (N_1898,N_59,N_625);
or U1899 (N_1899,N_922,N_250);
nand U1900 (N_1900,N_902,N_658);
nand U1901 (N_1901,N_84,N_507);
or U1902 (N_1902,N_971,N_360);
nand U1903 (N_1903,N_520,N_769);
nand U1904 (N_1904,N_648,N_952);
and U1905 (N_1905,N_830,N_930);
nand U1906 (N_1906,N_947,N_188);
nor U1907 (N_1907,N_932,N_532);
and U1908 (N_1908,N_778,N_425);
and U1909 (N_1909,N_944,N_629);
nand U1910 (N_1910,N_508,N_652);
nor U1911 (N_1911,N_564,N_272);
or U1912 (N_1912,N_832,N_527);
xor U1913 (N_1913,N_407,N_959);
nand U1914 (N_1914,N_2,N_749);
nand U1915 (N_1915,N_413,N_644);
nor U1916 (N_1916,N_56,N_414);
or U1917 (N_1917,N_832,N_113);
nand U1918 (N_1918,N_316,N_133);
or U1919 (N_1919,N_776,N_239);
or U1920 (N_1920,N_885,N_673);
nor U1921 (N_1921,N_182,N_351);
nand U1922 (N_1922,N_468,N_418);
nor U1923 (N_1923,N_528,N_9);
and U1924 (N_1924,N_283,N_687);
xor U1925 (N_1925,N_778,N_758);
nand U1926 (N_1926,N_549,N_87);
or U1927 (N_1927,N_87,N_125);
nand U1928 (N_1928,N_427,N_670);
and U1929 (N_1929,N_64,N_435);
nand U1930 (N_1930,N_514,N_553);
or U1931 (N_1931,N_779,N_196);
or U1932 (N_1932,N_493,N_333);
nor U1933 (N_1933,N_767,N_421);
and U1934 (N_1934,N_693,N_9);
or U1935 (N_1935,N_14,N_279);
nor U1936 (N_1936,N_748,N_413);
and U1937 (N_1937,N_317,N_201);
nor U1938 (N_1938,N_788,N_439);
and U1939 (N_1939,N_781,N_652);
nand U1940 (N_1940,N_110,N_10);
xnor U1941 (N_1941,N_532,N_862);
nand U1942 (N_1942,N_209,N_649);
nand U1943 (N_1943,N_220,N_955);
nor U1944 (N_1944,N_64,N_150);
or U1945 (N_1945,N_933,N_313);
nor U1946 (N_1946,N_271,N_766);
nand U1947 (N_1947,N_460,N_687);
or U1948 (N_1948,N_840,N_250);
nand U1949 (N_1949,N_203,N_985);
or U1950 (N_1950,N_245,N_135);
and U1951 (N_1951,N_607,N_272);
or U1952 (N_1952,N_131,N_692);
nand U1953 (N_1953,N_849,N_205);
and U1954 (N_1954,N_884,N_286);
xnor U1955 (N_1955,N_255,N_81);
nor U1956 (N_1956,N_431,N_734);
and U1957 (N_1957,N_4,N_305);
xnor U1958 (N_1958,N_402,N_590);
nor U1959 (N_1959,N_530,N_94);
or U1960 (N_1960,N_954,N_801);
or U1961 (N_1961,N_278,N_230);
nand U1962 (N_1962,N_106,N_988);
or U1963 (N_1963,N_87,N_31);
nor U1964 (N_1964,N_281,N_506);
or U1965 (N_1965,N_315,N_621);
nor U1966 (N_1966,N_512,N_992);
or U1967 (N_1967,N_499,N_932);
nor U1968 (N_1968,N_368,N_231);
nor U1969 (N_1969,N_710,N_437);
or U1970 (N_1970,N_450,N_274);
and U1971 (N_1971,N_313,N_664);
or U1972 (N_1972,N_169,N_474);
or U1973 (N_1973,N_209,N_842);
xnor U1974 (N_1974,N_741,N_687);
xor U1975 (N_1975,N_358,N_795);
and U1976 (N_1976,N_828,N_331);
nand U1977 (N_1977,N_665,N_357);
nand U1978 (N_1978,N_267,N_480);
and U1979 (N_1979,N_915,N_117);
xnor U1980 (N_1980,N_304,N_971);
nor U1981 (N_1981,N_823,N_199);
and U1982 (N_1982,N_647,N_726);
nand U1983 (N_1983,N_38,N_959);
and U1984 (N_1984,N_624,N_724);
and U1985 (N_1985,N_131,N_372);
and U1986 (N_1986,N_913,N_391);
or U1987 (N_1987,N_393,N_812);
and U1988 (N_1988,N_514,N_988);
and U1989 (N_1989,N_949,N_575);
nor U1990 (N_1990,N_5,N_100);
nor U1991 (N_1991,N_117,N_120);
or U1992 (N_1992,N_758,N_570);
or U1993 (N_1993,N_504,N_886);
and U1994 (N_1994,N_898,N_987);
nor U1995 (N_1995,N_888,N_444);
and U1996 (N_1996,N_896,N_200);
or U1997 (N_1997,N_811,N_506);
xor U1998 (N_1998,N_198,N_733);
nor U1999 (N_1999,N_125,N_141);
or U2000 (N_2000,N_1841,N_1079);
or U2001 (N_2001,N_1758,N_1929);
nand U2002 (N_2002,N_1838,N_1702);
nand U2003 (N_2003,N_1052,N_1212);
or U2004 (N_2004,N_1798,N_1021);
and U2005 (N_2005,N_1107,N_1770);
and U2006 (N_2006,N_1144,N_1966);
nand U2007 (N_2007,N_1100,N_1587);
and U2008 (N_2008,N_1179,N_1069);
nand U2009 (N_2009,N_1258,N_1676);
and U2010 (N_2010,N_1771,N_1589);
nand U2011 (N_2011,N_1633,N_1506);
or U2012 (N_2012,N_1397,N_1572);
nand U2013 (N_2013,N_1973,N_1960);
nor U2014 (N_2014,N_1666,N_1140);
and U2015 (N_2015,N_1224,N_1034);
or U2016 (N_2016,N_1521,N_1690);
nand U2017 (N_2017,N_1169,N_1201);
and U2018 (N_2018,N_1090,N_1428);
nand U2019 (N_2019,N_1736,N_1080);
and U2020 (N_2020,N_1136,N_1714);
or U2021 (N_2021,N_1309,N_1543);
or U2022 (N_2022,N_1157,N_1256);
and U2023 (N_2023,N_1989,N_1307);
and U2024 (N_2024,N_1265,N_1259);
nor U2025 (N_2025,N_1434,N_1796);
nor U2026 (N_2026,N_1363,N_1708);
and U2027 (N_2027,N_1367,N_1723);
or U2028 (N_2028,N_1431,N_1767);
or U2029 (N_2029,N_1848,N_1815);
or U2030 (N_2030,N_1358,N_1691);
or U2031 (N_2031,N_1790,N_1583);
nand U2032 (N_2032,N_1246,N_1555);
nor U2033 (N_2033,N_1113,N_1284);
or U2034 (N_2034,N_1772,N_1406);
and U2035 (N_2035,N_1316,N_1834);
and U2036 (N_2036,N_1833,N_1025);
nand U2037 (N_2037,N_1131,N_1682);
or U2038 (N_2038,N_1049,N_1922);
nor U2039 (N_2039,N_1083,N_1882);
nor U2040 (N_2040,N_1002,N_1713);
nand U2041 (N_2041,N_1400,N_1409);
or U2042 (N_2042,N_1156,N_1740);
or U2043 (N_2043,N_1031,N_1963);
nand U2044 (N_2044,N_1374,N_1875);
and U2045 (N_2045,N_1361,N_1436);
or U2046 (N_2046,N_1219,N_1077);
and U2047 (N_2047,N_1383,N_1119);
or U2048 (N_2048,N_1563,N_1500);
or U2049 (N_2049,N_1171,N_1896);
or U2050 (N_2050,N_1485,N_1032);
and U2051 (N_2051,N_1540,N_1218);
and U2052 (N_2052,N_1186,N_1151);
nand U2053 (N_2053,N_1920,N_1782);
nand U2054 (N_2054,N_1961,N_1055);
nor U2055 (N_2055,N_1104,N_1884);
nand U2056 (N_2056,N_1202,N_1451);
nor U2057 (N_2057,N_1338,N_1108);
nor U2058 (N_2058,N_1921,N_1611);
nor U2059 (N_2059,N_1362,N_1698);
nand U2060 (N_2060,N_1864,N_1480);
nand U2061 (N_2061,N_1588,N_1162);
and U2062 (N_2062,N_1483,N_1250);
and U2063 (N_2063,N_1347,N_1948);
and U2064 (N_2064,N_1757,N_1412);
or U2065 (N_2065,N_1011,N_1554);
nor U2066 (N_2066,N_1445,N_1659);
nand U2067 (N_2067,N_1733,N_1275);
or U2068 (N_2068,N_1334,N_1649);
and U2069 (N_2069,N_1881,N_1597);
nor U2070 (N_2070,N_1170,N_1674);
nand U2071 (N_2071,N_1575,N_1797);
nor U2072 (N_2072,N_1773,N_1139);
and U2073 (N_2073,N_1840,N_1203);
nor U2074 (N_2074,N_1695,N_1949);
or U2075 (N_2075,N_1335,N_1780);
nand U2076 (N_2076,N_1868,N_1035);
nand U2077 (N_2077,N_1985,N_1135);
or U2078 (N_2078,N_1742,N_1152);
and U2079 (N_2079,N_1784,N_1376);
or U2080 (N_2080,N_1274,N_1125);
or U2081 (N_2081,N_1624,N_1082);
nor U2082 (N_2082,N_1356,N_1054);
and U2083 (N_2083,N_1225,N_1228);
nand U2084 (N_2084,N_1579,N_1769);
nand U2085 (N_2085,N_1290,N_1147);
nand U2086 (N_2086,N_1298,N_1000);
nand U2087 (N_2087,N_1972,N_1626);
and U2088 (N_2088,N_1822,N_1574);
nand U2089 (N_2089,N_1941,N_1635);
and U2090 (N_2090,N_1053,N_1689);
or U2091 (N_2091,N_1737,N_1877);
and U2092 (N_2092,N_1405,N_1026);
or U2093 (N_2093,N_1014,N_1093);
nor U2094 (N_2094,N_1092,N_1600);
or U2095 (N_2095,N_1515,N_1775);
nor U2096 (N_2096,N_1590,N_1109);
nand U2097 (N_2097,N_1295,N_1291);
nand U2098 (N_2098,N_1852,N_1824);
or U2099 (N_2099,N_1622,N_1384);
nand U2100 (N_2100,N_1488,N_1242);
nor U2101 (N_2101,N_1793,N_1806);
or U2102 (N_2102,N_1399,N_1191);
nor U2103 (N_2103,N_1296,N_1519);
nor U2104 (N_2104,N_1925,N_1774);
xor U2105 (N_2105,N_1394,N_1876);
nand U2106 (N_2106,N_1816,N_1892);
and U2107 (N_2107,N_1208,N_1024);
and U2108 (N_2108,N_1102,N_1509);
and U2109 (N_2109,N_1781,N_1177);
or U2110 (N_2110,N_1042,N_1438);
nand U2111 (N_2111,N_1990,N_1762);
or U2112 (N_2112,N_1282,N_1235);
nand U2113 (N_2113,N_1819,N_1879);
nand U2114 (N_2114,N_1680,N_1971);
or U2115 (N_2115,N_1988,N_1992);
and U2116 (N_2116,N_1283,N_1732);
and U2117 (N_2117,N_1305,N_1349);
or U2118 (N_2118,N_1491,N_1752);
nor U2119 (N_2119,N_1463,N_1914);
or U2120 (N_2120,N_1878,N_1594);
or U2121 (N_2121,N_1905,N_1580);
or U2122 (N_2122,N_1684,N_1748);
and U2123 (N_2123,N_1312,N_1755);
or U2124 (N_2124,N_1127,N_1598);
or U2125 (N_2125,N_1655,N_1663);
nand U2126 (N_2126,N_1789,N_1984);
nor U2127 (N_2127,N_1422,N_1413);
nor U2128 (N_2128,N_1210,N_1226);
or U2129 (N_2129,N_1023,N_1814);
or U2130 (N_2130,N_1716,N_1459);
or U2131 (N_2131,N_1541,N_1527);
or U2132 (N_2132,N_1846,N_1919);
and U2133 (N_2133,N_1621,N_1869);
or U2134 (N_2134,N_1371,N_1074);
nor U2135 (N_2135,N_1350,N_1280);
and U2136 (N_2136,N_1469,N_1458);
nand U2137 (N_2137,N_1322,N_1811);
and U2138 (N_2138,N_1160,N_1526);
nor U2139 (N_2139,N_1936,N_1658);
xor U2140 (N_2140,N_1545,N_1013);
nand U2141 (N_2141,N_1452,N_1324);
or U2142 (N_2142,N_1453,N_1874);
nor U2143 (N_2143,N_1724,N_1730);
and U2144 (N_2144,N_1880,N_1620);
and U2145 (N_2145,N_1951,N_1918);
nor U2146 (N_2146,N_1234,N_1533);
nor U2147 (N_2147,N_1665,N_1373);
and U2148 (N_2148,N_1681,N_1262);
or U2149 (N_2149,N_1154,N_1206);
nor U2150 (N_2150,N_1101,N_1381);
or U2151 (N_2151,N_1516,N_1553);
nand U2152 (N_2152,N_1245,N_1071);
nand U2153 (N_2153,N_1576,N_1940);
nand U2154 (N_2154,N_1244,N_1289);
nor U2155 (N_2155,N_1184,N_1567);
xnor U2156 (N_2156,N_1703,N_1474);
nand U2157 (N_2157,N_1308,N_1717);
or U2158 (N_2158,N_1027,N_1530);
and U2159 (N_2159,N_1236,N_1067);
and U2160 (N_2160,N_1986,N_1855);
and U2161 (N_2161,N_1634,N_1022);
nand U2162 (N_2162,N_1222,N_1660);
nor U2163 (N_2163,N_1970,N_1872);
or U2164 (N_2164,N_1043,N_1496);
nor U2165 (N_2165,N_1562,N_1685);
and U2166 (N_2166,N_1697,N_1865);
nor U2167 (N_2167,N_1860,N_1435);
and U2168 (N_2168,N_1085,N_1099);
and U2169 (N_2169,N_1686,N_1327);
and U2170 (N_2170,N_1639,N_1417);
nor U2171 (N_2171,N_1299,N_1803);
and U2172 (N_2172,N_1999,N_1954);
nor U2173 (N_2173,N_1552,N_1075);
or U2174 (N_2174,N_1835,N_1938);
xnor U2175 (N_2175,N_1292,N_1277);
or U2176 (N_2176,N_1839,N_1895);
nand U2177 (N_2177,N_1694,N_1087);
nor U2178 (N_2178,N_1336,N_1549);
and U2179 (N_2179,N_1411,N_1913);
nand U2180 (N_2180,N_1243,N_1965);
nand U2181 (N_2181,N_1706,N_1486);
nor U2182 (N_2182,N_1903,N_1754);
and U2183 (N_2183,N_1566,N_1030);
and U2184 (N_2184,N_1492,N_1517);
nor U2185 (N_2185,N_1227,N_1640);
nand U2186 (N_2186,N_1612,N_1204);
nand U2187 (N_2187,N_1785,N_1181);
xnor U2188 (N_2188,N_1433,N_1904);
nor U2189 (N_2189,N_1176,N_1270);
nor U2190 (N_2190,N_1461,N_1651);
and U2191 (N_2191,N_1637,N_1539);
nand U2192 (N_2192,N_1328,N_1481);
or U2193 (N_2193,N_1707,N_1871);
nand U2194 (N_2194,N_1489,N_1462);
nand U2195 (N_2195,N_1098,N_1375);
nor U2196 (N_2196,N_1173,N_1126);
or U2197 (N_2197,N_1393,N_1091);
and U2198 (N_2198,N_1163,N_1033);
or U2199 (N_2199,N_1110,N_1189);
nor U2200 (N_2200,N_1040,N_1573);
nor U2201 (N_2201,N_1821,N_1370);
xor U2202 (N_2202,N_1380,N_1546);
nor U2203 (N_2203,N_1536,N_1502);
and U2204 (N_2204,N_1595,N_1609);
and U2205 (N_2205,N_1508,N_1858);
and U2206 (N_2206,N_1130,N_1669);
and U2207 (N_2207,N_1942,N_1190);
nand U2208 (N_2208,N_1355,N_1894);
nor U2209 (N_2209,N_1143,N_1047);
nor U2210 (N_2210,N_1642,N_1410);
and U2211 (N_2211,N_1060,N_1885);
or U2212 (N_2212,N_1494,N_1269);
and U2213 (N_2213,N_1995,N_1571);
nor U2214 (N_2214,N_1512,N_1746);
nor U2215 (N_2215,N_1631,N_1801);
or U2216 (N_2216,N_1267,N_1252);
nand U2217 (N_2217,N_1537,N_1072);
nand U2218 (N_2218,N_1388,N_1873);
and U2219 (N_2219,N_1808,N_1018);
or U2220 (N_2220,N_1357,N_1667);
and U2221 (N_2221,N_1472,N_1661);
nor U2222 (N_2222,N_1331,N_1231);
nor U2223 (N_2223,N_1711,N_1182);
and U2224 (N_2224,N_1854,N_1997);
nand U2225 (N_2225,N_1271,N_1809);
and U2226 (N_2226,N_1619,N_1365);
and U2227 (N_2227,N_1968,N_1128);
nor U2228 (N_2228,N_1983,N_1395);
nor U2229 (N_2229,N_1342,N_1439);
nand U2230 (N_2230,N_1741,N_1120);
and U2231 (N_2231,N_1129,N_1542);
nand U2232 (N_2232,N_1215,N_1715);
nor U2233 (N_2233,N_1476,N_1323);
or U2234 (N_2234,N_1825,N_1856);
nand U2235 (N_2235,N_1933,N_1029);
nand U2236 (N_2236,N_1550,N_1240);
nand U2237 (N_2237,N_1247,N_1578);
and U2238 (N_2238,N_1263,N_1321);
nand U2239 (N_2239,N_1149,N_1504);
and U2240 (N_2240,N_1310,N_1205);
nor U2241 (N_2241,N_1443,N_1890);
or U2242 (N_2242,N_1828,N_1705);
or U2243 (N_2243,N_1041,N_1337);
and U2244 (N_2244,N_1065,N_1786);
or U2245 (N_2245,N_1664,N_1341);
or U2246 (N_2246,N_1981,N_1910);
nor U2247 (N_2247,N_1487,N_1241);
and U2248 (N_2248,N_1721,N_1863);
nand U2249 (N_2249,N_1939,N_1534);
xnor U2250 (N_2250,N_1427,N_1223);
or U2251 (N_2251,N_1297,N_1329);
nor U2252 (N_2252,N_1407,N_1001);
or U2253 (N_2253,N_1340,N_1844);
and U2254 (N_2254,N_1471,N_1582);
nor U2255 (N_2255,N_1103,N_1165);
nand U2256 (N_2256,N_1759,N_1617);
nand U2257 (N_2257,N_1192,N_1490);
nor U2258 (N_2258,N_1194,N_1294);
nand U2259 (N_2259,N_1548,N_1729);
or U2260 (N_2260,N_1012,N_1264);
or U2261 (N_2261,N_1673,N_1800);
or U2262 (N_2262,N_1636,N_1853);
and U2263 (N_2263,N_1301,N_1314);
nand U2264 (N_2264,N_1947,N_1532);
and U2265 (N_2265,N_1187,N_1657);
or U2266 (N_2266,N_1048,N_1004);
nor U2267 (N_2267,N_1088,N_1996);
or U2268 (N_2268,N_1449,N_1086);
and U2269 (N_2269,N_1339,N_1134);
nor U2270 (N_2270,N_1306,N_1286);
or U2271 (N_2271,N_1006,N_1348);
nand U2272 (N_2272,N_1095,N_1912);
or U2273 (N_2273,N_1710,N_1429);
nand U2274 (N_2274,N_1261,N_1020);
nand U2275 (N_2275,N_1056,N_1569);
and U2276 (N_2276,N_1776,N_1902);
nand U2277 (N_2277,N_1836,N_1112);
nand U2278 (N_2278,N_1805,N_1221);
or U2279 (N_2279,N_1867,N_1505);
and U2280 (N_2280,N_1911,N_1039);
or U2281 (N_2281,N_1473,N_1503);
nor U2282 (N_2282,N_1213,N_1899);
nand U2283 (N_2283,N_1401,N_1368);
nor U2284 (N_2284,N_1354,N_1254);
and U2285 (N_2285,N_1010,N_1420);
nor U2286 (N_2286,N_1081,N_1584);
nor U2287 (N_2287,N_1084,N_1209);
nand U2288 (N_2288,N_1994,N_1416);
and U2289 (N_2289,N_1618,N_1288);
xor U2290 (N_2290,N_1217,N_1607);
nand U2291 (N_2291,N_1843,N_1253);
nand U2292 (N_2292,N_1330,N_1313);
and U2293 (N_2293,N_1544,N_1302);
nand U2294 (N_2294,N_1830,N_1106);
or U2295 (N_2295,N_1638,N_1118);
and U2296 (N_2296,N_1058,N_1722);
nor U2297 (N_2297,N_1565,N_1870);
nor U2298 (N_2298,N_1564,N_1200);
nor U2299 (N_2299,N_1279,N_1538);
nand U2300 (N_2300,N_1096,N_1470);
nor U2301 (N_2301,N_1076,N_1391);
or U2302 (N_2302,N_1662,N_1479);
or U2303 (N_2303,N_1482,N_1671);
nand U2304 (N_2304,N_1237,N_1761);
nand U2305 (N_2305,N_1560,N_1248);
and U2306 (N_2306,N_1851,N_1211);
or U2307 (N_2307,N_1753,N_1728);
nand U2308 (N_2308,N_1141,N_1688);
nor U2309 (N_2309,N_1807,N_1017);
nand U2310 (N_2310,N_1514,N_1117);
or U2311 (N_2311,N_1137,N_1377);
nor U2312 (N_2312,N_1064,N_1003);
nand U2313 (N_2313,N_1352,N_1063);
and U2314 (N_2314,N_1734,N_1382);
or U2315 (N_2315,N_1628,N_1008);
nor U2316 (N_2316,N_1278,N_1557);
or U2317 (N_2317,N_1944,N_1826);
and U2318 (N_2318,N_1440,N_1709);
nor U2319 (N_2319,N_1111,N_1561);
nor U2320 (N_2320,N_1180,N_1608);
and U2321 (N_2321,N_1178,N_1007);
or U2322 (N_2322,N_1791,N_1955);
nor U2323 (N_2323,N_1158,N_1887);
nor U2324 (N_2324,N_1677,N_1326);
and U2325 (N_2325,N_1656,N_1727);
or U2326 (N_2326,N_1498,N_1332);
or U2327 (N_2327,N_1132,N_1764);
nand U2328 (N_2328,N_1820,N_1168);
or U2329 (N_2329,N_1518,N_1456);
nor U2330 (N_2330,N_1842,N_1345);
and U2331 (N_2331,N_1794,N_1418);
and U2332 (N_2332,N_1847,N_1898);
nor U2333 (N_2333,N_1568,N_1699);
nor U2334 (N_2334,N_1603,N_1585);
nand U2335 (N_2335,N_1744,N_1447);
nand U2336 (N_2336,N_1344,N_1037);
and U2337 (N_2337,N_1059,N_1028);
nand U2338 (N_2338,N_1934,N_1251);
nand U2339 (N_2339,N_1946,N_1950);
nor U2340 (N_2340,N_1760,N_1317);
nor U2341 (N_2341,N_1991,N_1005);
nand U2342 (N_2342,N_1943,N_1045);
or U2343 (N_2343,N_1398,N_1195);
or U2344 (N_2344,N_1792,N_1450);
nor U2345 (N_2345,N_1679,N_1813);
and U2346 (N_2346,N_1507,N_1862);
and U2347 (N_2347,N_1756,N_1351);
and U2348 (N_2348,N_1146,N_1378);
nand U2349 (N_2349,N_1610,N_1493);
or U2350 (N_2350,N_1718,N_1094);
nor U2351 (N_2351,N_1229,N_1387);
and U2352 (N_2352,N_1446,N_1731);
nor U2353 (N_2353,N_1893,N_1325);
nand U2354 (N_2354,N_1379,N_1959);
xor U2355 (N_2355,N_1467,N_1672);
and U2356 (N_2356,N_1057,N_1592);
and U2357 (N_2357,N_1167,N_1523);
nor U2358 (N_2358,N_1061,N_1886);
nor U2359 (N_2359,N_1883,N_1935);
and U2360 (N_2360,N_1645,N_1632);
nand U2361 (N_2361,N_1799,N_1788);
or U2362 (N_2362,N_1531,N_1964);
and U2363 (N_2363,N_1460,N_1926);
nor U2364 (N_2364,N_1923,N_1425);
or U2365 (N_2365,N_1304,N_1977);
or U2366 (N_2366,N_1625,N_1745);
or U2367 (N_2367,N_1696,N_1148);
nand U2368 (N_2368,N_1272,N_1802);
nor U2369 (N_2369,N_1457,N_1372);
nor U2370 (N_2370,N_1535,N_1551);
xnor U2371 (N_2371,N_1359,N_1596);
and U2372 (N_2372,N_1787,N_1817);
or U2373 (N_2373,N_1627,N_1524);
and U2374 (N_2374,N_1866,N_1408);
nand U2375 (N_2375,N_1924,N_1046);
or U2376 (N_2376,N_1980,N_1581);
nor U2377 (N_2377,N_1392,N_1646);
nor U2378 (N_2378,N_1448,N_1888);
or U2379 (N_2379,N_1525,N_1464);
and U2380 (N_2380,N_1454,N_1547);
nand U2381 (N_2381,N_1174,N_1138);
or U2382 (N_2382,N_1166,N_1068);
nor U2383 (N_2383,N_1155,N_1386);
or U2384 (N_2384,N_1593,N_1232);
and U2385 (N_2385,N_1268,N_1993);
nand U2386 (N_2386,N_1937,N_1750);
nand U2387 (N_2387,N_1164,N_1257);
nand U2388 (N_2388,N_1601,N_1315);
nand U2389 (N_2389,N_1570,N_1804);
and U2390 (N_2390,N_1987,N_1693);
or U2391 (N_2391,N_1444,N_1906);
nor U2392 (N_2392,N_1038,N_1749);
nor U2393 (N_2393,N_1604,N_1908);
and U2394 (N_2394,N_1930,N_1832);
and U2395 (N_2395,N_1123,N_1145);
nand U2396 (N_2396,N_1115,N_1073);
or U2397 (N_2397,N_1396,N_1743);
and U2398 (N_2398,N_1931,N_1404);
nor U2399 (N_2399,N_1795,N_1974);
nand U2400 (N_2400,N_1777,N_1738);
or U2401 (N_2401,N_1239,N_1692);
or U2402 (N_2402,N_1150,N_1653);
or U2403 (N_2403,N_1207,N_1050);
or U2404 (N_2404,N_1293,N_1105);
nand U2405 (N_2405,N_1441,N_1962);
nand U2406 (N_2406,N_1605,N_1078);
or U2407 (N_2407,N_1917,N_1122);
and U2408 (N_2408,N_1630,N_1285);
or U2409 (N_2409,N_1066,N_1818);
nand U2410 (N_2410,N_1779,N_1648);
and U2411 (N_2411,N_1916,N_1153);
nor U2412 (N_2412,N_1199,N_1810);
and U2413 (N_2413,N_1586,N_1238);
or U2414 (N_2414,N_1214,N_1982);
and U2415 (N_2415,N_1193,N_1366);
and U2416 (N_2416,N_1495,N_1513);
nor U2417 (N_2417,N_1455,N_1114);
or U2418 (N_2418,N_1421,N_1683);
nor U2419 (N_2419,N_1629,N_1124);
and U2420 (N_2420,N_1390,N_1556);
and U2421 (N_2421,N_1089,N_1142);
nor U2422 (N_2422,N_1829,N_1499);
nor U2423 (N_2423,N_1320,N_1812);
nor U2424 (N_2424,N_1303,N_1121);
and U2425 (N_2425,N_1185,N_1281);
and U2426 (N_2426,N_1998,N_1650);
and U2427 (N_2427,N_1465,N_1602);
nand U2428 (N_2428,N_1319,N_1712);
nand U2429 (N_2429,N_1778,N_1389);
nor U2430 (N_2430,N_1528,N_1343);
nand U2431 (N_2431,N_1850,N_1466);
nor U2432 (N_2432,N_1747,N_1837);
nand U2433 (N_2433,N_1070,N_1701);
nand U2434 (N_2434,N_1558,N_1196);
and U2435 (N_2435,N_1360,N_1402);
and U2436 (N_2436,N_1720,N_1385);
or U2437 (N_2437,N_1197,N_1019);
nand U2438 (N_2438,N_1953,N_1654);
or U2439 (N_2439,N_1364,N_1675);
nor U2440 (N_2440,N_1520,N_1249);
and U2441 (N_2441,N_1051,N_1415);
nand U2442 (N_2442,N_1591,N_1932);
nor U2443 (N_2443,N_1423,N_1900);
and U2444 (N_2444,N_1907,N_1751);
and U2445 (N_2445,N_1432,N_1857);
nor U2446 (N_2446,N_1198,N_1188);
and U2447 (N_2447,N_1845,N_1353);
nor U2448 (N_2448,N_1260,N_1172);
and U2449 (N_2449,N_1015,N_1009);
nand U2450 (N_2450,N_1735,N_1097);
nand U2451 (N_2451,N_1159,N_1062);
or U2452 (N_2452,N_1497,N_1958);
nor U2453 (N_2453,N_1036,N_1599);
or U2454 (N_2454,N_1700,N_1901);
and U2455 (N_2455,N_1957,N_1670);
or U2456 (N_2456,N_1969,N_1529);
and U2457 (N_2457,N_1273,N_1927);
or U2458 (N_2458,N_1623,N_1719);
nor U2459 (N_2459,N_1976,N_1255);
nor U2460 (N_2460,N_1511,N_1823);
or U2461 (N_2461,N_1403,N_1928);
and U2462 (N_2462,N_1501,N_1766);
nand U2463 (N_2463,N_1945,N_1644);
nor U2464 (N_2464,N_1311,N_1442);
nor U2465 (N_2465,N_1510,N_1175);
or U2466 (N_2466,N_1652,N_1704);
and U2467 (N_2467,N_1559,N_1468);
nor U2468 (N_2468,N_1230,N_1116);
and U2469 (N_2469,N_1419,N_1909);
nor U2470 (N_2470,N_1016,N_1889);
or U2471 (N_2471,N_1739,N_1161);
xor U2472 (N_2472,N_1726,N_1216);
nor U2473 (N_2473,N_1967,N_1827);
and U2474 (N_2474,N_1369,N_1266);
nand U2475 (N_2475,N_1276,N_1783);
nor U2476 (N_2476,N_1424,N_1831);
nand U2477 (N_2477,N_1133,N_1430);
and U2478 (N_2478,N_1956,N_1915);
or U2479 (N_2479,N_1346,N_1859);
nand U2480 (N_2480,N_1765,N_1615);
nor U2481 (N_2481,N_1414,N_1437);
nand U2482 (N_2482,N_1220,N_1478);
and U2483 (N_2483,N_1687,N_1849);
or U2484 (N_2484,N_1725,N_1768);
nor U2485 (N_2485,N_1484,N_1975);
nand U2486 (N_2486,N_1333,N_1287);
or U2487 (N_2487,N_1891,N_1044);
nor U2488 (N_2488,N_1475,N_1643);
or U2489 (N_2489,N_1641,N_1979);
or U2490 (N_2490,N_1897,N_1318);
or U2491 (N_2491,N_1678,N_1861);
and U2492 (N_2492,N_1668,N_1577);
and U2493 (N_2493,N_1763,N_1477);
and U2494 (N_2494,N_1233,N_1978);
nor U2495 (N_2495,N_1614,N_1952);
or U2496 (N_2496,N_1183,N_1522);
nand U2497 (N_2497,N_1426,N_1616);
nand U2498 (N_2498,N_1300,N_1647);
and U2499 (N_2499,N_1606,N_1613);
xor U2500 (N_2500,N_1650,N_1611);
nor U2501 (N_2501,N_1983,N_1034);
and U2502 (N_2502,N_1559,N_1624);
or U2503 (N_2503,N_1820,N_1963);
nor U2504 (N_2504,N_1305,N_1897);
nor U2505 (N_2505,N_1227,N_1706);
or U2506 (N_2506,N_1707,N_1011);
and U2507 (N_2507,N_1941,N_1016);
nand U2508 (N_2508,N_1431,N_1592);
nand U2509 (N_2509,N_1061,N_1183);
or U2510 (N_2510,N_1490,N_1045);
and U2511 (N_2511,N_1663,N_1064);
nand U2512 (N_2512,N_1691,N_1553);
nand U2513 (N_2513,N_1705,N_1895);
nor U2514 (N_2514,N_1707,N_1121);
or U2515 (N_2515,N_1695,N_1223);
and U2516 (N_2516,N_1855,N_1518);
nand U2517 (N_2517,N_1251,N_1590);
xor U2518 (N_2518,N_1451,N_1705);
and U2519 (N_2519,N_1164,N_1779);
nor U2520 (N_2520,N_1661,N_1901);
nor U2521 (N_2521,N_1931,N_1701);
xnor U2522 (N_2522,N_1055,N_1449);
nand U2523 (N_2523,N_1350,N_1877);
or U2524 (N_2524,N_1052,N_1241);
and U2525 (N_2525,N_1618,N_1037);
and U2526 (N_2526,N_1021,N_1633);
nand U2527 (N_2527,N_1701,N_1376);
and U2528 (N_2528,N_1987,N_1738);
nand U2529 (N_2529,N_1575,N_1350);
nand U2530 (N_2530,N_1902,N_1522);
nor U2531 (N_2531,N_1450,N_1978);
or U2532 (N_2532,N_1391,N_1781);
and U2533 (N_2533,N_1029,N_1140);
and U2534 (N_2534,N_1898,N_1069);
and U2535 (N_2535,N_1191,N_1806);
or U2536 (N_2536,N_1783,N_1412);
xnor U2537 (N_2537,N_1166,N_1039);
or U2538 (N_2538,N_1005,N_1471);
and U2539 (N_2539,N_1376,N_1162);
or U2540 (N_2540,N_1045,N_1481);
and U2541 (N_2541,N_1334,N_1827);
or U2542 (N_2542,N_1644,N_1794);
nand U2543 (N_2543,N_1716,N_1473);
or U2544 (N_2544,N_1524,N_1134);
nor U2545 (N_2545,N_1174,N_1087);
or U2546 (N_2546,N_1459,N_1020);
nand U2547 (N_2547,N_1107,N_1774);
or U2548 (N_2548,N_1070,N_1861);
nor U2549 (N_2549,N_1546,N_1289);
and U2550 (N_2550,N_1845,N_1965);
nand U2551 (N_2551,N_1508,N_1465);
nor U2552 (N_2552,N_1770,N_1182);
or U2553 (N_2553,N_1560,N_1763);
nand U2554 (N_2554,N_1040,N_1398);
nor U2555 (N_2555,N_1110,N_1848);
nor U2556 (N_2556,N_1682,N_1334);
xor U2557 (N_2557,N_1355,N_1566);
nand U2558 (N_2558,N_1017,N_1745);
or U2559 (N_2559,N_1840,N_1791);
and U2560 (N_2560,N_1590,N_1862);
nand U2561 (N_2561,N_1221,N_1068);
or U2562 (N_2562,N_1243,N_1019);
nand U2563 (N_2563,N_1801,N_1987);
nor U2564 (N_2564,N_1246,N_1731);
xnor U2565 (N_2565,N_1936,N_1982);
nor U2566 (N_2566,N_1174,N_1992);
nand U2567 (N_2567,N_1555,N_1051);
nor U2568 (N_2568,N_1117,N_1050);
or U2569 (N_2569,N_1713,N_1290);
or U2570 (N_2570,N_1210,N_1013);
nor U2571 (N_2571,N_1107,N_1450);
nand U2572 (N_2572,N_1527,N_1841);
and U2573 (N_2573,N_1028,N_1606);
or U2574 (N_2574,N_1146,N_1048);
nor U2575 (N_2575,N_1377,N_1988);
nand U2576 (N_2576,N_1023,N_1689);
nand U2577 (N_2577,N_1703,N_1018);
nand U2578 (N_2578,N_1195,N_1188);
nand U2579 (N_2579,N_1766,N_1653);
nand U2580 (N_2580,N_1932,N_1355);
xor U2581 (N_2581,N_1515,N_1672);
nand U2582 (N_2582,N_1350,N_1998);
nor U2583 (N_2583,N_1429,N_1376);
or U2584 (N_2584,N_1988,N_1969);
or U2585 (N_2585,N_1070,N_1772);
and U2586 (N_2586,N_1059,N_1435);
or U2587 (N_2587,N_1550,N_1392);
and U2588 (N_2588,N_1002,N_1174);
nand U2589 (N_2589,N_1349,N_1135);
nand U2590 (N_2590,N_1668,N_1425);
nor U2591 (N_2591,N_1762,N_1002);
and U2592 (N_2592,N_1011,N_1766);
nand U2593 (N_2593,N_1788,N_1021);
or U2594 (N_2594,N_1592,N_1346);
nor U2595 (N_2595,N_1809,N_1179);
or U2596 (N_2596,N_1092,N_1191);
nor U2597 (N_2597,N_1277,N_1813);
or U2598 (N_2598,N_1553,N_1355);
or U2599 (N_2599,N_1134,N_1263);
and U2600 (N_2600,N_1182,N_1210);
nand U2601 (N_2601,N_1929,N_1349);
and U2602 (N_2602,N_1707,N_1426);
or U2603 (N_2603,N_1075,N_1301);
nand U2604 (N_2604,N_1912,N_1637);
and U2605 (N_2605,N_1969,N_1962);
nand U2606 (N_2606,N_1885,N_1296);
or U2607 (N_2607,N_1140,N_1047);
nor U2608 (N_2608,N_1213,N_1112);
and U2609 (N_2609,N_1688,N_1091);
or U2610 (N_2610,N_1328,N_1635);
or U2611 (N_2611,N_1830,N_1743);
and U2612 (N_2612,N_1208,N_1676);
nor U2613 (N_2613,N_1745,N_1103);
nor U2614 (N_2614,N_1808,N_1820);
nand U2615 (N_2615,N_1816,N_1082);
nor U2616 (N_2616,N_1855,N_1924);
or U2617 (N_2617,N_1261,N_1408);
or U2618 (N_2618,N_1262,N_1724);
nand U2619 (N_2619,N_1509,N_1792);
nor U2620 (N_2620,N_1697,N_1500);
and U2621 (N_2621,N_1672,N_1311);
or U2622 (N_2622,N_1559,N_1760);
and U2623 (N_2623,N_1268,N_1502);
nor U2624 (N_2624,N_1100,N_1634);
or U2625 (N_2625,N_1278,N_1556);
or U2626 (N_2626,N_1607,N_1617);
and U2627 (N_2627,N_1187,N_1926);
and U2628 (N_2628,N_1821,N_1620);
and U2629 (N_2629,N_1551,N_1756);
nor U2630 (N_2630,N_1586,N_1026);
nor U2631 (N_2631,N_1757,N_1601);
xor U2632 (N_2632,N_1646,N_1699);
xor U2633 (N_2633,N_1819,N_1364);
nor U2634 (N_2634,N_1276,N_1124);
or U2635 (N_2635,N_1865,N_1308);
nand U2636 (N_2636,N_1103,N_1442);
or U2637 (N_2637,N_1772,N_1422);
nand U2638 (N_2638,N_1793,N_1366);
or U2639 (N_2639,N_1821,N_1835);
or U2640 (N_2640,N_1305,N_1723);
and U2641 (N_2641,N_1392,N_1505);
and U2642 (N_2642,N_1254,N_1806);
nand U2643 (N_2643,N_1099,N_1976);
and U2644 (N_2644,N_1485,N_1729);
nor U2645 (N_2645,N_1496,N_1172);
nor U2646 (N_2646,N_1983,N_1380);
or U2647 (N_2647,N_1823,N_1772);
nor U2648 (N_2648,N_1727,N_1035);
nand U2649 (N_2649,N_1107,N_1273);
nor U2650 (N_2650,N_1327,N_1034);
and U2651 (N_2651,N_1228,N_1763);
or U2652 (N_2652,N_1079,N_1835);
nand U2653 (N_2653,N_1391,N_1551);
or U2654 (N_2654,N_1319,N_1924);
nor U2655 (N_2655,N_1521,N_1995);
or U2656 (N_2656,N_1831,N_1853);
or U2657 (N_2657,N_1649,N_1111);
nand U2658 (N_2658,N_1598,N_1139);
nand U2659 (N_2659,N_1496,N_1171);
and U2660 (N_2660,N_1449,N_1830);
nor U2661 (N_2661,N_1360,N_1235);
and U2662 (N_2662,N_1798,N_1757);
nand U2663 (N_2663,N_1883,N_1531);
or U2664 (N_2664,N_1739,N_1652);
xnor U2665 (N_2665,N_1796,N_1190);
xnor U2666 (N_2666,N_1861,N_1995);
nand U2667 (N_2667,N_1233,N_1740);
nand U2668 (N_2668,N_1816,N_1377);
nand U2669 (N_2669,N_1491,N_1395);
nand U2670 (N_2670,N_1885,N_1373);
and U2671 (N_2671,N_1002,N_1926);
and U2672 (N_2672,N_1300,N_1061);
nand U2673 (N_2673,N_1410,N_1452);
nand U2674 (N_2674,N_1908,N_1483);
and U2675 (N_2675,N_1449,N_1464);
nor U2676 (N_2676,N_1409,N_1155);
nand U2677 (N_2677,N_1929,N_1634);
nor U2678 (N_2678,N_1817,N_1243);
or U2679 (N_2679,N_1241,N_1233);
nor U2680 (N_2680,N_1961,N_1369);
nand U2681 (N_2681,N_1006,N_1176);
nor U2682 (N_2682,N_1676,N_1119);
or U2683 (N_2683,N_1875,N_1190);
or U2684 (N_2684,N_1873,N_1346);
xor U2685 (N_2685,N_1922,N_1951);
or U2686 (N_2686,N_1819,N_1689);
nand U2687 (N_2687,N_1074,N_1852);
and U2688 (N_2688,N_1921,N_1362);
nand U2689 (N_2689,N_1562,N_1845);
nand U2690 (N_2690,N_1848,N_1584);
nor U2691 (N_2691,N_1853,N_1491);
or U2692 (N_2692,N_1391,N_1297);
and U2693 (N_2693,N_1860,N_1394);
nand U2694 (N_2694,N_1499,N_1359);
nand U2695 (N_2695,N_1021,N_1248);
or U2696 (N_2696,N_1579,N_1822);
xnor U2697 (N_2697,N_1901,N_1279);
or U2698 (N_2698,N_1573,N_1589);
nor U2699 (N_2699,N_1040,N_1286);
nand U2700 (N_2700,N_1126,N_1879);
nor U2701 (N_2701,N_1023,N_1322);
nor U2702 (N_2702,N_1090,N_1959);
or U2703 (N_2703,N_1821,N_1294);
and U2704 (N_2704,N_1791,N_1612);
and U2705 (N_2705,N_1387,N_1976);
nand U2706 (N_2706,N_1144,N_1746);
nor U2707 (N_2707,N_1252,N_1367);
and U2708 (N_2708,N_1017,N_1432);
or U2709 (N_2709,N_1629,N_1327);
nor U2710 (N_2710,N_1180,N_1793);
and U2711 (N_2711,N_1610,N_1970);
and U2712 (N_2712,N_1063,N_1505);
or U2713 (N_2713,N_1724,N_1816);
nor U2714 (N_2714,N_1078,N_1185);
and U2715 (N_2715,N_1931,N_1136);
nor U2716 (N_2716,N_1680,N_1701);
nand U2717 (N_2717,N_1212,N_1664);
nand U2718 (N_2718,N_1542,N_1843);
nand U2719 (N_2719,N_1433,N_1324);
and U2720 (N_2720,N_1773,N_1009);
nand U2721 (N_2721,N_1617,N_1803);
nor U2722 (N_2722,N_1849,N_1461);
and U2723 (N_2723,N_1891,N_1619);
nor U2724 (N_2724,N_1524,N_1333);
or U2725 (N_2725,N_1694,N_1568);
or U2726 (N_2726,N_1510,N_1950);
or U2727 (N_2727,N_1171,N_1602);
and U2728 (N_2728,N_1231,N_1749);
nand U2729 (N_2729,N_1227,N_1092);
or U2730 (N_2730,N_1852,N_1876);
and U2731 (N_2731,N_1975,N_1237);
or U2732 (N_2732,N_1592,N_1110);
nand U2733 (N_2733,N_1287,N_1450);
or U2734 (N_2734,N_1711,N_1997);
nor U2735 (N_2735,N_1677,N_1474);
or U2736 (N_2736,N_1222,N_1230);
and U2737 (N_2737,N_1243,N_1463);
nand U2738 (N_2738,N_1091,N_1718);
and U2739 (N_2739,N_1490,N_1163);
nor U2740 (N_2740,N_1184,N_1233);
nor U2741 (N_2741,N_1462,N_1036);
nor U2742 (N_2742,N_1979,N_1786);
or U2743 (N_2743,N_1913,N_1858);
and U2744 (N_2744,N_1047,N_1911);
nand U2745 (N_2745,N_1824,N_1418);
nor U2746 (N_2746,N_1062,N_1357);
and U2747 (N_2747,N_1518,N_1170);
or U2748 (N_2748,N_1314,N_1432);
and U2749 (N_2749,N_1856,N_1751);
xor U2750 (N_2750,N_1497,N_1435);
and U2751 (N_2751,N_1328,N_1912);
xor U2752 (N_2752,N_1075,N_1444);
xor U2753 (N_2753,N_1189,N_1608);
nand U2754 (N_2754,N_1797,N_1700);
nand U2755 (N_2755,N_1786,N_1233);
or U2756 (N_2756,N_1300,N_1442);
nor U2757 (N_2757,N_1068,N_1664);
nand U2758 (N_2758,N_1518,N_1282);
nor U2759 (N_2759,N_1317,N_1623);
nor U2760 (N_2760,N_1026,N_1156);
nor U2761 (N_2761,N_1529,N_1915);
or U2762 (N_2762,N_1278,N_1776);
nand U2763 (N_2763,N_1043,N_1339);
nor U2764 (N_2764,N_1227,N_1370);
and U2765 (N_2765,N_1840,N_1492);
or U2766 (N_2766,N_1505,N_1631);
and U2767 (N_2767,N_1947,N_1898);
nor U2768 (N_2768,N_1410,N_1687);
nor U2769 (N_2769,N_1457,N_1975);
nor U2770 (N_2770,N_1399,N_1789);
and U2771 (N_2771,N_1603,N_1392);
and U2772 (N_2772,N_1064,N_1891);
and U2773 (N_2773,N_1849,N_1379);
nand U2774 (N_2774,N_1987,N_1564);
or U2775 (N_2775,N_1151,N_1204);
or U2776 (N_2776,N_1880,N_1433);
or U2777 (N_2777,N_1967,N_1672);
nand U2778 (N_2778,N_1981,N_1646);
nand U2779 (N_2779,N_1705,N_1405);
and U2780 (N_2780,N_1148,N_1623);
or U2781 (N_2781,N_1291,N_1079);
nor U2782 (N_2782,N_1685,N_1875);
and U2783 (N_2783,N_1933,N_1562);
or U2784 (N_2784,N_1059,N_1898);
or U2785 (N_2785,N_1559,N_1672);
and U2786 (N_2786,N_1864,N_1910);
nand U2787 (N_2787,N_1679,N_1307);
or U2788 (N_2788,N_1625,N_1922);
nor U2789 (N_2789,N_1713,N_1916);
or U2790 (N_2790,N_1554,N_1156);
or U2791 (N_2791,N_1626,N_1275);
nor U2792 (N_2792,N_1336,N_1320);
and U2793 (N_2793,N_1781,N_1830);
or U2794 (N_2794,N_1923,N_1278);
nor U2795 (N_2795,N_1686,N_1683);
nand U2796 (N_2796,N_1030,N_1731);
and U2797 (N_2797,N_1375,N_1054);
or U2798 (N_2798,N_1899,N_1407);
and U2799 (N_2799,N_1753,N_1277);
or U2800 (N_2800,N_1070,N_1961);
and U2801 (N_2801,N_1956,N_1944);
and U2802 (N_2802,N_1118,N_1218);
nor U2803 (N_2803,N_1787,N_1392);
nand U2804 (N_2804,N_1730,N_1565);
or U2805 (N_2805,N_1595,N_1791);
nor U2806 (N_2806,N_1563,N_1247);
nor U2807 (N_2807,N_1703,N_1330);
nor U2808 (N_2808,N_1190,N_1512);
nand U2809 (N_2809,N_1637,N_1080);
nand U2810 (N_2810,N_1243,N_1080);
or U2811 (N_2811,N_1635,N_1251);
or U2812 (N_2812,N_1312,N_1379);
and U2813 (N_2813,N_1180,N_1591);
nand U2814 (N_2814,N_1038,N_1571);
and U2815 (N_2815,N_1420,N_1450);
nor U2816 (N_2816,N_1432,N_1316);
nor U2817 (N_2817,N_1890,N_1326);
nand U2818 (N_2818,N_1678,N_1966);
nor U2819 (N_2819,N_1134,N_1846);
nor U2820 (N_2820,N_1329,N_1698);
and U2821 (N_2821,N_1617,N_1964);
or U2822 (N_2822,N_1645,N_1693);
nand U2823 (N_2823,N_1942,N_1743);
or U2824 (N_2824,N_1608,N_1103);
and U2825 (N_2825,N_1376,N_1775);
and U2826 (N_2826,N_1106,N_1334);
and U2827 (N_2827,N_1202,N_1816);
nand U2828 (N_2828,N_1502,N_1281);
nand U2829 (N_2829,N_1609,N_1209);
nor U2830 (N_2830,N_1352,N_1322);
and U2831 (N_2831,N_1193,N_1828);
nand U2832 (N_2832,N_1845,N_1900);
nand U2833 (N_2833,N_1342,N_1097);
nor U2834 (N_2834,N_1730,N_1327);
and U2835 (N_2835,N_1882,N_1329);
nand U2836 (N_2836,N_1696,N_1885);
and U2837 (N_2837,N_1412,N_1410);
nor U2838 (N_2838,N_1156,N_1262);
or U2839 (N_2839,N_1924,N_1070);
and U2840 (N_2840,N_1219,N_1562);
nor U2841 (N_2841,N_1652,N_1574);
nor U2842 (N_2842,N_1754,N_1090);
nor U2843 (N_2843,N_1052,N_1548);
nand U2844 (N_2844,N_1772,N_1603);
nor U2845 (N_2845,N_1220,N_1979);
or U2846 (N_2846,N_1914,N_1832);
and U2847 (N_2847,N_1615,N_1666);
and U2848 (N_2848,N_1998,N_1789);
nor U2849 (N_2849,N_1883,N_1809);
nand U2850 (N_2850,N_1485,N_1478);
nand U2851 (N_2851,N_1236,N_1891);
nor U2852 (N_2852,N_1424,N_1574);
nand U2853 (N_2853,N_1007,N_1449);
nor U2854 (N_2854,N_1990,N_1386);
or U2855 (N_2855,N_1476,N_1063);
nor U2856 (N_2856,N_1465,N_1430);
and U2857 (N_2857,N_1216,N_1758);
and U2858 (N_2858,N_1748,N_1264);
or U2859 (N_2859,N_1177,N_1467);
or U2860 (N_2860,N_1900,N_1099);
or U2861 (N_2861,N_1630,N_1858);
and U2862 (N_2862,N_1398,N_1414);
or U2863 (N_2863,N_1338,N_1351);
nand U2864 (N_2864,N_1665,N_1319);
and U2865 (N_2865,N_1004,N_1928);
and U2866 (N_2866,N_1633,N_1113);
nand U2867 (N_2867,N_1046,N_1010);
and U2868 (N_2868,N_1038,N_1584);
nor U2869 (N_2869,N_1112,N_1006);
or U2870 (N_2870,N_1027,N_1026);
nor U2871 (N_2871,N_1611,N_1125);
nor U2872 (N_2872,N_1755,N_1984);
nand U2873 (N_2873,N_1887,N_1282);
or U2874 (N_2874,N_1610,N_1616);
and U2875 (N_2875,N_1837,N_1552);
or U2876 (N_2876,N_1359,N_1296);
nor U2877 (N_2877,N_1195,N_1942);
and U2878 (N_2878,N_1815,N_1273);
and U2879 (N_2879,N_1425,N_1938);
or U2880 (N_2880,N_1448,N_1205);
and U2881 (N_2881,N_1095,N_1786);
nand U2882 (N_2882,N_1269,N_1539);
nor U2883 (N_2883,N_1005,N_1739);
and U2884 (N_2884,N_1086,N_1193);
nand U2885 (N_2885,N_1717,N_1171);
nand U2886 (N_2886,N_1454,N_1782);
nor U2887 (N_2887,N_1084,N_1706);
and U2888 (N_2888,N_1031,N_1312);
xnor U2889 (N_2889,N_1992,N_1693);
xor U2890 (N_2890,N_1363,N_1219);
or U2891 (N_2891,N_1869,N_1956);
xnor U2892 (N_2892,N_1030,N_1813);
and U2893 (N_2893,N_1842,N_1824);
or U2894 (N_2894,N_1845,N_1338);
or U2895 (N_2895,N_1086,N_1641);
nand U2896 (N_2896,N_1365,N_1201);
nor U2897 (N_2897,N_1040,N_1067);
nand U2898 (N_2898,N_1313,N_1736);
or U2899 (N_2899,N_1233,N_1414);
nand U2900 (N_2900,N_1410,N_1167);
nand U2901 (N_2901,N_1142,N_1161);
and U2902 (N_2902,N_1626,N_1418);
nor U2903 (N_2903,N_1233,N_1643);
and U2904 (N_2904,N_1934,N_1401);
nor U2905 (N_2905,N_1073,N_1634);
and U2906 (N_2906,N_1805,N_1661);
nand U2907 (N_2907,N_1863,N_1965);
or U2908 (N_2908,N_1391,N_1144);
and U2909 (N_2909,N_1093,N_1527);
nor U2910 (N_2910,N_1523,N_1268);
nand U2911 (N_2911,N_1901,N_1937);
and U2912 (N_2912,N_1722,N_1640);
or U2913 (N_2913,N_1176,N_1344);
nand U2914 (N_2914,N_1115,N_1358);
or U2915 (N_2915,N_1694,N_1935);
nand U2916 (N_2916,N_1319,N_1799);
nand U2917 (N_2917,N_1488,N_1178);
and U2918 (N_2918,N_1406,N_1384);
and U2919 (N_2919,N_1883,N_1632);
nand U2920 (N_2920,N_1671,N_1399);
and U2921 (N_2921,N_1738,N_1289);
nor U2922 (N_2922,N_1779,N_1158);
nand U2923 (N_2923,N_1120,N_1318);
or U2924 (N_2924,N_1097,N_1966);
or U2925 (N_2925,N_1328,N_1362);
and U2926 (N_2926,N_1523,N_1907);
nand U2927 (N_2927,N_1436,N_1133);
nor U2928 (N_2928,N_1838,N_1710);
and U2929 (N_2929,N_1815,N_1779);
and U2930 (N_2930,N_1094,N_1547);
nor U2931 (N_2931,N_1411,N_1689);
nor U2932 (N_2932,N_1829,N_1149);
or U2933 (N_2933,N_1719,N_1533);
nand U2934 (N_2934,N_1966,N_1100);
nor U2935 (N_2935,N_1700,N_1025);
nor U2936 (N_2936,N_1737,N_1859);
or U2937 (N_2937,N_1636,N_1939);
and U2938 (N_2938,N_1108,N_1677);
nor U2939 (N_2939,N_1166,N_1861);
and U2940 (N_2940,N_1448,N_1909);
and U2941 (N_2941,N_1596,N_1740);
xnor U2942 (N_2942,N_1852,N_1269);
nand U2943 (N_2943,N_1752,N_1018);
and U2944 (N_2944,N_1430,N_1012);
and U2945 (N_2945,N_1477,N_1291);
or U2946 (N_2946,N_1779,N_1978);
nor U2947 (N_2947,N_1135,N_1243);
and U2948 (N_2948,N_1740,N_1524);
xnor U2949 (N_2949,N_1564,N_1595);
and U2950 (N_2950,N_1778,N_1504);
and U2951 (N_2951,N_1719,N_1188);
and U2952 (N_2952,N_1659,N_1976);
or U2953 (N_2953,N_1755,N_1254);
nor U2954 (N_2954,N_1259,N_1629);
and U2955 (N_2955,N_1750,N_1113);
nor U2956 (N_2956,N_1526,N_1387);
nor U2957 (N_2957,N_1043,N_1602);
or U2958 (N_2958,N_1203,N_1247);
or U2959 (N_2959,N_1099,N_1067);
or U2960 (N_2960,N_1653,N_1582);
and U2961 (N_2961,N_1071,N_1419);
and U2962 (N_2962,N_1733,N_1658);
nand U2963 (N_2963,N_1046,N_1002);
nor U2964 (N_2964,N_1705,N_1850);
and U2965 (N_2965,N_1751,N_1823);
or U2966 (N_2966,N_1088,N_1664);
or U2967 (N_2967,N_1903,N_1156);
and U2968 (N_2968,N_1411,N_1087);
and U2969 (N_2969,N_1048,N_1966);
nor U2970 (N_2970,N_1309,N_1411);
or U2971 (N_2971,N_1380,N_1134);
nor U2972 (N_2972,N_1504,N_1805);
or U2973 (N_2973,N_1695,N_1660);
and U2974 (N_2974,N_1058,N_1129);
or U2975 (N_2975,N_1475,N_1007);
nor U2976 (N_2976,N_1282,N_1828);
and U2977 (N_2977,N_1061,N_1661);
nand U2978 (N_2978,N_1124,N_1147);
nor U2979 (N_2979,N_1532,N_1421);
nor U2980 (N_2980,N_1024,N_1789);
or U2981 (N_2981,N_1816,N_1272);
nor U2982 (N_2982,N_1055,N_1335);
nand U2983 (N_2983,N_1397,N_1636);
and U2984 (N_2984,N_1519,N_1818);
nor U2985 (N_2985,N_1178,N_1190);
nor U2986 (N_2986,N_1275,N_1910);
and U2987 (N_2987,N_1215,N_1471);
and U2988 (N_2988,N_1010,N_1915);
or U2989 (N_2989,N_1383,N_1854);
xnor U2990 (N_2990,N_1335,N_1326);
and U2991 (N_2991,N_1802,N_1875);
and U2992 (N_2992,N_1193,N_1416);
xor U2993 (N_2993,N_1183,N_1893);
nand U2994 (N_2994,N_1930,N_1749);
nand U2995 (N_2995,N_1911,N_1726);
nand U2996 (N_2996,N_1949,N_1127);
and U2997 (N_2997,N_1098,N_1767);
nor U2998 (N_2998,N_1361,N_1472);
and U2999 (N_2999,N_1755,N_1060);
xnor U3000 (N_3000,N_2103,N_2607);
or U3001 (N_3001,N_2734,N_2049);
nor U3002 (N_3002,N_2909,N_2838);
or U3003 (N_3003,N_2966,N_2153);
nor U3004 (N_3004,N_2030,N_2656);
nand U3005 (N_3005,N_2148,N_2368);
or U3006 (N_3006,N_2835,N_2256);
and U3007 (N_3007,N_2226,N_2700);
and U3008 (N_3008,N_2866,N_2144);
nor U3009 (N_3009,N_2090,N_2419);
or U3010 (N_3010,N_2619,N_2766);
and U3011 (N_3011,N_2324,N_2091);
nor U3012 (N_3012,N_2793,N_2377);
nand U3013 (N_3013,N_2764,N_2265);
xor U3014 (N_3014,N_2503,N_2666);
or U3015 (N_3015,N_2326,N_2232);
or U3016 (N_3016,N_2356,N_2597);
and U3017 (N_3017,N_2385,N_2338);
nor U3018 (N_3018,N_2916,N_2970);
nor U3019 (N_3019,N_2512,N_2874);
nor U3020 (N_3020,N_2689,N_2977);
nor U3021 (N_3021,N_2576,N_2114);
nand U3022 (N_3022,N_2271,N_2981);
or U3023 (N_3023,N_2476,N_2540);
nand U3024 (N_3024,N_2509,N_2831);
nand U3025 (N_3025,N_2146,N_2985);
and U3026 (N_3026,N_2520,N_2038);
nand U3027 (N_3027,N_2094,N_2541);
and U3028 (N_3028,N_2648,N_2051);
nand U3029 (N_3029,N_2382,N_2446);
or U3030 (N_3030,N_2312,N_2273);
nand U3031 (N_3031,N_2078,N_2341);
and U3032 (N_3032,N_2658,N_2486);
and U3033 (N_3033,N_2829,N_2089);
or U3034 (N_3034,N_2622,N_2842);
or U3035 (N_3035,N_2505,N_2818);
nand U3036 (N_3036,N_2754,N_2650);
nand U3037 (N_3037,N_2283,N_2757);
or U3038 (N_3038,N_2009,N_2404);
nor U3039 (N_3039,N_2388,N_2363);
nor U3040 (N_3040,N_2275,N_2287);
or U3041 (N_3041,N_2302,N_2834);
or U3042 (N_3042,N_2875,N_2591);
nand U3043 (N_3043,N_2187,N_2889);
nand U3044 (N_3044,N_2353,N_2612);
and U3045 (N_3045,N_2483,N_2696);
nand U3046 (N_3046,N_2641,N_2344);
or U3047 (N_3047,N_2037,N_2109);
or U3048 (N_3048,N_2647,N_2913);
nor U3049 (N_3049,N_2034,N_2726);
nand U3050 (N_3050,N_2182,N_2280);
nand U3051 (N_3051,N_2203,N_2274);
and U3052 (N_3052,N_2065,N_2295);
and U3053 (N_3053,N_2452,N_2570);
nand U3054 (N_3054,N_2224,N_2730);
or U3055 (N_3055,N_2905,N_2460);
nor U3056 (N_3056,N_2347,N_2426);
nand U3057 (N_3057,N_2887,N_2635);
nand U3058 (N_3058,N_2473,N_2801);
nor U3059 (N_3059,N_2120,N_2911);
nor U3060 (N_3060,N_2624,N_2096);
nand U3061 (N_3061,N_2351,N_2539);
and U3062 (N_3062,N_2674,N_2490);
nand U3063 (N_3063,N_2603,N_2327);
or U3064 (N_3064,N_2346,N_2147);
and U3065 (N_3065,N_2467,N_2405);
or U3066 (N_3066,N_2093,N_2627);
and U3067 (N_3067,N_2787,N_2514);
or U3068 (N_3068,N_2593,N_2684);
or U3069 (N_3069,N_2851,N_2279);
nand U3070 (N_3070,N_2814,N_2912);
and U3071 (N_3071,N_2738,N_2447);
nor U3072 (N_3072,N_2343,N_2507);
nor U3073 (N_3073,N_2334,N_2546);
or U3074 (N_3074,N_2417,N_2588);
nor U3075 (N_3075,N_2972,N_2104);
or U3076 (N_3076,N_2762,N_2340);
xor U3077 (N_3077,N_2599,N_2944);
nand U3078 (N_3078,N_2322,N_2310);
or U3079 (N_3079,N_2974,N_2886);
or U3080 (N_3080,N_2501,N_2435);
nand U3081 (N_3081,N_2806,N_2075);
or U3082 (N_3082,N_2841,N_2748);
nand U3083 (N_3083,N_2703,N_2823);
and U3084 (N_3084,N_2554,N_2995);
and U3085 (N_3085,N_2837,N_2113);
xor U3086 (N_3086,N_2769,N_2087);
nand U3087 (N_3087,N_2918,N_2025);
and U3088 (N_3088,N_2016,N_2844);
and U3089 (N_3089,N_2252,N_2739);
and U3090 (N_3090,N_2943,N_2240);
nand U3091 (N_3091,N_2391,N_2527);
nor U3092 (N_3092,N_2167,N_2931);
nand U3093 (N_3093,N_2686,N_2048);
nand U3094 (N_3094,N_2522,N_2142);
and U3095 (N_3095,N_2006,N_2197);
or U3096 (N_3096,N_2425,N_2745);
nand U3097 (N_3097,N_2044,N_2538);
and U3098 (N_3098,N_2796,N_2238);
nor U3099 (N_3099,N_2967,N_2053);
or U3100 (N_3100,N_2156,N_2415);
nor U3101 (N_3101,N_2784,N_2459);
nor U3102 (N_3102,N_2297,N_2794);
nor U3103 (N_3103,N_2457,N_2646);
nand U3104 (N_3104,N_2106,N_2750);
nand U3105 (N_3105,N_2410,N_2565);
nor U3106 (N_3106,N_2481,N_2077);
nand U3107 (N_3107,N_2448,N_2953);
and U3108 (N_3108,N_2139,N_2836);
nor U3109 (N_3109,N_2433,N_2100);
nor U3110 (N_3110,N_2468,N_2592);
and U3111 (N_3111,N_2561,N_2384);
or U3112 (N_3112,N_2744,N_2278);
nand U3113 (N_3113,N_2598,N_2121);
or U3114 (N_3114,N_2880,N_2062);
and U3115 (N_3115,N_2581,N_2615);
xor U3116 (N_3116,N_2804,N_2097);
or U3117 (N_3117,N_2403,N_2978);
or U3118 (N_3118,N_2208,N_2492);
or U3119 (N_3119,N_2186,N_2019);
nand U3120 (N_3120,N_2463,N_2129);
or U3121 (N_3121,N_2408,N_2021);
nand U3122 (N_3122,N_2680,N_2763);
or U3123 (N_3123,N_2337,N_2239);
nand U3124 (N_3124,N_2637,N_2999);
nor U3125 (N_3125,N_2939,N_2811);
and U3126 (N_3126,N_2920,N_2262);
nand U3127 (N_3127,N_2218,N_2737);
or U3128 (N_3128,N_2946,N_2493);
or U3129 (N_3129,N_2079,N_2979);
or U3130 (N_3130,N_2155,N_2535);
or U3131 (N_3131,N_2907,N_2852);
nor U3132 (N_3132,N_2994,N_2000);
and U3133 (N_3133,N_2269,N_2487);
or U3134 (N_3134,N_2454,N_2498);
nand U3135 (N_3135,N_2050,N_2679);
nor U3136 (N_3136,N_2128,N_2135);
and U3137 (N_3137,N_2123,N_2160);
or U3138 (N_3138,N_2869,N_2475);
and U3139 (N_3139,N_2589,N_2349);
nor U3140 (N_3140,N_2854,N_2042);
and U3141 (N_3141,N_2372,N_2817);
or U3142 (N_3142,N_2098,N_2013);
or U3143 (N_3143,N_2193,N_2028);
and U3144 (N_3144,N_2675,N_2747);
nor U3145 (N_3145,N_2345,N_2017);
or U3146 (N_3146,N_2162,N_2761);
and U3147 (N_3147,N_2253,N_2717);
and U3148 (N_3148,N_2740,N_2845);
nor U3149 (N_3149,N_2657,N_2178);
and U3150 (N_3150,N_2753,N_2248);
nor U3151 (N_3151,N_2168,N_2477);
nor U3152 (N_3152,N_2354,N_2800);
or U3153 (N_3153,N_2722,N_2716);
nor U3154 (N_3154,N_2428,N_2792);
nand U3155 (N_3155,N_2936,N_2685);
nand U3156 (N_3156,N_2848,N_2413);
nor U3157 (N_3157,N_2832,N_2101);
nand U3158 (N_3158,N_2430,N_2870);
and U3159 (N_3159,N_2318,N_2192);
nor U3160 (N_3160,N_2115,N_2315);
nor U3161 (N_3161,N_2640,N_2059);
nand U3162 (N_3162,N_2623,N_2865);
or U3163 (N_3163,N_2665,N_2298);
and U3164 (N_3164,N_2258,N_2267);
or U3165 (N_3165,N_2471,N_2213);
or U3166 (N_3166,N_2373,N_2032);
nor U3167 (N_3167,N_2742,N_2055);
nor U3168 (N_3168,N_2949,N_2449);
nand U3169 (N_3169,N_2583,N_2444);
or U3170 (N_3170,N_2102,N_2709);
nand U3171 (N_3171,N_2469,N_2900);
and U3172 (N_3172,N_2394,N_2626);
and U3173 (N_3173,N_2910,N_2940);
nand U3174 (N_3174,N_2361,N_2618);
nor U3175 (N_3175,N_2960,N_2462);
xnor U3176 (N_3176,N_2140,N_2383);
nand U3177 (N_3177,N_2521,N_2973);
or U3178 (N_3178,N_2234,N_2644);
nand U3179 (N_3179,N_2491,N_2270);
or U3180 (N_3180,N_2692,N_2350);
nor U3181 (N_3181,N_2791,N_2779);
and U3182 (N_3182,N_2152,N_2617);
nand U3183 (N_3183,N_2321,N_2932);
and U3184 (N_3184,N_2751,N_2195);
nor U3185 (N_3185,N_2012,N_2442);
and U3186 (N_3186,N_2878,N_2897);
and U3187 (N_3187,N_2003,N_2330);
nand U3188 (N_3188,N_2743,N_2529);
or U3189 (N_3189,N_2859,N_2688);
nor U3190 (N_3190,N_2694,N_2702);
nor U3191 (N_3191,N_2506,N_2690);
and U3192 (N_3192,N_2370,N_2500);
or U3193 (N_3193,N_2456,N_2798);
nor U3194 (N_3194,N_2277,N_2357);
and U3195 (N_3195,N_2759,N_2400);
nor U3196 (N_3196,N_2282,N_2241);
nor U3197 (N_3197,N_2873,N_2867);
nor U3198 (N_3198,N_2510,N_2579);
and U3199 (N_3199,N_2336,N_2227);
nand U3200 (N_3200,N_2707,N_2802);
nand U3201 (N_3201,N_2063,N_2407);
nand U3202 (N_3202,N_2333,N_2711);
and U3203 (N_3203,N_2633,N_2803);
and U3204 (N_3204,N_2921,N_2437);
and U3205 (N_3205,N_2249,N_2790);
and U3206 (N_3206,N_2497,N_2902);
or U3207 (N_3207,N_2668,N_2472);
or U3208 (N_3208,N_2553,N_2574);
or U3209 (N_3209,N_2645,N_2821);
xor U3210 (N_3210,N_2504,N_2934);
nand U3211 (N_3211,N_2933,N_2774);
and U3212 (N_3212,N_2209,N_2780);
nand U3213 (N_3213,N_2876,N_2560);
or U3214 (N_3214,N_2638,N_2888);
nand U3215 (N_3215,N_2221,N_2057);
or U3216 (N_3216,N_2184,N_2201);
and U3217 (N_3217,N_2673,N_2714);
and U3218 (N_3218,N_2247,N_2223);
nor U3219 (N_3219,N_2935,N_2547);
or U3220 (N_3220,N_2732,N_2534);
nand U3221 (N_3221,N_2022,N_2849);
and U3222 (N_3222,N_2060,N_2375);
and U3223 (N_3223,N_2728,N_2489);
or U3224 (N_3224,N_2568,N_2290);
nor U3225 (N_3225,N_2177,N_2171);
or U3226 (N_3226,N_2358,N_2996);
nor U3227 (N_3227,N_2020,N_2567);
nand U3228 (N_3228,N_2450,N_2133);
and U3229 (N_3229,N_2216,N_2975);
and U3230 (N_3230,N_2136,N_2231);
xnor U3231 (N_3231,N_2092,N_2004);
nand U3232 (N_3232,N_2421,N_2924);
nand U3233 (N_3233,N_2785,N_2422);
and U3234 (N_3234,N_2643,N_2533);
nand U3235 (N_3235,N_2432,N_2304);
or U3236 (N_3236,N_2608,N_2291);
or U3237 (N_3237,N_2537,N_2392);
or U3238 (N_3238,N_2519,N_2724);
and U3239 (N_3239,N_2395,N_2308);
nand U3240 (N_3240,N_2122,N_2040);
or U3241 (N_3241,N_2074,N_2157);
nand U3242 (N_3242,N_2894,N_2856);
or U3243 (N_3243,N_2896,N_2788);
or U3244 (N_3244,N_2323,N_2143);
nand U3245 (N_3245,N_2664,N_2190);
or U3246 (N_3246,N_2963,N_2479);
nor U3247 (N_3247,N_2993,N_2331);
and U3248 (N_3248,N_2551,N_2513);
nand U3249 (N_3249,N_2652,N_2495);
or U3250 (N_3250,N_2969,N_2332);
xnor U3251 (N_3251,N_2399,N_2884);
or U3252 (N_3252,N_2515,N_2531);
nor U3253 (N_3253,N_2199,N_2263);
and U3254 (N_3254,N_2923,N_2927);
nand U3255 (N_3255,N_2289,N_2789);
and U3256 (N_3256,N_2393,N_2169);
or U3257 (N_3257,N_2107,N_2095);
nand U3258 (N_3258,N_2015,N_2138);
nor U3259 (N_3259,N_2613,N_2161);
nor U3260 (N_3260,N_2134,N_2555);
and U3261 (N_3261,N_2071,N_2957);
nand U3262 (N_3262,N_2339,N_2301);
nor U3263 (N_3263,N_2914,N_2816);
nor U3264 (N_3264,N_2954,N_2145);
and U3265 (N_3265,N_2438,N_2670);
or U3266 (N_3266,N_2891,N_2198);
or U3267 (N_3267,N_2982,N_2655);
or U3268 (N_3268,N_2526,N_2584);
nor U3269 (N_3269,N_2217,N_2125);
and U3270 (N_3270,N_2200,N_2243);
xnor U3271 (N_3271,N_2137,N_2296);
nand U3272 (N_3272,N_2843,N_2215);
or U3273 (N_3273,N_2904,N_2118);
or U3274 (N_3274,N_2868,N_2132);
nor U3275 (N_3275,N_2369,N_2947);
nor U3276 (N_3276,N_2795,N_2528);
nor U3277 (N_3277,N_2154,N_2853);
and U3278 (N_3278,N_2445,N_2381);
and U3279 (N_3279,N_2600,N_2205);
nand U3280 (N_3280,N_2112,N_2434);
nand U3281 (N_3281,N_2485,N_2839);
or U3282 (N_3282,N_2536,N_2228);
or U3283 (N_3283,N_2611,N_2713);
xor U3284 (N_3284,N_2461,N_2586);
nor U3285 (N_3285,N_2299,N_2770);
xnor U3286 (N_3286,N_2928,N_2746);
nor U3287 (N_3287,N_2237,N_2799);
nand U3288 (N_3288,N_2698,N_2488);
or U3289 (N_3289,N_2731,N_2039);
or U3290 (N_3290,N_2986,N_2108);
or U3291 (N_3291,N_2950,N_2305);
nor U3292 (N_3292,N_2458,N_2628);
and U3293 (N_3293,N_2482,N_2056);
or U3294 (N_3294,N_2261,N_2701);
nand U3295 (N_3295,N_2041,N_2710);
and U3296 (N_3296,N_2244,N_2313);
or U3297 (N_3297,N_2725,N_2671);
and U3298 (N_3298,N_2348,N_2174);
nand U3299 (N_3299,N_2508,N_2777);
nor U3300 (N_3300,N_2235,N_2890);
xor U3301 (N_3301,N_2704,N_2119);
and U3302 (N_3302,N_2691,N_2066);
nand U3303 (N_3303,N_2782,N_2046);
or U3304 (N_3304,N_2523,N_2983);
nand U3305 (N_3305,N_2001,N_2951);
nand U3306 (N_3306,N_2266,N_2773);
and U3307 (N_3307,N_2809,N_2727);
nand U3308 (N_3308,N_2429,N_2797);
and U3309 (N_3309,N_2952,N_2516);
nor U3310 (N_3310,N_2320,N_2557);
or U3311 (N_3311,N_2176,N_2110);
nand U3312 (N_3312,N_2436,N_2260);
nor U3313 (N_3313,N_2511,N_2396);
nand U3314 (N_3314,N_2272,N_2465);
nand U3315 (N_3315,N_2807,N_2319);
or U3316 (N_3316,N_2002,N_2903);
nor U3317 (N_3317,N_2958,N_2230);
nand U3318 (N_3318,N_2259,N_2687);
or U3319 (N_3319,N_2948,N_2307);
nand U3320 (N_3320,N_2602,N_2478);
and U3321 (N_3321,N_2359,N_2676);
nand U3322 (N_3322,N_2172,N_2822);
and U3323 (N_3323,N_2376,N_2860);
or U3324 (N_3324,N_2300,N_2833);
nand U3325 (N_3325,N_2654,N_2810);
nand U3326 (N_3326,N_2882,N_2517);
and U3327 (N_3327,N_2758,N_2412);
and U3328 (N_3328,N_2556,N_2081);
nand U3329 (N_3329,N_2086,N_2961);
or U3330 (N_3330,N_2634,N_2767);
nor U3331 (N_3331,N_2827,N_2008);
or U3332 (N_3332,N_2585,N_2830);
nand U3333 (N_3333,N_2639,N_2968);
or U3334 (N_3334,N_2058,N_2861);
and U3335 (N_3335,N_2054,N_2678);
or U3336 (N_3336,N_2552,N_2151);
and U3337 (N_3337,N_2276,N_2938);
or U3338 (N_3338,N_2605,N_2219);
nand U3339 (N_3339,N_2206,N_2695);
nor U3340 (N_3340,N_2989,N_2772);
or U3341 (N_3341,N_2294,N_2677);
nand U3342 (N_3342,N_2942,N_2862);
nor U3343 (N_3343,N_2202,N_2250);
nor U3344 (N_3344,N_2316,N_2825);
nor U3345 (N_3345,N_2893,N_2594);
and U3346 (N_3346,N_2877,N_2719);
or U3347 (N_3347,N_2033,N_2416);
nor U3348 (N_3348,N_2311,N_2755);
and U3349 (N_3349,N_2466,N_2706);
and U3350 (N_3350,N_2741,N_2616);
nor U3351 (N_3351,N_2669,N_2998);
or U3352 (N_3352,N_2418,N_2901);
and U3353 (N_3353,N_2693,N_2898);
nand U3354 (N_3354,N_2127,N_2211);
nor U3355 (N_3355,N_2614,N_2518);
nand U3356 (N_3356,N_2378,N_2858);
or U3357 (N_3357,N_2715,N_2024);
nand U3358 (N_3358,N_2220,N_2783);
and U3359 (N_3359,N_2464,N_2281);
or U3360 (N_3360,N_2962,N_2812);
nand U3361 (N_3361,N_2293,N_2064);
and U3362 (N_3362,N_2029,N_2188);
and U3363 (N_3363,N_2007,N_2180);
nor U3364 (N_3364,N_2937,N_2011);
nor U3365 (N_3365,N_2035,N_2246);
nand U3366 (N_3366,N_2661,N_2288);
or U3367 (N_3367,N_2440,N_2204);
nand U3368 (N_3368,N_2660,N_2729);
nand U3369 (N_3369,N_2264,N_2683);
nand U3370 (N_3370,N_2328,N_2760);
xor U3371 (N_3371,N_2663,N_2047);
or U3372 (N_3372,N_2023,N_2045);
nand U3373 (N_3373,N_2181,N_2229);
nor U3374 (N_3374,N_2105,N_2752);
nor U3375 (N_3375,N_2212,N_2362);
or U3376 (N_3376,N_2257,N_2544);
and U3377 (N_3377,N_2596,N_2031);
or U3378 (N_3378,N_2329,N_2871);
or U3379 (N_3379,N_2131,N_2292);
and U3380 (N_3380,N_2926,N_2580);
and U3381 (N_3381,N_2820,N_2380);
nor U3382 (N_3382,N_2563,N_2242);
and U3383 (N_3383,N_2411,N_2636);
nor U3384 (N_3384,N_2254,N_2718);
or U3385 (N_3385,N_2183,N_2451);
and U3386 (N_3386,N_2899,N_2582);
nand U3387 (N_3387,N_2915,N_2965);
and U3388 (N_3388,N_2813,N_2499);
xnor U3389 (N_3389,N_2595,N_2141);
or U3390 (N_3390,N_2335,N_2632);
nand U3391 (N_3391,N_2987,N_2117);
and U3392 (N_3392,N_2964,N_2991);
nand U3393 (N_3393,N_2808,N_2578);
and U3394 (N_3394,N_2524,N_2149);
nor U3395 (N_3395,N_2420,N_2620);
or U3396 (N_3396,N_2771,N_2409);
nand U3397 (N_3397,N_2530,N_2721);
or U3398 (N_3398,N_2572,N_2325);
and U3399 (N_3399,N_2708,N_2571);
or U3400 (N_3400,N_2443,N_2945);
nor U3401 (N_3401,N_2371,N_2662);
xnor U3402 (N_3402,N_2532,N_2883);
nor U3403 (N_3403,N_2562,N_2398);
and U3404 (N_3404,N_2885,N_2955);
and U3405 (N_3405,N_2525,N_2667);
nand U3406 (N_3406,N_2749,N_2917);
nand U3407 (N_3407,N_2401,N_2303);
nand U3408 (N_3408,N_2659,N_2036);
nand U3409 (N_3409,N_2052,N_2824);
xor U3410 (N_3410,N_2402,N_2360);
nor U3411 (N_3411,N_2158,N_2681);
or U3412 (N_3412,N_2815,N_2175);
and U3413 (N_3413,N_2439,N_2159);
or U3414 (N_3414,N_2018,N_2210);
or U3415 (N_3415,N_2756,N_2621);
nand U3416 (N_3416,N_2855,N_2251);
and U3417 (N_3417,N_2406,N_2379);
or U3418 (N_3418,N_2355,N_2268);
and U3419 (N_3419,N_2245,N_2083);
nand U3420 (N_3420,N_2971,N_2712);
nor U3421 (N_3421,N_2941,N_2697);
nor U3422 (N_3422,N_2390,N_2863);
nand U3423 (N_3423,N_2082,N_2455);
and U3424 (N_3424,N_2374,N_2805);
or U3425 (N_3425,N_2189,N_2786);
or U3426 (N_3426,N_2781,N_2850);
nand U3427 (N_3427,N_2630,N_2566);
and U3428 (N_3428,N_2494,N_2352);
or U3429 (N_3429,N_2366,N_2179);
nand U3430 (N_3430,N_2069,N_2705);
nor U3431 (N_3431,N_2919,N_2061);
or U3432 (N_3432,N_2881,N_2984);
or U3433 (N_3433,N_2496,N_2389);
nor U3434 (N_3434,N_2606,N_2587);
and U3435 (N_3435,N_2906,N_2550);
nor U3436 (N_3436,N_2545,N_2959);
nor U3437 (N_3437,N_2930,N_2474);
xnor U3438 (N_3438,N_2424,N_2126);
nand U3439 (N_3439,N_2191,N_2609);
or U3440 (N_3440,N_2828,N_2990);
nand U3441 (N_3441,N_2768,N_2651);
nand U3442 (N_3442,N_2733,N_2776);
nor U3443 (N_3443,N_2342,N_2601);
nand U3444 (N_3444,N_2558,N_2765);
nand U3445 (N_3445,N_2085,N_2173);
and U3446 (N_3446,N_2625,N_2367);
nor U3447 (N_3447,N_2778,N_2222);
or U3448 (N_3448,N_2604,N_2387);
and U3449 (N_3449,N_2872,N_2014);
nand U3450 (N_3450,N_2699,N_2847);
or U3451 (N_3451,N_2099,N_2925);
or U3452 (N_3452,N_2010,N_2427);
nand U3453 (N_3453,N_2116,N_2286);
nand U3454 (N_3454,N_2736,N_2164);
nor U3455 (N_3455,N_2543,N_2577);
and U3456 (N_3456,N_2067,N_2559);
nand U3457 (N_3457,N_2185,N_2441);
nor U3458 (N_3458,N_2775,N_2629);
and U3459 (N_3459,N_2956,N_2480);
nor U3460 (N_3460,N_2988,N_2072);
or U3461 (N_3461,N_2027,N_2976);
or U3462 (N_3462,N_2233,N_2255);
nand U3463 (N_3463,N_2165,N_2214);
nand U3464 (N_3464,N_2364,N_2895);
nor U3465 (N_3465,N_2929,N_2317);
nor U3466 (N_3466,N_2470,N_2484);
and U3467 (N_3467,N_2682,N_2076);
nor U3468 (N_3468,N_2631,N_2084);
nand U3469 (N_3469,N_2194,N_2124);
nand U3470 (N_3470,N_2386,N_2992);
nand U3471 (N_3471,N_2314,N_2542);
or U3472 (N_3472,N_2573,N_2819);
and U3473 (N_3473,N_2908,N_2163);
nand U3474 (N_3474,N_2864,N_2225);
nor U3475 (N_3475,N_2569,N_2026);
or U3476 (N_3476,N_2564,N_2548);
nor U3477 (N_3477,N_2170,N_2735);
nand U3478 (N_3478,N_2166,N_2610);
nor U3479 (N_3479,N_2309,N_2840);
and U3480 (N_3480,N_2005,N_2892);
or U3481 (N_3481,N_2088,N_2073);
nand U3482 (N_3482,N_2590,N_2070);
and U3483 (N_3483,N_2653,N_2720);
or U3484 (N_3484,N_2080,N_2826);
or U3485 (N_3485,N_2453,N_2549);
or U3486 (N_3486,N_2846,N_2431);
nand U3487 (N_3487,N_2068,N_2980);
nand U3488 (N_3488,N_2642,N_2043);
nand U3489 (N_3489,N_2397,N_2236);
and U3490 (N_3490,N_2997,N_2723);
nor U3491 (N_3491,N_2130,N_2414);
nand U3492 (N_3492,N_2879,N_2111);
or U3493 (N_3493,N_2365,N_2284);
nand U3494 (N_3494,N_2285,N_2306);
xnor U3495 (N_3495,N_2423,N_2672);
nor U3496 (N_3496,N_2150,N_2196);
nor U3497 (N_3497,N_2922,N_2207);
nor U3498 (N_3498,N_2575,N_2502);
or U3499 (N_3499,N_2649,N_2857);
nor U3500 (N_3500,N_2678,N_2122);
and U3501 (N_3501,N_2648,N_2794);
nand U3502 (N_3502,N_2226,N_2443);
or U3503 (N_3503,N_2007,N_2281);
and U3504 (N_3504,N_2899,N_2865);
nand U3505 (N_3505,N_2091,N_2194);
or U3506 (N_3506,N_2887,N_2091);
nand U3507 (N_3507,N_2602,N_2512);
nand U3508 (N_3508,N_2424,N_2031);
nor U3509 (N_3509,N_2376,N_2980);
and U3510 (N_3510,N_2321,N_2492);
xor U3511 (N_3511,N_2130,N_2331);
or U3512 (N_3512,N_2438,N_2322);
and U3513 (N_3513,N_2735,N_2919);
nor U3514 (N_3514,N_2238,N_2386);
nand U3515 (N_3515,N_2826,N_2679);
and U3516 (N_3516,N_2083,N_2811);
or U3517 (N_3517,N_2712,N_2588);
or U3518 (N_3518,N_2888,N_2031);
nand U3519 (N_3519,N_2723,N_2114);
nand U3520 (N_3520,N_2658,N_2182);
or U3521 (N_3521,N_2367,N_2712);
nor U3522 (N_3522,N_2194,N_2924);
and U3523 (N_3523,N_2152,N_2996);
nand U3524 (N_3524,N_2645,N_2565);
or U3525 (N_3525,N_2963,N_2316);
nor U3526 (N_3526,N_2249,N_2714);
nor U3527 (N_3527,N_2545,N_2460);
nand U3528 (N_3528,N_2272,N_2928);
nor U3529 (N_3529,N_2848,N_2733);
nor U3530 (N_3530,N_2391,N_2440);
and U3531 (N_3531,N_2872,N_2576);
nand U3532 (N_3532,N_2348,N_2872);
or U3533 (N_3533,N_2134,N_2028);
or U3534 (N_3534,N_2637,N_2069);
or U3535 (N_3535,N_2339,N_2211);
and U3536 (N_3536,N_2695,N_2527);
xor U3537 (N_3537,N_2412,N_2439);
or U3538 (N_3538,N_2081,N_2894);
nor U3539 (N_3539,N_2219,N_2207);
or U3540 (N_3540,N_2374,N_2396);
and U3541 (N_3541,N_2055,N_2726);
and U3542 (N_3542,N_2413,N_2983);
and U3543 (N_3543,N_2708,N_2092);
nand U3544 (N_3544,N_2504,N_2640);
nand U3545 (N_3545,N_2545,N_2835);
or U3546 (N_3546,N_2722,N_2000);
and U3547 (N_3547,N_2452,N_2774);
nor U3548 (N_3548,N_2732,N_2106);
nor U3549 (N_3549,N_2130,N_2427);
nand U3550 (N_3550,N_2607,N_2757);
nor U3551 (N_3551,N_2992,N_2228);
nor U3552 (N_3552,N_2587,N_2171);
nand U3553 (N_3553,N_2569,N_2340);
nor U3554 (N_3554,N_2280,N_2392);
or U3555 (N_3555,N_2894,N_2779);
or U3556 (N_3556,N_2737,N_2732);
and U3557 (N_3557,N_2223,N_2124);
nor U3558 (N_3558,N_2935,N_2740);
or U3559 (N_3559,N_2635,N_2462);
or U3560 (N_3560,N_2704,N_2631);
nand U3561 (N_3561,N_2642,N_2474);
nor U3562 (N_3562,N_2907,N_2698);
nor U3563 (N_3563,N_2018,N_2711);
or U3564 (N_3564,N_2641,N_2631);
nor U3565 (N_3565,N_2067,N_2850);
or U3566 (N_3566,N_2477,N_2882);
and U3567 (N_3567,N_2834,N_2536);
or U3568 (N_3568,N_2444,N_2569);
nand U3569 (N_3569,N_2348,N_2715);
nor U3570 (N_3570,N_2143,N_2446);
nor U3571 (N_3571,N_2594,N_2920);
nor U3572 (N_3572,N_2955,N_2530);
nor U3573 (N_3573,N_2581,N_2113);
nor U3574 (N_3574,N_2626,N_2847);
or U3575 (N_3575,N_2490,N_2171);
and U3576 (N_3576,N_2427,N_2076);
nand U3577 (N_3577,N_2340,N_2852);
nor U3578 (N_3578,N_2740,N_2335);
nor U3579 (N_3579,N_2945,N_2184);
and U3580 (N_3580,N_2434,N_2582);
and U3581 (N_3581,N_2984,N_2983);
or U3582 (N_3582,N_2720,N_2476);
and U3583 (N_3583,N_2304,N_2069);
or U3584 (N_3584,N_2371,N_2915);
or U3585 (N_3585,N_2836,N_2970);
or U3586 (N_3586,N_2260,N_2592);
or U3587 (N_3587,N_2080,N_2655);
and U3588 (N_3588,N_2302,N_2886);
nor U3589 (N_3589,N_2737,N_2162);
or U3590 (N_3590,N_2988,N_2813);
and U3591 (N_3591,N_2252,N_2016);
nor U3592 (N_3592,N_2216,N_2836);
nand U3593 (N_3593,N_2670,N_2710);
nor U3594 (N_3594,N_2321,N_2313);
nor U3595 (N_3595,N_2867,N_2695);
or U3596 (N_3596,N_2766,N_2746);
or U3597 (N_3597,N_2822,N_2890);
or U3598 (N_3598,N_2213,N_2055);
or U3599 (N_3599,N_2076,N_2511);
or U3600 (N_3600,N_2611,N_2878);
or U3601 (N_3601,N_2591,N_2175);
or U3602 (N_3602,N_2411,N_2200);
nor U3603 (N_3603,N_2633,N_2360);
or U3604 (N_3604,N_2217,N_2739);
and U3605 (N_3605,N_2978,N_2639);
nand U3606 (N_3606,N_2096,N_2740);
nor U3607 (N_3607,N_2918,N_2229);
nor U3608 (N_3608,N_2734,N_2918);
or U3609 (N_3609,N_2295,N_2020);
nor U3610 (N_3610,N_2605,N_2053);
nor U3611 (N_3611,N_2363,N_2062);
nand U3612 (N_3612,N_2697,N_2155);
nor U3613 (N_3613,N_2738,N_2157);
nand U3614 (N_3614,N_2924,N_2423);
or U3615 (N_3615,N_2671,N_2376);
or U3616 (N_3616,N_2298,N_2644);
or U3617 (N_3617,N_2344,N_2876);
nor U3618 (N_3618,N_2875,N_2367);
nor U3619 (N_3619,N_2381,N_2601);
nor U3620 (N_3620,N_2097,N_2660);
nand U3621 (N_3621,N_2039,N_2583);
or U3622 (N_3622,N_2895,N_2525);
nor U3623 (N_3623,N_2801,N_2746);
and U3624 (N_3624,N_2728,N_2095);
nor U3625 (N_3625,N_2605,N_2412);
nand U3626 (N_3626,N_2506,N_2598);
and U3627 (N_3627,N_2039,N_2304);
or U3628 (N_3628,N_2252,N_2426);
or U3629 (N_3629,N_2316,N_2336);
or U3630 (N_3630,N_2292,N_2708);
or U3631 (N_3631,N_2504,N_2952);
nand U3632 (N_3632,N_2384,N_2487);
nand U3633 (N_3633,N_2150,N_2665);
or U3634 (N_3634,N_2721,N_2367);
nor U3635 (N_3635,N_2235,N_2721);
nand U3636 (N_3636,N_2825,N_2225);
or U3637 (N_3637,N_2648,N_2946);
and U3638 (N_3638,N_2913,N_2180);
or U3639 (N_3639,N_2793,N_2897);
and U3640 (N_3640,N_2574,N_2512);
and U3641 (N_3641,N_2432,N_2958);
nor U3642 (N_3642,N_2511,N_2678);
or U3643 (N_3643,N_2694,N_2631);
and U3644 (N_3644,N_2881,N_2452);
and U3645 (N_3645,N_2992,N_2689);
and U3646 (N_3646,N_2031,N_2355);
and U3647 (N_3647,N_2374,N_2976);
or U3648 (N_3648,N_2323,N_2481);
and U3649 (N_3649,N_2757,N_2136);
and U3650 (N_3650,N_2983,N_2361);
nor U3651 (N_3651,N_2011,N_2770);
or U3652 (N_3652,N_2634,N_2159);
or U3653 (N_3653,N_2416,N_2709);
nand U3654 (N_3654,N_2393,N_2427);
and U3655 (N_3655,N_2923,N_2893);
nand U3656 (N_3656,N_2819,N_2860);
or U3657 (N_3657,N_2736,N_2632);
nand U3658 (N_3658,N_2568,N_2030);
or U3659 (N_3659,N_2665,N_2152);
and U3660 (N_3660,N_2426,N_2909);
or U3661 (N_3661,N_2666,N_2113);
nand U3662 (N_3662,N_2637,N_2293);
and U3663 (N_3663,N_2111,N_2569);
and U3664 (N_3664,N_2315,N_2098);
nor U3665 (N_3665,N_2574,N_2461);
nor U3666 (N_3666,N_2949,N_2086);
and U3667 (N_3667,N_2098,N_2437);
or U3668 (N_3668,N_2235,N_2599);
nor U3669 (N_3669,N_2127,N_2958);
nand U3670 (N_3670,N_2354,N_2143);
nand U3671 (N_3671,N_2785,N_2605);
and U3672 (N_3672,N_2988,N_2606);
nor U3673 (N_3673,N_2269,N_2237);
and U3674 (N_3674,N_2998,N_2886);
or U3675 (N_3675,N_2145,N_2110);
nor U3676 (N_3676,N_2737,N_2933);
nand U3677 (N_3677,N_2124,N_2013);
nor U3678 (N_3678,N_2010,N_2766);
nand U3679 (N_3679,N_2503,N_2192);
and U3680 (N_3680,N_2992,N_2192);
or U3681 (N_3681,N_2363,N_2621);
nor U3682 (N_3682,N_2324,N_2563);
and U3683 (N_3683,N_2225,N_2953);
and U3684 (N_3684,N_2196,N_2040);
or U3685 (N_3685,N_2831,N_2944);
nor U3686 (N_3686,N_2560,N_2710);
and U3687 (N_3687,N_2281,N_2535);
nand U3688 (N_3688,N_2203,N_2682);
nand U3689 (N_3689,N_2793,N_2331);
or U3690 (N_3690,N_2444,N_2727);
or U3691 (N_3691,N_2845,N_2270);
nand U3692 (N_3692,N_2404,N_2324);
and U3693 (N_3693,N_2800,N_2028);
nor U3694 (N_3694,N_2170,N_2703);
nand U3695 (N_3695,N_2682,N_2619);
nand U3696 (N_3696,N_2139,N_2783);
and U3697 (N_3697,N_2617,N_2879);
and U3698 (N_3698,N_2838,N_2327);
nand U3699 (N_3699,N_2184,N_2106);
nor U3700 (N_3700,N_2726,N_2701);
nor U3701 (N_3701,N_2194,N_2926);
nand U3702 (N_3702,N_2354,N_2099);
or U3703 (N_3703,N_2977,N_2560);
nand U3704 (N_3704,N_2788,N_2015);
nor U3705 (N_3705,N_2226,N_2678);
and U3706 (N_3706,N_2086,N_2396);
and U3707 (N_3707,N_2704,N_2791);
nand U3708 (N_3708,N_2419,N_2180);
nand U3709 (N_3709,N_2057,N_2102);
and U3710 (N_3710,N_2415,N_2416);
nor U3711 (N_3711,N_2742,N_2175);
nor U3712 (N_3712,N_2972,N_2468);
nor U3713 (N_3713,N_2983,N_2392);
xor U3714 (N_3714,N_2575,N_2258);
or U3715 (N_3715,N_2329,N_2155);
nand U3716 (N_3716,N_2030,N_2011);
nor U3717 (N_3717,N_2330,N_2595);
nand U3718 (N_3718,N_2534,N_2585);
xor U3719 (N_3719,N_2822,N_2404);
or U3720 (N_3720,N_2373,N_2797);
nor U3721 (N_3721,N_2392,N_2103);
nand U3722 (N_3722,N_2842,N_2097);
nor U3723 (N_3723,N_2576,N_2642);
xor U3724 (N_3724,N_2560,N_2913);
and U3725 (N_3725,N_2812,N_2116);
nor U3726 (N_3726,N_2298,N_2065);
or U3727 (N_3727,N_2944,N_2941);
and U3728 (N_3728,N_2767,N_2443);
nand U3729 (N_3729,N_2261,N_2270);
nand U3730 (N_3730,N_2859,N_2302);
nor U3731 (N_3731,N_2156,N_2809);
nand U3732 (N_3732,N_2995,N_2388);
or U3733 (N_3733,N_2896,N_2217);
and U3734 (N_3734,N_2585,N_2176);
nand U3735 (N_3735,N_2884,N_2204);
nand U3736 (N_3736,N_2646,N_2816);
and U3737 (N_3737,N_2324,N_2008);
nor U3738 (N_3738,N_2216,N_2424);
xnor U3739 (N_3739,N_2994,N_2599);
nor U3740 (N_3740,N_2071,N_2473);
and U3741 (N_3741,N_2933,N_2821);
and U3742 (N_3742,N_2552,N_2498);
and U3743 (N_3743,N_2895,N_2403);
nor U3744 (N_3744,N_2617,N_2085);
nor U3745 (N_3745,N_2676,N_2513);
nor U3746 (N_3746,N_2243,N_2127);
or U3747 (N_3747,N_2648,N_2247);
nand U3748 (N_3748,N_2333,N_2514);
and U3749 (N_3749,N_2646,N_2676);
or U3750 (N_3750,N_2726,N_2767);
and U3751 (N_3751,N_2659,N_2218);
or U3752 (N_3752,N_2411,N_2601);
or U3753 (N_3753,N_2807,N_2766);
nor U3754 (N_3754,N_2657,N_2600);
or U3755 (N_3755,N_2349,N_2182);
nor U3756 (N_3756,N_2739,N_2430);
nand U3757 (N_3757,N_2415,N_2140);
and U3758 (N_3758,N_2452,N_2870);
and U3759 (N_3759,N_2782,N_2650);
nand U3760 (N_3760,N_2418,N_2896);
or U3761 (N_3761,N_2485,N_2096);
nor U3762 (N_3762,N_2947,N_2917);
nor U3763 (N_3763,N_2553,N_2769);
nand U3764 (N_3764,N_2277,N_2665);
and U3765 (N_3765,N_2534,N_2524);
or U3766 (N_3766,N_2117,N_2975);
nor U3767 (N_3767,N_2554,N_2672);
nor U3768 (N_3768,N_2952,N_2532);
nor U3769 (N_3769,N_2033,N_2050);
nand U3770 (N_3770,N_2792,N_2692);
nor U3771 (N_3771,N_2104,N_2587);
nor U3772 (N_3772,N_2057,N_2444);
and U3773 (N_3773,N_2210,N_2860);
or U3774 (N_3774,N_2088,N_2242);
or U3775 (N_3775,N_2770,N_2021);
nor U3776 (N_3776,N_2590,N_2750);
nor U3777 (N_3777,N_2280,N_2984);
nand U3778 (N_3778,N_2667,N_2643);
or U3779 (N_3779,N_2463,N_2188);
nor U3780 (N_3780,N_2084,N_2342);
nor U3781 (N_3781,N_2542,N_2938);
or U3782 (N_3782,N_2205,N_2386);
nor U3783 (N_3783,N_2568,N_2100);
or U3784 (N_3784,N_2547,N_2422);
and U3785 (N_3785,N_2572,N_2385);
nor U3786 (N_3786,N_2199,N_2705);
nor U3787 (N_3787,N_2702,N_2655);
xnor U3788 (N_3788,N_2661,N_2546);
nor U3789 (N_3789,N_2331,N_2394);
xnor U3790 (N_3790,N_2825,N_2788);
or U3791 (N_3791,N_2589,N_2012);
or U3792 (N_3792,N_2795,N_2193);
or U3793 (N_3793,N_2917,N_2999);
nor U3794 (N_3794,N_2226,N_2077);
xor U3795 (N_3795,N_2214,N_2530);
and U3796 (N_3796,N_2239,N_2513);
nor U3797 (N_3797,N_2026,N_2379);
or U3798 (N_3798,N_2674,N_2407);
nand U3799 (N_3799,N_2647,N_2928);
and U3800 (N_3800,N_2825,N_2967);
nor U3801 (N_3801,N_2441,N_2765);
or U3802 (N_3802,N_2263,N_2817);
or U3803 (N_3803,N_2783,N_2104);
or U3804 (N_3804,N_2701,N_2807);
and U3805 (N_3805,N_2763,N_2882);
or U3806 (N_3806,N_2326,N_2400);
and U3807 (N_3807,N_2208,N_2875);
and U3808 (N_3808,N_2031,N_2279);
or U3809 (N_3809,N_2163,N_2823);
nand U3810 (N_3810,N_2145,N_2198);
and U3811 (N_3811,N_2813,N_2252);
or U3812 (N_3812,N_2379,N_2068);
nand U3813 (N_3813,N_2337,N_2060);
nand U3814 (N_3814,N_2989,N_2967);
and U3815 (N_3815,N_2168,N_2306);
nand U3816 (N_3816,N_2230,N_2390);
or U3817 (N_3817,N_2736,N_2147);
nor U3818 (N_3818,N_2903,N_2254);
and U3819 (N_3819,N_2194,N_2511);
and U3820 (N_3820,N_2153,N_2208);
and U3821 (N_3821,N_2198,N_2370);
xnor U3822 (N_3822,N_2334,N_2650);
nand U3823 (N_3823,N_2651,N_2483);
nor U3824 (N_3824,N_2106,N_2420);
nor U3825 (N_3825,N_2303,N_2363);
nor U3826 (N_3826,N_2137,N_2681);
nand U3827 (N_3827,N_2082,N_2398);
nand U3828 (N_3828,N_2089,N_2611);
nor U3829 (N_3829,N_2560,N_2073);
xor U3830 (N_3830,N_2852,N_2709);
nand U3831 (N_3831,N_2162,N_2289);
nand U3832 (N_3832,N_2727,N_2327);
nand U3833 (N_3833,N_2069,N_2106);
or U3834 (N_3834,N_2412,N_2831);
and U3835 (N_3835,N_2244,N_2465);
or U3836 (N_3836,N_2866,N_2008);
and U3837 (N_3837,N_2552,N_2123);
and U3838 (N_3838,N_2663,N_2592);
or U3839 (N_3839,N_2782,N_2698);
nor U3840 (N_3840,N_2240,N_2786);
nor U3841 (N_3841,N_2288,N_2460);
nor U3842 (N_3842,N_2397,N_2703);
and U3843 (N_3843,N_2353,N_2689);
nor U3844 (N_3844,N_2147,N_2822);
and U3845 (N_3845,N_2774,N_2647);
and U3846 (N_3846,N_2775,N_2103);
nor U3847 (N_3847,N_2244,N_2095);
nor U3848 (N_3848,N_2778,N_2010);
and U3849 (N_3849,N_2521,N_2390);
and U3850 (N_3850,N_2385,N_2680);
nor U3851 (N_3851,N_2303,N_2283);
or U3852 (N_3852,N_2223,N_2162);
nor U3853 (N_3853,N_2058,N_2279);
nor U3854 (N_3854,N_2502,N_2178);
nor U3855 (N_3855,N_2675,N_2029);
nor U3856 (N_3856,N_2479,N_2778);
nor U3857 (N_3857,N_2496,N_2986);
nor U3858 (N_3858,N_2922,N_2505);
nand U3859 (N_3859,N_2213,N_2971);
nor U3860 (N_3860,N_2873,N_2765);
nand U3861 (N_3861,N_2699,N_2815);
nor U3862 (N_3862,N_2058,N_2791);
and U3863 (N_3863,N_2987,N_2151);
nor U3864 (N_3864,N_2269,N_2864);
or U3865 (N_3865,N_2128,N_2994);
nor U3866 (N_3866,N_2023,N_2905);
nor U3867 (N_3867,N_2656,N_2809);
and U3868 (N_3868,N_2300,N_2109);
or U3869 (N_3869,N_2707,N_2379);
nor U3870 (N_3870,N_2503,N_2161);
or U3871 (N_3871,N_2872,N_2720);
nor U3872 (N_3872,N_2816,N_2841);
and U3873 (N_3873,N_2605,N_2795);
and U3874 (N_3874,N_2319,N_2101);
or U3875 (N_3875,N_2200,N_2317);
nor U3876 (N_3876,N_2733,N_2827);
nand U3877 (N_3877,N_2035,N_2906);
nor U3878 (N_3878,N_2427,N_2021);
and U3879 (N_3879,N_2347,N_2082);
nor U3880 (N_3880,N_2741,N_2608);
or U3881 (N_3881,N_2280,N_2289);
nor U3882 (N_3882,N_2092,N_2445);
nor U3883 (N_3883,N_2740,N_2267);
nand U3884 (N_3884,N_2944,N_2776);
nor U3885 (N_3885,N_2982,N_2571);
and U3886 (N_3886,N_2677,N_2765);
or U3887 (N_3887,N_2901,N_2647);
or U3888 (N_3888,N_2257,N_2054);
nor U3889 (N_3889,N_2530,N_2178);
nor U3890 (N_3890,N_2441,N_2014);
nand U3891 (N_3891,N_2418,N_2788);
nor U3892 (N_3892,N_2541,N_2994);
nor U3893 (N_3893,N_2725,N_2273);
nor U3894 (N_3894,N_2892,N_2303);
and U3895 (N_3895,N_2937,N_2305);
and U3896 (N_3896,N_2415,N_2995);
nand U3897 (N_3897,N_2972,N_2045);
nor U3898 (N_3898,N_2480,N_2870);
and U3899 (N_3899,N_2709,N_2066);
nand U3900 (N_3900,N_2000,N_2088);
and U3901 (N_3901,N_2244,N_2101);
xor U3902 (N_3902,N_2517,N_2083);
and U3903 (N_3903,N_2380,N_2542);
and U3904 (N_3904,N_2520,N_2679);
nand U3905 (N_3905,N_2300,N_2084);
and U3906 (N_3906,N_2101,N_2879);
or U3907 (N_3907,N_2385,N_2566);
or U3908 (N_3908,N_2272,N_2165);
xor U3909 (N_3909,N_2678,N_2591);
nor U3910 (N_3910,N_2542,N_2269);
nor U3911 (N_3911,N_2893,N_2053);
nand U3912 (N_3912,N_2362,N_2819);
and U3913 (N_3913,N_2601,N_2199);
and U3914 (N_3914,N_2699,N_2621);
nand U3915 (N_3915,N_2407,N_2787);
or U3916 (N_3916,N_2188,N_2555);
xor U3917 (N_3917,N_2973,N_2998);
or U3918 (N_3918,N_2558,N_2887);
and U3919 (N_3919,N_2588,N_2347);
nor U3920 (N_3920,N_2150,N_2137);
and U3921 (N_3921,N_2806,N_2157);
nor U3922 (N_3922,N_2771,N_2056);
and U3923 (N_3923,N_2239,N_2320);
nor U3924 (N_3924,N_2206,N_2379);
and U3925 (N_3925,N_2849,N_2549);
and U3926 (N_3926,N_2598,N_2211);
nand U3927 (N_3927,N_2498,N_2712);
nand U3928 (N_3928,N_2051,N_2511);
and U3929 (N_3929,N_2181,N_2947);
and U3930 (N_3930,N_2927,N_2504);
and U3931 (N_3931,N_2114,N_2654);
nand U3932 (N_3932,N_2104,N_2328);
nor U3933 (N_3933,N_2699,N_2586);
nand U3934 (N_3934,N_2777,N_2841);
nand U3935 (N_3935,N_2735,N_2712);
and U3936 (N_3936,N_2349,N_2677);
and U3937 (N_3937,N_2500,N_2527);
nand U3938 (N_3938,N_2850,N_2554);
nor U3939 (N_3939,N_2707,N_2352);
nand U3940 (N_3940,N_2892,N_2235);
and U3941 (N_3941,N_2084,N_2627);
and U3942 (N_3942,N_2855,N_2943);
nand U3943 (N_3943,N_2908,N_2951);
and U3944 (N_3944,N_2991,N_2668);
nor U3945 (N_3945,N_2474,N_2233);
or U3946 (N_3946,N_2346,N_2357);
or U3947 (N_3947,N_2617,N_2761);
nand U3948 (N_3948,N_2704,N_2446);
nor U3949 (N_3949,N_2316,N_2912);
or U3950 (N_3950,N_2396,N_2497);
nor U3951 (N_3951,N_2399,N_2067);
or U3952 (N_3952,N_2642,N_2561);
nand U3953 (N_3953,N_2342,N_2564);
and U3954 (N_3954,N_2562,N_2355);
nor U3955 (N_3955,N_2983,N_2725);
and U3956 (N_3956,N_2506,N_2376);
nor U3957 (N_3957,N_2128,N_2561);
nand U3958 (N_3958,N_2377,N_2373);
and U3959 (N_3959,N_2648,N_2541);
and U3960 (N_3960,N_2607,N_2998);
nor U3961 (N_3961,N_2131,N_2266);
nand U3962 (N_3962,N_2643,N_2008);
or U3963 (N_3963,N_2359,N_2836);
or U3964 (N_3964,N_2573,N_2337);
or U3965 (N_3965,N_2962,N_2515);
nand U3966 (N_3966,N_2679,N_2229);
and U3967 (N_3967,N_2101,N_2235);
and U3968 (N_3968,N_2406,N_2672);
or U3969 (N_3969,N_2291,N_2087);
and U3970 (N_3970,N_2939,N_2739);
nand U3971 (N_3971,N_2840,N_2543);
nand U3972 (N_3972,N_2826,N_2067);
nand U3973 (N_3973,N_2883,N_2620);
or U3974 (N_3974,N_2324,N_2397);
nand U3975 (N_3975,N_2282,N_2122);
nand U3976 (N_3976,N_2763,N_2327);
nand U3977 (N_3977,N_2592,N_2253);
nand U3978 (N_3978,N_2548,N_2830);
and U3979 (N_3979,N_2377,N_2708);
nor U3980 (N_3980,N_2156,N_2466);
or U3981 (N_3981,N_2898,N_2466);
and U3982 (N_3982,N_2825,N_2607);
and U3983 (N_3983,N_2931,N_2030);
or U3984 (N_3984,N_2124,N_2255);
nor U3985 (N_3985,N_2486,N_2219);
and U3986 (N_3986,N_2261,N_2269);
nor U3987 (N_3987,N_2256,N_2128);
or U3988 (N_3988,N_2312,N_2060);
nand U3989 (N_3989,N_2134,N_2533);
and U3990 (N_3990,N_2347,N_2739);
nand U3991 (N_3991,N_2953,N_2652);
and U3992 (N_3992,N_2924,N_2233);
nand U3993 (N_3993,N_2504,N_2780);
nand U3994 (N_3994,N_2588,N_2507);
nor U3995 (N_3995,N_2995,N_2935);
nand U3996 (N_3996,N_2839,N_2125);
nor U3997 (N_3997,N_2725,N_2027);
nor U3998 (N_3998,N_2472,N_2374);
and U3999 (N_3999,N_2205,N_2123);
nor U4000 (N_4000,N_3091,N_3568);
nor U4001 (N_4001,N_3592,N_3368);
nand U4002 (N_4002,N_3652,N_3215);
nor U4003 (N_4003,N_3617,N_3935);
nand U4004 (N_4004,N_3209,N_3114);
and U4005 (N_4005,N_3983,N_3884);
or U4006 (N_4006,N_3280,N_3126);
nand U4007 (N_4007,N_3943,N_3538);
and U4008 (N_4008,N_3129,N_3377);
or U4009 (N_4009,N_3949,N_3974);
nand U4010 (N_4010,N_3885,N_3536);
or U4011 (N_4011,N_3214,N_3840);
or U4012 (N_4012,N_3515,N_3271);
or U4013 (N_4013,N_3781,N_3729);
nor U4014 (N_4014,N_3450,N_3939);
and U4015 (N_4015,N_3934,N_3494);
or U4016 (N_4016,N_3422,N_3995);
nand U4017 (N_4017,N_3531,N_3276);
xnor U4018 (N_4018,N_3660,N_3644);
and U4019 (N_4019,N_3703,N_3875);
nor U4020 (N_4020,N_3680,N_3095);
nand U4021 (N_4021,N_3544,N_3292);
nand U4022 (N_4022,N_3951,N_3820);
nor U4023 (N_4023,N_3487,N_3208);
or U4024 (N_4024,N_3321,N_3927);
nor U4025 (N_4025,N_3355,N_3527);
nor U4026 (N_4026,N_3365,N_3948);
and U4027 (N_4027,N_3014,N_3107);
or U4028 (N_4028,N_3813,N_3818);
nand U4029 (N_4029,N_3438,N_3746);
or U4030 (N_4030,N_3491,N_3678);
nand U4031 (N_4031,N_3191,N_3728);
or U4032 (N_4032,N_3685,N_3655);
or U4033 (N_4033,N_3203,N_3798);
nand U4034 (N_4034,N_3077,N_3941);
or U4035 (N_4035,N_3334,N_3518);
nor U4036 (N_4036,N_3714,N_3398);
nand U4037 (N_4037,N_3325,N_3111);
and U4038 (N_4038,N_3539,N_3643);
nor U4039 (N_4039,N_3912,N_3869);
and U4040 (N_4040,N_3137,N_3453);
nand U4041 (N_4041,N_3289,N_3360);
nand U4042 (N_4042,N_3754,N_3174);
and U4043 (N_4043,N_3513,N_3201);
or U4044 (N_4044,N_3026,N_3525);
and U4045 (N_4045,N_3353,N_3339);
nor U4046 (N_4046,N_3159,N_3767);
and U4047 (N_4047,N_3222,N_3615);
nor U4048 (N_4048,N_3488,N_3141);
nand U4049 (N_4049,N_3633,N_3027);
and U4050 (N_4050,N_3390,N_3199);
or U4051 (N_4051,N_3895,N_3665);
nand U4052 (N_4052,N_3822,N_3247);
or U4053 (N_4053,N_3439,N_3435);
nor U4054 (N_4054,N_3018,N_3792);
or U4055 (N_4055,N_3661,N_3385);
and U4056 (N_4056,N_3184,N_3128);
and U4057 (N_4057,N_3032,N_3379);
and U4058 (N_4058,N_3606,N_3858);
or U4059 (N_4059,N_3079,N_3192);
or U4060 (N_4060,N_3521,N_3853);
or U4061 (N_4061,N_3268,N_3735);
and U4062 (N_4062,N_3666,N_3483);
or U4063 (N_4063,N_3534,N_3696);
nand U4064 (N_4064,N_3473,N_3601);
nor U4065 (N_4065,N_3337,N_3374);
and U4066 (N_4066,N_3082,N_3641);
or U4067 (N_4067,N_3358,N_3413);
or U4068 (N_4068,N_3631,N_3711);
nand U4069 (N_4069,N_3153,N_3252);
nand U4070 (N_4070,N_3824,N_3973);
or U4071 (N_4071,N_3731,N_3348);
nor U4072 (N_4072,N_3849,N_3019);
nor U4073 (N_4073,N_3761,N_3725);
or U4074 (N_4074,N_3784,N_3050);
or U4075 (N_4075,N_3833,N_3636);
and U4076 (N_4076,N_3599,N_3257);
nand U4077 (N_4077,N_3419,N_3647);
nor U4078 (N_4078,N_3877,N_3844);
xor U4079 (N_4079,N_3476,N_3477);
or U4080 (N_4080,N_3359,N_3412);
or U4081 (N_4081,N_3284,N_3426);
or U4082 (N_4082,N_3857,N_3765);
nand U4083 (N_4083,N_3656,N_3421);
nand U4084 (N_4084,N_3607,N_3965);
and U4085 (N_4085,N_3352,N_3492);
or U4086 (N_4086,N_3382,N_3416);
nand U4087 (N_4087,N_3320,N_3024);
or U4088 (N_4088,N_3505,N_3464);
nor U4089 (N_4089,N_3418,N_3575);
nor U4090 (N_4090,N_3845,N_3627);
nand U4091 (N_4091,N_3256,N_3381);
and U4092 (N_4092,N_3996,N_3751);
nand U4093 (N_4093,N_3386,N_3445);
nor U4094 (N_4094,N_3241,N_3094);
or U4095 (N_4095,N_3688,N_3790);
or U4096 (N_4096,N_3902,N_3580);
and U4097 (N_4097,N_3530,N_3806);
or U4098 (N_4098,N_3296,N_3261);
xor U4099 (N_4099,N_3611,N_3344);
and U4100 (N_4100,N_3238,N_3682);
and U4101 (N_4101,N_3290,N_3231);
or U4102 (N_4102,N_3747,N_3179);
or U4103 (N_4103,N_3340,N_3710);
nor U4104 (N_4104,N_3451,N_3740);
nor U4105 (N_4105,N_3994,N_3171);
xnor U4106 (N_4106,N_3783,N_3712);
nor U4107 (N_4107,N_3506,N_3039);
nor U4108 (N_4108,N_3403,N_3275);
and U4109 (N_4109,N_3038,N_3345);
nor U4110 (N_4110,N_3613,N_3304);
nand U4111 (N_4111,N_3883,N_3232);
and U4112 (N_4112,N_3303,N_3136);
and U4113 (N_4113,N_3975,N_3173);
nand U4114 (N_4114,N_3210,N_3444);
nor U4115 (N_4115,N_3429,N_3910);
nor U4116 (N_4116,N_3187,N_3063);
nor U4117 (N_4117,N_3244,N_3075);
or U4118 (N_4118,N_3100,N_3855);
and U4119 (N_4119,N_3831,N_3763);
and U4120 (N_4120,N_3431,N_3604);
and U4121 (N_4121,N_3332,N_3808);
xnor U4122 (N_4122,N_3677,N_3088);
and U4123 (N_4123,N_3499,N_3070);
nor U4124 (N_4124,N_3559,N_3990);
or U4125 (N_4125,N_3931,N_3762);
nand U4126 (N_4126,N_3594,N_3102);
nor U4127 (N_4127,N_3131,N_3417);
nor U4128 (N_4128,N_3484,N_3624);
and U4129 (N_4129,N_3732,N_3981);
nand U4130 (N_4130,N_3928,N_3501);
nor U4131 (N_4131,N_3356,N_3821);
and U4132 (N_4132,N_3291,N_3906);
nor U4133 (N_4133,N_3794,N_3228);
or U4134 (N_4134,N_3850,N_3964);
or U4135 (N_4135,N_3540,N_3157);
or U4136 (N_4136,N_3098,N_3814);
or U4137 (N_4137,N_3793,N_3579);
nor U4138 (N_4138,N_3148,N_3985);
nor U4139 (N_4139,N_3908,N_3519);
or U4140 (N_4140,N_3589,N_3218);
and U4141 (N_4141,N_3898,N_3581);
nand U4142 (N_4142,N_3860,N_3968);
nand U4143 (N_4143,N_3090,N_3523);
nor U4144 (N_4144,N_3512,N_3913);
nand U4145 (N_4145,N_3625,N_3260);
nand U4146 (N_4146,N_3901,N_3073);
xnor U4147 (N_4147,N_3447,N_3852);
and U4148 (N_4148,N_3741,N_3759);
nor U4149 (N_4149,N_3915,N_3395);
nor U4150 (N_4150,N_3470,N_3460);
and U4151 (N_4151,N_3800,N_3757);
or U4152 (N_4152,N_3255,N_3378);
and U4153 (N_4153,N_3329,N_3726);
and U4154 (N_4154,N_3086,N_3893);
nand U4155 (N_4155,N_3286,N_3502);
or U4156 (N_4156,N_3616,N_3701);
or U4157 (N_4157,N_3122,N_3892);
nor U4158 (N_4158,N_3467,N_3245);
nand U4159 (N_4159,N_3497,N_3341);
nor U4160 (N_4160,N_3971,N_3957);
or U4161 (N_4161,N_3671,N_3002);
nand U4162 (N_4162,N_3772,N_3380);
and U4163 (N_4163,N_3586,N_3917);
and U4164 (N_4164,N_3240,N_3155);
nand U4165 (N_4165,N_3197,N_3015);
or U4166 (N_4166,N_3768,N_3163);
and U4167 (N_4167,N_3557,N_3654);
nor U4168 (N_4168,N_3376,N_3988);
and U4169 (N_4169,N_3999,N_3319);
and U4170 (N_4170,N_3442,N_3554);
or U4171 (N_4171,N_3393,N_3524);
and U4172 (N_4172,N_3269,N_3425);
or U4173 (N_4173,N_3897,N_3614);
nand U4174 (N_4174,N_3135,N_3707);
and U4175 (N_4175,N_3862,N_3236);
nand U4176 (N_4176,N_3874,N_3391);
or U4177 (N_4177,N_3550,N_3495);
and U4178 (N_4178,N_3387,N_3817);
nand U4179 (N_4179,N_3206,N_3097);
and U4180 (N_4180,N_3582,N_3738);
and U4181 (N_4181,N_3574,N_3577);
nor U4182 (N_4182,N_3803,N_3634);
and U4183 (N_4183,N_3828,N_3904);
and U4184 (N_4184,N_3169,N_3561);
and U4185 (N_4185,N_3055,N_3318);
nand U4186 (N_4186,N_3936,N_3733);
and U4187 (N_4187,N_3944,N_3016);
nand U4188 (N_4188,N_3593,N_3327);
and U4189 (N_4189,N_3013,N_3590);
nand U4190 (N_4190,N_3051,N_3202);
or U4191 (N_4191,N_3773,N_3096);
nand U4192 (N_4192,N_3062,N_3791);
or U4193 (N_4193,N_3558,N_3388);
nand U4194 (N_4194,N_3724,N_3270);
or U4195 (N_4195,N_3645,N_3000);
nand U4196 (N_4196,N_3695,N_3690);
nor U4197 (N_4197,N_3775,N_3144);
nor U4198 (N_4198,N_3437,N_3500);
nor U4199 (N_4199,N_3363,N_3493);
or U4200 (N_4200,N_3583,N_3743);
or U4201 (N_4201,N_3342,N_3952);
and U4202 (N_4202,N_3886,N_3839);
and U4203 (N_4203,N_3890,N_3399);
nand U4204 (N_4204,N_3749,N_3409);
nand U4205 (N_4205,N_3121,N_3190);
nor U4206 (N_4206,N_3151,N_3816);
nand U4207 (N_4207,N_3003,N_3720);
nor U4208 (N_4208,N_3258,N_3408);
nand U4209 (N_4209,N_3116,N_3675);
and U4210 (N_4210,N_3044,N_3123);
nand U4211 (N_4211,N_3030,N_3668);
or U4212 (N_4212,N_3204,N_3942);
nor U4213 (N_4213,N_3310,N_3597);
nand U4214 (N_4214,N_3861,N_3864);
and U4215 (N_4215,N_3980,N_3150);
nor U4216 (N_4216,N_3600,N_3838);
and U4217 (N_4217,N_3306,N_3804);
nor U4218 (N_4218,N_3715,N_3043);
nor U4219 (N_4219,N_3237,N_3972);
and U4220 (N_4220,N_3008,N_3516);
nand U4221 (N_4221,N_3357,N_3313);
or U4222 (N_4222,N_3925,N_3452);
nand U4223 (N_4223,N_3650,N_3533);
or U4224 (N_4224,N_3630,N_3737);
and U4225 (N_4225,N_3713,N_3991);
nand U4226 (N_4226,N_3955,N_3087);
xnor U4227 (N_4227,N_3481,N_3730);
nor U4228 (N_4228,N_3056,N_3074);
and U4229 (N_4229,N_3273,N_3958);
and U4230 (N_4230,N_3588,N_3653);
nand U4231 (N_4231,N_3347,N_3177);
nor U4232 (N_4232,N_3428,N_3555);
or U4233 (N_4233,N_3560,N_3946);
and U4234 (N_4234,N_3145,N_3287);
nor U4235 (N_4235,N_3708,N_3045);
xnor U4236 (N_4236,N_3672,N_3295);
nor U4237 (N_4237,N_3367,N_3785);
and U4238 (N_4238,N_3702,N_3940);
nand U4239 (N_4239,N_3246,N_3219);
nand U4240 (N_4240,N_3127,N_3520);
and U4241 (N_4241,N_3632,N_3022);
and U4242 (N_4242,N_3970,N_3160);
or U4243 (N_4243,N_3982,N_3101);
nor U4244 (N_4244,N_3278,N_3830);
nand U4245 (N_4245,N_3338,N_3311);
nor U4246 (N_4246,N_3716,N_3528);
and U4247 (N_4247,N_3081,N_3189);
and U4248 (N_4248,N_3400,N_3143);
and U4249 (N_4249,N_3001,N_3254);
and U4250 (N_4250,N_3529,N_3262);
nor U4251 (N_4251,N_3693,N_3549);
and U4252 (N_4252,N_3253,N_3036);
nand U4253 (N_4253,N_3508,N_3446);
and U4254 (N_4254,N_3788,N_3683);
or U4255 (N_4255,N_3349,N_3774);
xnor U4256 (N_4256,N_3796,N_3216);
or U4257 (N_4257,N_3182,N_3023);
nand U4258 (N_4258,N_3124,N_3921);
nand U4259 (N_4259,N_3322,N_3224);
and U4260 (N_4260,N_3595,N_3078);
nor U4261 (N_4261,N_3891,N_3938);
nor U4262 (N_4262,N_3109,N_3308);
nor U4263 (N_4263,N_3134,N_3293);
nand U4264 (N_4264,N_3674,N_3361);
nor U4265 (N_4265,N_3571,N_3778);
nor U4266 (N_4266,N_3040,N_3681);
nand U4267 (N_4267,N_3220,N_3548);
and U4268 (N_4268,N_3234,N_3061);
or U4269 (N_4269,N_3642,N_3007);
nor U4270 (N_4270,N_3805,N_3465);
nand U4271 (N_4271,N_3602,N_3384);
or U4272 (N_4272,N_3842,N_3119);
nand U4273 (N_4273,N_3552,N_3221);
nor U4274 (N_4274,N_3542,N_3006);
or U4275 (N_4275,N_3919,N_3829);
nand U4276 (N_4276,N_3156,N_3166);
and U4277 (N_4277,N_3049,N_3758);
and U4278 (N_4278,N_3383,N_3541);
nor U4279 (N_4279,N_3037,N_3401);
and U4280 (N_4280,N_3612,N_3092);
or U4281 (N_4281,N_3866,N_3371);
nand U4282 (N_4282,N_3066,N_3727);
xor U4283 (N_4283,N_3054,N_3510);
and U4284 (N_4284,N_3835,N_3937);
and U4285 (N_4285,N_3423,N_3212);
or U4286 (N_4286,N_3887,N_3468);
nor U4287 (N_4287,N_3354,N_3503);
and U4288 (N_4288,N_3362,N_3670);
or U4289 (N_4289,N_3264,N_3563);
or U4290 (N_4290,N_3277,N_3640);
nand U4291 (N_4291,N_3099,N_3879);
and U4292 (N_4292,N_3432,N_3198);
and U4293 (N_4293,N_3230,N_3474);
nand U4294 (N_4294,N_3300,N_3139);
or U4295 (N_4295,N_3578,N_3689);
nor U4296 (N_4296,N_3158,N_3479);
or U4297 (N_4297,N_3165,N_3837);
nor U4298 (N_4298,N_3526,N_3251);
or U4299 (N_4299,N_3691,N_3011);
or U4300 (N_4300,N_3553,N_3605);
and U4301 (N_4301,N_3977,N_3882);
nor U4302 (N_4302,N_3142,N_3415);
or U4303 (N_4303,N_3795,N_3229);
nor U4304 (N_4304,N_3797,N_3807);
and U4305 (N_4305,N_3461,N_3265);
nor U4306 (N_4306,N_3048,N_3744);
and U4307 (N_4307,N_3181,N_3623);
nand U4308 (N_4308,N_3427,N_3603);
or U4309 (N_4309,N_3889,N_3802);
nand U4310 (N_4310,N_3279,N_3718);
and U4311 (N_4311,N_3776,N_3926);
or U4312 (N_4312,N_3962,N_3809);
and U4313 (N_4313,N_3755,N_3164);
or U4314 (N_4314,N_3414,N_3335);
nand U4315 (N_4315,N_3351,N_3454);
nor U4316 (N_4316,N_3175,N_3108);
nor U4317 (N_4317,N_3004,N_3125);
and U4318 (N_4318,N_3694,N_3462);
and U4319 (N_4319,N_3152,N_3294);
nand U4320 (N_4320,N_3847,N_3020);
or U4321 (N_4321,N_3243,N_3899);
nor U4322 (N_4322,N_3517,N_3424);
or U4323 (N_4323,N_3084,N_3281);
nand U4324 (N_4324,N_3932,N_3080);
and U4325 (N_4325,N_3113,N_3485);
nand U4326 (N_4326,N_3771,N_3992);
or U4327 (N_4327,N_3396,N_3609);
or U4328 (N_4328,N_3748,N_3411);
and U4329 (N_4329,N_3639,N_3047);
nand U4330 (N_4330,N_3779,N_3878);
nand U4331 (N_4331,N_3021,N_3679);
nand U4332 (N_4332,N_3005,N_3811);
and U4333 (N_4333,N_3213,N_3698);
and U4334 (N_4334,N_3035,N_3226);
xnor U4335 (N_4335,N_3498,N_3140);
and U4336 (N_4336,N_3865,N_3967);
and U4337 (N_4337,N_3118,N_3596);
nor U4338 (N_4338,N_3619,N_3194);
or U4339 (N_4339,N_3333,N_3556);
nor U4340 (N_4340,N_3402,N_3282);
and U4341 (N_4341,N_3343,N_3176);
and U4342 (N_4342,N_3350,N_3819);
nor U4343 (N_4343,N_3172,N_3188);
xnor U4344 (N_4344,N_3721,N_3914);
or U4345 (N_4345,N_3907,N_3193);
nor U4346 (N_4346,N_3638,N_3302);
or U4347 (N_4347,N_3288,N_3305);
and U4348 (N_4348,N_3881,N_3285);
or U4349 (N_4349,N_3433,N_3394);
nand U4350 (N_4350,N_3966,N_3430);
nand U4351 (N_4351,N_3659,N_3998);
and U4352 (N_4352,N_3871,N_3489);
nand U4353 (N_4353,N_3083,N_3610);
nand U4354 (N_4354,N_3532,N_3834);
and U4355 (N_4355,N_3138,N_3239);
or U4356 (N_4356,N_3598,N_3103);
or U4357 (N_4357,N_3205,N_3186);
nand U4358 (N_4358,N_3922,N_3770);
nand U4359 (N_4359,N_3764,N_3537);
and U4360 (N_4360,N_3584,N_3217);
nand U4361 (N_4361,N_3826,N_3298);
nand U4362 (N_4362,N_3183,N_3168);
or U4363 (N_4363,N_3449,N_3832);
and U4364 (N_4364,N_3328,N_3976);
nor U4365 (N_4365,N_3064,N_3567);
nand U4366 (N_4366,N_3331,N_3905);
or U4367 (N_4367,N_3918,N_3250);
nor U4368 (N_4368,N_3662,N_3566);
nor U4369 (N_4369,N_3407,N_3509);
nand U4370 (N_4370,N_3149,N_3736);
nor U4371 (N_4371,N_3545,N_3315);
or U4372 (N_4372,N_3185,N_3397);
and U4373 (N_4373,N_3233,N_3562);
nor U4374 (N_4374,N_3041,N_3072);
nand U4375 (N_4375,N_3069,N_3060);
nand U4376 (N_4376,N_3456,N_3872);
or U4377 (N_4377,N_3112,N_3903);
and U4378 (N_4378,N_3272,N_3330);
nor U4379 (N_4379,N_3207,N_3745);
xor U4380 (N_4380,N_3565,N_3455);
or U4381 (N_4381,N_3211,N_3507);
nor U4382 (N_4382,N_3734,N_3511);
and U4383 (N_4383,N_3434,N_3009);
and U4384 (N_4384,N_3753,N_3259);
nor U4385 (N_4385,N_3742,N_3723);
and U4386 (N_4386,N_3389,N_3564);
nand U4387 (N_4387,N_3167,N_3370);
nor U4388 (N_4388,N_3482,N_3490);
or U4389 (N_4389,N_3916,N_3405);
and U4390 (N_4390,N_3993,N_3686);
nand U4391 (N_4391,N_3267,N_3900);
and U4392 (N_4392,N_3618,N_3873);
nor U4393 (N_4393,N_3104,N_3441);
nand U4394 (N_4394,N_3752,N_3105);
nand U4395 (N_4395,N_3366,N_3046);
or U4396 (N_4396,N_3458,N_3894);
and U4397 (N_4397,N_3876,N_3547);
nor U4398 (N_4398,N_3297,N_3225);
nand U4399 (N_4399,N_3572,N_3896);
nor U4400 (N_4400,N_3719,N_3420);
and U4401 (N_4401,N_3722,N_3963);
and U4402 (N_4402,N_3989,N_3651);
nand U4403 (N_4403,N_3249,N_3573);
nand U4404 (N_4404,N_3274,N_3859);
and U4405 (N_4405,N_3504,N_3868);
nor U4406 (N_4406,N_3132,N_3546);
nor U4407 (N_4407,N_3375,N_3443);
nand U4408 (N_4408,N_3827,N_3635);
nand U4409 (N_4409,N_3475,N_3010);
nand U4410 (N_4410,N_3115,N_3283);
or U4411 (N_4411,N_3486,N_3620);
nor U4412 (N_4412,N_3266,N_3042);
and U4413 (N_4413,N_3130,N_3029);
and U4414 (N_4414,N_3480,N_3033);
and U4415 (N_4415,N_3836,N_3782);
nand U4416 (N_4416,N_3825,N_3629);
and U4417 (N_4417,N_3664,N_3930);
or U4418 (N_4418,N_3314,N_3496);
nand U4419 (N_4419,N_3697,N_3017);
nand U4420 (N_4420,N_3848,N_3961);
and U4421 (N_4421,N_3323,N_3769);
nand U4422 (N_4422,N_3025,N_3178);
and U4423 (N_4423,N_3570,N_3888);
and U4424 (N_4424,N_3841,N_3404);
and U4425 (N_4425,N_3801,N_3705);
and U4426 (N_4426,N_3076,N_3522);
nand U4427 (N_4427,N_3856,N_3463);
nand U4428 (N_4428,N_3622,N_3760);
and U4429 (N_4429,N_3823,N_3110);
nor U4430 (N_4430,N_3923,N_3756);
nor U4431 (N_4431,N_3997,N_3669);
nor U4432 (N_4432,N_3789,N_3154);
nand U4433 (N_4433,N_3200,N_3777);
nand U4434 (N_4434,N_3704,N_3543);
or U4435 (N_4435,N_3945,N_3471);
and U4436 (N_4436,N_3863,N_3960);
nand U4437 (N_4437,N_3956,N_3089);
nor U4438 (N_4438,N_3846,N_3684);
nor U4439 (N_4439,N_3920,N_3626);
or U4440 (N_4440,N_3373,N_3478);
or U4441 (N_4441,N_3780,N_3787);
or U4442 (N_4442,N_3706,N_3929);
or U4443 (N_4443,N_3309,N_3059);
nand U4444 (N_4444,N_3301,N_3223);
nor U4445 (N_4445,N_3459,N_3242);
nand U4446 (N_4446,N_3621,N_3709);
nand U4447 (N_4447,N_3587,N_3067);
or U4448 (N_4448,N_3117,N_3068);
nand U4449 (N_4449,N_3569,N_3436);
or U4450 (N_4450,N_3053,N_3440);
or U4451 (N_4451,N_3648,N_3448);
nand U4452 (N_4452,N_3161,N_3933);
and U4453 (N_4453,N_3472,N_3954);
nand U4454 (N_4454,N_3608,N_3576);
nor U4455 (N_4455,N_3263,N_3316);
and U4456 (N_4456,N_3034,N_3085);
or U4457 (N_4457,N_3248,N_3146);
and U4458 (N_4458,N_3180,N_3854);
and U4459 (N_4459,N_3364,N_3120);
or U4460 (N_4460,N_3299,N_3317);
and U4461 (N_4461,N_3799,N_3810);
and U4462 (N_4462,N_3466,N_3924);
and U4463 (N_4463,N_3687,N_3312);
and U4464 (N_4464,N_3766,N_3667);
nor U4465 (N_4465,N_3815,N_3699);
nor U4466 (N_4466,N_3700,N_3880);
or U4467 (N_4467,N_3843,N_3984);
xnor U4468 (N_4468,N_3646,N_3392);
nand U4469 (N_4469,N_3551,N_3867);
nand U4470 (N_4470,N_3978,N_3133);
nor U4471 (N_4471,N_3739,N_3028);
xnor U4472 (N_4472,N_3057,N_3065);
nand U4473 (N_4473,N_3324,N_3870);
or U4474 (N_4474,N_3093,N_3372);
nor U4475 (N_4475,N_3195,N_3469);
or U4476 (N_4476,N_3147,N_3947);
nor U4477 (N_4477,N_3717,N_3969);
and U4478 (N_4478,N_3170,N_3346);
or U4479 (N_4479,N_3658,N_3786);
nor U4480 (N_4480,N_3227,N_3196);
and U4481 (N_4481,N_3326,N_3406);
xor U4482 (N_4482,N_3410,N_3457);
or U4483 (N_4483,N_3012,N_3909);
nor U4484 (N_4484,N_3986,N_3307);
nor U4485 (N_4485,N_3235,N_3987);
or U4486 (N_4486,N_3336,N_3676);
or U4487 (N_4487,N_3637,N_3750);
or U4488 (N_4488,N_3628,N_3514);
and U4489 (N_4489,N_3535,N_3162);
and U4490 (N_4490,N_3851,N_3911);
xor U4491 (N_4491,N_3663,N_3106);
or U4492 (N_4492,N_3812,N_3673);
or U4493 (N_4493,N_3979,N_3959);
nand U4494 (N_4494,N_3071,N_3585);
or U4495 (N_4495,N_3052,N_3369);
xnor U4496 (N_4496,N_3649,N_3058);
and U4497 (N_4497,N_3591,N_3692);
and U4498 (N_4498,N_3950,N_3953);
or U4499 (N_4499,N_3031,N_3657);
or U4500 (N_4500,N_3220,N_3171);
nand U4501 (N_4501,N_3608,N_3607);
and U4502 (N_4502,N_3372,N_3262);
nand U4503 (N_4503,N_3450,N_3373);
nor U4504 (N_4504,N_3185,N_3390);
or U4505 (N_4505,N_3322,N_3835);
nor U4506 (N_4506,N_3788,N_3052);
nand U4507 (N_4507,N_3033,N_3511);
nand U4508 (N_4508,N_3929,N_3952);
nor U4509 (N_4509,N_3476,N_3289);
or U4510 (N_4510,N_3813,N_3125);
nor U4511 (N_4511,N_3680,N_3929);
nor U4512 (N_4512,N_3028,N_3946);
nor U4513 (N_4513,N_3453,N_3748);
nand U4514 (N_4514,N_3035,N_3928);
and U4515 (N_4515,N_3718,N_3894);
or U4516 (N_4516,N_3415,N_3842);
nor U4517 (N_4517,N_3343,N_3302);
nor U4518 (N_4518,N_3693,N_3465);
or U4519 (N_4519,N_3589,N_3374);
nand U4520 (N_4520,N_3196,N_3596);
and U4521 (N_4521,N_3047,N_3124);
and U4522 (N_4522,N_3605,N_3664);
nand U4523 (N_4523,N_3425,N_3311);
nand U4524 (N_4524,N_3866,N_3187);
nor U4525 (N_4525,N_3871,N_3583);
and U4526 (N_4526,N_3751,N_3842);
or U4527 (N_4527,N_3365,N_3851);
or U4528 (N_4528,N_3683,N_3258);
or U4529 (N_4529,N_3191,N_3551);
and U4530 (N_4530,N_3934,N_3707);
and U4531 (N_4531,N_3834,N_3188);
nor U4532 (N_4532,N_3365,N_3777);
nand U4533 (N_4533,N_3839,N_3555);
or U4534 (N_4534,N_3292,N_3507);
nand U4535 (N_4535,N_3625,N_3356);
or U4536 (N_4536,N_3083,N_3595);
nand U4537 (N_4537,N_3914,N_3436);
or U4538 (N_4538,N_3354,N_3513);
or U4539 (N_4539,N_3722,N_3341);
nand U4540 (N_4540,N_3399,N_3683);
nand U4541 (N_4541,N_3581,N_3586);
nand U4542 (N_4542,N_3905,N_3649);
nand U4543 (N_4543,N_3547,N_3303);
and U4544 (N_4544,N_3182,N_3213);
nor U4545 (N_4545,N_3143,N_3883);
or U4546 (N_4546,N_3127,N_3700);
or U4547 (N_4547,N_3796,N_3144);
or U4548 (N_4548,N_3883,N_3817);
nor U4549 (N_4549,N_3193,N_3525);
xor U4550 (N_4550,N_3969,N_3319);
nand U4551 (N_4551,N_3519,N_3697);
nor U4552 (N_4552,N_3034,N_3671);
or U4553 (N_4553,N_3798,N_3794);
and U4554 (N_4554,N_3514,N_3992);
or U4555 (N_4555,N_3637,N_3005);
nand U4556 (N_4556,N_3601,N_3606);
xnor U4557 (N_4557,N_3166,N_3931);
nand U4558 (N_4558,N_3609,N_3046);
nand U4559 (N_4559,N_3032,N_3286);
nand U4560 (N_4560,N_3954,N_3518);
and U4561 (N_4561,N_3631,N_3571);
and U4562 (N_4562,N_3727,N_3793);
nor U4563 (N_4563,N_3062,N_3422);
nor U4564 (N_4564,N_3492,N_3886);
nor U4565 (N_4565,N_3916,N_3447);
or U4566 (N_4566,N_3581,N_3148);
nor U4567 (N_4567,N_3509,N_3989);
nand U4568 (N_4568,N_3857,N_3535);
and U4569 (N_4569,N_3675,N_3770);
or U4570 (N_4570,N_3017,N_3476);
or U4571 (N_4571,N_3095,N_3030);
nand U4572 (N_4572,N_3105,N_3438);
and U4573 (N_4573,N_3620,N_3959);
and U4574 (N_4574,N_3520,N_3497);
nand U4575 (N_4575,N_3857,N_3143);
xor U4576 (N_4576,N_3043,N_3813);
or U4577 (N_4577,N_3500,N_3256);
and U4578 (N_4578,N_3496,N_3435);
nand U4579 (N_4579,N_3199,N_3742);
nor U4580 (N_4580,N_3690,N_3063);
or U4581 (N_4581,N_3308,N_3991);
or U4582 (N_4582,N_3787,N_3031);
nor U4583 (N_4583,N_3235,N_3608);
or U4584 (N_4584,N_3040,N_3579);
and U4585 (N_4585,N_3808,N_3131);
nor U4586 (N_4586,N_3550,N_3524);
nor U4587 (N_4587,N_3554,N_3510);
and U4588 (N_4588,N_3672,N_3973);
nor U4589 (N_4589,N_3480,N_3381);
and U4590 (N_4590,N_3011,N_3427);
nand U4591 (N_4591,N_3786,N_3248);
nor U4592 (N_4592,N_3922,N_3487);
or U4593 (N_4593,N_3101,N_3204);
or U4594 (N_4594,N_3116,N_3368);
nor U4595 (N_4595,N_3409,N_3398);
nand U4596 (N_4596,N_3871,N_3385);
and U4597 (N_4597,N_3869,N_3491);
or U4598 (N_4598,N_3799,N_3312);
nand U4599 (N_4599,N_3836,N_3690);
or U4600 (N_4600,N_3687,N_3689);
nor U4601 (N_4601,N_3244,N_3755);
nand U4602 (N_4602,N_3969,N_3474);
or U4603 (N_4603,N_3654,N_3758);
or U4604 (N_4604,N_3406,N_3591);
or U4605 (N_4605,N_3063,N_3565);
nand U4606 (N_4606,N_3556,N_3706);
nor U4607 (N_4607,N_3168,N_3698);
and U4608 (N_4608,N_3450,N_3314);
xor U4609 (N_4609,N_3726,N_3649);
nor U4610 (N_4610,N_3131,N_3556);
or U4611 (N_4611,N_3917,N_3402);
and U4612 (N_4612,N_3521,N_3294);
nor U4613 (N_4613,N_3539,N_3349);
nor U4614 (N_4614,N_3699,N_3023);
or U4615 (N_4615,N_3261,N_3131);
or U4616 (N_4616,N_3196,N_3775);
and U4617 (N_4617,N_3226,N_3186);
or U4618 (N_4618,N_3787,N_3099);
nand U4619 (N_4619,N_3734,N_3769);
nand U4620 (N_4620,N_3922,N_3634);
and U4621 (N_4621,N_3188,N_3255);
and U4622 (N_4622,N_3969,N_3241);
nor U4623 (N_4623,N_3903,N_3595);
or U4624 (N_4624,N_3106,N_3985);
nand U4625 (N_4625,N_3009,N_3556);
nor U4626 (N_4626,N_3844,N_3487);
nor U4627 (N_4627,N_3353,N_3657);
nor U4628 (N_4628,N_3250,N_3700);
nand U4629 (N_4629,N_3931,N_3188);
nor U4630 (N_4630,N_3123,N_3546);
and U4631 (N_4631,N_3088,N_3914);
and U4632 (N_4632,N_3457,N_3306);
nand U4633 (N_4633,N_3060,N_3269);
and U4634 (N_4634,N_3479,N_3255);
and U4635 (N_4635,N_3215,N_3505);
nor U4636 (N_4636,N_3614,N_3019);
or U4637 (N_4637,N_3665,N_3705);
nand U4638 (N_4638,N_3473,N_3533);
nor U4639 (N_4639,N_3736,N_3439);
and U4640 (N_4640,N_3659,N_3172);
or U4641 (N_4641,N_3686,N_3469);
or U4642 (N_4642,N_3596,N_3289);
xor U4643 (N_4643,N_3389,N_3789);
or U4644 (N_4644,N_3770,N_3261);
and U4645 (N_4645,N_3148,N_3992);
nand U4646 (N_4646,N_3171,N_3475);
and U4647 (N_4647,N_3906,N_3557);
and U4648 (N_4648,N_3956,N_3986);
and U4649 (N_4649,N_3007,N_3278);
and U4650 (N_4650,N_3348,N_3324);
nand U4651 (N_4651,N_3273,N_3692);
and U4652 (N_4652,N_3440,N_3319);
nand U4653 (N_4653,N_3031,N_3188);
and U4654 (N_4654,N_3644,N_3931);
and U4655 (N_4655,N_3219,N_3647);
or U4656 (N_4656,N_3300,N_3299);
or U4657 (N_4657,N_3034,N_3967);
and U4658 (N_4658,N_3915,N_3984);
nand U4659 (N_4659,N_3317,N_3133);
and U4660 (N_4660,N_3318,N_3991);
nand U4661 (N_4661,N_3306,N_3924);
and U4662 (N_4662,N_3820,N_3176);
or U4663 (N_4663,N_3791,N_3211);
xor U4664 (N_4664,N_3737,N_3637);
or U4665 (N_4665,N_3772,N_3455);
or U4666 (N_4666,N_3010,N_3401);
nor U4667 (N_4667,N_3531,N_3316);
nand U4668 (N_4668,N_3154,N_3159);
nor U4669 (N_4669,N_3797,N_3434);
nand U4670 (N_4670,N_3019,N_3139);
nand U4671 (N_4671,N_3833,N_3979);
nand U4672 (N_4672,N_3347,N_3854);
nand U4673 (N_4673,N_3770,N_3839);
xnor U4674 (N_4674,N_3888,N_3202);
xor U4675 (N_4675,N_3704,N_3892);
nor U4676 (N_4676,N_3736,N_3328);
nor U4677 (N_4677,N_3997,N_3130);
and U4678 (N_4678,N_3639,N_3429);
and U4679 (N_4679,N_3220,N_3292);
and U4680 (N_4680,N_3091,N_3317);
nand U4681 (N_4681,N_3398,N_3818);
and U4682 (N_4682,N_3165,N_3728);
and U4683 (N_4683,N_3166,N_3574);
or U4684 (N_4684,N_3466,N_3119);
and U4685 (N_4685,N_3413,N_3280);
or U4686 (N_4686,N_3893,N_3129);
nor U4687 (N_4687,N_3555,N_3640);
nand U4688 (N_4688,N_3788,N_3535);
nor U4689 (N_4689,N_3246,N_3138);
nand U4690 (N_4690,N_3358,N_3165);
or U4691 (N_4691,N_3283,N_3003);
or U4692 (N_4692,N_3788,N_3429);
or U4693 (N_4693,N_3420,N_3508);
or U4694 (N_4694,N_3488,N_3257);
nand U4695 (N_4695,N_3124,N_3736);
nand U4696 (N_4696,N_3867,N_3528);
nor U4697 (N_4697,N_3971,N_3955);
nand U4698 (N_4698,N_3285,N_3476);
or U4699 (N_4699,N_3000,N_3414);
nand U4700 (N_4700,N_3258,N_3753);
or U4701 (N_4701,N_3911,N_3520);
or U4702 (N_4702,N_3236,N_3288);
or U4703 (N_4703,N_3013,N_3427);
and U4704 (N_4704,N_3214,N_3786);
xnor U4705 (N_4705,N_3296,N_3458);
nand U4706 (N_4706,N_3155,N_3865);
and U4707 (N_4707,N_3346,N_3953);
or U4708 (N_4708,N_3532,N_3579);
and U4709 (N_4709,N_3914,N_3615);
nand U4710 (N_4710,N_3391,N_3008);
or U4711 (N_4711,N_3589,N_3136);
nand U4712 (N_4712,N_3808,N_3670);
nor U4713 (N_4713,N_3448,N_3412);
nor U4714 (N_4714,N_3894,N_3908);
nand U4715 (N_4715,N_3805,N_3631);
or U4716 (N_4716,N_3376,N_3842);
or U4717 (N_4717,N_3433,N_3024);
nand U4718 (N_4718,N_3115,N_3083);
nor U4719 (N_4719,N_3098,N_3473);
nand U4720 (N_4720,N_3378,N_3881);
or U4721 (N_4721,N_3156,N_3692);
and U4722 (N_4722,N_3075,N_3760);
nand U4723 (N_4723,N_3716,N_3522);
nand U4724 (N_4724,N_3473,N_3419);
nor U4725 (N_4725,N_3102,N_3279);
and U4726 (N_4726,N_3447,N_3553);
nand U4727 (N_4727,N_3880,N_3515);
or U4728 (N_4728,N_3715,N_3926);
nor U4729 (N_4729,N_3701,N_3808);
and U4730 (N_4730,N_3079,N_3797);
nor U4731 (N_4731,N_3823,N_3789);
nor U4732 (N_4732,N_3448,N_3889);
nand U4733 (N_4733,N_3109,N_3500);
nor U4734 (N_4734,N_3932,N_3185);
nor U4735 (N_4735,N_3278,N_3192);
or U4736 (N_4736,N_3220,N_3831);
xnor U4737 (N_4737,N_3798,N_3780);
nor U4738 (N_4738,N_3003,N_3476);
and U4739 (N_4739,N_3523,N_3980);
and U4740 (N_4740,N_3218,N_3192);
nand U4741 (N_4741,N_3672,N_3985);
and U4742 (N_4742,N_3631,N_3543);
and U4743 (N_4743,N_3617,N_3470);
and U4744 (N_4744,N_3146,N_3653);
and U4745 (N_4745,N_3772,N_3892);
nor U4746 (N_4746,N_3174,N_3455);
or U4747 (N_4747,N_3785,N_3605);
nor U4748 (N_4748,N_3089,N_3599);
nand U4749 (N_4749,N_3184,N_3412);
nand U4750 (N_4750,N_3380,N_3970);
or U4751 (N_4751,N_3062,N_3606);
nand U4752 (N_4752,N_3324,N_3251);
or U4753 (N_4753,N_3628,N_3470);
nand U4754 (N_4754,N_3942,N_3316);
nor U4755 (N_4755,N_3909,N_3689);
xnor U4756 (N_4756,N_3349,N_3155);
and U4757 (N_4757,N_3880,N_3594);
nand U4758 (N_4758,N_3070,N_3551);
or U4759 (N_4759,N_3366,N_3657);
and U4760 (N_4760,N_3641,N_3292);
nand U4761 (N_4761,N_3159,N_3522);
nand U4762 (N_4762,N_3198,N_3767);
or U4763 (N_4763,N_3883,N_3235);
nor U4764 (N_4764,N_3562,N_3227);
and U4765 (N_4765,N_3592,N_3861);
nor U4766 (N_4766,N_3038,N_3773);
and U4767 (N_4767,N_3953,N_3126);
nand U4768 (N_4768,N_3819,N_3402);
nand U4769 (N_4769,N_3736,N_3413);
and U4770 (N_4770,N_3620,N_3433);
nand U4771 (N_4771,N_3952,N_3316);
nor U4772 (N_4772,N_3564,N_3662);
nand U4773 (N_4773,N_3443,N_3078);
nand U4774 (N_4774,N_3082,N_3206);
and U4775 (N_4775,N_3374,N_3385);
nor U4776 (N_4776,N_3192,N_3802);
nand U4777 (N_4777,N_3966,N_3006);
or U4778 (N_4778,N_3550,N_3862);
xnor U4779 (N_4779,N_3593,N_3534);
or U4780 (N_4780,N_3335,N_3953);
nand U4781 (N_4781,N_3539,N_3412);
nand U4782 (N_4782,N_3614,N_3158);
nor U4783 (N_4783,N_3141,N_3351);
nand U4784 (N_4784,N_3782,N_3767);
and U4785 (N_4785,N_3488,N_3715);
and U4786 (N_4786,N_3713,N_3738);
nor U4787 (N_4787,N_3192,N_3249);
and U4788 (N_4788,N_3336,N_3520);
nand U4789 (N_4789,N_3609,N_3064);
nand U4790 (N_4790,N_3501,N_3232);
nor U4791 (N_4791,N_3541,N_3929);
nor U4792 (N_4792,N_3691,N_3476);
nor U4793 (N_4793,N_3989,N_3637);
nor U4794 (N_4794,N_3569,N_3638);
and U4795 (N_4795,N_3231,N_3157);
nand U4796 (N_4796,N_3900,N_3650);
nand U4797 (N_4797,N_3725,N_3373);
nand U4798 (N_4798,N_3633,N_3538);
nand U4799 (N_4799,N_3897,N_3202);
or U4800 (N_4800,N_3778,N_3029);
or U4801 (N_4801,N_3786,N_3063);
and U4802 (N_4802,N_3751,N_3734);
nor U4803 (N_4803,N_3977,N_3062);
nor U4804 (N_4804,N_3959,N_3156);
and U4805 (N_4805,N_3206,N_3622);
nand U4806 (N_4806,N_3294,N_3038);
and U4807 (N_4807,N_3896,N_3420);
nor U4808 (N_4808,N_3845,N_3774);
xnor U4809 (N_4809,N_3655,N_3448);
and U4810 (N_4810,N_3562,N_3478);
and U4811 (N_4811,N_3511,N_3701);
nor U4812 (N_4812,N_3224,N_3785);
and U4813 (N_4813,N_3048,N_3050);
and U4814 (N_4814,N_3447,N_3259);
and U4815 (N_4815,N_3786,N_3231);
nor U4816 (N_4816,N_3479,N_3645);
and U4817 (N_4817,N_3949,N_3001);
nor U4818 (N_4818,N_3462,N_3879);
and U4819 (N_4819,N_3701,N_3235);
nand U4820 (N_4820,N_3731,N_3027);
nor U4821 (N_4821,N_3199,N_3439);
and U4822 (N_4822,N_3283,N_3482);
and U4823 (N_4823,N_3016,N_3396);
or U4824 (N_4824,N_3626,N_3027);
nand U4825 (N_4825,N_3883,N_3772);
and U4826 (N_4826,N_3113,N_3959);
and U4827 (N_4827,N_3782,N_3434);
nor U4828 (N_4828,N_3744,N_3168);
nand U4829 (N_4829,N_3616,N_3808);
xnor U4830 (N_4830,N_3360,N_3109);
nor U4831 (N_4831,N_3510,N_3307);
nand U4832 (N_4832,N_3578,N_3221);
or U4833 (N_4833,N_3320,N_3776);
nand U4834 (N_4834,N_3768,N_3421);
and U4835 (N_4835,N_3804,N_3534);
nor U4836 (N_4836,N_3821,N_3580);
nand U4837 (N_4837,N_3519,N_3347);
nand U4838 (N_4838,N_3249,N_3931);
nor U4839 (N_4839,N_3673,N_3125);
or U4840 (N_4840,N_3776,N_3463);
nor U4841 (N_4841,N_3249,N_3531);
nand U4842 (N_4842,N_3275,N_3170);
nor U4843 (N_4843,N_3951,N_3718);
xor U4844 (N_4844,N_3318,N_3989);
nor U4845 (N_4845,N_3016,N_3390);
nor U4846 (N_4846,N_3435,N_3213);
nor U4847 (N_4847,N_3416,N_3417);
and U4848 (N_4848,N_3555,N_3175);
nand U4849 (N_4849,N_3512,N_3797);
or U4850 (N_4850,N_3224,N_3570);
nor U4851 (N_4851,N_3219,N_3375);
nand U4852 (N_4852,N_3002,N_3282);
and U4853 (N_4853,N_3716,N_3398);
nor U4854 (N_4854,N_3607,N_3774);
or U4855 (N_4855,N_3988,N_3151);
and U4856 (N_4856,N_3666,N_3567);
or U4857 (N_4857,N_3886,N_3832);
or U4858 (N_4858,N_3335,N_3092);
nor U4859 (N_4859,N_3349,N_3884);
or U4860 (N_4860,N_3290,N_3848);
nor U4861 (N_4861,N_3983,N_3651);
or U4862 (N_4862,N_3496,N_3887);
or U4863 (N_4863,N_3425,N_3515);
nand U4864 (N_4864,N_3903,N_3793);
nor U4865 (N_4865,N_3898,N_3231);
and U4866 (N_4866,N_3842,N_3854);
nand U4867 (N_4867,N_3412,N_3485);
or U4868 (N_4868,N_3786,N_3953);
or U4869 (N_4869,N_3842,N_3530);
nor U4870 (N_4870,N_3048,N_3460);
nor U4871 (N_4871,N_3599,N_3618);
and U4872 (N_4872,N_3303,N_3784);
nor U4873 (N_4873,N_3476,N_3833);
xor U4874 (N_4874,N_3287,N_3419);
or U4875 (N_4875,N_3074,N_3342);
and U4876 (N_4876,N_3215,N_3453);
nand U4877 (N_4877,N_3071,N_3698);
nand U4878 (N_4878,N_3630,N_3502);
nor U4879 (N_4879,N_3012,N_3736);
nor U4880 (N_4880,N_3971,N_3574);
and U4881 (N_4881,N_3163,N_3208);
nand U4882 (N_4882,N_3839,N_3026);
nor U4883 (N_4883,N_3106,N_3095);
nor U4884 (N_4884,N_3529,N_3321);
and U4885 (N_4885,N_3623,N_3369);
and U4886 (N_4886,N_3680,N_3084);
nand U4887 (N_4887,N_3688,N_3547);
and U4888 (N_4888,N_3370,N_3527);
and U4889 (N_4889,N_3050,N_3759);
nand U4890 (N_4890,N_3143,N_3372);
nand U4891 (N_4891,N_3825,N_3731);
nor U4892 (N_4892,N_3529,N_3010);
nand U4893 (N_4893,N_3301,N_3966);
and U4894 (N_4894,N_3521,N_3655);
nand U4895 (N_4895,N_3689,N_3355);
nand U4896 (N_4896,N_3101,N_3935);
and U4897 (N_4897,N_3144,N_3938);
and U4898 (N_4898,N_3474,N_3775);
nor U4899 (N_4899,N_3773,N_3368);
nand U4900 (N_4900,N_3612,N_3421);
and U4901 (N_4901,N_3943,N_3130);
or U4902 (N_4902,N_3836,N_3295);
nor U4903 (N_4903,N_3281,N_3423);
nand U4904 (N_4904,N_3273,N_3676);
or U4905 (N_4905,N_3802,N_3293);
nand U4906 (N_4906,N_3904,N_3175);
nor U4907 (N_4907,N_3046,N_3414);
or U4908 (N_4908,N_3884,N_3371);
nor U4909 (N_4909,N_3403,N_3967);
and U4910 (N_4910,N_3745,N_3864);
and U4911 (N_4911,N_3109,N_3690);
and U4912 (N_4912,N_3815,N_3162);
or U4913 (N_4913,N_3032,N_3719);
or U4914 (N_4914,N_3568,N_3008);
nand U4915 (N_4915,N_3645,N_3996);
and U4916 (N_4916,N_3294,N_3836);
nor U4917 (N_4917,N_3428,N_3683);
nand U4918 (N_4918,N_3888,N_3763);
nand U4919 (N_4919,N_3037,N_3245);
nand U4920 (N_4920,N_3327,N_3502);
or U4921 (N_4921,N_3550,N_3139);
nand U4922 (N_4922,N_3435,N_3307);
or U4923 (N_4923,N_3954,N_3745);
and U4924 (N_4924,N_3951,N_3545);
nor U4925 (N_4925,N_3386,N_3177);
nor U4926 (N_4926,N_3415,N_3021);
or U4927 (N_4927,N_3892,N_3282);
and U4928 (N_4928,N_3688,N_3342);
nor U4929 (N_4929,N_3412,N_3254);
or U4930 (N_4930,N_3407,N_3200);
and U4931 (N_4931,N_3277,N_3253);
or U4932 (N_4932,N_3004,N_3297);
or U4933 (N_4933,N_3925,N_3269);
nor U4934 (N_4934,N_3427,N_3151);
nor U4935 (N_4935,N_3481,N_3971);
nor U4936 (N_4936,N_3421,N_3486);
nand U4937 (N_4937,N_3255,N_3519);
or U4938 (N_4938,N_3099,N_3124);
and U4939 (N_4939,N_3652,N_3439);
nand U4940 (N_4940,N_3592,N_3340);
or U4941 (N_4941,N_3788,N_3113);
or U4942 (N_4942,N_3235,N_3033);
and U4943 (N_4943,N_3601,N_3954);
and U4944 (N_4944,N_3368,N_3529);
nor U4945 (N_4945,N_3847,N_3786);
nand U4946 (N_4946,N_3590,N_3358);
nand U4947 (N_4947,N_3656,N_3186);
nand U4948 (N_4948,N_3685,N_3513);
and U4949 (N_4949,N_3400,N_3707);
and U4950 (N_4950,N_3717,N_3094);
and U4951 (N_4951,N_3362,N_3960);
nand U4952 (N_4952,N_3936,N_3206);
and U4953 (N_4953,N_3926,N_3598);
and U4954 (N_4954,N_3678,N_3888);
xnor U4955 (N_4955,N_3303,N_3586);
and U4956 (N_4956,N_3361,N_3893);
nor U4957 (N_4957,N_3215,N_3563);
or U4958 (N_4958,N_3190,N_3301);
nor U4959 (N_4959,N_3316,N_3686);
and U4960 (N_4960,N_3501,N_3312);
nor U4961 (N_4961,N_3180,N_3286);
nor U4962 (N_4962,N_3162,N_3649);
nand U4963 (N_4963,N_3945,N_3171);
nand U4964 (N_4964,N_3028,N_3121);
or U4965 (N_4965,N_3480,N_3242);
nor U4966 (N_4966,N_3764,N_3038);
and U4967 (N_4967,N_3869,N_3767);
and U4968 (N_4968,N_3115,N_3354);
or U4969 (N_4969,N_3425,N_3879);
nand U4970 (N_4970,N_3704,N_3151);
or U4971 (N_4971,N_3595,N_3989);
or U4972 (N_4972,N_3686,N_3226);
and U4973 (N_4973,N_3824,N_3025);
and U4974 (N_4974,N_3098,N_3898);
and U4975 (N_4975,N_3808,N_3813);
nor U4976 (N_4976,N_3318,N_3163);
or U4977 (N_4977,N_3666,N_3406);
xnor U4978 (N_4978,N_3291,N_3168);
and U4979 (N_4979,N_3282,N_3218);
and U4980 (N_4980,N_3863,N_3194);
nor U4981 (N_4981,N_3546,N_3894);
nor U4982 (N_4982,N_3455,N_3783);
nand U4983 (N_4983,N_3470,N_3859);
and U4984 (N_4984,N_3534,N_3438);
nand U4985 (N_4985,N_3816,N_3927);
nand U4986 (N_4986,N_3224,N_3954);
or U4987 (N_4987,N_3861,N_3044);
nand U4988 (N_4988,N_3267,N_3718);
nor U4989 (N_4989,N_3220,N_3624);
or U4990 (N_4990,N_3746,N_3317);
nand U4991 (N_4991,N_3488,N_3461);
nand U4992 (N_4992,N_3968,N_3782);
or U4993 (N_4993,N_3694,N_3121);
nand U4994 (N_4994,N_3042,N_3679);
nor U4995 (N_4995,N_3402,N_3784);
nor U4996 (N_4996,N_3514,N_3020);
nor U4997 (N_4997,N_3104,N_3978);
or U4998 (N_4998,N_3451,N_3043);
and U4999 (N_4999,N_3575,N_3152);
and UO_0 (O_0,N_4671,N_4319);
or UO_1 (O_1,N_4793,N_4920);
or UO_2 (O_2,N_4923,N_4395);
or UO_3 (O_3,N_4289,N_4107);
or UO_4 (O_4,N_4742,N_4729);
nand UO_5 (O_5,N_4869,N_4199);
xor UO_6 (O_6,N_4785,N_4104);
or UO_7 (O_7,N_4495,N_4596);
and UO_8 (O_8,N_4875,N_4816);
and UO_9 (O_9,N_4953,N_4050);
xor UO_10 (O_10,N_4633,N_4681);
nor UO_11 (O_11,N_4666,N_4523);
nor UO_12 (O_12,N_4113,N_4743);
nor UO_13 (O_13,N_4763,N_4685);
or UO_14 (O_14,N_4547,N_4583);
nor UO_15 (O_15,N_4739,N_4692);
nor UO_16 (O_16,N_4250,N_4718);
nor UO_17 (O_17,N_4654,N_4570);
nor UO_18 (O_18,N_4323,N_4995);
nor UO_19 (O_19,N_4391,N_4438);
or UO_20 (O_20,N_4860,N_4463);
xnor UO_21 (O_21,N_4094,N_4112);
or UO_22 (O_22,N_4118,N_4960);
nor UO_23 (O_23,N_4440,N_4795);
or UO_24 (O_24,N_4769,N_4908);
nor UO_25 (O_25,N_4624,N_4322);
nor UO_26 (O_26,N_4864,N_4677);
nand UO_27 (O_27,N_4032,N_4011);
and UO_28 (O_28,N_4569,N_4880);
nand UO_29 (O_29,N_4727,N_4884);
and UO_30 (O_30,N_4997,N_4179);
nor UO_31 (O_31,N_4225,N_4932);
or UO_32 (O_32,N_4499,N_4702);
nor UO_33 (O_33,N_4367,N_4068);
and UO_34 (O_34,N_4600,N_4881);
nand UO_35 (O_35,N_4934,N_4837);
and UO_36 (O_36,N_4160,N_4886);
or UO_37 (O_37,N_4196,N_4525);
and UO_38 (O_38,N_4990,N_4811);
and UO_39 (O_39,N_4812,N_4784);
xnor UO_40 (O_40,N_4268,N_4445);
or UO_41 (O_41,N_4360,N_4972);
or UO_42 (O_42,N_4758,N_4650);
nand UO_43 (O_43,N_4631,N_4406);
or UO_44 (O_44,N_4296,N_4500);
and UO_45 (O_45,N_4899,N_4086);
nand UO_46 (O_46,N_4204,N_4925);
nor UO_47 (O_47,N_4079,N_4771);
nor UO_48 (O_48,N_4386,N_4018);
nor UO_49 (O_49,N_4961,N_4124);
or UO_50 (O_50,N_4272,N_4511);
and UO_51 (O_51,N_4081,N_4189);
nand UO_52 (O_52,N_4279,N_4798);
and UO_53 (O_53,N_4248,N_4023);
nor UO_54 (O_54,N_4400,N_4016);
nand UO_55 (O_55,N_4276,N_4530);
nor UO_56 (O_56,N_4167,N_4158);
nand UO_57 (O_57,N_4721,N_4355);
and UO_58 (O_58,N_4574,N_4859);
and UO_59 (O_59,N_4197,N_4797);
nor UO_60 (O_60,N_4384,N_4558);
or UO_61 (O_61,N_4205,N_4143);
or UO_62 (O_62,N_4168,N_4903);
or UO_63 (O_63,N_4682,N_4794);
and UO_64 (O_64,N_4683,N_4416);
nand UO_65 (O_65,N_4078,N_4116);
nand UO_66 (O_66,N_4031,N_4173);
nand UO_67 (O_67,N_4183,N_4576);
or UO_68 (O_68,N_4064,N_4477);
nor UO_69 (O_69,N_4099,N_4985);
and UO_70 (O_70,N_4640,N_4310);
or UO_71 (O_71,N_4620,N_4324);
and UO_72 (O_72,N_4806,N_4441);
nor UO_73 (O_73,N_4870,N_4084);
nand UO_74 (O_74,N_4447,N_4106);
nand UO_75 (O_75,N_4835,N_4820);
and UO_76 (O_76,N_4460,N_4177);
and UO_77 (O_77,N_4539,N_4220);
nor UO_78 (O_78,N_4898,N_4212);
nand UO_79 (O_79,N_4863,N_4637);
nand UO_80 (O_80,N_4470,N_4579);
and UO_81 (O_81,N_4625,N_4365);
or UO_82 (O_82,N_4745,N_4328);
nand UO_83 (O_83,N_4442,N_4255);
nor UO_84 (O_84,N_4096,N_4832);
and UO_85 (O_85,N_4595,N_4396);
nand UO_86 (O_86,N_4809,N_4194);
and UO_87 (O_87,N_4644,N_4782);
or UO_88 (O_88,N_4227,N_4534);
and UO_89 (O_89,N_4805,N_4280);
and UO_90 (O_90,N_4978,N_4484);
nand UO_91 (O_91,N_4325,N_4675);
and UO_92 (O_92,N_4175,N_4370);
and UO_93 (O_93,N_4580,N_4592);
or UO_94 (O_94,N_4235,N_4374);
and UO_95 (O_95,N_4402,N_4730);
xnor UO_96 (O_96,N_4012,N_4819);
and UO_97 (O_97,N_4623,N_4895);
nor UO_98 (O_98,N_4706,N_4329);
nand UO_99 (O_99,N_4561,N_4088);
or UO_100 (O_100,N_4418,N_4823);
nor UO_101 (O_101,N_4469,N_4824);
or UO_102 (O_102,N_4028,N_4709);
and UO_103 (O_103,N_4425,N_4332);
nand UO_104 (O_104,N_4215,N_4493);
and UO_105 (O_105,N_4528,N_4836);
nand UO_106 (O_106,N_4853,N_4548);
nand UO_107 (O_107,N_4145,N_4055);
or UO_108 (O_108,N_4343,N_4213);
nor UO_109 (O_109,N_4737,N_4956);
nand UO_110 (O_110,N_4589,N_4750);
nand UO_111 (O_111,N_4919,N_4751);
or UO_112 (O_112,N_4756,N_4258);
nor UO_113 (O_113,N_4532,N_4764);
nor UO_114 (O_114,N_4065,N_4556);
and UO_115 (O_115,N_4480,N_4348);
nand UO_116 (O_116,N_4606,N_4059);
or UO_117 (O_117,N_4133,N_4999);
nor UO_118 (O_118,N_4292,N_4566);
and UO_119 (O_119,N_4083,N_4185);
nand UO_120 (O_120,N_4070,N_4672);
and UO_121 (O_121,N_4904,N_4544);
or UO_122 (O_122,N_4444,N_4714);
nor UO_123 (O_123,N_4981,N_4388);
nand UO_124 (O_124,N_4260,N_4135);
and UO_125 (O_125,N_4987,N_4221);
nor UO_126 (O_126,N_4253,N_4399);
nand UO_127 (O_127,N_4555,N_4776);
and UO_128 (O_128,N_4728,N_4263);
or UO_129 (O_129,N_4788,N_4379);
and UO_130 (O_130,N_4153,N_4567);
nor UO_131 (O_131,N_4652,N_4791);
nand UO_132 (O_132,N_4696,N_4646);
nor UO_133 (O_133,N_4757,N_4636);
nand UO_134 (O_134,N_4915,N_4546);
and UO_135 (O_135,N_4607,N_4264);
and UO_136 (O_136,N_4103,N_4927);
and UO_137 (O_137,N_4005,N_4377);
or UO_138 (O_138,N_4410,N_4862);
or UO_139 (O_139,N_4778,N_4186);
and UO_140 (O_140,N_4694,N_4344);
or UO_141 (O_141,N_4282,N_4598);
xor UO_142 (O_142,N_4019,N_4342);
nor UO_143 (O_143,N_4542,N_4170);
nand UO_144 (O_144,N_4269,N_4412);
nand UO_145 (O_145,N_4049,N_4270);
and UO_146 (O_146,N_4452,N_4614);
and UO_147 (O_147,N_4354,N_4218);
nor UO_148 (O_148,N_4643,N_4715);
or UO_149 (O_149,N_4419,N_4732);
and UO_150 (O_150,N_4467,N_4735);
or UO_151 (O_151,N_4662,N_4320);
or UO_152 (O_152,N_4491,N_4826);
and UO_153 (O_153,N_4717,N_4004);
nand UO_154 (O_154,N_4628,N_4125);
or UO_155 (O_155,N_4922,N_4108);
nand UO_156 (O_156,N_4973,N_4290);
nand UO_157 (O_157,N_4146,N_4102);
and UO_158 (O_158,N_4283,N_4411);
or UO_159 (O_159,N_4959,N_4335);
nand UO_160 (O_160,N_4473,N_4844);
or UO_161 (O_161,N_4131,N_4907);
or UO_162 (O_162,N_4201,N_4286);
or UO_163 (O_163,N_4381,N_4306);
and UO_164 (O_164,N_4257,N_4132);
nor UO_165 (O_165,N_4955,N_4334);
nand UO_166 (O_166,N_4349,N_4510);
xor UO_167 (O_167,N_4439,N_4963);
nand UO_168 (O_168,N_4725,N_4462);
xor UO_169 (O_169,N_4856,N_4380);
and UO_170 (O_170,N_4450,N_4026);
or UO_171 (O_171,N_4298,N_4184);
and UO_172 (O_172,N_4770,N_4436);
xor UO_173 (O_173,N_4098,N_4817);
nand UO_174 (O_174,N_4243,N_4670);
nand UO_175 (O_175,N_4256,N_4188);
nand UO_176 (O_176,N_4573,N_4383);
or UO_177 (O_177,N_4376,N_4033);
nand UO_178 (O_178,N_4851,N_4315);
nor UO_179 (O_179,N_4497,N_4581);
or UO_180 (O_180,N_4610,N_4378);
and UO_181 (O_181,N_4341,N_4195);
and UO_182 (O_182,N_4488,N_4203);
nor UO_183 (O_183,N_4317,N_4803);
or UO_184 (O_184,N_4456,N_4868);
xnor UO_185 (O_185,N_4695,N_4490);
nor UO_186 (O_186,N_4597,N_4362);
and UO_187 (O_187,N_4615,N_4137);
nor UO_188 (O_188,N_4707,N_4274);
nor UO_189 (O_189,N_4375,N_4267);
nor UO_190 (O_190,N_4455,N_4871);
or UO_191 (O_191,N_4039,N_4941);
nand UO_192 (O_192,N_4829,N_4846);
and UO_193 (O_193,N_4563,N_4437);
nand UO_194 (O_194,N_4746,N_4611);
and UO_195 (O_195,N_4691,N_4842);
nor UO_196 (O_196,N_4855,N_4529);
xor UO_197 (O_197,N_4236,N_4048);
nor UO_198 (O_198,N_4085,N_4568);
and UO_199 (O_199,N_4513,N_4924);
nor UO_200 (O_200,N_4407,N_4427);
xnor UO_201 (O_201,N_4277,N_4524);
nor UO_202 (O_202,N_4123,N_4674);
nor UO_203 (O_203,N_4850,N_4629);
nand UO_204 (O_204,N_4466,N_4664);
or UO_205 (O_205,N_4711,N_4009);
and UO_206 (O_206,N_4635,N_4434);
or UO_207 (O_207,N_4936,N_4752);
and UO_208 (O_208,N_4479,N_4134);
or UO_209 (O_209,N_4509,N_4551);
or UO_210 (O_210,N_4553,N_4810);
or UO_211 (O_211,N_4024,N_4653);
nand UO_212 (O_212,N_4001,N_4219);
nand UO_213 (O_213,N_4474,N_4559);
and UO_214 (O_214,N_4390,N_4288);
nand UO_215 (O_215,N_4678,N_4578);
nand UO_216 (O_216,N_4082,N_4190);
nand UO_217 (O_217,N_4408,N_4266);
nand UO_218 (O_218,N_4147,N_4430);
and UO_219 (O_219,N_4359,N_4216);
nand UO_220 (O_220,N_4062,N_4814);
nand UO_221 (O_221,N_4517,N_4127);
or UO_222 (O_222,N_4373,N_4804);
nor UO_223 (O_223,N_4295,N_4057);
nand UO_224 (O_224,N_4502,N_4779);
or UO_225 (O_225,N_4389,N_4545);
nand UO_226 (O_226,N_4991,N_4605);
nand UO_227 (O_227,N_4159,N_4854);
nand UO_228 (O_228,N_4882,N_4223);
nand UO_229 (O_229,N_4661,N_4187);
or UO_230 (O_230,N_4777,N_4461);
or UO_231 (O_231,N_4647,N_4166);
nand UO_232 (O_232,N_4965,N_4364);
xnor UO_233 (O_233,N_4465,N_4345);
and UO_234 (O_234,N_4822,N_4852);
or UO_235 (O_235,N_4003,N_4565);
nor UO_236 (O_236,N_4040,N_4831);
or UO_237 (O_237,N_4808,N_4246);
or UO_238 (O_238,N_4487,N_4202);
or UO_239 (O_239,N_4571,N_4352);
or UO_240 (O_240,N_4152,N_4948);
nor UO_241 (O_241,N_4818,N_4686);
and UO_242 (O_242,N_4989,N_4849);
nor UO_243 (O_243,N_4262,N_4535);
nand UO_244 (O_244,N_4587,N_4519);
and UO_245 (O_245,N_4156,N_4287);
nand UO_246 (O_246,N_4021,N_4312);
and UO_247 (O_247,N_4657,N_4585);
and UO_248 (O_248,N_4608,N_4697);
nand UO_249 (O_249,N_4802,N_4748);
nand UO_250 (O_250,N_4526,N_4609);
or UO_251 (O_251,N_4140,N_4921);
or UO_252 (O_252,N_4414,N_4020);
nor UO_253 (O_253,N_4014,N_4792);
nor UO_254 (O_254,N_4401,N_4387);
nand UO_255 (O_255,N_4731,N_4993);
or UO_256 (O_256,N_4353,N_4942);
or UO_257 (O_257,N_4845,N_4540);
or UO_258 (O_258,N_4006,N_4035);
and UO_259 (O_259,N_4954,N_4431);
nand UO_260 (O_260,N_4182,N_4966);
nor UO_261 (O_261,N_4045,N_4138);
nand UO_262 (O_262,N_4541,N_4155);
or UO_263 (O_263,N_4626,N_4673);
and UO_264 (O_264,N_4192,N_4962);
and UO_265 (O_265,N_4949,N_4889);
nor UO_266 (O_266,N_4929,N_4211);
or UO_267 (O_267,N_4351,N_4668);
nor UO_268 (O_268,N_4872,N_4952);
or UO_269 (O_269,N_4453,N_4733);
and UO_270 (O_270,N_4928,N_4760);
nor UO_271 (O_271,N_4483,N_4476);
nor UO_272 (O_272,N_4887,N_4612);
or UO_273 (O_273,N_4178,N_4834);
nand UO_274 (O_274,N_4828,N_4913);
nor UO_275 (O_275,N_4753,N_4848);
nand UO_276 (O_276,N_4301,N_4141);
nand UO_277 (O_277,N_4744,N_4238);
or UO_278 (O_278,N_4428,N_4122);
or UO_279 (O_279,N_4911,N_4117);
nand UO_280 (O_280,N_4554,N_4841);
nor UO_281 (O_281,N_4121,N_4361);
nand UO_282 (O_282,N_4549,N_4054);
or UO_283 (O_283,N_4052,N_4577);
nor UO_284 (O_284,N_4939,N_4339);
nand UO_285 (O_285,N_4200,N_4126);
or UO_286 (O_286,N_4056,N_4066);
or UO_287 (O_287,N_4457,N_4734);
nor UO_288 (O_288,N_4813,N_4067);
nor UO_289 (O_289,N_4226,N_4594);
and UO_290 (O_290,N_4092,N_4508);
nor UO_291 (O_291,N_4773,N_4232);
nor UO_292 (O_292,N_4689,N_4244);
and UO_293 (O_293,N_4910,N_4240);
nor UO_294 (O_294,N_4632,N_4642);
and UO_295 (O_295,N_4494,N_4129);
and UO_296 (O_296,N_4356,N_4930);
or UO_297 (O_297,N_4172,N_4634);
nand UO_298 (O_298,N_4759,N_4552);
nor UO_299 (O_299,N_4489,N_4789);
and UO_300 (O_300,N_4582,N_4766);
or UO_301 (O_301,N_4180,N_4007);
and UO_302 (O_302,N_4520,N_4327);
or UO_303 (O_303,N_4368,N_4307);
and UO_304 (O_304,N_4982,N_4485);
or UO_305 (O_305,N_4747,N_4900);
nand UO_306 (O_306,N_4091,N_4041);
xnor UO_307 (O_307,N_4575,N_4537);
xor UO_308 (O_308,N_4933,N_4665);
or UO_309 (O_309,N_4780,N_4712);
nor UO_310 (O_310,N_4648,N_4772);
nand UO_311 (O_311,N_4230,N_4053);
and UO_312 (O_312,N_4658,N_4036);
nor UO_313 (O_313,N_4247,N_4504);
nor UO_314 (O_314,N_4382,N_4060);
and UO_315 (O_315,N_4423,N_4627);
nor UO_316 (O_316,N_4839,N_4420);
nor UO_317 (O_317,N_4432,N_4917);
nor UO_318 (O_318,N_4801,N_4284);
nand UO_319 (O_319,N_4522,N_4840);
nand UO_320 (O_320,N_4821,N_4892);
or UO_321 (O_321,N_4090,N_4481);
nand UO_322 (O_322,N_4720,N_4120);
nand UO_323 (O_323,N_4278,N_4741);
nor UO_324 (O_324,N_4755,N_4075);
nor UO_325 (O_325,N_4890,N_4660);
and UO_326 (O_326,N_4017,N_4825);
nor UO_327 (O_327,N_4224,N_4478);
or UO_328 (O_328,N_4687,N_4800);
and UO_329 (O_329,N_4340,N_4710);
nand UO_330 (O_330,N_4861,N_4655);
or UO_331 (O_331,N_4969,N_4506);
and UO_332 (O_332,N_4701,N_4472);
xnor UO_333 (O_333,N_4193,N_4905);
and UO_334 (O_334,N_4372,N_4252);
and UO_335 (O_335,N_4590,N_4151);
nor UO_336 (O_336,N_4433,N_4207);
or UO_337 (O_337,N_4562,N_4983);
nor UO_338 (O_338,N_4429,N_4231);
nor UO_339 (O_339,N_4946,N_4937);
and UO_340 (O_340,N_4459,N_4943);
or UO_341 (O_341,N_4303,N_4074);
nor UO_342 (O_342,N_4774,N_4259);
or UO_343 (O_343,N_4297,N_4971);
or UO_344 (O_344,N_4063,N_4191);
nand UO_345 (O_345,N_4069,N_4149);
or UO_346 (O_346,N_4891,N_4938);
and UO_347 (O_347,N_4331,N_4699);
nand UO_348 (O_348,N_4815,N_4154);
nand UO_349 (O_349,N_4030,N_4350);
nand UO_350 (O_350,N_4667,N_4783);
nand UO_351 (O_351,N_4931,N_4726);
nor UO_352 (O_352,N_4304,N_4669);
and UO_353 (O_353,N_4454,N_4398);
and UO_354 (O_354,N_4616,N_4369);
nor UO_355 (O_355,N_4790,N_4700);
xor UO_356 (O_356,N_4073,N_4680);
or UO_357 (O_357,N_4176,N_4271);
nor UO_358 (O_358,N_4042,N_4409);
and UO_359 (O_359,N_4393,N_4874);
nor UO_360 (O_360,N_4603,N_4516);
nand UO_361 (O_361,N_4945,N_4162);
xnor UO_362 (O_362,N_4940,N_4181);
and UO_363 (O_363,N_4613,N_4237);
and UO_364 (O_364,N_4977,N_4765);
and UO_365 (O_365,N_4617,N_4443);
nand UO_366 (O_366,N_4013,N_4639);
nor UO_367 (O_367,N_4164,N_4171);
nand UO_368 (O_368,N_4451,N_4857);
or UO_369 (O_369,N_4165,N_4958);
or UO_370 (O_370,N_4208,N_4724);
or UO_371 (O_371,N_4169,N_4101);
or UO_372 (O_372,N_4984,N_4486);
nand UO_373 (O_373,N_4308,N_4405);
or UO_374 (O_374,N_4338,N_4796);
and UO_375 (O_375,N_4471,N_4787);
nor UO_376 (O_376,N_4139,N_4584);
nor UO_377 (O_377,N_4630,N_4110);
and UO_378 (O_378,N_4265,N_4641);
or UO_379 (O_379,N_4501,N_4034);
or UO_380 (O_380,N_4698,N_4496);
nand UO_381 (O_381,N_4002,N_4847);
nor UO_382 (O_382,N_4119,N_4944);
nor UO_383 (O_383,N_4521,N_4302);
nor UO_384 (O_384,N_4309,N_4560);
and UO_385 (O_385,N_4543,N_4649);
nand UO_386 (O_386,N_4449,N_4008);
and UO_387 (O_387,N_4622,N_4229);
nand UO_388 (O_388,N_4051,N_4588);
nand UO_389 (O_389,N_4217,N_4676);
and UO_390 (O_390,N_4507,N_4980);
and UO_391 (O_391,N_4736,N_4448);
or UO_392 (O_392,N_4417,N_4704);
and UO_393 (O_393,N_4762,N_4533);
xor UO_394 (O_394,N_4046,N_4027);
nand UO_395 (O_395,N_4878,N_4951);
nand UO_396 (O_396,N_4291,N_4975);
or UO_397 (O_397,N_4080,N_4705);
nand UO_398 (O_398,N_4740,N_4865);
nand UO_399 (O_399,N_4174,N_4888);
and UO_400 (O_400,N_4058,N_4906);
nor UO_401 (O_401,N_4115,N_4464);
and UO_402 (O_402,N_4974,N_4209);
and UO_403 (O_403,N_4210,N_4397);
nand UO_404 (O_404,N_4093,N_4404);
nor UO_405 (O_405,N_4071,N_4572);
or UO_406 (O_406,N_4087,N_4458);
or UO_407 (O_407,N_4557,N_4206);
nand UO_408 (O_408,N_4619,N_4371);
or UO_409 (O_409,N_4316,N_4300);
nand UO_410 (O_410,N_4249,N_4294);
xor UO_411 (O_411,N_4621,N_4314);
and UO_412 (O_412,N_4144,N_4077);
nand UO_413 (O_413,N_4593,N_4475);
or UO_414 (O_414,N_4843,N_4254);
and UO_415 (O_415,N_4114,N_4498);
or UO_416 (O_416,N_4337,N_4047);
and UO_417 (O_417,N_4688,N_4894);
nand UO_418 (O_418,N_4311,N_4967);
and UO_419 (O_419,N_4468,N_4357);
or UO_420 (O_420,N_4708,N_4514);
or UO_421 (O_421,N_4947,N_4893);
and UO_422 (O_422,N_4935,N_4347);
nand UO_423 (O_423,N_4128,N_4044);
nand UO_424 (O_424,N_4749,N_4363);
nor UO_425 (O_425,N_4879,N_4330);
xor UO_426 (O_426,N_4111,N_4723);
nor UO_427 (O_427,N_4105,N_4781);
and UO_428 (O_428,N_4392,N_4979);
or UO_429 (O_429,N_4305,N_4902);
nand UO_430 (O_430,N_4994,N_4503);
nand UO_431 (O_431,N_4299,N_4768);
or UO_432 (O_432,N_4222,N_4022);
nor UO_433 (O_433,N_4964,N_4318);
or UO_434 (O_434,N_4645,N_4358);
and UO_435 (O_435,N_4713,N_4015);
nor UO_436 (O_436,N_4988,N_4738);
nand UO_437 (O_437,N_4719,N_4415);
nand UO_438 (O_438,N_4245,N_4394);
or UO_439 (O_439,N_4157,N_4076);
nor UO_440 (O_440,N_4422,N_4916);
nand UO_441 (O_441,N_4421,N_4109);
or UO_442 (O_442,N_4061,N_4986);
nand UO_443 (O_443,N_4482,N_4827);
nor UO_444 (O_444,N_4638,N_4161);
and UO_445 (O_445,N_4333,N_4536);
or UO_446 (O_446,N_4866,N_4996);
and UO_447 (O_447,N_4550,N_4914);
nand UO_448 (O_448,N_4873,N_4950);
nor UO_449 (O_449,N_4926,N_4130);
and UO_450 (O_450,N_4693,N_4876);
xor UO_451 (O_451,N_4604,N_4761);
and UO_452 (O_452,N_4807,N_4492);
nand UO_453 (O_453,N_4601,N_4043);
nor UO_454 (O_454,N_4656,N_4599);
nor UO_455 (O_455,N_4992,N_4918);
nor UO_456 (O_456,N_4512,N_4403);
nand UO_457 (O_457,N_4591,N_4029);
and UO_458 (O_458,N_4957,N_4321);
nor UO_459 (O_459,N_4242,N_4722);
nor UO_460 (O_460,N_4912,N_4366);
nand UO_461 (O_461,N_4163,N_4010);
nand UO_462 (O_462,N_4901,N_4037);
nand UO_463 (O_463,N_4786,N_4602);
nor UO_464 (O_464,N_4518,N_4976);
or UO_465 (O_465,N_4703,N_4767);
or UO_466 (O_466,N_4150,N_4233);
nand UO_467 (O_467,N_4885,N_4775);
nor UO_468 (O_468,N_4426,N_4136);
nor UO_469 (O_469,N_4293,N_4659);
nor UO_470 (O_470,N_4000,N_4089);
or UO_471 (O_471,N_4097,N_4385);
nor UO_472 (O_472,N_4538,N_4285);
or UO_473 (O_473,N_4833,N_4446);
and UO_474 (O_474,N_4413,N_4716);
or UO_475 (O_475,N_4830,N_4663);
nor UO_476 (O_476,N_4228,N_4586);
and UO_477 (O_477,N_4867,N_4313);
or UO_478 (O_478,N_4038,N_4838);
or UO_479 (O_479,N_4998,N_4326);
or UO_480 (O_480,N_4241,N_4025);
nand UO_481 (O_481,N_4346,N_4281);
or UO_482 (O_482,N_4148,N_4435);
and UO_483 (O_483,N_4100,N_4897);
nand UO_484 (O_484,N_4234,N_4858);
and UO_485 (O_485,N_4754,N_4690);
nor UO_486 (O_486,N_4877,N_4531);
or UO_487 (O_487,N_4198,N_4251);
and UO_488 (O_488,N_4142,N_4095);
or UO_489 (O_489,N_4336,N_4505);
nand UO_490 (O_490,N_4651,N_4679);
and UO_491 (O_491,N_4275,N_4883);
or UO_492 (O_492,N_4515,N_4618);
and UO_493 (O_493,N_4214,N_4072);
nand UO_494 (O_494,N_4968,N_4239);
nand UO_495 (O_495,N_4684,N_4527);
and UO_496 (O_496,N_4896,N_4799);
nand UO_497 (O_497,N_4970,N_4261);
and UO_498 (O_498,N_4909,N_4273);
and UO_499 (O_499,N_4564,N_4424);
nand UO_500 (O_500,N_4454,N_4261);
nor UO_501 (O_501,N_4640,N_4419);
nor UO_502 (O_502,N_4541,N_4322);
nor UO_503 (O_503,N_4304,N_4240);
and UO_504 (O_504,N_4139,N_4187);
or UO_505 (O_505,N_4792,N_4046);
and UO_506 (O_506,N_4880,N_4540);
or UO_507 (O_507,N_4171,N_4945);
and UO_508 (O_508,N_4581,N_4018);
nor UO_509 (O_509,N_4740,N_4096);
nand UO_510 (O_510,N_4121,N_4417);
xnor UO_511 (O_511,N_4787,N_4116);
nor UO_512 (O_512,N_4305,N_4226);
or UO_513 (O_513,N_4541,N_4676);
nand UO_514 (O_514,N_4741,N_4137);
nand UO_515 (O_515,N_4164,N_4142);
nand UO_516 (O_516,N_4750,N_4733);
nor UO_517 (O_517,N_4839,N_4127);
and UO_518 (O_518,N_4823,N_4563);
nand UO_519 (O_519,N_4560,N_4818);
nor UO_520 (O_520,N_4468,N_4591);
xor UO_521 (O_521,N_4819,N_4646);
nand UO_522 (O_522,N_4172,N_4302);
or UO_523 (O_523,N_4067,N_4198);
nor UO_524 (O_524,N_4123,N_4544);
nor UO_525 (O_525,N_4322,N_4267);
and UO_526 (O_526,N_4437,N_4810);
and UO_527 (O_527,N_4517,N_4514);
nor UO_528 (O_528,N_4455,N_4988);
and UO_529 (O_529,N_4473,N_4379);
nor UO_530 (O_530,N_4673,N_4388);
or UO_531 (O_531,N_4102,N_4668);
nand UO_532 (O_532,N_4032,N_4607);
nand UO_533 (O_533,N_4639,N_4218);
or UO_534 (O_534,N_4590,N_4376);
nor UO_535 (O_535,N_4454,N_4019);
and UO_536 (O_536,N_4891,N_4673);
or UO_537 (O_537,N_4040,N_4824);
nor UO_538 (O_538,N_4266,N_4820);
or UO_539 (O_539,N_4662,N_4428);
nand UO_540 (O_540,N_4072,N_4966);
nor UO_541 (O_541,N_4719,N_4922);
or UO_542 (O_542,N_4459,N_4085);
or UO_543 (O_543,N_4278,N_4096);
or UO_544 (O_544,N_4364,N_4522);
nand UO_545 (O_545,N_4536,N_4200);
nand UO_546 (O_546,N_4210,N_4622);
nor UO_547 (O_547,N_4863,N_4741);
and UO_548 (O_548,N_4422,N_4808);
or UO_549 (O_549,N_4278,N_4832);
and UO_550 (O_550,N_4309,N_4991);
or UO_551 (O_551,N_4825,N_4429);
nand UO_552 (O_552,N_4393,N_4192);
nand UO_553 (O_553,N_4272,N_4869);
nor UO_554 (O_554,N_4759,N_4546);
nand UO_555 (O_555,N_4073,N_4576);
nand UO_556 (O_556,N_4635,N_4765);
or UO_557 (O_557,N_4220,N_4908);
and UO_558 (O_558,N_4136,N_4002);
xor UO_559 (O_559,N_4230,N_4246);
or UO_560 (O_560,N_4905,N_4081);
nand UO_561 (O_561,N_4753,N_4828);
nand UO_562 (O_562,N_4644,N_4077);
nand UO_563 (O_563,N_4186,N_4670);
or UO_564 (O_564,N_4358,N_4198);
and UO_565 (O_565,N_4867,N_4072);
nand UO_566 (O_566,N_4476,N_4867);
nand UO_567 (O_567,N_4390,N_4876);
nand UO_568 (O_568,N_4468,N_4178);
nor UO_569 (O_569,N_4554,N_4849);
or UO_570 (O_570,N_4926,N_4132);
nor UO_571 (O_571,N_4750,N_4119);
and UO_572 (O_572,N_4412,N_4028);
and UO_573 (O_573,N_4953,N_4387);
nand UO_574 (O_574,N_4675,N_4309);
and UO_575 (O_575,N_4635,N_4464);
nor UO_576 (O_576,N_4224,N_4296);
nor UO_577 (O_577,N_4438,N_4299);
nand UO_578 (O_578,N_4279,N_4936);
or UO_579 (O_579,N_4787,N_4295);
nand UO_580 (O_580,N_4619,N_4596);
nor UO_581 (O_581,N_4329,N_4825);
nand UO_582 (O_582,N_4697,N_4893);
and UO_583 (O_583,N_4902,N_4410);
nand UO_584 (O_584,N_4864,N_4559);
nand UO_585 (O_585,N_4699,N_4945);
nand UO_586 (O_586,N_4764,N_4446);
nand UO_587 (O_587,N_4297,N_4762);
nor UO_588 (O_588,N_4741,N_4115);
nand UO_589 (O_589,N_4345,N_4249);
nand UO_590 (O_590,N_4054,N_4978);
nor UO_591 (O_591,N_4725,N_4887);
nor UO_592 (O_592,N_4294,N_4900);
or UO_593 (O_593,N_4459,N_4270);
and UO_594 (O_594,N_4485,N_4910);
or UO_595 (O_595,N_4107,N_4782);
and UO_596 (O_596,N_4841,N_4253);
nor UO_597 (O_597,N_4308,N_4555);
nand UO_598 (O_598,N_4024,N_4886);
nor UO_599 (O_599,N_4652,N_4868);
nand UO_600 (O_600,N_4658,N_4671);
nand UO_601 (O_601,N_4997,N_4010);
and UO_602 (O_602,N_4695,N_4683);
and UO_603 (O_603,N_4654,N_4760);
or UO_604 (O_604,N_4464,N_4074);
nor UO_605 (O_605,N_4041,N_4264);
and UO_606 (O_606,N_4786,N_4432);
nand UO_607 (O_607,N_4419,N_4815);
nand UO_608 (O_608,N_4319,N_4751);
nand UO_609 (O_609,N_4437,N_4239);
or UO_610 (O_610,N_4141,N_4531);
or UO_611 (O_611,N_4913,N_4641);
nand UO_612 (O_612,N_4859,N_4943);
nand UO_613 (O_613,N_4115,N_4850);
and UO_614 (O_614,N_4447,N_4378);
and UO_615 (O_615,N_4879,N_4756);
nor UO_616 (O_616,N_4780,N_4245);
or UO_617 (O_617,N_4313,N_4437);
nand UO_618 (O_618,N_4336,N_4556);
xor UO_619 (O_619,N_4386,N_4686);
xnor UO_620 (O_620,N_4181,N_4461);
or UO_621 (O_621,N_4439,N_4944);
nor UO_622 (O_622,N_4076,N_4920);
and UO_623 (O_623,N_4210,N_4953);
nor UO_624 (O_624,N_4851,N_4064);
nor UO_625 (O_625,N_4319,N_4926);
nand UO_626 (O_626,N_4580,N_4355);
nor UO_627 (O_627,N_4904,N_4132);
or UO_628 (O_628,N_4771,N_4130);
or UO_629 (O_629,N_4854,N_4389);
nor UO_630 (O_630,N_4982,N_4529);
nor UO_631 (O_631,N_4036,N_4952);
nor UO_632 (O_632,N_4802,N_4693);
nor UO_633 (O_633,N_4143,N_4009);
nand UO_634 (O_634,N_4580,N_4590);
nor UO_635 (O_635,N_4349,N_4745);
and UO_636 (O_636,N_4602,N_4046);
and UO_637 (O_637,N_4458,N_4980);
nor UO_638 (O_638,N_4121,N_4978);
or UO_639 (O_639,N_4161,N_4798);
and UO_640 (O_640,N_4786,N_4485);
nand UO_641 (O_641,N_4922,N_4016);
nand UO_642 (O_642,N_4794,N_4577);
or UO_643 (O_643,N_4429,N_4758);
or UO_644 (O_644,N_4379,N_4358);
and UO_645 (O_645,N_4874,N_4319);
nor UO_646 (O_646,N_4492,N_4405);
and UO_647 (O_647,N_4711,N_4063);
nand UO_648 (O_648,N_4418,N_4626);
or UO_649 (O_649,N_4848,N_4507);
nand UO_650 (O_650,N_4753,N_4954);
xor UO_651 (O_651,N_4158,N_4085);
nor UO_652 (O_652,N_4884,N_4847);
nor UO_653 (O_653,N_4193,N_4959);
nor UO_654 (O_654,N_4294,N_4360);
nor UO_655 (O_655,N_4919,N_4377);
nor UO_656 (O_656,N_4126,N_4961);
nand UO_657 (O_657,N_4370,N_4948);
and UO_658 (O_658,N_4715,N_4543);
and UO_659 (O_659,N_4942,N_4602);
or UO_660 (O_660,N_4967,N_4144);
nand UO_661 (O_661,N_4481,N_4390);
and UO_662 (O_662,N_4200,N_4847);
and UO_663 (O_663,N_4082,N_4971);
nand UO_664 (O_664,N_4197,N_4385);
nor UO_665 (O_665,N_4584,N_4026);
and UO_666 (O_666,N_4934,N_4548);
or UO_667 (O_667,N_4596,N_4608);
or UO_668 (O_668,N_4715,N_4869);
and UO_669 (O_669,N_4270,N_4613);
nand UO_670 (O_670,N_4685,N_4976);
nor UO_671 (O_671,N_4819,N_4631);
nor UO_672 (O_672,N_4893,N_4739);
or UO_673 (O_673,N_4076,N_4702);
nor UO_674 (O_674,N_4088,N_4815);
nand UO_675 (O_675,N_4791,N_4048);
nand UO_676 (O_676,N_4804,N_4676);
nor UO_677 (O_677,N_4733,N_4527);
and UO_678 (O_678,N_4595,N_4606);
or UO_679 (O_679,N_4881,N_4019);
and UO_680 (O_680,N_4873,N_4255);
nand UO_681 (O_681,N_4337,N_4424);
and UO_682 (O_682,N_4347,N_4078);
nor UO_683 (O_683,N_4428,N_4638);
nor UO_684 (O_684,N_4526,N_4200);
nand UO_685 (O_685,N_4288,N_4448);
nor UO_686 (O_686,N_4598,N_4196);
and UO_687 (O_687,N_4648,N_4421);
nor UO_688 (O_688,N_4285,N_4279);
nor UO_689 (O_689,N_4155,N_4128);
or UO_690 (O_690,N_4889,N_4716);
and UO_691 (O_691,N_4055,N_4071);
xnor UO_692 (O_692,N_4184,N_4539);
and UO_693 (O_693,N_4138,N_4979);
or UO_694 (O_694,N_4184,N_4212);
or UO_695 (O_695,N_4192,N_4211);
nor UO_696 (O_696,N_4672,N_4524);
and UO_697 (O_697,N_4261,N_4848);
or UO_698 (O_698,N_4531,N_4903);
or UO_699 (O_699,N_4985,N_4777);
nor UO_700 (O_700,N_4695,N_4247);
and UO_701 (O_701,N_4548,N_4899);
nor UO_702 (O_702,N_4292,N_4583);
or UO_703 (O_703,N_4151,N_4988);
and UO_704 (O_704,N_4191,N_4616);
nor UO_705 (O_705,N_4953,N_4353);
and UO_706 (O_706,N_4088,N_4669);
or UO_707 (O_707,N_4423,N_4912);
and UO_708 (O_708,N_4630,N_4884);
nor UO_709 (O_709,N_4362,N_4739);
nand UO_710 (O_710,N_4340,N_4884);
nand UO_711 (O_711,N_4224,N_4887);
or UO_712 (O_712,N_4070,N_4898);
nor UO_713 (O_713,N_4655,N_4928);
nor UO_714 (O_714,N_4716,N_4538);
and UO_715 (O_715,N_4059,N_4296);
nor UO_716 (O_716,N_4497,N_4333);
or UO_717 (O_717,N_4765,N_4407);
or UO_718 (O_718,N_4629,N_4606);
nand UO_719 (O_719,N_4181,N_4665);
xnor UO_720 (O_720,N_4375,N_4977);
nand UO_721 (O_721,N_4271,N_4979);
and UO_722 (O_722,N_4117,N_4662);
nor UO_723 (O_723,N_4601,N_4008);
or UO_724 (O_724,N_4355,N_4791);
nand UO_725 (O_725,N_4780,N_4142);
nand UO_726 (O_726,N_4948,N_4664);
and UO_727 (O_727,N_4500,N_4075);
or UO_728 (O_728,N_4800,N_4071);
nand UO_729 (O_729,N_4037,N_4644);
or UO_730 (O_730,N_4035,N_4369);
or UO_731 (O_731,N_4490,N_4267);
nand UO_732 (O_732,N_4282,N_4303);
nand UO_733 (O_733,N_4631,N_4963);
or UO_734 (O_734,N_4545,N_4546);
and UO_735 (O_735,N_4992,N_4719);
nor UO_736 (O_736,N_4793,N_4485);
and UO_737 (O_737,N_4344,N_4402);
nor UO_738 (O_738,N_4450,N_4682);
and UO_739 (O_739,N_4586,N_4989);
and UO_740 (O_740,N_4662,N_4869);
or UO_741 (O_741,N_4456,N_4816);
nand UO_742 (O_742,N_4425,N_4859);
and UO_743 (O_743,N_4671,N_4366);
nand UO_744 (O_744,N_4192,N_4048);
nor UO_745 (O_745,N_4076,N_4323);
or UO_746 (O_746,N_4839,N_4829);
or UO_747 (O_747,N_4897,N_4624);
or UO_748 (O_748,N_4097,N_4177);
and UO_749 (O_749,N_4460,N_4790);
nor UO_750 (O_750,N_4575,N_4822);
nand UO_751 (O_751,N_4587,N_4424);
or UO_752 (O_752,N_4208,N_4857);
nor UO_753 (O_753,N_4064,N_4841);
nand UO_754 (O_754,N_4156,N_4440);
and UO_755 (O_755,N_4843,N_4380);
or UO_756 (O_756,N_4991,N_4932);
and UO_757 (O_757,N_4540,N_4260);
and UO_758 (O_758,N_4519,N_4255);
nor UO_759 (O_759,N_4362,N_4022);
and UO_760 (O_760,N_4790,N_4166);
nor UO_761 (O_761,N_4161,N_4072);
and UO_762 (O_762,N_4032,N_4869);
nor UO_763 (O_763,N_4434,N_4809);
and UO_764 (O_764,N_4613,N_4036);
and UO_765 (O_765,N_4694,N_4597);
and UO_766 (O_766,N_4960,N_4341);
and UO_767 (O_767,N_4300,N_4781);
nor UO_768 (O_768,N_4018,N_4421);
or UO_769 (O_769,N_4847,N_4790);
and UO_770 (O_770,N_4904,N_4830);
and UO_771 (O_771,N_4750,N_4832);
and UO_772 (O_772,N_4447,N_4498);
nand UO_773 (O_773,N_4058,N_4310);
nor UO_774 (O_774,N_4696,N_4924);
nand UO_775 (O_775,N_4712,N_4071);
or UO_776 (O_776,N_4489,N_4275);
or UO_777 (O_777,N_4197,N_4757);
or UO_778 (O_778,N_4459,N_4138);
and UO_779 (O_779,N_4066,N_4917);
nor UO_780 (O_780,N_4296,N_4225);
and UO_781 (O_781,N_4226,N_4921);
nor UO_782 (O_782,N_4802,N_4901);
nor UO_783 (O_783,N_4244,N_4360);
nand UO_784 (O_784,N_4859,N_4626);
nand UO_785 (O_785,N_4703,N_4305);
nor UO_786 (O_786,N_4423,N_4130);
nand UO_787 (O_787,N_4854,N_4380);
or UO_788 (O_788,N_4345,N_4712);
nor UO_789 (O_789,N_4540,N_4180);
nor UO_790 (O_790,N_4323,N_4070);
or UO_791 (O_791,N_4037,N_4984);
or UO_792 (O_792,N_4105,N_4029);
nor UO_793 (O_793,N_4855,N_4633);
xnor UO_794 (O_794,N_4680,N_4035);
and UO_795 (O_795,N_4415,N_4208);
and UO_796 (O_796,N_4085,N_4345);
or UO_797 (O_797,N_4762,N_4832);
or UO_798 (O_798,N_4001,N_4747);
nor UO_799 (O_799,N_4415,N_4079);
or UO_800 (O_800,N_4753,N_4308);
and UO_801 (O_801,N_4782,N_4031);
nand UO_802 (O_802,N_4215,N_4694);
nor UO_803 (O_803,N_4540,N_4751);
nand UO_804 (O_804,N_4884,N_4530);
or UO_805 (O_805,N_4026,N_4562);
and UO_806 (O_806,N_4415,N_4055);
and UO_807 (O_807,N_4840,N_4547);
nor UO_808 (O_808,N_4151,N_4657);
nor UO_809 (O_809,N_4604,N_4074);
and UO_810 (O_810,N_4736,N_4637);
and UO_811 (O_811,N_4730,N_4759);
nor UO_812 (O_812,N_4475,N_4272);
nor UO_813 (O_813,N_4249,N_4853);
xnor UO_814 (O_814,N_4750,N_4972);
nand UO_815 (O_815,N_4301,N_4648);
nor UO_816 (O_816,N_4854,N_4390);
nand UO_817 (O_817,N_4813,N_4097);
or UO_818 (O_818,N_4754,N_4406);
or UO_819 (O_819,N_4527,N_4827);
and UO_820 (O_820,N_4803,N_4342);
nand UO_821 (O_821,N_4119,N_4345);
nor UO_822 (O_822,N_4406,N_4901);
and UO_823 (O_823,N_4276,N_4461);
and UO_824 (O_824,N_4759,N_4994);
nand UO_825 (O_825,N_4905,N_4833);
or UO_826 (O_826,N_4008,N_4658);
and UO_827 (O_827,N_4382,N_4641);
nor UO_828 (O_828,N_4273,N_4288);
nor UO_829 (O_829,N_4819,N_4962);
nand UO_830 (O_830,N_4086,N_4229);
and UO_831 (O_831,N_4189,N_4607);
or UO_832 (O_832,N_4756,N_4557);
nor UO_833 (O_833,N_4835,N_4906);
and UO_834 (O_834,N_4008,N_4524);
nand UO_835 (O_835,N_4527,N_4162);
nand UO_836 (O_836,N_4840,N_4382);
nand UO_837 (O_837,N_4218,N_4474);
and UO_838 (O_838,N_4150,N_4891);
nor UO_839 (O_839,N_4210,N_4084);
or UO_840 (O_840,N_4692,N_4311);
and UO_841 (O_841,N_4669,N_4410);
xor UO_842 (O_842,N_4515,N_4419);
nand UO_843 (O_843,N_4206,N_4968);
nor UO_844 (O_844,N_4851,N_4886);
nor UO_845 (O_845,N_4247,N_4690);
or UO_846 (O_846,N_4261,N_4162);
and UO_847 (O_847,N_4819,N_4640);
nor UO_848 (O_848,N_4952,N_4498);
or UO_849 (O_849,N_4037,N_4589);
and UO_850 (O_850,N_4764,N_4594);
nor UO_851 (O_851,N_4898,N_4299);
nor UO_852 (O_852,N_4074,N_4327);
or UO_853 (O_853,N_4324,N_4543);
or UO_854 (O_854,N_4349,N_4736);
nor UO_855 (O_855,N_4679,N_4390);
or UO_856 (O_856,N_4896,N_4916);
or UO_857 (O_857,N_4007,N_4919);
and UO_858 (O_858,N_4139,N_4951);
and UO_859 (O_859,N_4227,N_4014);
and UO_860 (O_860,N_4791,N_4496);
or UO_861 (O_861,N_4871,N_4769);
xnor UO_862 (O_862,N_4539,N_4455);
or UO_863 (O_863,N_4455,N_4524);
nand UO_864 (O_864,N_4167,N_4735);
and UO_865 (O_865,N_4660,N_4688);
and UO_866 (O_866,N_4194,N_4337);
and UO_867 (O_867,N_4437,N_4352);
nor UO_868 (O_868,N_4261,N_4996);
and UO_869 (O_869,N_4177,N_4355);
nand UO_870 (O_870,N_4326,N_4155);
and UO_871 (O_871,N_4189,N_4513);
nand UO_872 (O_872,N_4871,N_4157);
nor UO_873 (O_873,N_4137,N_4148);
nor UO_874 (O_874,N_4245,N_4901);
nor UO_875 (O_875,N_4606,N_4829);
nor UO_876 (O_876,N_4574,N_4501);
and UO_877 (O_877,N_4811,N_4231);
nand UO_878 (O_878,N_4895,N_4312);
or UO_879 (O_879,N_4403,N_4875);
and UO_880 (O_880,N_4650,N_4115);
and UO_881 (O_881,N_4707,N_4125);
and UO_882 (O_882,N_4379,N_4387);
nor UO_883 (O_883,N_4243,N_4220);
or UO_884 (O_884,N_4605,N_4610);
nor UO_885 (O_885,N_4772,N_4739);
nor UO_886 (O_886,N_4285,N_4979);
and UO_887 (O_887,N_4039,N_4997);
nand UO_888 (O_888,N_4564,N_4598);
nor UO_889 (O_889,N_4259,N_4468);
nand UO_890 (O_890,N_4259,N_4186);
or UO_891 (O_891,N_4499,N_4190);
nor UO_892 (O_892,N_4982,N_4877);
nor UO_893 (O_893,N_4155,N_4607);
nor UO_894 (O_894,N_4963,N_4147);
nand UO_895 (O_895,N_4068,N_4134);
or UO_896 (O_896,N_4153,N_4075);
and UO_897 (O_897,N_4952,N_4781);
nand UO_898 (O_898,N_4724,N_4614);
nand UO_899 (O_899,N_4974,N_4778);
and UO_900 (O_900,N_4939,N_4595);
or UO_901 (O_901,N_4618,N_4398);
nor UO_902 (O_902,N_4499,N_4508);
nor UO_903 (O_903,N_4089,N_4046);
or UO_904 (O_904,N_4053,N_4609);
or UO_905 (O_905,N_4232,N_4710);
and UO_906 (O_906,N_4658,N_4339);
nor UO_907 (O_907,N_4524,N_4070);
and UO_908 (O_908,N_4342,N_4271);
nand UO_909 (O_909,N_4984,N_4193);
nor UO_910 (O_910,N_4657,N_4624);
and UO_911 (O_911,N_4726,N_4382);
nand UO_912 (O_912,N_4136,N_4559);
or UO_913 (O_913,N_4167,N_4829);
nor UO_914 (O_914,N_4038,N_4157);
nand UO_915 (O_915,N_4530,N_4272);
nor UO_916 (O_916,N_4911,N_4931);
or UO_917 (O_917,N_4248,N_4874);
xor UO_918 (O_918,N_4761,N_4976);
nor UO_919 (O_919,N_4448,N_4772);
or UO_920 (O_920,N_4299,N_4945);
or UO_921 (O_921,N_4977,N_4640);
nor UO_922 (O_922,N_4283,N_4444);
nor UO_923 (O_923,N_4203,N_4018);
or UO_924 (O_924,N_4536,N_4599);
nand UO_925 (O_925,N_4325,N_4775);
nand UO_926 (O_926,N_4720,N_4163);
nand UO_927 (O_927,N_4455,N_4353);
nand UO_928 (O_928,N_4585,N_4588);
nor UO_929 (O_929,N_4410,N_4242);
or UO_930 (O_930,N_4630,N_4660);
nor UO_931 (O_931,N_4076,N_4241);
nor UO_932 (O_932,N_4895,N_4149);
nand UO_933 (O_933,N_4546,N_4439);
nand UO_934 (O_934,N_4020,N_4843);
or UO_935 (O_935,N_4795,N_4245);
or UO_936 (O_936,N_4411,N_4214);
nand UO_937 (O_937,N_4193,N_4329);
or UO_938 (O_938,N_4660,N_4498);
and UO_939 (O_939,N_4596,N_4853);
nand UO_940 (O_940,N_4999,N_4709);
and UO_941 (O_941,N_4673,N_4347);
nand UO_942 (O_942,N_4876,N_4444);
nor UO_943 (O_943,N_4769,N_4365);
and UO_944 (O_944,N_4936,N_4099);
nand UO_945 (O_945,N_4417,N_4099);
nand UO_946 (O_946,N_4046,N_4925);
nand UO_947 (O_947,N_4008,N_4151);
or UO_948 (O_948,N_4497,N_4255);
or UO_949 (O_949,N_4266,N_4358);
nand UO_950 (O_950,N_4070,N_4308);
nand UO_951 (O_951,N_4902,N_4651);
nor UO_952 (O_952,N_4574,N_4548);
and UO_953 (O_953,N_4866,N_4875);
nor UO_954 (O_954,N_4188,N_4288);
and UO_955 (O_955,N_4591,N_4833);
nor UO_956 (O_956,N_4889,N_4452);
or UO_957 (O_957,N_4317,N_4441);
or UO_958 (O_958,N_4507,N_4079);
nand UO_959 (O_959,N_4431,N_4993);
or UO_960 (O_960,N_4715,N_4634);
nand UO_961 (O_961,N_4235,N_4528);
or UO_962 (O_962,N_4523,N_4043);
nand UO_963 (O_963,N_4688,N_4464);
or UO_964 (O_964,N_4506,N_4355);
and UO_965 (O_965,N_4433,N_4705);
or UO_966 (O_966,N_4569,N_4026);
nor UO_967 (O_967,N_4563,N_4568);
nand UO_968 (O_968,N_4587,N_4259);
nand UO_969 (O_969,N_4947,N_4263);
nor UO_970 (O_970,N_4720,N_4679);
and UO_971 (O_971,N_4098,N_4749);
nand UO_972 (O_972,N_4125,N_4317);
or UO_973 (O_973,N_4860,N_4641);
nand UO_974 (O_974,N_4111,N_4508);
or UO_975 (O_975,N_4575,N_4887);
and UO_976 (O_976,N_4986,N_4792);
nand UO_977 (O_977,N_4171,N_4943);
or UO_978 (O_978,N_4966,N_4607);
nand UO_979 (O_979,N_4827,N_4288);
and UO_980 (O_980,N_4281,N_4828);
nand UO_981 (O_981,N_4219,N_4423);
nand UO_982 (O_982,N_4372,N_4464);
xor UO_983 (O_983,N_4809,N_4638);
and UO_984 (O_984,N_4386,N_4339);
or UO_985 (O_985,N_4396,N_4446);
nand UO_986 (O_986,N_4450,N_4424);
or UO_987 (O_987,N_4611,N_4367);
and UO_988 (O_988,N_4067,N_4313);
or UO_989 (O_989,N_4339,N_4790);
or UO_990 (O_990,N_4954,N_4295);
nand UO_991 (O_991,N_4935,N_4467);
nand UO_992 (O_992,N_4517,N_4226);
nor UO_993 (O_993,N_4053,N_4270);
and UO_994 (O_994,N_4998,N_4191);
or UO_995 (O_995,N_4220,N_4038);
nor UO_996 (O_996,N_4014,N_4703);
nand UO_997 (O_997,N_4454,N_4828);
nand UO_998 (O_998,N_4091,N_4375);
and UO_999 (O_999,N_4231,N_4520);
endmodule