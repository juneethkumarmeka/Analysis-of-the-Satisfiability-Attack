module basic_500_3000_500_50_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_436,In_13);
and U1 (N_1,In_104,In_475);
nand U2 (N_2,In_413,In_490);
and U3 (N_3,In_170,In_169);
or U4 (N_4,In_88,In_183);
or U5 (N_5,In_155,In_288);
nand U6 (N_6,In_497,In_319);
or U7 (N_7,In_146,In_215);
and U8 (N_8,In_52,In_495);
or U9 (N_9,In_37,In_164);
xnor U10 (N_10,In_381,In_453);
nand U11 (N_11,In_347,In_270);
nand U12 (N_12,In_289,In_305);
xnor U13 (N_13,In_236,In_247);
and U14 (N_14,In_228,In_130);
and U15 (N_15,In_12,In_244);
nor U16 (N_16,In_158,In_229);
nand U17 (N_17,In_486,In_129);
nand U18 (N_18,In_121,In_120);
and U19 (N_19,In_78,In_338);
or U20 (N_20,In_156,In_85);
and U21 (N_21,In_177,In_202);
xor U22 (N_22,In_14,In_329);
and U23 (N_23,In_160,In_246);
or U24 (N_24,In_137,In_439);
or U25 (N_25,In_191,In_362);
or U26 (N_26,In_340,In_252);
and U27 (N_27,In_293,In_421);
or U28 (N_28,In_352,In_400);
nor U29 (N_29,In_326,In_374);
or U30 (N_30,In_61,In_282);
or U31 (N_31,In_272,In_141);
nand U32 (N_32,In_300,In_150);
xor U33 (N_33,In_101,In_111);
xor U34 (N_34,In_212,In_240);
nor U35 (N_35,In_344,In_380);
or U36 (N_36,In_368,In_455);
nor U37 (N_37,In_280,In_356);
xor U38 (N_38,In_234,In_67);
or U39 (N_39,In_10,In_124);
xnor U40 (N_40,In_309,In_286);
nand U41 (N_41,In_378,In_437);
and U42 (N_42,In_242,In_103);
nand U43 (N_43,In_446,In_379);
nor U44 (N_44,In_408,In_335);
and U45 (N_45,In_245,In_306);
or U46 (N_46,In_197,In_96);
and U47 (N_47,In_256,In_87);
and U48 (N_48,In_71,In_287);
and U49 (N_49,In_154,In_302);
nor U50 (N_50,In_366,In_79);
or U51 (N_51,In_296,In_72);
xnor U52 (N_52,In_136,In_114);
xor U53 (N_53,In_369,In_435);
and U54 (N_54,In_310,In_251);
nor U55 (N_55,In_98,In_449);
or U56 (N_56,In_377,In_55);
and U57 (N_57,In_94,In_152);
nor U58 (N_58,In_291,In_482);
xnor U59 (N_59,In_20,In_48);
and U60 (N_60,In_97,In_263);
xnor U61 (N_61,In_6,In_307);
or U62 (N_62,N_27,In_483);
and U63 (N_63,In_469,In_468);
nor U64 (N_64,In_123,In_303);
or U65 (N_65,In_91,N_9);
nand U66 (N_66,In_144,In_203);
or U67 (N_67,N_21,N_35);
xor U68 (N_68,In_450,In_117);
or U69 (N_69,In_2,In_56);
nor U70 (N_70,N_31,In_195);
xor U71 (N_71,In_151,In_334);
nand U72 (N_72,In_180,In_418);
nand U73 (N_73,In_32,N_4);
nand U74 (N_74,N_8,In_53);
nand U75 (N_75,In_443,In_69);
nor U76 (N_76,In_28,In_273);
nand U77 (N_77,In_54,In_29);
nor U78 (N_78,In_190,In_386);
nor U79 (N_79,In_162,In_159);
xor U80 (N_80,In_488,In_447);
xor U81 (N_81,In_161,In_66);
or U82 (N_82,In_385,In_253);
or U83 (N_83,In_312,In_138);
nand U84 (N_84,In_233,In_11);
nor U85 (N_85,In_58,In_208);
nand U86 (N_86,In_115,In_354);
and U87 (N_87,N_56,In_188);
nor U88 (N_88,N_40,In_39);
and U89 (N_89,In_186,In_370);
or U90 (N_90,N_19,In_285);
or U91 (N_91,In_393,In_485);
xor U92 (N_92,In_178,N_26);
xnor U93 (N_93,N_25,In_142);
or U94 (N_94,In_358,In_339);
nor U95 (N_95,In_214,In_49);
nand U96 (N_96,In_82,N_41);
or U97 (N_97,In_411,In_70);
xor U98 (N_98,In_281,In_412);
and U99 (N_99,In_360,In_193);
nand U100 (N_100,In_390,In_399);
or U101 (N_101,In_403,N_52);
and U102 (N_102,In_398,In_119);
or U103 (N_103,In_131,In_239);
and U104 (N_104,N_6,In_147);
or U105 (N_105,In_425,In_409);
nor U106 (N_106,In_187,In_36);
and U107 (N_107,In_81,In_462);
nor U108 (N_108,In_185,In_128);
nor U109 (N_109,In_218,In_149);
and U110 (N_110,In_265,In_254);
or U111 (N_111,N_7,In_496);
nand U112 (N_112,In_417,N_45);
nand U113 (N_113,In_416,In_423);
or U114 (N_114,In_241,N_13);
or U115 (N_115,In_461,In_51);
nor U116 (N_116,In_176,In_313);
xnor U117 (N_117,In_471,In_168);
nor U118 (N_118,In_41,In_24);
nand U119 (N_119,In_127,In_118);
xor U120 (N_120,N_44,In_116);
xor U121 (N_121,In_80,In_15);
nand U122 (N_122,N_70,In_456);
xnor U123 (N_123,In_480,In_93);
or U124 (N_124,N_66,N_62);
or U125 (N_125,In_392,In_424);
or U126 (N_126,In_199,In_383);
xnor U127 (N_127,N_72,N_73);
or U128 (N_128,In_126,In_179);
and U129 (N_129,N_17,In_62);
nor U130 (N_130,In_258,N_88);
and U131 (N_131,N_117,In_477);
and U132 (N_132,In_57,In_325);
nand U133 (N_133,In_181,In_9);
nor U134 (N_134,In_414,In_46);
nor U135 (N_135,In_295,In_232);
nor U136 (N_136,N_84,In_442);
nor U137 (N_137,In_132,In_262);
or U138 (N_138,In_341,N_42);
and U139 (N_139,In_75,In_298);
nor U140 (N_140,In_259,N_2);
xor U141 (N_141,In_27,In_478);
or U142 (N_142,In_311,N_3);
and U143 (N_143,In_153,N_80);
xnor U144 (N_144,In_394,In_207);
nor U145 (N_145,In_444,In_322);
nor U146 (N_146,In_60,N_71);
or U147 (N_147,In_34,In_292);
or U148 (N_148,In_107,In_64);
xor U149 (N_149,In_174,In_493);
nor U150 (N_150,In_472,N_77);
nor U151 (N_151,In_200,In_38);
and U152 (N_152,In_431,N_63);
xor U153 (N_153,N_58,In_261);
xor U154 (N_154,In_430,In_125);
nand U155 (N_155,N_92,In_112);
nor U156 (N_156,In_166,N_5);
xnor U157 (N_157,In_276,In_299);
and U158 (N_158,N_82,N_75);
nand U159 (N_159,In_110,In_221);
nor U160 (N_160,In_106,N_64);
xnor U161 (N_161,In_42,In_134);
or U162 (N_162,In_460,N_94);
or U163 (N_163,In_315,In_135);
nor U164 (N_164,In_422,In_372);
xnor U165 (N_165,In_109,N_114);
nor U166 (N_166,In_84,In_491);
nand U167 (N_167,N_39,In_90);
xor U168 (N_168,In_209,In_463);
xor U169 (N_169,N_87,In_50);
or U170 (N_170,N_29,In_357);
nor U171 (N_171,N_86,In_382);
or U172 (N_172,In_458,In_448);
and U173 (N_173,In_225,In_182);
and U174 (N_174,In_184,In_459);
xor U175 (N_175,In_30,In_434);
and U176 (N_176,In_314,In_77);
and U177 (N_177,In_31,In_337);
xnor U178 (N_178,N_54,In_316);
xnor U179 (N_179,N_22,In_17);
nand U180 (N_180,In_328,N_61);
nand U181 (N_181,In_465,In_391);
xnor U182 (N_182,N_98,N_131);
nor U183 (N_183,In_1,N_89);
or U184 (N_184,In_33,N_107);
or U185 (N_185,N_104,N_158);
nand U186 (N_186,In_321,N_30);
nor U187 (N_187,In_264,N_59);
or U188 (N_188,In_257,N_157);
xnor U189 (N_189,N_164,In_25);
or U190 (N_190,N_134,In_405);
xor U191 (N_191,In_238,In_330);
xor U192 (N_192,N_142,N_169);
xor U193 (N_193,In_301,In_196);
or U194 (N_194,In_499,In_139);
and U195 (N_195,In_359,N_160);
and U196 (N_196,In_226,In_349);
or U197 (N_197,N_10,N_99);
nor U198 (N_198,In_324,N_67);
nor U199 (N_199,In_432,In_133);
nor U200 (N_200,N_48,N_47);
or U201 (N_201,In_5,N_118);
and U202 (N_202,In_420,N_110);
nand U203 (N_203,In_397,In_364);
nor U204 (N_204,In_343,N_85);
nor U205 (N_205,In_220,N_14);
and U206 (N_206,N_100,N_141);
nor U207 (N_207,In_426,N_128);
nand U208 (N_208,In_248,N_132);
or U209 (N_209,In_277,In_205);
and U210 (N_210,N_171,In_74);
xnor U211 (N_211,N_123,N_116);
or U212 (N_212,N_150,In_428);
nor U213 (N_213,In_275,In_363);
nor U214 (N_214,N_168,In_375);
nor U215 (N_215,N_83,N_51);
nor U216 (N_216,In_95,N_20);
nor U217 (N_217,In_223,In_407);
nor U218 (N_218,In_65,N_46);
nand U219 (N_219,In_192,In_317);
and U220 (N_220,In_86,In_278);
and U221 (N_221,N_161,N_156);
nand U222 (N_222,N_32,In_165);
or U223 (N_223,N_109,In_355);
and U224 (N_224,In_140,N_93);
or U225 (N_225,In_108,N_121);
nor U226 (N_226,In_213,N_127);
and U227 (N_227,In_83,In_473);
nor U228 (N_228,In_402,In_63);
or U229 (N_229,In_249,N_176);
and U230 (N_230,In_206,In_323);
nor U231 (N_231,In_384,In_255);
nand U232 (N_232,In_4,In_243);
xor U233 (N_233,N_148,N_149);
xor U234 (N_234,N_167,In_367);
nand U235 (N_235,In_451,In_452);
and U236 (N_236,N_102,In_476);
nand U237 (N_237,In_204,N_60);
nor U238 (N_238,In_318,N_170);
xnor U239 (N_239,In_7,N_81);
nand U240 (N_240,N_198,N_108);
nor U241 (N_241,N_124,N_188);
xor U242 (N_242,In_470,In_73);
xor U243 (N_243,N_126,In_173);
or U244 (N_244,In_8,In_492);
or U245 (N_245,N_213,In_175);
xor U246 (N_246,N_178,In_353);
nor U247 (N_247,In_113,N_208);
nand U248 (N_248,In_100,N_234);
or U249 (N_249,N_140,In_267);
nand U250 (N_250,N_101,In_331);
nand U251 (N_251,N_115,N_207);
nor U252 (N_252,In_487,In_283);
xor U253 (N_253,N_236,N_34);
nor U254 (N_254,In_294,N_209);
and U255 (N_255,In_404,In_237);
or U256 (N_256,N_90,In_327);
xor U257 (N_257,N_214,N_112);
or U258 (N_258,In_16,N_139);
xor U259 (N_259,N_189,In_260);
or U260 (N_260,In_148,In_68);
and U261 (N_261,N_129,N_230);
and U262 (N_262,In_410,In_336);
and U263 (N_263,In_224,N_136);
and U264 (N_264,In_467,In_44);
or U265 (N_265,N_12,In_433);
or U266 (N_266,N_190,N_155);
nor U267 (N_267,In_489,N_222);
nand U268 (N_268,N_18,N_196);
xnor U269 (N_269,In_346,N_36);
nand U270 (N_270,In_201,N_147);
and U271 (N_271,In_89,N_144);
nor U272 (N_272,In_219,In_498);
nor U273 (N_273,N_203,In_479);
nor U274 (N_274,N_76,N_216);
xnor U275 (N_275,N_165,N_65);
xnor U276 (N_276,In_454,In_396);
xnor U277 (N_277,N_231,N_229);
xor U278 (N_278,In_429,N_137);
xor U279 (N_279,In_406,N_177);
xor U280 (N_280,In_59,In_304);
nand U281 (N_281,In_395,In_350);
nand U282 (N_282,In_122,In_211);
nand U283 (N_283,In_279,In_40);
nor U284 (N_284,N_119,In_19);
nand U285 (N_285,In_345,N_111);
and U286 (N_286,N_152,In_376);
nand U287 (N_287,In_216,In_333);
xor U288 (N_288,In_157,N_184);
nand U289 (N_289,In_415,In_222);
xnor U290 (N_290,In_320,N_57);
nand U291 (N_291,N_38,In_427);
nor U292 (N_292,N_163,N_219);
nand U293 (N_293,N_69,In_474);
nand U294 (N_294,In_171,In_231);
xnor U295 (N_295,N_224,In_388);
nand U296 (N_296,In_230,In_348);
nand U297 (N_297,N_215,In_290);
or U298 (N_298,N_210,N_146);
nor U299 (N_299,N_206,In_438);
and U300 (N_300,N_195,N_239);
or U301 (N_301,N_221,N_24);
and U302 (N_302,N_295,In_464);
and U303 (N_303,In_189,N_299);
nor U304 (N_304,N_228,In_167);
or U305 (N_305,N_74,In_332);
nand U306 (N_306,In_250,N_251);
and U307 (N_307,N_223,N_194);
and U308 (N_308,N_280,In_284);
nor U309 (N_309,N_266,In_194);
nand U310 (N_310,N_252,N_151);
nor U311 (N_311,N_106,N_218);
nor U312 (N_312,N_37,N_293);
nor U313 (N_313,N_91,N_276);
and U314 (N_314,N_284,N_23);
nor U315 (N_315,N_285,N_217);
xor U316 (N_316,N_133,N_288);
nand U317 (N_317,N_237,N_296);
nand U318 (N_318,In_198,N_245);
xnor U319 (N_319,N_200,N_179);
and U320 (N_320,N_247,N_175);
xor U321 (N_321,N_277,In_297);
nand U322 (N_322,In_102,N_153);
xor U323 (N_323,In_163,In_361);
nand U324 (N_324,N_264,In_457);
nand U325 (N_325,N_244,N_95);
or U326 (N_326,In_445,N_254);
xnor U327 (N_327,N_253,In_0);
xnor U328 (N_328,In_365,In_419);
or U329 (N_329,In_441,N_53);
nand U330 (N_330,N_113,N_130);
nor U331 (N_331,N_16,N_267);
and U332 (N_332,N_182,N_1);
nand U333 (N_333,N_241,In_76);
nand U334 (N_334,N_273,N_271);
or U335 (N_335,In_342,N_290);
xnor U336 (N_336,N_242,N_181);
nand U337 (N_337,N_49,In_217);
xnor U338 (N_338,In_274,In_271);
nand U339 (N_339,In_35,In_440);
xor U340 (N_340,N_270,N_211);
xor U341 (N_341,N_105,N_268);
nand U342 (N_342,N_238,In_268);
and U343 (N_343,N_192,N_235);
or U344 (N_344,N_281,N_278);
and U345 (N_345,In_47,N_249);
or U346 (N_346,N_78,N_11);
xor U347 (N_347,In_18,In_23);
nand U348 (N_348,N_201,N_265);
nor U349 (N_349,N_97,N_291);
nor U350 (N_350,N_261,N_187);
nand U351 (N_351,In_22,N_255);
nand U352 (N_352,N_257,In_308);
and U353 (N_353,N_232,N_240);
or U354 (N_354,N_246,N_103);
nand U355 (N_355,In_235,In_351);
or U356 (N_356,N_287,N_28);
nand U357 (N_357,In_172,N_263);
and U358 (N_358,N_202,N_186);
nor U359 (N_359,N_212,N_183);
and U360 (N_360,In_266,N_122);
xnor U361 (N_361,N_145,In_401);
and U362 (N_362,N_303,N_322);
nor U363 (N_363,N_333,N_316);
and U364 (N_364,N_225,N_248);
xnor U365 (N_365,N_256,N_283);
or U366 (N_366,N_301,N_300);
or U367 (N_367,N_43,N_358);
nor U368 (N_368,In_21,N_180);
nand U369 (N_369,N_185,N_346);
nand U370 (N_370,In_494,N_338);
or U371 (N_371,N_313,In_210);
and U372 (N_372,In_389,N_272);
nor U373 (N_373,N_205,In_373);
and U374 (N_374,N_220,N_325);
xor U375 (N_375,N_310,N_259);
xor U376 (N_376,In_481,N_354);
nor U377 (N_377,N_306,N_309);
and U378 (N_378,N_197,N_135);
or U379 (N_379,N_345,N_274);
and U380 (N_380,N_0,N_226);
and U381 (N_381,N_351,In_371);
or U382 (N_382,N_191,N_143);
and U383 (N_383,N_138,In_45);
xnor U384 (N_384,N_243,N_279);
or U385 (N_385,In_26,N_342);
and U386 (N_386,N_233,N_314);
or U387 (N_387,N_312,N_305);
nand U388 (N_388,N_359,N_341);
xnor U389 (N_389,N_327,N_340);
xnor U390 (N_390,N_292,N_347);
or U391 (N_391,N_125,In_269);
nor U392 (N_392,N_357,N_162);
xor U393 (N_393,N_302,N_258);
and U394 (N_394,N_337,N_286);
nor U395 (N_395,N_174,N_318);
or U396 (N_396,N_298,N_320);
and U397 (N_397,N_353,N_311);
xor U398 (N_398,N_355,N_308);
xnor U399 (N_399,N_172,N_294);
xor U400 (N_400,N_329,N_260);
xor U401 (N_401,N_315,N_159);
nor U402 (N_402,N_68,N_250);
nand U403 (N_403,N_326,N_227);
or U404 (N_404,N_335,N_269);
or U405 (N_405,N_348,N_356);
or U406 (N_406,N_324,In_99);
nand U407 (N_407,N_352,In_43);
or U408 (N_408,N_50,N_323);
nand U409 (N_409,N_282,In_92);
xnor U410 (N_410,N_297,N_33);
xnor U411 (N_411,N_319,N_79);
nor U412 (N_412,In_227,N_344);
nand U413 (N_413,N_204,N_166);
nand U414 (N_414,N_350,In_105);
and U415 (N_415,N_321,N_330);
and U416 (N_416,N_317,N_289);
or U417 (N_417,In_3,N_343);
xnor U418 (N_418,N_199,N_96);
nor U419 (N_419,N_334,In_387);
nor U420 (N_420,N_382,N_417);
nand U421 (N_421,N_328,N_419);
and U422 (N_422,N_415,N_362);
and U423 (N_423,N_120,N_385);
xnor U424 (N_424,In_145,N_413);
and U425 (N_425,N_360,N_275);
xor U426 (N_426,N_388,N_332);
or U427 (N_427,N_383,N_365);
nor U428 (N_428,N_399,N_387);
or U429 (N_429,N_395,In_466);
nor U430 (N_430,N_400,N_389);
nand U431 (N_431,N_307,N_411);
or U432 (N_432,N_374,N_416);
xnor U433 (N_433,N_418,N_336);
nor U434 (N_434,N_369,N_366);
nor U435 (N_435,In_143,N_404);
nand U436 (N_436,N_394,In_484);
nor U437 (N_437,N_401,N_154);
xor U438 (N_438,N_55,N_173);
or U439 (N_439,N_339,N_349);
xnor U440 (N_440,N_409,N_368);
nand U441 (N_441,N_361,N_402);
nand U442 (N_442,N_392,N_397);
and U443 (N_443,N_414,N_412);
nor U444 (N_444,N_380,N_370);
or U445 (N_445,N_15,N_403);
and U446 (N_446,N_384,N_410);
or U447 (N_447,N_405,N_364);
or U448 (N_448,N_378,N_393);
xnor U449 (N_449,N_386,N_375);
or U450 (N_450,N_371,N_331);
and U451 (N_451,N_377,N_363);
or U452 (N_452,N_372,N_367);
nand U453 (N_453,N_193,N_407);
xor U454 (N_454,N_390,N_381);
nor U455 (N_455,N_391,N_406);
xnor U456 (N_456,N_373,N_379);
xnor U457 (N_457,N_398,N_396);
nand U458 (N_458,N_262,N_304);
xor U459 (N_459,N_376,N_408);
nand U460 (N_460,N_378,N_398);
or U461 (N_461,N_120,N_408);
xnor U462 (N_462,N_391,N_349);
nor U463 (N_463,N_275,N_389);
or U464 (N_464,N_364,N_403);
or U465 (N_465,N_398,N_55);
or U466 (N_466,N_275,N_368);
nor U467 (N_467,N_386,N_368);
nand U468 (N_468,N_366,N_414);
xnor U469 (N_469,N_369,N_405);
or U470 (N_470,N_154,N_375);
nand U471 (N_471,N_401,N_370);
and U472 (N_472,N_55,N_392);
and U473 (N_473,N_360,N_394);
or U474 (N_474,N_398,N_371);
nor U475 (N_475,N_407,N_392);
nand U476 (N_476,N_395,N_331);
or U477 (N_477,N_388,N_385);
or U478 (N_478,N_383,In_466);
xnor U479 (N_479,N_375,In_466);
or U480 (N_480,N_438,N_462);
nand U481 (N_481,N_435,N_479);
xnor U482 (N_482,N_456,N_461);
and U483 (N_483,N_434,N_463);
or U484 (N_484,N_420,N_437);
and U485 (N_485,N_430,N_422);
and U486 (N_486,N_428,N_455);
nand U487 (N_487,N_476,N_471);
nor U488 (N_488,N_449,N_429);
or U489 (N_489,N_425,N_431);
or U490 (N_490,N_472,N_424);
nor U491 (N_491,N_477,N_446);
and U492 (N_492,N_460,N_454);
or U493 (N_493,N_453,N_465);
and U494 (N_494,N_423,N_436);
and U495 (N_495,N_426,N_473);
nand U496 (N_496,N_433,N_464);
nor U497 (N_497,N_442,N_469);
nor U498 (N_498,N_440,N_448);
xnor U499 (N_499,N_475,N_474);
nor U500 (N_500,N_458,N_467);
and U501 (N_501,N_444,N_427);
nand U502 (N_502,N_468,N_445);
xnor U503 (N_503,N_450,N_470);
or U504 (N_504,N_441,N_457);
xnor U505 (N_505,N_478,N_452);
nor U506 (N_506,N_432,N_459);
xnor U507 (N_507,N_443,N_421);
xor U508 (N_508,N_466,N_451);
nand U509 (N_509,N_439,N_447);
and U510 (N_510,N_475,N_473);
and U511 (N_511,N_477,N_439);
nor U512 (N_512,N_444,N_423);
nor U513 (N_513,N_479,N_437);
nand U514 (N_514,N_451,N_453);
or U515 (N_515,N_436,N_424);
nor U516 (N_516,N_443,N_429);
and U517 (N_517,N_427,N_451);
or U518 (N_518,N_479,N_434);
xnor U519 (N_519,N_456,N_427);
and U520 (N_520,N_459,N_427);
or U521 (N_521,N_437,N_465);
nand U522 (N_522,N_444,N_458);
or U523 (N_523,N_438,N_439);
nor U524 (N_524,N_430,N_464);
nor U525 (N_525,N_460,N_467);
nand U526 (N_526,N_437,N_464);
nor U527 (N_527,N_464,N_445);
nor U528 (N_528,N_436,N_469);
xor U529 (N_529,N_460,N_424);
xnor U530 (N_530,N_447,N_456);
nor U531 (N_531,N_462,N_456);
or U532 (N_532,N_460,N_453);
nand U533 (N_533,N_430,N_435);
nand U534 (N_534,N_461,N_451);
nand U535 (N_535,N_438,N_478);
or U536 (N_536,N_462,N_439);
or U537 (N_537,N_420,N_476);
nor U538 (N_538,N_449,N_476);
nand U539 (N_539,N_477,N_461);
nor U540 (N_540,N_502,N_520);
nor U541 (N_541,N_523,N_529);
and U542 (N_542,N_498,N_519);
and U543 (N_543,N_482,N_492);
nor U544 (N_544,N_538,N_512);
nand U545 (N_545,N_525,N_531);
or U546 (N_546,N_528,N_522);
xnor U547 (N_547,N_494,N_527);
and U548 (N_548,N_509,N_535);
nor U549 (N_549,N_537,N_485);
nor U550 (N_550,N_514,N_493);
or U551 (N_551,N_488,N_517);
xor U552 (N_552,N_486,N_481);
and U553 (N_553,N_500,N_501);
or U554 (N_554,N_484,N_483);
nand U555 (N_555,N_489,N_480);
nand U556 (N_556,N_504,N_524);
xor U557 (N_557,N_497,N_539);
nand U558 (N_558,N_526,N_532);
nand U559 (N_559,N_518,N_511);
nor U560 (N_560,N_521,N_515);
nand U561 (N_561,N_516,N_513);
xnor U562 (N_562,N_534,N_507);
and U563 (N_563,N_505,N_495);
nand U564 (N_564,N_490,N_496);
nand U565 (N_565,N_499,N_508);
nor U566 (N_566,N_491,N_530);
nor U567 (N_567,N_503,N_536);
or U568 (N_568,N_506,N_533);
xnor U569 (N_569,N_487,N_510);
or U570 (N_570,N_507,N_491);
xnor U571 (N_571,N_486,N_539);
or U572 (N_572,N_521,N_484);
xnor U573 (N_573,N_504,N_487);
or U574 (N_574,N_497,N_503);
and U575 (N_575,N_524,N_499);
nor U576 (N_576,N_502,N_539);
and U577 (N_577,N_504,N_522);
and U578 (N_578,N_495,N_535);
nand U579 (N_579,N_515,N_526);
nor U580 (N_580,N_489,N_482);
nand U581 (N_581,N_529,N_481);
nand U582 (N_582,N_484,N_480);
xor U583 (N_583,N_539,N_531);
nand U584 (N_584,N_494,N_528);
and U585 (N_585,N_502,N_524);
or U586 (N_586,N_490,N_505);
xor U587 (N_587,N_513,N_518);
nand U588 (N_588,N_523,N_491);
and U589 (N_589,N_485,N_490);
nand U590 (N_590,N_516,N_510);
nand U591 (N_591,N_500,N_486);
or U592 (N_592,N_532,N_533);
xor U593 (N_593,N_506,N_528);
xnor U594 (N_594,N_508,N_485);
xor U595 (N_595,N_508,N_534);
or U596 (N_596,N_498,N_535);
or U597 (N_597,N_539,N_524);
nor U598 (N_598,N_535,N_511);
nor U599 (N_599,N_492,N_531);
xnor U600 (N_600,N_561,N_558);
nor U601 (N_601,N_563,N_583);
or U602 (N_602,N_552,N_543);
and U603 (N_603,N_573,N_545);
and U604 (N_604,N_581,N_591);
nand U605 (N_605,N_553,N_575);
or U606 (N_606,N_541,N_571);
xor U607 (N_607,N_579,N_577);
and U608 (N_608,N_549,N_588);
and U609 (N_609,N_594,N_576);
nand U610 (N_610,N_572,N_584);
and U611 (N_611,N_578,N_587);
xnor U612 (N_612,N_568,N_547);
and U613 (N_613,N_570,N_598);
nor U614 (N_614,N_574,N_586);
xor U615 (N_615,N_544,N_592);
nand U616 (N_616,N_567,N_540);
nor U617 (N_617,N_546,N_569);
or U618 (N_618,N_590,N_562);
and U619 (N_619,N_554,N_560);
and U620 (N_620,N_582,N_556);
and U621 (N_621,N_548,N_580);
and U622 (N_622,N_550,N_566);
nor U623 (N_623,N_564,N_559);
and U624 (N_624,N_593,N_585);
nor U625 (N_625,N_565,N_596);
and U626 (N_626,N_599,N_595);
nor U627 (N_627,N_555,N_597);
xnor U628 (N_628,N_557,N_551);
nand U629 (N_629,N_589,N_542);
and U630 (N_630,N_553,N_560);
and U631 (N_631,N_550,N_556);
or U632 (N_632,N_598,N_564);
xor U633 (N_633,N_568,N_543);
nor U634 (N_634,N_583,N_540);
or U635 (N_635,N_599,N_597);
xnor U636 (N_636,N_555,N_591);
nand U637 (N_637,N_556,N_578);
nand U638 (N_638,N_593,N_561);
or U639 (N_639,N_585,N_548);
nand U640 (N_640,N_597,N_556);
xor U641 (N_641,N_587,N_574);
and U642 (N_642,N_548,N_562);
nor U643 (N_643,N_558,N_565);
nor U644 (N_644,N_551,N_544);
nor U645 (N_645,N_593,N_555);
and U646 (N_646,N_570,N_587);
nor U647 (N_647,N_591,N_547);
xnor U648 (N_648,N_566,N_549);
xor U649 (N_649,N_554,N_591);
or U650 (N_650,N_579,N_549);
nor U651 (N_651,N_574,N_575);
and U652 (N_652,N_546,N_580);
xor U653 (N_653,N_570,N_557);
or U654 (N_654,N_563,N_552);
and U655 (N_655,N_587,N_543);
and U656 (N_656,N_581,N_588);
and U657 (N_657,N_598,N_557);
xor U658 (N_658,N_566,N_579);
nand U659 (N_659,N_565,N_587);
nand U660 (N_660,N_632,N_657);
xor U661 (N_661,N_646,N_617);
nor U662 (N_662,N_643,N_620);
or U663 (N_663,N_658,N_653);
xnor U664 (N_664,N_639,N_603);
or U665 (N_665,N_605,N_608);
nand U666 (N_666,N_648,N_638);
xor U667 (N_667,N_629,N_654);
nor U668 (N_668,N_610,N_613);
and U669 (N_669,N_618,N_627);
or U670 (N_670,N_623,N_606);
nand U671 (N_671,N_649,N_607);
or U672 (N_672,N_636,N_650);
nor U673 (N_673,N_626,N_614);
or U674 (N_674,N_656,N_628);
xor U675 (N_675,N_642,N_615);
nor U676 (N_676,N_635,N_619);
and U677 (N_677,N_645,N_602);
nor U678 (N_678,N_634,N_600);
and U679 (N_679,N_601,N_651);
and U680 (N_680,N_630,N_624);
and U681 (N_681,N_647,N_621);
nor U682 (N_682,N_611,N_625);
or U683 (N_683,N_641,N_622);
and U684 (N_684,N_644,N_655);
xnor U685 (N_685,N_640,N_633);
and U686 (N_686,N_631,N_612);
or U687 (N_687,N_637,N_659);
xor U688 (N_688,N_604,N_609);
nor U689 (N_689,N_616,N_652);
nand U690 (N_690,N_650,N_646);
or U691 (N_691,N_653,N_610);
and U692 (N_692,N_642,N_631);
and U693 (N_693,N_653,N_633);
or U694 (N_694,N_622,N_642);
or U695 (N_695,N_631,N_633);
nor U696 (N_696,N_610,N_646);
xnor U697 (N_697,N_604,N_606);
and U698 (N_698,N_649,N_646);
and U699 (N_699,N_625,N_654);
nor U700 (N_700,N_622,N_613);
nor U701 (N_701,N_657,N_620);
xnor U702 (N_702,N_645,N_603);
or U703 (N_703,N_607,N_611);
and U704 (N_704,N_617,N_659);
or U705 (N_705,N_645,N_618);
nor U706 (N_706,N_638,N_613);
xor U707 (N_707,N_628,N_641);
and U708 (N_708,N_608,N_650);
or U709 (N_709,N_609,N_623);
and U710 (N_710,N_656,N_605);
nor U711 (N_711,N_626,N_604);
nand U712 (N_712,N_635,N_610);
nand U713 (N_713,N_606,N_621);
or U714 (N_714,N_621,N_645);
xor U715 (N_715,N_646,N_654);
nor U716 (N_716,N_625,N_620);
xnor U717 (N_717,N_626,N_632);
nand U718 (N_718,N_636,N_621);
nor U719 (N_719,N_613,N_607);
nor U720 (N_720,N_689,N_711);
nand U721 (N_721,N_662,N_668);
and U722 (N_722,N_695,N_715);
nand U723 (N_723,N_660,N_690);
nor U724 (N_724,N_708,N_702);
or U725 (N_725,N_688,N_703);
nand U726 (N_726,N_683,N_704);
and U727 (N_727,N_684,N_710);
nand U728 (N_728,N_693,N_701);
nor U729 (N_729,N_677,N_670);
xnor U730 (N_730,N_681,N_705);
nand U731 (N_731,N_709,N_682);
and U732 (N_732,N_706,N_676);
and U733 (N_733,N_718,N_696);
or U734 (N_734,N_713,N_673);
xor U735 (N_735,N_666,N_719);
nand U736 (N_736,N_672,N_669);
nor U737 (N_737,N_686,N_714);
and U738 (N_738,N_692,N_712);
nand U739 (N_739,N_717,N_678);
and U740 (N_740,N_697,N_716);
or U741 (N_741,N_698,N_707);
or U742 (N_742,N_665,N_661);
and U743 (N_743,N_679,N_664);
and U744 (N_744,N_675,N_663);
nand U745 (N_745,N_680,N_674);
xor U746 (N_746,N_667,N_687);
or U747 (N_747,N_700,N_691);
or U748 (N_748,N_699,N_694);
nor U749 (N_749,N_671,N_685);
nor U750 (N_750,N_660,N_716);
nor U751 (N_751,N_707,N_708);
and U752 (N_752,N_699,N_676);
or U753 (N_753,N_679,N_691);
and U754 (N_754,N_704,N_684);
xnor U755 (N_755,N_712,N_684);
xnor U756 (N_756,N_706,N_674);
nand U757 (N_757,N_662,N_714);
and U758 (N_758,N_677,N_686);
nand U759 (N_759,N_711,N_683);
xnor U760 (N_760,N_662,N_686);
nand U761 (N_761,N_675,N_688);
and U762 (N_762,N_663,N_713);
or U763 (N_763,N_709,N_686);
xor U764 (N_764,N_660,N_717);
or U765 (N_765,N_692,N_695);
nand U766 (N_766,N_709,N_691);
nor U767 (N_767,N_699,N_687);
xor U768 (N_768,N_695,N_675);
or U769 (N_769,N_678,N_714);
and U770 (N_770,N_700,N_660);
nand U771 (N_771,N_687,N_665);
and U772 (N_772,N_706,N_675);
xor U773 (N_773,N_680,N_708);
nand U774 (N_774,N_703,N_661);
xnor U775 (N_775,N_686,N_719);
or U776 (N_776,N_718,N_707);
xnor U777 (N_777,N_701,N_677);
nor U778 (N_778,N_693,N_698);
or U779 (N_779,N_717,N_681);
xnor U780 (N_780,N_749,N_768);
xnor U781 (N_781,N_762,N_772);
or U782 (N_782,N_743,N_742);
xor U783 (N_783,N_758,N_751);
or U784 (N_784,N_741,N_731);
xor U785 (N_785,N_723,N_750);
nor U786 (N_786,N_766,N_767);
nand U787 (N_787,N_771,N_748);
nand U788 (N_788,N_756,N_778);
and U789 (N_789,N_757,N_769);
or U790 (N_790,N_732,N_739);
or U791 (N_791,N_755,N_775);
nand U792 (N_792,N_759,N_738);
and U793 (N_793,N_726,N_720);
and U794 (N_794,N_740,N_752);
xnor U795 (N_795,N_727,N_754);
xor U796 (N_796,N_746,N_736);
nor U797 (N_797,N_765,N_721);
or U798 (N_798,N_735,N_725);
xnor U799 (N_799,N_724,N_770);
nor U800 (N_800,N_774,N_761);
nand U801 (N_801,N_776,N_744);
or U802 (N_802,N_779,N_753);
and U803 (N_803,N_745,N_734);
xor U804 (N_804,N_760,N_773);
and U805 (N_805,N_747,N_777);
xnor U806 (N_806,N_764,N_737);
nand U807 (N_807,N_763,N_728);
xnor U808 (N_808,N_733,N_729);
and U809 (N_809,N_722,N_730);
nand U810 (N_810,N_753,N_758);
or U811 (N_811,N_757,N_740);
and U812 (N_812,N_747,N_743);
xor U813 (N_813,N_727,N_749);
nand U814 (N_814,N_765,N_750);
nand U815 (N_815,N_751,N_720);
nor U816 (N_816,N_766,N_749);
and U817 (N_817,N_777,N_725);
or U818 (N_818,N_777,N_768);
nor U819 (N_819,N_720,N_767);
and U820 (N_820,N_739,N_755);
xnor U821 (N_821,N_723,N_735);
nor U822 (N_822,N_746,N_761);
and U823 (N_823,N_741,N_758);
nor U824 (N_824,N_757,N_775);
or U825 (N_825,N_759,N_748);
nand U826 (N_826,N_773,N_778);
and U827 (N_827,N_752,N_730);
nand U828 (N_828,N_730,N_777);
or U829 (N_829,N_720,N_763);
and U830 (N_830,N_753,N_742);
and U831 (N_831,N_721,N_770);
xor U832 (N_832,N_762,N_771);
xnor U833 (N_833,N_758,N_767);
xor U834 (N_834,N_762,N_779);
or U835 (N_835,N_769,N_749);
nor U836 (N_836,N_764,N_745);
and U837 (N_837,N_764,N_723);
nand U838 (N_838,N_722,N_754);
nand U839 (N_839,N_746,N_763);
nor U840 (N_840,N_792,N_832);
or U841 (N_841,N_816,N_801);
or U842 (N_842,N_824,N_826);
xnor U843 (N_843,N_789,N_833);
nand U844 (N_844,N_784,N_812);
xnor U845 (N_845,N_829,N_796);
xnor U846 (N_846,N_811,N_785);
nand U847 (N_847,N_839,N_825);
and U848 (N_848,N_783,N_787);
nor U849 (N_849,N_813,N_834);
and U850 (N_850,N_800,N_802);
nand U851 (N_851,N_797,N_814);
nor U852 (N_852,N_818,N_805);
nand U853 (N_853,N_804,N_803);
and U854 (N_854,N_809,N_837);
and U855 (N_855,N_831,N_795);
or U856 (N_856,N_791,N_808);
xor U857 (N_857,N_781,N_830);
xnor U858 (N_858,N_819,N_782);
nor U859 (N_859,N_788,N_828);
and U860 (N_860,N_790,N_823);
and U861 (N_861,N_815,N_806);
and U862 (N_862,N_835,N_838);
nor U863 (N_863,N_794,N_780);
nor U864 (N_864,N_820,N_836);
xnor U865 (N_865,N_786,N_810);
and U866 (N_866,N_817,N_827);
and U867 (N_867,N_807,N_793);
or U868 (N_868,N_799,N_821);
nand U869 (N_869,N_798,N_822);
xor U870 (N_870,N_797,N_792);
or U871 (N_871,N_800,N_827);
and U872 (N_872,N_832,N_825);
and U873 (N_873,N_797,N_837);
nand U874 (N_874,N_834,N_803);
or U875 (N_875,N_791,N_805);
or U876 (N_876,N_804,N_797);
and U877 (N_877,N_805,N_822);
nor U878 (N_878,N_835,N_791);
xnor U879 (N_879,N_829,N_788);
and U880 (N_880,N_798,N_783);
xnor U881 (N_881,N_823,N_836);
nor U882 (N_882,N_784,N_814);
or U883 (N_883,N_800,N_833);
xnor U884 (N_884,N_794,N_787);
or U885 (N_885,N_783,N_820);
and U886 (N_886,N_808,N_804);
xnor U887 (N_887,N_795,N_790);
and U888 (N_888,N_837,N_820);
nor U889 (N_889,N_784,N_780);
and U890 (N_890,N_835,N_787);
nand U891 (N_891,N_801,N_793);
nor U892 (N_892,N_783,N_806);
or U893 (N_893,N_798,N_835);
nand U894 (N_894,N_814,N_817);
xor U895 (N_895,N_784,N_809);
and U896 (N_896,N_825,N_814);
xnor U897 (N_897,N_797,N_781);
nor U898 (N_898,N_812,N_787);
nand U899 (N_899,N_815,N_790);
xor U900 (N_900,N_847,N_897);
or U901 (N_901,N_854,N_888);
or U902 (N_902,N_845,N_846);
nor U903 (N_903,N_883,N_859);
nand U904 (N_904,N_844,N_873);
nand U905 (N_905,N_877,N_858);
nor U906 (N_906,N_841,N_868);
nor U907 (N_907,N_887,N_867);
or U908 (N_908,N_857,N_885);
nand U909 (N_909,N_860,N_892);
and U910 (N_910,N_842,N_886);
nand U911 (N_911,N_889,N_849);
and U912 (N_912,N_865,N_862);
and U913 (N_913,N_855,N_894);
and U914 (N_914,N_851,N_856);
nor U915 (N_915,N_881,N_874);
or U916 (N_916,N_890,N_848);
and U917 (N_917,N_863,N_896);
xor U918 (N_918,N_875,N_869);
or U919 (N_919,N_871,N_872);
nor U920 (N_920,N_853,N_870);
xnor U921 (N_921,N_899,N_843);
nor U922 (N_922,N_895,N_882);
nor U923 (N_923,N_878,N_866);
xnor U924 (N_924,N_884,N_879);
or U925 (N_925,N_861,N_880);
nand U926 (N_926,N_852,N_891);
nand U927 (N_927,N_864,N_898);
or U928 (N_928,N_893,N_840);
xor U929 (N_929,N_876,N_850);
xnor U930 (N_930,N_857,N_868);
nand U931 (N_931,N_843,N_889);
nor U932 (N_932,N_849,N_844);
xor U933 (N_933,N_840,N_881);
nor U934 (N_934,N_881,N_852);
nor U935 (N_935,N_869,N_861);
nand U936 (N_936,N_896,N_840);
and U937 (N_937,N_882,N_862);
and U938 (N_938,N_898,N_895);
nand U939 (N_939,N_885,N_845);
nand U940 (N_940,N_886,N_880);
xnor U941 (N_941,N_872,N_840);
or U942 (N_942,N_881,N_879);
or U943 (N_943,N_880,N_876);
or U944 (N_944,N_845,N_873);
nor U945 (N_945,N_854,N_899);
or U946 (N_946,N_881,N_871);
and U947 (N_947,N_880,N_841);
nor U948 (N_948,N_853,N_855);
nor U949 (N_949,N_850,N_886);
nand U950 (N_950,N_849,N_881);
xor U951 (N_951,N_899,N_882);
or U952 (N_952,N_845,N_878);
nor U953 (N_953,N_840,N_869);
or U954 (N_954,N_877,N_856);
and U955 (N_955,N_844,N_862);
nand U956 (N_956,N_885,N_869);
and U957 (N_957,N_889,N_896);
nand U958 (N_958,N_879,N_848);
and U959 (N_959,N_845,N_877);
xor U960 (N_960,N_929,N_910);
and U961 (N_961,N_947,N_954);
nor U962 (N_962,N_911,N_923);
nor U963 (N_963,N_956,N_926);
nand U964 (N_964,N_914,N_953);
nand U965 (N_965,N_915,N_925);
xnor U966 (N_966,N_957,N_904);
and U967 (N_967,N_935,N_934);
nor U968 (N_968,N_931,N_941);
nor U969 (N_969,N_959,N_903);
or U970 (N_970,N_950,N_908);
or U971 (N_971,N_939,N_919);
xor U972 (N_972,N_940,N_955);
and U973 (N_973,N_949,N_937);
or U974 (N_974,N_921,N_906);
and U975 (N_975,N_924,N_952);
and U976 (N_976,N_951,N_912);
nor U977 (N_977,N_930,N_902);
nand U978 (N_978,N_913,N_900);
or U979 (N_979,N_945,N_933);
xor U980 (N_980,N_943,N_938);
xor U981 (N_981,N_928,N_936);
and U982 (N_982,N_948,N_916);
nor U983 (N_983,N_927,N_917);
nand U984 (N_984,N_922,N_946);
and U985 (N_985,N_942,N_932);
nand U986 (N_986,N_907,N_918);
xor U987 (N_987,N_920,N_901);
nor U988 (N_988,N_905,N_944);
xor U989 (N_989,N_909,N_958);
or U990 (N_990,N_936,N_906);
or U991 (N_991,N_924,N_915);
and U992 (N_992,N_944,N_952);
nand U993 (N_993,N_940,N_958);
nand U994 (N_994,N_903,N_948);
or U995 (N_995,N_924,N_946);
nand U996 (N_996,N_949,N_911);
nor U997 (N_997,N_927,N_919);
nand U998 (N_998,N_926,N_943);
nor U999 (N_999,N_934,N_921);
and U1000 (N_1000,N_929,N_903);
and U1001 (N_1001,N_954,N_913);
nand U1002 (N_1002,N_916,N_915);
xor U1003 (N_1003,N_921,N_936);
or U1004 (N_1004,N_954,N_934);
nand U1005 (N_1005,N_952,N_927);
nor U1006 (N_1006,N_942,N_950);
or U1007 (N_1007,N_951,N_906);
nand U1008 (N_1008,N_924,N_901);
nor U1009 (N_1009,N_949,N_914);
and U1010 (N_1010,N_902,N_943);
nor U1011 (N_1011,N_904,N_930);
or U1012 (N_1012,N_940,N_951);
nand U1013 (N_1013,N_906,N_916);
nor U1014 (N_1014,N_929,N_955);
xor U1015 (N_1015,N_952,N_905);
nor U1016 (N_1016,N_921,N_920);
nor U1017 (N_1017,N_957,N_959);
xnor U1018 (N_1018,N_944,N_903);
xor U1019 (N_1019,N_916,N_918);
or U1020 (N_1020,N_1016,N_1006);
nor U1021 (N_1021,N_971,N_997);
nor U1022 (N_1022,N_1007,N_964);
xor U1023 (N_1023,N_995,N_990);
nor U1024 (N_1024,N_996,N_998);
xor U1025 (N_1025,N_1015,N_993);
and U1026 (N_1026,N_1014,N_962);
nand U1027 (N_1027,N_979,N_999);
and U1028 (N_1028,N_1017,N_1011);
nand U1029 (N_1029,N_985,N_987);
nor U1030 (N_1030,N_1010,N_961);
xnor U1031 (N_1031,N_994,N_1008);
and U1032 (N_1032,N_982,N_991);
or U1033 (N_1033,N_972,N_1009);
and U1034 (N_1034,N_960,N_1013);
xnor U1035 (N_1035,N_989,N_980);
xnor U1036 (N_1036,N_992,N_1019);
and U1037 (N_1037,N_1001,N_981);
nor U1038 (N_1038,N_988,N_975);
nor U1039 (N_1039,N_965,N_1002);
or U1040 (N_1040,N_1018,N_970);
nand U1041 (N_1041,N_1012,N_974);
nand U1042 (N_1042,N_978,N_968);
and U1043 (N_1043,N_976,N_1003);
nor U1044 (N_1044,N_1000,N_967);
nand U1045 (N_1045,N_969,N_983);
nand U1046 (N_1046,N_1004,N_984);
nand U1047 (N_1047,N_973,N_966);
or U1048 (N_1048,N_963,N_986);
xor U1049 (N_1049,N_977,N_1005);
and U1050 (N_1050,N_964,N_1005);
and U1051 (N_1051,N_970,N_995);
and U1052 (N_1052,N_1009,N_1010);
nand U1053 (N_1053,N_994,N_1010);
nor U1054 (N_1054,N_989,N_987);
nor U1055 (N_1055,N_1000,N_989);
or U1056 (N_1056,N_1009,N_983);
nand U1057 (N_1057,N_979,N_1004);
nor U1058 (N_1058,N_995,N_997);
xnor U1059 (N_1059,N_990,N_986);
nand U1060 (N_1060,N_981,N_973);
nor U1061 (N_1061,N_962,N_982);
and U1062 (N_1062,N_991,N_986);
and U1063 (N_1063,N_993,N_1016);
nand U1064 (N_1064,N_970,N_1004);
nand U1065 (N_1065,N_1003,N_1012);
xnor U1066 (N_1066,N_1001,N_985);
nor U1067 (N_1067,N_987,N_1018);
nor U1068 (N_1068,N_991,N_981);
or U1069 (N_1069,N_998,N_1009);
nor U1070 (N_1070,N_968,N_982);
nor U1071 (N_1071,N_1011,N_1013);
nand U1072 (N_1072,N_1015,N_998);
nand U1073 (N_1073,N_980,N_974);
xor U1074 (N_1074,N_969,N_971);
and U1075 (N_1075,N_977,N_963);
or U1076 (N_1076,N_989,N_993);
nand U1077 (N_1077,N_965,N_1018);
xor U1078 (N_1078,N_1011,N_1001);
or U1079 (N_1079,N_982,N_1019);
or U1080 (N_1080,N_1071,N_1061);
nor U1081 (N_1081,N_1047,N_1052);
and U1082 (N_1082,N_1073,N_1022);
xnor U1083 (N_1083,N_1027,N_1036);
or U1084 (N_1084,N_1032,N_1056);
nor U1085 (N_1085,N_1028,N_1063);
or U1086 (N_1086,N_1023,N_1029);
xnor U1087 (N_1087,N_1045,N_1039);
and U1088 (N_1088,N_1079,N_1026);
or U1089 (N_1089,N_1078,N_1030);
nor U1090 (N_1090,N_1051,N_1066);
nor U1091 (N_1091,N_1062,N_1037);
nor U1092 (N_1092,N_1049,N_1074);
and U1093 (N_1093,N_1058,N_1053);
xnor U1094 (N_1094,N_1064,N_1059);
xor U1095 (N_1095,N_1033,N_1025);
nand U1096 (N_1096,N_1043,N_1067);
nand U1097 (N_1097,N_1034,N_1072);
nand U1098 (N_1098,N_1060,N_1075);
and U1099 (N_1099,N_1070,N_1031);
and U1100 (N_1100,N_1044,N_1041);
nor U1101 (N_1101,N_1050,N_1077);
nor U1102 (N_1102,N_1057,N_1069);
or U1103 (N_1103,N_1021,N_1035);
and U1104 (N_1104,N_1065,N_1076);
xor U1105 (N_1105,N_1038,N_1048);
nor U1106 (N_1106,N_1046,N_1024);
xnor U1107 (N_1107,N_1068,N_1055);
nand U1108 (N_1108,N_1042,N_1054);
and U1109 (N_1109,N_1040,N_1020);
nor U1110 (N_1110,N_1048,N_1051);
nor U1111 (N_1111,N_1029,N_1021);
xnor U1112 (N_1112,N_1056,N_1039);
nand U1113 (N_1113,N_1072,N_1060);
and U1114 (N_1114,N_1038,N_1067);
xnor U1115 (N_1115,N_1033,N_1026);
nand U1116 (N_1116,N_1029,N_1064);
and U1117 (N_1117,N_1078,N_1055);
nand U1118 (N_1118,N_1031,N_1077);
or U1119 (N_1119,N_1020,N_1028);
and U1120 (N_1120,N_1025,N_1021);
nor U1121 (N_1121,N_1028,N_1070);
nor U1122 (N_1122,N_1067,N_1030);
nand U1123 (N_1123,N_1065,N_1026);
xnor U1124 (N_1124,N_1048,N_1037);
or U1125 (N_1125,N_1065,N_1046);
xnor U1126 (N_1126,N_1042,N_1069);
xnor U1127 (N_1127,N_1044,N_1021);
xnor U1128 (N_1128,N_1068,N_1063);
and U1129 (N_1129,N_1070,N_1025);
and U1130 (N_1130,N_1020,N_1071);
xor U1131 (N_1131,N_1063,N_1066);
or U1132 (N_1132,N_1044,N_1042);
nor U1133 (N_1133,N_1059,N_1022);
nor U1134 (N_1134,N_1055,N_1065);
nor U1135 (N_1135,N_1033,N_1050);
nor U1136 (N_1136,N_1028,N_1037);
nand U1137 (N_1137,N_1037,N_1029);
or U1138 (N_1138,N_1077,N_1055);
xnor U1139 (N_1139,N_1030,N_1051);
or U1140 (N_1140,N_1120,N_1092);
or U1141 (N_1141,N_1081,N_1137);
and U1142 (N_1142,N_1087,N_1112);
nand U1143 (N_1143,N_1096,N_1098);
and U1144 (N_1144,N_1116,N_1095);
xor U1145 (N_1145,N_1136,N_1097);
and U1146 (N_1146,N_1089,N_1090);
or U1147 (N_1147,N_1086,N_1080);
and U1148 (N_1148,N_1102,N_1129);
or U1149 (N_1149,N_1133,N_1131);
or U1150 (N_1150,N_1106,N_1093);
nand U1151 (N_1151,N_1099,N_1117);
or U1152 (N_1152,N_1108,N_1082);
or U1153 (N_1153,N_1119,N_1113);
or U1154 (N_1154,N_1115,N_1083);
xnor U1155 (N_1155,N_1094,N_1128);
and U1156 (N_1156,N_1104,N_1139);
or U1157 (N_1157,N_1123,N_1101);
xnor U1158 (N_1158,N_1132,N_1103);
nor U1159 (N_1159,N_1135,N_1121);
nand U1160 (N_1160,N_1107,N_1088);
or U1161 (N_1161,N_1084,N_1122);
nor U1162 (N_1162,N_1134,N_1126);
xor U1163 (N_1163,N_1091,N_1105);
or U1164 (N_1164,N_1114,N_1138);
nand U1165 (N_1165,N_1111,N_1130);
xnor U1166 (N_1166,N_1127,N_1125);
nand U1167 (N_1167,N_1109,N_1110);
xnor U1168 (N_1168,N_1100,N_1085);
and U1169 (N_1169,N_1124,N_1118);
nor U1170 (N_1170,N_1132,N_1108);
nor U1171 (N_1171,N_1088,N_1122);
and U1172 (N_1172,N_1134,N_1097);
nor U1173 (N_1173,N_1093,N_1088);
xor U1174 (N_1174,N_1109,N_1139);
or U1175 (N_1175,N_1117,N_1107);
nor U1176 (N_1176,N_1104,N_1117);
nor U1177 (N_1177,N_1120,N_1106);
nor U1178 (N_1178,N_1098,N_1125);
nor U1179 (N_1179,N_1120,N_1094);
or U1180 (N_1180,N_1127,N_1129);
and U1181 (N_1181,N_1128,N_1092);
and U1182 (N_1182,N_1089,N_1106);
and U1183 (N_1183,N_1095,N_1137);
nand U1184 (N_1184,N_1119,N_1087);
and U1185 (N_1185,N_1123,N_1136);
xor U1186 (N_1186,N_1114,N_1106);
nor U1187 (N_1187,N_1118,N_1088);
nor U1188 (N_1188,N_1098,N_1134);
nor U1189 (N_1189,N_1088,N_1123);
or U1190 (N_1190,N_1111,N_1087);
and U1191 (N_1191,N_1085,N_1094);
nor U1192 (N_1192,N_1084,N_1118);
or U1193 (N_1193,N_1086,N_1129);
nor U1194 (N_1194,N_1099,N_1125);
nor U1195 (N_1195,N_1132,N_1128);
nand U1196 (N_1196,N_1102,N_1088);
or U1197 (N_1197,N_1087,N_1127);
xnor U1198 (N_1198,N_1104,N_1124);
nand U1199 (N_1199,N_1129,N_1107);
or U1200 (N_1200,N_1143,N_1150);
or U1201 (N_1201,N_1175,N_1179);
nor U1202 (N_1202,N_1148,N_1185);
xor U1203 (N_1203,N_1162,N_1161);
nor U1204 (N_1204,N_1173,N_1169);
nand U1205 (N_1205,N_1168,N_1198);
or U1206 (N_1206,N_1191,N_1140);
xnor U1207 (N_1207,N_1172,N_1153);
and U1208 (N_1208,N_1186,N_1194);
xor U1209 (N_1209,N_1157,N_1199);
and U1210 (N_1210,N_1151,N_1189);
xor U1211 (N_1211,N_1171,N_1178);
nand U1212 (N_1212,N_1197,N_1166);
and U1213 (N_1213,N_1159,N_1180);
or U1214 (N_1214,N_1184,N_1156);
xnor U1215 (N_1215,N_1158,N_1149);
or U1216 (N_1216,N_1190,N_1155);
nor U1217 (N_1217,N_1182,N_1174);
nand U1218 (N_1218,N_1163,N_1145);
nor U1219 (N_1219,N_1141,N_1165);
or U1220 (N_1220,N_1187,N_1147);
nand U1221 (N_1221,N_1146,N_1160);
or U1222 (N_1222,N_1181,N_1144);
nand U1223 (N_1223,N_1176,N_1188);
and U1224 (N_1224,N_1152,N_1154);
and U1225 (N_1225,N_1193,N_1167);
or U1226 (N_1226,N_1164,N_1192);
nor U1227 (N_1227,N_1196,N_1183);
xor U1228 (N_1228,N_1195,N_1177);
nand U1229 (N_1229,N_1170,N_1142);
xor U1230 (N_1230,N_1165,N_1168);
nor U1231 (N_1231,N_1183,N_1164);
or U1232 (N_1232,N_1166,N_1199);
or U1233 (N_1233,N_1163,N_1187);
or U1234 (N_1234,N_1147,N_1197);
xor U1235 (N_1235,N_1183,N_1140);
nand U1236 (N_1236,N_1150,N_1160);
nor U1237 (N_1237,N_1181,N_1178);
and U1238 (N_1238,N_1198,N_1176);
or U1239 (N_1239,N_1161,N_1177);
nor U1240 (N_1240,N_1146,N_1193);
and U1241 (N_1241,N_1155,N_1177);
xnor U1242 (N_1242,N_1187,N_1186);
nor U1243 (N_1243,N_1180,N_1146);
xnor U1244 (N_1244,N_1153,N_1197);
nand U1245 (N_1245,N_1172,N_1189);
xnor U1246 (N_1246,N_1190,N_1141);
nand U1247 (N_1247,N_1180,N_1142);
nor U1248 (N_1248,N_1144,N_1192);
and U1249 (N_1249,N_1142,N_1199);
xnor U1250 (N_1250,N_1149,N_1165);
nand U1251 (N_1251,N_1145,N_1150);
nor U1252 (N_1252,N_1199,N_1172);
or U1253 (N_1253,N_1162,N_1177);
and U1254 (N_1254,N_1167,N_1159);
and U1255 (N_1255,N_1180,N_1194);
xor U1256 (N_1256,N_1174,N_1146);
or U1257 (N_1257,N_1169,N_1194);
xnor U1258 (N_1258,N_1169,N_1149);
xor U1259 (N_1259,N_1196,N_1190);
nand U1260 (N_1260,N_1251,N_1248);
xor U1261 (N_1261,N_1244,N_1213);
or U1262 (N_1262,N_1235,N_1229);
and U1263 (N_1263,N_1258,N_1204);
nand U1264 (N_1264,N_1205,N_1200);
nand U1265 (N_1265,N_1259,N_1253);
or U1266 (N_1266,N_1233,N_1246);
or U1267 (N_1267,N_1236,N_1241);
or U1268 (N_1268,N_1218,N_1247);
xnor U1269 (N_1269,N_1223,N_1219);
nand U1270 (N_1270,N_1227,N_1255);
nand U1271 (N_1271,N_1254,N_1217);
or U1272 (N_1272,N_1203,N_1221);
and U1273 (N_1273,N_1222,N_1225);
nand U1274 (N_1274,N_1206,N_1228);
or U1275 (N_1275,N_1202,N_1207);
xnor U1276 (N_1276,N_1210,N_1256);
xnor U1277 (N_1277,N_1215,N_1250);
or U1278 (N_1278,N_1242,N_1245);
nand U1279 (N_1279,N_1237,N_1214);
nor U1280 (N_1280,N_1232,N_1211);
or U1281 (N_1281,N_1234,N_1226);
nor U1282 (N_1282,N_1224,N_1238);
nand U1283 (N_1283,N_1230,N_1252);
nor U1284 (N_1284,N_1240,N_1239);
xor U1285 (N_1285,N_1208,N_1231);
or U1286 (N_1286,N_1216,N_1220);
or U1287 (N_1287,N_1201,N_1209);
nand U1288 (N_1288,N_1243,N_1257);
xor U1289 (N_1289,N_1249,N_1212);
nand U1290 (N_1290,N_1246,N_1227);
xnor U1291 (N_1291,N_1255,N_1252);
or U1292 (N_1292,N_1246,N_1202);
nand U1293 (N_1293,N_1215,N_1213);
nand U1294 (N_1294,N_1239,N_1214);
nand U1295 (N_1295,N_1237,N_1251);
or U1296 (N_1296,N_1234,N_1235);
or U1297 (N_1297,N_1257,N_1215);
nor U1298 (N_1298,N_1248,N_1255);
nand U1299 (N_1299,N_1207,N_1232);
nand U1300 (N_1300,N_1244,N_1209);
or U1301 (N_1301,N_1238,N_1244);
or U1302 (N_1302,N_1218,N_1205);
and U1303 (N_1303,N_1205,N_1252);
xnor U1304 (N_1304,N_1205,N_1237);
and U1305 (N_1305,N_1222,N_1226);
nor U1306 (N_1306,N_1212,N_1246);
and U1307 (N_1307,N_1225,N_1232);
and U1308 (N_1308,N_1222,N_1208);
or U1309 (N_1309,N_1219,N_1220);
or U1310 (N_1310,N_1244,N_1250);
nor U1311 (N_1311,N_1216,N_1228);
or U1312 (N_1312,N_1244,N_1253);
and U1313 (N_1313,N_1220,N_1207);
or U1314 (N_1314,N_1204,N_1229);
nor U1315 (N_1315,N_1252,N_1254);
xnor U1316 (N_1316,N_1242,N_1240);
nand U1317 (N_1317,N_1251,N_1235);
xnor U1318 (N_1318,N_1229,N_1255);
xor U1319 (N_1319,N_1234,N_1216);
xnor U1320 (N_1320,N_1312,N_1277);
and U1321 (N_1321,N_1317,N_1286);
nand U1322 (N_1322,N_1267,N_1301);
and U1323 (N_1323,N_1290,N_1319);
nor U1324 (N_1324,N_1306,N_1272);
nand U1325 (N_1325,N_1310,N_1316);
nand U1326 (N_1326,N_1289,N_1307);
nand U1327 (N_1327,N_1268,N_1287);
xor U1328 (N_1328,N_1271,N_1280);
xor U1329 (N_1329,N_1284,N_1302);
nor U1330 (N_1330,N_1288,N_1283);
nand U1331 (N_1331,N_1295,N_1314);
xnor U1332 (N_1332,N_1273,N_1260);
nor U1333 (N_1333,N_1276,N_1298);
and U1334 (N_1334,N_1297,N_1270);
nand U1335 (N_1335,N_1305,N_1285);
and U1336 (N_1336,N_1269,N_1278);
nand U1337 (N_1337,N_1261,N_1282);
nor U1338 (N_1338,N_1264,N_1315);
nor U1339 (N_1339,N_1275,N_1318);
nor U1340 (N_1340,N_1303,N_1262);
nand U1341 (N_1341,N_1309,N_1281);
xor U1342 (N_1342,N_1291,N_1292);
or U1343 (N_1343,N_1294,N_1279);
xor U1344 (N_1344,N_1266,N_1311);
and U1345 (N_1345,N_1263,N_1313);
xor U1346 (N_1346,N_1299,N_1300);
or U1347 (N_1347,N_1274,N_1265);
or U1348 (N_1348,N_1293,N_1304);
nor U1349 (N_1349,N_1296,N_1308);
nor U1350 (N_1350,N_1291,N_1280);
nor U1351 (N_1351,N_1307,N_1291);
or U1352 (N_1352,N_1262,N_1270);
and U1353 (N_1353,N_1262,N_1305);
or U1354 (N_1354,N_1283,N_1297);
nor U1355 (N_1355,N_1279,N_1285);
and U1356 (N_1356,N_1299,N_1281);
nor U1357 (N_1357,N_1319,N_1273);
nor U1358 (N_1358,N_1302,N_1264);
xnor U1359 (N_1359,N_1317,N_1268);
nand U1360 (N_1360,N_1277,N_1294);
nand U1361 (N_1361,N_1297,N_1316);
xnor U1362 (N_1362,N_1289,N_1299);
nand U1363 (N_1363,N_1313,N_1270);
xnor U1364 (N_1364,N_1319,N_1303);
nor U1365 (N_1365,N_1269,N_1316);
and U1366 (N_1366,N_1312,N_1303);
xnor U1367 (N_1367,N_1281,N_1285);
or U1368 (N_1368,N_1293,N_1262);
nand U1369 (N_1369,N_1272,N_1316);
nand U1370 (N_1370,N_1303,N_1281);
and U1371 (N_1371,N_1301,N_1317);
xnor U1372 (N_1372,N_1306,N_1260);
and U1373 (N_1373,N_1312,N_1278);
nor U1374 (N_1374,N_1283,N_1273);
xor U1375 (N_1375,N_1288,N_1296);
or U1376 (N_1376,N_1281,N_1287);
nor U1377 (N_1377,N_1264,N_1265);
or U1378 (N_1378,N_1306,N_1288);
and U1379 (N_1379,N_1285,N_1308);
xor U1380 (N_1380,N_1364,N_1348);
and U1381 (N_1381,N_1325,N_1322);
or U1382 (N_1382,N_1343,N_1326);
nand U1383 (N_1383,N_1356,N_1353);
and U1384 (N_1384,N_1369,N_1354);
xor U1385 (N_1385,N_1320,N_1344);
nor U1386 (N_1386,N_1361,N_1335);
nor U1387 (N_1387,N_1345,N_1355);
and U1388 (N_1388,N_1372,N_1370);
xnor U1389 (N_1389,N_1330,N_1346);
or U1390 (N_1390,N_1349,N_1332);
xnor U1391 (N_1391,N_1340,N_1378);
xor U1392 (N_1392,N_1352,N_1360);
xnor U1393 (N_1393,N_1337,N_1347);
nand U1394 (N_1394,N_1365,N_1321);
nand U1395 (N_1395,N_1375,N_1367);
or U1396 (N_1396,N_1363,N_1351);
nor U1397 (N_1397,N_1376,N_1331);
nor U1398 (N_1398,N_1373,N_1368);
nand U1399 (N_1399,N_1359,N_1333);
nor U1400 (N_1400,N_1327,N_1377);
nand U1401 (N_1401,N_1323,N_1336);
xor U1402 (N_1402,N_1362,N_1374);
and U1403 (N_1403,N_1328,N_1324);
nor U1404 (N_1404,N_1366,N_1350);
nand U1405 (N_1405,N_1334,N_1329);
nand U1406 (N_1406,N_1342,N_1357);
or U1407 (N_1407,N_1338,N_1379);
nor U1408 (N_1408,N_1371,N_1341);
nor U1409 (N_1409,N_1339,N_1358);
and U1410 (N_1410,N_1339,N_1355);
nor U1411 (N_1411,N_1330,N_1342);
nand U1412 (N_1412,N_1336,N_1350);
and U1413 (N_1413,N_1338,N_1331);
and U1414 (N_1414,N_1326,N_1371);
nand U1415 (N_1415,N_1334,N_1378);
or U1416 (N_1416,N_1377,N_1329);
xnor U1417 (N_1417,N_1332,N_1374);
xor U1418 (N_1418,N_1371,N_1368);
nor U1419 (N_1419,N_1363,N_1369);
xor U1420 (N_1420,N_1338,N_1324);
and U1421 (N_1421,N_1375,N_1348);
or U1422 (N_1422,N_1365,N_1375);
xor U1423 (N_1423,N_1349,N_1366);
or U1424 (N_1424,N_1356,N_1352);
xnor U1425 (N_1425,N_1338,N_1352);
or U1426 (N_1426,N_1338,N_1372);
nand U1427 (N_1427,N_1362,N_1358);
xor U1428 (N_1428,N_1364,N_1355);
xor U1429 (N_1429,N_1348,N_1365);
or U1430 (N_1430,N_1337,N_1322);
xnor U1431 (N_1431,N_1359,N_1351);
nand U1432 (N_1432,N_1321,N_1359);
and U1433 (N_1433,N_1369,N_1340);
xor U1434 (N_1434,N_1343,N_1344);
and U1435 (N_1435,N_1326,N_1333);
or U1436 (N_1436,N_1353,N_1354);
and U1437 (N_1437,N_1376,N_1357);
xnor U1438 (N_1438,N_1369,N_1373);
xor U1439 (N_1439,N_1355,N_1349);
xnor U1440 (N_1440,N_1410,N_1391);
and U1441 (N_1441,N_1401,N_1390);
xor U1442 (N_1442,N_1432,N_1411);
xor U1443 (N_1443,N_1397,N_1439);
nand U1444 (N_1444,N_1400,N_1394);
and U1445 (N_1445,N_1438,N_1398);
xor U1446 (N_1446,N_1429,N_1393);
xnor U1447 (N_1447,N_1419,N_1430);
xor U1448 (N_1448,N_1396,N_1431);
nand U1449 (N_1449,N_1381,N_1406);
xor U1450 (N_1450,N_1412,N_1437);
nand U1451 (N_1451,N_1428,N_1424);
or U1452 (N_1452,N_1414,N_1409);
and U1453 (N_1453,N_1385,N_1402);
nand U1454 (N_1454,N_1380,N_1416);
and U1455 (N_1455,N_1404,N_1382);
and U1456 (N_1456,N_1415,N_1434);
nand U1457 (N_1457,N_1425,N_1427);
nor U1458 (N_1458,N_1405,N_1433);
nor U1459 (N_1459,N_1383,N_1421);
or U1460 (N_1460,N_1388,N_1392);
nor U1461 (N_1461,N_1436,N_1423);
nor U1462 (N_1462,N_1389,N_1407);
or U1463 (N_1463,N_1387,N_1420);
nor U1464 (N_1464,N_1422,N_1426);
nand U1465 (N_1465,N_1418,N_1399);
nand U1466 (N_1466,N_1408,N_1413);
and U1467 (N_1467,N_1435,N_1386);
xor U1468 (N_1468,N_1384,N_1403);
xor U1469 (N_1469,N_1417,N_1395);
xor U1470 (N_1470,N_1381,N_1434);
xnor U1471 (N_1471,N_1392,N_1419);
nand U1472 (N_1472,N_1403,N_1422);
xor U1473 (N_1473,N_1408,N_1415);
nand U1474 (N_1474,N_1431,N_1392);
or U1475 (N_1475,N_1428,N_1413);
or U1476 (N_1476,N_1402,N_1399);
nor U1477 (N_1477,N_1413,N_1393);
or U1478 (N_1478,N_1403,N_1433);
nand U1479 (N_1479,N_1415,N_1428);
or U1480 (N_1480,N_1402,N_1394);
nor U1481 (N_1481,N_1418,N_1402);
and U1482 (N_1482,N_1397,N_1433);
or U1483 (N_1483,N_1422,N_1439);
or U1484 (N_1484,N_1430,N_1439);
nand U1485 (N_1485,N_1396,N_1388);
nor U1486 (N_1486,N_1432,N_1395);
and U1487 (N_1487,N_1419,N_1424);
and U1488 (N_1488,N_1436,N_1394);
nor U1489 (N_1489,N_1427,N_1382);
nor U1490 (N_1490,N_1414,N_1438);
nand U1491 (N_1491,N_1403,N_1392);
nand U1492 (N_1492,N_1413,N_1426);
and U1493 (N_1493,N_1439,N_1410);
nor U1494 (N_1494,N_1387,N_1427);
nor U1495 (N_1495,N_1388,N_1384);
and U1496 (N_1496,N_1393,N_1384);
nand U1497 (N_1497,N_1414,N_1408);
xnor U1498 (N_1498,N_1426,N_1382);
or U1499 (N_1499,N_1400,N_1427);
nor U1500 (N_1500,N_1496,N_1479);
xor U1501 (N_1501,N_1492,N_1497);
and U1502 (N_1502,N_1440,N_1477);
nor U1503 (N_1503,N_1453,N_1470);
nor U1504 (N_1504,N_1490,N_1484);
nand U1505 (N_1505,N_1494,N_1459);
xor U1506 (N_1506,N_1476,N_1473);
or U1507 (N_1507,N_1474,N_1461);
xnor U1508 (N_1508,N_1451,N_1485);
nand U1509 (N_1509,N_1462,N_1463);
nand U1510 (N_1510,N_1450,N_1493);
or U1511 (N_1511,N_1442,N_1452);
or U1512 (N_1512,N_1458,N_1481);
xnor U1513 (N_1513,N_1469,N_1489);
xor U1514 (N_1514,N_1471,N_1454);
or U1515 (N_1515,N_1483,N_1447);
or U1516 (N_1516,N_1441,N_1468);
and U1517 (N_1517,N_1443,N_1460);
nor U1518 (N_1518,N_1475,N_1449);
and U1519 (N_1519,N_1448,N_1482);
nor U1520 (N_1520,N_1495,N_1486);
nor U1521 (N_1521,N_1456,N_1472);
nor U1522 (N_1522,N_1464,N_1499);
or U1523 (N_1523,N_1445,N_1480);
nand U1524 (N_1524,N_1457,N_1498);
and U1525 (N_1525,N_1467,N_1444);
or U1526 (N_1526,N_1478,N_1446);
xor U1527 (N_1527,N_1487,N_1466);
nor U1528 (N_1528,N_1488,N_1465);
nand U1529 (N_1529,N_1491,N_1455);
xor U1530 (N_1530,N_1475,N_1466);
or U1531 (N_1531,N_1450,N_1490);
xnor U1532 (N_1532,N_1462,N_1484);
and U1533 (N_1533,N_1464,N_1456);
nor U1534 (N_1534,N_1481,N_1457);
and U1535 (N_1535,N_1478,N_1494);
xnor U1536 (N_1536,N_1444,N_1441);
nor U1537 (N_1537,N_1451,N_1484);
nor U1538 (N_1538,N_1489,N_1483);
or U1539 (N_1539,N_1466,N_1459);
nor U1540 (N_1540,N_1462,N_1477);
xnor U1541 (N_1541,N_1499,N_1473);
xnor U1542 (N_1542,N_1441,N_1455);
or U1543 (N_1543,N_1452,N_1490);
nor U1544 (N_1544,N_1465,N_1475);
and U1545 (N_1545,N_1496,N_1480);
nor U1546 (N_1546,N_1483,N_1454);
or U1547 (N_1547,N_1488,N_1457);
nand U1548 (N_1548,N_1487,N_1494);
nand U1549 (N_1549,N_1493,N_1471);
nor U1550 (N_1550,N_1482,N_1477);
and U1551 (N_1551,N_1457,N_1466);
nor U1552 (N_1552,N_1468,N_1447);
nor U1553 (N_1553,N_1454,N_1453);
and U1554 (N_1554,N_1456,N_1482);
nor U1555 (N_1555,N_1480,N_1465);
and U1556 (N_1556,N_1456,N_1462);
nor U1557 (N_1557,N_1446,N_1494);
nor U1558 (N_1558,N_1494,N_1443);
nand U1559 (N_1559,N_1463,N_1497);
nand U1560 (N_1560,N_1528,N_1510);
and U1561 (N_1561,N_1519,N_1500);
nor U1562 (N_1562,N_1538,N_1545);
and U1563 (N_1563,N_1516,N_1534);
nor U1564 (N_1564,N_1509,N_1546);
nor U1565 (N_1565,N_1548,N_1541);
nor U1566 (N_1566,N_1524,N_1557);
and U1567 (N_1567,N_1540,N_1523);
nor U1568 (N_1568,N_1549,N_1556);
and U1569 (N_1569,N_1552,N_1535);
and U1570 (N_1570,N_1505,N_1507);
nand U1571 (N_1571,N_1544,N_1512);
or U1572 (N_1572,N_1543,N_1514);
xor U1573 (N_1573,N_1547,N_1526);
or U1574 (N_1574,N_1517,N_1522);
xor U1575 (N_1575,N_1530,N_1532);
nand U1576 (N_1576,N_1529,N_1515);
or U1577 (N_1577,N_1555,N_1525);
xnor U1578 (N_1578,N_1542,N_1527);
nor U1579 (N_1579,N_1536,N_1539);
or U1580 (N_1580,N_1531,N_1513);
xnor U1581 (N_1581,N_1504,N_1559);
xor U1582 (N_1582,N_1511,N_1521);
nand U1583 (N_1583,N_1533,N_1506);
or U1584 (N_1584,N_1550,N_1518);
and U1585 (N_1585,N_1537,N_1508);
nor U1586 (N_1586,N_1558,N_1503);
and U1587 (N_1587,N_1553,N_1554);
nand U1588 (N_1588,N_1501,N_1520);
and U1589 (N_1589,N_1551,N_1502);
or U1590 (N_1590,N_1551,N_1515);
nand U1591 (N_1591,N_1536,N_1511);
xor U1592 (N_1592,N_1531,N_1534);
and U1593 (N_1593,N_1551,N_1520);
nand U1594 (N_1594,N_1539,N_1535);
and U1595 (N_1595,N_1554,N_1548);
and U1596 (N_1596,N_1513,N_1520);
and U1597 (N_1597,N_1558,N_1537);
nand U1598 (N_1598,N_1535,N_1551);
nand U1599 (N_1599,N_1515,N_1549);
nor U1600 (N_1600,N_1506,N_1522);
xor U1601 (N_1601,N_1558,N_1500);
nor U1602 (N_1602,N_1533,N_1521);
or U1603 (N_1603,N_1515,N_1544);
nor U1604 (N_1604,N_1554,N_1522);
xnor U1605 (N_1605,N_1531,N_1554);
and U1606 (N_1606,N_1517,N_1514);
and U1607 (N_1607,N_1503,N_1516);
nand U1608 (N_1608,N_1545,N_1539);
and U1609 (N_1609,N_1520,N_1552);
nand U1610 (N_1610,N_1536,N_1551);
nand U1611 (N_1611,N_1526,N_1532);
and U1612 (N_1612,N_1507,N_1525);
and U1613 (N_1613,N_1543,N_1538);
xnor U1614 (N_1614,N_1548,N_1505);
or U1615 (N_1615,N_1523,N_1528);
nand U1616 (N_1616,N_1514,N_1547);
or U1617 (N_1617,N_1517,N_1503);
nand U1618 (N_1618,N_1538,N_1551);
nand U1619 (N_1619,N_1508,N_1528);
nand U1620 (N_1620,N_1598,N_1608);
xor U1621 (N_1621,N_1603,N_1594);
nand U1622 (N_1622,N_1592,N_1571);
nand U1623 (N_1623,N_1602,N_1584);
xnor U1624 (N_1624,N_1610,N_1585);
xor U1625 (N_1625,N_1586,N_1580);
or U1626 (N_1626,N_1611,N_1613);
and U1627 (N_1627,N_1617,N_1591);
nor U1628 (N_1628,N_1609,N_1576);
nor U1629 (N_1629,N_1616,N_1561);
xor U1630 (N_1630,N_1612,N_1593);
xnor U1631 (N_1631,N_1600,N_1601);
xnor U1632 (N_1632,N_1578,N_1574);
nor U1633 (N_1633,N_1618,N_1582);
or U1634 (N_1634,N_1572,N_1565);
nor U1635 (N_1635,N_1595,N_1564);
or U1636 (N_1636,N_1583,N_1563);
nand U1637 (N_1637,N_1570,N_1607);
or U1638 (N_1638,N_1614,N_1596);
and U1639 (N_1639,N_1562,N_1599);
xor U1640 (N_1640,N_1581,N_1568);
xor U1641 (N_1641,N_1577,N_1589);
nor U1642 (N_1642,N_1579,N_1569);
or U1643 (N_1643,N_1587,N_1590);
xnor U1644 (N_1644,N_1597,N_1619);
or U1645 (N_1645,N_1560,N_1606);
nor U1646 (N_1646,N_1604,N_1575);
nor U1647 (N_1647,N_1605,N_1615);
nand U1648 (N_1648,N_1588,N_1573);
and U1649 (N_1649,N_1566,N_1567);
and U1650 (N_1650,N_1574,N_1583);
nor U1651 (N_1651,N_1577,N_1593);
or U1652 (N_1652,N_1565,N_1571);
nand U1653 (N_1653,N_1605,N_1583);
or U1654 (N_1654,N_1577,N_1562);
nand U1655 (N_1655,N_1575,N_1605);
and U1656 (N_1656,N_1604,N_1586);
and U1657 (N_1657,N_1613,N_1562);
and U1658 (N_1658,N_1567,N_1578);
xor U1659 (N_1659,N_1571,N_1609);
and U1660 (N_1660,N_1582,N_1611);
xor U1661 (N_1661,N_1573,N_1587);
nor U1662 (N_1662,N_1561,N_1565);
or U1663 (N_1663,N_1616,N_1614);
and U1664 (N_1664,N_1591,N_1563);
and U1665 (N_1665,N_1574,N_1604);
or U1666 (N_1666,N_1575,N_1609);
nor U1667 (N_1667,N_1607,N_1609);
xor U1668 (N_1668,N_1601,N_1616);
xnor U1669 (N_1669,N_1585,N_1596);
and U1670 (N_1670,N_1602,N_1560);
nor U1671 (N_1671,N_1575,N_1603);
nor U1672 (N_1672,N_1580,N_1595);
nor U1673 (N_1673,N_1563,N_1569);
or U1674 (N_1674,N_1607,N_1619);
xor U1675 (N_1675,N_1580,N_1594);
xor U1676 (N_1676,N_1606,N_1597);
nand U1677 (N_1677,N_1564,N_1608);
or U1678 (N_1678,N_1567,N_1575);
nand U1679 (N_1679,N_1572,N_1602);
xor U1680 (N_1680,N_1649,N_1678);
xnor U1681 (N_1681,N_1646,N_1640);
and U1682 (N_1682,N_1662,N_1675);
and U1683 (N_1683,N_1664,N_1635);
and U1684 (N_1684,N_1658,N_1665);
nand U1685 (N_1685,N_1671,N_1630);
nor U1686 (N_1686,N_1634,N_1627);
or U1687 (N_1687,N_1623,N_1629);
and U1688 (N_1688,N_1676,N_1622);
nor U1689 (N_1689,N_1666,N_1621);
or U1690 (N_1690,N_1626,N_1642);
xor U1691 (N_1691,N_1641,N_1661);
and U1692 (N_1692,N_1648,N_1632);
and U1693 (N_1693,N_1636,N_1653);
nand U1694 (N_1694,N_1638,N_1633);
or U1695 (N_1695,N_1669,N_1625);
or U1696 (N_1696,N_1659,N_1652);
or U1697 (N_1697,N_1677,N_1667);
or U1698 (N_1698,N_1631,N_1663);
nor U1699 (N_1699,N_1645,N_1672);
and U1700 (N_1700,N_1670,N_1668);
and U1701 (N_1701,N_1624,N_1647);
xor U1702 (N_1702,N_1674,N_1650);
or U1703 (N_1703,N_1644,N_1660);
nand U1704 (N_1704,N_1637,N_1656);
and U1705 (N_1705,N_1655,N_1654);
xor U1706 (N_1706,N_1679,N_1651);
nand U1707 (N_1707,N_1620,N_1643);
nand U1708 (N_1708,N_1639,N_1628);
nand U1709 (N_1709,N_1657,N_1673);
nor U1710 (N_1710,N_1658,N_1661);
nor U1711 (N_1711,N_1620,N_1652);
nor U1712 (N_1712,N_1642,N_1645);
nor U1713 (N_1713,N_1628,N_1670);
xor U1714 (N_1714,N_1649,N_1629);
nand U1715 (N_1715,N_1621,N_1677);
nand U1716 (N_1716,N_1650,N_1679);
or U1717 (N_1717,N_1641,N_1642);
and U1718 (N_1718,N_1623,N_1643);
and U1719 (N_1719,N_1671,N_1667);
nor U1720 (N_1720,N_1663,N_1658);
or U1721 (N_1721,N_1653,N_1668);
nor U1722 (N_1722,N_1677,N_1637);
and U1723 (N_1723,N_1632,N_1629);
xor U1724 (N_1724,N_1674,N_1641);
and U1725 (N_1725,N_1643,N_1621);
nand U1726 (N_1726,N_1642,N_1663);
or U1727 (N_1727,N_1624,N_1676);
xor U1728 (N_1728,N_1676,N_1648);
and U1729 (N_1729,N_1630,N_1620);
nand U1730 (N_1730,N_1665,N_1675);
nor U1731 (N_1731,N_1628,N_1678);
and U1732 (N_1732,N_1655,N_1679);
or U1733 (N_1733,N_1650,N_1651);
and U1734 (N_1734,N_1660,N_1666);
nor U1735 (N_1735,N_1650,N_1672);
nor U1736 (N_1736,N_1665,N_1667);
and U1737 (N_1737,N_1645,N_1638);
xnor U1738 (N_1738,N_1655,N_1668);
and U1739 (N_1739,N_1626,N_1635);
xor U1740 (N_1740,N_1720,N_1733);
xor U1741 (N_1741,N_1710,N_1688);
and U1742 (N_1742,N_1709,N_1715);
nor U1743 (N_1743,N_1735,N_1736);
nand U1744 (N_1744,N_1724,N_1725);
nand U1745 (N_1745,N_1699,N_1701);
or U1746 (N_1746,N_1703,N_1738);
nor U1747 (N_1747,N_1719,N_1732);
or U1748 (N_1748,N_1718,N_1682);
nand U1749 (N_1749,N_1729,N_1692);
and U1750 (N_1750,N_1687,N_1722);
nand U1751 (N_1751,N_1684,N_1690);
and U1752 (N_1752,N_1728,N_1705);
and U1753 (N_1753,N_1712,N_1698);
nor U1754 (N_1754,N_1723,N_1714);
nor U1755 (N_1755,N_1739,N_1704);
nand U1756 (N_1756,N_1691,N_1716);
nor U1757 (N_1757,N_1702,N_1727);
xnor U1758 (N_1758,N_1708,N_1685);
xor U1759 (N_1759,N_1713,N_1731);
nand U1760 (N_1760,N_1695,N_1681);
and U1761 (N_1761,N_1726,N_1683);
nor U1762 (N_1762,N_1706,N_1730);
xor U1763 (N_1763,N_1711,N_1694);
or U1764 (N_1764,N_1721,N_1734);
xor U1765 (N_1765,N_1700,N_1707);
and U1766 (N_1766,N_1717,N_1696);
nand U1767 (N_1767,N_1737,N_1680);
or U1768 (N_1768,N_1689,N_1697);
or U1769 (N_1769,N_1686,N_1693);
and U1770 (N_1770,N_1713,N_1680);
and U1771 (N_1771,N_1728,N_1721);
nand U1772 (N_1772,N_1733,N_1696);
and U1773 (N_1773,N_1684,N_1729);
and U1774 (N_1774,N_1706,N_1716);
xor U1775 (N_1775,N_1733,N_1702);
and U1776 (N_1776,N_1723,N_1683);
or U1777 (N_1777,N_1725,N_1710);
nor U1778 (N_1778,N_1695,N_1705);
and U1779 (N_1779,N_1681,N_1727);
nor U1780 (N_1780,N_1732,N_1737);
and U1781 (N_1781,N_1718,N_1726);
and U1782 (N_1782,N_1716,N_1697);
xor U1783 (N_1783,N_1723,N_1726);
xor U1784 (N_1784,N_1735,N_1695);
and U1785 (N_1785,N_1681,N_1717);
xnor U1786 (N_1786,N_1706,N_1721);
xnor U1787 (N_1787,N_1697,N_1700);
nand U1788 (N_1788,N_1705,N_1696);
or U1789 (N_1789,N_1695,N_1686);
and U1790 (N_1790,N_1736,N_1688);
or U1791 (N_1791,N_1689,N_1691);
nand U1792 (N_1792,N_1705,N_1684);
xnor U1793 (N_1793,N_1690,N_1701);
nor U1794 (N_1794,N_1718,N_1699);
nor U1795 (N_1795,N_1722,N_1704);
xnor U1796 (N_1796,N_1718,N_1739);
nor U1797 (N_1797,N_1731,N_1701);
nor U1798 (N_1798,N_1701,N_1719);
and U1799 (N_1799,N_1736,N_1710);
nor U1800 (N_1800,N_1756,N_1798);
or U1801 (N_1801,N_1763,N_1743);
or U1802 (N_1802,N_1796,N_1794);
nor U1803 (N_1803,N_1783,N_1761);
and U1804 (N_1804,N_1775,N_1740);
nand U1805 (N_1805,N_1766,N_1781);
nand U1806 (N_1806,N_1773,N_1771);
or U1807 (N_1807,N_1790,N_1770);
xnor U1808 (N_1808,N_1777,N_1753);
and U1809 (N_1809,N_1779,N_1742);
nand U1810 (N_1810,N_1769,N_1755);
nor U1811 (N_1811,N_1789,N_1749);
or U1812 (N_1812,N_1741,N_1746);
nor U1813 (N_1813,N_1754,N_1776);
nor U1814 (N_1814,N_1764,N_1758);
or U1815 (N_1815,N_1786,N_1791);
nor U1816 (N_1816,N_1747,N_1778);
and U1817 (N_1817,N_1784,N_1767);
or U1818 (N_1818,N_1780,N_1745);
nand U1819 (N_1819,N_1760,N_1762);
and U1820 (N_1820,N_1795,N_1785);
or U1821 (N_1821,N_1757,N_1799);
or U1822 (N_1822,N_1772,N_1768);
xor U1823 (N_1823,N_1793,N_1748);
nand U1824 (N_1824,N_1765,N_1752);
nor U1825 (N_1825,N_1792,N_1759);
nand U1826 (N_1826,N_1744,N_1782);
or U1827 (N_1827,N_1774,N_1797);
xor U1828 (N_1828,N_1788,N_1750);
or U1829 (N_1829,N_1787,N_1751);
or U1830 (N_1830,N_1764,N_1799);
or U1831 (N_1831,N_1776,N_1779);
nand U1832 (N_1832,N_1797,N_1753);
nand U1833 (N_1833,N_1785,N_1781);
nor U1834 (N_1834,N_1783,N_1794);
and U1835 (N_1835,N_1783,N_1753);
and U1836 (N_1836,N_1768,N_1780);
xnor U1837 (N_1837,N_1773,N_1745);
and U1838 (N_1838,N_1757,N_1796);
nand U1839 (N_1839,N_1787,N_1786);
nand U1840 (N_1840,N_1769,N_1758);
or U1841 (N_1841,N_1793,N_1784);
xnor U1842 (N_1842,N_1785,N_1787);
and U1843 (N_1843,N_1763,N_1798);
xnor U1844 (N_1844,N_1782,N_1790);
nor U1845 (N_1845,N_1798,N_1751);
or U1846 (N_1846,N_1744,N_1745);
xnor U1847 (N_1847,N_1764,N_1777);
or U1848 (N_1848,N_1765,N_1796);
xor U1849 (N_1849,N_1794,N_1760);
or U1850 (N_1850,N_1740,N_1759);
or U1851 (N_1851,N_1776,N_1767);
or U1852 (N_1852,N_1766,N_1741);
nand U1853 (N_1853,N_1774,N_1760);
xor U1854 (N_1854,N_1790,N_1791);
and U1855 (N_1855,N_1768,N_1793);
nor U1856 (N_1856,N_1782,N_1768);
or U1857 (N_1857,N_1745,N_1770);
or U1858 (N_1858,N_1745,N_1766);
xnor U1859 (N_1859,N_1764,N_1776);
or U1860 (N_1860,N_1812,N_1831);
nand U1861 (N_1861,N_1838,N_1826);
nand U1862 (N_1862,N_1825,N_1842);
or U1863 (N_1863,N_1832,N_1859);
and U1864 (N_1864,N_1833,N_1823);
nand U1865 (N_1865,N_1804,N_1817);
nand U1866 (N_1866,N_1837,N_1805);
xor U1867 (N_1867,N_1858,N_1815);
and U1868 (N_1868,N_1813,N_1836);
or U1869 (N_1869,N_1811,N_1843);
nand U1870 (N_1870,N_1807,N_1819);
and U1871 (N_1871,N_1809,N_1818);
xor U1872 (N_1872,N_1839,N_1834);
and U1873 (N_1873,N_1855,N_1853);
and U1874 (N_1874,N_1822,N_1846);
xor U1875 (N_1875,N_1829,N_1830);
and U1876 (N_1876,N_1810,N_1814);
nand U1877 (N_1877,N_1821,N_1835);
xnor U1878 (N_1878,N_1856,N_1828);
xnor U1879 (N_1879,N_1816,N_1802);
or U1880 (N_1880,N_1851,N_1806);
and U1881 (N_1881,N_1845,N_1841);
nor U1882 (N_1882,N_1849,N_1857);
nor U1883 (N_1883,N_1820,N_1840);
or U1884 (N_1884,N_1801,N_1852);
nand U1885 (N_1885,N_1800,N_1850);
xor U1886 (N_1886,N_1808,N_1847);
nor U1887 (N_1887,N_1803,N_1827);
and U1888 (N_1888,N_1848,N_1824);
nand U1889 (N_1889,N_1844,N_1854);
nand U1890 (N_1890,N_1836,N_1855);
xnor U1891 (N_1891,N_1852,N_1807);
xor U1892 (N_1892,N_1850,N_1805);
or U1893 (N_1893,N_1838,N_1832);
and U1894 (N_1894,N_1814,N_1818);
nand U1895 (N_1895,N_1832,N_1847);
nand U1896 (N_1896,N_1822,N_1830);
or U1897 (N_1897,N_1850,N_1811);
nor U1898 (N_1898,N_1852,N_1857);
xor U1899 (N_1899,N_1843,N_1800);
or U1900 (N_1900,N_1844,N_1848);
nor U1901 (N_1901,N_1818,N_1853);
xor U1902 (N_1902,N_1848,N_1833);
nand U1903 (N_1903,N_1817,N_1859);
nor U1904 (N_1904,N_1851,N_1837);
nor U1905 (N_1905,N_1835,N_1805);
nand U1906 (N_1906,N_1806,N_1822);
and U1907 (N_1907,N_1844,N_1805);
or U1908 (N_1908,N_1827,N_1833);
nand U1909 (N_1909,N_1802,N_1839);
nand U1910 (N_1910,N_1806,N_1827);
or U1911 (N_1911,N_1851,N_1801);
and U1912 (N_1912,N_1809,N_1819);
and U1913 (N_1913,N_1811,N_1803);
nand U1914 (N_1914,N_1851,N_1835);
nor U1915 (N_1915,N_1816,N_1804);
nor U1916 (N_1916,N_1859,N_1803);
xor U1917 (N_1917,N_1839,N_1846);
nand U1918 (N_1918,N_1815,N_1809);
nor U1919 (N_1919,N_1805,N_1851);
nand U1920 (N_1920,N_1899,N_1866);
and U1921 (N_1921,N_1883,N_1870);
nor U1922 (N_1922,N_1908,N_1919);
xor U1923 (N_1923,N_1873,N_1867);
or U1924 (N_1924,N_1918,N_1868);
nor U1925 (N_1925,N_1891,N_1879);
xnor U1926 (N_1926,N_1865,N_1915);
nand U1927 (N_1927,N_1905,N_1881);
nor U1928 (N_1928,N_1896,N_1888);
nand U1929 (N_1929,N_1894,N_1869);
and U1930 (N_1930,N_1861,N_1911);
or U1931 (N_1931,N_1890,N_1886);
nor U1932 (N_1932,N_1917,N_1889);
nand U1933 (N_1933,N_1916,N_1862);
and U1934 (N_1934,N_1904,N_1912);
xnor U1935 (N_1935,N_1903,N_1878);
nor U1936 (N_1936,N_1885,N_1892);
xor U1937 (N_1937,N_1864,N_1874);
or U1938 (N_1938,N_1876,N_1887);
nor U1939 (N_1939,N_1863,N_1910);
and U1940 (N_1940,N_1897,N_1875);
or U1941 (N_1941,N_1882,N_1909);
nand U1942 (N_1942,N_1880,N_1884);
xor U1943 (N_1943,N_1895,N_1902);
nand U1944 (N_1944,N_1898,N_1907);
nand U1945 (N_1945,N_1901,N_1872);
nor U1946 (N_1946,N_1871,N_1860);
or U1947 (N_1947,N_1914,N_1913);
nor U1948 (N_1948,N_1877,N_1900);
or U1949 (N_1949,N_1893,N_1906);
nand U1950 (N_1950,N_1894,N_1914);
xor U1951 (N_1951,N_1907,N_1912);
or U1952 (N_1952,N_1888,N_1861);
xor U1953 (N_1953,N_1890,N_1873);
and U1954 (N_1954,N_1915,N_1894);
xnor U1955 (N_1955,N_1879,N_1860);
nand U1956 (N_1956,N_1917,N_1913);
nand U1957 (N_1957,N_1896,N_1892);
and U1958 (N_1958,N_1878,N_1874);
nand U1959 (N_1959,N_1904,N_1884);
or U1960 (N_1960,N_1892,N_1862);
nor U1961 (N_1961,N_1877,N_1890);
nand U1962 (N_1962,N_1895,N_1887);
or U1963 (N_1963,N_1888,N_1907);
or U1964 (N_1964,N_1903,N_1919);
and U1965 (N_1965,N_1889,N_1887);
nand U1966 (N_1966,N_1883,N_1898);
nor U1967 (N_1967,N_1867,N_1910);
nand U1968 (N_1968,N_1868,N_1872);
and U1969 (N_1969,N_1912,N_1860);
nor U1970 (N_1970,N_1919,N_1914);
nand U1971 (N_1971,N_1911,N_1885);
or U1972 (N_1972,N_1884,N_1910);
xor U1973 (N_1973,N_1911,N_1894);
and U1974 (N_1974,N_1876,N_1913);
xnor U1975 (N_1975,N_1891,N_1919);
or U1976 (N_1976,N_1917,N_1899);
xor U1977 (N_1977,N_1902,N_1882);
nor U1978 (N_1978,N_1903,N_1901);
or U1979 (N_1979,N_1898,N_1886);
or U1980 (N_1980,N_1929,N_1930);
or U1981 (N_1981,N_1968,N_1928);
xor U1982 (N_1982,N_1953,N_1954);
xnor U1983 (N_1983,N_1950,N_1971);
and U1984 (N_1984,N_1975,N_1972);
and U1985 (N_1985,N_1966,N_1962);
and U1986 (N_1986,N_1926,N_1932);
nor U1987 (N_1987,N_1936,N_1959);
nor U1988 (N_1988,N_1969,N_1927);
nor U1989 (N_1989,N_1958,N_1947);
nand U1990 (N_1990,N_1921,N_1925);
and U1991 (N_1991,N_1940,N_1976);
and U1992 (N_1992,N_1964,N_1978);
nor U1993 (N_1993,N_1931,N_1956);
or U1994 (N_1994,N_1979,N_1938);
or U1995 (N_1995,N_1949,N_1963);
nand U1996 (N_1996,N_1957,N_1961);
or U1997 (N_1997,N_1955,N_1946);
or U1998 (N_1998,N_1948,N_1977);
or U1999 (N_1999,N_1967,N_1943);
xnor U2000 (N_2000,N_1944,N_1920);
nand U2001 (N_2001,N_1952,N_1933);
and U2002 (N_2002,N_1945,N_1960);
nor U2003 (N_2003,N_1942,N_1935);
nand U2004 (N_2004,N_1974,N_1941);
and U2005 (N_2005,N_1922,N_1951);
or U2006 (N_2006,N_1923,N_1924);
nand U2007 (N_2007,N_1973,N_1970);
and U2008 (N_2008,N_1934,N_1965);
nand U2009 (N_2009,N_1939,N_1937);
xor U2010 (N_2010,N_1966,N_1951);
or U2011 (N_2011,N_1958,N_1920);
or U2012 (N_2012,N_1927,N_1963);
nor U2013 (N_2013,N_1962,N_1931);
nand U2014 (N_2014,N_1940,N_1950);
xor U2015 (N_2015,N_1972,N_1924);
xnor U2016 (N_2016,N_1956,N_1951);
nand U2017 (N_2017,N_1933,N_1947);
nor U2018 (N_2018,N_1941,N_1924);
nand U2019 (N_2019,N_1955,N_1953);
nand U2020 (N_2020,N_1971,N_1922);
nor U2021 (N_2021,N_1962,N_1945);
nor U2022 (N_2022,N_1952,N_1924);
nor U2023 (N_2023,N_1964,N_1948);
xnor U2024 (N_2024,N_1960,N_1961);
nor U2025 (N_2025,N_1978,N_1938);
and U2026 (N_2026,N_1928,N_1926);
xor U2027 (N_2027,N_1958,N_1972);
xnor U2028 (N_2028,N_1923,N_1971);
nor U2029 (N_2029,N_1927,N_1931);
and U2030 (N_2030,N_1967,N_1964);
nor U2031 (N_2031,N_1963,N_1951);
and U2032 (N_2032,N_1944,N_1958);
and U2033 (N_2033,N_1948,N_1958);
or U2034 (N_2034,N_1929,N_1944);
xor U2035 (N_2035,N_1956,N_1943);
nand U2036 (N_2036,N_1923,N_1934);
nand U2037 (N_2037,N_1975,N_1974);
nand U2038 (N_2038,N_1922,N_1973);
nor U2039 (N_2039,N_1948,N_1965);
xor U2040 (N_2040,N_1984,N_1997);
nor U2041 (N_2041,N_1999,N_2024);
nand U2042 (N_2042,N_1980,N_1992);
or U2043 (N_2043,N_2008,N_1998);
xnor U2044 (N_2044,N_2022,N_1986);
or U2045 (N_2045,N_2016,N_1985);
nand U2046 (N_2046,N_2027,N_2030);
and U2047 (N_2047,N_1993,N_2009);
nand U2048 (N_2048,N_2029,N_2037);
xor U2049 (N_2049,N_2028,N_2015);
nor U2050 (N_2050,N_2036,N_2026);
nand U2051 (N_2051,N_1987,N_2034);
nor U2052 (N_2052,N_1996,N_1995);
and U2053 (N_2053,N_2023,N_2011);
and U2054 (N_2054,N_2038,N_2014);
nor U2055 (N_2055,N_2000,N_2032);
xor U2056 (N_2056,N_2003,N_2020);
xor U2057 (N_2057,N_1982,N_1991);
nand U2058 (N_2058,N_1994,N_1990);
or U2059 (N_2059,N_2012,N_2013);
xor U2060 (N_2060,N_2021,N_2002);
nand U2061 (N_2061,N_2007,N_2006);
xor U2062 (N_2062,N_2001,N_2004);
or U2063 (N_2063,N_1988,N_2031);
or U2064 (N_2064,N_2017,N_2035);
nand U2065 (N_2065,N_1983,N_2019);
xor U2066 (N_2066,N_2039,N_1981);
xnor U2067 (N_2067,N_1989,N_2025);
or U2068 (N_2068,N_2010,N_2033);
nand U2069 (N_2069,N_2005,N_2018);
nor U2070 (N_2070,N_1985,N_2034);
and U2071 (N_2071,N_2008,N_1987);
xor U2072 (N_2072,N_2028,N_1991);
nand U2073 (N_2073,N_2039,N_2002);
or U2074 (N_2074,N_1996,N_1997);
xnor U2075 (N_2075,N_2011,N_1981);
or U2076 (N_2076,N_1992,N_1999);
or U2077 (N_2077,N_2039,N_2015);
nand U2078 (N_2078,N_1997,N_2037);
and U2079 (N_2079,N_2011,N_1991);
nand U2080 (N_2080,N_2011,N_2026);
nor U2081 (N_2081,N_2009,N_2006);
or U2082 (N_2082,N_2026,N_2008);
and U2083 (N_2083,N_2011,N_2020);
nor U2084 (N_2084,N_1991,N_2036);
or U2085 (N_2085,N_2034,N_1981);
nor U2086 (N_2086,N_2007,N_2016);
or U2087 (N_2087,N_1989,N_2031);
and U2088 (N_2088,N_2016,N_1996);
or U2089 (N_2089,N_2002,N_2007);
nor U2090 (N_2090,N_2001,N_2019);
and U2091 (N_2091,N_1981,N_2005);
and U2092 (N_2092,N_2008,N_1982);
and U2093 (N_2093,N_2012,N_2016);
xnor U2094 (N_2094,N_1986,N_2013);
or U2095 (N_2095,N_1985,N_2011);
xnor U2096 (N_2096,N_2032,N_1987);
or U2097 (N_2097,N_2035,N_1992);
nand U2098 (N_2098,N_2000,N_1998);
nand U2099 (N_2099,N_2037,N_2022);
and U2100 (N_2100,N_2050,N_2074);
or U2101 (N_2101,N_2097,N_2088);
nand U2102 (N_2102,N_2084,N_2049);
nand U2103 (N_2103,N_2078,N_2040);
and U2104 (N_2104,N_2092,N_2071);
xor U2105 (N_2105,N_2099,N_2043);
nand U2106 (N_2106,N_2058,N_2093);
or U2107 (N_2107,N_2048,N_2052);
and U2108 (N_2108,N_2094,N_2087);
and U2109 (N_2109,N_2055,N_2063);
and U2110 (N_2110,N_2095,N_2065);
and U2111 (N_2111,N_2072,N_2046);
xor U2112 (N_2112,N_2076,N_2067);
nand U2113 (N_2113,N_2069,N_2091);
nand U2114 (N_2114,N_2096,N_2047);
nand U2115 (N_2115,N_2068,N_2090);
xor U2116 (N_2116,N_2051,N_2070);
or U2117 (N_2117,N_2082,N_2061);
or U2118 (N_2118,N_2042,N_2075);
or U2119 (N_2119,N_2057,N_2059);
or U2120 (N_2120,N_2044,N_2080);
and U2121 (N_2121,N_2054,N_2089);
nand U2122 (N_2122,N_2073,N_2079);
nand U2123 (N_2123,N_2045,N_2085);
or U2124 (N_2124,N_2053,N_2041);
nand U2125 (N_2125,N_2064,N_2098);
or U2126 (N_2126,N_2077,N_2081);
xor U2127 (N_2127,N_2083,N_2086);
nand U2128 (N_2128,N_2062,N_2066);
or U2129 (N_2129,N_2060,N_2056);
and U2130 (N_2130,N_2050,N_2060);
nand U2131 (N_2131,N_2042,N_2086);
nand U2132 (N_2132,N_2073,N_2093);
or U2133 (N_2133,N_2084,N_2061);
nor U2134 (N_2134,N_2094,N_2079);
and U2135 (N_2135,N_2097,N_2095);
nor U2136 (N_2136,N_2068,N_2093);
or U2137 (N_2137,N_2063,N_2083);
xnor U2138 (N_2138,N_2046,N_2084);
and U2139 (N_2139,N_2061,N_2053);
xor U2140 (N_2140,N_2099,N_2066);
xnor U2141 (N_2141,N_2063,N_2041);
nor U2142 (N_2142,N_2080,N_2096);
nor U2143 (N_2143,N_2089,N_2057);
and U2144 (N_2144,N_2095,N_2080);
or U2145 (N_2145,N_2087,N_2049);
and U2146 (N_2146,N_2088,N_2049);
nand U2147 (N_2147,N_2088,N_2070);
xnor U2148 (N_2148,N_2060,N_2041);
and U2149 (N_2149,N_2072,N_2060);
xor U2150 (N_2150,N_2062,N_2058);
or U2151 (N_2151,N_2095,N_2092);
or U2152 (N_2152,N_2059,N_2061);
or U2153 (N_2153,N_2079,N_2088);
or U2154 (N_2154,N_2099,N_2069);
and U2155 (N_2155,N_2049,N_2094);
xnor U2156 (N_2156,N_2082,N_2046);
and U2157 (N_2157,N_2053,N_2062);
xnor U2158 (N_2158,N_2071,N_2050);
nand U2159 (N_2159,N_2059,N_2068);
and U2160 (N_2160,N_2142,N_2152);
nor U2161 (N_2161,N_2151,N_2131);
nor U2162 (N_2162,N_2155,N_2130);
and U2163 (N_2163,N_2128,N_2149);
nor U2164 (N_2164,N_2119,N_2102);
and U2165 (N_2165,N_2129,N_2106);
and U2166 (N_2166,N_2110,N_2157);
nor U2167 (N_2167,N_2100,N_2120);
and U2168 (N_2168,N_2144,N_2134);
nor U2169 (N_2169,N_2146,N_2103);
nor U2170 (N_2170,N_2121,N_2114);
nand U2171 (N_2171,N_2116,N_2112);
nand U2172 (N_2172,N_2104,N_2115);
and U2173 (N_2173,N_2127,N_2118);
xnor U2174 (N_2174,N_2147,N_2137);
or U2175 (N_2175,N_2133,N_2126);
nor U2176 (N_2176,N_2125,N_2124);
and U2177 (N_2177,N_2111,N_2141);
or U2178 (N_2178,N_2101,N_2143);
or U2179 (N_2179,N_2153,N_2113);
and U2180 (N_2180,N_2136,N_2154);
nor U2181 (N_2181,N_2123,N_2135);
nand U2182 (N_2182,N_2122,N_2148);
nor U2183 (N_2183,N_2117,N_2158);
nor U2184 (N_2184,N_2159,N_2156);
and U2185 (N_2185,N_2145,N_2105);
or U2186 (N_2186,N_2139,N_2132);
or U2187 (N_2187,N_2140,N_2109);
and U2188 (N_2188,N_2138,N_2108);
nor U2189 (N_2189,N_2107,N_2150);
and U2190 (N_2190,N_2119,N_2158);
or U2191 (N_2191,N_2138,N_2143);
nand U2192 (N_2192,N_2151,N_2101);
and U2193 (N_2193,N_2116,N_2110);
xnor U2194 (N_2194,N_2137,N_2159);
nand U2195 (N_2195,N_2123,N_2118);
nor U2196 (N_2196,N_2138,N_2103);
and U2197 (N_2197,N_2138,N_2133);
and U2198 (N_2198,N_2120,N_2124);
and U2199 (N_2199,N_2151,N_2136);
or U2200 (N_2200,N_2109,N_2103);
nand U2201 (N_2201,N_2128,N_2154);
nand U2202 (N_2202,N_2118,N_2114);
xor U2203 (N_2203,N_2133,N_2119);
and U2204 (N_2204,N_2138,N_2146);
or U2205 (N_2205,N_2131,N_2136);
and U2206 (N_2206,N_2134,N_2150);
and U2207 (N_2207,N_2149,N_2139);
nor U2208 (N_2208,N_2155,N_2119);
or U2209 (N_2209,N_2140,N_2125);
and U2210 (N_2210,N_2139,N_2101);
nand U2211 (N_2211,N_2107,N_2125);
nand U2212 (N_2212,N_2128,N_2106);
nor U2213 (N_2213,N_2100,N_2156);
or U2214 (N_2214,N_2147,N_2122);
nand U2215 (N_2215,N_2157,N_2125);
or U2216 (N_2216,N_2140,N_2100);
nor U2217 (N_2217,N_2158,N_2105);
and U2218 (N_2218,N_2112,N_2123);
nor U2219 (N_2219,N_2122,N_2110);
or U2220 (N_2220,N_2181,N_2207);
xnor U2221 (N_2221,N_2165,N_2174);
xor U2222 (N_2222,N_2188,N_2211);
nand U2223 (N_2223,N_2217,N_2162);
or U2224 (N_2224,N_2176,N_2189);
or U2225 (N_2225,N_2187,N_2219);
nand U2226 (N_2226,N_2205,N_2175);
nor U2227 (N_2227,N_2194,N_2214);
or U2228 (N_2228,N_2163,N_2201);
and U2229 (N_2229,N_2198,N_2178);
xor U2230 (N_2230,N_2192,N_2161);
nor U2231 (N_2231,N_2185,N_2203);
nor U2232 (N_2232,N_2166,N_2186);
or U2233 (N_2233,N_2177,N_2170);
xor U2234 (N_2234,N_2218,N_2200);
and U2235 (N_2235,N_2179,N_2184);
nor U2236 (N_2236,N_2204,N_2171);
xnor U2237 (N_2237,N_2167,N_2206);
xor U2238 (N_2238,N_2169,N_2199);
and U2239 (N_2239,N_2164,N_2182);
nor U2240 (N_2240,N_2173,N_2208);
nand U2241 (N_2241,N_2195,N_2160);
nor U2242 (N_2242,N_2212,N_2190);
nand U2243 (N_2243,N_2193,N_2172);
nand U2244 (N_2244,N_2196,N_2209);
or U2245 (N_2245,N_2180,N_2183);
or U2246 (N_2246,N_2191,N_2202);
xor U2247 (N_2247,N_2168,N_2213);
nand U2248 (N_2248,N_2215,N_2216);
nor U2249 (N_2249,N_2197,N_2210);
xnor U2250 (N_2250,N_2172,N_2216);
and U2251 (N_2251,N_2202,N_2194);
or U2252 (N_2252,N_2204,N_2201);
xnor U2253 (N_2253,N_2188,N_2208);
xor U2254 (N_2254,N_2179,N_2208);
and U2255 (N_2255,N_2202,N_2195);
xor U2256 (N_2256,N_2203,N_2194);
nand U2257 (N_2257,N_2178,N_2202);
nor U2258 (N_2258,N_2179,N_2173);
nor U2259 (N_2259,N_2176,N_2173);
nor U2260 (N_2260,N_2197,N_2209);
or U2261 (N_2261,N_2176,N_2208);
or U2262 (N_2262,N_2175,N_2203);
nand U2263 (N_2263,N_2186,N_2177);
or U2264 (N_2264,N_2179,N_2216);
and U2265 (N_2265,N_2201,N_2211);
xnor U2266 (N_2266,N_2168,N_2177);
nor U2267 (N_2267,N_2184,N_2208);
or U2268 (N_2268,N_2189,N_2208);
nand U2269 (N_2269,N_2217,N_2203);
nor U2270 (N_2270,N_2160,N_2216);
or U2271 (N_2271,N_2183,N_2184);
xor U2272 (N_2272,N_2203,N_2197);
nand U2273 (N_2273,N_2213,N_2183);
nand U2274 (N_2274,N_2211,N_2215);
nor U2275 (N_2275,N_2163,N_2194);
and U2276 (N_2276,N_2189,N_2169);
or U2277 (N_2277,N_2204,N_2214);
xnor U2278 (N_2278,N_2202,N_2170);
nand U2279 (N_2279,N_2203,N_2174);
nand U2280 (N_2280,N_2251,N_2271);
nand U2281 (N_2281,N_2256,N_2261);
and U2282 (N_2282,N_2264,N_2241);
and U2283 (N_2283,N_2228,N_2274);
nor U2284 (N_2284,N_2222,N_2268);
nand U2285 (N_2285,N_2279,N_2239);
nand U2286 (N_2286,N_2224,N_2266);
xnor U2287 (N_2287,N_2221,N_2240);
nor U2288 (N_2288,N_2269,N_2238);
xnor U2289 (N_2289,N_2257,N_2233);
nand U2290 (N_2290,N_2225,N_2248);
nand U2291 (N_2291,N_2237,N_2254);
xnor U2292 (N_2292,N_2245,N_2236);
nor U2293 (N_2293,N_2232,N_2273);
or U2294 (N_2294,N_2276,N_2270);
nand U2295 (N_2295,N_2267,N_2259);
and U2296 (N_2296,N_2253,N_2246);
and U2297 (N_2297,N_2226,N_2247);
and U2298 (N_2298,N_2249,N_2223);
nor U2299 (N_2299,N_2220,N_2258);
or U2300 (N_2300,N_2231,N_2229);
nand U2301 (N_2301,N_2242,N_2265);
xnor U2302 (N_2302,N_2227,N_2243);
or U2303 (N_2303,N_2255,N_2272);
and U2304 (N_2304,N_2275,N_2277);
and U2305 (N_2305,N_2250,N_2262);
nor U2306 (N_2306,N_2260,N_2234);
nand U2307 (N_2307,N_2278,N_2252);
or U2308 (N_2308,N_2235,N_2230);
nor U2309 (N_2309,N_2244,N_2263);
or U2310 (N_2310,N_2258,N_2224);
or U2311 (N_2311,N_2242,N_2263);
nor U2312 (N_2312,N_2270,N_2220);
and U2313 (N_2313,N_2234,N_2220);
xnor U2314 (N_2314,N_2266,N_2257);
or U2315 (N_2315,N_2238,N_2222);
xnor U2316 (N_2316,N_2238,N_2266);
nand U2317 (N_2317,N_2252,N_2275);
or U2318 (N_2318,N_2252,N_2262);
or U2319 (N_2319,N_2267,N_2261);
or U2320 (N_2320,N_2260,N_2258);
nand U2321 (N_2321,N_2225,N_2234);
or U2322 (N_2322,N_2223,N_2221);
and U2323 (N_2323,N_2262,N_2231);
xnor U2324 (N_2324,N_2262,N_2263);
or U2325 (N_2325,N_2245,N_2256);
and U2326 (N_2326,N_2235,N_2275);
or U2327 (N_2327,N_2265,N_2232);
nand U2328 (N_2328,N_2258,N_2226);
xor U2329 (N_2329,N_2235,N_2241);
nor U2330 (N_2330,N_2223,N_2239);
nand U2331 (N_2331,N_2253,N_2261);
nor U2332 (N_2332,N_2228,N_2223);
nand U2333 (N_2333,N_2249,N_2272);
or U2334 (N_2334,N_2235,N_2270);
or U2335 (N_2335,N_2262,N_2249);
and U2336 (N_2336,N_2255,N_2244);
or U2337 (N_2337,N_2278,N_2254);
xnor U2338 (N_2338,N_2220,N_2241);
nor U2339 (N_2339,N_2250,N_2222);
or U2340 (N_2340,N_2293,N_2339);
or U2341 (N_2341,N_2296,N_2303);
or U2342 (N_2342,N_2292,N_2291);
nand U2343 (N_2343,N_2298,N_2304);
nor U2344 (N_2344,N_2335,N_2281);
xnor U2345 (N_2345,N_2300,N_2329);
nor U2346 (N_2346,N_2280,N_2320);
or U2347 (N_2347,N_2317,N_2308);
xor U2348 (N_2348,N_2316,N_2336);
nand U2349 (N_2349,N_2330,N_2326);
nor U2350 (N_2350,N_2299,N_2319);
and U2351 (N_2351,N_2338,N_2318);
xnor U2352 (N_2352,N_2302,N_2295);
nor U2353 (N_2353,N_2334,N_2287);
nand U2354 (N_2354,N_2301,N_2297);
xor U2355 (N_2355,N_2337,N_2288);
nand U2356 (N_2356,N_2311,N_2289);
xnor U2357 (N_2357,N_2309,N_2328);
xnor U2358 (N_2358,N_2314,N_2331);
nand U2359 (N_2359,N_2305,N_2307);
nand U2360 (N_2360,N_2332,N_2333);
nor U2361 (N_2361,N_2294,N_2324);
nor U2362 (N_2362,N_2282,N_2322);
and U2363 (N_2363,N_2323,N_2283);
nand U2364 (N_2364,N_2306,N_2285);
nand U2365 (N_2365,N_2315,N_2313);
nand U2366 (N_2366,N_2327,N_2290);
nand U2367 (N_2367,N_2284,N_2286);
and U2368 (N_2368,N_2321,N_2325);
nand U2369 (N_2369,N_2310,N_2312);
and U2370 (N_2370,N_2290,N_2313);
nand U2371 (N_2371,N_2304,N_2308);
or U2372 (N_2372,N_2318,N_2302);
nor U2373 (N_2373,N_2308,N_2331);
nand U2374 (N_2374,N_2295,N_2303);
nor U2375 (N_2375,N_2281,N_2289);
nor U2376 (N_2376,N_2289,N_2304);
xor U2377 (N_2377,N_2297,N_2330);
nor U2378 (N_2378,N_2328,N_2320);
xor U2379 (N_2379,N_2294,N_2305);
nor U2380 (N_2380,N_2317,N_2338);
nor U2381 (N_2381,N_2288,N_2309);
nand U2382 (N_2382,N_2338,N_2298);
nor U2383 (N_2383,N_2290,N_2312);
or U2384 (N_2384,N_2318,N_2309);
nor U2385 (N_2385,N_2335,N_2319);
nand U2386 (N_2386,N_2333,N_2295);
nand U2387 (N_2387,N_2283,N_2312);
xnor U2388 (N_2388,N_2336,N_2296);
or U2389 (N_2389,N_2293,N_2302);
or U2390 (N_2390,N_2286,N_2289);
xor U2391 (N_2391,N_2286,N_2318);
or U2392 (N_2392,N_2282,N_2333);
nand U2393 (N_2393,N_2300,N_2318);
nand U2394 (N_2394,N_2328,N_2300);
xnor U2395 (N_2395,N_2306,N_2310);
xor U2396 (N_2396,N_2294,N_2315);
or U2397 (N_2397,N_2291,N_2303);
nand U2398 (N_2398,N_2332,N_2330);
and U2399 (N_2399,N_2296,N_2293);
or U2400 (N_2400,N_2371,N_2356);
nor U2401 (N_2401,N_2392,N_2372);
xnor U2402 (N_2402,N_2376,N_2397);
and U2403 (N_2403,N_2389,N_2370);
xnor U2404 (N_2404,N_2355,N_2394);
or U2405 (N_2405,N_2358,N_2386);
and U2406 (N_2406,N_2360,N_2362);
or U2407 (N_2407,N_2348,N_2365);
xnor U2408 (N_2408,N_2393,N_2343);
xor U2409 (N_2409,N_2347,N_2388);
and U2410 (N_2410,N_2344,N_2382);
xnor U2411 (N_2411,N_2399,N_2380);
xnor U2412 (N_2412,N_2366,N_2341);
nor U2413 (N_2413,N_2345,N_2398);
or U2414 (N_2414,N_2342,N_2391);
and U2415 (N_2415,N_2379,N_2346);
xnor U2416 (N_2416,N_2384,N_2353);
nand U2417 (N_2417,N_2340,N_2390);
and U2418 (N_2418,N_2350,N_2373);
or U2419 (N_2419,N_2361,N_2368);
or U2420 (N_2420,N_2367,N_2375);
nor U2421 (N_2421,N_2387,N_2381);
and U2422 (N_2422,N_2396,N_2357);
xor U2423 (N_2423,N_2364,N_2385);
xnor U2424 (N_2424,N_2374,N_2383);
xor U2425 (N_2425,N_2395,N_2352);
and U2426 (N_2426,N_2363,N_2369);
or U2427 (N_2427,N_2349,N_2351);
nor U2428 (N_2428,N_2378,N_2377);
or U2429 (N_2429,N_2359,N_2354);
nor U2430 (N_2430,N_2370,N_2369);
and U2431 (N_2431,N_2371,N_2340);
nor U2432 (N_2432,N_2357,N_2397);
or U2433 (N_2433,N_2387,N_2360);
xor U2434 (N_2434,N_2372,N_2357);
and U2435 (N_2435,N_2382,N_2353);
nand U2436 (N_2436,N_2355,N_2364);
or U2437 (N_2437,N_2391,N_2395);
nand U2438 (N_2438,N_2391,N_2371);
nand U2439 (N_2439,N_2354,N_2387);
nor U2440 (N_2440,N_2353,N_2365);
or U2441 (N_2441,N_2396,N_2342);
or U2442 (N_2442,N_2372,N_2345);
and U2443 (N_2443,N_2352,N_2349);
xor U2444 (N_2444,N_2391,N_2392);
nand U2445 (N_2445,N_2372,N_2361);
and U2446 (N_2446,N_2350,N_2399);
nand U2447 (N_2447,N_2351,N_2373);
xor U2448 (N_2448,N_2354,N_2383);
and U2449 (N_2449,N_2399,N_2386);
nand U2450 (N_2450,N_2352,N_2350);
xnor U2451 (N_2451,N_2359,N_2363);
xor U2452 (N_2452,N_2384,N_2341);
or U2453 (N_2453,N_2350,N_2395);
or U2454 (N_2454,N_2397,N_2362);
and U2455 (N_2455,N_2374,N_2386);
and U2456 (N_2456,N_2348,N_2361);
xnor U2457 (N_2457,N_2377,N_2347);
xor U2458 (N_2458,N_2364,N_2369);
or U2459 (N_2459,N_2388,N_2387);
or U2460 (N_2460,N_2406,N_2421);
nor U2461 (N_2461,N_2451,N_2400);
or U2462 (N_2462,N_2441,N_2440);
nor U2463 (N_2463,N_2402,N_2416);
or U2464 (N_2464,N_2425,N_2439);
and U2465 (N_2465,N_2444,N_2448);
and U2466 (N_2466,N_2424,N_2430);
or U2467 (N_2467,N_2438,N_2420);
nor U2468 (N_2468,N_2429,N_2442);
or U2469 (N_2469,N_2418,N_2428);
or U2470 (N_2470,N_2456,N_2422);
xnor U2471 (N_2471,N_2401,N_2407);
or U2472 (N_2472,N_2431,N_2458);
or U2473 (N_2473,N_2405,N_2454);
xnor U2474 (N_2474,N_2433,N_2445);
nand U2475 (N_2475,N_2447,N_2452);
or U2476 (N_2476,N_2414,N_2426);
xor U2477 (N_2477,N_2443,N_2427);
nor U2478 (N_2478,N_2419,N_2449);
nand U2479 (N_2479,N_2403,N_2450);
nand U2480 (N_2480,N_2455,N_2434);
nand U2481 (N_2481,N_2459,N_2411);
and U2482 (N_2482,N_2457,N_2423);
and U2483 (N_2483,N_2409,N_2413);
or U2484 (N_2484,N_2435,N_2453);
xnor U2485 (N_2485,N_2412,N_2437);
or U2486 (N_2486,N_2404,N_2410);
nor U2487 (N_2487,N_2436,N_2446);
nand U2488 (N_2488,N_2408,N_2417);
xnor U2489 (N_2489,N_2432,N_2415);
nand U2490 (N_2490,N_2433,N_2438);
or U2491 (N_2491,N_2409,N_2420);
nand U2492 (N_2492,N_2411,N_2407);
nand U2493 (N_2493,N_2407,N_2425);
or U2494 (N_2494,N_2437,N_2447);
xor U2495 (N_2495,N_2449,N_2416);
and U2496 (N_2496,N_2416,N_2446);
or U2497 (N_2497,N_2458,N_2447);
and U2498 (N_2498,N_2421,N_2400);
or U2499 (N_2499,N_2454,N_2434);
and U2500 (N_2500,N_2449,N_2436);
nand U2501 (N_2501,N_2407,N_2428);
nand U2502 (N_2502,N_2433,N_2441);
and U2503 (N_2503,N_2432,N_2405);
nand U2504 (N_2504,N_2423,N_2434);
nand U2505 (N_2505,N_2442,N_2405);
nor U2506 (N_2506,N_2432,N_2409);
and U2507 (N_2507,N_2446,N_2425);
nor U2508 (N_2508,N_2450,N_2408);
or U2509 (N_2509,N_2437,N_2400);
or U2510 (N_2510,N_2446,N_2401);
nand U2511 (N_2511,N_2441,N_2429);
and U2512 (N_2512,N_2440,N_2449);
or U2513 (N_2513,N_2402,N_2412);
nor U2514 (N_2514,N_2422,N_2416);
nand U2515 (N_2515,N_2417,N_2413);
xor U2516 (N_2516,N_2406,N_2422);
and U2517 (N_2517,N_2424,N_2440);
nor U2518 (N_2518,N_2451,N_2405);
nor U2519 (N_2519,N_2400,N_2458);
nor U2520 (N_2520,N_2495,N_2460);
nand U2521 (N_2521,N_2485,N_2500);
xnor U2522 (N_2522,N_2475,N_2499);
nor U2523 (N_2523,N_2506,N_2479);
xor U2524 (N_2524,N_2502,N_2461);
and U2525 (N_2525,N_2512,N_2519);
or U2526 (N_2526,N_2473,N_2464);
xnor U2527 (N_2527,N_2476,N_2463);
xnor U2528 (N_2528,N_2504,N_2517);
nand U2529 (N_2529,N_2468,N_2507);
nor U2530 (N_2530,N_2472,N_2505);
xnor U2531 (N_2531,N_2466,N_2513);
nor U2532 (N_2532,N_2491,N_2501);
nor U2533 (N_2533,N_2489,N_2469);
and U2534 (N_2534,N_2465,N_2471);
nand U2535 (N_2535,N_2470,N_2508);
or U2536 (N_2536,N_2511,N_2510);
or U2537 (N_2537,N_2490,N_2487);
and U2538 (N_2538,N_2480,N_2483);
and U2539 (N_2539,N_2498,N_2488);
or U2540 (N_2540,N_2474,N_2478);
nand U2541 (N_2541,N_2516,N_2515);
nand U2542 (N_2542,N_2503,N_2462);
nor U2543 (N_2543,N_2518,N_2481);
and U2544 (N_2544,N_2484,N_2514);
or U2545 (N_2545,N_2467,N_2509);
nor U2546 (N_2546,N_2477,N_2493);
nor U2547 (N_2547,N_2494,N_2492);
or U2548 (N_2548,N_2486,N_2482);
nand U2549 (N_2549,N_2496,N_2497);
nor U2550 (N_2550,N_2497,N_2473);
and U2551 (N_2551,N_2490,N_2479);
and U2552 (N_2552,N_2495,N_2514);
xnor U2553 (N_2553,N_2484,N_2496);
nor U2554 (N_2554,N_2502,N_2486);
and U2555 (N_2555,N_2466,N_2461);
nand U2556 (N_2556,N_2512,N_2484);
nor U2557 (N_2557,N_2478,N_2469);
or U2558 (N_2558,N_2512,N_2478);
xor U2559 (N_2559,N_2480,N_2513);
xor U2560 (N_2560,N_2475,N_2466);
and U2561 (N_2561,N_2488,N_2468);
nand U2562 (N_2562,N_2499,N_2506);
nor U2563 (N_2563,N_2483,N_2516);
or U2564 (N_2564,N_2513,N_2503);
nand U2565 (N_2565,N_2470,N_2498);
xor U2566 (N_2566,N_2467,N_2488);
nand U2567 (N_2567,N_2465,N_2494);
and U2568 (N_2568,N_2506,N_2475);
xor U2569 (N_2569,N_2485,N_2486);
nand U2570 (N_2570,N_2478,N_2468);
nor U2571 (N_2571,N_2473,N_2489);
nand U2572 (N_2572,N_2500,N_2470);
nand U2573 (N_2573,N_2510,N_2482);
xor U2574 (N_2574,N_2513,N_2502);
xnor U2575 (N_2575,N_2509,N_2519);
nor U2576 (N_2576,N_2490,N_2517);
nand U2577 (N_2577,N_2475,N_2514);
and U2578 (N_2578,N_2511,N_2514);
or U2579 (N_2579,N_2489,N_2474);
xor U2580 (N_2580,N_2553,N_2523);
and U2581 (N_2581,N_2528,N_2569);
or U2582 (N_2582,N_2529,N_2546);
or U2583 (N_2583,N_2551,N_2575);
or U2584 (N_2584,N_2572,N_2563);
xor U2585 (N_2585,N_2559,N_2547);
and U2586 (N_2586,N_2527,N_2576);
and U2587 (N_2587,N_2567,N_2554);
or U2588 (N_2588,N_2548,N_2561);
nand U2589 (N_2589,N_2550,N_2525);
nand U2590 (N_2590,N_2571,N_2557);
xor U2591 (N_2591,N_2524,N_2552);
nand U2592 (N_2592,N_2564,N_2573);
nand U2593 (N_2593,N_2560,N_2566);
and U2594 (N_2594,N_2574,N_2544);
or U2595 (N_2595,N_2577,N_2558);
or U2596 (N_2596,N_2568,N_2570);
nand U2597 (N_2597,N_2578,N_2533);
nor U2598 (N_2598,N_2536,N_2555);
nand U2599 (N_2599,N_2549,N_2539);
nor U2600 (N_2600,N_2542,N_2526);
xnor U2601 (N_2601,N_2537,N_2535);
or U2602 (N_2602,N_2540,N_2545);
nor U2603 (N_2603,N_2556,N_2562);
or U2604 (N_2604,N_2534,N_2520);
nand U2605 (N_2605,N_2531,N_2521);
nand U2606 (N_2606,N_2579,N_2538);
nor U2607 (N_2607,N_2541,N_2532);
nor U2608 (N_2608,N_2522,N_2565);
nand U2609 (N_2609,N_2543,N_2530);
and U2610 (N_2610,N_2559,N_2554);
or U2611 (N_2611,N_2565,N_2556);
nand U2612 (N_2612,N_2536,N_2523);
and U2613 (N_2613,N_2570,N_2524);
xnor U2614 (N_2614,N_2557,N_2544);
xnor U2615 (N_2615,N_2530,N_2558);
xnor U2616 (N_2616,N_2535,N_2545);
nand U2617 (N_2617,N_2557,N_2567);
or U2618 (N_2618,N_2534,N_2575);
nand U2619 (N_2619,N_2574,N_2528);
nand U2620 (N_2620,N_2574,N_2558);
nor U2621 (N_2621,N_2563,N_2573);
nor U2622 (N_2622,N_2570,N_2565);
or U2623 (N_2623,N_2553,N_2522);
and U2624 (N_2624,N_2540,N_2533);
nor U2625 (N_2625,N_2577,N_2543);
xnor U2626 (N_2626,N_2541,N_2539);
nand U2627 (N_2627,N_2537,N_2573);
or U2628 (N_2628,N_2551,N_2525);
and U2629 (N_2629,N_2521,N_2535);
nand U2630 (N_2630,N_2523,N_2567);
xnor U2631 (N_2631,N_2540,N_2570);
xor U2632 (N_2632,N_2576,N_2545);
or U2633 (N_2633,N_2559,N_2555);
xnor U2634 (N_2634,N_2538,N_2546);
nor U2635 (N_2635,N_2561,N_2556);
xnor U2636 (N_2636,N_2527,N_2525);
or U2637 (N_2637,N_2526,N_2536);
and U2638 (N_2638,N_2529,N_2549);
or U2639 (N_2639,N_2526,N_2568);
nor U2640 (N_2640,N_2600,N_2636);
xor U2641 (N_2641,N_2585,N_2599);
xor U2642 (N_2642,N_2622,N_2592);
nor U2643 (N_2643,N_2607,N_2618);
and U2644 (N_2644,N_2634,N_2605);
nor U2645 (N_2645,N_2609,N_2614);
and U2646 (N_2646,N_2587,N_2586);
and U2647 (N_2647,N_2594,N_2632);
or U2648 (N_2648,N_2626,N_2603);
nand U2649 (N_2649,N_2610,N_2629);
and U2650 (N_2650,N_2598,N_2619);
and U2651 (N_2651,N_2584,N_2581);
nor U2652 (N_2652,N_2593,N_2608);
nor U2653 (N_2653,N_2620,N_2639);
nor U2654 (N_2654,N_2613,N_2580);
and U2655 (N_2655,N_2623,N_2589);
nor U2656 (N_2656,N_2596,N_2637);
or U2657 (N_2657,N_2588,N_2597);
nor U2658 (N_2658,N_2621,N_2635);
xnor U2659 (N_2659,N_2615,N_2628);
and U2660 (N_2660,N_2631,N_2604);
or U2661 (N_2661,N_2630,N_2617);
and U2662 (N_2662,N_2633,N_2582);
and U2663 (N_2663,N_2616,N_2624);
nand U2664 (N_2664,N_2611,N_2595);
and U2665 (N_2665,N_2591,N_2590);
nand U2666 (N_2666,N_2627,N_2606);
or U2667 (N_2667,N_2602,N_2625);
and U2668 (N_2668,N_2601,N_2583);
or U2669 (N_2669,N_2612,N_2638);
or U2670 (N_2670,N_2635,N_2607);
nand U2671 (N_2671,N_2638,N_2583);
nand U2672 (N_2672,N_2621,N_2639);
nand U2673 (N_2673,N_2587,N_2596);
and U2674 (N_2674,N_2597,N_2614);
and U2675 (N_2675,N_2638,N_2616);
or U2676 (N_2676,N_2613,N_2627);
nor U2677 (N_2677,N_2597,N_2602);
or U2678 (N_2678,N_2621,N_2634);
nor U2679 (N_2679,N_2630,N_2629);
xnor U2680 (N_2680,N_2632,N_2599);
or U2681 (N_2681,N_2606,N_2624);
nor U2682 (N_2682,N_2629,N_2597);
xnor U2683 (N_2683,N_2620,N_2635);
nor U2684 (N_2684,N_2615,N_2609);
xnor U2685 (N_2685,N_2586,N_2623);
nor U2686 (N_2686,N_2582,N_2600);
or U2687 (N_2687,N_2585,N_2636);
or U2688 (N_2688,N_2610,N_2599);
nand U2689 (N_2689,N_2607,N_2608);
nand U2690 (N_2690,N_2593,N_2616);
xor U2691 (N_2691,N_2598,N_2638);
or U2692 (N_2692,N_2614,N_2636);
xnor U2693 (N_2693,N_2629,N_2627);
nand U2694 (N_2694,N_2586,N_2632);
and U2695 (N_2695,N_2619,N_2635);
and U2696 (N_2696,N_2580,N_2609);
nand U2697 (N_2697,N_2599,N_2613);
nand U2698 (N_2698,N_2638,N_2622);
or U2699 (N_2699,N_2617,N_2636);
xor U2700 (N_2700,N_2659,N_2664);
nand U2701 (N_2701,N_2641,N_2660);
and U2702 (N_2702,N_2694,N_2646);
nand U2703 (N_2703,N_2665,N_2662);
nand U2704 (N_2704,N_2681,N_2698);
and U2705 (N_2705,N_2674,N_2667);
xnor U2706 (N_2706,N_2657,N_2666);
nand U2707 (N_2707,N_2692,N_2686);
or U2708 (N_2708,N_2658,N_2649);
and U2709 (N_2709,N_2689,N_2679);
xor U2710 (N_2710,N_2672,N_2697);
or U2711 (N_2711,N_2684,N_2685);
or U2712 (N_2712,N_2647,N_2661);
nand U2713 (N_2713,N_2648,N_2656);
and U2714 (N_2714,N_2696,N_2695);
nor U2715 (N_2715,N_2640,N_2699);
xnor U2716 (N_2716,N_2671,N_2691);
nor U2717 (N_2717,N_2680,N_2687);
nand U2718 (N_2718,N_2669,N_2655);
and U2719 (N_2719,N_2653,N_2682);
xnor U2720 (N_2720,N_2645,N_2654);
and U2721 (N_2721,N_2690,N_2652);
xnor U2722 (N_2722,N_2688,N_2650);
nor U2723 (N_2723,N_2677,N_2678);
or U2724 (N_2724,N_2643,N_2644);
nand U2725 (N_2725,N_2642,N_2693);
nor U2726 (N_2726,N_2663,N_2676);
xnor U2727 (N_2727,N_2683,N_2673);
xor U2728 (N_2728,N_2668,N_2675);
nand U2729 (N_2729,N_2651,N_2670);
xnor U2730 (N_2730,N_2683,N_2684);
nor U2731 (N_2731,N_2644,N_2653);
or U2732 (N_2732,N_2669,N_2644);
nand U2733 (N_2733,N_2647,N_2682);
or U2734 (N_2734,N_2645,N_2699);
xnor U2735 (N_2735,N_2672,N_2650);
nor U2736 (N_2736,N_2683,N_2650);
nand U2737 (N_2737,N_2656,N_2699);
xnor U2738 (N_2738,N_2682,N_2698);
nand U2739 (N_2739,N_2668,N_2644);
nor U2740 (N_2740,N_2644,N_2670);
nor U2741 (N_2741,N_2655,N_2692);
nand U2742 (N_2742,N_2688,N_2680);
nand U2743 (N_2743,N_2647,N_2652);
and U2744 (N_2744,N_2657,N_2654);
and U2745 (N_2745,N_2677,N_2646);
nand U2746 (N_2746,N_2698,N_2655);
xnor U2747 (N_2747,N_2667,N_2676);
nand U2748 (N_2748,N_2666,N_2640);
nand U2749 (N_2749,N_2683,N_2654);
nor U2750 (N_2750,N_2672,N_2674);
and U2751 (N_2751,N_2691,N_2680);
xor U2752 (N_2752,N_2697,N_2661);
and U2753 (N_2753,N_2666,N_2651);
nand U2754 (N_2754,N_2663,N_2680);
and U2755 (N_2755,N_2666,N_2660);
xnor U2756 (N_2756,N_2691,N_2660);
nor U2757 (N_2757,N_2690,N_2693);
nor U2758 (N_2758,N_2647,N_2674);
or U2759 (N_2759,N_2673,N_2686);
nand U2760 (N_2760,N_2741,N_2748);
xor U2761 (N_2761,N_2732,N_2733);
xnor U2762 (N_2762,N_2708,N_2736);
and U2763 (N_2763,N_2705,N_2709);
or U2764 (N_2764,N_2707,N_2717);
nand U2765 (N_2765,N_2716,N_2718);
nor U2766 (N_2766,N_2711,N_2702);
nand U2767 (N_2767,N_2720,N_2751);
nor U2768 (N_2768,N_2747,N_2759);
xnor U2769 (N_2769,N_2738,N_2719);
and U2770 (N_2770,N_2737,N_2726);
or U2771 (N_2771,N_2706,N_2710);
nor U2772 (N_2772,N_2725,N_2727);
or U2773 (N_2773,N_2712,N_2722);
and U2774 (N_2774,N_2701,N_2743);
nand U2775 (N_2775,N_2703,N_2704);
nor U2776 (N_2776,N_2729,N_2745);
nand U2777 (N_2777,N_2735,N_2721);
nand U2778 (N_2778,N_2746,N_2730);
nor U2779 (N_2779,N_2728,N_2755);
nor U2780 (N_2780,N_2749,N_2740);
xor U2781 (N_2781,N_2714,N_2734);
and U2782 (N_2782,N_2753,N_2724);
nor U2783 (N_2783,N_2723,N_2713);
or U2784 (N_2784,N_2758,N_2715);
nor U2785 (N_2785,N_2731,N_2700);
and U2786 (N_2786,N_2742,N_2756);
and U2787 (N_2787,N_2750,N_2757);
xnor U2788 (N_2788,N_2739,N_2752);
nand U2789 (N_2789,N_2754,N_2744);
nor U2790 (N_2790,N_2749,N_2756);
and U2791 (N_2791,N_2731,N_2738);
or U2792 (N_2792,N_2722,N_2733);
and U2793 (N_2793,N_2757,N_2738);
and U2794 (N_2794,N_2749,N_2746);
nor U2795 (N_2795,N_2727,N_2704);
nand U2796 (N_2796,N_2725,N_2735);
or U2797 (N_2797,N_2754,N_2742);
or U2798 (N_2798,N_2749,N_2726);
xnor U2799 (N_2799,N_2740,N_2741);
nor U2800 (N_2800,N_2743,N_2711);
nand U2801 (N_2801,N_2715,N_2742);
nor U2802 (N_2802,N_2754,N_2711);
and U2803 (N_2803,N_2726,N_2744);
and U2804 (N_2804,N_2718,N_2733);
nand U2805 (N_2805,N_2734,N_2723);
nand U2806 (N_2806,N_2742,N_2700);
and U2807 (N_2807,N_2741,N_2750);
nand U2808 (N_2808,N_2713,N_2759);
nor U2809 (N_2809,N_2737,N_2725);
and U2810 (N_2810,N_2719,N_2706);
xnor U2811 (N_2811,N_2753,N_2721);
and U2812 (N_2812,N_2750,N_2724);
or U2813 (N_2813,N_2723,N_2743);
or U2814 (N_2814,N_2701,N_2741);
and U2815 (N_2815,N_2739,N_2751);
nand U2816 (N_2816,N_2725,N_2721);
or U2817 (N_2817,N_2739,N_2711);
nand U2818 (N_2818,N_2759,N_2738);
nor U2819 (N_2819,N_2738,N_2732);
nor U2820 (N_2820,N_2797,N_2776);
and U2821 (N_2821,N_2761,N_2771);
nand U2822 (N_2822,N_2769,N_2788);
nor U2823 (N_2823,N_2793,N_2780);
xnor U2824 (N_2824,N_2803,N_2790);
or U2825 (N_2825,N_2775,N_2765);
nand U2826 (N_2826,N_2777,N_2784);
nand U2827 (N_2827,N_2812,N_2807);
xnor U2828 (N_2828,N_2763,N_2782);
nand U2829 (N_2829,N_2785,N_2798);
or U2830 (N_2830,N_2813,N_2770);
and U2831 (N_2831,N_2815,N_2773);
xnor U2832 (N_2832,N_2809,N_2791);
nand U2833 (N_2833,N_2760,N_2801);
nand U2834 (N_2834,N_2814,N_2778);
and U2835 (N_2835,N_2764,N_2800);
or U2836 (N_2836,N_2819,N_2817);
and U2837 (N_2837,N_2796,N_2772);
or U2838 (N_2838,N_2794,N_2789);
or U2839 (N_2839,N_2802,N_2804);
or U2840 (N_2840,N_2781,N_2767);
nand U2841 (N_2841,N_2810,N_2766);
nand U2842 (N_2842,N_2816,N_2806);
and U2843 (N_2843,N_2799,N_2811);
nand U2844 (N_2844,N_2787,N_2762);
nor U2845 (N_2845,N_2779,N_2783);
nand U2846 (N_2846,N_2774,N_2795);
or U2847 (N_2847,N_2818,N_2805);
nor U2848 (N_2848,N_2786,N_2792);
xor U2849 (N_2849,N_2768,N_2808);
and U2850 (N_2850,N_2809,N_2766);
and U2851 (N_2851,N_2776,N_2795);
xnor U2852 (N_2852,N_2782,N_2772);
xnor U2853 (N_2853,N_2809,N_2799);
xor U2854 (N_2854,N_2772,N_2763);
and U2855 (N_2855,N_2816,N_2795);
nand U2856 (N_2856,N_2809,N_2761);
nor U2857 (N_2857,N_2806,N_2780);
and U2858 (N_2858,N_2808,N_2793);
nor U2859 (N_2859,N_2790,N_2818);
and U2860 (N_2860,N_2762,N_2819);
nand U2861 (N_2861,N_2790,N_2771);
nor U2862 (N_2862,N_2791,N_2771);
nor U2863 (N_2863,N_2796,N_2780);
nor U2864 (N_2864,N_2770,N_2817);
or U2865 (N_2865,N_2814,N_2809);
or U2866 (N_2866,N_2787,N_2773);
nand U2867 (N_2867,N_2769,N_2767);
or U2868 (N_2868,N_2796,N_2779);
nor U2869 (N_2869,N_2811,N_2789);
nor U2870 (N_2870,N_2770,N_2784);
nand U2871 (N_2871,N_2765,N_2764);
nor U2872 (N_2872,N_2810,N_2804);
and U2873 (N_2873,N_2774,N_2779);
and U2874 (N_2874,N_2779,N_2773);
nor U2875 (N_2875,N_2819,N_2777);
or U2876 (N_2876,N_2776,N_2798);
and U2877 (N_2877,N_2806,N_2762);
and U2878 (N_2878,N_2804,N_2796);
xor U2879 (N_2879,N_2791,N_2766);
nand U2880 (N_2880,N_2829,N_2840);
and U2881 (N_2881,N_2870,N_2859);
nand U2882 (N_2882,N_2866,N_2856);
or U2883 (N_2883,N_2855,N_2825);
or U2884 (N_2884,N_2867,N_2847);
nor U2885 (N_2885,N_2833,N_2852);
or U2886 (N_2886,N_2853,N_2874);
nand U2887 (N_2887,N_2872,N_2834);
and U2888 (N_2888,N_2845,N_2846);
nor U2889 (N_2889,N_2832,N_2841);
or U2890 (N_2890,N_2828,N_2843);
and U2891 (N_2891,N_2826,N_2851);
nor U2892 (N_2892,N_2862,N_2842);
or U2893 (N_2893,N_2863,N_2850);
nor U2894 (N_2894,N_2830,N_2854);
xnor U2895 (N_2895,N_2821,N_2824);
and U2896 (N_2896,N_2836,N_2844);
and U2897 (N_2897,N_2875,N_2868);
or U2898 (N_2898,N_2860,N_2869);
or U2899 (N_2899,N_2865,N_2858);
nand U2900 (N_2900,N_2827,N_2835);
and U2901 (N_2901,N_2857,N_2822);
nor U2902 (N_2902,N_2873,N_2876);
nor U2903 (N_2903,N_2861,N_2838);
and U2904 (N_2904,N_2879,N_2871);
xnor U2905 (N_2905,N_2823,N_2839);
nor U2906 (N_2906,N_2837,N_2820);
xor U2907 (N_2907,N_2831,N_2848);
or U2908 (N_2908,N_2849,N_2864);
xnor U2909 (N_2909,N_2878,N_2877);
nor U2910 (N_2910,N_2822,N_2877);
nand U2911 (N_2911,N_2870,N_2833);
or U2912 (N_2912,N_2823,N_2861);
and U2913 (N_2913,N_2828,N_2846);
and U2914 (N_2914,N_2836,N_2853);
nor U2915 (N_2915,N_2841,N_2874);
xnor U2916 (N_2916,N_2852,N_2832);
xor U2917 (N_2917,N_2836,N_2856);
and U2918 (N_2918,N_2863,N_2834);
nand U2919 (N_2919,N_2876,N_2867);
and U2920 (N_2920,N_2853,N_2828);
or U2921 (N_2921,N_2835,N_2874);
and U2922 (N_2922,N_2858,N_2822);
and U2923 (N_2923,N_2820,N_2865);
xor U2924 (N_2924,N_2838,N_2820);
xor U2925 (N_2925,N_2876,N_2859);
and U2926 (N_2926,N_2859,N_2829);
nand U2927 (N_2927,N_2854,N_2860);
nor U2928 (N_2928,N_2856,N_2830);
and U2929 (N_2929,N_2839,N_2857);
xnor U2930 (N_2930,N_2865,N_2842);
or U2931 (N_2931,N_2876,N_2878);
and U2932 (N_2932,N_2832,N_2839);
nand U2933 (N_2933,N_2844,N_2873);
or U2934 (N_2934,N_2842,N_2827);
and U2935 (N_2935,N_2865,N_2860);
and U2936 (N_2936,N_2844,N_2858);
nor U2937 (N_2937,N_2874,N_2823);
nand U2938 (N_2938,N_2841,N_2861);
xor U2939 (N_2939,N_2838,N_2833);
or U2940 (N_2940,N_2902,N_2921);
and U2941 (N_2941,N_2925,N_2884);
or U2942 (N_2942,N_2909,N_2908);
nor U2943 (N_2943,N_2919,N_2913);
nor U2944 (N_2944,N_2892,N_2934);
nor U2945 (N_2945,N_2895,N_2910);
nand U2946 (N_2946,N_2929,N_2880);
or U2947 (N_2947,N_2915,N_2927);
and U2948 (N_2948,N_2914,N_2905);
nand U2949 (N_2949,N_2897,N_2907);
or U2950 (N_2950,N_2899,N_2893);
nor U2951 (N_2951,N_2922,N_2900);
xor U2952 (N_2952,N_2932,N_2917);
or U2953 (N_2953,N_2916,N_2911);
xor U2954 (N_2954,N_2933,N_2920);
or U2955 (N_2955,N_2938,N_2918);
and U2956 (N_2956,N_2891,N_2901);
nor U2957 (N_2957,N_2898,N_2939);
nor U2958 (N_2958,N_2887,N_2883);
and U2959 (N_2959,N_2928,N_2936);
nor U2960 (N_2960,N_2923,N_2935);
or U2961 (N_2961,N_2926,N_2903);
nor U2962 (N_2962,N_2924,N_2882);
or U2963 (N_2963,N_2937,N_2906);
nor U2964 (N_2964,N_2931,N_2912);
and U2965 (N_2965,N_2886,N_2889);
nor U2966 (N_2966,N_2885,N_2930);
nor U2967 (N_2967,N_2904,N_2896);
xor U2968 (N_2968,N_2881,N_2890);
nor U2969 (N_2969,N_2894,N_2888);
xnor U2970 (N_2970,N_2934,N_2884);
nand U2971 (N_2971,N_2910,N_2930);
and U2972 (N_2972,N_2931,N_2907);
xor U2973 (N_2973,N_2915,N_2938);
nand U2974 (N_2974,N_2893,N_2925);
nand U2975 (N_2975,N_2928,N_2886);
or U2976 (N_2976,N_2891,N_2907);
xor U2977 (N_2977,N_2932,N_2928);
and U2978 (N_2978,N_2919,N_2911);
nand U2979 (N_2979,N_2919,N_2903);
xor U2980 (N_2980,N_2891,N_2911);
and U2981 (N_2981,N_2927,N_2935);
and U2982 (N_2982,N_2919,N_2882);
xnor U2983 (N_2983,N_2925,N_2923);
or U2984 (N_2984,N_2938,N_2916);
or U2985 (N_2985,N_2928,N_2920);
and U2986 (N_2986,N_2886,N_2909);
nand U2987 (N_2987,N_2919,N_2917);
nor U2988 (N_2988,N_2893,N_2916);
and U2989 (N_2989,N_2884,N_2881);
nor U2990 (N_2990,N_2892,N_2909);
nor U2991 (N_2991,N_2898,N_2924);
nand U2992 (N_2992,N_2929,N_2912);
xor U2993 (N_2993,N_2937,N_2929);
or U2994 (N_2994,N_2906,N_2899);
nor U2995 (N_2995,N_2885,N_2907);
or U2996 (N_2996,N_2893,N_2900);
nor U2997 (N_2997,N_2883,N_2884);
nor U2998 (N_2998,N_2929,N_2902);
nand U2999 (N_2999,N_2920,N_2931);
and UO_0 (O_0,N_2955,N_2948);
or UO_1 (O_1,N_2990,N_2952);
nor UO_2 (O_2,N_2947,N_2970);
or UO_3 (O_3,N_2941,N_2996);
nor UO_4 (O_4,N_2979,N_2968);
and UO_5 (O_5,N_2956,N_2950);
or UO_6 (O_6,N_2991,N_2974);
and UO_7 (O_7,N_2945,N_2980);
or UO_8 (O_8,N_2957,N_2983);
nand UO_9 (O_9,N_2982,N_2997);
nor UO_10 (O_10,N_2972,N_2961);
nor UO_11 (O_11,N_2964,N_2989);
or UO_12 (O_12,N_2973,N_2943);
and UO_13 (O_13,N_2986,N_2954);
xnor UO_14 (O_14,N_2962,N_2969);
nand UO_15 (O_15,N_2966,N_2953);
or UO_16 (O_16,N_2975,N_2958);
xnor UO_17 (O_17,N_2960,N_2959);
and UO_18 (O_18,N_2951,N_2971);
and UO_19 (O_19,N_2981,N_2963);
nor UO_20 (O_20,N_2965,N_2993);
and UO_21 (O_21,N_2994,N_2977);
xor UO_22 (O_22,N_2940,N_2946);
nor UO_23 (O_23,N_2988,N_2985);
xnor UO_24 (O_24,N_2949,N_2998);
and UO_25 (O_25,N_2967,N_2987);
xnor UO_26 (O_26,N_2984,N_2978);
xnor UO_27 (O_27,N_2999,N_2976);
nor UO_28 (O_28,N_2992,N_2942);
xor UO_29 (O_29,N_2995,N_2944);
xor UO_30 (O_30,N_2949,N_2971);
and UO_31 (O_31,N_2970,N_2948);
or UO_32 (O_32,N_2976,N_2975);
or UO_33 (O_33,N_2997,N_2946);
xor UO_34 (O_34,N_2999,N_2987);
or UO_35 (O_35,N_2972,N_2948);
xnor UO_36 (O_36,N_2959,N_2973);
or UO_37 (O_37,N_2947,N_2964);
nand UO_38 (O_38,N_2983,N_2988);
and UO_39 (O_39,N_2976,N_2950);
xnor UO_40 (O_40,N_2979,N_2953);
or UO_41 (O_41,N_2972,N_2987);
xor UO_42 (O_42,N_2986,N_2943);
nor UO_43 (O_43,N_2969,N_2942);
xnor UO_44 (O_44,N_2995,N_2991);
nor UO_45 (O_45,N_2971,N_2999);
or UO_46 (O_46,N_2944,N_2954);
nand UO_47 (O_47,N_2941,N_2969);
or UO_48 (O_48,N_2981,N_2991);
and UO_49 (O_49,N_2979,N_2978);
and UO_50 (O_50,N_2993,N_2995);
nand UO_51 (O_51,N_2973,N_2992);
nor UO_52 (O_52,N_2943,N_2964);
or UO_53 (O_53,N_2991,N_2962);
nor UO_54 (O_54,N_2983,N_2952);
xor UO_55 (O_55,N_2951,N_2969);
nand UO_56 (O_56,N_2970,N_2943);
or UO_57 (O_57,N_2941,N_2944);
and UO_58 (O_58,N_2982,N_2957);
and UO_59 (O_59,N_2979,N_2981);
nand UO_60 (O_60,N_2974,N_2995);
nand UO_61 (O_61,N_2945,N_2970);
nand UO_62 (O_62,N_2969,N_2943);
xnor UO_63 (O_63,N_2976,N_2949);
xnor UO_64 (O_64,N_2948,N_2988);
and UO_65 (O_65,N_2970,N_2956);
xor UO_66 (O_66,N_2958,N_2972);
nor UO_67 (O_67,N_2943,N_2995);
and UO_68 (O_68,N_2945,N_2941);
or UO_69 (O_69,N_2993,N_2951);
or UO_70 (O_70,N_2958,N_2945);
xnor UO_71 (O_71,N_2964,N_2969);
nor UO_72 (O_72,N_2999,N_2982);
or UO_73 (O_73,N_2993,N_2950);
nor UO_74 (O_74,N_2979,N_2988);
nor UO_75 (O_75,N_2977,N_2973);
nor UO_76 (O_76,N_2977,N_2957);
and UO_77 (O_77,N_2949,N_2943);
nor UO_78 (O_78,N_2977,N_2988);
nor UO_79 (O_79,N_2946,N_2953);
xnor UO_80 (O_80,N_2984,N_2979);
or UO_81 (O_81,N_2962,N_2946);
xnor UO_82 (O_82,N_2944,N_2998);
xor UO_83 (O_83,N_2955,N_2994);
nand UO_84 (O_84,N_2975,N_2995);
xor UO_85 (O_85,N_2990,N_2964);
nand UO_86 (O_86,N_2958,N_2981);
or UO_87 (O_87,N_2968,N_2959);
xor UO_88 (O_88,N_2960,N_2984);
nand UO_89 (O_89,N_2957,N_2954);
or UO_90 (O_90,N_2954,N_2987);
or UO_91 (O_91,N_2976,N_2986);
and UO_92 (O_92,N_2963,N_2992);
and UO_93 (O_93,N_2971,N_2991);
nor UO_94 (O_94,N_2981,N_2982);
nor UO_95 (O_95,N_2983,N_2940);
nand UO_96 (O_96,N_2945,N_2995);
and UO_97 (O_97,N_2955,N_2954);
nand UO_98 (O_98,N_2977,N_2965);
xnor UO_99 (O_99,N_2940,N_2975);
nor UO_100 (O_100,N_2995,N_2965);
xor UO_101 (O_101,N_2994,N_2970);
nand UO_102 (O_102,N_2965,N_2941);
xor UO_103 (O_103,N_2957,N_2976);
or UO_104 (O_104,N_2979,N_2955);
nor UO_105 (O_105,N_2980,N_2965);
or UO_106 (O_106,N_2998,N_2988);
nor UO_107 (O_107,N_2985,N_2942);
nor UO_108 (O_108,N_2952,N_2951);
nor UO_109 (O_109,N_2955,N_2963);
nor UO_110 (O_110,N_2998,N_2996);
nor UO_111 (O_111,N_2985,N_2964);
nand UO_112 (O_112,N_2950,N_2999);
or UO_113 (O_113,N_2985,N_2941);
nor UO_114 (O_114,N_2977,N_2967);
and UO_115 (O_115,N_2958,N_2999);
or UO_116 (O_116,N_2991,N_2990);
and UO_117 (O_117,N_2979,N_2985);
or UO_118 (O_118,N_2967,N_2980);
or UO_119 (O_119,N_2990,N_2956);
nor UO_120 (O_120,N_2966,N_2984);
xnor UO_121 (O_121,N_2989,N_2952);
nand UO_122 (O_122,N_2970,N_2951);
nand UO_123 (O_123,N_2989,N_2996);
or UO_124 (O_124,N_2997,N_2942);
nor UO_125 (O_125,N_2955,N_2953);
or UO_126 (O_126,N_2975,N_2949);
or UO_127 (O_127,N_2989,N_2995);
nor UO_128 (O_128,N_2964,N_2970);
nor UO_129 (O_129,N_2985,N_2971);
xor UO_130 (O_130,N_2986,N_2993);
nor UO_131 (O_131,N_2976,N_2947);
and UO_132 (O_132,N_2994,N_2967);
nor UO_133 (O_133,N_2946,N_2942);
and UO_134 (O_134,N_2942,N_2977);
xor UO_135 (O_135,N_2990,N_2975);
and UO_136 (O_136,N_2965,N_2978);
nor UO_137 (O_137,N_2960,N_2989);
nand UO_138 (O_138,N_2995,N_2940);
nand UO_139 (O_139,N_2987,N_2948);
nand UO_140 (O_140,N_2972,N_2997);
or UO_141 (O_141,N_2999,N_2966);
or UO_142 (O_142,N_2947,N_2991);
nand UO_143 (O_143,N_2969,N_2985);
and UO_144 (O_144,N_2943,N_2991);
and UO_145 (O_145,N_2979,N_2994);
or UO_146 (O_146,N_2965,N_2972);
nor UO_147 (O_147,N_2981,N_2944);
and UO_148 (O_148,N_2949,N_2951);
and UO_149 (O_149,N_2985,N_2989);
nor UO_150 (O_150,N_2976,N_2984);
xor UO_151 (O_151,N_2942,N_2956);
xnor UO_152 (O_152,N_2968,N_2997);
xor UO_153 (O_153,N_2997,N_2989);
and UO_154 (O_154,N_2955,N_2960);
or UO_155 (O_155,N_2997,N_2983);
xor UO_156 (O_156,N_2958,N_2969);
or UO_157 (O_157,N_2970,N_2993);
and UO_158 (O_158,N_2961,N_2993);
xor UO_159 (O_159,N_2955,N_2965);
or UO_160 (O_160,N_2976,N_2942);
or UO_161 (O_161,N_2974,N_2990);
or UO_162 (O_162,N_2976,N_2966);
or UO_163 (O_163,N_2980,N_2947);
xor UO_164 (O_164,N_2961,N_2959);
nor UO_165 (O_165,N_2970,N_2942);
nor UO_166 (O_166,N_2941,N_2999);
xor UO_167 (O_167,N_2994,N_2973);
or UO_168 (O_168,N_2992,N_2978);
and UO_169 (O_169,N_2993,N_2974);
nor UO_170 (O_170,N_2960,N_2946);
and UO_171 (O_171,N_2972,N_2988);
nor UO_172 (O_172,N_2959,N_2987);
nor UO_173 (O_173,N_2969,N_2988);
nand UO_174 (O_174,N_2980,N_2940);
or UO_175 (O_175,N_2943,N_2976);
or UO_176 (O_176,N_2951,N_2972);
nand UO_177 (O_177,N_2940,N_2961);
or UO_178 (O_178,N_2953,N_2950);
and UO_179 (O_179,N_2947,N_2993);
nand UO_180 (O_180,N_2960,N_2945);
and UO_181 (O_181,N_2962,N_2945);
nor UO_182 (O_182,N_2985,N_2977);
nand UO_183 (O_183,N_2987,N_2983);
nor UO_184 (O_184,N_2972,N_2978);
nand UO_185 (O_185,N_2955,N_2949);
nor UO_186 (O_186,N_2948,N_2947);
nor UO_187 (O_187,N_2950,N_2974);
or UO_188 (O_188,N_2999,N_2993);
nor UO_189 (O_189,N_2993,N_2980);
or UO_190 (O_190,N_2956,N_2946);
or UO_191 (O_191,N_2943,N_2996);
nand UO_192 (O_192,N_2967,N_2955);
and UO_193 (O_193,N_2948,N_2994);
or UO_194 (O_194,N_2987,N_2977);
or UO_195 (O_195,N_2978,N_2953);
nand UO_196 (O_196,N_2992,N_2956);
or UO_197 (O_197,N_2997,N_2978);
xnor UO_198 (O_198,N_2993,N_2984);
and UO_199 (O_199,N_2955,N_2964);
nor UO_200 (O_200,N_2967,N_2969);
nand UO_201 (O_201,N_2986,N_2990);
nor UO_202 (O_202,N_2944,N_2955);
and UO_203 (O_203,N_2984,N_2998);
nand UO_204 (O_204,N_2975,N_2969);
nor UO_205 (O_205,N_2962,N_2971);
nand UO_206 (O_206,N_2991,N_2992);
and UO_207 (O_207,N_2961,N_2971);
nor UO_208 (O_208,N_2964,N_2956);
or UO_209 (O_209,N_2959,N_2988);
and UO_210 (O_210,N_2964,N_2948);
nor UO_211 (O_211,N_2989,N_2992);
nand UO_212 (O_212,N_2971,N_2992);
nor UO_213 (O_213,N_2945,N_2979);
xnor UO_214 (O_214,N_2952,N_2986);
and UO_215 (O_215,N_2957,N_2981);
or UO_216 (O_216,N_2978,N_2985);
nor UO_217 (O_217,N_2965,N_2947);
xnor UO_218 (O_218,N_2962,N_2944);
or UO_219 (O_219,N_2972,N_2999);
nor UO_220 (O_220,N_2985,N_2949);
xnor UO_221 (O_221,N_2964,N_2940);
and UO_222 (O_222,N_2996,N_2961);
nor UO_223 (O_223,N_2973,N_2976);
or UO_224 (O_224,N_2975,N_2964);
xor UO_225 (O_225,N_2952,N_2944);
nor UO_226 (O_226,N_2942,N_2993);
xor UO_227 (O_227,N_2965,N_2984);
nand UO_228 (O_228,N_2979,N_2989);
or UO_229 (O_229,N_2977,N_2989);
nor UO_230 (O_230,N_2992,N_2968);
or UO_231 (O_231,N_2948,N_2958);
xnor UO_232 (O_232,N_2999,N_2943);
nand UO_233 (O_233,N_2957,N_2979);
nand UO_234 (O_234,N_2990,N_2994);
nand UO_235 (O_235,N_2953,N_2987);
or UO_236 (O_236,N_2957,N_2969);
nor UO_237 (O_237,N_2991,N_2960);
or UO_238 (O_238,N_2967,N_2972);
nor UO_239 (O_239,N_2999,N_2992);
xor UO_240 (O_240,N_2943,N_2946);
xor UO_241 (O_241,N_2982,N_2950);
nor UO_242 (O_242,N_2980,N_2941);
xnor UO_243 (O_243,N_2958,N_2946);
and UO_244 (O_244,N_2969,N_2996);
nand UO_245 (O_245,N_2984,N_2967);
nor UO_246 (O_246,N_2951,N_2943);
nand UO_247 (O_247,N_2988,N_2950);
nand UO_248 (O_248,N_2998,N_2954);
xnor UO_249 (O_249,N_2968,N_2988);
and UO_250 (O_250,N_2954,N_2999);
nand UO_251 (O_251,N_2971,N_2980);
and UO_252 (O_252,N_2944,N_2964);
and UO_253 (O_253,N_2948,N_2979);
nor UO_254 (O_254,N_2961,N_2974);
or UO_255 (O_255,N_2966,N_2998);
nand UO_256 (O_256,N_2958,N_2982);
nand UO_257 (O_257,N_2979,N_2982);
nand UO_258 (O_258,N_2957,N_2944);
nand UO_259 (O_259,N_2985,N_2945);
or UO_260 (O_260,N_2988,N_2973);
nor UO_261 (O_261,N_2978,N_2952);
nand UO_262 (O_262,N_2984,N_2956);
nor UO_263 (O_263,N_2969,N_2944);
and UO_264 (O_264,N_2976,N_2960);
xnor UO_265 (O_265,N_2973,N_2956);
nand UO_266 (O_266,N_2990,N_2971);
and UO_267 (O_267,N_2978,N_2970);
or UO_268 (O_268,N_2946,N_2989);
nand UO_269 (O_269,N_2973,N_2984);
nor UO_270 (O_270,N_2956,N_2951);
xnor UO_271 (O_271,N_2962,N_2940);
xnor UO_272 (O_272,N_2976,N_2985);
nor UO_273 (O_273,N_2983,N_2984);
nand UO_274 (O_274,N_2988,N_2970);
nand UO_275 (O_275,N_2971,N_2953);
and UO_276 (O_276,N_2988,N_2994);
nand UO_277 (O_277,N_2966,N_2951);
or UO_278 (O_278,N_2990,N_2948);
xor UO_279 (O_279,N_2984,N_2964);
nand UO_280 (O_280,N_2979,N_2963);
xor UO_281 (O_281,N_2991,N_2978);
and UO_282 (O_282,N_2962,N_2993);
or UO_283 (O_283,N_2951,N_2955);
nand UO_284 (O_284,N_2981,N_2959);
xnor UO_285 (O_285,N_2986,N_2991);
or UO_286 (O_286,N_2974,N_2992);
and UO_287 (O_287,N_2950,N_2965);
and UO_288 (O_288,N_2993,N_2969);
xnor UO_289 (O_289,N_2973,N_2969);
nor UO_290 (O_290,N_2995,N_2942);
xnor UO_291 (O_291,N_2983,N_2982);
and UO_292 (O_292,N_2982,N_2965);
and UO_293 (O_293,N_2994,N_2975);
nand UO_294 (O_294,N_2996,N_2940);
xor UO_295 (O_295,N_2942,N_2962);
nand UO_296 (O_296,N_2974,N_2940);
xor UO_297 (O_297,N_2990,N_2995);
xor UO_298 (O_298,N_2951,N_2995);
and UO_299 (O_299,N_2960,N_2982);
xnor UO_300 (O_300,N_2987,N_2973);
and UO_301 (O_301,N_2962,N_2954);
xnor UO_302 (O_302,N_2973,N_2951);
nand UO_303 (O_303,N_2968,N_2941);
nand UO_304 (O_304,N_2995,N_2958);
nand UO_305 (O_305,N_2947,N_2952);
and UO_306 (O_306,N_2963,N_2941);
nor UO_307 (O_307,N_2973,N_2966);
and UO_308 (O_308,N_2987,N_2965);
or UO_309 (O_309,N_2955,N_2993);
or UO_310 (O_310,N_2956,N_2987);
xnor UO_311 (O_311,N_2960,N_2980);
or UO_312 (O_312,N_2994,N_2957);
nor UO_313 (O_313,N_2990,N_2953);
or UO_314 (O_314,N_2942,N_2966);
xnor UO_315 (O_315,N_2985,N_2954);
xor UO_316 (O_316,N_2960,N_2941);
xor UO_317 (O_317,N_2990,N_2967);
and UO_318 (O_318,N_2970,N_2982);
and UO_319 (O_319,N_2947,N_2944);
xor UO_320 (O_320,N_2954,N_2943);
nand UO_321 (O_321,N_2953,N_2988);
xnor UO_322 (O_322,N_2941,N_2967);
xnor UO_323 (O_323,N_2964,N_2965);
xnor UO_324 (O_324,N_2976,N_2963);
nand UO_325 (O_325,N_2973,N_2947);
nand UO_326 (O_326,N_2990,N_2954);
nand UO_327 (O_327,N_2969,N_2946);
or UO_328 (O_328,N_2978,N_2946);
nor UO_329 (O_329,N_2942,N_2991);
nor UO_330 (O_330,N_2952,N_2977);
or UO_331 (O_331,N_2958,N_2984);
and UO_332 (O_332,N_2950,N_2969);
or UO_333 (O_333,N_2940,N_2989);
nand UO_334 (O_334,N_2962,N_2983);
nand UO_335 (O_335,N_2973,N_2989);
nor UO_336 (O_336,N_2994,N_2983);
or UO_337 (O_337,N_2993,N_2966);
and UO_338 (O_338,N_2956,N_2941);
and UO_339 (O_339,N_2945,N_2989);
nand UO_340 (O_340,N_2999,N_2994);
or UO_341 (O_341,N_2965,N_2973);
nand UO_342 (O_342,N_2969,N_2966);
or UO_343 (O_343,N_2963,N_2951);
nand UO_344 (O_344,N_2985,N_2961);
nand UO_345 (O_345,N_2974,N_2942);
or UO_346 (O_346,N_2963,N_2946);
nand UO_347 (O_347,N_2956,N_2999);
nand UO_348 (O_348,N_2951,N_2965);
or UO_349 (O_349,N_2998,N_2942);
nor UO_350 (O_350,N_2971,N_2972);
nor UO_351 (O_351,N_2983,N_2972);
xnor UO_352 (O_352,N_2978,N_2998);
or UO_353 (O_353,N_2959,N_2978);
or UO_354 (O_354,N_2950,N_2943);
and UO_355 (O_355,N_2968,N_2951);
or UO_356 (O_356,N_2977,N_2997);
nand UO_357 (O_357,N_2953,N_2960);
or UO_358 (O_358,N_2981,N_2964);
nor UO_359 (O_359,N_2979,N_2969);
and UO_360 (O_360,N_2984,N_2943);
nand UO_361 (O_361,N_2996,N_2945);
and UO_362 (O_362,N_2969,N_2992);
nand UO_363 (O_363,N_2964,N_2976);
xor UO_364 (O_364,N_2985,N_2943);
xor UO_365 (O_365,N_2961,N_2978);
xnor UO_366 (O_366,N_2968,N_2971);
and UO_367 (O_367,N_2981,N_2978);
xnor UO_368 (O_368,N_2954,N_2948);
nand UO_369 (O_369,N_2993,N_2991);
nand UO_370 (O_370,N_2971,N_2989);
xor UO_371 (O_371,N_2959,N_2992);
and UO_372 (O_372,N_2979,N_2995);
or UO_373 (O_373,N_2946,N_2957);
xor UO_374 (O_374,N_2946,N_2991);
or UO_375 (O_375,N_2954,N_2988);
xnor UO_376 (O_376,N_2948,N_2942);
and UO_377 (O_377,N_2948,N_2991);
and UO_378 (O_378,N_2945,N_2963);
and UO_379 (O_379,N_2957,N_2988);
xnor UO_380 (O_380,N_2942,N_2971);
and UO_381 (O_381,N_2983,N_2985);
nor UO_382 (O_382,N_2997,N_2965);
nand UO_383 (O_383,N_2964,N_2950);
or UO_384 (O_384,N_2968,N_2962);
and UO_385 (O_385,N_2986,N_2982);
nand UO_386 (O_386,N_2973,N_2953);
xor UO_387 (O_387,N_2974,N_2988);
or UO_388 (O_388,N_2991,N_2955);
xnor UO_389 (O_389,N_2983,N_2944);
xnor UO_390 (O_390,N_2942,N_2958);
and UO_391 (O_391,N_2951,N_2984);
nor UO_392 (O_392,N_2954,N_2968);
nand UO_393 (O_393,N_2985,N_2997);
or UO_394 (O_394,N_2983,N_2966);
nand UO_395 (O_395,N_2951,N_2961);
nand UO_396 (O_396,N_2943,N_2947);
or UO_397 (O_397,N_2991,N_2967);
and UO_398 (O_398,N_2957,N_2997);
xnor UO_399 (O_399,N_2990,N_2959);
or UO_400 (O_400,N_2984,N_2974);
xor UO_401 (O_401,N_2956,N_2994);
nand UO_402 (O_402,N_2995,N_2956);
xor UO_403 (O_403,N_2975,N_2987);
and UO_404 (O_404,N_2959,N_2957);
nor UO_405 (O_405,N_2946,N_2971);
or UO_406 (O_406,N_2975,N_2980);
nand UO_407 (O_407,N_2948,N_2999);
nand UO_408 (O_408,N_2979,N_2986);
and UO_409 (O_409,N_2988,N_2987);
nand UO_410 (O_410,N_2954,N_2949);
and UO_411 (O_411,N_2969,N_2997);
nand UO_412 (O_412,N_2968,N_2977);
nor UO_413 (O_413,N_2978,N_2999);
and UO_414 (O_414,N_2983,N_2959);
or UO_415 (O_415,N_2957,N_2966);
and UO_416 (O_416,N_2958,N_2961);
or UO_417 (O_417,N_2961,N_2943);
xor UO_418 (O_418,N_2987,N_2991);
nand UO_419 (O_419,N_2986,N_2974);
xnor UO_420 (O_420,N_2995,N_2968);
xor UO_421 (O_421,N_2993,N_2944);
and UO_422 (O_422,N_2954,N_2966);
or UO_423 (O_423,N_2951,N_2976);
xor UO_424 (O_424,N_2997,N_2941);
nand UO_425 (O_425,N_2952,N_2972);
and UO_426 (O_426,N_2965,N_2967);
or UO_427 (O_427,N_2975,N_2941);
xnor UO_428 (O_428,N_2993,N_2977);
and UO_429 (O_429,N_2972,N_2945);
or UO_430 (O_430,N_2958,N_2998);
nand UO_431 (O_431,N_2966,N_2979);
xnor UO_432 (O_432,N_2947,N_2950);
nand UO_433 (O_433,N_2991,N_2966);
nand UO_434 (O_434,N_2968,N_2956);
nand UO_435 (O_435,N_2983,N_2961);
nand UO_436 (O_436,N_2960,N_2975);
and UO_437 (O_437,N_2997,N_2948);
and UO_438 (O_438,N_2957,N_2990);
nand UO_439 (O_439,N_2970,N_2968);
or UO_440 (O_440,N_2970,N_2944);
and UO_441 (O_441,N_2971,N_2958);
xor UO_442 (O_442,N_2981,N_2956);
xor UO_443 (O_443,N_2967,N_2982);
and UO_444 (O_444,N_2994,N_2974);
or UO_445 (O_445,N_2994,N_2940);
xor UO_446 (O_446,N_2943,N_2953);
xnor UO_447 (O_447,N_2950,N_2977);
xor UO_448 (O_448,N_2997,N_2998);
and UO_449 (O_449,N_2978,N_2943);
xnor UO_450 (O_450,N_2976,N_2992);
xnor UO_451 (O_451,N_2963,N_2983);
or UO_452 (O_452,N_2957,N_2995);
xor UO_453 (O_453,N_2963,N_2990);
nand UO_454 (O_454,N_2995,N_2949);
and UO_455 (O_455,N_2956,N_2996);
xnor UO_456 (O_456,N_2949,N_2961);
or UO_457 (O_457,N_2974,N_2957);
xnor UO_458 (O_458,N_2973,N_2962);
xor UO_459 (O_459,N_2964,N_2994);
or UO_460 (O_460,N_2946,N_2984);
or UO_461 (O_461,N_2992,N_2994);
nand UO_462 (O_462,N_2991,N_2945);
nor UO_463 (O_463,N_2987,N_2984);
nor UO_464 (O_464,N_2992,N_2952);
nor UO_465 (O_465,N_2941,N_2966);
nor UO_466 (O_466,N_2970,N_2958);
nand UO_467 (O_467,N_2987,N_2940);
nor UO_468 (O_468,N_2976,N_2994);
and UO_469 (O_469,N_2973,N_2991);
and UO_470 (O_470,N_2954,N_2960);
nand UO_471 (O_471,N_2976,N_2968);
and UO_472 (O_472,N_2975,N_2993);
and UO_473 (O_473,N_2978,N_2989);
nor UO_474 (O_474,N_2991,N_2961);
nor UO_475 (O_475,N_2982,N_2966);
and UO_476 (O_476,N_2968,N_2965);
xor UO_477 (O_477,N_2982,N_2993);
or UO_478 (O_478,N_2975,N_2985);
nand UO_479 (O_479,N_2957,N_2967);
xnor UO_480 (O_480,N_2972,N_2998);
xnor UO_481 (O_481,N_2961,N_2946);
nor UO_482 (O_482,N_2997,N_2970);
or UO_483 (O_483,N_2966,N_2968);
nand UO_484 (O_484,N_2947,N_2958);
nand UO_485 (O_485,N_2961,N_2988);
nor UO_486 (O_486,N_2972,N_2991);
or UO_487 (O_487,N_2964,N_2946);
and UO_488 (O_488,N_2956,N_2965);
nor UO_489 (O_489,N_2964,N_2953);
nor UO_490 (O_490,N_2960,N_2952);
xnor UO_491 (O_491,N_2961,N_2994);
xor UO_492 (O_492,N_2963,N_2975);
and UO_493 (O_493,N_2969,N_2947);
and UO_494 (O_494,N_2992,N_2986);
or UO_495 (O_495,N_2974,N_2949);
nor UO_496 (O_496,N_2945,N_2998);
xor UO_497 (O_497,N_2963,N_2995);
nor UO_498 (O_498,N_2943,N_2948);
xor UO_499 (O_499,N_2998,N_2961);
endmodule