module basic_1000_10000_1500_5_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_0,In_267);
or U1 (N_1,In_994,In_335);
nand U2 (N_2,In_913,In_266);
nor U3 (N_3,In_864,In_923);
or U4 (N_4,In_808,In_964);
and U5 (N_5,In_793,In_287);
nor U6 (N_6,In_324,In_201);
nor U7 (N_7,In_722,In_355);
and U8 (N_8,In_34,In_907);
nand U9 (N_9,In_40,In_55);
nand U10 (N_10,In_498,In_777);
and U11 (N_11,In_1,In_929);
or U12 (N_12,In_865,In_566);
nor U13 (N_13,In_223,In_998);
or U14 (N_14,In_354,In_131);
nand U15 (N_15,In_203,In_749);
and U16 (N_16,In_129,In_323);
nor U17 (N_17,In_825,In_692);
nand U18 (N_18,In_547,In_155);
or U19 (N_19,In_684,In_352);
or U20 (N_20,In_384,In_948);
xnor U21 (N_21,In_270,In_814);
or U22 (N_22,In_123,In_659);
and U23 (N_23,In_960,In_197);
nor U24 (N_24,In_532,In_363);
or U25 (N_25,In_405,In_748);
and U26 (N_26,In_370,In_971);
and U27 (N_27,In_503,In_318);
or U28 (N_28,In_506,In_185);
or U29 (N_29,In_407,In_641);
and U30 (N_30,In_141,In_778);
or U31 (N_31,In_169,In_963);
nand U32 (N_32,In_480,In_952);
nand U33 (N_33,In_11,In_481);
or U34 (N_34,In_837,In_773);
or U35 (N_35,In_242,In_983);
nand U36 (N_36,In_877,In_950);
and U37 (N_37,In_918,In_982);
and U38 (N_38,In_632,In_424);
nand U39 (N_39,In_365,In_48);
nor U40 (N_40,In_130,In_309);
nand U41 (N_41,In_658,In_465);
nor U42 (N_42,In_797,In_235);
or U43 (N_43,In_263,In_174);
or U44 (N_44,In_920,In_179);
or U45 (N_45,In_184,In_711);
or U46 (N_46,In_327,In_935);
or U47 (N_47,In_359,In_910);
nand U48 (N_48,In_151,In_701);
xnor U49 (N_49,In_124,In_905);
nor U50 (N_50,In_953,In_975);
or U51 (N_51,In_829,In_22);
or U52 (N_52,In_602,In_727);
nor U53 (N_53,In_332,In_482);
nor U54 (N_54,In_436,In_210);
and U55 (N_55,In_887,In_746);
nand U56 (N_56,In_931,In_614);
nor U57 (N_57,In_928,In_820);
nor U58 (N_58,In_858,In_13);
nand U59 (N_59,In_233,In_400);
and U60 (N_60,In_981,In_799);
nor U61 (N_61,In_431,In_536);
nand U62 (N_62,In_285,In_574);
and U63 (N_63,In_810,In_468);
nor U64 (N_64,In_144,In_888);
xor U65 (N_65,In_795,In_484);
nand U66 (N_66,In_968,In_885);
and U67 (N_67,In_588,In_551);
nor U68 (N_68,In_107,In_417);
nor U69 (N_69,In_709,In_71);
nand U70 (N_70,In_30,In_261);
or U71 (N_71,In_416,In_522);
nand U72 (N_72,In_554,In_898);
nand U73 (N_73,In_337,In_163);
nand U74 (N_74,In_544,In_739);
or U75 (N_75,In_956,In_694);
nor U76 (N_76,In_310,In_500);
nand U77 (N_77,In_138,In_903);
and U78 (N_78,In_446,In_98);
or U79 (N_79,In_967,In_507);
or U80 (N_80,In_700,In_183);
or U81 (N_81,In_895,In_325);
nand U82 (N_82,In_136,In_474);
nand U83 (N_83,In_863,In_651);
nor U84 (N_84,In_200,In_630);
or U85 (N_85,In_281,In_220);
or U86 (N_86,In_853,In_404);
or U87 (N_87,In_996,In_788);
nand U88 (N_88,In_565,In_284);
nor U89 (N_89,In_445,In_294);
nor U90 (N_90,In_550,In_985);
nand U91 (N_91,In_139,In_234);
or U92 (N_92,In_957,In_342);
nand U93 (N_93,In_82,In_378);
and U94 (N_94,In_784,In_635);
or U95 (N_95,In_954,In_598);
or U96 (N_96,In_891,In_254);
or U97 (N_97,In_487,In_610);
nor U98 (N_98,In_977,In_856);
or U99 (N_99,In_356,In_27);
nor U100 (N_100,In_580,In_763);
nand U101 (N_101,In_36,In_575);
nor U102 (N_102,In_271,In_361);
xor U103 (N_103,In_24,In_938);
and U104 (N_104,In_851,In_840);
nand U105 (N_105,In_54,In_67);
and U106 (N_106,In_389,In_186);
nand U107 (N_107,In_501,In_742);
nor U108 (N_108,In_539,In_785);
and U109 (N_109,In_428,In_674);
or U110 (N_110,In_666,In_120);
nor U111 (N_111,In_198,In_529);
or U112 (N_112,In_690,In_707);
or U113 (N_113,In_549,In_677);
or U114 (N_114,In_644,In_958);
nor U115 (N_115,In_463,In_319);
xor U116 (N_116,In_754,In_766);
xnor U117 (N_117,In_473,In_329);
xnor U118 (N_118,In_505,In_341);
and U119 (N_119,In_542,In_304);
or U120 (N_120,In_798,In_984);
and U121 (N_121,In_495,In_401);
and U122 (N_122,In_317,In_687);
or U123 (N_123,In_857,In_939);
and U124 (N_124,In_872,In_768);
nand U125 (N_125,In_879,In_555);
nand U126 (N_126,In_257,In_801);
or U127 (N_127,In_670,In_892);
or U128 (N_128,In_31,In_615);
or U129 (N_129,In_483,In_278);
and U130 (N_130,In_455,In_292);
and U131 (N_131,In_53,In_275);
and U132 (N_132,In_740,In_158);
or U133 (N_133,In_274,In_188);
or U134 (N_134,In_770,In_75);
or U135 (N_135,In_812,In_936);
nor U136 (N_136,In_52,In_32);
or U137 (N_137,In_245,In_221);
or U138 (N_138,In_37,In_940);
nand U139 (N_139,In_18,In_86);
and U140 (N_140,In_252,In_328);
xnor U141 (N_141,In_458,In_77);
nand U142 (N_142,In_695,In_624);
and U143 (N_143,In_564,In_375);
nand U144 (N_144,In_121,In_525);
and U145 (N_145,In_597,In_927);
nand U146 (N_146,In_85,In_15);
nor U147 (N_147,In_909,In_38);
nor U148 (N_148,In_461,In_642);
or U149 (N_149,In_349,In_921);
xor U150 (N_150,In_741,In_567);
nand U151 (N_151,In_213,In_623);
xor U152 (N_152,In_225,In_914);
and U153 (N_153,In_492,In_576);
nor U154 (N_154,In_866,In_586);
xnor U155 (N_155,In_875,In_358);
nand U156 (N_156,In_496,In_16);
nor U157 (N_157,In_966,In_678);
xor U158 (N_158,In_861,In_391);
nand U159 (N_159,In_710,In_942);
and U160 (N_160,In_886,In_448);
xnor U161 (N_161,In_511,In_326);
xor U162 (N_162,In_764,In_970);
or U163 (N_163,In_673,In_787);
or U164 (N_164,In_870,In_871);
xnor U165 (N_165,In_421,In_330);
nor U166 (N_166,In_541,In_519);
nor U167 (N_167,In_753,In_896);
or U168 (N_168,In_125,In_313);
nand U169 (N_169,In_691,In_504);
xnor U170 (N_170,In_732,In_59);
and U171 (N_171,In_862,In_944);
nand U172 (N_172,In_20,In_637);
and U173 (N_173,In_170,In_699);
or U174 (N_174,In_582,In_973);
or U175 (N_175,In_530,In_58);
nand U176 (N_176,In_403,In_789);
nand U177 (N_177,In_729,In_548);
or U178 (N_178,In_388,In_934);
nand U179 (N_179,In_260,In_546);
nor U180 (N_180,In_250,In_301);
nand U181 (N_181,In_643,In_608);
nand U182 (N_182,In_29,In_884);
nand U183 (N_183,In_290,In_959);
nand U184 (N_184,In_676,In_828);
or U185 (N_185,In_414,In_173);
and U186 (N_186,In_802,In_847);
nand U187 (N_187,In_600,In_704);
nand U188 (N_188,In_122,In_925);
and U189 (N_189,In_272,In_51);
or U190 (N_190,In_491,In_241);
xor U191 (N_191,In_584,In_372);
nor U192 (N_192,In_962,In_843);
and U193 (N_193,In_663,In_119);
nand U194 (N_194,In_955,In_227);
xnor U195 (N_195,In_974,In_104);
or U196 (N_196,In_73,In_626);
and U197 (N_197,In_848,In_535);
or U198 (N_198,In_559,In_418);
nand U199 (N_199,In_890,In_762);
nor U200 (N_200,In_779,In_50);
xor U201 (N_201,In_145,In_737);
nor U202 (N_202,In_110,In_805);
or U203 (N_203,In_114,In_490);
or U204 (N_204,In_256,In_279);
xnor U205 (N_205,In_723,In_478);
and U206 (N_206,In_297,In_65);
nand U207 (N_207,In_395,In_288);
and U208 (N_208,In_81,In_719);
nor U209 (N_209,In_399,In_322);
or U210 (N_210,In_207,In_581);
xnor U211 (N_211,In_744,In_154);
or U212 (N_212,In_61,In_930);
or U213 (N_213,In_613,In_108);
nor U214 (N_214,In_611,In_599);
nor U215 (N_215,In_331,In_190);
or U216 (N_216,In_650,In_538);
and U217 (N_217,In_572,In_760);
nand U218 (N_218,In_56,In_187);
or U219 (N_219,In_721,In_751);
nand U220 (N_220,In_655,In_606);
nand U221 (N_221,In_873,In_238);
and U222 (N_222,In_628,In_49);
and U223 (N_223,In_860,In_889);
nor U224 (N_224,In_380,In_752);
nand U225 (N_225,In_444,In_406);
nor U226 (N_226,In_743,In_621);
nand U227 (N_227,In_915,In_912);
nand U228 (N_228,In_993,In_579);
and U229 (N_229,In_874,In_443);
or U230 (N_230,In_282,In_681);
or U231 (N_231,In_855,In_259);
and U232 (N_232,In_652,In_502);
xor U233 (N_233,In_293,In_657);
nor U234 (N_234,In_410,In_181);
and U235 (N_235,In_685,In_800);
nor U236 (N_236,In_593,In_987);
nand U237 (N_237,In_427,In_215);
nor U238 (N_238,In_452,In_537);
or U239 (N_239,In_577,In_647);
and U240 (N_240,In_570,In_782);
or U241 (N_241,In_922,In_826);
or U242 (N_242,In_883,In_774);
nand U243 (N_243,In_617,In_348);
nor U244 (N_244,In_305,In_553);
or U245 (N_245,In_373,In_786);
nor U246 (N_246,In_587,In_645);
or U247 (N_247,In_791,In_96);
and U248 (N_248,In_589,In_750);
or U249 (N_249,In_19,In_196);
and U250 (N_250,In_453,In_845);
nand U251 (N_251,In_720,In_790);
xnor U252 (N_252,In_594,In_730);
nor U253 (N_253,In_265,In_671);
nor U254 (N_254,In_216,In_368);
nor U255 (N_255,In_454,In_69);
nand U256 (N_256,In_633,In_94);
nand U257 (N_257,In_457,In_253);
nand U258 (N_258,In_543,In_426);
nor U259 (N_259,In_276,In_804);
nor U260 (N_260,In_303,In_346);
or U261 (N_261,In_150,In_489);
and U262 (N_262,In_239,In_702);
or U263 (N_263,In_683,In_409);
and U264 (N_264,In_941,In_316);
nor U265 (N_265,In_965,In_47);
or U266 (N_266,In_943,In_514);
nor U267 (N_267,In_419,In_88);
and U268 (N_268,In_631,In_9);
or U269 (N_269,In_714,In_618);
or U270 (N_270,In_258,In_464);
xor U271 (N_271,In_60,In_78);
nor U272 (N_272,In_758,In_485);
nor U273 (N_273,In_733,In_39);
nand U274 (N_274,In_343,In_35);
and U275 (N_275,In_470,In_376);
xnor U276 (N_276,In_634,In_609);
nand U277 (N_277,In_182,In_243);
xnor U278 (N_278,In_134,In_757);
nor U279 (N_279,In_604,In_79);
nor U280 (N_280,In_781,In_653);
nand U281 (N_281,In_299,In_148);
nor U282 (N_282,In_622,In_402);
nand U283 (N_283,In_980,In_693);
and U284 (N_284,In_441,In_63);
or U285 (N_285,In_244,In_423);
nor U286 (N_286,In_988,In_979);
and U287 (N_287,In_161,In_806);
xnor U288 (N_288,In_472,In_780);
and U289 (N_289,In_57,In_509);
or U290 (N_290,In_515,In_989);
nor U291 (N_291,In_240,In_229);
nor U292 (N_292,In_715,In_153);
nand U293 (N_293,In_901,In_300);
or U294 (N_294,In_708,In_841);
or U295 (N_295,In_412,In_911);
nand U296 (N_296,In_42,In_717);
nand U297 (N_297,In_456,In_705);
xor U298 (N_298,In_99,In_377);
nand U299 (N_299,In_237,In_510);
nand U300 (N_300,In_25,In_745);
nand U301 (N_301,In_118,In_601);
nand U302 (N_302,In_269,In_759);
nor U303 (N_303,In_435,In_596);
nand U304 (N_304,In_512,In_919);
or U305 (N_305,In_199,In_236);
or U306 (N_306,In_852,In_859);
xnor U307 (N_307,In_545,In_135);
and U308 (N_308,In_398,In_7);
nor U309 (N_309,In_209,In_675);
nand U310 (N_310,In_809,In_291);
nor U311 (N_311,In_698,In_14);
and U312 (N_312,In_947,In_442);
or U313 (N_313,In_202,In_807);
or U314 (N_314,In_756,In_152);
or U315 (N_315,In_924,In_682);
nand U316 (N_316,In_568,In_383);
or U317 (N_317,In_603,In_823);
or U318 (N_318,In_854,In_619);
nor U319 (N_319,In_513,In_353);
or U320 (N_320,In_595,In_616);
nand U321 (N_321,In_390,In_280);
nor U322 (N_322,In_206,In_140);
and U323 (N_323,In_493,In_508);
nand U324 (N_324,In_45,In_433);
and U325 (N_325,In_83,In_128);
nand U326 (N_326,In_661,In_916);
and U327 (N_327,In_712,In_881);
or U328 (N_328,In_44,In_667);
nand U329 (N_329,In_822,In_17);
nor U330 (N_330,In_264,In_164);
nor U331 (N_331,In_605,In_249);
nand U332 (N_332,In_33,In_697);
or U333 (N_333,In_385,In_102);
nand U334 (N_334,In_106,In_524);
nand U335 (N_335,In_109,In_990);
and U336 (N_336,In_408,In_262);
nor U337 (N_337,In_434,In_897);
xor U338 (N_338,In_429,In_629);
nand U339 (N_339,In_439,In_724);
nor U340 (N_340,In_307,In_248);
xnor U341 (N_341,In_146,In_451);
nand U342 (N_342,In_10,In_339);
or U343 (N_343,In_450,In_344);
nand U344 (N_344,In_80,In_563);
and U345 (N_345,In_394,In_23);
nor U346 (N_346,In_747,In_469);
or U347 (N_347,In_101,In_413);
or U348 (N_348,In_133,In_231);
and U349 (N_349,In_571,In_298);
nand U350 (N_350,In_999,In_171);
nor U351 (N_351,In_127,In_76);
or U352 (N_352,In_771,In_842);
nand U353 (N_353,In_351,In_821);
xor U354 (N_354,In_516,In_46);
xor U355 (N_355,In_783,In_718);
nand U356 (N_356,In_374,In_371);
nor U357 (N_357,In_725,In_112);
xor U358 (N_358,In_816,In_558);
or U359 (N_359,In_247,In_165);
nand U360 (N_360,In_302,In_835);
or U361 (N_361,In_569,In_180);
nor U362 (N_362,In_66,In_649);
nand U363 (N_363,In_672,In_459);
nor U364 (N_364,In_4,In_159);
or U365 (N_365,In_393,In_103);
or U366 (N_366,In_41,In_591);
or U367 (N_367,In_396,In_893);
nand U368 (N_368,In_899,In_876);
or U369 (N_369,In_156,In_97);
and U370 (N_370,In_345,In_562);
nor U371 (N_371,In_904,In_830);
nand U372 (N_372,In_100,In_268);
nor U373 (N_373,In_43,In_607);
and U374 (N_374,In_437,In_583);
or U375 (N_375,In_177,In_357);
and U376 (N_376,In_908,In_976);
or U377 (N_377,In_665,In_868);
or U378 (N_378,In_639,In_204);
xnor U379 (N_379,In_533,In_517);
xor U380 (N_380,In_132,In_648);
or U381 (N_381,In_84,In_308);
nor U382 (N_382,In_526,In_590);
nand U383 (N_383,In_26,In_475);
and U384 (N_384,In_230,In_178);
or U385 (N_385,In_573,In_289);
nor U386 (N_386,In_882,In_447);
or U387 (N_387,In_668,In_420);
nor U388 (N_388,In_350,In_926);
nand U389 (N_389,In_314,In_226);
nand U390 (N_390,In_321,In_422);
xor U391 (N_391,In_552,In_246);
and U392 (N_392,In_834,In_728);
nor U393 (N_393,In_74,In_126);
nor U394 (N_394,In_713,In_726);
and U395 (N_395,In_21,In_906);
or U396 (N_396,In_578,In_969);
or U397 (N_397,In_194,In_286);
or U398 (N_398,In_902,In_311);
or U399 (N_399,In_765,In_933);
or U400 (N_400,In_776,In_386);
nor U401 (N_401,In_193,In_162);
nand U402 (N_402,In_646,In_731);
nor U403 (N_403,In_315,In_775);
or U404 (N_404,In_736,In_937);
and U405 (N_405,In_105,In_794);
nor U406 (N_406,In_831,In_340);
or U407 (N_407,In_612,In_460);
and U408 (N_408,In_392,In_827);
or U409 (N_409,In_360,In_523);
nand U410 (N_410,In_338,In_277);
xor U411 (N_411,In_143,In_900);
nand U412 (N_412,In_620,In_160);
and U413 (N_413,In_440,In_767);
xnor U414 (N_414,In_415,In_222);
nor U415 (N_415,In_6,In_662);
nor U416 (N_416,In_12,In_479);
nand U417 (N_417,In_208,In_149);
or U418 (N_418,In_664,In_62);
and U419 (N_419,In_425,In_991);
and U420 (N_420,In_494,In_90);
nand U421 (N_421,In_362,In_471);
nor U422 (N_422,In_364,In_585);
and U423 (N_423,In_336,In_157);
or U424 (N_424,In_846,In_817);
nor U425 (N_425,In_467,In_867);
or U426 (N_426,In_894,In_844);
nand U427 (N_427,In_366,In_534);
or U428 (N_428,In_518,In_992);
nand U429 (N_429,In_686,In_849);
nor U430 (N_430,In_560,In_836);
or U431 (N_431,In_951,In_195);
and U432 (N_432,In_486,In_669);
nand U433 (N_433,In_219,In_217);
nand U434 (N_434,In_528,In_166);
nand U435 (N_435,In_679,In_755);
nand U436 (N_436,In_312,In_932);
nand U437 (N_437,In_769,In_772);
nor U438 (N_438,In_716,In_869);
and U439 (N_439,In_995,In_462);
xor U440 (N_440,In_382,In_228);
or U441 (N_441,In_172,In_557);
and U442 (N_442,In_488,In_438);
nand U443 (N_443,In_689,In_476);
or U444 (N_444,In_115,In_232);
nor U445 (N_445,In_411,In_499);
xnor U446 (N_446,In_636,In_218);
nor U447 (N_447,In_379,In_833);
nand U448 (N_448,In_625,In_703);
and U449 (N_449,In_95,In_273);
and U450 (N_450,In_986,In_997);
xnor U451 (N_451,In_815,In_68);
nor U452 (N_452,In_497,In_397);
nand U453 (N_453,In_283,In_792);
nor U454 (N_454,In_214,In_654);
and U455 (N_455,In_432,In_93);
or U456 (N_456,In_333,In_92);
and U457 (N_457,In_761,In_295);
nor U458 (N_458,In_211,In_521);
or U459 (N_459,In_819,In_192);
and U460 (N_460,In_175,In_878);
nor U461 (N_461,In_660,In_527);
and U462 (N_462,In_320,In_255);
nor U463 (N_463,In_592,In_347);
nand U464 (N_464,In_638,In_191);
nand U465 (N_465,In_189,In_70);
and U466 (N_466,In_961,In_738);
and U467 (N_467,In_477,In_466);
and U468 (N_468,In_2,In_89);
or U469 (N_469,In_838,In_449);
and U470 (N_470,In_387,In_978);
nor U471 (N_471,In_680,In_176);
nor U472 (N_472,In_832,In_706);
nor U473 (N_473,In_205,In_531);
nand U474 (N_474,In_796,In_824);
and U475 (N_475,In_3,In_556);
or U476 (N_476,In_87,In_111);
or U477 (N_477,In_627,In_839);
or U478 (N_478,In_520,In_367);
nand U479 (N_479,In_251,In_880);
and U480 (N_480,In_640,In_167);
nor U481 (N_481,In_735,In_696);
or U482 (N_482,In_381,In_91);
and U483 (N_483,In_917,In_561);
nor U484 (N_484,In_212,In_224);
nand U485 (N_485,In_137,In_656);
xor U486 (N_486,In_813,In_147);
nand U487 (N_487,In_946,In_5);
xor U488 (N_488,In_850,In_734);
and U489 (N_489,In_306,In_540);
and U490 (N_490,In_430,In_688);
and U491 (N_491,In_116,In_8);
nor U492 (N_492,In_296,In_945);
nand U493 (N_493,In_142,In_972);
or U494 (N_494,In_64,In_811);
xnor U495 (N_495,In_949,In_369);
nor U496 (N_496,In_818,In_113);
and U497 (N_497,In_72,In_117);
nand U498 (N_498,In_334,In_168);
or U499 (N_499,In_803,In_28);
nand U500 (N_500,In_568,In_275);
and U501 (N_501,In_683,In_6);
and U502 (N_502,In_766,In_615);
nand U503 (N_503,In_82,In_601);
nand U504 (N_504,In_608,In_310);
or U505 (N_505,In_357,In_205);
xnor U506 (N_506,In_653,In_60);
and U507 (N_507,In_102,In_623);
xnor U508 (N_508,In_911,In_980);
nand U509 (N_509,In_238,In_882);
or U510 (N_510,In_387,In_603);
or U511 (N_511,In_137,In_842);
nor U512 (N_512,In_729,In_931);
xnor U513 (N_513,In_168,In_227);
and U514 (N_514,In_428,In_41);
nand U515 (N_515,In_727,In_252);
nor U516 (N_516,In_330,In_238);
xnor U517 (N_517,In_397,In_780);
nor U518 (N_518,In_416,In_348);
nor U519 (N_519,In_857,In_874);
or U520 (N_520,In_718,In_604);
or U521 (N_521,In_354,In_589);
and U522 (N_522,In_632,In_725);
and U523 (N_523,In_381,In_651);
or U524 (N_524,In_970,In_621);
or U525 (N_525,In_94,In_410);
or U526 (N_526,In_782,In_755);
or U527 (N_527,In_66,In_864);
and U528 (N_528,In_467,In_122);
nor U529 (N_529,In_290,In_730);
nor U530 (N_530,In_496,In_646);
and U531 (N_531,In_425,In_760);
xor U532 (N_532,In_743,In_185);
xnor U533 (N_533,In_980,In_416);
and U534 (N_534,In_712,In_977);
and U535 (N_535,In_933,In_902);
or U536 (N_536,In_770,In_601);
or U537 (N_537,In_65,In_828);
and U538 (N_538,In_434,In_386);
and U539 (N_539,In_272,In_9);
nor U540 (N_540,In_166,In_45);
nor U541 (N_541,In_796,In_117);
and U542 (N_542,In_496,In_761);
nor U543 (N_543,In_448,In_902);
and U544 (N_544,In_279,In_641);
and U545 (N_545,In_211,In_544);
and U546 (N_546,In_244,In_167);
or U547 (N_547,In_851,In_505);
nor U548 (N_548,In_271,In_537);
or U549 (N_549,In_159,In_407);
nor U550 (N_550,In_697,In_57);
nor U551 (N_551,In_33,In_184);
nand U552 (N_552,In_377,In_71);
or U553 (N_553,In_96,In_418);
and U554 (N_554,In_638,In_802);
nor U555 (N_555,In_301,In_425);
xnor U556 (N_556,In_415,In_544);
and U557 (N_557,In_282,In_801);
or U558 (N_558,In_404,In_896);
nand U559 (N_559,In_651,In_173);
nor U560 (N_560,In_571,In_618);
or U561 (N_561,In_576,In_490);
nor U562 (N_562,In_429,In_670);
or U563 (N_563,In_595,In_291);
nor U564 (N_564,In_558,In_459);
nand U565 (N_565,In_192,In_655);
or U566 (N_566,In_232,In_996);
or U567 (N_567,In_132,In_967);
nand U568 (N_568,In_657,In_772);
nor U569 (N_569,In_384,In_988);
xor U570 (N_570,In_131,In_308);
nand U571 (N_571,In_660,In_140);
and U572 (N_572,In_704,In_362);
nand U573 (N_573,In_981,In_94);
or U574 (N_574,In_859,In_152);
and U575 (N_575,In_98,In_813);
nor U576 (N_576,In_556,In_481);
xor U577 (N_577,In_608,In_728);
or U578 (N_578,In_969,In_385);
xnor U579 (N_579,In_798,In_932);
or U580 (N_580,In_724,In_740);
nor U581 (N_581,In_16,In_563);
and U582 (N_582,In_893,In_614);
and U583 (N_583,In_183,In_930);
nand U584 (N_584,In_738,In_474);
nand U585 (N_585,In_678,In_683);
nand U586 (N_586,In_343,In_692);
xnor U587 (N_587,In_586,In_999);
nand U588 (N_588,In_395,In_279);
nor U589 (N_589,In_622,In_701);
xnor U590 (N_590,In_663,In_550);
or U591 (N_591,In_139,In_199);
or U592 (N_592,In_832,In_335);
or U593 (N_593,In_935,In_855);
nand U594 (N_594,In_515,In_679);
and U595 (N_595,In_272,In_750);
and U596 (N_596,In_857,In_126);
or U597 (N_597,In_743,In_930);
nor U598 (N_598,In_76,In_633);
or U599 (N_599,In_836,In_20);
nand U600 (N_600,In_775,In_181);
and U601 (N_601,In_360,In_269);
or U602 (N_602,In_368,In_438);
nand U603 (N_603,In_755,In_304);
nor U604 (N_604,In_128,In_801);
nor U605 (N_605,In_773,In_233);
nor U606 (N_606,In_336,In_196);
nor U607 (N_607,In_858,In_845);
and U608 (N_608,In_300,In_342);
and U609 (N_609,In_797,In_607);
nor U610 (N_610,In_490,In_292);
and U611 (N_611,In_442,In_830);
and U612 (N_612,In_699,In_575);
nor U613 (N_613,In_196,In_547);
nand U614 (N_614,In_433,In_742);
and U615 (N_615,In_841,In_637);
nand U616 (N_616,In_73,In_274);
or U617 (N_617,In_623,In_702);
nor U618 (N_618,In_887,In_556);
and U619 (N_619,In_101,In_12);
nor U620 (N_620,In_654,In_325);
and U621 (N_621,In_839,In_838);
or U622 (N_622,In_619,In_447);
nand U623 (N_623,In_626,In_325);
nor U624 (N_624,In_771,In_652);
or U625 (N_625,In_235,In_743);
or U626 (N_626,In_108,In_275);
nor U627 (N_627,In_257,In_344);
nor U628 (N_628,In_824,In_612);
nand U629 (N_629,In_80,In_582);
and U630 (N_630,In_595,In_974);
xnor U631 (N_631,In_259,In_647);
and U632 (N_632,In_903,In_652);
xnor U633 (N_633,In_330,In_340);
and U634 (N_634,In_383,In_734);
nor U635 (N_635,In_874,In_826);
xnor U636 (N_636,In_985,In_94);
nor U637 (N_637,In_302,In_195);
nor U638 (N_638,In_190,In_929);
and U639 (N_639,In_500,In_750);
nor U640 (N_640,In_419,In_80);
or U641 (N_641,In_682,In_417);
and U642 (N_642,In_506,In_64);
xor U643 (N_643,In_596,In_905);
and U644 (N_644,In_215,In_925);
nand U645 (N_645,In_921,In_175);
or U646 (N_646,In_738,In_475);
nand U647 (N_647,In_712,In_482);
or U648 (N_648,In_838,In_405);
or U649 (N_649,In_593,In_678);
and U650 (N_650,In_885,In_267);
nor U651 (N_651,In_601,In_405);
and U652 (N_652,In_994,In_617);
and U653 (N_653,In_125,In_440);
or U654 (N_654,In_196,In_442);
nand U655 (N_655,In_899,In_15);
nand U656 (N_656,In_534,In_98);
and U657 (N_657,In_975,In_391);
nor U658 (N_658,In_264,In_528);
nor U659 (N_659,In_870,In_29);
xor U660 (N_660,In_37,In_424);
nor U661 (N_661,In_91,In_476);
or U662 (N_662,In_283,In_795);
nor U663 (N_663,In_928,In_285);
xor U664 (N_664,In_60,In_111);
nor U665 (N_665,In_792,In_286);
or U666 (N_666,In_777,In_842);
and U667 (N_667,In_776,In_468);
and U668 (N_668,In_283,In_308);
or U669 (N_669,In_436,In_207);
nand U670 (N_670,In_567,In_375);
nand U671 (N_671,In_599,In_580);
xor U672 (N_672,In_671,In_667);
nand U673 (N_673,In_248,In_810);
and U674 (N_674,In_395,In_232);
and U675 (N_675,In_927,In_720);
or U676 (N_676,In_509,In_881);
and U677 (N_677,In_237,In_155);
or U678 (N_678,In_566,In_240);
and U679 (N_679,In_967,In_317);
or U680 (N_680,In_410,In_424);
or U681 (N_681,In_339,In_964);
nor U682 (N_682,In_319,In_618);
nor U683 (N_683,In_592,In_969);
nor U684 (N_684,In_447,In_131);
nand U685 (N_685,In_393,In_241);
nor U686 (N_686,In_974,In_924);
nor U687 (N_687,In_433,In_394);
nor U688 (N_688,In_500,In_521);
xor U689 (N_689,In_846,In_453);
and U690 (N_690,In_414,In_812);
or U691 (N_691,In_161,In_750);
or U692 (N_692,In_241,In_687);
xnor U693 (N_693,In_115,In_990);
or U694 (N_694,In_310,In_793);
or U695 (N_695,In_416,In_765);
nor U696 (N_696,In_454,In_672);
or U697 (N_697,In_473,In_271);
nand U698 (N_698,In_226,In_175);
or U699 (N_699,In_125,In_941);
xor U700 (N_700,In_233,In_198);
and U701 (N_701,In_135,In_394);
xor U702 (N_702,In_589,In_831);
or U703 (N_703,In_822,In_294);
and U704 (N_704,In_952,In_293);
xor U705 (N_705,In_573,In_807);
and U706 (N_706,In_316,In_893);
nor U707 (N_707,In_830,In_323);
or U708 (N_708,In_330,In_580);
nand U709 (N_709,In_353,In_10);
nor U710 (N_710,In_765,In_54);
and U711 (N_711,In_367,In_961);
or U712 (N_712,In_792,In_813);
nor U713 (N_713,In_341,In_0);
nor U714 (N_714,In_181,In_431);
and U715 (N_715,In_718,In_49);
nor U716 (N_716,In_628,In_955);
and U717 (N_717,In_380,In_624);
and U718 (N_718,In_110,In_341);
nand U719 (N_719,In_851,In_783);
or U720 (N_720,In_694,In_308);
and U721 (N_721,In_758,In_674);
or U722 (N_722,In_769,In_29);
and U723 (N_723,In_495,In_388);
xor U724 (N_724,In_992,In_142);
nor U725 (N_725,In_498,In_946);
xnor U726 (N_726,In_981,In_849);
nor U727 (N_727,In_451,In_788);
or U728 (N_728,In_228,In_27);
and U729 (N_729,In_47,In_428);
nor U730 (N_730,In_834,In_367);
and U731 (N_731,In_467,In_747);
and U732 (N_732,In_64,In_949);
and U733 (N_733,In_445,In_896);
xnor U734 (N_734,In_828,In_985);
xor U735 (N_735,In_952,In_700);
nand U736 (N_736,In_795,In_263);
nand U737 (N_737,In_573,In_124);
nand U738 (N_738,In_912,In_204);
or U739 (N_739,In_434,In_83);
nand U740 (N_740,In_888,In_555);
nor U741 (N_741,In_226,In_830);
nand U742 (N_742,In_379,In_607);
nor U743 (N_743,In_530,In_293);
nand U744 (N_744,In_689,In_797);
nor U745 (N_745,In_658,In_998);
and U746 (N_746,In_64,In_992);
and U747 (N_747,In_308,In_997);
xor U748 (N_748,In_397,In_498);
or U749 (N_749,In_345,In_132);
and U750 (N_750,In_479,In_153);
nand U751 (N_751,In_746,In_812);
and U752 (N_752,In_131,In_414);
or U753 (N_753,In_764,In_426);
or U754 (N_754,In_26,In_565);
and U755 (N_755,In_52,In_219);
nor U756 (N_756,In_162,In_868);
xnor U757 (N_757,In_778,In_286);
and U758 (N_758,In_262,In_137);
nor U759 (N_759,In_61,In_890);
nand U760 (N_760,In_21,In_755);
and U761 (N_761,In_620,In_694);
and U762 (N_762,In_108,In_583);
nand U763 (N_763,In_791,In_135);
nor U764 (N_764,In_709,In_341);
or U765 (N_765,In_220,In_491);
nand U766 (N_766,In_71,In_181);
nor U767 (N_767,In_839,In_334);
and U768 (N_768,In_547,In_734);
nor U769 (N_769,In_260,In_490);
nor U770 (N_770,In_820,In_977);
nor U771 (N_771,In_183,In_927);
and U772 (N_772,In_770,In_533);
or U773 (N_773,In_532,In_144);
and U774 (N_774,In_944,In_687);
nand U775 (N_775,In_825,In_424);
nand U776 (N_776,In_609,In_258);
xnor U777 (N_777,In_711,In_991);
and U778 (N_778,In_980,In_52);
nor U779 (N_779,In_857,In_242);
and U780 (N_780,In_992,In_903);
and U781 (N_781,In_979,In_656);
nor U782 (N_782,In_440,In_970);
and U783 (N_783,In_332,In_396);
nor U784 (N_784,In_544,In_794);
or U785 (N_785,In_251,In_489);
or U786 (N_786,In_225,In_297);
xnor U787 (N_787,In_359,In_736);
and U788 (N_788,In_641,In_671);
and U789 (N_789,In_822,In_110);
or U790 (N_790,In_111,In_517);
and U791 (N_791,In_626,In_335);
nand U792 (N_792,In_698,In_132);
nand U793 (N_793,In_750,In_751);
nor U794 (N_794,In_835,In_708);
or U795 (N_795,In_444,In_292);
nand U796 (N_796,In_901,In_598);
or U797 (N_797,In_867,In_373);
nor U798 (N_798,In_619,In_422);
xor U799 (N_799,In_399,In_626);
or U800 (N_800,In_395,In_135);
and U801 (N_801,In_323,In_668);
xnor U802 (N_802,In_24,In_249);
nor U803 (N_803,In_715,In_641);
or U804 (N_804,In_509,In_337);
nand U805 (N_805,In_438,In_171);
or U806 (N_806,In_207,In_771);
nor U807 (N_807,In_191,In_819);
and U808 (N_808,In_344,In_598);
or U809 (N_809,In_416,In_940);
xor U810 (N_810,In_329,In_558);
or U811 (N_811,In_726,In_638);
nand U812 (N_812,In_390,In_552);
nand U813 (N_813,In_76,In_782);
nand U814 (N_814,In_120,In_509);
nor U815 (N_815,In_992,In_614);
xnor U816 (N_816,In_976,In_624);
and U817 (N_817,In_582,In_846);
or U818 (N_818,In_512,In_884);
or U819 (N_819,In_923,In_390);
nor U820 (N_820,In_644,In_82);
or U821 (N_821,In_40,In_407);
nand U822 (N_822,In_91,In_251);
or U823 (N_823,In_326,In_863);
and U824 (N_824,In_935,In_562);
and U825 (N_825,In_268,In_592);
nand U826 (N_826,In_885,In_496);
and U827 (N_827,In_45,In_232);
and U828 (N_828,In_872,In_213);
and U829 (N_829,In_272,In_873);
and U830 (N_830,In_555,In_641);
nor U831 (N_831,In_768,In_704);
nor U832 (N_832,In_992,In_886);
nor U833 (N_833,In_335,In_278);
and U834 (N_834,In_396,In_977);
and U835 (N_835,In_406,In_858);
nand U836 (N_836,In_430,In_279);
and U837 (N_837,In_166,In_663);
nor U838 (N_838,In_416,In_774);
and U839 (N_839,In_585,In_654);
nand U840 (N_840,In_557,In_556);
nor U841 (N_841,In_48,In_874);
or U842 (N_842,In_344,In_937);
or U843 (N_843,In_290,In_538);
nand U844 (N_844,In_731,In_584);
and U845 (N_845,In_159,In_764);
nand U846 (N_846,In_755,In_136);
nand U847 (N_847,In_909,In_58);
nor U848 (N_848,In_377,In_277);
nor U849 (N_849,In_371,In_775);
nand U850 (N_850,In_68,In_898);
or U851 (N_851,In_239,In_175);
and U852 (N_852,In_884,In_912);
or U853 (N_853,In_571,In_720);
nor U854 (N_854,In_342,In_780);
nor U855 (N_855,In_880,In_847);
or U856 (N_856,In_948,In_367);
nand U857 (N_857,In_773,In_383);
xnor U858 (N_858,In_539,In_309);
and U859 (N_859,In_690,In_170);
nor U860 (N_860,In_351,In_702);
nand U861 (N_861,In_441,In_725);
nor U862 (N_862,In_985,In_177);
nor U863 (N_863,In_136,In_177);
nor U864 (N_864,In_459,In_335);
nand U865 (N_865,In_610,In_558);
nand U866 (N_866,In_390,In_958);
and U867 (N_867,In_472,In_985);
nor U868 (N_868,In_846,In_985);
and U869 (N_869,In_823,In_120);
nand U870 (N_870,In_49,In_427);
nand U871 (N_871,In_667,In_880);
and U872 (N_872,In_408,In_295);
or U873 (N_873,In_611,In_828);
nor U874 (N_874,In_735,In_651);
and U875 (N_875,In_846,In_241);
or U876 (N_876,In_130,In_340);
and U877 (N_877,In_5,In_701);
and U878 (N_878,In_602,In_619);
or U879 (N_879,In_743,In_761);
or U880 (N_880,In_852,In_503);
or U881 (N_881,In_401,In_301);
xnor U882 (N_882,In_653,In_919);
xor U883 (N_883,In_348,In_125);
or U884 (N_884,In_165,In_366);
nor U885 (N_885,In_138,In_553);
nor U886 (N_886,In_981,In_248);
nand U887 (N_887,In_283,In_711);
nor U888 (N_888,In_554,In_729);
nor U889 (N_889,In_827,In_518);
nor U890 (N_890,In_717,In_177);
and U891 (N_891,In_550,In_77);
nor U892 (N_892,In_464,In_418);
and U893 (N_893,In_839,In_723);
nor U894 (N_894,In_790,In_99);
or U895 (N_895,In_715,In_497);
or U896 (N_896,In_272,In_340);
nor U897 (N_897,In_157,In_197);
or U898 (N_898,In_149,In_154);
xor U899 (N_899,In_185,In_748);
xnor U900 (N_900,In_29,In_921);
xor U901 (N_901,In_63,In_866);
nand U902 (N_902,In_710,In_964);
xor U903 (N_903,In_361,In_638);
and U904 (N_904,In_993,In_435);
or U905 (N_905,In_9,In_582);
nand U906 (N_906,In_489,In_604);
and U907 (N_907,In_578,In_110);
nand U908 (N_908,In_110,In_766);
or U909 (N_909,In_418,In_853);
nand U910 (N_910,In_773,In_545);
or U911 (N_911,In_790,In_602);
or U912 (N_912,In_379,In_871);
and U913 (N_913,In_509,In_265);
nand U914 (N_914,In_488,In_832);
and U915 (N_915,In_1,In_139);
xor U916 (N_916,In_17,In_946);
nor U917 (N_917,In_562,In_989);
and U918 (N_918,In_502,In_639);
and U919 (N_919,In_558,In_926);
and U920 (N_920,In_840,In_757);
and U921 (N_921,In_68,In_491);
nor U922 (N_922,In_752,In_847);
nand U923 (N_923,In_561,In_776);
nand U924 (N_924,In_646,In_819);
and U925 (N_925,In_222,In_735);
nand U926 (N_926,In_574,In_20);
nand U927 (N_927,In_704,In_51);
and U928 (N_928,In_17,In_339);
and U929 (N_929,In_944,In_617);
or U930 (N_930,In_383,In_650);
xnor U931 (N_931,In_377,In_471);
and U932 (N_932,In_173,In_462);
nand U933 (N_933,In_846,In_826);
nor U934 (N_934,In_443,In_10);
and U935 (N_935,In_193,In_319);
nor U936 (N_936,In_472,In_91);
nor U937 (N_937,In_846,In_78);
and U938 (N_938,In_844,In_940);
nor U939 (N_939,In_920,In_243);
nor U940 (N_940,In_919,In_275);
and U941 (N_941,In_815,In_465);
xnor U942 (N_942,In_913,In_90);
and U943 (N_943,In_859,In_7);
nor U944 (N_944,In_899,In_70);
nor U945 (N_945,In_872,In_419);
nand U946 (N_946,In_666,In_191);
nand U947 (N_947,In_493,In_428);
and U948 (N_948,In_464,In_413);
nor U949 (N_949,In_718,In_269);
or U950 (N_950,In_406,In_21);
nor U951 (N_951,In_400,In_414);
and U952 (N_952,In_260,In_973);
and U953 (N_953,In_766,In_864);
and U954 (N_954,In_723,In_949);
and U955 (N_955,In_862,In_285);
and U956 (N_956,In_498,In_554);
or U957 (N_957,In_680,In_607);
nand U958 (N_958,In_657,In_554);
or U959 (N_959,In_831,In_236);
nand U960 (N_960,In_13,In_228);
nor U961 (N_961,In_551,In_91);
nor U962 (N_962,In_470,In_522);
nand U963 (N_963,In_333,In_135);
nor U964 (N_964,In_268,In_785);
or U965 (N_965,In_553,In_297);
or U966 (N_966,In_792,In_237);
and U967 (N_967,In_927,In_429);
nor U968 (N_968,In_673,In_498);
or U969 (N_969,In_840,In_925);
nor U970 (N_970,In_620,In_420);
or U971 (N_971,In_815,In_202);
nand U972 (N_972,In_160,In_657);
nand U973 (N_973,In_717,In_404);
or U974 (N_974,In_720,In_39);
xor U975 (N_975,In_934,In_462);
or U976 (N_976,In_686,In_87);
and U977 (N_977,In_426,In_959);
or U978 (N_978,In_793,In_202);
nor U979 (N_979,In_897,In_499);
xnor U980 (N_980,In_201,In_674);
and U981 (N_981,In_267,In_332);
nand U982 (N_982,In_157,In_254);
nor U983 (N_983,In_888,In_962);
nor U984 (N_984,In_902,In_501);
nand U985 (N_985,In_50,In_493);
nor U986 (N_986,In_286,In_573);
nor U987 (N_987,In_675,In_796);
nand U988 (N_988,In_422,In_604);
or U989 (N_989,In_850,In_900);
and U990 (N_990,In_941,In_824);
and U991 (N_991,In_433,In_719);
nor U992 (N_992,In_124,In_644);
or U993 (N_993,In_797,In_756);
and U994 (N_994,In_233,In_373);
and U995 (N_995,In_318,In_325);
or U996 (N_996,In_234,In_577);
or U997 (N_997,In_542,In_635);
nor U998 (N_998,In_599,In_988);
nand U999 (N_999,In_26,In_450);
and U1000 (N_1000,In_707,In_998);
nand U1001 (N_1001,In_86,In_999);
and U1002 (N_1002,In_872,In_914);
nand U1003 (N_1003,In_945,In_619);
and U1004 (N_1004,In_463,In_537);
or U1005 (N_1005,In_641,In_699);
or U1006 (N_1006,In_186,In_409);
nand U1007 (N_1007,In_207,In_69);
or U1008 (N_1008,In_696,In_651);
nor U1009 (N_1009,In_248,In_381);
xor U1010 (N_1010,In_368,In_904);
xor U1011 (N_1011,In_982,In_987);
and U1012 (N_1012,In_539,In_489);
nand U1013 (N_1013,In_754,In_200);
and U1014 (N_1014,In_572,In_465);
nor U1015 (N_1015,In_309,In_89);
nor U1016 (N_1016,In_971,In_114);
nor U1017 (N_1017,In_701,In_939);
nor U1018 (N_1018,In_358,In_298);
nand U1019 (N_1019,In_395,In_495);
nor U1020 (N_1020,In_821,In_126);
nand U1021 (N_1021,In_799,In_381);
and U1022 (N_1022,In_897,In_250);
or U1023 (N_1023,In_882,In_23);
or U1024 (N_1024,In_508,In_679);
or U1025 (N_1025,In_915,In_271);
nor U1026 (N_1026,In_56,In_62);
and U1027 (N_1027,In_549,In_314);
nor U1028 (N_1028,In_912,In_919);
and U1029 (N_1029,In_322,In_388);
or U1030 (N_1030,In_361,In_573);
and U1031 (N_1031,In_975,In_385);
and U1032 (N_1032,In_966,In_142);
and U1033 (N_1033,In_702,In_9);
or U1034 (N_1034,In_383,In_417);
and U1035 (N_1035,In_740,In_227);
nor U1036 (N_1036,In_172,In_257);
nor U1037 (N_1037,In_990,In_735);
or U1038 (N_1038,In_361,In_599);
or U1039 (N_1039,In_171,In_741);
nor U1040 (N_1040,In_519,In_758);
nand U1041 (N_1041,In_993,In_526);
xor U1042 (N_1042,In_211,In_67);
nor U1043 (N_1043,In_137,In_27);
nor U1044 (N_1044,In_450,In_851);
and U1045 (N_1045,In_559,In_857);
or U1046 (N_1046,In_774,In_682);
and U1047 (N_1047,In_787,In_512);
nand U1048 (N_1048,In_295,In_800);
nor U1049 (N_1049,In_688,In_655);
or U1050 (N_1050,In_987,In_306);
xnor U1051 (N_1051,In_486,In_281);
and U1052 (N_1052,In_95,In_20);
nand U1053 (N_1053,In_315,In_264);
and U1054 (N_1054,In_761,In_990);
nor U1055 (N_1055,In_734,In_963);
and U1056 (N_1056,In_387,In_929);
and U1057 (N_1057,In_548,In_422);
and U1058 (N_1058,In_286,In_802);
nand U1059 (N_1059,In_292,In_891);
and U1060 (N_1060,In_73,In_72);
and U1061 (N_1061,In_258,In_514);
or U1062 (N_1062,In_165,In_378);
xor U1063 (N_1063,In_761,In_691);
and U1064 (N_1064,In_800,In_648);
or U1065 (N_1065,In_836,In_488);
nand U1066 (N_1066,In_169,In_922);
nand U1067 (N_1067,In_507,In_993);
and U1068 (N_1068,In_144,In_701);
xnor U1069 (N_1069,In_744,In_243);
xnor U1070 (N_1070,In_867,In_956);
nor U1071 (N_1071,In_847,In_624);
nand U1072 (N_1072,In_903,In_186);
and U1073 (N_1073,In_508,In_929);
or U1074 (N_1074,In_816,In_344);
nor U1075 (N_1075,In_838,In_91);
or U1076 (N_1076,In_569,In_238);
xnor U1077 (N_1077,In_305,In_349);
and U1078 (N_1078,In_429,In_998);
and U1079 (N_1079,In_274,In_374);
or U1080 (N_1080,In_411,In_537);
or U1081 (N_1081,In_29,In_61);
nor U1082 (N_1082,In_202,In_7);
or U1083 (N_1083,In_46,In_847);
nor U1084 (N_1084,In_926,In_426);
nor U1085 (N_1085,In_485,In_89);
nand U1086 (N_1086,In_380,In_615);
xor U1087 (N_1087,In_604,In_162);
and U1088 (N_1088,In_249,In_63);
nor U1089 (N_1089,In_472,In_587);
or U1090 (N_1090,In_738,In_677);
nor U1091 (N_1091,In_694,In_33);
and U1092 (N_1092,In_475,In_753);
nor U1093 (N_1093,In_835,In_892);
or U1094 (N_1094,In_614,In_617);
nand U1095 (N_1095,In_736,In_469);
nand U1096 (N_1096,In_585,In_534);
and U1097 (N_1097,In_845,In_92);
nand U1098 (N_1098,In_543,In_632);
or U1099 (N_1099,In_8,In_542);
nand U1100 (N_1100,In_935,In_745);
or U1101 (N_1101,In_790,In_707);
and U1102 (N_1102,In_178,In_796);
nor U1103 (N_1103,In_561,In_89);
xnor U1104 (N_1104,In_934,In_83);
nand U1105 (N_1105,In_976,In_696);
or U1106 (N_1106,In_898,In_938);
and U1107 (N_1107,In_669,In_804);
nor U1108 (N_1108,In_529,In_28);
nand U1109 (N_1109,In_714,In_800);
and U1110 (N_1110,In_169,In_452);
and U1111 (N_1111,In_548,In_734);
nor U1112 (N_1112,In_656,In_770);
nand U1113 (N_1113,In_500,In_290);
or U1114 (N_1114,In_51,In_471);
or U1115 (N_1115,In_806,In_581);
nand U1116 (N_1116,In_331,In_961);
nand U1117 (N_1117,In_226,In_527);
nor U1118 (N_1118,In_980,In_80);
nor U1119 (N_1119,In_929,In_477);
nor U1120 (N_1120,In_214,In_373);
and U1121 (N_1121,In_530,In_111);
xor U1122 (N_1122,In_858,In_527);
and U1123 (N_1123,In_767,In_961);
nand U1124 (N_1124,In_179,In_95);
and U1125 (N_1125,In_410,In_635);
nor U1126 (N_1126,In_39,In_671);
nor U1127 (N_1127,In_952,In_365);
nand U1128 (N_1128,In_986,In_184);
nor U1129 (N_1129,In_57,In_874);
nand U1130 (N_1130,In_294,In_960);
nor U1131 (N_1131,In_973,In_50);
nor U1132 (N_1132,In_642,In_336);
nor U1133 (N_1133,In_497,In_72);
nand U1134 (N_1134,In_806,In_390);
nand U1135 (N_1135,In_101,In_575);
xnor U1136 (N_1136,In_327,In_774);
or U1137 (N_1137,In_716,In_899);
nor U1138 (N_1138,In_456,In_869);
and U1139 (N_1139,In_774,In_975);
and U1140 (N_1140,In_428,In_309);
or U1141 (N_1141,In_234,In_846);
nand U1142 (N_1142,In_57,In_290);
or U1143 (N_1143,In_404,In_376);
and U1144 (N_1144,In_713,In_960);
and U1145 (N_1145,In_103,In_953);
xor U1146 (N_1146,In_62,In_640);
and U1147 (N_1147,In_296,In_67);
and U1148 (N_1148,In_275,In_685);
nor U1149 (N_1149,In_609,In_432);
nand U1150 (N_1150,In_783,In_478);
nand U1151 (N_1151,In_309,In_869);
nor U1152 (N_1152,In_54,In_201);
and U1153 (N_1153,In_363,In_156);
or U1154 (N_1154,In_155,In_931);
nor U1155 (N_1155,In_194,In_510);
or U1156 (N_1156,In_783,In_53);
or U1157 (N_1157,In_133,In_761);
and U1158 (N_1158,In_817,In_856);
or U1159 (N_1159,In_86,In_846);
nor U1160 (N_1160,In_951,In_569);
and U1161 (N_1161,In_660,In_874);
nor U1162 (N_1162,In_58,In_9);
nand U1163 (N_1163,In_85,In_202);
nand U1164 (N_1164,In_739,In_253);
and U1165 (N_1165,In_316,In_586);
nand U1166 (N_1166,In_572,In_509);
and U1167 (N_1167,In_49,In_979);
and U1168 (N_1168,In_526,In_71);
xor U1169 (N_1169,In_387,In_73);
and U1170 (N_1170,In_332,In_23);
nor U1171 (N_1171,In_155,In_478);
nand U1172 (N_1172,In_226,In_402);
xnor U1173 (N_1173,In_435,In_625);
or U1174 (N_1174,In_751,In_39);
and U1175 (N_1175,In_578,In_119);
nor U1176 (N_1176,In_312,In_830);
or U1177 (N_1177,In_327,In_196);
or U1178 (N_1178,In_275,In_853);
nand U1179 (N_1179,In_490,In_1);
nor U1180 (N_1180,In_765,In_863);
and U1181 (N_1181,In_307,In_139);
or U1182 (N_1182,In_807,In_138);
nand U1183 (N_1183,In_693,In_679);
nor U1184 (N_1184,In_935,In_120);
and U1185 (N_1185,In_830,In_753);
nor U1186 (N_1186,In_892,In_879);
nor U1187 (N_1187,In_311,In_609);
and U1188 (N_1188,In_952,In_610);
nor U1189 (N_1189,In_583,In_763);
or U1190 (N_1190,In_372,In_638);
and U1191 (N_1191,In_385,In_668);
or U1192 (N_1192,In_787,In_666);
nor U1193 (N_1193,In_523,In_609);
and U1194 (N_1194,In_64,In_465);
and U1195 (N_1195,In_844,In_905);
or U1196 (N_1196,In_39,In_596);
or U1197 (N_1197,In_618,In_563);
and U1198 (N_1198,In_739,In_235);
or U1199 (N_1199,In_922,In_717);
or U1200 (N_1200,In_537,In_403);
nor U1201 (N_1201,In_921,In_926);
or U1202 (N_1202,In_425,In_422);
or U1203 (N_1203,In_94,In_889);
xnor U1204 (N_1204,In_292,In_153);
and U1205 (N_1205,In_861,In_844);
nor U1206 (N_1206,In_191,In_988);
and U1207 (N_1207,In_976,In_29);
or U1208 (N_1208,In_787,In_552);
or U1209 (N_1209,In_791,In_315);
nor U1210 (N_1210,In_760,In_217);
xnor U1211 (N_1211,In_981,In_57);
and U1212 (N_1212,In_631,In_12);
nand U1213 (N_1213,In_752,In_979);
nand U1214 (N_1214,In_94,In_738);
xnor U1215 (N_1215,In_916,In_834);
and U1216 (N_1216,In_137,In_543);
nor U1217 (N_1217,In_439,In_234);
xnor U1218 (N_1218,In_40,In_299);
nand U1219 (N_1219,In_345,In_524);
nand U1220 (N_1220,In_492,In_857);
nor U1221 (N_1221,In_261,In_456);
or U1222 (N_1222,In_691,In_742);
nand U1223 (N_1223,In_607,In_828);
nor U1224 (N_1224,In_470,In_333);
xnor U1225 (N_1225,In_848,In_844);
nand U1226 (N_1226,In_956,In_642);
and U1227 (N_1227,In_827,In_420);
nand U1228 (N_1228,In_984,In_41);
nor U1229 (N_1229,In_402,In_793);
or U1230 (N_1230,In_288,In_35);
nand U1231 (N_1231,In_570,In_532);
or U1232 (N_1232,In_789,In_22);
nand U1233 (N_1233,In_240,In_701);
nor U1234 (N_1234,In_953,In_702);
nand U1235 (N_1235,In_336,In_806);
and U1236 (N_1236,In_479,In_427);
or U1237 (N_1237,In_531,In_864);
and U1238 (N_1238,In_281,In_213);
nor U1239 (N_1239,In_255,In_978);
or U1240 (N_1240,In_105,In_442);
or U1241 (N_1241,In_643,In_155);
nor U1242 (N_1242,In_166,In_770);
and U1243 (N_1243,In_523,In_722);
nor U1244 (N_1244,In_881,In_638);
and U1245 (N_1245,In_600,In_28);
or U1246 (N_1246,In_786,In_617);
nand U1247 (N_1247,In_635,In_482);
nand U1248 (N_1248,In_253,In_369);
and U1249 (N_1249,In_402,In_295);
nor U1250 (N_1250,In_348,In_820);
nand U1251 (N_1251,In_257,In_271);
and U1252 (N_1252,In_473,In_132);
and U1253 (N_1253,In_682,In_14);
and U1254 (N_1254,In_293,In_869);
nor U1255 (N_1255,In_422,In_485);
nor U1256 (N_1256,In_610,In_58);
nor U1257 (N_1257,In_919,In_9);
nand U1258 (N_1258,In_397,In_186);
nand U1259 (N_1259,In_11,In_583);
nand U1260 (N_1260,In_938,In_316);
xnor U1261 (N_1261,In_2,In_79);
nor U1262 (N_1262,In_612,In_315);
nand U1263 (N_1263,In_129,In_327);
nor U1264 (N_1264,In_875,In_142);
and U1265 (N_1265,In_318,In_38);
and U1266 (N_1266,In_583,In_904);
or U1267 (N_1267,In_559,In_618);
or U1268 (N_1268,In_669,In_284);
nor U1269 (N_1269,In_940,In_444);
and U1270 (N_1270,In_822,In_255);
nand U1271 (N_1271,In_187,In_508);
nor U1272 (N_1272,In_132,In_815);
nand U1273 (N_1273,In_291,In_11);
or U1274 (N_1274,In_613,In_842);
or U1275 (N_1275,In_127,In_285);
nand U1276 (N_1276,In_418,In_771);
nand U1277 (N_1277,In_231,In_254);
and U1278 (N_1278,In_42,In_455);
nor U1279 (N_1279,In_892,In_308);
nand U1280 (N_1280,In_449,In_731);
and U1281 (N_1281,In_433,In_297);
nor U1282 (N_1282,In_330,In_630);
xnor U1283 (N_1283,In_337,In_637);
nor U1284 (N_1284,In_865,In_756);
nand U1285 (N_1285,In_718,In_806);
xnor U1286 (N_1286,In_440,In_4);
nand U1287 (N_1287,In_626,In_272);
xnor U1288 (N_1288,In_75,In_286);
xor U1289 (N_1289,In_903,In_564);
and U1290 (N_1290,In_316,In_948);
or U1291 (N_1291,In_430,In_116);
nor U1292 (N_1292,In_412,In_288);
or U1293 (N_1293,In_667,In_862);
xor U1294 (N_1294,In_898,In_40);
nand U1295 (N_1295,In_314,In_787);
nand U1296 (N_1296,In_969,In_115);
nand U1297 (N_1297,In_576,In_51);
or U1298 (N_1298,In_837,In_755);
nand U1299 (N_1299,In_862,In_558);
or U1300 (N_1300,In_776,In_603);
nor U1301 (N_1301,In_449,In_221);
and U1302 (N_1302,In_809,In_162);
xnor U1303 (N_1303,In_46,In_146);
or U1304 (N_1304,In_263,In_546);
and U1305 (N_1305,In_684,In_189);
xnor U1306 (N_1306,In_947,In_546);
nor U1307 (N_1307,In_433,In_558);
nand U1308 (N_1308,In_520,In_15);
nand U1309 (N_1309,In_42,In_183);
nand U1310 (N_1310,In_468,In_725);
or U1311 (N_1311,In_416,In_484);
nor U1312 (N_1312,In_437,In_133);
and U1313 (N_1313,In_390,In_922);
nand U1314 (N_1314,In_794,In_108);
nand U1315 (N_1315,In_104,In_607);
nand U1316 (N_1316,In_369,In_97);
and U1317 (N_1317,In_441,In_473);
or U1318 (N_1318,In_523,In_533);
or U1319 (N_1319,In_605,In_398);
and U1320 (N_1320,In_994,In_892);
nand U1321 (N_1321,In_345,In_979);
nor U1322 (N_1322,In_232,In_865);
nand U1323 (N_1323,In_859,In_278);
nor U1324 (N_1324,In_130,In_752);
xnor U1325 (N_1325,In_50,In_836);
and U1326 (N_1326,In_500,In_531);
and U1327 (N_1327,In_32,In_203);
nand U1328 (N_1328,In_829,In_155);
or U1329 (N_1329,In_335,In_732);
xor U1330 (N_1330,In_173,In_297);
nor U1331 (N_1331,In_796,In_74);
nand U1332 (N_1332,In_905,In_704);
or U1333 (N_1333,In_492,In_35);
and U1334 (N_1334,In_723,In_131);
and U1335 (N_1335,In_931,In_230);
nor U1336 (N_1336,In_649,In_184);
and U1337 (N_1337,In_690,In_151);
nand U1338 (N_1338,In_161,In_307);
and U1339 (N_1339,In_344,In_95);
or U1340 (N_1340,In_13,In_180);
nand U1341 (N_1341,In_572,In_817);
nor U1342 (N_1342,In_639,In_718);
and U1343 (N_1343,In_127,In_27);
and U1344 (N_1344,In_127,In_162);
and U1345 (N_1345,In_492,In_348);
nand U1346 (N_1346,In_793,In_260);
nor U1347 (N_1347,In_25,In_405);
nor U1348 (N_1348,In_484,In_308);
nor U1349 (N_1349,In_142,In_624);
nor U1350 (N_1350,In_811,In_296);
or U1351 (N_1351,In_801,In_605);
nand U1352 (N_1352,In_973,In_970);
nor U1353 (N_1353,In_328,In_726);
nand U1354 (N_1354,In_846,In_261);
and U1355 (N_1355,In_496,In_767);
nand U1356 (N_1356,In_572,In_507);
or U1357 (N_1357,In_612,In_701);
or U1358 (N_1358,In_462,In_505);
xor U1359 (N_1359,In_566,In_986);
nand U1360 (N_1360,In_274,In_137);
nand U1361 (N_1361,In_931,In_732);
or U1362 (N_1362,In_888,In_518);
and U1363 (N_1363,In_552,In_23);
nor U1364 (N_1364,In_374,In_858);
or U1365 (N_1365,In_664,In_502);
or U1366 (N_1366,In_613,In_827);
nor U1367 (N_1367,In_954,In_334);
nand U1368 (N_1368,In_23,In_762);
nand U1369 (N_1369,In_448,In_643);
and U1370 (N_1370,In_749,In_910);
nand U1371 (N_1371,In_37,In_41);
or U1372 (N_1372,In_520,In_766);
xnor U1373 (N_1373,In_253,In_227);
nand U1374 (N_1374,In_103,In_201);
or U1375 (N_1375,In_866,In_564);
and U1376 (N_1376,In_695,In_653);
or U1377 (N_1377,In_90,In_60);
or U1378 (N_1378,In_31,In_105);
and U1379 (N_1379,In_79,In_130);
or U1380 (N_1380,In_143,In_959);
xnor U1381 (N_1381,In_122,In_784);
nand U1382 (N_1382,In_144,In_320);
xor U1383 (N_1383,In_181,In_243);
and U1384 (N_1384,In_559,In_490);
xnor U1385 (N_1385,In_710,In_130);
and U1386 (N_1386,In_109,In_345);
xnor U1387 (N_1387,In_357,In_338);
or U1388 (N_1388,In_201,In_113);
nor U1389 (N_1389,In_368,In_373);
nor U1390 (N_1390,In_566,In_275);
nand U1391 (N_1391,In_746,In_959);
or U1392 (N_1392,In_238,In_629);
nor U1393 (N_1393,In_623,In_347);
nor U1394 (N_1394,In_921,In_561);
and U1395 (N_1395,In_906,In_744);
nor U1396 (N_1396,In_457,In_14);
and U1397 (N_1397,In_715,In_719);
and U1398 (N_1398,In_512,In_385);
or U1399 (N_1399,In_668,In_620);
nor U1400 (N_1400,In_976,In_846);
and U1401 (N_1401,In_43,In_171);
or U1402 (N_1402,In_640,In_664);
nand U1403 (N_1403,In_871,In_81);
and U1404 (N_1404,In_855,In_596);
nand U1405 (N_1405,In_911,In_933);
nand U1406 (N_1406,In_184,In_662);
nor U1407 (N_1407,In_668,In_438);
or U1408 (N_1408,In_10,In_316);
nand U1409 (N_1409,In_717,In_693);
nand U1410 (N_1410,In_641,In_218);
or U1411 (N_1411,In_235,In_826);
nor U1412 (N_1412,In_377,In_922);
or U1413 (N_1413,In_532,In_995);
or U1414 (N_1414,In_644,In_743);
and U1415 (N_1415,In_103,In_387);
nor U1416 (N_1416,In_371,In_824);
or U1417 (N_1417,In_13,In_544);
nand U1418 (N_1418,In_151,In_61);
and U1419 (N_1419,In_407,In_94);
nand U1420 (N_1420,In_31,In_338);
xor U1421 (N_1421,In_434,In_465);
and U1422 (N_1422,In_317,In_108);
nor U1423 (N_1423,In_752,In_219);
nor U1424 (N_1424,In_912,In_839);
and U1425 (N_1425,In_774,In_991);
and U1426 (N_1426,In_731,In_218);
and U1427 (N_1427,In_698,In_921);
nor U1428 (N_1428,In_866,In_611);
or U1429 (N_1429,In_843,In_870);
or U1430 (N_1430,In_78,In_318);
or U1431 (N_1431,In_166,In_150);
or U1432 (N_1432,In_572,In_823);
or U1433 (N_1433,In_136,In_542);
nor U1434 (N_1434,In_923,In_417);
nor U1435 (N_1435,In_742,In_856);
nand U1436 (N_1436,In_557,In_730);
nor U1437 (N_1437,In_784,In_124);
or U1438 (N_1438,In_825,In_561);
or U1439 (N_1439,In_723,In_935);
nor U1440 (N_1440,In_866,In_986);
nand U1441 (N_1441,In_207,In_26);
and U1442 (N_1442,In_788,In_992);
nand U1443 (N_1443,In_797,In_483);
or U1444 (N_1444,In_168,In_396);
or U1445 (N_1445,In_974,In_200);
nor U1446 (N_1446,In_144,In_229);
xnor U1447 (N_1447,In_962,In_178);
nor U1448 (N_1448,In_208,In_603);
and U1449 (N_1449,In_469,In_81);
and U1450 (N_1450,In_843,In_294);
and U1451 (N_1451,In_68,In_593);
xnor U1452 (N_1452,In_830,In_359);
nor U1453 (N_1453,In_735,In_766);
or U1454 (N_1454,In_555,In_639);
or U1455 (N_1455,In_907,In_864);
or U1456 (N_1456,In_935,In_503);
nor U1457 (N_1457,In_771,In_351);
or U1458 (N_1458,In_608,In_260);
xor U1459 (N_1459,In_472,In_284);
or U1460 (N_1460,In_627,In_148);
xnor U1461 (N_1461,In_516,In_358);
nand U1462 (N_1462,In_35,In_366);
and U1463 (N_1463,In_305,In_406);
nand U1464 (N_1464,In_677,In_408);
and U1465 (N_1465,In_709,In_211);
nor U1466 (N_1466,In_619,In_374);
or U1467 (N_1467,In_124,In_988);
or U1468 (N_1468,In_522,In_263);
nor U1469 (N_1469,In_446,In_870);
nand U1470 (N_1470,In_638,In_500);
nand U1471 (N_1471,In_339,In_441);
nand U1472 (N_1472,In_148,In_676);
xor U1473 (N_1473,In_66,In_188);
or U1474 (N_1474,In_383,In_472);
nand U1475 (N_1475,In_275,In_384);
nand U1476 (N_1476,In_540,In_81);
nand U1477 (N_1477,In_446,In_900);
and U1478 (N_1478,In_831,In_407);
nand U1479 (N_1479,In_326,In_752);
or U1480 (N_1480,In_688,In_438);
or U1481 (N_1481,In_911,In_690);
nor U1482 (N_1482,In_565,In_974);
or U1483 (N_1483,In_431,In_749);
nor U1484 (N_1484,In_123,In_498);
nand U1485 (N_1485,In_748,In_805);
xnor U1486 (N_1486,In_462,In_366);
nand U1487 (N_1487,In_565,In_834);
or U1488 (N_1488,In_514,In_684);
or U1489 (N_1489,In_527,In_440);
or U1490 (N_1490,In_145,In_580);
nor U1491 (N_1491,In_55,In_958);
or U1492 (N_1492,In_631,In_769);
nor U1493 (N_1493,In_773,In_284);
nor U1494 (N_1494,In_313,In_355);
nand U1495 (N_1495,In_695,In_460);
or U1496 (N_1496,In_471,In_709);
or U1497 (N_1497,In_453,In_409);
nor U1498 (N_1498,In_758,In_522);
nand U1499 (N_1499,In_226,In_131);
nand U1500 (N_1500,In_656,In_487);
and U1501 (N_1501,In_660,In_869);
nand U1502 (N_1502,In_90,In_943);
or U1503 (N_1503,In_120,In_872);
nor U1504 (N_1504,In_55,In_63);
nor U1505 (N_1505,In_947,In_181);
nand U1506 (N_1506,In_713,In_755);
nor U1507 (N_1507,In_541,In_806);
or U1508 (N_1508,In_356,In_722);
nand U1509 (N_1509,In_980,In_72);
nand U1510 (N_1510,In_141,In_918);
nor U1511 (N_1511,In_690,In_594);
nand U1512 (N_1512,In_115,In_465);
nand U1513 (N_1513,In_120,In_108);
or U1514 (N_1514,In_837,In_941);
and U1515 (N_1515,In_567,In_58);
and U1516 (N_1516,In_676,In_902);
nor U1517 (N_1517,In_487,In_126);
and U1518 (N_1518,In_515,In_183);
and U1519 (N_1519,In_560,In_156);
or U1520 (N_1520,In_981,In_517);
or U1521 (N_1521,In_759,In_303);
nand U1522 (N_1522,In_248,In_780);
nor U1523 (N_1523,In_321,In_325);
nor U1524 (N_1524,In_463,In_663);
nand U1525 (N_1525,In_816,In_678);
or U1526 (N_1526,In_845,In_739);
nand U1527 (N_1527,In_282,In_872);
or U1528 (N_1528,In_369,In_752);
and U1529 (N_1529,In_939,In_247);
nand U1530 (N_1530,In_537,In_998);
xor U1531 (N_1531,In_522,In_437);
nand U1532 (N_1532,In_450,In_657);
nor U1533 (N_1533,In_497,In_743);
and U1534 (N_1534,In_528,In_148);
nor U1535 (N_1535,In_494,In_423);
nand U1536 (N_1536,In_171,In_84);
nor U1537 (N_1537,In_562,In_141);
and U1538 (N_1538,In_92,In_660);
nand U1539 (N_1539,In_602,In_823);
and U1540 (N_1540,In_23,In_103);
or U1541 (N_1541,In_543,In_701);
nand U1542 (N_1542,In_720,In_575);
or U1543 (N_1543,In_857,In_201);
or U1544 (N_1544,In_503,In_547);
nor U1545 (N_1545,In_635,In_525);
or U1546 (N_1546,In_402,In_129);
or U1547 (N_1547,In_802,In_561);
or U1548 (N_1548,In_195,In_984);
nand U1549 (N_1549,In_687,In_517);
nand U1550 (N_1550,In_147,In_43);
and U1551 (N_1551,In_668,In_276);
nor U1552 (N_1552,In_828,In_864);
nor U1553 (N_1553,In_994,In_917);
xor U1554 (N_1554,In_797,In_208);
and U1555 (N_1555,In_566,In_389);
nor U1556 (N_1556,In_709,In_523);
or U1557 (N_1557,In_15,In_298);
or U1558 (N_1558,In_658,In_639);
and U1559 (N_1559,In_841,In_707);
xnor U1560 (N_1560,In_547,In_73);
or U1561 (N_1561,In_100,In_155);
nand U1562 (N_1562,In_866,In_617);
nor U1563 (N_1563,In_550,In_907);
and U1564 (N_1564,In_899,In_445);
nand U1565 (N_1565,In_43,In_638);
nand U1566 (N_1566,In_792,In_924);
and U1567 (N_1567,In_758,In_833);
or U1568 (N_1568,In_201,In_980);
nand U1569 (N_1569,In_589,In_696);
and U1570 (N_1570,In_456,In_895);
or U1571 (N_1571,In_298,In_972);
nand U1572 (N_1572,In_843,In_770);
and U1573 (N_1573,In_659,In_714);
and U1574 (N_1574,In_947,In_548);
or U1575 (N_1575,In_266,In_554);
or U1576 (N_1576,In_513,In_607);
nor U1577 (N_1577,In_651,In_180);
xnor U1578 (N_1578,In_461,In_455);
and U1579 (N_1579,In_541,In_842);
or U1580 (N_1580,In_298,In_237);
or U1581 (N_1581,In_146,In_390);
nor U1582 (N_1582,In_826,In_53);
xor U1583 (N_1583,In_797,In_710);
or U1584 (N_1584,In_993,In_710);
nand U1585 (N_1585,In_941,In_421);
xnor U1586 (N_1586,In_792,In_616);
xnor U1587 (N_1587,In_442,In_863);
or U1588 (N_1588,In_859,In_999);
or U1589 (N_1589,In_58,In_0);
nand U1590 (N_1590,In_389,In_676);
or U1591 (N_1591,In_863,In_998);
nor U1592 (N_1592,In_351,In_960);
or U1593 (N_1593,In_313,In_966);
and U1594 (N_1594,In_393,In_435);
and U1595 (N_1595,In_72,In_411);
or U1596 (N_1596,In_131,In_709);
nor U1597 (N_1597,In_202,In_501);
or U1598 (N_1598,In_251,In_874);
nand U1599 (N_1599,In_279,In_448);
or U1600 (N_1600,In_906,In_299);
or U1601 (N_1601,In_75,In_264);
nor U1602 (N_1602,In_228,In_816);
and U1603 (N_1603,In_439,In_494);
and U1604 (N_1604,In_537,In_235);
or U1605 (N_1605,In_724,In_192);
nor U1606 (N_1606,In_997,In_356);
nor U1607 (N_1607,In_356,In_416);
and U1608 (N_1608,In_6,In_611);
xor U1609 (N_1609,In_756,In_549);
nand U1610 (N_1610,In_16,In_37);
or U1611 (N_1611,In_963,In_365);
xnor U1612 (N_1612,In_663,In_283);
nand U1613 (N_1613,In_397,In_894);
nand U1614 (N_1614,In_625,In_114);
and U1615 (N_1615,In_702,In_733);
xnor U1616 (N_1616,In_716,In_406);
nor U1617 (N_1617,In_461,In_588);
and U1618 (N_1618,In_992,In_644);
and U1619 (N_1619,In_363,In_288);
and U1620 (N_1620,In_112,In_849);
or U1621 (N_1621,In_700,In_412);
nor U1622 (N_1622,In_983,In_36);
nor U1623 (N_1623,In_557,In_761);
or U1624 (N_1624,In_307,In_34);
and U1625 (N_1625,In_458,In_291);
xor U1626 (N_1626,In_6,In_942);
and U1627 (N_1627,In_364,In_572);
or U1628 (N_1628,In_520,In_620);
and U1629 (N_1629,In_477,In_224);
nand U1630 (N_1630,In_337,In_295);
nand U1631 (N_1631,In_194,In_402);
or U1632 (N_1632,In_579,In_996);
nand U1633 (N_1633,In_625,In_112);
or U1634 (N_1634,In_697,In_566);
and U1635 (N_1635,In_824,In_80);
and U1636 (N_1636,In_594,In_108);
or U1637 (N_1637,In_477,In_586);
or U1638 (N_1638,In_316,In_646);
nor U1639 (N_1639,In_877,In_924);
and U1640 (N_1640,In_554,In_616);
nand U1641 (N_1641,In_789,In_217);
or U1642 (N_1642,In_517,In_356);
nor U1643 (N_1643,In_287,In_201);
xnor U1644 (N_1644,In_971,In_39);
nand U1645 (N_1645,In_563,In_92);
nand U1646 (N_1646,In_662,In_692);
xnor U1647 (N_1647,In_841,In_626);
nor U1648 (N_1648,In_368,In_705);
nor U1649 (N_1649,In_471,In_978);
nand U1650 (N_1650,In_943,In_809);
nand U1651 (N_1651,In_903,In_770);
nand U1652 (N_1652,In_672,In_696);
nand U1653 (N_1653,In_358,In_843);
or U1654 (N_1654,In_71,In_647);
nand U1655 (N_1655,In_767,In_533);
xor U1656 (N_1656,In_916,In_137);
nor U1657 (N_1657,In_601,In_22);
nor U1658 (N_1658,In_928,In_699);
nor U1659 (N_1659,In_157,In_393);
and U1660 (N_1660,In_128,In_903);
or U1661 (N_1661,In_829,In_960);
nor U1662 (N_1662,In_466,In_262);
and U1663 (N_1663,In_624,In_411);
nand U1664 (N_1664,In_222,In_791);
and U1665 (N_1665,In_149,In_739);
or U1666 (N_1666,In_679,In_293);
nor U1667 (N_1667,In_657,In_70);
or U1668 (N_1668,In_787,In_271);
and U1669 (N_1669,In_866,In_142);
xor U1670 (N_1670,In_795,In_209);
and U1671 (N_1671,In_599,In_113);
nor U1672 (N_1672,In_512,In_192);
nor U1673 (N_1673,In_811,In_932);
and U1674 (N_1674,In_39,In_89);
nor U1675 (N_1675,In_541,In_657);
and U1676 (N_1676,In_305,In_870);
and U1677 (N_1677,In_187,In_925);
or U1678 (N_1678,In_226,In_62);
nor U1679 (N_1679,In_259,In_240);
nand U1680 (N_1680,In_895,In_465);
nand U1681 (N_1681,In_156,In_966);
nor U1682 (N_1682,In_562,In_931);
and U1683 (N_1683,In_531,In_636);
nor U1684 (N_1684,In_921,In_196);
nand U1685 (N_1685,In_465,In_497);
xor U1686 (N_1686,In_632,In_991);
and U1687 (N_1687,In_699,In_327);
and U1688 (N_1688,In_571,In_818);
or U1689 (N_1689,In_536,In_991);
nor U1690 (N_1690,In_893,In_486);
nor U1691 (N_1691,In_66,In_803);
and U1692 (N_1692,In_499,In_164);
nand U1693 (N_1693,In_91,In_620);
nor U1694 (N_1694,In_655,In_132);
or U1695 (N_1695,In_291,In_76);
nor U1696 (N_1696,In_483,In_701);
nor U1697 (N_1697,In_971,In_158);
nor U1698 (N_1698,In_374,In_49);
and U1699 (N_1699,In_585,In_948);
and U1700 (N_1700,In_419,In_554);
nand U1701 (N_1701,In_180,In_843);
nor U1702 (N_1702,In_74,In_848);
or U1703 (N_1703,In_89,In_849);
and U1704 (N_1704,In_204,In_117);
and U1705 (N_1705,In_372,In_552);
nand U1706 (N_1706,In_963,In_916);
nor U1707 (N_1707,In_456,In_496);
and U1708 (N_1708,In_62,In_95);
nand U1709 (N_1709,In_644,In_574);
and U1710 (N_1710,In_280,In_286);
and U1711 (N_1711,In_580,In_416);
nand U1712 (N_1712,In_494,In_580);
nand U1713 (N_1713,In_900,In_350);
nand U1714 (N_1714,In_269,In_8);
or U1715 (N_1715,In_408,In_975);
nor U1716 (N_1716,In_812,In_625);
nand U1717 (N_1717,In_525,In_845);
nor U1718 (N_1718,In_167,In_998);
or U1719 (N_1719,In_386,In_779);
nor U1720 (N_1720,In_50,In_268);
or U1721 (N_1721,In_43,In_260);
or U1722 (N_1722,In_492,In_627);
nor U1723 (N_1723,In_58,In_165);
or U1724 (N_1724,In_14,In_98);
nand U1725 (N_1725,In_181,In_237);
nor U1726 (N_1726,In_385,In_712);
and U1727 (N_1727,In_935,In_691);
nand U1728 (N_1728,In_918,In_38);
nand U1729 (N_1729,In_794,In_739);
and U1730 (N_1730,In_997,In_335);
nor U1731 (N_1731,In_963,In_583);
nor U1732 (N_1732,In_146,In_23);
or U1733 (N_1733,In_430,In_620);
nor U1734 (N_1734,In_979,In_137);
and U1735 (N_1735,In_776,In_627);
nand U1736 (N_1736,In_56,In_898);
nor U1737 (N_1737,In_833,In_19);
and U1738 (N_1738,In_610,In_759);
or U1739 (N_1739,In_106,In_161);
xor U1740 (N_1740,In_359,In_972);
or U1741 (N_1741,In_785,In_809);
nand U1742 (N_1742,In_917,In_708);
nand U1743 (N_1743,In_4,In_502);
nor U1744 (N_1744,In_796,In_681);
and U1745 (N_1745,In_599,In_768);
nand U1746 (N_1746,In_265,In_663);
or U1747 (N_1747,In_32,In_806);
nor U1748 (N_1748,In_392,In_672);
nor U1749 (N_1749,In_766,In_94);
nand U1750 (N_1750,In_749,In_210);
or U1751 (N_1751,In_974,In_290);
or U1752 (N_1752,In_771,In_72);
and U1753 (N_1753,In_744,In_327);
xor U1754 (N_1754,In_288,In_170);
and U1755 (N_1755,In_412,In_540);
nor U1756 (N_1756,In_477,In_547);
or U1757 (N_1757,In_606,In_46);
nor U1758 (N_1758,In_633,In_207);
xor U1759 (N_1759,In_141,In_494);
xor U1760 (N_1760,In_948,In_283);
nor U1761 (N_1761,In_327,In_38);
or U1762 (N_1762,In_205,In_392);
or U1763 (N_1763,In_153,In_419);
and U1764 (N_1764,In_362,In_356);
or U1765 (N_1765,In_887,In_908);
or U1766 (N_1766,In_512,In_83);
nand U1767 (N_1767,In_512,In_922);
nor U1768 (N_1768,In_564,In_694);
and U1769 (N_1769,In_154,In_150);
and U1770 (N_1770,In_309,In_341);
and U1771 (N_1771,In_845,In_623);
and U1772 (N_1772,In_759,In_435);
nor U1773 (N_1773,In_492,In_961);
nand U1774 (N_1774,In_0,In_408);
and U1775 (N_1775,In_410,In_570);
nand U1776 (N_1776,In_961,In_786);
xnor U1777 (N_1777,In_612,In_215);
or U1778 (N_1778,In_420,In_332);
nand U1779 (N_1779,In_910,In_648);
nor U1780 (N_1780,In_916,In_391);
or U1781 (N_1781,In_295,In_575);
and U1782 (N_1782,In_16,In_811);
nor U1783 (N_1783,In_674,In_829);
and U1784 (N_1784,In_381,In_766);
or U1785 (N_1785,In_560,In_518);
and U1786 (N_1786,In_51,In_857);
nand U1787 (N_1787,In_483,In_394);
and U1788 (N_1788,In_442,In_547);
or U1789 (N_1789,In_490,In_740);
nor U1790 (N_1790,In_683,In_762);
or U1791 (N_1791,In_672,In_574);
or U1792 (N_1792,In_980,In_309);
nor U1793 (N_1793,In_250,In_921);
xor U1794 (N_1794,In_640,In_584);
xor U1795 (N_1795,In_601,In_343);
and U1796 (N_1796,In_867,In_754);
or U1797 (N_1797,In_599,In_466);
or U1798 (N_1798,In_125,In_984);
nand U1799 (N_1799,In_976,In_926);
or U1800 (N_1800,In_588,In_704);
or U1801 (N_1801,In_527,In_338);
xnor U1802 (N_1802,In_878,In_372);
nand U1803 (N_1803,In_305,In_692);
or U1804 (N_1804,In_359,In_353);
nand U1805 (N_1805,In_466,In_561);
and U1806 (N_1806,In_770,In_891);
nor U1807 (N_1807,In_933,In_696);
xor U1808 (N_1808,In_233,In_811);
nor U1809 (N_1809,In_606,In_637);
and U1810 (N_1810,In_494,In_289);
nor U1811 (N_1811,In_49,In_337);
or U1812 (N_1812,In_144,In_677);
and U1813 (N_1813,In_84,In_611);
nand U1814 (N_1814,In_888,In_645);
xnor U1815 (N_1815,In_242,In_897);
and U1816 (N_1816,In_730,In_411);
or U1817 (N_1817,In_188,In_463);
nand U1818 (N_1818,In_850,In_480);
nand U1819 (N_1819,In_703,In_928);
nand U1820 (N_1820,In_715,In_400);
or U1821 (N_1821,In_803,In_340);
and U1822 (N_1822,In_892,In_658);
nor U1823 (N_1823,In_453,In_922);
nand U1824 (N_1824,In_626,In_116);
or U1825 (N_1825,In_406,In_248);
xor U1826 (N_1826,In_648,In_274);
nand U1827 (N_1827,In_935,In_141);
or U1828 (N_1828,In_132,In_213);
and U1829 (N_1829,In_719,In_821);
nand U1830 (N_1830,In_5,In_307);
nor U1831 (N_1831,In_666,In_767);
nor U1832 (N_1832,In_580,In_921);
nand U1833 (N_1833,In_692,In_412);
or U1834 (N_1834,In_996,In_227);
nand U1835 (N_1835,In_818,In_372);
or U1836 (N_1836,In_303,In_590);
or U1837 (N_1837,In_552,In_240);
or U1838 (N_1838,In_307,In_88);
xnor U1839 (N_1839,In_530,In_76);
or U1840 (N_1840,In_447,In_278);
nor U1841 (N_1841,In_658,In_520);
nand U1842 (N_1842,In_368,In_163);
and U1843 (N_1843,In_326,In_304);
nor U1844 (N_1844,In_277,In_586);
nor U1845 (N_1845,In_834,In_479);
nor U1846 (N_1846,In_516,In_990);
nand U1847 (N_1847,In_70,In_178);
nand U1848 (N_1848,In_137,In_181);
and U1849 (N_1849,In_386,In_431);
nand U1850 (N_1850,In_591,In_753);
and U1851 (N_1851,In_347,In_662);
nor U1852 (N_1852,In_413,In_84);
and U1853 (N_1853,In_445,In_675);
and U1854 (N_1854,In_643,In_166);
and U1855 (N_1855,In_813,In_255);
nand U1856 (N_1856,In_512,In_393);
nand U1857 (N_1857,In_243,In_313);
and U1858 (N_1858,In_257,In_58);
nor U1859 (N_1859,In_889,In_116);
or U1860 (N_1860,In_365,In_573);
or U1861 (N_1861,In_922,In_832);
xor U1862 (N_1862,In_779,In_41);
nor U1863 (N_1863,In_185,In_413);
or U1864 (N_1864,In_48,In_170);
nand U1865 (N_1865,In_87,In_414);
or U1866 (N_1866,In_541,In_565);
nand U1867 (N_1867,In_373,In_608);
and U1868 (N_1868,In_893,In_131);
nand U1869 (N_1869,In_132,In_423);
nand U1870 (N_1870,In_163,In_461);
or U1871 (N_1871,In_987,In_95);
and U1872 (N_1872,In_551,In_358);
nand U1873 (N_1873,In_604,In_668);
xor U1874 (N_1874,In_23,In_145);
nand U1875 (N_1875,In_853,In_294);
nand U1876 (N_1876,In_284,In_722);
and U1877 (N_1877,In_120,In_817);
nand U1878 (N_1878,In_752,In_17);
nand U1879 (N_1879,In_586,In_998);
nor U1880 (N_1880,In_16,In_119);
and U1881 (N_1881,In_905,In_523);
or U1882 (N_1882,In_535,In_938);
or U1883 (N_1883,In_702,In_350);
or U1884 (N_1884,In_316,In_97);
nand U1885 (N_1885,In_528,In_397);
nor U1886 (N_1886,In_977,In_718);
nor U1887 (N_1887,In_870,In_923);
xnor U1888 (N_1888,In_153,In_683);
nand U1889 (N_1889,In_348,In_380);
nand U1890 (N_1890,In_442,In_400);
or U1891 (N_1891,In_135,In_534);
nand U1892 (N_1892,In_213,In_708);
nor U1893 (N_1893,In_228,In_309);
nand U1894 (N_1894,In_312,In_122);
or U1895 (N_1895,In_336,In_70);
xor U1896 (N_1896,In_945,In_749);
xor U1897 (N_1897,In_285,In_74);
or U1898 (N_1898,In_747,In_159);
and U1899 (N_1899,In_646,In_268);
nor U1900 (N_1900,In_892,In_473);
nor U1901 (N_1901,In_195,In_167);
and U1902 (N_1902,In_764,In_136);
nor U1903 (N_1903,In_672,In_603);
or U1904 (N_1904,In_998,In_871);
nor U1905 (N_1905,In_218,In_550);
xnor U1906 (N_1906,In_235,In_343);
and U1907 (N_1907,In_464,In_596);
and U1908 (N_1908,In_348,In_962);
nor U1909 (N_1909,In_905,In_768);
and U1910 (N_1910,In_80,In_202);
and U1911 (N_1911,In_69,In_478);
or U1912 (N_1912,In_763,In_803);
nor U1913 (N_1913,In_434,In_106);
xor U1914 (N_1914,In_568,In_683);
xor U1915 (N_1915,In_933,In_137);
nand U1916 (N_1916,In_314,In_776);
nor U1917 (N_1917,In_711,In_219);
nand U1918 (N_1918,In_725,In_544);
nor U1919 (N_1919,In_629,In_192);
xnor U1920 (N_1920,In_784,In_219);
nor U1921 (N_1921,In_826,In_204);
or U1922 (N_1922,In_297,In_284);
nor U1923 (N_1923,In_863,In_213);
and U1924 (N_1924,In_787,In_732);
or U1925 (N_1925,In_78,In_46);
nor U1926 (N_1926,In_196,In_890);
and U1927 (N_1927,In_207,In_985);
xnor U1928 (N_1928,In_520,In_330);
or U1929 (N_1929,In_103,In_747);
and U1930 (N_1930,In_238,In_160);
and U1931 (N_1931,In_921,In_894);
nand U1932 (N_1932,In_332,In_707);
nor U1933 (N_1933,In_908,In_730);
or U1934 (N_1934,In_11,In_411);
nor U1935 (N_1935,In_959,In_306);
or U1936 (N_1936,In_756,In_502);
and U1937 (N_1937,In_242,In_312);
or U1938 (N_1938,In_589,In_997);
nand U1939 (N_1939,In_520,In_864);
or U1940 (N_1940,In_57,In_850);
and U1941 (N_1941,In_42,In_379);
or U1942 (N_1942,In_798,In_881);
nand U1943 (N_1943,In_445,In_608);
nor U1944 (N_1944,In_145,In_382);
or U1945 (N_1945,In_847,In_253);
or U1946 (N_1946,In_996,In_169);
nor U1947 (N_1947,In_921,In_115);
nand U1948 (N_1948,In_970,In_353);
or U1949 (N_1949,In_448,In_619);
or U1950 (N_1950,In_150,In_4);
or U1951 (N_1951,In_35,In_175);
nor U1952 (N_1952,In_74,In_644);
or U1953 (N_1953,In_705,In_992);
nor U1954 (N_1954,In_579,In_178);
and U1955 (N_1955,In_106,In_758);
nand U1956 (N_1956,In_851,In_554);
or U1957 (N_1957,In_255,In_408);
nor U1958 (N_1958,In_487,In_446);
nand U1959 (N_1959,In_77,In_0);
or U1960 (N_1960,In_789,In_211);
nand U1961 (N_1961,In_873,In_888);
and U1962 (N_1962,In_720,In_209);
nand U1963 (N_1963,In_329,In_568);
and U1964 (N_1964,In_784,In_864);
or U1965 (N_1965,In_163,In_796);
and U1966 (N_1966,In_813,In_354);
nor U1967 (N_1967,In_351,In_324);
or U1968 (N_1968,In_977,In_848);
nor U1969 (N_1969,In_886,In_487);
or U1970 (N_1970,In_622,In_9);
nand U1971 (N_1971,In_582,In_547);
and U1972 (N_1972,In_573,In_282);
nor U1973 (N_1973,In_847,In_263);
xor U1974 (N_1974,In_945,In_573);
and U1975 (N_1975,In_330,In_375);
nand U1976 (N_1976,In_827,In_418);
nand U1977 (N_1977,In_65,In_764);
or U1978 (N_1978,In_934,In_147);
nor U1979 (N_1979,In_14,In_759);
nor U1980 (N_1980,In_238,In_337);
nand U1981 (N_1981,In_70,In_261);
nor U1982 (N_1982,In_876,In_726);
and U1983 (N_1983,In_95,In_301);
or U1984 (N_1984,In_860,In_747);
or U1985 (N_1985,In_873,In_127);
nand U1986 (N_1986,In_4,In_179);
or U1987 (N_1987,In_279,In_290);
nand U1988 (N_1988,In_557,In_122);
nor U1989 (N_1989,In_320,In_827);
and U1990 (N_1990,In_827,In_319);
nand U1991 (N_1991,In_683,In_475);
or U1992 (N_1992,In_944,In_541);
nor U1993 (N_1993,In_99,In_272);
nand U1994 (N_1994,In_625,In_871);
and U1995 (N_1995,In_177,In_223);
and U1996 (N_1996,In_695,In_465);
nor U1997 (N_1997,In_776,In_124);
nor U1998 (N_1998,In_824,In_120);
nand U1999 (N_1999,In_170,In_707);
xor U2000 (N_2000,N_938,N_1522);
and U2001 (N_2001,N_869,N_1626);
and U2002 (N_2002,N_926,N_1964);
xor U2003 (N_2003,N_1351,N_581);
xnor U2004 (N_2004,N_107,N_444);
and U2005 (N_2005,N_597,N_1142);
nor U2006 (N_2006,N_93,N_474);
and U2007 (N_2007,N_1380,N_775);
and U2008 (N_2008,N_1776,N_1105);
and U2009 (N_2009,N_913,N_1622);
and U2010 (N_2010,N_1940,N_545);
nor U2011 (N_2011,N_1917,N_864);
nor U2012 (N_2012,N_1901,N_1580);
or U2013 (N_2013,N_219,N_615);
and U2014 (N_2014,N_1437,N_164);
nor U2015 (N_2015,N_1914,N_376);
xnor U2016 (N_2016,N_1609,N_524);
nand U2017 (N_2017,N_690,N_1500);
nor U2018 (N_2018,N_147,N_807);
nand U2019 (N_2019,N_240,N_361);
nor U2020 (N_2020,N_1002,N_553);
xor U2021 (N_2021,N_290,N_539);
and U2022 (N_2022,N_1990,N_1100);
and U2023 (N_2023,N_908,N_1666);
nand U2024 (N_2024,N_1853,N_15);
nand U2025 (N_2025,N_1548,N_985);
nor U2026 (N_2026,N_99,N_1256);
or U2027 (N_2027,N_892,N_1905);
and U2028 (N_2028,N_1126,N_69);
and U2029 (N_2029,N_1368,N_3);
xnor U2030 (N_2030,N_664,N_243);
and U2031 (N_2031,N_962,N_1504);
xor U2032 (N_2032,N_1510,N_1751);
nor U2033 (N_2033,N_1306,N_114);
nor U2034 (N_2034,N_883,N_1341);
xor U2035 (N_2035,N_188,N_56);
or U2036 (N_2036,N_673,N_1801);
nand U2037 (N_2037,N_1922,N_126);
xor U2038 (N_2038,N_1319,N_874);
or U2039 (N_2039,N_591,N_1070);
nor U2040 (N_2040,N_1201,N_412);
xnor U2041 (N_2041,N_1680,N_856);
xor U2042 (N_2042,N_1684,N_1952);
and U2043 (N_2043,N_1307,N_1218);
and U2044 (N_2044,N_1779,N_1619);
and U2045 (N_2045,N_1902,N_1975);
nand U2046 (N_2046,N_385,N_1452);
nor U2047 (N_2047,N_478,N_1515);
nand U2048 (N_2048,N_1178,N_1007);
or U2049 (N_2049,N_50,N_1832);
and U2050 (N_2050,N_1967,N_55);
nand U2051 (N_2051,N_1140,N_1054);
nand U2052 (N_2052,N_975,N_1294);
nand U2053 (N_2053,N_277,N_564);
nor U2054 (N_2054,N_101,N_369);
nor U2055 (N_2055,N_537,N_781);
nand U2056 (N_2056,N_1644,N_1222);
nand U2057 (N_2057,N_245,N_843);
and U2058 (N_2058,N_1577,N_1998);
or U2059 (N_2059,N_991,N_170);
nor U2060 (N_2060,N_464,N_161);
nor U2061 (N_2061,N_1717,N_1014);
and U2062 (N_2062,N_1193,N_1027);
or U2063 (N_2063,N_401,N_432);
and U2064 (N_2064,N_1327,N_259);
nor U2065 (N_2065,N_530,N_496);
or U2066 (N_2066,N_1291,N_275);
nor U2067 (N_2067,N_197,N_642);
nand U2068 (N_2068,N_1004,N_1093);
nand U2069 (N_2069,N_779,N_386);
or U2070 (N_2070,N_1470,N_185);
xor U2071 (N_2071,N_291,N_1512);
and U2072 (N_2072,N_945,N_839);
or U2073 (N_2073,N_1524,N_1486);
or U2074 (N_2074,N_1325,N_1314);
nand U2075 (N_2075,N_1558,N_77);
nor U2076 (N_2076,N_98,N_1814);
nand U2077 (N_2077,N_1671,N_454);
and U2078 (N_2078,N_1395,N_1704);
and U2079 (N_2079,N_1163,N_980);
nor U2080 (N_2080,N_1273,N_878);
nand U2081 (N_2081,N_492,N_441);
nand U2082 (N_2082,N_611,N_175);
nand U2083 (N_2083,N_284,N_999);
nand U2084 (N_2084,N_208,N_381);
or U2085 (N_2085,N_907,N_557);
xnor U2086 (N_2086,N_254,N_1980);
nand U2087 (N_2087,N_313,N_1710);
xnor U2088 (N_2088,N_1048,N_1157);
nand U2089 (N_2089,N_1979,N_967);
or U2090 (N_2090,N_933,N_439);
xnor U2091 (N_2091,N_155,N_1383);
and U2092 (N_2092,N_1816,N_260);
or U2093 (N_2093,N_42,N_505);
nor U2094 (N_2094,N_176,N_647);
nor U2095 (N_2095,N_605,N_124);
nand U2096 (N_2096,N_1421,N_61);
or U2097 (N_2097,N_1931,N_1603);
or U2098 (N_2098,N_1764,N_1670);
or U2099 (N_2099,N_1389,N_1090);
nor U2100 (N_2100,N_1624,N_1542);
and U2101 (N_2101,N_1363,N_1232);
nand U2102 (N_2102,N_650,N_1336);
nor U2103 (N_2103,N_763,N_1274);
xnor U2104 (N_2104,N_1230,N_1258);
xor U2105 (N_2105,N_1555,N_927);
xnor U2106 (N_2106,N_22,N_136);
nand U2107 (N_2107,N_1191,N_267);
nand U2108 (N_2108,N_630,N_901);
or U2109 (N_2109,N_418,N_483);
nor U2110 (N_2110,N_702,N_6);
nor U2111 (N_2111,N_696,N_726);
and U2112 (N_2112,N_893,N_1691);
nor U2113 (N_2113,N_1071,N_1834);
and U2114 (N_2114,N_1244,N_223);
nor U2115 (N_2115,N_787,N_421);
nand U2116 (N_2116,N_1849,N_1117);
and U2117 (N_2117,N_1777,N_1183);
and U2118 (N_2118,N_954,N_1479);
or U2119 (N_2119,N_1811,N_470);
and U2120 (N_2120,N_210,N_1173);
or U2121 (N_2121,N_1873,N_1496);
nor U2122 (N_2122,N_1487,N_1761);
nor U2123 (N_2123,N_1049,N_881);
and U2124 (N_2124,N_1502,N_1094);
or U2125 (N_2125,N_863,N_287);
and U2126 (N_2126,N_1259,N_187);
and U2127 (N_2127,N_1360,N_773);
nand U2128 (N_2128,N_1417,N_1628);
or U2129 (N_2129,N_1883,N_1392);
nand U2130 (N_2130,N_449,N_366);
nor U2131 (N_2131,N_1313,N_1428);
and U2132 (N_2132,N_1694,N_472);
nand U2133 (N_2133,N_1768,N_959);
or U2134 (N_2134,N_1974,N_251);
nor U2135 (N_2135,N_18,N_1983);
and U2136 (N_2136,N_1842,N_709);
nand U2137 (N_2137,N_1771,N_915);
or U2138 (N_2138,N_1175,N_555);
nand U2139 (N_2139,N_728,N_1495);
xnor U2140 (N_2140,N_744,N_675);
and U2141 (N_2141,N_390,N_105);
nor U2142 (N_2142,N_1848,N_1077);
or U2143 (N_2143,N_289,N_937);
nor U2144 (N_2144,N_1404,N_522);
nor U2145 (N_2145,N_1455,N_956);
nand U2146 (N_2146,N_1858,N_95);
and U2147 (N_2147,N_34,N_297);
and U2148 (N_2148,N_1583,N_1478);
nand U2149 (N_2149,N_1135,N_867);
or U2150 (N_2150,N_1016,N_784);
and U2151 (N_2151,N_1330,N_1593);
nor U2152 (N_2152,N_976,N_1910);
nand U2153 (N_2153,N_765,N_508);
or U2154 (N_2154,N_1119,N_894);
or U2155 (N_2155,N_868,N_94);
and U2156 (N_2156,N_565,N_182);
nand U2157 (N_2157,N_1614,N_1145);
nand U2158 (N_2158,N_1243,N_579);
and U2159 (N_2159,N_792,N_1571);
and U2160 (N_2160,N_1878,N_1862);
or U2161 (N_2161,N_1997,N_405);
xnor U2162 (N_2162,N_1630,N_1869);
and U2163 (N_2163,N_1774,N_1652);
nand U2164 (N_2164,N_710,N_1097);
nor U2165 (N_2165,N_1362,N_48);
xor U2166 (N_2166,N_317,N_355);
or U2167 (N_2167,N_139,N_311);
and U2168 (N_2168,N_104,N_1210);
nor U2169 (N_2169,N_875,N_809);
and U2170 (N_2170,N_1015,N_1525);
and U2171 (N_2171,N_337,N_1889);
and U2172 (N_2172,N_207,N_1466);
and U2173 (N_2173,N_1503,N_944);
and U2174 (N_2174,N_1633,N_1023);
nor U2175 (N_2175,N_1800,N_1326);
nand U2176 (N_2176,N_580,N_1084);
xor U2177 (N_2177,N_1066,N_1059);
or U2178 (N_2178,N_1456,N_523);
or U2179 (N_2179,N_26,N_700);
nor U2180 (N_2180,N_1535,N_745);
nor U2181 (N_2181,N_1903,N_145);
and U2182 (N_2182,N_1859,N_1067);
and U2183 (N_2183,N_1445,N_1198);
xnor U2184 (N_2184,N_183,N_1591);
nor U2185 (N_2185,N_435,N_320);
or U2186 (N_2186,N_1870,N_391);
nand U2187 (N_2187,N_72,N_733);
nor U2188 (N_2188,N_641,N_742);
nor U2189 (N_2189,N_1890,N_613);
xnor U2190 (N_2190,N_1984,N_886);
or U2191 (N_2191,N_903,N_739);
or U2192 (N_2192,N_1220,N_683);
nor U2193 (N_2193,N_1449,N_1053);
xnor U2194 (N_2194,N_998,N_1925);
nand U2195 (N_2195,N_129,N_1891);
nor U2196 (N_2196,N_870,N_417);
and U2197 (N_2197,N_65,N_905);
or U2198 (N_2198,N_1523,N_1594);
and U2199 (N_2199,N_1729,N_237);
and U2200 (N_2200,N_443,N_1034);
nor U2201 (N_2201,N_968,N_339);
xnor U2202 (N_2202,N_46,N_764);
and U2203 (N_2203,N_84,N_626);
and U2204 (N_2204,N_1242,N_670);
nor U2205 (N_2205,N_704,N_1480);
nor U2206 (N_2206,N_137,N_1755);
nand U2207 (N_2207,N_1909,N_1010);
nor U2208 (N_2208,N_1440,N_1130);
xor U2209 (N_2209,N_1753,N_1513);
or U2210 (N_2210,N_794,N_1699);
and U2211 (N_2211,N_828,N_1020);
and U2212 (N_2212,N_1118,N_1683);
nor U2213 (N_2213,N_218,N_1397);
nand U2214 (N_2214,N_285,N_268);
or U2215 (N_2215,N_1200,N_399);
and U2216 (N_2216,N_1492,N_900);
nand U2217 (N_2217,N_1531,N_1528);
xnor U2218 (N_2218,N_785,N_526);
nor U2219 (N_2219,N_1822,N_184);
and U2220 (N_2220,N_1155,N_648);
xnor U2221 (N_2221,N_1018,N_177);
or U2222 (N_2222,N_460,N_1752);
nor U2223 (N_2223,N_592,N_1038);
nand U2224 (N_2224,N_1186,N_1866);
or U2225 (N_2225,N_606,N_952);
nand U2226 (N_2226,N_762,N_1969);
nand U2227 (N_2227,N_1340,N_769);
nor U2228 (N_2228,N_1672,N_821);
nor U2229 (N_2229,N_947,N_20);
xor U2230 (N_2230,N_1098,N_378);
nor U2231 (N_2231,N_1782,N_1374);
xor U2232 (N_2232,N_639,N_1621);
xor U2233 (N_2233,N_1876,N_1673);
nand U2234 (N_2234,N_1199,N_1475);
nand U2235 (N_2235,N_1977,N_1095);
xor U2236 (N_2236,N_1387,N_1143);
nor U2237 (N_2237,N_1391,N_583);
xor U2238 (N_2238,N_877,N_1134);
nand U2239 (N_2239,N_117,N_315);
or U2240 (N_2240,N_1563,N_1216);
nand U2241 (N_2241,N_940,N_1951);
or U2242 (N_2242,N_970,N_64);
or U2243 (N_2243,N_1564,N_961);
and U2244 (N_2244,N_1530,N_1572);
or U2245 (N_2245,N_271,N_157);
and U2246 (N_2246,N_142,N_981);
nor U2247 (N_2247,N_1506,N_1716);
nand U2248 (N_2248,N_1260,N_574);
and U2249 (N_2249,N_1120,N_485);
and U2250 (N_2250,N_1723,N_389);
nand U2251 (N_2251,N_844,N_1806);
and U2252 (N_2252,N_63,N_517);
or U2253 (N_2253,N_992,N_236);
and U2254 (N_2254,N_358,N_249);
xor U2255 (N_2255,N_788,N_1802);
nand U2256 (N_2256,N_91,N_616);
or U2257 (N_2257,N_1152,N_1176);
and U2258 (N_2258,N_322,N_860);
or U2259 (N_2259,N_708,N_397);
xnor U2260 (N_2260,N_603,N_1103);
nor U2261 (N_2261,N_582,N_1182);
and U2262 (N_2262,N_73,N_578);
or U2263 (N_2263,N_1133,N_1714);
and U2264 (N_2264,N_487,N_1843);
nor U2265 (N_2265,N_1436,N_1857);
nor U2266 (N_2266,N_621,N_1649);
or U2267 (N_2267,N_644,N_1308);
and U2268 (N_2268,N_1278,N_1426);
or U2269 (N_2269,N_608,N_836);
nor U2270 (N_2270,N_459,N_1044);
and U2271 (N_2271,N_1003,N_832);
or U2272 (N_2272,N_774,N_215);
nor U2273 (N_2273,N_547,N_720);
and U2274 (N_2274,N_1772,N_1992);
and U2275 (N_2275,N_786,N_620);
nand U2276 (N_2276,N_80,N_425);
nand U2277 (N_2277,N_1676,N_1312);
or U2278 (N_2278,N_1927,N_1116);
nor U2279 (N_2279,N_576,N_1787);
nor U2280 (N_2280,N_1301,N_248);
xor U2281 (N_2281,N_989,N_910);
or U2282 (N_2282,N_224,N_1352);
nand U2283 (N_2283,N_14,N_51);
or U2284 (N_2284,N_402,N_543);
nor U2285 (N_2285,N_1433,N_1179);
and U2286 (N_2286,N_1401,N_423);
or U2287 (N_2287,N_1646,N_1557);
or U2288 (N_2288,N_1618,N_1290);
nor U2289 (N_2289,N_1447,N_1907);
nand U2290 (N_2290,N_588,N_292);
or U2291 (N_2291,N_1544,N_632);
and U2292 (N_2292,N_178,N_1737);
nor U2293 (N_2293,N_1211,N_780);
nand U2294 (N_2294,N_1289,N_1375);
and U2295 (N_2295,N_727,N_717);
xnor U2296 (N_2296,N_1919,N_1300);
or U2297 (N_2297,N_738,N_855);
xnor U2298 (N_2298,N_1386,N_1229);
nand U2299 (N_2299,N_1149,N_1129);
or U2300 (N_2300,N_1584,N_1272);
and U2301 (N_2301,N_367,N_1598);
and U2302 (N_2302,N_13,N_885);
and U2303 (N_2303,N_468,N_1678);
or U2304 (N_2304,N_997,N_891);
or U2305 (N_2305,N_946,N_1904);
or U2306 (N_2306,N_1682,N_1473);
nor U2307 (N_2307,N_923,N_1420);
nand U2308 (N_2308,N_1617,N_33);
and U2309 (N_2309,N_206,N_607);
or U2310 (N_2310,N_234,N_1139);
or U2311 (N_2311,N_1187,N_808);
and U2312 (N_2312,N_1600,N_1819);
or U2313 (N_2313,N_590,N_1110);
and U2314 (N_2314,N_1916,N_345);
nand U2315 (N_2315,N_1713,N_1477);
nor U2316 (N_2316,N_1681,N_481);
nor U2317 (N_2317,N_988,N_1575);
and U2318 (N_2318,N_408,N_887);
nor U2319 (N_2319,N_192,N_1322);
xor U2320 (N_2320,N_1329,N_186);
nand U2321 (N_2321,N_1342,N_228);
nand U2322 (N_2322,N_1263,N_293);
and U2323 (N_2323,N_637,N_711);
nand U2324 (N_2324,N_698,N_450);
or U2325 (N_2325,N_445,N_1749);
or U2326 (N_2326,N_1275,N_40);
nor U2327 (N_2327,N_798,N_463);
nor U2328 (N_2328,N_571,N_1978);
nand U2329 (N_2329,N_81,N_174);
or U2330 (N_2330,N_1605,N_370);
nor U2331 (N_2331,N_1852,N_643);
or U2332 (N_2332,N_1061,N_1269);
nor U2333 (N_2333,N_419,N_199);
and U2334 (N_2334,N_1485,N_1039);
nor U2335 (N_2335,N_1921,N_382);
and U2336 (N_2336,N_318,N_667);
nor U2337 (N_2337,N_150,N_495);
or U2338 (N_2338,N_825,N_1727);
or U2339 (N_2339,N_422,N_1724);
nor U2340 (N_2340,N_306,N_1611);
and U2341 (N_2341,N_1788,N_39);
and U2342 (N_2342,N_71,N_519);
nor U2343 (N_2343,N_1136,N_707);
nand U2344 (N_2344,N_1585,N_1606);
nor U2345 (N_2345,N_761,N_209);
or U2346 (N_2346,N_1830,N_802);
xor U2347 (N_2347,N_1223,N_740);
and U2348 (N_2348,N_309,N_890);
or U2349 (N_2349,N_851,N_1196);
and U2350 (N_2350,N_627,N_1730);
nor U2351 (N_2351,N_1913,N_235);
or U2352 (N_2352,N_214,N_1692);
or U2353 (N_2353,N_803,N_1385);
or U2354 (N_2354,N_1958,N_593);
nand U2355 (N_2355,N_1250,N_41);
or U2356 (N_2356,N_755,N_820);
or U2357 (N_2357,N_1028,N_873);
nand U2358 (N_2358,N_1328,N_872);
xnor U2359 (N_2359,N_958,N_1868);
and U2360 (N_2360,N_1482,N_895);
and U2361 (N_2361,N_1252,N_252);
nand U2362 (N_2362,N_840,N_159);
nor U2363 (N_2363,N_68,N_655);
nand U2364 (N_2364,N_1035,N_1740);
nor U2365 (N_2365,N_973,N_685);
nor U2366 (N_2366,N_969,N_200);
nor U2367 (N_2367,N_167,N_943);
nand U2368 (N_2368,N_1156,N_1347);
and U2369 (N_2369,N_244,N_680);
and U2370 (N_2370,N_1659,N_1172);
nand U2371 (N_2371,N_1655,N_1180);
or U2372 (N_2372,N_1316,N_49);
and U2373 (N_2373,N_1219,N_471);
or U2374 (N_2374,N_796,N_96);
or U2375 (N_2375,N_1108,N_888);
nor U2376 (N_2376,N_230,N_279);
or U2377 (N_2377,N_1726,N_541);
and U2378 (N_2378,N_377,N_1928);
nand U2379 (N_2379,N_350,N_1851);
xor U2380 (N_2380,N_684,N_1005);
nand U2381 (N_2381,N_584,N_609);
or U2382 (N_2382,N_1826,N_846);
or U2383 (N_2383,N_1864,N_269);
and U2384 (N_2384,N_1497,N_272);
and U2385 (N_2385,N_1770,N_749);
and U2386 (N_2386,N_323,N_1359);
xor U2387 (N_2387,N_817,N_1378);
nor U2388 (N_2388,N_1871,N_1062);
nor U2389 (N_2389,N_1001,N_1960);
or U2390 (N_2390,N_1656,N_1254);
or U2391 (N_2391,N_1642,N_1657);
nor U2392 (N_2392,N_1321,N_1547);
xnor U2393 (N_2393,N_633,N_879);
and U2394 (N_2394,N_1817,N_1450);
and U2395 (N_2395,N_841,N_876);
and U2396 (N_2396,N_924,N_697);
xnor U2397 (N_2397,N_149,N_1267);
nor U2398 (N_2398,N_17,N_127);
or U2399 (N_2399,N_1625,N_1698);
or U2400 (N_2400,N_1950,N_79);
and U2401 (N_2401,N_1171,N_420);
nor U2402 (N_2402,N_978,N_1879);
xnor U2403 (N_2403,N_131,N_1912);
and U2404 (N_2404,N_53,N_861);
nor U2405 (N_2405,N_1367,N_356);
nor U2406 (N_2406,N_392,N_1246);
nand U2407 (N_2407,N_70,N_1343);
nor U2408 (N_2408,N_987,N_1778);
nand U2409 (N_2409,N_516,N_1356);
or U2410 (N_2410,N_5,N_518);
xor U2411 (N_2411,N_651,N_1836);
and U2412 (N_2412,N_1856,N_737);
nor U2413 (N_2413,N_1235,N_1797);
and U2414 (N_2414,N_407,N_437);
or U2415 (N_2415,N_455,N_1460);
or U2416 (N_2416,N_343,N_715);
nand U2417 (N_2417,N_1651,N_1861);
nand U2418 (N_2418,N_949,N_484);
nand U2419 (N_2419,N_1712,N_1215);
or U2420 (N_2420,N_815,N_857);
or U2421 (N_2421,N_1932,N_829);
and U2422 (N_2422,N_212,N_270);
nand U2423 (N_2423,N_457,N_920);
and U2424 (N_2424,N_1590,N_520);
nand U2425 (N_2425,N_1111,N_1058);
nor U2426 (N_2426,N_357,N_1277);
and U2427 (N_2427,N_213,N_1635);
nor U2428 (N_2428,N_1760,N_406);
xor U2429 (N_2429,N_1794,N_566);
or U2430 (N_2430,N_993,N_1151);
and U2431 (N_2431,N_398,N_301);
xnor U2432 (N_2432,N_990,N_1501);
or U2433 (N_2433,N_1364,N_957);
nor U2434 (N_2434,N_1505,N_1442);
or U2435 (N_2435,N_173,N_859);
xor U2436 (N_2436,N_222,N_1376);
nor U2437 (N_2437,N_181,N_546);
xnor U2438 (N_2438,N_466,N_953);
and U2439 (N_2439,N_160,N_835);
and U2440 (N_2440,N_882,N_563);
or U2441 (N_2441,N_672,N_941);
xnor U2442 (N_2442,N_85,N_100);
nand U2443 (N_2443,N_1262,N_16);
xnor U2444 (N_2444,N_1446,N_1773);
nor U2445 (N_2445,N_734,N_1435);
and U2446 (N_2446,N_1805,N_329);
nand U2447 (N_2447,N_1177,N_8);
nand U2448 (N_2448,N_1037,N_865);
or U2449 (N_2449,N_1551,N_917);
xnor U2450 (N_2450,N_1884,N_701);
or U2451 (N_2451,N_344,N_1780);
nor U2452 (N_2452,N_805,N_128);
or U2453 (N_2453,N_1996,N_795);
or U2454 (N_2454,N_1241,N_548);
nand U2455 (N_2455,N_262,N_884);
nor U2456 (N_2456,N_1754,N_1169);
nor U2457 (N_2457,N_556,N_1721);
nor U2458 (N_2458,N_1334,N_1715);
and U2459 (N_2459,N_1693,N_87);
and U2460 (N_2460,N_1346,N_1205);
xnor U2461 (N_2461,N_661,N_1285);
nor U2462 (N_2462,N_812,N_335);
or U2463 (N_2463,N_671,N_1102);
or U2464 (N_2464,N_964,N_451);
xnor U2465 (N_2465,N_1029,N_1231);
xnor U2466 (N_2466,N_1379,N_1520);
and U2467 (N_2467,N_148,N_1315);
xnor U2468 (N_2468,N_965,N_304);
and U2469 (N_2469,N_1578,N_1454);
and U2470 (N_2470,N_111,N_121);
nor U2471 (N_2471,N_902,N_653);
and U2472 (N_2472,N_333,N_814);
nor U2473 (N_2473,N_1565,N_845);
or U2474 (N_2474,N_30,N_372);
or U2475 (N_2475,N_1875,N_1534);
nor U2476 (N_2476,N_1769,N_612);
and U2477 (N_2477,N_1045,N_1517);
nor U2478 (N_2478,N_1465,N_1377);
nand U2479 (N_2479,N_629,N_1763);
or U2480 (N_2480,N_1813,N_904);
and U2481 (N_2481,N_486,N_365);
and U2482 (N_2482,N_1365,N_247);
and U2483 (N_2483,N_1798,N_1137);
nor U2484 (N_2484,N_799,N_1677);
nor U2485 (N_2485,N_1224,N_1011);
and U2486 (N_2486,N_654,N_404);
nand U2487 (N_2487,N_501,N_1170);
or U2488 (N_2488,N_1481,N_1213);
and U2489 (N_2489,N_427,N_929);
and U2490 (N_2490,N_433,N_1664);
and U2491 (N_2491,N_165,N_816);
nor U2492 (N_2492,N_67,N_1867);
or U2493 (N_2493,N_32,N_666);
nor U2494 (N_2494,N_102,N_1488);
or U2495 (N_2495,N_1393,N_225);
nor U2496 (N_2496,N_898,N_1238);
nor U2497 (N_2497,N_760,N_716);
or U2498 (N_2498,N_138,N_595);
nor U2499 (N_2499,N_528,N_103);
nand U2500 (N_2500,N_1491,N_682);
and U2501 (N_2501,N_11,N_1138);
nand U2502 (N_2502,N_669,N_925);
or U2503 (N_2503,N_772,N_1537);
nor U2504 (N_2504,N_1767,N_677);
nand U2505 (N_2505,N_1731,N_371);
xnor U2506 (N_2506,N_205,N_1150);
and U2507 (N_2507,N_587,N_656);
and U2508 (N_2508,N_273,N_411);
or U2509 (N_2509,N_1561,N_153);
xor U2510 (N_2510,N_1926,N_303);
nand U2511 (N_2511,N_179,N_233);
nand U2512 (N_2512,N_1665,N_1493);
and U2513 (N_2513,N_573,N_1918);
or U2514 (N_2514,N_1793,N_135);
nand U2515 (N_2515,N_848,N_782);
and U2516 (N_2516,N_753,N_45);
nor U2517 (N_2517,N_112,N_211);
nand U2518 (N_2518,N_1350,N_527);
or U2519 (N_2519,N_1089,N_1920);
or U2520 (N_2520,N_108,N_1299);
or U2521 (N_2521,N_1128,N_1214);
or U2522 (N_2522,N_241,N_899);
or U2523 (N_2523,N_1893,N_931);
xor U2524 (N_2524,N_379,N_1886);
xor U2525 (N_2525,N_1845,N_2);
or U2526 (N_2526,N_456,N_189);
nand U2527 (N_2527,N_1144,N_364);
or U2528 (N_2528,N_752,N_842);
nand U2529 (N_2529,N_1679,N_1756);
or U2530 (N_2530,N_1934,N_434);
nor U2531 (N_2531,N_1463,N_4);
xnor U2532 (N_2532,N_797,N_741);
xnor U2533 (N_2533,N_826,N_1438);
nand U2534 (N_2534,N_1911,N_996);
and U2535 (N_2535,N_266,N_963);
nand U2536 (N_2536,N_1131,N_1168);
nor U2537 (N_2537,N_1616,N_1711);
nor U2538 (N_2538,N_1947,N_134);
and U2539 (N_2539,N_1532,N_889);
or U2540 (N_2540,N_1837,N_1707);
and U2541 (N_2541,N_28,N_146);
and U2542 (N_2542,N_568,N_1212);
or U2543 (N_2543,N_1448,N_930);
nor U2544 (N_2544,N_635,N_368);
nor U2545 (N_2545,N_1645,N_724);
nor U2546 (N_2546,N_257,N_1400);
nand U2547 (N_2547,N_1153,N_436);
and U2548 (N_2548,N_995,N_854);
nand U2549 (N_2549,N_1750,N_47);
or U2550 (N_2550,N_1441,N_935);
nor U2551 (N_2551,N_1271,N_1647);
or U2552 (N_2552,N_1390,N_1073);
nand U2553 (N_2553,N_393,N_572);
nor U2554 (N_2554,N_1576,N_1101);
or U2555 (N_2555,N_866,N_388);
and U2556 (N_2556,N_1047,N_1908);
nand U2557 (N_2557,N_1279,N_1613);
nor U2558 (N_2558,N_163,N_1874);
xor U2559 (N_2559,N_511,N_1791);
and U2560 (N_2560,N_125,N_1141);
or U2561 (N_2561,N_261,N_1184);
nand U2562 (N_2562,N_1738,N_628);
and U2563 (N_2563,N_1999,N_201);
nor U2564 (N_2564,N_1471,N_1443);
nor U2565 (N_2565,N_410,N_531);
nand U2566 (N_2566,N_453,N_1550);
nand U2567 (N_2567,N_1159,N_1012);
and U2568 (N_2568,N_1042,N_1718);
nand U2569 (N_2569,N_512,N_1796);
nand U2570 (N_2570,N_767,N_850);
and U2571 (N_2571,N_674,N_932);
nor U2572 (N_2572,N_1546,N_220);
or U2573 (N_2573,N_922,N_1317);
nand U2574 (N_2574,N_400,N_1043);
and U2575 (N_2575,N_721,N_636);
nand U2576 (N_2576,N_83,N_831);
or U2577 (N_2577,N_490,N_1303);
xor U2578 (N_2578,N_1489,N_1668);
nor U2579 (N_2579,N_1971,N_1236);
xor U2580 (N_2580,N_1596,N_1248);
nand U2581 (N_2581,N_180,N_1451);
and U2582 (N_2582,N_1024,N_759);
or U2583 (N_2583,N_1310,N_156);
nand U2584 (N_2584,N_1742,N_1146);
nand U2585 (N_2585,N_387,N_977);
nor U2586 (N_2586,N_554,N_1688);
and U2587 (N_2587,N_950,N_1406);
or U2588 (N_2588,N_1663,N_1298);
nor U2589 (N_2589,N_811,N_1939);
and U2590 (N_2590,N_239,N_1892);
xnor U2591 (N_2591,N_1549,N_122);
or U2592 (N_2592,N_1188,N_1860);
nor U2593 (N_2593,N_676,N_328);
nor U2594 (N_2594,N_1511,N_314);
or U2595 (N_2595,N_438,N_1021);
nor U2596 (N_2596,N_204,N_1620);
and U2597 (N_2597,N_1792,N_1416);
or U2598 (N_2598,N_880,N_416);
or U2599 (N_2599,N_770,N_1507);
or U2600 (N_2600,N_169,N_1431);
nor U2601 (N_2601,N_1000,N_1784);
or U2602 (N_2602,N_43,N_1009);
and U2603 (N_2603,N_631,N_1955);
or U2604 (N_2604,N_1610,N_983);
xor U2605 (N_2605,N_1569,N_1831);
or U2606 (N_2606,N_428,N_1762);
and U2607 (N_2607,N_1653,N_1739);
or U2608 (N_2608,N_1345,N_1439);
and U2609 (N_2609,N_1494,N_446);
nor U2610 (N_2610,N_723,N_1556);
and U2611 (N_2611,N_1354,N_469);
nand U2612 (N_2612,N_231,N_570);
or U2613 (N_2613,N_1372,N_625);
nand U2614 (N_2614,N_1462,N_1976);
nand U2615 (N_2615,N_619,N_88);
and U2616 (N_2616,N_1076,N_1181);
nand U2617 (N_2617,N_1399,N_1013);
or U2618 (N_2618,N_380,N_1923);
or U2619 (N_2619,N_113,N_296);
xor U2620 (N_2620,N_1559,N_515);
nor U2621 (N_2621,N_1643,N_1288);
and U2622 (N_2622,N_1339,N_193);
nand U2623 (N_2623,N_1669,N_1945);
nor U2624 (N_2624,N_1206,N_1946);
nand U2625 (N_2625,N_1846,N_689);
nand U2626 (N_2626,N_1746,N_1612);
or U2627 (N_2627,N_1121,N_1369);
nand U2628 (N_2628,N_645,N_1757);
or U2629 (N_2629,N_409,N_1687);
or U2630 (N_2630,N_514,N_431);
xor U2631 (N_2631,N_525,N_1017);
nand U2632 (N_2632,N_375,N_1415);
nand U2633 (N_2633,N_1541,N_766);
nor U2634 (N_2634,N_1785,N_1708);
nand U2635 (N_2635,N_1965,N_1304);
and U2636 (N_2636,N_1006,N_693);
nand U2637 (N_2637,N_29,N_1160);
and U2638 (N_2638,N_918,N_52);
nor U2639 (N_2639,N_415,N_373);
nor U2640 (N_2640,N_1228,N_27);
or U2641 (N_2641,N_489,N_747);
and U2642 (N_2642,N_818,N_1264);
nand U2643 (N_2643,N_349,N_133);
or U2644 (N_2644,N_1125,N_1207);
and U2645 (N_2645,N_1662,N_1667);
nand U2646 (N_2646,N_1432,N_1970);
nand U2647 (N_2647,N_1949,N_1748);
and U2648 (N_2648,N_106,N_374);
and U2649 (N_2649,N_1924,N_1533);
nand U2650 (N_2650,N_714,N_1991);
or U2651 (N_2651,N_60,N_1759);
and U2652 (N_2652,N_1783,N_1185);
xor U2653 (N_2653,N_810,N_253);
or U2654 (N_2654,N_1203,N_21);
or U2655 (N_2655,N_1732,N_806);
or U2656 (N_2656,N_359,N_256);
nand U2657 (N_2657,N_586,N_1197);
and U2658 (N_2658,N_1064,N_614);
nand U2659 (N_2659,N_198,N_610);
xnor U2660 (N_2660,N_348,N_1069);
nand U2661 (N_2661,N_1981,N_1935);
nand U2662 (N_2662,N_1113,N_1589);
nor U2663 (N_2663,N_1388,N_1282);
or U2664 (N_2664,N_838,N_1689);
or U2665 (N_2665,N_1765,N_1804);
or U2666 (N_2666,N_1057,N_1174);
and U2667 (N_2667,N_396,N_984);
or U2668 (N_2668,N_141,N_1943);
nor U2669 (N_2669,N_757,N_722);
and U2670 (N_2670,N_713,N_1209);
nor U2671 (N_2671,N_120,N_413);
nand U2672 (N_2672,N_1899,N_1795);
nand U2673 (N_2673,N_1529,N_1434);
nand U2674 (N_2674,N_679,N_1060);
and U2675 (N_2675,N_363,N_242);
or U2676 (N_2676,N_1292,N_353);
nor U2677 (N_2677,N_542,N_330);
and U2678 (N_2678,N_1457,N_1995);
nor U2679 (N_2679,N_283,N_263);
or U2680 (N_2680,N_1962,N_1963);
or U2681 (N_2681,N_771,N_1744);
nand U2682 (N_2682,N_649,N_1936);
nand U2683 (N_2683,N_302,N_1166);
nand U2684 (N_2684,N_1579,N_1332);
and U2685 (N_2685,N_1430,N_1286);
nor U2686 (N_2686,N_1468,N_1320);
xor U2687 (N_2687,N_897,N_1821);
xnor U2688 (N_2688,N_538,N_331);
and U2689 (N_2689,N_561,N_1281);
nor U2690 (N_2690,N_858,N_498);
or U2691 (N_2691,N_1335,N_544);
xnor U2692 (N_2692,N_37,N_1781);
nor U2693 (N_2693,N_325,N_338);
nand U2694 (N_2694,N_1190,N_1855);
or U2695 (N_2695,N_1877,N_663);
and U2696 (N_2696,N_1587,N_1287);
or U2697 (N_2697,N_585,N_1818);
nand U2698 (N_2698,N_217,N_1881);
and U2699 (N_2699,N_533,N_1032);
nand U2700 (N_2700,N_1728,N_1414);
or U2701 (N_2701,N_783,N_1233);
xnor U2702 (N_2702,N_1424,N_521);
or U2703 (N_2703,N_1835,N_623);
or U2704 (N_2704,N_1355,N_1825);
nand U2705 (N_2705,N_1245,N_662);
xor U2706 (N_2706,N_44,N_1709);
or U2707 (N_2707,N_1833,N_712);
and U2708 (N_2708,N_1789,N_1249);
nor U2709 (N_2709,N_979,N_1472);
nand U2710 (N_2710,N_916,N_1050);
nor U2711 (N_2711,N_1394,N_1968);
or U2712 (N_2712,N_659,N_694);
nand U2713 (N_2713,N_1295,N_1743);
nor U2714 (N_2714,N_1253,N_488);
nor U2715 (N_2715,N_326,N_1539);
nor U2716 (N_2716,N_732,N_250);
or U2717 (N_2717,N_1885,N_1637);
nand U2718 (N_2718,N_982,N_1240);
and U2719 (N_2719,N_1953,N_1959);
or U2720 (N_2720,N_540,N_1602);
and U2721 (N_2721,N_634,N_912);
nor U2722 (N_2722,N_281,N_1675);
or U2723 (N_2723,N_1810,N_706);
and U2724 (N_2724,N_506,N_862);
or U2725 (N_2725,N_1695,N_699);
or U2726 (N_2726,N_168,N_500);
nor U2727 (N_2727,N_754,N_731);
and U2728 (N_2728,N_58,N_504);
and U2729 (N_2729,N_1650,N_23);
or U2730 (N_2730,N_871,N_936);
or U2731 (N_2731,N_1107,N_778);
and U2732 (N_2732,N_691,N_229);
and U2733 (N_2733,N_1608,N_960);
nand U2734 (N_2734,N_1036,N_226);
nand U2735 (N_2735,N_1607,N_638);
and U2736 (N_2736,N_1148,N_1453);
and U2737 (N_2737,N_1056,N_1381);
xor U2738 (N_2738,N_640,N_646);
nor U2739 (N_2739,N_1040,N_191);
xor U2740 (N_2740,N_598,N_1686);
or U2741 (N_2741,N_54,N_123);
or U2742 (N_2742,N_467,N_1019);
and U2743 (N_2743,N_1055,N_1357);
nor U2744 (N_2744,N_692,N_194);
and U2745 (N_2745,N_971,N_1597);
nand U2746 (N_2746,N_1519,N_1674);
and U2747 (N_2747,N_1,N_19);
nand U2748 (N_2748,N_1641,N_575);
or U2749 (N_2749,N_1333,N_955);
nand U2750 (N_2750,N_1648,N_92);
nand U2751 (N_2751,N_1079,N_342);
xnor U2752 (N_2752,N_1154,N_1733);
and U2753 (N_2753,N_1829,N_300);
or U2754 (N_2754,N_110,N_972);
and U2755 (N_2755,N_62,N_1562);
nand U2756 (N_2756,N_1411,N_919);
nor U2757 (N_2757,N_1948,N_1540);
nor U2758 (N_2758,N_974,N_1988);
or U2759 (N_2759,N_1701,N_1022);
nor U2760 (N_2760,N_140,N_600);
nor U2761 (N_2761,N_1498,N_1956);
or U2762 (N_2762,N_1349,N_1601);
or U2763 (N_2763,N_1972,N_768);
nor U2764 (N_2764,N_1217,N_1444);
nand U2765 (N_2765,N_827,N_1099);
and U2766 (N_2766,N_801,N_686);
nand U2767 (N_2767,N_1296,N_1944);
and U2768 (N_2768,N_321,N_562);
xor U2769 (N_2769,N_1595,N_1632);
or U2770 (N_2770,N_718,N_1894);
nor U2771 (N_2771,N_119,N_1553);
nand U2772 (N_2772,N_1900,N_1418);
xor U2773 (N_2773,N_1164,N_265);
xor U2774 (N_2774,N_1104,N_509);
nand U2775 (N_2775,N_695,N_535);
nand U2776 (N_2776,N_31,N_424);
or U2777 (N_2777,N_1132,N_1030);
nor U2778 (N_2778,N_529,N_1766);
xnor U2779 (N_2779,N_729,N_1790);
nand U2780 (N_2780,N_276,N_1734);
nor U2781 (N_2781,N_1514,N_1469);
or U2782 (N_2782,N_116,N_246);
nor U2783 (N_2783,N_196,N_1823);
nor U2784 (N_2784,N_1545,N_1895);
or U2785 (N_2785,N_558,N_1839);
xnor U2786 (N_2786,N_494,N_130);
xor U2787 (N_2787,N_1706,N_1192);
or U2788 (N_2788,N_1266,N_849);
nand U2789 (N_2789,N_324,N_1270);
nand U2790 (N_2790,N_921,N_577);
nand U2791 (N_2791,N_475,N_1091);
or U2792 (N_2792,N_914,N_1408);
or U2793 (N_2793,N_1046,N_1309);
nand U2794 (N_2794,N_74,N_1075);
nand U2795 (N_2795,N_1827,N_499);
and U2796 (N_2796,N_822,N_1251);
nor U2797 (N_2797,N_1703,N_1933);
nor U2798 (N_2798,N_430,N_1973);
nor U2799 (N_2799,N_552,N_440);
nor U2800 (N_2800,N_1409,N_601);
and U2801 (N_2801,N_461,N_1068);
xor U2802 (N_2802,N_1490,N_1031);
nand U2803 (N_2803,N_1654,N_227);
or U2804 (N_2804,N_1114,N_503);
and U2805 (N_2805,N_789,N_1162);
and U2806 (N_2806,N_1838,N_1700);
or U2807 (N_2807,N_939,N_1373);
or U2808 (N_2808,N_1382,N_1165);
and U2809 (N_2809,N_800,N_1745);
nor U2810 (N_2810,N_1106,N_906);
and U2811 (N_2811,N_109,N_202);
nor U2812 (N_2812,N_1741,N_288);
and U2813 (N_2813,N_1085,N_660);
or U2814 (N_2814,N_824,N_491);
nand U2815 (N_2815,N_1467,N_1560);
nor U2816 (N_2816,N_559,N_1631);
and U2817 (N_2817,N_813,N_319);
and U2818 (N_2818,N_476,N_751);
nor U2819 (N_2819,N_480,N_550);
nand U2820 (N_2820,N_1937,N_510);
nand U2821 (N_2821,N_1226,N_1461);
or U2822 (N_2822,N_166,N_1808);
and U2823 (N_2823,N_1065,N_0);
nand U2824 (N_2824,N_1586,N_618);
xor U2825 (N_2825,N_151,N_1427);
nand U2826 (N_2826,N_1204,N_1690);
nor U2827 (N_2827,N_896,N_1239);
xor U2828 (N_2828,N_82,N_76);
nor U2829 (N_2829,N_1574,N_1484);
xor U2830 (N_2830,N_278,N_1305);
and U2831 (N_2831,N_9,N_1122);
nand U2832 (N_2832,N_143,N_1112);
or U2833 (N_2833,N_688,N_1265);
or U2834 (N_2834,N_1221,N_1280);
and U2835 (N_2835,N_830,N_216);
nand U2836 (N_2836,N_1088,N_294);
nor U2837 (N_2837,N_1661,N_569);
and U2838 (N_2838,N_928,N_1660);
nor U2839 (N_2839,N_1284,N_986);
nand U2840 (N_2840,N_681,N_994);
and U2841 (N_2841,N_1985,N_1994);
nor U2842 (N_2842,N_1293,N_298);
and U2843 (N_2843,N_966,N_10);
xnor U2844 (N_2844,N_948,N_1092);
or U2845 (N_2845,N_171,N_144);
nor U2846 (N_2846,N_1581,N_1124);
nor U2847 (N_2847,N_599,N_1705);
nor U2848 (N_2848,N_1915,N_1237);
nand U2849 (N_2849,N_1604,N_1087);
xor U2850 (N_2850,N_429,N_305);
nor U2851 (N_2851,N_479,N_1930);
and U2852 (N_2852,N_255,N_951);
xor U2853 (N_2853,N_1627,N_911);
xor U2854 (N_2854,N_1850,N_299);
xnor U2855 (N_2855,N_1865,N_1423);
nand U2856 (N_2856,N_1599,N_1938);
nand U2857 (N_2857,N_1208,N_776);
xnor U2858 (N_2858,N_162,N_334);
nor U2859 (N_2859,N_414,N_1371);
and U2860 (N_2860,N_758,N_332);
nand U2861 (N_2861,N_852,N_1358);
or U2862 (N_2862,N_1052,N_1986);
or U2863 (N_2863,N_942,N_1195);
or U2864 (N_2864,N_394,N_1521);
nor U2865 (N_2865,N_793,N_703);
nor U2866 (N_2866,N_426,N_403);
and U2867 (N_2867,N_791,N_624);
nor U2868 (N_2868,N_1844,N_274);
nor U2869 (N_2869,N_1929,N_1518);
nor U2870 (N_2870,N_1872,N_1370);
and U2871 (N_2871,N_1615,N_203);
nand U2872 (N_2872,N_1147,N_1261);
xnor U2873 (N_2873,N_1353,N_1234);
and U2874 (N_2874,N_316,N_536);
xnor U2875 (N_2875,N_756,N_307);
nand U2876 (N_2876,N_1941,N_1276);
nor U2877 (N_2877,N_1078,N_38);
nor U2878 (N_2878,N_258,N_1422);
xnor U2879 (N_2879,N_1161,N_622);
or U2880 (N_2880,N_493,N_1158);
nand U2881 (N_2881,N_360,N_190);
and U2882 (N_2882,N_746,N_282);
nor U2883 (N_2883,N_596,N_1025);
xor U2884 (N_2884,N_1636,N_658);
nor U2885 (N_2885,N_1348,N_1247);
and U2886 (N_2886,N_1634,N_1194);
and U2887 (N_2887,N_59,N_750);
and U2888 (N_2888,N_1993,N_1403);
or U2889 (N_2889,N_1623,N_1719);
or U2890 (N_2890,N_132,N_340);
nor U2891 (N_2891,N_1888,N_1083);
and U2892 (N_2892,N_1297,N_1775);
and U2893 (N_2893,N_1516,N_1366);
and U2894 (N_2894,N_1898,N_1202);
nand U2895 (N_2895,N_312,N_1189);
xnor U2896 (N_2896,N_1906,N_90);
nand U2897 (N_2897,N_668,N_308);
or U2898 (N_2898,N_1966,N_1527);
nor U2899 (N_2899,N_1640,N_1008);
nor U2900 (N_2900,N_1685,N_1026);
nor U2901 (N_2901,N_1227,N_777);
nor U2902 (N_2902,N_154,N_560);
nand U2903 (N_2903,N_66,N_1509);
nor U2904 (N_2904,N_346,N_1338);
or U2905 (N_2905,N_1987,N_1225);
nand U2906 (N_2906,N_833,N_513);
nor U2907 (N_2907,N_1080,N_452);
nand U2908 (N_2908,N_172,N_1786);
nor U2909 (N_2909,N_35,N_1459);
and U2910 (N_2910,N_853,N_1554);
nor U2911 (N_2911,N_362,N_1989);
or U2912 (N_2912,N_1051,N_458);
or U2913 (N_2913,N_1961,N_1526);
nand U2914 (N_2914,N_1384,N_1735);
nand U2915 (N_2915,N_1567,N_75);
or U2916 (N_2916,N_804,N_1697);
and U2917 (N_2917,N_86,N_1897);
nor U2918 (N_2918,N_78,N_1425);
nor U2919 (N_2919,N_1302,N_310);
nor U2920 (N_2920,N_847,N_1127);
and U2921 (N_2921,N_1543,N_347);
and U2922 (N_2922,N_549,N_743);
nand U2923 (N_2923,N_1592,N_934);
xnor U2924 (N_2924,N_57,N_1568);
and U2925 (N_2925,N_725,N_1982);
and U2926 (N_2926,N_602,N_1323);
or U2927 (N_2927,N_551,N_730);
nand U2928 (N_2928,N_118,N_1268);
or U2929 (N_2929,N_823,N_89);
or U2930 (N_2930,N_351,N_7);
nor U2931 (N_2931,N_25,N_1344);
or U2932 (N_2932,N_617,N_657);
and U2933 (N_2933,N_1074,N_1410);
or U2934 (N_2934,N_735,N_534);
or U2935 (N_2935,N_1318,N_1799);
xnor U2936 (N_2936,N_1807,N_1499);
nand U2937 (N_2937,N_295,N_1255);
and U2938 (N_2938,N_1082,N_1629);
xor U2939 (N_2939,N_502,N_1896);
xor U2940 (N_2940,N_1402,N_834);
nand U2941 (N_2941,N_594,N_158);
or U2942 (N_2942,N_1324,N_1854);
or U2943 (N_2943,N_719,N_1412);
xnor U2944 (N_2944,N_1123,N_687);
nand U2945 (N_2945,N_1033,N_462);
nor U2946 (N_2946,N_280,N_1464);
xnor U2947 (N_2947,N_1720,N_1840);
nor U2948 (N_2948,N_1722,N_1847);
and U2949 (N_2949,N_264,N_395);
or U2950 (N_2950,N_1812,N_482);
and U2951 (N_2951,N_1538,N_1407);
and U2952 (N_2952,N_819,N_1758);
nand U2953 (N_2953,N_1570,N_652);
and U2954 (N_2954,N_1115,N_1283);
nor U2955 (N_2955,N_1736,N_1882);
or U2956 (N_2956,N_736,N_1419);
and U2957 (N_2957,N_604,N_12);
nor U2958 (N_2958,N_1096,N_1696);
nand U2959 (N_2959,N_1398,N_1257);
and U2960 (N_2960,N_384,N_748);
nor U2961 (N_2961,N_477,N_497);
nand U2962 (N_2962,N_442,N_1405);
nor U2963 (N_2963,N_465,N_232);
nor U2964 (N_2964,N_1887,N_473);
xnor U2965 (N_2965,N_447,N_790);
nor U2966 (N_2966,N_1582,N_1552);
or U2967 (N_2967,N_1566,N_1809);
and U2968 (N_2968,N_705,N_1041);
nor U2969 (N_2969,N_909,N_1573);
and U2970 (N_2970,N_448,N_152);
nor U2971 (N_2971,N_665,N_1725);
nand U2972 (N_2972,N_1815,N_1820);
and U2973 (N_2973,N_1337,N_1747);
nor U2974 (N_2974,N_1429,N_36);
or U2975 (N_2975,N_1483,N_1361);
nand U2976 (N_2976,N_327,N_341);
and U2977 (N_2977,N_336,N_1803);
or U2978 (N_2978,N_1841,N_1942);
and U2979 (N_2979,N_383,N_1508);
and U2980 (N_2980,N_567,N_1413);
xor U2981 (N_2981,N_507,N_678);
nor U2982 (N_2982,N_221,N_1311);
nor U2983 (N_2983,N_1639,N_1536);
xor U2984 (N_2984,N_532,N_1957);
nand U2985 (N_2985,N_1081,N_238);
and U2986 (N_2986,N_1063,N_1638);
nor U2987 (N_2987,N_1086,N_1863);
and U2988 (N_2988,N_837,N_97);
nor U2989 (N_2989,N_1331,N_1109);
or U2990 (N_2990,N_1167,N_1880);
nand U2991 (N_2991,N_195,N_115);
or U2992 (N_2992,N_1474,N_1824);
nand U2993 (N_2993,N_352,N_1072);
or U2994 (N_2994,N_24,N_1588);
or U2995 (N_2995,N_1954,N_1828);
or U2996 (N_2996,N_1658,N_1476);
or U2997 (N_2997,N_354,N_1458);
nor U2998 (N_2998,N_1702,N_286);
and U2999 (N_2999,N_589,N_1396);
xnor U3000 (N_3000,N_351,N_1851);
nand U3001 (N_3001,N_1907,N_277);
nand U3002 (N_3002,N_1293,N_505);
or U3003 (N_3003,N_462,N_456);
nor U3004 (N_3004,N_584,N_1725);
or U3005 (N_3005,N_406,N_1054);
nor U3006 (N_3006,N_1622,N_1586);
or U3007 (N_3007,N_427,N_730);
and U3008 (N_3008,N_1720,N_765);
nand U3009 (N_3009,N_1429,N_1844);
or U3010 (N_3010,N_630,N_258);
xor U3011 (N_3011,N_1034,N_39);
or U3012 (N_3012,N_231,N_1632);
and U3013 (N_3013,N_1951,N_865);
nor U3014 (N_3014,N_1782,N_1206);
or U3015 (N_3015,N_1029,N_970);
nor U3016 (N_3016,N_1427,N_473);
nand U3017 (N_3017,N_1303,N_162);
nand U3018 (N_3018,N_139,N_467);
nor U3019 (N_3019,N_1691,N_1898);
and U3020 (N_3020,N_738,N_1841);
nor U3021 (N_3021,N_325,N_34);
nand U3022 (N_3022,N_389,N_540);
xor U3023 (N_3023,N_1070,N_657);
or U3024 (N_3024,N_30,N_476);
nand U3025 (N_3025,N_1159,N_1320);
xor U3026 (N_3026,N_694,N_742);
xnor U3027 (N_3027,N_1747,N_319);
nand U3028 (N_3028,N_331,N_1745);
nand U3029 (N_3029,N_1195,N_626);
and U3030 (N_3030,N_449,N_958);
nand U3031 (N_3031,N_273,N_1661);
xnor U3032 (N_3032,N_193,N_339);
nand U3033 (N_3033,N_851,N_525);
or U3034 (N_3034,N_1660,N_1652);
nand U3035 (N_3035,N_841,N_1692);
xnor U3036 (N_3036,N_644,N_974);
xnor U3037 (N_3037,N_755,N_1796);
nand U3038 (N_3038,N_1823,N_448);
nand U3039 (N_3039,N_1393,N_1361);
or U3040 (N_3040,N_1502,N_1445);
nand U3041 (N_3041,N_1913,N_1728);
nor U3042 (N_3042,N_1241,N_461);
nand U3043 (N_3043,N_1431,N_1955);
nor U3044 (N_3044,N_1206,N_1519);
and U3045 (N_3045,N_932,N_1291);
nor U3046 (N_3046,N_979,N_236);
nor U3047 (N_3047,N_1118,N_286);
xor U3048 (N_3048,N_210,N_861);
or U3049 (N_3049,N_1663,N_1193);
and U3050 (N_3050,N_159,N_383);
nand U3051 (N_3051,N_113,N_1514);
and U3052 (N_3052,N_1859,N_899);
nor U3053 (N_3053,N_1066,N_419);
nand U3054 (N_3054,N_217,N_1409);
and U3055 (N_3055,N_1300,N_575);
and U3056 (N_3056,N_567,N_551);
nor U3057 (N_3057,N_1189,N_1009);
nand U3058 (N_3058,N_654,N_1377);
nand U3059 (N_3059,N_1685,N_696);
or U3060 (N_3060,N_1617,N_1828);
nand U3061 (N_3061,N_868,N_514);
nor U3062 (N_3062,N_1593,N_816);
or U3063 (N_3063,N_1140,N_394);
nor U3064 (N_3064,N_1451,N_1575);
nor U3065 (N_3065,N_1200,N_1437);
nand U3066 (N_3066,N_137,N_1188);
nand U3067 (N_3067,N_1952,N_1555);
nor U3068 (N_3068,N_1930,N_551);
or U3069 (N_3069,N_1807,N_820);
nand U3070 (N_3070,N_404,N_13);
or U3071 (N_3071,N_349,N_388);
and U3072 (N_3072,N_1326,N_1480);
or U3073 (N_3073,N_382,N_1183);
or U3074 (N_3074,N_913,N_220);
or U3075 (N_3075,N_998,N_223);
and U3076 (N_3076,N_631,N_1492);
nand U3077 (N_3077,N_847,N_1514);
nor U3078 (N_3078,N_1653,N_513);
or U3079 (N_3079,N_588,N_474);
nand U3080 (N_3080,N_80,N_1536);
or U3081 (N_3081,N_1067,N_637);
xor U3082 (N_3082,N_260,N_521);
nor U3083 (N_3083,N_552,N_1954);
nor U3084 (N_3084,N_901,N_668);
nor U3085 (N_3085,N_253,N_1273);
nand U3086 (N_3086,N_599,N_516);
nor U3087 (N_3087,N_957,N_560);
and U3088 (N_3088,N_711,N_1810);
or U3089 (N_3089,N_957,N_1175);
and U3090 (N_3090,N_760,N_1417);
and U3091 (N_3091,N_858,N_1336);
nor U3092 (N_3092,N_895,N_1459);
nand U3093 (N_3093,N_1688,N_188);
nor U3094 (N_3094,N_681,N_45);
nor U3095 (N_3095,N_30,N_1623);
xor U3096 (N_3096,N_962,N_1580);
and U3097 (N_3097,N_552,N_1177);
nor U3098 (N_3098,N_317,N_489);
or U3099 (N_3099,N_1629,N_1525);
nor U3100 (N_3100,N_1367,N_1827);
or U3101 (N_3101,N_598,N_520);
nand U3102 (N_3102,N_565,N_1387);
xor U3103 (N_3103,N_359,N_1725);
nand U3104 (N_3104,N_1890,N_1157);
and U3105 (N_3105,N_1949,N_1368);
nor U3106 (N_3106,N_176,N_766);
and U3107 (N_3107,N_33,N_853);
and U3108 (N_3108,N_1510,N_421);
nor U3109 (N_3109,N_154,N_1034);
nand U3110 (N_3110,N_1754,N_1512);
nor U3111 (N_3111,N_589,N_1079);
and U3112 (N_3112,N_1160,N_1676);
and U3113 (N_3113,N_7,N_508);
or U3114 (N_3114,N_1191,N_1237);
xnor U3115 (N_3115,N_517,N_1307);
nand U3116 (N_3116,N_1205,N_439);
nand U3117 (N_3117,N_128,N_653);
nand U3118 (N_3118,N_1172,N_291);
nand U3119 (N_3119,N_1739,N_1184);
nand U3120 (N_3120,N_23,N_620);
or U3121 (N_3121,N_1070,N_504);
nor U3122 (N_3122,N_1837,N_1726);
or U3123 (N_3123,N_1008,N_1819);
or U3124 (N_3124,N_115,N_990);
nor U3125 (N_3125,N_582,N_1825);
nand U3126 (N_3126,N_1417,N_1674);
and U3127 (N_3127,N_150,N_1856);
nor U3128 (N_3128,N_394,N_822);
nand U3129 (N_3129,N_314,N_1979);
nor U3130 (N_3130,N_1010,N_1315);
nand U3131 (N_3131,N_1795,N_1568);
nand U3132 (N_3132,N_103,N_1829);
or U3133 (N_3133,N_1209,N_706);
or U3134 (N_3134,N_1788,N_1990);
and U3135 (N_3135,N_89,N_785);
and U3136 (N_3136,N_1649,N_659);
nand U3137 (N_3137,N_379,N_798);
nor U3138 (N_3138,N_1658,N_835);
or U3139 (N_3139,N_571,N_1349);
nor U3140 (N_3140,N_1859,N_631);
nand U3141 (N_3141,N_573,N_509);
nand U3142 (N_3142,N_1446,N_1454);
nor U3143 (N_3143,N_913,N_1786);
or U3144 (N_3144,N_487,N_963);
nor U3145 (N_3145,N_1387,N_1716);
nor U3146 (N_3146,N_1290,N_1448);
nor U3147 (N_3147,N_105,N_1231);
and U3148 (N_3148,N_329,N_1324);
nand U3149 (N_3149,N_130,N_1148);
and U3150 (N_3150,N_680,N_1573);
nor U3151 (N_3151,N_1678,N_750);
or U3152 (N_3152,N_553,N_735);
and U3153 (N_3153,N_780,N_820);
and U3154 (N_3154,N_576,N_1541);
or U3155 (N_3155,N_1870,N_1432);
nor U3156 (N_3156,N_580,N_277);
or U3157 (N_3157,N_1141,N_831);
and U3158 (N_3158,N_1959,N_748);
nand U3159 (N_3159,N_1558,N_1062);
nor U3160 (N_3160,N_851,N_1426);
and U3161 (N_3161,N_1044,N_1481);
and U3162 (N_3162,N_908,N_1730);
or U3163 (N_3163,N_474,N_526);
xor U3164 (N_3164,N_762,N_1598);
or U3165 (N_3165,N_1834,N_1699);
xor U3166 (N_3166,N_201,N_1472);
nor U3167 (N_3167,N_838,N_1767);
nand U3168 (N_3168,N_132,N_1809);
nand U3169 (N_3169,N_622,N_887);
nand U3170 (N_3170,N_785,N_1888);
nand U3171 (N_3171,N_890,N_1514);
nor U3172 (N_3172,N_1333,N_147);
and U3173 (N_3173,N_1184,N_1401);
and U3174 (N_3174,N_603,N_1417);
or U3175 (N_3175,N_880,N_1281);
and U3176 (N_3176,N_1325,N_1336);
or U3177 (N_3177,N_1034,N_918);
nand U3178 (N_3178,N_334,N_1222);
nand U3179 (N_3179,N_834,N_32);
or U3180 (N_3180,N_1692,N_343);
xnor U3181 (N_3181,N_1319,N_1033);
or U3182 (N_3182,N_1280,N_1918);
nand U3183 (N_3183,N_512,N_1159);
xnor U3184 (N_3184,N_976,N_1113);
nor U3185 (N_3185,N_163,N_1325);
nand U3186 (N_3186,N_499,N_600);
nand U3187 (N_3187,N_310,N_24);
and U3188 (N_3188,N_923,N_150);
nand U3189 (N_3189,N_704,N_284);
and U3190 (N_3190,N_973,N_841);
and U3191 (N_3191,N_895,N_491);
nor U3192 (N_3192,N_1439,N_833);
and U3193 (N_3193,N_1336,N_914);
nand U3194 (N_3194,N_587,N_1005);
nor U3195 (N_3195,N_1115,N_555);
xor U3196 (N_3196,N_1277,N_758);
or U3197 (N_3197,N_1228,N_282);
or U3198 (N_3198,N_506,N_109);
nand U3199 (N_3199,N_561,N_1044);
or U3200 (N_3200,N_874,N_749);
nand U3201 (N_3201,N_1580,N_1433);
and U3202 (N_3202,N_1072,N_900);
and U3203 (N_3203,N_452,N_1064);
and U3204 (N_3204,N_491,N_1107);
xnor U3205 (N_3205,N_597,N_693);
nor U3206 (N_3206,N_1300,N_1234);
nand U3207 (N_3207,N_1739,N_1331);
nand U3208 (N_3208,N_1934,N_1922);
nor U3209 (N_3209,N_1752,N_1849);
nor U3210 (N_3210,N_690,N_873);
nor U3211 (N_3211,N_1974,N_855);
and U3212 (N_3212,N_1105,N_1337);
or U3213 (N_3213,N_1503,N_109);
or U3214 (N_3214,N_1498,N_1792);
nand U3215 (N_3215,N_639,N_954);
nor U3216 (N_3216,N_1890,N_98);
and U3217 (N_3217,N_1627,N_1386);
nand U3218 (N_3218,N_1357,N_25);
and U3219 (N_3219,N_1538,N_1774);
nand U3220 (N_3220,N_1655,N_702);
or U3221 (N_3221,N_308,N_99);
nor U3222 (N_3222,N_1417,N_1219);
nor U3223 (N_3223,N_777,N_1119);
nand U3224 (N_3224,N_389,N_1099);
nor U3225 (N_3225,N_1600,N_786);
nand U3226 (N_3226,N_563,N_1846);
nand U3227 (N_3227,N_582,N_1303);
nor U3228 (N_3228,N_1666,N_1911);
or U3229 (N_3229,N_184,N_737);
or U3230 (N_3230,N_434,N_802);
and U3231 (N_3231,N_1686,N_896);
nand U3232 (N_3232,N_1980,N_325);
or U3233 (N_3233,N_1581,N_285);
nand U3234 (N_3234,N_1019,N_501);
nand U3235 (N_3235,N_404,N_1279);
nand U3236 (N_3236,N_112,N_161);
xnor U3237 (N_3237,N_1538,N_810);
nor U3238 (N_3238,N_1783,N_1927);
xnor U3239 (N_3239,N_1900,N_1088);
or U3240 (N_3240,N_62,N_1584);
xnor U3241 (N_3241,N_1047,N_380);
nand U3242 (N_3242,N_1848,N_371);
and U3243 (N_3243,N_1696,N_878);
and U3244 (N_3244,N_1146,N_1087);
nand U3245 (N_3245,N_1493,N_760);
or U3246 (N_3246,N_1147,N_685);
xor U3247 (N_3247,N_1706,N_150);
nor U3248 (N_3248,N_1008,N_166);
nor U3249 (N_3249,N_1953,N_194);
nor U3250 (N_3250,N_777,N_1131);
or U3251 (N_3251,N_1354,N_1195);
nor U3252 (N_3252,N_21,N_126);
xnor U3253 (N_3253,N_1807,N_617);
and U3254 (N_3254,N_513,N_404);
or U3255 (N_3255,N_1593,N_598);
nor U3256 (N_3256,N_1015,N_1931);
xor U3257 (N_3257,N_1065,N_1286);
nor U3258 (N_3258,N_1142,N_1429);
xor U3259 (N_3259,N_1098,N_749);
nor U3260 (N_3260,N_1903,N_1438);
and U3261 (N_3261,N_763,N_1935);
nor U3262 (N_3262,N_1727,N_220);
xnor U3263 (N_3263,N_209,N_249);
and U3264 (N_3264,N_1408,N_679);
or U3265 (N_3265,N_1018,N_1128);
nor U3266 (N_3266,N_204,N_1375);
or U3267 (N_3267,N_1831,N_413);
nand U3268 (N_3268,N_1814,N_1698);
nand U3269 (N_3269,N_1202,N_413);
nand U3270 (N_3270,N_1469,N_1589);
nor U3271 (N_3271,N_928,N_988);
xnor U3272 (N_3272,N_1717,N_1375);
and U3273 (N_3273,N_128,N_270);
and U3274 (N_3274,N_450,N_11);
and U3275 (N_3275,N_255,N_1692);
or U3276 (N_3276,N_577,N_1978);
nor U3277 (N_3277,N_436,N_1628);
and U3278 (N_3278,N_1258,N_800);
xnor U3279 (N_3279,N_175,N_772);
nand U3280 (N_3280,N_788,N_1989);
nand U3281 (N_3281,N_1525,N_430);
or U3282 (N_3282,N_98,N_147);
nor U3283 (N_3283,N_986,N_498);
and U3284 (N_3284,N_824,N_571);
nand U3285 (N_3285,N_7,N_1462);
and U3286 (N_3286,N_720,N_1252);
and U3287 (N_3287,N_50,N_820);
nand U3288 (N_3288,N_1417,N_778);
and U3289 (N_3289,N_110,N_98);
and U3290 (N_3290,N_1877,N_923);
or U3291 (N_3291,N_1607,N_715);
or U3292 (N_3292,N_1891,N_1458);
xor U3293 (N_3293,N_1975,N_580);
and U3294 (N_3294,N_1055,N_1227);
nor U3295 (N_3295,N_1519,N_1279);
and U3296 (N_3296,N_1655,N_337);
nor U3297 (N_3297,N_863,N_840);
nor U3298 (N_3298,N_492,N_1586);
and U3299 (N_3299,N_1731,N_1568);
nor U3300 (N_3300,N_624,N_1666);
nand U3301 (N_3301,N_223,N_499);
nand U3302 (N_3302,N_990,N_23);
xnor U3303 (N_3303,N_1864,N_712);
xnor U3304 (N_3304,N_51,N_1589);
nor U3305 (N_3305,N_755,N_30);
or U3306 (N_3306,N_425,N_1591);
or U3307 (N_3307,N_538,N_279);
nand U3308 (N_3308,N_863,N_617);
and U3309 (N_3309,N_314,N_1251);
or U3310 (N_3310,N_1563,N_1547);
or U3311 (N_3311,N_1849,N_1995);
xnor U3312 (N_3312,N_929,N_279);
xnor U3313 (N_3313,N_654,N_603);
nor U3314 (N_3314,N_264,N_1782);
nand U3315 (N_3315,N_1039,N_1069);
nand U3316 (N_3316,N_582,N_1041);
and U3317 (N_3317,N_1379,N_1498);
nand U3318 (N_3318,N_722,N_1878);
nor U3319 (N_3319,N_107,N_651);
nor U3320 (N_3320,N_551,N_1631);
or U3321 (N_3321,N_1618,N_225);
xor U3322 (N_3322,N_1653,N_1524);
or U3323 (N_3323,N_1943,N_431);
and U3324 (N_3324,N_894,N_538);
xor U3325 (N_3325,N_748,N_330);
nand U3326 (N_3326,N_1607,N_1160);
nand U3327 (N_3327,N_139,N_1627);
nor U3328 (N_3328,N_1043,N_54);
or U3329 (N_3329,N_801,N_1601);
xor U3330 (N_3330,N_1930,N_250);
nand U3331 (N_3331,N_1748,N_735);
nor U3332 (N_3332,N_1159,N_237);
or U3333 (N_3333,N_38,N_247);
or U3334 (N_3334,N_216,N_723);
nor U3335 (N_3335,N_1164,N_922);
nand U3336 (N_3336,N_571,N_1251);
nand U3337 (N_3337,N_4,N_64);
or U3338 (N_3338,N_1892,N_992);
nand U3339 (N_3339,N_842,N_1205);
nand U3340 (N_3340,N_1668,N_1627);
nand U3341 (N_3341,N_1355,N_1153);
or U3342 (N_3342,N_467,N_678);
nor U3343 (N_3343,N_514,N_565);
nor U3344 (N_3344,N_9,N_297);
nand U3345 (N_3345,N_1001,N_1903);
and U3346 (N_3346,N_181,N_726);
and U3347 (N_3347,N_418,N_579);
nor U3348 (N_3348,N_937,N_1541);
xor U3349 (N_3349,N_1121,N_1983);
and U3350 (N_3350,N_1923,N_354);
xnor U3351 (N_3351,N_292,N_373);
and U3352 (N_3352,N_1553,N_1012);
nand U3353 (N_3353,N_956,N_1448);
nor U3354 (N_3354,N_1664,N_1172);
nand U3355 (N_3355,N_1599,N_316);
xnor U3356 (N_3356,N_1089,N_1217);
nor U3357 (N_3357,N_1189,N_1259);
nor U3358 (N_3358,N_1302,N_555);
or U3359 (N_3359,N_1642,N_1342);
nand U3360 (N_3360,N_2,N_1005);
nor U3361 (N_3361,N_1611,N_314);
and U3362 (N_3362,N_924,N_1659);
nand U3363 (N_3363,N_1441,N_1270);
xor U3364 (N_3364,N_225,N_29);
and U3365 (N_3365,N_864,N_401);
and U3366 (N_3366,N_1607,N_317);
and U3367 (N_3367,N_1686,N_1329);
or U3368 (N_3368,N_954,N_1423);
nand U3369 (N_3369,N_1414,N_746);
or U3370 (N_3370,N_1977,N_1446);
and U3371 (N_3371,N_1949,N_1279);
and U3372 (N_3372,N_193,N_587);
and U3373 (N_3373,N_661,N_1407);
and U3374 (N_3374,N_1850,N_659);
nand U3375 (N_3375,N_345,N_1652);
nand U3376 (N_3376,N_484,N_49);
nand U3377 (N_3377,N_1845,N_1062);
xnor U3378 (N_3378,N_1663,N_366);
nor U3379 (N_3379,N_845,N_1653);
xnor U3380 (N_3380,N_1189,N_1939);
or U3381 (N_3381,N_57,N_622);
or U3382 (N_3382,N_1571,N_1860);
and U3383 (N_3383,N_475,N_500);
nand U3384 (N_3384,N_1036,N_1400);
nor U3385 (N_3385,N_1905,N_819);
nand U3386 (N_3386,N_675,N_1513);
nor U3387 (N_3387,N_1878,N_1143);
xor U3388 (N_3388,N_792,N_498);
or U3389 (N_3389,N_635,N_1069);
xnor U3390 (N_3390,N_1030,N_935);
nand U3391 (N_3391,N_1696,N_1727);
nand U3392 (N_3392,N_995,N_161);
nor U3393 (N_3393,N_696,N_1751);
or U3394 (N_3394,N_1905,N_759);
and U3395 (N_3395,N_1792,N_386);
nor U3396 (N_3396,N_1089,N_155);
and U3397 (N_3397,N_736,N_757);
and U3398 (N_3398,N_1765,N_564);
xor U3399 (N_3399,N_529,N_1039);
or U3400 (N_3400,N_1176,N_32);
and U3401 (N_3401,N_302,N_1878);
or U3402 (N_3402,N_454,N_1608);
and U3403 (N_3403,N_1095,N_245);
nor U3404 (N_3404,N_1298,N_1981);
nor U3405 (N_3405,N_597,N_1529);
or U3406 (N_3406,N_286,N_1648);
or U3407 (N_3407,N_1670,N_1192);
nand U3408 (N_3408,N_1718,N_1218);
or U3409 (N_3409,N_704,N_1609);
nor U3410 (N_3410,N_203,N_1758);
and U3411 (N_3411,N_766,N_804);
xor U3412 (N_3412,N_1133,N_1498);
or U3413 (N_3413,N_1613,N_850);
and U3414 (N_3414,N_722,N_42);
or U3415 (N_3415,N_533,N_1299);
nand U3416 (N_3416,N_1873,N_284);
and U3417 (N_3417,N_1967,N_1876);
nor U3418 (N_3418,N_1769,N_801);
nor U3419 (N_3419,N_318,N_1252);
nand U3420 (N_3420,N_1621,N_1564);
and U3421 (N_3421,N_918,N_425);
or U3422 (N_3422,N_690,N_1239);
and U3423 (N_3423,N_569,N_1207);
nor U3424 (N_3424,N_1322,N_802);
and U3425 (N_3425,N_1873,N_775);
or U3426 (N_3426,N_631,N_597);
or U3427 (N_3427,N_700,N_202);
and U3428 (N_3428,N_741,N_387);
nor U3429 (N_3429,N_222,N_430);
nor U3430 (N_3430,N_1120,N_1758);
and U3431 (N_3431,N_1001,N_738);
or U3432 (N_3432,N_569,N_1728);
nor U3433 (N_3433,N_994,N_357);
and U3434 (N_3434,N_1305,N_1417);
and U3435 (N_3435,N_43,N_1758);
and U3436 (N_3436,N_1456,N_1369);
nor U3437 (N_3437,N_601,N_173);
nor U3438 (N_3438,N_409,N_1368);
nor U3439 (N_3439,N_1464,N_1202);
and U3440 (N_3440,N_1863,N_1532);
and U3441 (N_3441,N_492,N_193);
xnor U3442 (N_3442,N_1872,N_1339);
and U3443 (N_3443,N_250,N_985);
or U3444 (N_3444,N_162,N_1843);
xnor U3445 (N_3445,N_1353,N_1772);
or U3446 (N_3446,N_1595,N_619);
xor U3447 (N_3447,N_1175,N_1516);
xnor U3448 (N_3448,N_844,N_173);
nand U3449 (N_3449,N_1060,N_471);
or U3450 (N_3450,N_179,N_1909);
nand U3451 (N_3451,N_763,N_1226);
or U3452 (N_3452,N_1470,N_1280);
nand U3453 (N_3453,N_363,N_684);
nor U3454 (N_3454,N_351,N_1804);
xnor U3455 (N_3455,N_987,N_674);
nand U3456 (N_3456,N_493,N_741);
and U3457 (N_3457,N_172,N_1744);
nand U3458 (N_3458,N_1848,N_137);
nand U3459 (N_3459,N_148,N_1936);
xor U3460 (N_3460,N_47,N_125);
and U3461 (N_3461,N_479,N_1526);
nor U3462 (N_3462,N_281,N_1197);
nand U3463 (N_3463,N_1426,N_227);
or U3464 (N_3464,N_504,N_224);
nand U3465 (N_3465,N_137,N_1100);
nand U3466 (N_3466,N_815,N_88);
or U3467 (N_3467,N_899,N_1386);
and U3468 (N_3468,N_298,N_1573);
and U3469 (N_3469,N_405,N_102);
nor U3470 (N_3470,N_243,N_561);
or U3471 (N_3471,N_717,N_1361);
xnor U3472 (N_3472,N_1453,N_1524);
or U3473 (N_3473,N_1793,N_1280);
nor U3474 (N_3474,N_58,N_1348);
xor U3475 (N_3475,N_182,N_659);
nor U3476 (N_3476,N_1093,N_1451);
or U3477 (N_3477,N_1077,N_1920);
nand U3478 (N_3478,N_193,N_968);
nor U3479 (N_3479,N_1031,N_1839);
and U3480 (N_3480,N_36,N_1297);
nor U3481 (N_3481,N_34,N_678);
and U3482 (N_3482,N_1036,N_37);
and U3483 (N_3483,N_1100,N_71);
or U3484 (N_3484,N_1936,N_924);
nand U3485 (N_3485,N_283,N_108);
nand U3486 (N_3486,N_922,N_1728);
or U3487 (N_3487,N_1680,N_0);
and U3488 (N_3488,N_623,N_128);
xor U3489 (N_3489,N_810,N_1007);
and U3490 (N_3490,N_1323,N_1141);
or U3491 (N_3491,N_1590,N_1541);
nand U3492 (N_3492,N_255,N_269);
and U3493 (N_3493,N_699,N_457);
or U3494 (N_3494,N_613,N_594);
xnor U3495 (N_3495,N_1721,N_121);
xnor U3496 (N_3496,N_37,N_293);
nand U3497 (N_3497,N_234,N_746);
nor U3498 (N_3498,N_1400,N_1238);
and U3499 (N_3499,N_64,N_403);
xor U3500 (N_3500,N_283,N_1388);
and U3501 (N_3501,N_108,N_314);
and U3502 (N_3502,N_74,N_1949);
or U3503 (N_3503,N_190,N_1615);
nor U3504 (N_3504,N_654,N_1246);
nor U3505 (N_3505,N_1047,N_316);
xnor U3506 (N_3506,N_933,N_244);
nand U3507 (N_3507,N_1236,N_44);
xor U3508 (N_3508,N_484,N_1827);
nand U3509 (N_3509,N_827,N_21);
nand U3510 (N_3510,N_224,N_1687);
nor U3511 (N_3511,N_1859,N_909);
nand U3512 (N_3512,N_751,N_383);
or U3513 (N_3513,N_350,N_1546);
xnor U3514 (N_3514,N_72,N_1233);
and U3515 (N_3515,N_490,N_1344);
or U3516 (N_3516,N_456,N_1890);
nand U3517 (N_3517,N_914,N_1277);
and U3518 (N_3518,N_1888,N_513);
or U3519 (N_3519,N_720,N_762);
or U3520 (N_3520,N_1506,N_1839);
and U3521 (N_3521,N_1571,N_1189);
or U3522 (N_3522,N_202,N_1701);
xnor U3523 (N_3523,N_26,N_675);
or U3524 (N_3524,N_1447,N_186);
nor U3525 (N_3525,N_474,N_635);
nand U3526 (N_3526,N_1853,N_140);
nand U3527 (N_3527,N_1823,N_1886);
nand U3528 (N_3528,N_1434,N_356);
nor U3529 (N_3529,N_1333,N_1167);
xnor U3530 (N_3530,N_876,N_899);
or U3531 (N_3531,N_1429,N_224);
or U3532 (N_3532,N_1413,N_241);
nand U3533 (N_3533,N_421,N_647);
nor U3534 (N_3534,N_1645,N_1302);
nand U3535 (N_3535,N_1571,N_1537);
nor U3536 (N_3536,N_1843,N_912);
and U3537 (N_3537,N_296,N_1458);
or U3538 (N_3538,N_1538,N_240);
and U3539 (N_3539,N_1914,N_1016);
xnor U3540 (N_3540,N_1240,N_833);
nor U3541 (N_3541,N_1359,N_443);
nand U3542 (N_3542,N_1110,N_821);
xnor U3543 (N_3543,N_218,N_1815);
nor U3544 (N_3544,N_1945,N_526);
nand U3545 (N_3545,N_1026,N_1191);
nand U3546 (N_3546,N_1353,N_1355);
or U3547 (N_3547,N_849,N_673);
nand U3548 (N_3548,N_349,N_248);
or U3549 (N_3549,N_1642,N_1159);
and U3550 (N_3550,N_969,N_1897);
and U3551 (N_3551,N_1440,N_1645);
or U3552 (N_3552,N_1945,N_530);
nor U3553 (N_3553,N_1067,N_1184);
nor U3554 (N_3554,N_1226,N_1275);
or U3555 (N_3555,N_1849,N_1765);
or U3556 (N_3556,N_249,N_1012);
and U3557 (N_3557,N_1381,N_1344);
or U3558 (N_3558,N_240,N_118);
and U3559 (N_3559,N_1934,N_326);
nand U3560 (N_3560,N_421,N_796);
or U3561 (N_3561,N_501,N_1386);
nor U3562 (N_3562,N_932,N_777);
and U3563 (N_3563,N_806,N_1052);
or U3564 (N_3564,N_64,N_104);
nor U3565 (N_3565,N_547,N_761);
nor U3566 (N_3566,N_274,N_123);
nand U3567 (N_3567,N_273,N_1322);
nor U3568 (N_3568,N_1778,N_1213);
nor U3569 (N_3569,N_1343,N_800);
or U3570 (N_3570,N_516,N_1064);
xor U3571 (N_3571,N_1124,N_184);
nor U3572 (N_3572,N_1783,N_1288);
and U3573 (N_3573,N_1102,N_460);
and U3574 (N_3574,N_805,N_798);
nor U3575 (N_3575,N_977,N_1993);
nand U3576 (N_3576,N_1131,N_761);
and U3577 (N_3577,N_440,N_373);
nor U3578 (N_3578,N_1958,N_946);
or U3579 (N_3579,N_1038,N_1897);
and U3580 (N_3580,N_273,N_1249);
nand U3581 (N_3581,N_1310,N_1957);
or U3582 (N_3582,N_1266,N_1427);
nor U3583 (N_3583,N_1270,N_1188);
nor U3584 (N_3584,N_1768,N_822);
nand U3585 (N_3585,N_60,N_450);
and U3586 (N_3586,N_1855,N_837);
or U3587 (N_3587,N_1959,N_738);
and U3588 (N_3588,N_1250,N_863);
and U3589 (N_3589,N_1646,N_337);
nand U3590 (N_3590,N_1466,N_284);
nor U3591 (N_3591,N_1504,N_1326);
xnor U3592 (N_3592,N_657,N_1144);
nor U3593 (N_3593,N_46,N_1571);
nand U3594 (N_3594,N_985,N_1976);
and U3595 (N_3595,N_1024,N_540);
nand U3596 (N_3596,N_373,N_1225);
or U3597 (N_3597,N_1359,N_1285);
and U3598 (N_3598,N_1206,N_5);
xor U3599 (N_3599,N_299,N_737);
and U3600 (N_3600,N_442,N_1800);
nor U3601 (N_3601,N_1202,N_900);
nand U3602 (N_3602,N_506,N_1595);
or U3603 (N_3603,N_1264,N_152);
nand U3604 (N_3604,N_282,N_1436);
nand U3605 (N_3605,N_750,N_1670);
nor U3606 (N_3606,N_1643,N_422);
nor U3607 (N_3607,N_344,N_1068);
xnor U3608 (N_3608,N_1670,N_334);
xor U3609 (N_3609,N_1674,N_632);
nor U3610 (N_3610,N_1547,N_1711);
or U3611 (N_3611,N_732,N_1200);
or U3612 (N_3612,N_864,N_1347);
nand U3613 (N_3613,N_1153,N_356);
or U3614 (N_3614,N_324,N_1624);
and U3615 (N_3615,N_1268,N_1047);
or U3616 (N_3616,N_1496,N_43);
or U3617 (N_3617,N_311,N_1075);
nor U3618 (N_3618,N_1939,N_1612);
nand U3619 (N_3619,N_1698,N_1973);
nand U3620 (N_3620,N_745,N_1680);
nor U3621 (N_3621,N_1544,N_1054);
nand U3622 (N_3622,N_980,N_1423);
and U3623 (N_3623,N_1005,N_949);
nand U3624 (N_3624,N_736,N_245);
nor U3625 (N_3625,N_362,N_1716);
or U3626 (N_3626,N_1179,N_1839);
and U3627 (N_3627,N_1458,N_631);
or U3628 (N_3628,N_1878,N_1249);
nor U3629 (N_3629,N_1783,N_1107);
xnor U3630 (N_3630,N_317,N_389);
nor U3631 (N_3631,N_1321,N_1926);
or U3632 (N_3632,N_1447,N_38);
nand U3633 (N_3633,N_1793,N_1428);
or U3634 (N_3634,N_402,N_1993);
nor U3635 (N_3635,N_1824,N_1277);
or U3636 (N_3636,N_1158,N_1622);
nor U3637 (N_3637,N_1295,N_636);
nand U3638 (N_3638,N_1549,N_1640);
xor U3639 (N_3639,N_359,N_329);
or U3640 (N_3640,N_827,N_570);
and U3641 (N_3641,N_1905,N_1042);
nor U3642 (N_3642,N_1468,N_1898);
and U3643 (N_3643,N_311,N_1570);
and U3644 (N_3644,N_386,N_200);
and U3645 (N_3645,N_657,N_1385);
nor U3646 (N_3646,N_159,N_963);
and U3647 (N_3647,N_889,N_771);
and U3648 (N_3648,N_1406,N_406);
or U3649 (N_3649,N_1810,N_46);
nand U3650 (N_3650,N_206,N_342);
nand U3651 (N_3651,N_732,N_1114);
or U3652 (N_3652,N_1961,N_409);
nand U3653 (N_3653,N_1626,N_981);
nor U3654 (N_3654,N_1896,N_1857);
or U3655 (N_3655,N_228,N_1693);
and U3656 (N_3656,N_1555,N_1463);
and U3657 (N_3657,N_1274,N_1756);
and U3658 (N_3658,N_1200,N_350);
xor U3659 (N_3659,N_1800,N_991);
nor U3660 (N_3660,N_1019,N_341);
nor U3661 (N_3661,N_204,N_880);
and U3662 (N_3662,N_422,N_271);
or U3663 (N_3663,N_1115,N_506);
or U3664 (N_3664,N_622,N_1087);
nand U3665 (N_3665,N_290,N_1817);
nor U3666 (N_3666,N_1683,N_1233);
xnor U3667 (N_3667,N_545,N_1579);
and U3668 (N_3668,N_1555,N_390);
nor U3669 (N_3669,N_430,N_1922);
nor U3670 (N_3670,N_175,N_707);
nor U3671 (N_3671,N_1633,N_1356);
or U3672 (N_3672,N_1386,N_1446);
and U3673 (N_3673,N_246,N_1140);
nand U3674 (N_3674,N_1239,N_1500);
xor U3675 (N_3675,N_1774,N_1843);
and U3676 (N_3676,N_1195,N_999);
nor U3677 (N_3677,N_509,N_1833);
and U3678 (N_3678,N_898,N_970);
and U3679 (N_3679,N_1873,N_1249);
nand U3680 (N_3680,N_1082,N_1513);
nand U3681 (N_3681,N_1945,N_1445);
and U3682 (N_3682,N_1979,N_13);
and U3683 (N_3683,N_841,N_1281);
nor U3684 (N_3684,N_555,N_57);
and U3685 (N_3685,N_1783,N_526);
and U3686 (N_3686,N_1118,N_615);
nand U3687 (N_3687,N_306,N_1582);
and U3688 (N_3688,N_261,N_1180);
or U3689 (N_3689,N_990,N_1243);
or U3690 (N_3690,N_72,N_650);
and U3691 (N_3691,N_167,N_1034);
nor U3692 (N_3692,N_1357,N_1889);
xnor U3693 (N_3693,N_35,N_973);
and U3694 (N_3694,N_490,N_1449);
or U3695 (N_3695,N_422,N_214);
and U3696 (N_3696,N_1782,N_41);
nor U3697 (N_3697,N_1636,N_369);
and U3698 (N_3698,N_1469,N_1357);
xor U3699 (N_3699,N_1388,N_797);
nand U3700 (N_3700,N_1474,N_463);
xor U3701 (N_3701,N_1093,N_355);
nor U3702 (N_3702,N_1358,N_1071);
or U3703 (N_3703,N_1788,N_834);
or U3704 (N_3704,N_435,N_1048);
nand U3705 (N_3705,N_230,N_1168);
nor U3706 (N_3706,N_1703,N_227);
and U3707 (N_3707,N_183,N_1025);
and U3708 (N_3708,N_416,N_1867);
nand U3709 (N_3709,N_872,N_15);
nand U3710 (N_3710,N_795,N_1862);
and U3711 (N_3711,N_1610,N_379);
nor U3712 (N_3712,N_114,N_1679);
or U3713 (N_3713,N_727,N_99);
and U3714 (N_3714,N_1981,N_136);
or U3715 (N_3715,N_389,N_470);
xnor U3716 (N_3716,N_1057,N_128);
and U3717 (N_3717,N_165,N_1809);
nand U3718 (N_3718,N_172,N_501);
nor U3719 (N_3719,N_954,N_1239);
nand U3720 (N_3720,N_1940,N_114);
or U3721 (N_3721,N_1157,N_1202);
nand U3722 (N_3722,N_977,N_1570);
xor U3723 (N_3723,N_963,N_391);
or U3724 (N_3724,N_308,N_134);
nor U3725 (N_3725,N_1214,N_454);
and U3726 (N_3726,N_84,N_1129);
and U3727 (N_3727,N_1027,N_583);
nand U3728 (N_3728,N_520,N_1904);
nor U3729 (N_3729,N_1452,N_231);
nor U3730 (N_3730,N_1912,N_1221);
or U3731 (N_3731,N_869,N_1440);
nor U3732 (N_3732,N_84,N_1505);
and U3733 (N_3733,N_306,N_826);
nor U3734 (N_3734,N_1975,N_720);
nor U3735 (N_3735,N_1828,N_899);
xor U3736 (N_3736,N_1607,N_619);
xor U3737 (N_3737,N_411,N_1289);
nor U3738 (N_3738,N_1559,N_1668);
and U3739 (N_3739,N_1903,N_1521);
nor U3740 (N_3740,N_104,N_702);
nand U3741 (N_3741,N_1436,N_974);
or U3742 (N_3742,N_1744,N_71);
nor U3743 (N_3743,N_1250,N_1159);
or U3744 (N_3744,N_1090,N_1829);
nor U3745 (N_3745,N_60,N_126);
or U3746 (N_3746,N_1262,N_729);
or U3747 (N_3747,N_1141,N_1140);
and U3748 (N_3748,N_1727,N_1167);
and U3749 (N_3749,N_1475,N_1690);
nor U3750 (N_3750,N_1543,N_300);
nor U3751 (N_3751,N_1864,N_981);
nor U3752 (N_3752,N_1254,N_988);
and U3753 (N_3753,N_1308,N_237);
nand U3754 (N_3754,N_1108,N_1198);
nand U3755 (N_3755,N_1200,N_1064);
or U3756 (N_3756,N_1716,N_406);
and U3757 (N_3757,N_1858,N_475);
nor U3758 (N_3758,N_625,N_1352);
nand U3759 (N_3759,N_1732,N_372);
nand U3760 (N_3760,N_369,N_1542);
nor U3761 (N_3761,N_1728,N_268);
and U3762 (N_3762,N_1178,N_889);
nand U3763 (N_3763,N_1737,N_368);
nor U3764 (N_3764,N_482,N_1030);
and U3765 (N_3765,N_1228,N_1216);
nor U3766 (N_3766,N_1922,N_1811);
and U3767 (N_3767,N_1943,N_1890);
and U3768 (N_3768,N_1543,N_628);
or U3769 (N_3769,N_1339,N_1294);
nor U3770 (N_3770,N_1426,N_244);
nor U3771 (N_3771,N_1577,N_162);
xor U3772 (N_3772,N_1705,N_841);
and U3773 (N_3773,N_235,N_1889);
nor U3774 (N_3774,N_1290,N_157);
or U3775 (N_3775,N_1721,N_1809);
or U3776 (N_3776,N_964,N_1945);
nand U3777 (N_3777,N_947,N_448);
and U3778 (N_3778,N_1604,N_156);
or U3779 (N_3779,N_588,N_144);
and U3780 (N_3780,N_1645,N_1592);
nor U3781 (N_3781,N_64,N_614);
and U3782 (N_3782,N_858,N_1567);
and U3783 (N_3783,N_528,N_1273);
nor U3784 (N_3784,N_696,N_1787);
and U3785 (N_3785,N_1443,N_313);
xnor U3786 (N_3786,N_1559,N_343);
or U3787 (N_3787,N_1955,N_1773);
xor U3788 (N_3788,N_398,N_208);
or U3789 (N_3789,N_700,N_739);
nand U3790 (N_3790,N_703,N_876);
xor U3791 (N_3791,N_1300,N_149);
xnor U3792 (N_3792,N_1023,N_582);
and U3793 (N_3793,N_1302,N_408);
nor U3794 (N_3794,N_1164,N_1795);
nand U3795 (N_3795,N_1374,N_424);
or U3796 (N_3796,N_875,N_854);
nand U3797 (N_3797,N_1807,N_1363);
nand U3798 (N_3798,N_1089,N_1299);
or U3799 (N_3799,N_1293,N_1849);
or U3800 (N_3800,N_549,N_1502);
and U3801 (N_3801,N_439,N_56);
or U3802 (N_3802,N_371,N_988);
or U3803 (N_3803,N_1126,N_51);
or U3804 (N_3804,N_1811,N_406);
nand U3805 (N_3805,N_139,N_785);
or U3806 (N_3806,N_1980,N_1215);
or U3807 (N_3807,N_1198,N_662);
xnor U3808 (N_3808,N_650,N_49);
or U3809 (N_3809,N_329,N_1311);
or U3810 (N_3810,N_227,N_1200);
xnor U3811 (N_3811,N_597,N_1420);
nand U3812 (N_3812,N_1944,N_291);
xnor U3813 (N_3813,N_938,N_1871);
nor U3814 (N_3814,N_1379,N_1667);
nor U3815 (N_3815,N_157,N_1630);
nand U3816 (N_3816,N_1504,N_1304);
or U3817 (N_3817,N_869,N_906);
or U3818 (N_3818,N_478,N_888);
nor U3819 (N_3819,N_1080,N_1914);
nand U3820 (N_3820,N_1963,N_1929);
nor U3821 (N_3821,N_1901,N_1771);
and U3822 (N_3822,N_1716,N_1911);
nor U3823 (N_3823,N_1842,N_1783);
nor U3824 (N_3824,N_404,N_225);
or U3825 (N_3825,N_539,N_756);
and U3826 (N_3826,N_101,N_1173);
nand U3827 (N_3827,N_247,N_246);
and U3828 (N_3828,N_1260,N_139);
or U3829 (N_3829,N_1861,N_221);
nor U3830 (N_3830,N_1735,N_806);
xnor U3831 (N_3831,N_1702,N_1435);
nand U3832 (N_3832,N_752,N_577);
or U3833 (N_3833,N_64,N_292);
nor U3834 (N_3834,N_1680,N_624);
and U3835 (N_3835,N_612,N_1747);
and U3836 (N_3836,N_111,N_1298);
nor U3837 (N_3837,N_601,N_84);
nand U3838 (N_3838,N_1609,N_684);
or U3839 (N_3839,N_1505,N_1725);
nor U3840 (N_3840,N_582,N_388);
or U3841 (N_3841,N_411,N_907);
or U3842 (N_3842,N_337,N_131);
or U3843 (N_3843,N_300,N_571);
or U3844 (N_3844,N_1726,N_1730);
xor U3845 (N_3845,N_1841,N_1417);
and U3846 (N_3846,N_1445,N_714);
nor U3847 (N_3847,N_1336,N_1171);
nor U3848 (N_3848,N_898,N_5);
or U3849 (N_3849,N_976,N_1706);
nand U3850 (N_3850,N_355,N_1349);
nand U3851 (N_3851,N_1368,N_1605);
or U3852 (N_3852,N_313,N_639);
nand U3853 (N_3853,N_1641,N_93);
or U3854 (N_3854,N_324,N_1178);
nand U3855 (N_3855,N_459,N_784);
and U3856 (N_3856,N_825,N_1692);
nor U3857 (N_3857,N_740,N_45);
or U3858 (N_3858,N_1642,N_375);
and U3859 (N_3859,N_321,N_1260);
and U3860 (N_3860,N_1067,N_1707);
xnor U3861 (N_3861,N_633,N_1320);
nand U3862 (N_3862,N_1935,N_442);
or U3863 (N_3863,N_896,N_1967);
or U3864 (N_3864,N_736,N_1879);
xor U3865 (N_3865,N_1333,N_375);
and U3866 (N_3866,N_687,N_496);
nand U3867 (N_3867,N_1096,N_1796);
or U3868 (N_3868,N_625,N_742);
nand U3869 (N_3869,N_655,N_390);
or U3870 (N_3870,N_687,N_860);
xor U3871 (N_3871,N_756,N_149);
nor U3872 (N_3872,N_1593,N_83);
and U3873 (N_3873,N_1514,N_1817);
xor U3874 (N_3874,N_636,N_1827);
nand U3875 (N_3875,N_910,N_874);
xnor U3876 (N_3876,N_208,N_1119);
nor U3877 (N_3877,N_1371,N_373);
nor U3878 (N_3878,N_668,N_1806);
and U3879 (N_3879,N_1567,N_854);
or U3880 (N_3880,N_1115,N_902);
nor U3881 (N_3881,N_156,N_1404);
or U3882 (N_3882,N_158,N_873);
nand U3883 (N_3883,N_1433,N_245);
or U3884 (N_3884,N_1294,N_1747);
nor U3885 (N_3885,N_719,N_1525);
nor U3886 (N_3886,N_1190,N_1684);
nand U3887 (N_3887,N_317,N_527);
and U3888 (N_3888,N_932,N_830);
nor U3889 (N_3889,N_190,N_1321);
or U3890 (N_3890,N_805,N_39);
or U3891 (N_3891,N_1658,N_575);
xor U3892 (N_3892,N_490,N_950);
or U3893 (N_3893,N_87,N_503);
nand U3894 (N_3894,N_1280,N_1555);
and U3895 (N_3895,N_466,N_1565);
or U3896 (N_3896,N_1106,N_1178);
nor U3897 (N_3897,N_1943,N_1412);
nand U3898 (N_3898,N_479,N_1369);
xor U3899 (N_3899,N_1170,N_1629);
nand U3900 (N_3900,N_743,N_882);
nand U3901 (N_3901,N_332,N_985);
and U3902 (N_3902,N_1207,N_1491);
nand U3903 (N_3903,N_394,N_556);
or U3904 (N_3904,N_1028,N_450);
or U3905 (N_3905,N_1287,N_6);
and U3906 (N_3906,N_1746,N_1876);
nand U3907 (N_3907,N_1944,N_1450);
xnor U3908 (N_3908,N_1476,N_1735);
or U3909 (N_3909,N_1309,N_111);
and U3910 (N_3910,N_670,N_1381);
and U3911 (N_3911,N_556,N_849);
nand U3912 (N_3912,N_1186,N_1043);
and U3913 (N_3913,N_1744,N_233);
nand U3914 (N_3914,N_767,N_753);
and U3915 (N_3915,N_542,N_1240);
and U3916 (N_3916,N_1654,N_59);
nand U3917 (N_3917,N_593,N_970);
nand U3918 (N_3918,N_310,N_1521);
or U3919 (N_3919,N_52,N_378);
xor U3920 (N_3920,N_469,N_1881);
and U3921 (N_3921,N_1046,N_566);
xor U3922 (N_3922,N_907,N_420);
or U3923 (N_3923,N_1827,N_43);
xor U3924 (N_3924,N_1285,N_1257);
nand U3925 (N_3925,N_985,N_852);
nor U3926 (N_3926,N_789,N_742);
xnor U3927 (N_3927,N_496,N_114);
and U3928 (N_3928,N_1376,N_1349);
nand U3929 (N_3929,N_1130,N_886);
and U3930 (N_3930,N_640,N_192);
nor U3931 (N_3931,N_1832,N_1681);
nand U3932 (N_3932,N_184,N_1091);
xor U3933 (N_3933,N_1898,N_1156);
nor U3934 (N_3934,N_417,N_967);
nor U3935 (N_3935,N_1581,N_1673);
and U3936 (N_3936,N_1170,N_630);
or U3937 (N_3937,N_197,N_742);
xor U3938 (N_3938,N_834,N_774);
nor U3939 (N_3939,N_966,N_1894);
nor U3940 (N_3940,N_1103,N_970);
or U3941 (N_3941,N_91,N_1125);
nor U3942 (N_3942,N_544,N_1611);
xnor U3943 (N_3943,N_1807,N_1531);
nor U3944 (N_3944,N_1114,N_337);
or U3945 (N_3945,N_8,N_258);
and U3946 (N_3946,N_1262,N_1022);
nor U3947 (N_3947,N_29,N_828);
nor U3948 (N_3948,N_602,N_435);
xor U3949 (N_3949,N_727,N_1446);
and U3950 (N_3950,N_331,N_765);
nand U3951 (N_3951,N_110,N_1662);
or U3952 (N_3952,N_934,N_564);
and U3953 (N_3953,N_18,N_1992);
and U3954 (N_3954,N_275,N_1705);
or U3955 (N_3955,N_259,N_1046);
and U3956 (N_3956,N_1841,N_536);
or U3957 (N_3957,N_406,N_1618);
xor U3958 (N_3958,N_1129,N_1866);
nand U3959 (N_3959,N_845,N_1347);
xor U3960 (N_3960,N_1485,N_1950);
or U3961 (N_3961,N_731,N_1010);
xor U3962 (N_3962,N_1054,N_1919);
or U3963 (N_3963,N_825,N_767);
xnor U3964 (N_3964,N_607,N_1082);
and U3965 (N_3965,N_173,N_1701);
and U3966 (N_3966,N_1013,N_581);
nand U3967 (N_3967,N_798,N_1031);
or U3968 (N_3968,N_429,N_1010);
or U3969 (N_3969,N_474,N_114);
nand U3970 (N_3970,N_982,N_1294);
or U3971 (N_3971,N_422,N_1666);
or U3972 (N_3972,N_398,N_1492);
nor U3973 (N_3973,N_999,N_277);
or U3974 (N_3974,N_835,N_1560);
nand U3975 (N_3975,N_1082,N_290);
or U3976 (N_3976,N_1025,N_1933);
or U3977 (N_3977,N_1010,N_161);
nand U3978 (N_3978,N_331,N_1306);
nor U3979 (N_3979,N_172,N_1319);
or U3980 (N_3980,N_497,N_1604);
and U3981 (N_3981,N_1365,N_590);
xor U3982 (N_3982,N_956,N_1964);
nand U3983 (N_3983,N_738,N_154);
or U3984 (N_3984,N_1328,N_634);
or U3985 (N_3985,N_668,N_225);
nor U3986 (N_3986,N_534,N_9);
nor U3987 (N_3987,N_845,N_1624);
xor U3988 (N_3988,N_1316,N_713);
nor U3989 (N_3989,N_1000,N_157);
nand U3990 (N_3990,N_897,N_1058);
and U3991 (N_3991,N_50,N_974);
nand U3992 (N_3992,N_948,N_1817);
and U3993 (N_3993,N_1828,N_593);
xnor U3994 (N_3994,N_841,N_1848);
and U3995 (N_3995,N_1913,N_1625);
and U3996 (N_3996,N_1437,N_1688);
or U3997 (N_3997,N_1339,N_788);
or U3998 (N_3998,N_1570,N_1130);
and U3999 (N_3999,N_320,N_12);
nor U4000 (N_4000,N_3314,N_2982);
or U4001 (N_4001,N_3776,N_2182);
and U4002 (N_4002,N_2050,N_3426);
and U4003 (N_4003,N_2996,N_2181);
nor U4004 (N_4004,N_3485,N_2142);
and U4005 (N_4005,N_2700,N_3040);
and U4006 (N_4006,N_2397,N_2192);
nor U4007 (N_4007,N_2878,N_2458);
nand U4008 (N_4008,N_3510,N_2058);
nor U4009 (N_4009,N_2619,N_3604);
nand U4010 (N_4010,N_2510,N_3172);
nand U4011 (N_4011,N_2798,N_3247);
nand U4012 (N_4012,N_3428,N_3998);
or U4013 (N_4013,N_3458,N_2896);
or U4014 (N_4014,N_2566,N_3561);
nor U4015 (N_4015,N_2825,N_2621);
xor U4016 (N_4016,N_3061,N_2833);
nand U4017 (N_4017,N_3204,N_3914);
nor U4018 (N_4018,N_2446,N_3448);
nor U4019 (N_4019,N_3926,N_3438);
and U4020 (N_4020,N_3697,N_3892);
and U4021 (N_4021,N_2095,N_3372);
nor U4022 (N_4022,N_2012,N_2416);
nor U4023 (N_4023,N_3359,N_2722);
xor U4024 (N_4024,N_3009,N_3355);
and U4025 (N_4025,N_3780,N_3553);
and U4026 (N_4026,N_3851,N_2190);
or U4027 (N_4027,N_3154,N_3045);
and U4028 (N_4028,N_2369,N_2539);
or U4029 (N_4029,N_2728,N_2334);
nand U4030 (N_4030,N_2780,N_3170);
xor U4031 (N_4031,N_2927,N_2959);
xnor U4032 (N_4032,N_2752,N_2315);
nand U4033 (N_4033,N_3232,N_3261);
xor U4034 (N_4034,N_3612,N_2212);
nand U4035 (N_4035,N_3953,N_2158);
or U4036 (N_4036,N_2877,N_3498);
nand U4037 (N_4037,N_2561,N_3843);
nor U4038 (N_4038,N_3169,N_2456);
nand U4039 (N_4039,N_3677,N_2802);
and U4040 (N_4040,N_3205,N_3797);
nor U4041 (N_4041,N_2884,N_3992);
nor U4042 (N_4042,N_3416,N_2588);
nand U4043 (N_4043,N_3222,N_3410);
or U4044 (N_4044,N_2267,N_2357);
or U4045 (N_4045,N_3971,N_3296);
nand U4046 (N_4046,N_2628,N_3579);
xor U4047 (N_4047,N_3075,N_3814);
xnor U4048 (N_4048,N_2252,N_3996);
or U4049 (N_4049,N_3624,N_3645);
and U4050 (N_4050,N_2944,N_3546);
or U4051 (N_4051,N_3837,N_2506);
and U4052 (N_4052,N_3093,N_3309);
nand U4053 (N_4053,N_2596,N_3186);
and U4054 (N_4054,N_2302,N_2536);
nand U4055 (N_4055,N_3351,N_2550);
or U4056 (N_4056,N_2143,N_3119);
nor U4057 (N_4057,N_2209,N_2865);
or U4058 (N_4058,N_3409,N_3921);
nor U4059 (N_4059,N_3631,N_2739);
and U4060 (N_4060,N_3421,N_3668);
or U4061 (N_4061,N_3722,N_2041);
or U4062 (N_4062,N_2636,N_3108);
nor U4063 (N_4063,N_3275,N_3392);
nor U4064 (N_4064,N_3103,N_2680);
and U4065 (N_4065,N_2056,N_2104);
xor U4066 (N_4066,N_3126,N_3765);
or U4067 (N_4067,N_2652,N_2358);
or U4068 (N_4068,N_2476,N_2605);
xor U4069 (N_4069,N_2467,N_2692);
and U4070 (N_4070,N_3331,N_2101);
and U4071 (N_4071,N_2303,N_2053);
xnor U4072 (N_4072,N_2795,N_2805);
nor U4073 (N_4073,N_3411,N_2349);
and U4074 (N_4074,N_3975,N_3181);
or U4075 (N_4075,N_2885,N_3603);
nand U4076 (N_4076,N_2340,N_2451);
or U4077 (N_4077,N_3818,N_3384);
or U4078 (N_4078,N_2293,N_2284);
or U4079 (N_4079,N_2983,N_3095);
or U4080 (N_4080,N_3618,N_3489);
and U4081 (N_4081,N_3539,N_2732);
xor U4082 (N_4082,N_3071,N_2200);
nor U4083 (N_4083,N_2077,N_3511);
nor U4084 (N_4084,N_2162,N_3019);
nand U4085 (N_4085,N_2133,N_3446);
nand U4086 (N_4086,N_2455,N_3667);
nand U4087 (N_4087,N_2491,N_2689);
and U4088 (N_4088,N_3687,N_2970);
and U4089 (N_4089,N_3209,N_3642);
xnor U4090 (N_4090,N_2583,N_2705);
nor U4091 (N_4091,N_2609,N_3820);
and U4092 (N_4092,N_2201,N_3889);
and U4093 (N_4093,N_2666,N_2599);
nand U4094 (N_4094,N_3969,N_2319);
xnor U4095 (N_4095,N_3400,N_2193);
or U4096 (N_4096,N_3349,N_2215);
and U4097 (N_4097,N_2102,N_3863);
or U4098 (N_4098,N_3110,N_3012);
nand U4099 (N_4099,N_2263,N_2850);
nand U4100 (N_4100,N_2399,N_2727);
nand U4101 (N_4101,N_3880,N_3360);
xor U4102 (N_4102,N_3724,N_2164);
nand U4103 (N_4103,N_3823,N_2714);
nand U4104 (N_4104,N_2866,N_2024);
nand U4105 (N_4105,N_2000,N_3982);
nand U4106 (N_4106,N_2625,N_3390);
nand U4107 (N_4107,N_2396,N_3799);
nand U4108 (N_4108,N_3201,N_3419);
nand U4109 (N_4109,N_3492,N_2317);
or U4110 (N_4110,N_2560,N_3264);
or U4111 (N_4111,N_2063,N_2634);
xor U4112 (N_4112,N_3871,N_2381);
or U4113 (N_4113,N_2097,N_3237);
nand U4114 (N_4114,N_2065,N_2137);
and U4115 (N_4115,N_3676,N_3699);
or U4116 (N_4116,N_3449,N_2330);
and U4117 (N_4117,N_3445,N_3918);
or U4118 (N_4118,N_2901,N_2250);
or U4119 (N_4119,N_3568,N_3565);
nand U4120 (N_4120,N_3938,N_2236);
xor U4121 (N_4121,N_2864,N_3875);
and U4122 (N_4122,N_2367,N_2219);
or U4123 (N_4123,N_3405,N_2743);
nand U4124 (N_4124,N_3233,N_2829);
or U4125 (N_4125,N_2568,N_2995);
or U4126 (N_4126,N_2635,N_2696);
nor U4127 (N_4127,N_2136,N_3277);
and U4128 (N_4128,N_3842,N_2059);
nand U4129 (N_4129,N_3589,N_2907);
xnor U4130 (N_4130,N_3235,N_2016);
nand U4131 (N_4131,N_3328,N_2614);
nor U4132 (N_4132,N_3902,N_2574);
and U4133 (N_4133,N_3096,N_2213);
nand U4134 (N_4134,N_3712,N_2346);
and U4135 (N_4135,N_3435,N_2486);
nor U4136 (N_4136,N_2520,N_2036);
xor U4137 (N_4137,N_2487,N_2433);
and U4138 (N_4138,N_3022,N_3109);
xor U4139 (N_4139,N_3753,N_3690);
nor U4140 (N_4140,N_2546,N_2003);
nor U4141 (N_4141,N_3081,N_3148);
or U4142 (N_4142,N_3933,N_3620);
nand U4143 (N_4143,N_2713,N_3861);
and U4144 (N_4144,N_2135,N_2686);
nor U4145 (N_4145,N_2814,N_2817);
xor U4146 (N_4146,N_2529,N_2662);
nand U4147 (N_4147,N_2572,N_2088);
nand U4148 (N_4148,N_3904,N_3771);
nor U4149 (N_4149,N_3060,N_2270);
nor U4150 (N_4150,N_3911,N_2894);
nand U4151 (N_4151,N_3475,N_3260);
and U4152 (N_4152,N_3361,N_2475);
xnor U4153 (N_4153,N_3466,N_3027);
nand U4154 (N_4154,N_3422,N_2023);
or U4155 (N_4155,N_3900,N_2961);
or U4156 (N_4156,N_2757,N_3582);
nand U4157 (N_4157,N_2177,N_2457);
or U4158 (N_4158,N_3218,N_3132);
nand U4159 (N_4159,N_2241,N_3014);
or U4160 (N_4160,N_2807,N_2993);
or U4161 (N_4161,N_2134,N_2294);
nor U4162 (N_4162,N_2984,N_2637);
xnor U4163 (N_4163,N_2698,N_3125);
and U4164 (N_4164,N_3718,N_3176);
nor U4165 (N_4165,N_2488,N_2060);
nand U4166 (N_4166,N_2300,N_3810);
and U4167 (N_4167,N_3236,N_2904);
xor U4168 (N_4168,N_2248,N_3318);
and U4169 (N_4169,N_2482,N_2266);
xor U4170 (N_4170,N_3393,N_2049);
or U4171 (N_4171,N_3369,N_3255);
or U4172 (N_4172,N_3219,N_3559);
nand U4173 (N_4173,N_3964,N_2590);
nand U4174 (N_4174,N_2554,N_3436);
nand U4175 (N_4175,N_3433,N_3832);
and U4176 (N_4176,N_2015,N_3520);
and U4177 (N_4177,N_3386,N_3594);
nor U4178 (N_4178,N_2924,N_2132);
and U4179 (N_4179,N_2292,N_3388);
and U4180 (N_4180,N_2775,N_2075);
and U4181 (N_4181,N_2933,N_2103);
or U4182 (N_4182,N_2830,N_2191);
and U4183 (N_4183,N_3816,N_2377);
xnor U4184 (N_4184,N_2110,N_3544);
or U4185 (N_4185,N_3437,N_2453);
and U4186 (N_4186,N_3171,N_2564);
nand U4187 (N_4187,N_2495,N_3610);
nand U4188 (N_4188,N_3703,N_2542);
nand U4189 (N_4189,N_3532,N_2563);
nand U4190 (N_4190,N_3827,N_3290);
nand U4191 (N_4191,N_2912,N_3663);
nand U4192 (N_4192,N_2932,N_3836);
nand U4193 (N_4193,N_3379,N_3795);
and U4194 (N_4194,N_2187,N_3270);
nor U4195 (N_4195,N_3143,N_2659);
xnor U4196 (N_4196,N_3202,N_2310);
xnor U4197 (N_4197,N_3876,N_3666);
or U4198 (N_4198,N_2422,N_2582);
nand U4199 (N_4199,N_2972,N_3670);
nand U4200 (N_4200,N_2316,N_2950);
nor U4201 (N_4201,N_2279,N_2255);
nand U4202 (N_4202,N_3640,N_2514);
or U4203 (N_4203,N_2028,N_3671);
and U4204 (N_4204,N_2083,N_2928);
nand U4205 (N_4205,N_3688,N_3145);
nor U4206 (N_4206,N_3987,N_3635);
xnor U4207 (N_4207,N_2172,N_2038);
nand U4208 (N_4208,N_3212,N_3175);
and U4209 (N_4209,N_2955,N_3330);
nor U4210 (N_4210,N_3121,N_3210);
xor U4211 (N_4211,N_3809,N_2818);
and U4212 (N_4212,N_3129,N_2918);
nand U4213 (N_4213,N_3211,N_3897);
nor U4214 (N_4214,N_3128,N_3800);
and U4215 (N_4215,N_3363,N_2111);
nor U4216 (N_4216,N_2759,N_2139);
xor U4217 (N_4217,N_3463,N_3808);
xnor U4218 (N_4218,N_2513,N_3960);
and U4219 (N_4219,N_2222,N_2871);
and U4220 (N_4220,N_3244,N_3710);
xor U4221 (N_4221,N_3378,N_3794);
nor U4222 (N_4222,N_2493,N_3404);
nand U4223 (N_4223,N_3460,N_2793);
nor U4224 (N_4224,N_2500,N_2677);
nand U4225 (N_4225,N_2120,N_2008);
nand U4226 (N_4226,N_2740,N_2979);
xor U4227 (N_4227,N_2254,N_3398);
nand U4228 (N_4228,N_3890,N_3069);
or U4229 (N_4229,N_3408,N_3841);
nor U4230 (N_4230,N_3134,N_3862);
nand U4231 (N_4231,N_2203,N_3333);
and U4232 (N_4232,N_2916,N_3420);
nor U4233 (N_4233,N_3826,N_2948);
nor U4234 (N_4234,N_2791,N_2708);
nor U4235 (N_4235,N_3374,N_2468);
or U4236 (N_4236,N_2234,N_3548);
and U4237 (N_4237,N_3227,N_2390);
or U4238 (N_4238,N_3705,N_2768);
nor U4239 (N_4239,N_2283,N_2719);
or U4240 (N_4240,N_3316,N_2820);
xnor U4241 (N_4241,N_3590,N_3158);
nand U4242 (N_4242,N_2039,N_2523);
or U4243 (N_4243,N_3630,N_2718);
nor U4244 (N_4244,N_3401,N_2681);
and U4245 (N_4245,N_2858,N_3951);
or U4246 (N_4246,N_2249,N_3326);
nand U4247 (N_4247,N_2951,N_3927);
nor U4248 (N_4248,N_2755,N_3908);
nand U4249 (N_4249,N_2031,N_3324);
or U4250 (N_4250,N_2620,N_2314);
or U4251 (N_4251,N_3523,N_3763);
or U4252 (N_4252,N_3573,N_2055);
nor U4253 (N_4253,N_3343,N_3097);
nor U4254 (N_4254,N_2400,N_3732);
or U4255 (N_4255,N_3530,N_3003);
nor U4256 (N_4256,N_3241,N_3519);
or U4257 (N_4257,N_2785,N_2675);
nand U4258 (N_4258,N_3284,N_2325);
and U4259 (N_4259,N_3524,N_2153);
nor U4260 (N_4260,N_2908,N_2929);
nand U4261 (N_4261,N_2240,N_3606);
xor U4262 (N_4262,N_2555,N_2812);
nand U4263 (N_4263,N_3111,N_3266);
or U4264 (N_4264,N_3439,N_2244);
xnor U4265 (N_4265,N_3067,N_3706);
nor U4266 (N_4266,N_2037,N_3660);
nor U4267 (N_4267,N_2227,N_2697);
nand U4268 (N_4268,N_2168,N_3016);
xnor U4269 (N_4269,N_3829,N_2471);
and U4270 (N_4270,N_3689,N_2741);
nor U4271 (N_4271,N_3425,N_3483);
or U4272 (N_4272,N_2761,N_2613);
and U4273 (N_4273,N_2532,N_3967);
xor U4274 (N_4274,N_2239,N_2524);
nand U4275 (N_4275,N_3074,N_2969);
nor U4276 (N_4276,N_3461,N_3293);
and U4277 (N_4277,N_2366,N_2099);
nand U4278 (N_4278,N_2264,N_2873);
or U4279 (N_4279,N_2849,N_2515);
xor U4280 (N_4280,N_2074,N_2521);
and U4281 (N_4281,N_2337,N_3955);
nand U4282 (N_4282,N_2886,N_3570);
nor U4283 (N_4283,N_3160,N_3038);
or U4284 (N_4284,N_2224,N_3627);
and U4285 (N_4285,N_3509,N_3299);
and U4286 (N_4286,N_3484,N_2679);
or U4287 (N_4287,N_3680,N_2570);
or U4288 (N_4288,N_3399,N_2956);
nor U4289 (N_4289,N_3010,N_2921);
nor U4290 (N_4290,N_3220,N_3518);
nand U4291 (N_4291,N_2046,N_2274);
nor U4292 (N_4292,N_2454,N_2067);
nand U4293 (N_4293,N_3099,N_2717);
nand U4294 (N_4294,N_3787,N_2939);
xor U4295 (N_4295,N_3298,N_3583);
nand U4296 (N_4296,N_3073,N_2986);
xnor U4297 (N_4297,N_2789,N_3749);
and U4298 (N_4298,N_3634,N_2556);
and U4299 (N_4299,N_3839,N_3123);
or U4300 (N_4300,N_3455,N_3602);
nor U4301 (N_4301,N_2845,N_2895);
nand U4302 (N_4302,N_2130,N_2331);
nor U4303 (N_4303,N_2040,N_3087);
nand U4304 (N_4304,N_3249,N_2832);
xnor U4305 (N_4305,N_2973,N_3543);
and U4306 (N_4306,N_2869,N_2149);
xnor U4307 (N_4307,N_2372,N_3427);
nor U4308 (N_4308,N_3526,N_2558);
nor U4309 (N_4309,N_3265,N_2695);
nor U4310 (N_4310,N_3711,N_3352);
nand U4311 (N_4311,N_3412,N_3114);
nor U4312 (N_4312,N_3286,N_2086);
and U4313 (N_4313,N_3740,N_3494);
and U4314 (N_4314,N_2954,N_3113);
and U4315 (N_4315,N_3868,N_3537);
nor U4316 (N_4316,N_3936,N_2449);
nor U4317 (N_4317,N_2345,N_2971);
or U4318 (N_4318,N_2230,N_3033);
xor U4319 (N_4319,N_3496,N_2257);
nand U4320 (N_4320,N_2112,N_2876);
nand U4321 (N_4321,N_3402,N_3057);
nand U4322 (N_4322,N_2750,N_3654);
nor U4323 (N_4323,N_2301,N_3403);
or U4324 (N_4324,N_3566,N_3869);
nand U4325 (N_4325,N_3536,N_3504);
or U4326 (N_4326,N_2952,N_3153);
and U4327 (N_4327,N_3886,N_2872);
nor U4328 (N_4328,N_3200,N_3848);
or U4329 (N_4329,N_2987,N_3741);
nor U4330 (N_4330,N_3834,N_2290);
nor U4331 (N_4331,N_2577,N_2184);
xnor U4332 (N_4332,N_2010,N_3646);
xor U4333 (N_4333,N_3801,N_3701);
and U4334 (N_4334,N_3824,N_2178);
nand U4335 (N_4335,N_3852,N_3694);
nand U4336 (N_4336,N_2167,N_2375);
or U4337 (N_4337,N_2004,N_2758);
nor U4338 (N_4338,N_3039,N_2512);
and U4339 (N_4339,N_2835,N_2914);
xor U4340 (N_4340,N_2720,N_2949);
nor U4341 (N_4341,N_2547,N_3752);
xor U4342 (N_4342,N_3004,N_3636);
and U4343 (N_4343,N_2808,N_2586);
nand U4344 (N_4344,N_2195,N_2352);
nand U4345 (N_4345,N_3184,N_3609);
xor U4346 (N_4346,N_3919,N_2034);
and U4347 (N_4347,N_2430,N_3207);
or U4348 (N_4348,N_2217,N_3025);
or U4349 (N_4349,N_3195,N_3600);
and U4350 (N_4350,N_2985,N_3613);
nand U4351 (N_4351,N_3507,N_2424);
nand U4352 (N_4352,N_3058,N_3082);
or U4353 (N_4353,N_2682,N_3203);
or U4354 (N_4354,N_2707,N_3441);
nor U4355 (N_4355,N_3116,N_3672);
or U4356 (N_4356,N_2962,N_3807);
nor U4357 (N_4357,N_2045,N_2980);
or U4358 (N_4358,N_3790,N_3424);
and U4359 (N_4359,N_3443,N_2745);
nor U4360 (N_4360,N_3358,N_3342);
or U4361 (N_4361,N_2623,N_2463);
nor U4362 (N_4362,N_2673,N_2839);
or U4363 (N_4363,N_2220,N_2093);
and U4364 (N_4364,N_2734,N_3055);
or U4365 (N_4365,N_3502,N_3118);
nand U4366 (N_4366,N_3135,N_2893);
or U4367 (N_4367,N_2981,N_3675);
nand U4368 (N_4368,N_3858,N_2660);
or U4369 (N_4369,N_2926,N_2612);
nor U4370 (N_4370,N_2883,N_3332);
or U4371 (N_4371,N_2837,N_2607);
nand U4372 (N_4372,N_2108,N_3070);
nand U4373 (N_4373,N_2261,N_3773);
nor U4374 (N_4374,N_3888,N_3246);
or U4375 (N_4375,N_2941,N_3648);
nor U4376 (N_4376,N_2490,N_3870);
nor U4377 (N_4377,N_2528,N_2800);
or U4378 (N_4378,N_3196,N_2942);
xor U4379 (N_4379,N_2070,N_3383);
and U4380 (N_4380,N_3357,N_2756);
or U4381 (N_4381,N_2033,N_2709);
xnor U4382 (N_4382,N_2671,N_2856);
nand U4383 (N_4383,N_3656,N_2790);
nand U4384 (N_4384,N_2199,N_2376);
nor U4385 (N_4385,N_3872,N_3943);
xnor U4386 (N_4386,N_2738,N_2502);
and U4387 (N_4387,N_3551,N_3307);
or U4388 (N_4388,N_2552,N_2185);
nand U4389 (N_4389,N_2062,N_2779);
or U4390 (N_4390,N_2503,N_3812);
or U4391 (N_4391,N_3860,N_3903);
or U4392 (N_4392,N_2988,N_2339);
or U4393 (N_4393,N_3981,N_3447);
xor U4394 (N_4394,N_2383,N_3731);
nor U4395 (N_4395,N_3729,N_2278);
xor U4396 (N_4396,N_2272,N_3101);
nand U4397 (N_4397,N_3853,N_3950);
and U4398 (N_4398,N_2801,N_3702);
nor U4399 (N_4399,N_3695,N_3490);
nor U4400 (N_4400,N_3774,N_2421);
and U4401 (N_4401,N_3089,N_2880);
nand U4402 (N_4402,N_3698,N_3844);
or U4403 (N_4403,N_2144,N_3238);
nand U4404 (N_4404,N_2764,N_2362);
nand U4405 (N_4405,N_2827,N_2898);
xnor U4406 (N_4406,N_3376,N_3213);
and U4407 (N_4407,N_2724,N_2540);
xor U4408 (N_4408,N_2892,N_2351);
nand U4409 (N_4409,N_2426,N_2589);
or U4410 (N_4410,N_3959,N_2138);
nor U4411 (N_4411,N_3757,N_2379);
nor U4412 (N_4412,N_2206,N_2151);
nor U4413 (N_4413,N_2418,N_3542);
nand U4414 (N_4414,N_3477,N_3292);
nor U4415 (N_4415,N_3183,N_2746);
nand U4416 (N_4416,N_3859,N_2013);
or U4417 (N_4417,N_2485,N_3616);
nor U4418 (N_4418,N_3174,N_3345);
and U4419 (N_4419,N_3065,N_3760);
nand U4420 (N_4420,N_2459,N_2911);
or U4421 (N_4421,N_2784,N_2079);
nand U4422 (N_4422,N_3337,N_3772);
nand U4423 (N_4423,N_3893,N_2836);
nand U4424 (N_4424,N_2440,N_3652);
or U4425 (N_4425,N_2654,N_3930);
nor U4426 (N_4426,N_3444,N_3821);
nand U4427 (N_4427,N_3017,N_3641);
nor U4428 (N_4428,N_3623,N_2176);
nand U4429 (N_4429,N_2196,N_3362);
nand U4430 (N_4430,N_2100,N_2022);
or U4431 (N_4431,N_2647,N_3397);
or U4432 (N_4432,N_3916,N_3693);
or U4433 (N_4433,N_2910,N_2018);
and U4434 (N_4434,N_2753,N_2683);
nand U4435 (N_4435,N_2649,N_2518);
nand U4436 (N_4436,N_2991,N_2179);
or U4437 (N_4437,N_3857,N_2762);
or U4438 (N_4438,N_3966,N_2810);
and U4439 (N_4439,N_3122,N_2668);
or U4440 (N_4440,N_3056,N_3550);
nor U4441 (N_4441,N_3736,N_3560);
and U4442 (N_4442,N_3091,N_3271);
xnor U4443 (N_4443,N_2963,N_3350);
nor U4444 (N_4444,N_2147,N_2676);
nand U4445 (N_4445,N_3997,N_2428);
or U4446 (N_4446,N_2006,N_3149);
xnor U4447 (N_4447,N_2145,N_3467);
nand U4448 (N_4448,N_2945,N_2389);
nand U4449 (N_4449,N_2822,N_3669);
or U4450 (N_4450,N_3323,N_2262);
or U4451 (N_4451,N_2776,N_2990);
or U4452 (N_4452,N_2615,N_3529);
nor U4453 (N_4453,N_3375,N_3214);
and U4454 (N_4454,N_2452,N_2842);
nand U4455 (N_4455,N_2541,N_3983);
nand U4456 (N_4456,N_2846,N_2285);
and U4457 (N_4457,N_3086,N_3051);
xnor U4458 (N_4458,N_2571,N_2651);
nor U4459 (N_4459,N_2868,N_3533);
nor U4460 (N_4460,N_3856,N_2477);
or U4461 (N_4461,N_3482,N_2348);
nand U4462 (N_4462,N_2297,N_2678);
nand U4463 (N_4463,N_3018,N_3381);
and U4464 (N_4464,N_2656,N_2843);
xor U4465 (N_4465,N_3304,N_2295);
nor U4466 (N_4466,N_2098,N_3514);
and U4467 (N_4467,N_3973,N_3341);
or U4468 (N_4468,N_2125,N_3313);
nand U4469 (N_4469,N_2394,N_2338);
and U4470 (N_4470,N_2976,N_3257);
xor U4471 (N_4471,N_2188,N_2595);
and U4472 (N_4472,N_2573,N_3571);
nand U4473 (N_4473,N_2639,N_3294);
nor U4474 (N_4474,N_2913,N_3217);
or U4475 (N_4475,N_3394,N_2298);
nand U4476 (N_4476,N_3804,N_3562);
and U4477 (N_4477,N_3054,N_2464);
or U4478 (N_4478,N_3961,N_2385);
nor U4479 (N_4479,N_3197,N_2860);
nand U4480 (N_4480,N_3758,N_3845);
nor U4481 (N_4481,N_3995,N_2169);
or U4482 (N_4482,N_3230,N_2781);
nor U4483 (N_4483,N_3479,N_2494);
and U4484 (N_4484,N_3474,N_2854);
and U4485 (N_4485,N_3389,N_2470);
or U4486 (N_4486,N_3288,N_2225);
nand U4487 (N_4487,N_3013,N_2043);
or U4488 (N_4488,N_3920,N_3180);
nand U4489 (N_4489,N_2531,N_2005);
nand U4490 (N_4490,N_2327,N_3813);
nand U4491 (N_4491,N_2862,N_3896);
and U4492 (N_4492,N_2797,N_3500);
or U4493 (N_4493,N_2173,N_3803);
or U4494 (N_4494,N_2092,N_3976);
or U4495 (N_4495,N_3162,N_3308);
xor U4496 (N_4496,N_3782,N_2189);
or U4497 (N_4497,N_2882,N_2794);
nand U4498 (N_4498,N_2344,N_3486);
nor U4499 (N_4499,N_3882,N_3569);
nor U4500 (N_4500,N_3878,N_2958);
xor U4501 (N_4501,N_2553,N_3598);
and U4502 (N_4502,N_3643,N_3759);
nor U4503 (N_4503,N_3686,N_2154);
and U4504 (N_4504,N_3280,N_2604);
nand U4505 (N_4505,N_2242,N_3506);
or U4506 (N_4506,N_3164,N_2533);
and U4507 (N_4507,N_3556,N_3413);
or U4508 (N_4508,N_3683,N_3182);
nor U4509 (N_4509,N_2118,N_3064);
or U4510 (N_4510,N_2824,N_3193);
xor U4511 (N_4511,N_3415,N_2505);
nor U4512 (N_4512,N_2165,N_2131);
and U4513 (N_4513,N_2624,N_3028);
nor U4514 (N_4514,N_2081,N_3855);
nor U4515 (N_4515,N_2064,N_3587);
and U4516 (N_4516,N_3768,N_2978);
and U4517 (N_4517,N_3516,N_2559);
or U4518 (N_4518,N_2940,N_3707);
or U4519 (N_4519,N_2296,N_3098);
nor U4520 (N_4520,N_2313,N_2047);
and U4521 (N_4521,N_2627,N_2852);
nor U4522 (N_4522,N_2057,N_3100);
nand U4523 (N_4523,N_2492,N_3440);
nand U4524 (N_4524,N_2321,N_3873);
nor U4525 (N_4525,N_2919,N_3713);
and U4526 (N_4526,N_3717,N_2966);
nand U4527 (N_4527,N_3796,N_2078);
or U4528 (N_4528,N_3285,N_2277);
or U4529 (N_4529,N_3334,N_3188);
or U4530 (N_4530,N_2140,N_3117);
nor U4531 (N_4531,N_3090,N_3312);
nand U4532 (N_4532,N_3198,N_2684);
and U4533 (N_4533,N_3747,N_2522);
xor U4534 (N_4534,N_2909,N_3572);
or U4535 (N_4535,N_3545,N_2460);
and U4536 (N_4536,N_3945,N_2026);
and U4537 (N_4537,N_3811,N_3946);
or U4538 (N_4538,N_3262,N_2054);
and U4539 (N_4539,N_2694,N_2126);
xor U4540 (N_4540,N_2186,N_2508);
or U4541 (N_4541,N_2875,N_2268);
nor U4542 (N_4542,N_3066,N_2364);
nand U4543 (N_4543,N_2419,N_3044);
or U4544 (N_4544,N_3306,N_3301);
and U4545 (N_4545,N_3788,N_2388);
xnor U4546 (N_4546,N_3231,N_2243);
nand U4547 (N_4547,N_2544,N_2930);
nand U4548 (N_4548,N_3963,N_2071);
nor U4549 (N_4549,N_3840,N_2899);
nor U4550 (N_4550,N_3748,N_2957);
nor U4551 (N_4551,N_2777,N_2967);
or U4552 (N_4552,N_2427,N_3470);
or U4553 (N_4553,N_2716,N_2404);
and U4554 (N_4554,N_3727,N_2391);
xor U4555 (N_4555,N_3558,N_3283);
nor U4556 (N_4556,N_2496,N_2943);
and U4557 (N_4557,N_3737,N_3248);
nand U4558 (N_4558,N_2584,N_3791);
or U4559 (N_4559,N_3456,N_2778);
xnor U4560 (N_4560,N_2343,N_2448);
nor U4561 (N_4561,N_3939,N_3273);
nor U4562 (N_4562,N_2436,N_2934);
or U4563 (N_4563,N_3607,N_2823);
nor U4564 (N_4564,N_3226,N_2197);
or U4565 (N_4565,N_2174,N_3320);
and U4566 (N_4566,N_3085,N_2403);
nor U4567 (N_4567,N_2735,N_2194);
nand U4568 (N_4568,N_3274,N_3608);
or U4569 (N_4569,N_3901,N_2897);
nand U4570 (N_4570,N_3166,N_2922);
or U4571 (N_4571,N_2114,N_2598);
or U4572 (N_4572,N_2373,N_2017);
nor U4573 (N_4573,N_2307,N_2259);
xor U4574 (N_4574,N_2549,N_2483);
xnor U4575 (N_4575,N_3835,N_3784);
nand U4576 (N_4576,N_3254,N_2640);
nor U4577 (N_4577,N_3977,N_2937);
and U4578 (N_4578,N_2906,N_3289);
or U4579 (N_4579,N_2170,N_2392);
xnor U4580 (N_4580,N_3021,N_3147);
and U4581 (N_4581,N_2335,N_3250);
and U4582 (N_4582,N_3726,N_3777);
nand U4583 (N_4583,N_3442,N_3999);
nand U4584 (N_4584,N_3347,N_3517);
nand U4585 (N_4585,N_3619,N_3682);
or U4586 (N_4586,N_2311,N_2674);
or U4587 (N_4587,N_3150,N_2107);
or U4588 (N_4588,N_3989,N_3317);
or U4589 (N_4589,N_2594,N_2851);
or U4590 (N_4590,N_3637,N_3647);
or U4591 (N_4591,N_2076,N_3315);
nor U4592 (N_4592,N_3673,N_2214);
nand U4593 (N_4593,N_3026,N_3850);
and U4594 (N_4594,N_3465,N_2626);
nor U4595 (N_4595,N_3761,N_2511);
or U4596 (N_4596,N_2269,N_3922);
nand U4597 (N_4597,N_2538,N_2387);
and U4598 (N_4598,N_2857,N_3281);
and U4599 (N_4599,N_3704,N_3535);
or U4600 (N_4600,N_3503,N_2417);
or U4601 (N_4601,N_3423,N_3015);
nor U4602 (N_4602,N_3036,N_2226);
nor U4603 (N_4603,N_2663,N_3168);
and U4604 (N_4604,N_3105,N_2336);
and U4605 (N_4605,N_2831,N_3001);
and U4606 (N_4606,N_3581,N_3785);
nor U4607 (N_4607,N_2998,N_2509);
or U4608 (N_4608,N_3563,N_3335);
and U4609 (N_4609,N_2657,N_3653);
and U4610 (N_4610,N_2867,N_3291);
or U4611 (N_4611,N_2638,N_2288);
nand U4612 (N_4612,N_3179,N_2581);
and U4613 (N_4613,N_3958,N_2617);
xor U4614 (N_4614,N_2374,N_2155);
or U4615 (N_4615,N_3194,N_2646);
or U4616 (N_4616,N_2308,N_3023);
nand U4617 (N_4617,N_2900,N_3078);
nand U4618 (N_4618,N_2413,N_2247);
and U4619 (N_4619,N_3034,N_3639);
and U4620 (N_4620,N_3008,N_3661);
and U4621 (N_4621,N_2815,N_2289);
xor U4622 (N_4622,N_3664,N_2089);
and U4623 (N_4623,N_3993,N_3302);
and U4624 (N_4624,N_3063,N_2699);
nand U4625 (N_4625,N_2163,N_2461);
and U4626 (N_4626,N_2122,N_2537);
xor U4627 (N_4627,N_2431,N_2611);
and U4628 (N_4628,N_2175,N_3567);
nor U4629 (N_4629,N_2408,N_2787);
or U4630 (N_4630,N_2445,N_3080);
nor U4631 (N_4631,N_3140,N_3225);
and U4632 (N_4632,N_2891,N_2410);
and U4633 (N_4633,N_3190,N_3905);
or U4634 (N_4634,N_2545,N_2870);
nor U4635 (N_4635,N_3030,N_3831);
nand U4636 (N_4636,N_2235,N_2691);
nand U4637 (N_4637,N_2765,N_2968);
or U4638 (N_4638,N_3866,N_3954);
nand U4639 (N_4639,N_2309,N_3659);
xor U4640 (N_4640,N_3138,N_2771);
nor U4641 (N_4641,N_3754,N_2587);
nand U4642 (N_4642,N_3894,N_3006);
nor U4643 (N_4643,N_2363,N_2042);
or U4644 (N_4644,N_2819,N_2811);
and U4645 (N_4645,N_2953,N_2965);
and U4646 (N_4646,N_2437,N_3157);
nand U4647 (N_4647,N_3547,N_3679);
nand U4648 (N_4648,N_2747,N_2606);
and U4649 (N_4649,N_3002,N_2393);
nand U4650 (N_4650,N_3493,N_2444);
nand U4651 (N_4651,N_2438,N_2600);
nand U4652 (N_4652,N_3041,N_2113);
and U4653 (N_4653,N_3730,N_2923);
xor U4654 (N_4654,N_2342,N_2286);
and U4655 (N_4655,N_2760,N_3931);
nand U4656 (N_4656,N_3733,N_3497);
or U4657 (N_4657,N_2848,N_3833);
nand U4658 (N_4658,N_2786,N_3256);
and U4659 (N_4659,N_3622,N_3450);
and U4660 (N_4660,N_2931,N_2504);
nor U4661 (N_4661,N_3513,N_3883);
nand U4662 (N_4662,N_3468,N_2774);
nand U4663 (N_4663,N_3629,N_2890);
nor U4664 (N_4664,N_2481,N_2799);
or U4665 (N_4665,N_2736,N_3371);
or U4666 (N_4666,N_3305,N_3899);
nand U4667 (N_4667,N_3591,N_3106);
or U4668 (N_4668,N_3079,N_2072);
or U4669 (N_4669,N_3414,N_2425);
and U4670 (N_4670,N_3528,N_2380);
nand U4671 (N_4671,N_2115,N_3329);
nor U4672 (N_4672,N_2543,N_3877);
or U4673 (N_4673,N_3986,N_2526);
nand U4674 (N_4674,N_3586,N_3136);
or U4675 (N_4675,N_2231,N_2443);
nor U4676 (N_4676,N_2406,N_2265);
and U4677 (N_4677,N_2610,N_2915);
xor U4678 (N_4678,N_3512,N_2672);
nand U4679 (N_4679,N_2593,N_2439);
and U4680 (N_4680,N_2754,N_2925);
and U4681 (N_4681,N_3681,N_2687);
or U4682 (N_4682,N_3956,N_2935);
nor U4683 (N_4683,N_3947,N_2863);
nand U4684 (N_4684,N_2567,N_2355);
and U4685 (N_4685,N_2080,N_3825);
xnor U4686 (N_4686,N_2826,N_3764);
nor U4687 (N_4687,N_2474,N_3356);
or U4688 (N_4688,N_2874,N_2557);
xnor U4689 (N_4689,N_3819,N_2763);
and U4690 (N_4690,N_3239,N_2304);
nand U4691 (N_4691,N_2535,N_2204);
nor U4692 (N_4692,N_2096,N_2021);
or U4693 (N_4693,N_3077,N_2974);
and U4694 (N_4694,N_2473,N_3685);
xor U4695 (N_4695,N_2580,N_3595);
nor U4696 (N_4696,N_2484,N_2578);
nand U4697 (N_4697,N_2398,N_3934);
nand U4698 (N_4698,N_3531,N_2917);
nor U4699 (N_4699,N_2629,N_2701);
nor U4700 (N_4700,N_3743,N_3806);
or U4701 (N_4701,N_2202,N_2938);
xor U4702 (N_4702,N_3593,N_2630);
xor U4703 (N_4703,N_2281,N_3895);
nand U4704 (N_4704,N_2642,N_3929);
and U4705 (N_4705,N_3734,N_2328);
or U4706 (N_4706,N_2090,N_3137);
nand U4707 (N_4707,N_2123,N_2702);
nand U4708 (N_4708,N_3798,N_3452);
xor U4709 (N_4709,N_2667,N_2975);
nor U4710 (N_4710,N_3037,N_2082);
or U4711 (N_4711,N_3940,N_2324);
nor U4712 (N_4712,N_3430,N_3650);
nor U4713 (N_4713,N_2828,N_3032);
nand U4714 (N_4714,N_2084,N_2888);
or U4715 (N_4715,N_3658,N_3665);
and U4716 (N_4716,N_3692,N_3364);
and U4717 (N_4717,N_3985,N_3913);
and U4718 (N_4718,N_2516,N_2507);
or U4719 (N_4719,N_2402,N_2232);
nand U4720 (N_4720,N_2670,N_3865);
nand U4721 (N_4721,N_2661,N_2844);
nor U4722 (N_4722,N_3472,N_3131);
and U4723 (N_4723,N_3024,N_3327);
xnor U4724 (N_4724,N_3662,N_3130);
nand U4725 (N_4725,N_3120,N_3259);
nor U4726 (N_4726,N_2148,N_3965);
nor U4727 (N_4727,N_3828,N_3980);
nand U4728 (N_4728,N_2608,N_2616);
nor U4729 (N_4729,N_2853,N_3891);
nor U4730 (N_4730,N_3501,N_2171);
nor U4731 (N_4731,N_3406,N_2347);
nor U4732 (N_4732,N_2129,N_3459);
nand U4733 (N_4733,N_3625,N_3912);
nor U4734 (N_4734,N_3368,N_2117);
nor U4735 (N_4735,N_3755,N_3322);
and U4736 (N_4736,N_3746,N_2447);
nand U4737 (N_4737,N_2479,N_2947);
nand U4738 (N_4738,N_3778,N_3112);
and U4739 (N_4739,N_3751,N_3793);
xor U4740 (N_4740,N_3221,N_2498);
and U4741 (N_4741,N_3417,N_3480);
and U4742 (N_4742,N_3303,N_3554);
xnor U4743 (N_4743,N_2579,N_2742);
xor U4744 (N_4744,N_3937,N_2730);
nand U4745 (N_4745,N_2469,N_3725);
nand U4746 (N_4746,N_2258,N_3165);
nor U4747 (N_4747,N_3354,N_2726);
nor U4748 (N_4748,N_2211,N_3907);
or U4749 (N_4749,N_3338,N_2519);
or U4750 (N_4750,N_2350,N_2405);
and U4751 (N_4751,N_2273,N_3380);
and U4752 (N_4752,N_2276,N_3854);
and U4753 (N_4753,N_2472,N_3578);
nor U4754 (N_4754,N_2840,N_2575);
xnor U4755 (N_4755,N_3615,N_3557);
and U4756 (N_4756,N_3750,N_3431);
nand U4757 (N_4757,N_3031,N_3208);
nand U4758 (N_4758,N_3770,N_3297);
nor U4759 (N_4759,N_3884,N_2706);
nand U4760 (N_4760,N_2977,N_2157);
or U4761 (N_4761,N_3802,N_3192);
nor U4762 (N_4762,N_3366,N_2994);
or U4763 (N_4763,N_2704,N_2664);
or U4764 (N_4764,N_3887,N_3525);
and U4765 (N_4765,N_2964,N_3552);
or U4766 (N_4766,N_2920,N_3508);
nor U4767 (N_4767,N_2782,N_2813);
or U4768 (N_4768,N_3781,N_3367);
nand U4769 (N_4769,N_2360,N_3146);
or U4770 (N_4770,N_2020,N_3849);
xnor U4771 (N_4771,N_2245,N_3744);
and U4772 (N_4772,N_3830,N_3053);
nor U4773 (N_4773,N_2238,N_2146);
xnor U4774 (N_4774,N_3133,N_3742);
xnor U4775 (N_4775,N_3151,N_3048);
nand U4776 (N_4776,N_3541,N_3473);
nor U4777 (N_4777,N_3278,N_3000);
and U4778 (N_4778,N_3783,N_2282);
nor U4779 (N_4779,N_3267,N_3577);
and U4780 (N_4780,N_2061,N_2223);
or U4781 (N_4781,N_2592,N_2002);
nand U4782 (N_4782,N_3059,N_3240);
nand U4783 (N_4783,N_3142,N_3555);
nor U4784 (N_4784,N_3935,N_3454);
nand U4785 (N_4785,N_3974,N_3046);
and U4786 (N_4786,N_3223,N_3295);
or U4787 (N_4787,N_3739,N_2371);
nor U4788 (N_4788,N_2412,N_2365);
nor U4789 (N_4789,N_2280,N_2435);
or U4790 (N_4790,N_2420,N_3738);
nor U4791 (N_4791,N_3007,N_2109);
or U4792 (N_4792,N_3084,N_2332);
and U4793 (N_4793,N_3377,N_3632);
or U4794 (N_4794,N_3144,N_3491);
and U4795 (N_4795,N_3769,N_2237);
nand U4796 (N_4796,N_2124,N_2166);
nand U4797 (N_4797,N_2009,N_3499);
and U4798 (N_4798,N_3321,N_3325);
nor U4799 (N_4799,N_2119,N_3924);
or U4800 (N_4800,N_2655,N_2803);
and U4801 (N_4801,N_2723,N_2690);
xnor U4802 (N_4802,N_2322,N_3102);
or U4803 (N_4803,N_2688,N_2216);
nor U4804 (N_4804,N_2305,N_2591);
and U4805 (N_4805,N_2207,N_3952);
nor U4806 (N_4806,N_3177,N_2601);
and U4807 (N_4807,N_2333,N_2210);
and U4808 (N_4808,N_3242,N_2029);
nand U4809 (N_4809,N_2035,N_3418);
or U4810 (N_4810,N_2353,N_3088);
nor U4811 (N_4811,N_2796,N_3588);
and U4812 (N_4812,N_2773,N_3779);
xnor U4813 (N_4813,N_2256,N_2407);
and U4814 (N_4814,N_3942,N_3786);
or U4815 (N_4815,N_3978,N_2441);
nand U4816 (N_4816,N_2881,N_3152);
xor U4817 (N_4817,N_3020,N_3611);
nor U4818 (N_4818,N_3716,N_3263);
and U4819 (N_4819,N_2749,N_2087);
nand U4820 (N_4820,N_3719,N_2887);
nand U4821 (N_4821,N_3994,N_3585);
and U4822 (N_4822,N_2121,N_3216);
nor U4823 (N_4823,N_3163,N_3229);
nor U4824 (N_4824,N_3191,N_3932);
nor U4825 (N_4825,N_3068,N_3432);
nor U4826 (N_4826,N_2855,N_3072);
or U4827 (N_4827,N_3407,N_3709);
or U4828 (N_4828,N_2879,N_2085);
and U4829 (N_4829,N_2159,N_2354);
xnor U4830 (N_4830,N_3674,N_3534);
nor U4831 (N_4831,N_3564,N_2602);
and U4832 (N_4832,N_2025,N_3049);
and U4833 (N_4833,N_2576,N_2415);
nor U4834 (N_4834,N_2816,N_2253);
and U4835 (N_4835,N_2299,N_3029);
and U4836 (N_4836,N_2766,N_3691);
or U4837 (N_4837,N_2525,N_2027);
nor U4838 (N_4838,N_3988,N_3644);
or U4839 (N_4839,N_2128,N_3276);
and U4840 (N_4840,N_3617,N_2094);
or U4841 (N_4841,N_2989,N_3453);
or U4842 (N_4842,N_2715,N_3970);
and U4843 (N_4843,N_2260,N_3684);
nor U4844 (N_4844,N_3300,N_3928);
xnor U4845 (N_4845,N_3253,N_2653);
or U4846 (N_4846,N_2685,N_2478);
or U4847 (N_4847,N_2048,N_3339);
nor U4848 (N_4848,N_2378,N_2068);
or U4849 (N_4849,N_3815,N_3864);
nand U4850 (N_4850,N_3495,N_3199);
nand U4851 (N_4851,N_3104,N_3979);
xnor U4852 (N_4852,N_2221,N_3269);
nand U4853 (N_4853,N_2669,N_3462);
nor U4854 (N_4854,N_3521,N_2480);
and U4855 (N_4855,N_3867,N_3139);
nor U4856 (N_4856,N_2275,N_3881);
or U4857 (N_4857,N_3310,N_3767);
nand U4858 (N_4858,N_3728,N_3941);
and U4859 (N_4859,N_2693,N_3538);
and U4860 (N_4860,N_2645,N_3540);
xnor U4861 (N_4861,N_2127,N_2792);
or U4862 (N_4862,N_3092,N_3915);
or U4863 (N_4863,N_2066,N_3159);
and U4864 (N_4864,N_3185,N_3282);
nand U4865 (N_4865,N_2218,N_2411);
and U4866 (N_4866,N_3141,N_3789);
nand U4867 (N_4867,N_3252,N_2838);
and U4868 (N_4868,N_3279,N_2462);
and U4869 (N_4869,N_2030,N_2641);
or U4870 (N_4870,N_3714,N_2534);
or U4871 (N_4871,N_2783,N_3910);
nand U4872 (N_4872,N_3817,N_3651);
nand U4873 (N_4873,N_2011,N_2936);
nor U4874 (N_4874,N_3792,N_3178);
nand U4875 (N_4875,N_2329,N_3584);
nand U4876 (N_4876,N_3700,N_2731);
xnor U4877 (N_4877,N_2359,N_2401);
and U4878 (N_4878,N_2644,N_2180);
or U4879 (N_4879,N_2903,N_3944);
nand U4880 (N_4880,N_3287,N_2001);
nor U4881 (N_4881,N_2729,N_2161);
xor U4882 (N_4882,N_3076,N_3925);
nand U4883 (N_4883,N_2597,N_2748);
and U4884 (N_4884,N_2517,N_2156);
or U4885 (N_4885,N_3161,N_2051);
nor U4886 (N_4886,N_2841,N_3457);
or U4887 (N_4887,N_2809,N_3156);
nand U4888 (N_4888,N_3766,N_3434);
xnor U4889 (N_4889,N_2497,N_2465);
or U4890 (N_4890,N_3481,N_3991);
nand U4891 (N_4891,N_3187,N_2450);
or U4892 (N_4892,N_2414,N_2527);
and U4893 (N_4893,N_3599,N_3948);
nor U4894 (N_4894,N_3173,N_2710);
nor U4895 (N_4895,N_2725,N_2356);
nand U4896 (N_4896,N_3124,N_2091);
and U4897 (N_4897,N_3258,N_3515);
and U4898 (N_4898,N_2712,N_3228);
or U4899 (N_4899,N_3614,N_3678);
nor U4900 (N_4900,N_3505,N_3655);
xor U4901 (N_4901,N_2069,N_3050);
nor U4902 (N_4902,N_2548,N_2499);
nor U4903 (N_4903,N_2287,N_2326);
nand U4904 (N_4904,N_3062,N_3596);
nor U4905 (N_4905,N_3708,N_3083);
nand U4906 (N_4906,N_2648,N_3745);
nor U4907 (N_4907,N_3805,N_3756);
and U4908 (N_4908,N_2769,N_2631);
nor U4909 (N_4909,N_2318,N_2106);
nor U4910 (N_4910,N_2116,N_2489);
or U4911 (N_4911,N_3268,N_2141);
nor U4912 (N_4912,N_3638,N_3471);
and U4913 (N_4913,N_2382,N_2847);
xnor U4914 (N_4914,N_3633,N_2821);
or U4915 (N_4915,N_2711,N_2341);
nor U4916 (N_4916,N_3469,N_2703);
xnor U4917 (N_4917,N_2105,N_3885);
or U4918 (N_4918,N_3382,N_3167);
nor U4919 (N_4919,N_3984,N_2429);
and U4920 (N_4920,N_3094,N_3906);
and U4921 (N_4921,N_2246,N_3234);
nand U4922 (N_4922,N_2228,N_3224);
and U4923 (N_4923,N_2770,N_3215);
nor U4924 (N_4924,N_2902,N_2737);
and U4925 (N_4925,N_3155,N_3847);
nand U4926 (N_4926,N_2271,N_2320);
xor U4927 (N_4927,N_2014,N_3626);
nand U4928 (N_4928,N_3775,N_2052);
xor U4929 (N_4929,N_3344,N_3476);
xnor U4930 (N_4930,N_2361,N_2370);
nand U4931 (N_4931,N_3879,N_2386);
nor U4932 (N_4932,N_2585,N_2562);
nor U4933 (N_4933,N_2409,N_2744);
and U4934 (N_4934,N_2603,N_3601);
and U4935 (N_4935,N_3990,N_3395);
or U4936 (N_4936,N_3657,N_2306);
nand U4937 (N_4937,N_2633,N_3319);
nor U4938 (N_4938,N_2861,N_2368);
nor U4939 (N_4939,N_3957,N_2032);
and U4940 (N_4940,N_3243,N_2569);
nor U4941 (N_4941,N_2395,N_2650);
nor U4942 (N_4942,N_2665,N_2721);
or U4943 (N_4943,N_3346,N_3245);
and U4944 (N_4944,N_3874,N_3365);
nand U4945 (N_4945,N_2772,N_3549);
or U4946 (N_4946,N_2565,N_2767);
nor U4947 (N_4947,N_3580,N_2233);
or U4948 (N_4948,N_3909,N_3923);
nor U4949 (N_4949,N_3035,N_2859);
or U4950 (N_4950,N_2751,N_3721);
nand U4951 (N_4951,N_3972,N_2618);
and U4952 (N_4952,N_3115,N_2044);
or U4953 (N_4953,N_3340,N_3464);
nor U4954 (N_4954,N_2205,N_3576);
nand U4955 (N_4955,N_3373,N_2946);
nor U4956 (N_4956,N_2432,N_3628);
xor U4957 (N_4957,N_3649,N_3605);
or U4958 (N_4958,N_2312,N_3336);
nor U4959 (N_4959,N_3370,N_2466);
nand U4960 (N_4960,N_3487,N_2251);
or U4961 (N_4961,N_2229,N_2208);
xnor U4962 (N_4962,N_3251,N_2019);
or U4963 (N_4963,N_3696,N_2960);
xnor U4964 (N_4964,N_3387,N_3107);
or U4965 (N_4965,N_2733,N_3846);
nand U4966 (N_4966,N_3949,N_2997);
or U4967 (N_4967,N_3575,N_2658);
or U4968 (N_4968,N_2992,N_3206);
and U4969 (N_4969,N_3715,N_3042);
xor U4970 (N_4970,N_2622,N_2530);
and U4971 (N_4971,N_2291,N_3723);
nand U4972 (N_4972,N_3522,N_3968);
or U4973 (N_4973,N_2643,N_3385);
or U4974 (N_4974,N_3574,N_3488);
or U4975 (N_4975,N_2160,N_2551);
and U4976 (N_4976,N_3311,N_2999);
and U4977 (N_4977,N_2905,N_3822);
nor U4978 (N_4978,N_2183,N_2788);
or U4979 (N_4979,N_3391,N_2323);
and U4980 (N_4980,N_3597,N_3189);
and U4981 (N_4981,N_3735,N_2501);
nor U4982 (N_4982,N_3127,N_3720);
and U4983 (N_4983,N_3043,N_2423);
or U4984 (N_4984,N_2150,N_2073);
xor U4985 (N_4985,N_2806,N_2804);
nand U4986 (N_4986,N_2384,N_2434);
or U4987 (N_4987,N_3011,N_3917);
or U4988 (N_4988,N_3272,N_2889);
nor U4989 (N_4989,N_2442,N_3396);
xor U4990 (N_4990,N_3962,N_3429);
and U4991 (N_4991,N_3838,N_2834);
or U4992 (N_4992,N_3451,N_3592);
nor U4993 (N_4993,N_3047,N_2198);
nand U4994 (N_4994,N_3898,N_3052);
and U4995 (N_4995,N_3353,N_3621);
nor U4996 (N_4996,N_3527,N_2007);
nand U4997 (N_4997,N_3762,N_3348);
and U4998 (N_4998,N_3005,N_3478);
or U4999 (N_4999,N_2632,N_2152);
nor U5000 (N_5000,N_2184,N_2168);
nor U5001 (N_5001,N_3521,N_3467);
and U5002 (N_5002,N_2446,N_3420);
or U5003 (N_5003,N_2429,N_3208);
and U5004 (N_5004,N_3275,N_2040);
nor U5005 (N_5005,N_3876,N_3166);
nand U5006 (N_5006,N_2416,N_2892);
nor U5007 (N_5007,N_2566,N_2010);
nor U5008 (N_5008,N_2380,N_3003);
nor U5009 (N_5009,N_3529,N_3434);
nor U5010 (N_5010,N_2211,N_3922);
or U5011 (N_5011,N_3913,N_3888);
and U5012 (N_5012,N_3126,N_2027);
and U5013 (N_5013,N_2551,N_2081);
and U5014 (N_5014,N_2843,N_2243);
nor U5015 (N_5015,N_2590,N_2489);
or U5016 (N_5016,N_2217,N_3146);
xnor U5017 (N_5017,N_3325,N_2418);
and U5018 (N_5018,N_3655,N_3345);
nand U5019 (N_5019,N_2683,N_2983);
nand U5020 (N_5020,N_3135,N_3164);
and U5021 (N_5021,N_3317,N_2909);
nor U5022 (N_5022,N_2189,N_3424);
xnor U5023 (N_5023,N_3557,N_3290);
nor U5024 (N_5024,N_3439,N_3925);
nand U5025 (N_5025,N_2572,N_2296);
and U5026 (N_5026,N_2640,N_2410);
and U5027 (N_5027,N_2291,N_2137);
nor U5028 (N_5028,N_2289,N_2383);
nor U5029 (N_5029,N_2881,N_3538);
nor U5030 (N_5030,N_3820,N_3501);
or U5031 (N_5031,N_2029,N_3707);
xnor U5032 (N_5032,N_3125,N_2281);
nor U5033 (N_5033,N_3524,N_2863);
or U5034 (N_5034,N_3917,N_2512);
xnor U5035 (N_5035,N_2930,N_3355);
nand U5036 (N_5036,N_2738,N_3562);
nand U5037 (N_5037,N_3584,N_3158);
and U5038 (N_5038,N_3943,N_2854);
and U5039 (N_5039,N_2950,N_3879);
nor U5040 (N_5040,N_3014,N_3751);
and U5041 (N_5041,N_2242,N_3612);
and U5042 (N_5042,N_2511,N_3542);
nand U5043 (N_5043,N_3299,N_3813);
nand U5044 (N_5044,N_2812,N_3008);
nor U5045 (N_5045,N_2739,N_2111);
or U5046 (N_5046,N_2476,N_3475);
and U5047 (N_5047,N_2855,N_2231);
nor U5048 (N_5048,N_2672,N_2634);
xor U5049 (N_5049,N_2944,N_2049);
xor U5050 (N_5050,N_3224,N_3469);
nand U5051 (N_5051,N_3918,N_2726);
nor U5052 (N_5052,N_2135,N_3495);
and U5053 (N_5053,N_3822,N_3406);
or U5054 (N_5054,N_2816,N_3300);
and U5055 (N_5055,N_2000,N_2304);
and U5056 (N_5056,N_3908,N_2313);
nor U5057 (N_5057,N_3266,N_2234);
and U5058 (N_5058,N_3432,N_3121);
and U5059 (N_5059,N_2113,N_3382);
nand U5060 (N_5060,N_3584,N_3765);
nor U5061 (N_5061,N_3206,N_2275);
or U5062 (N_5062,N_3553,N_3958);
or U5063 (N_5063,N_3104,N_2568);
nand U5064 (N_5064,N_3235,N_3244);
xor U5065 (N_5065,N_3857,N_3147);
nand U5066 (N_5066,N_3390,N_2713);
and U5067 (N_5067,N_2690,N_3046);
xor U5068 (N_5068,N_2042,N_3420);
nand U5069 (N_5069,N_2428,N_3599);
nor U5070 (N_5070,N_2284,N_2637);
nor U5071 (N_5071,N_2002,N_3012);
xor U5072 (N_5072,N_3299,N_2596);
nand U5073 (N_5073,N_2413,N_2507);
xnor U5074 (N_5074,N_2352,N_3281);
and U5075 (N_5075,N_3912,N_3895);
or U5076 (N_5076,N_2835,N_2200);
or U5077 (N_5077,N_2231,N_3105);
nand U5078 (N_5078,N_2449,N_2462);
nor U5079 (N_5079,N_2279,N_2349);
and U5080 (N_5080,N_3166,N_3197);
nor U5081 (N_5081,N_3032,N_2716);
xnor U5082 (N_5082,N_3690,N_3113);
xor U5083 (N_5083,N_2177,N_2195);
and U5084 (N_5084,N_3365,N_3410);
nor U5085 (N_5085,N_3443,N_2762);
nand U5086 (N_5086,N_2247,N_3264);
nand U5087 (N_5087,N_3756,N_3679);
or U5088 (N_5088,N_3999,N_2472);
nand U5089 (N_5089,N_3417,N_3804);
nor U5090 (N_5090,N_3496,N_2862);
or U5091 (N_5091,N_2661,N_2385);
nand U5092 (N_5092,N_3726,N_3327);
nor U5093 (N_5093,N_2222,N_2257);
and U5094 (N_5094,N_3068,N_3313);
nand U5095 (N_5095,N_2587,N_3318);
or U5096 (N_5096,N_3325,N_3754);
or U5097 (N_5097,N_3276,N_3325);
or U5098 (N_5098,N_3536,N_2140);
or U5099 (N_5099,N_3191,N_2487);
nor U5100 (N_5100,N_2192,N_2850);
nand U5101 (N_5101,N_3755,N_2880);
and U5102 (N_5102,N_3114,N_2819);
nor U5103 (N_5103,N_2156,N_2041);
and U5104 (N_5104,N_2103,N_2737);
xor U5105 (N_5105,N_2402,N_3587);
or U5106 (N_5106,N_2277,N_3042);
xor U5107 (N_5107,N_3951,N_2969);
and U5108 (N_5108,N_2515,N_3285);
and U5109 (N_5109,N_3270,N_3152);
or U5110 (N_5110,N_3577,N_3484);
nor U5111 (N_5111,N_2238,N_3562);
nor U5112 (N_5112,N_2772,N_3414);
and U5113 (N_5113,N_2489,N_2843);
nand U5114 (N_5114,N_2936,N_2882);
or U5115 (N_5115,N_3783,N_3275);
nor U5116 (N_5116,N_2107,N_2103);
and U5117 (N_5117,N_3433,N_2262);
xor U5118 (N_5118,N_2926,N_3005);
xnor U5119 (N_5119,N_3185,N_3047);
xor U5120 (N_5120,N_2864,N_2096);
or U5121 (N_5121,N_3158,N_3731);
and U5122 (N_5122,N_3428,N_2124);
or U5123 (N_5123,N_2622,N_3839);
nand U5124 (N_5124,N_2895,N_3067);
and U5125 (N_5125,N_2226,N_2140);
and U5126 (N_5126,N_2024,N_2430);
nand U5127 (N_5127,N_3134,N_2361);
nor U5128 (N_5128,N_2544,N_3113);
nor U5129 (N_5129,N_3578,N_3617);
and U5130 (N_5130,N_3707,N_3258);
or U5131 (N_5131,N_2639,N_3200);
and U5132 (N_5132,N_3034,N_2432);
xor U5133 (N_5133,N_2737,N_2118);
nor U5134 (N_5134,N_3033,N_3938);
nand U5135 (N_5135,N_3976,N_3196);
or U5136 (N_5136,N_3253,N_3210);
nor U5137 (N_5137,N_2491,N_2465);
or U5138 (N_5138,N_3265,N_2567);
nor U5139 (N_5139,N_3053,N_3153);
or U5140 (N_5140,N_2847,N_3362);
nand U5141 (N_5141,N_2557,N_3770);
or U5142 (N_5142,N_3389,N_2635);
and U5143 (N_5143,N_2483,N_2570);
or U5144 (N_5144,N_3638,N_3804);
nor U5145 (N_5145,N_3871,N_2840);
nor U5146 (N_5146,N_2193,N_3887);
nor U5147 (N_5147,N_3941,N_2769);
or U5148 (N_5148,N_3630,N_2099);
nor U5149 (N_5149,N_2270,N_3582);
and U5150 (N_5150,N_3309,N_2052);
or U5151 (N_5151,N_2094,N_3029);
nor U5152 (N_5152,N_2678,N_3613);
nand U5153 (N_5153,N_2874,N_2972);
nor U5154 (N_5154,N_3227,N_3166);
or U5155 (N_5155,N_2024,N_2730);
or U5156 (N_5156,N_3436,N_2864);
nor U5157 (N_5157,N_3577,N_2876);
and U5158 (N_5158,N_3794,N_3806);
nor U5159 (N_5159,N_2517,N_2908);
or U5160 (N_5160,N_2489,N_3554);
and U5161 (N_5161,N_3583,N_2490);
nor U5162 (N_5162,N_2450,N_2639);
nand U5163 (N_5163,N_2062,N_3079);
or U5164 (N_5164,N_3883,N_2626);
nor U5165 (N_5165,N_2079,N_2414);
nand U5166 (N_5166,N_3024,N_2807);
nor U5167 (N_5167,N_2887,N_3968);
and U5168 (N_5168,N_3873,N_3542);
and U5169 (N_5169,N_2928,N_2400);
nor U5170 (N_5170,N_2178,N_3128);
nand U5171 (N_5171,N_3725,N_3836);
and U5172 (N_5172,N_2235,N_3671);
or U5173 (N_5173,N_2214,N_2898);
nand U5174 (N_5174,N_3988,N_3566);
and U5175 (N_5175,N_3286,N_2468);
and U5176 (N_5176,N_2228,N_2403);
nand U5177 (N_5177,N_2405,N_2504);
nor U5178 (N_5178,N_2032,N_2924);
xnor U5179 (N_5179,N_2920,N_3349);
nor U5180 (N_5180,N_3255,N_3600);
and U5181 (N_5181,N_2545,N_2403);
or U5182 (N_5182,N_2270,N_2136);
nand U5183 (N_5183,N_2173,N_3632);
and U5184 (N_5184,N_3723,N_3318);
nand U5185 (N_5185,N_2570,N_2105);
or U5186 (N_5186,N_3937,N_3868);
nor U5187 (N_5187,N_3721,N_3489);
nor U5188 (N_5188,N_2230,N_3672);
or U5189 (N_5189,N_3549,N_2360);
or U5190 (N_5190,N_3308,N_2034);
and U5191 (N_5191,N_3124,N_3471);
nand U5192 (N_5192,N_3857,N_2375);
or U5193 (N_5193,N_3180,N_3480);
and U5194 (N_5194,N_2269,N_3118);
nand U5195 (N_5195,N_3382,N_2805);
nor U5196 (N_5196,N_3071,N_3088);
nor U5197 (N_5197,N_3685,N_2542);
nand U5198 (N_5198,N_3246,N_3404);
nor U5199 (N_5199,N_3162,N_2235);
nor U5200 (N_5200,N_2771,N_3162);
nor U5201 (N_5201,N_2464,N_2640);
or U5202 (N_5202,N_2087,N_3259);
and U5203 (N_5203,N_2525,N_2214);
and U5204 (N_5204,N_3902,N_3918);
nor U5205 (N_5205,N_3158,N_2696);
nand U5206 (N_5206,N_3030,N_3213);
or U5207 (N_5207,N_2279,N_2568);
and U5208 (N_5208,N_2881,N_2874);
and U5209 (N_5209,N_3179,N_3587);
nand U5210 (N_5210,N_2003,N_2322);
and U5211 (N_5211,N_3149,N_2111);
nand U5212 (N_5212,N_2560,N_3655);
nand U5213 (N_5213,N_2376,N_2825);
nor U5214 (N_5214,N_2557,N_2060);
nor U5215 (N_5215,N_3097,N_3943);
and U5216 (N_5216,N_3121,N_2615);
and U5217 (N_5217,N_3782,N_3520);
nand U5218 (N_5218,N_3552,N_2504);
and U5219 (N_5219,N_2893,N_3755);
nand U5220 (N_5220,N_2391,N_3034);
or U5221 (N_5221,N_2956,N_2208);
nor U5222 (N_5222,N_2536,N_3789);
or U5223 (N_5223,N_3556,N_3252);
and U5224 (N_5224,N_3364,N_3008);
and U5225 (N_5225,N_2635,N_3248);
or U5226 (N_5226,N_2719,N_2668);
and U5227 (N_5227,N_3489,N_2048);
or U5228 (N_5228,N_3576,N_3924);
xor U5229 (N_5229,N_2652,N_2750);
nand U5230 (N_5230,N_3983,N_3985);
and U5231 (N_5231,N_2728,N_3197);
nand U5232 (N_5232,N_3000,N_3910);
and U5233 (N_5233,N_3273,N_3426);
nand U5234 (N_5234,N_3023,N_3241);
nor U5235 (N_5235,N_2038,N_3836);
nand U5236 (N_5236,N_3431,N_2043);
xnor U5237 (N_5237,N_2441,N_2949);
xnor U5238 (N_5238,N_3518,N_2320);
and U5239 (N_5239,N_2379,N_3064);
xor U5240 (N_5240,N_3056,N_2263);
nand U5241 (N_5241,N_3154,N_2884);
nor U5242 (N_5242,N_3779,N_2103);
nand U5243 (N_5243,N_3373,N_3897);
xor U5244 (N_5244,N_3725,N_3400);
or U5245 (N_5245,N_2641,N_2226);
nand U5246 (N_5246,N_3678,N_2265);
or U5247 (N_5247,N_3299,N_2873);
nand U5248 (N_5248,N_3365,N_2273);
or U5249 (N_5249,N_2556,N_2114);
and U5250 (N_5250,N_2069,N_3235);
and U5251 (N_5251,N_3409,N_3957);
nor U5252 (N_5252,N_2610,N_3038);
and U5253 (N_5253,N_2956,N_2127);
nor U5254 (N_5254,N_2197,N_3663);
nand U5255 (N_5255,N_3994,N_2656);
nor U5256 (N_5256,N_2091,N_3349);
nand U5257 (N_5257,N_3246,N_2493);
nor U5258 (N_5258,N_3590,N_2589);
nand U5259 (N_5259,N_3474,N_2071);
and U5260 (N_5260,N_2204,N_3638);
or U5261 (N_5261,N_3735,N_2100);
or U5262 (N_5262,N_2362,N_2504);
xnor U5263 (N_5263,N_3199,N_2868);
nand U5264 (N_5264,N_2580,N_2485);
or U5265 (N_5265,N_2302,N_2919);
nor U5266 (N_5266,N_2589,N_2723);
and U5267 (N_5267,N_2230,N_3535);
nand U5268 (N_5268,N_3485,N_3594);
nor U5269 (N_5269,N_3484,N_3346);
and U5270 (N_5270,N_3460,N_3070);
or U5271 (N_5271,N_3666,N_3831);
nand U5272 (N_5272,N_2471,N_3627);
and U5273 (N_5273,N_3431,N_2228);
or U5274 (N_5274,N_2467,N_2165);
nor U5275 (N_5275,N_2843,N_3605);
nor U5276 (N_5276,N_2935,N_3773);
and U5277 (N_5277,N_3154,N_2871);
nand U5278 (N_5278,N_2263,N_2012);
or U5279 (N_5279,N_2244,N_2342);
nor U5280 (N_5280,N_2587,N_3994);
nor U5281 (N_5281,N_3673,N_2739);
and U5282 (N_5282,N_3563,N_2087);
xnor U5283 (N_5283,N_2955,N_2292);
nor U5284 (N_5284,N_2759,N_2503);
or U5285 (N_5285,N_3255,N_2496);
nor U5286 (N_5286,N_2763,N_2766);
or U5287 (N_5287,N_3370,N_2857);
nor U5288 (N_5288,N_2205,N_2110);
or U5289 (N_5289,N_3354,N_2510);
nor U5290 (N_5290,N_3601,N_3896);
or U5291 (N_5291,N_2194,N_2370);
and U5292 (N_5292,N_3893,N_3774);
xnor U5293 (N_5293,N_3727,N_3951);
and U5294 (N_5294,N_3796,N_3809);
and U5295 (N_5295,N_3526,N_3451);
nor U5296 (N_5296,N_2165,N_3805);
and U5297 (N_5297,N_3590,N_2735);
xor U5298 (N_5298,N_2867,N_3475);
and U5299 (N_5299,N_3136,N_3653);
nor U5300 (N_5300,N_2025,N_3278);
xor U5301 (N_5301,N_3164,N_3702);
nand U5302 (N_5302,N_2397,N_2798);
or U5303 (N_5303,N_2019,N_3003);
xnor U5304 (N_5304,N_2879,N_2384);
and U5305 (N_5305,N_3079,N_2565);
nand U5306 (N_5306,N_2913,N_2121);
nor U5307 (N_5307,N_3107,N_3528);
nor U5308 (N_5308,N_2740,N_2844);
nor U5309 (N_5309,N_2843,N_2908);
nor U5310 (N_5310,N_2864,N_3733);
and U5311 (N_5311,N_2495,N_2710);
and U5312 (N_5312,N_2488,N_3817);
nor U5313 (N_5313,N_2497,N_3090);
nor U5314 (N_5314,N_3828,N_2571);
and U5315 (N_5315,N_3919,N_2922);
or U5316 (N_5316,N_3490,N_2454);
xnor U5317 (N_5317,N_3720,N_3809);
nand U5318 (N_5318,N_3052,N_2999);
nor U5319 (N_5319,N_2397,N_2859);
nand U5320 (N_5320,N_3104,N_3570);
nand U5321 (N_5321,N_3698,N_3375);
nand U5322 (N_5322,N_2327,N_2056);
nor U5323 (N_5323,N_2869,N_2416);
nand U5324 (N_5324,N_3600,N_3583);
or U5325 (N_5325,N_3684,N_2872);
nor U5326 (N_5326,N_3351,N_3778);
nand U5327 (N_5327,N_3899,N_3173);
or U5328 (N_5328,N_3652,N_3319);
nand U5329 (N_5329,N_2407,N_2564);
or U5330 (N_5330,N_3633,N_2091);
nor U5331 (N_5331,N_3246,N_3201);
nand U5332 (N_5332,N_2836,N_3415);
nand U5333 (N_5333,N_3619,N_2742);
nand U5334 (N_5334,N_2209,N_3865);
and U5335 (N_5335,N_2376,N_2947);
and U5336 (N_5336,N_3481,N_3578);
nor U5337 (N_5337,N_2811,N_2871);
nor U5338 (N_5338,N_3235,N_2782);
or U5339 (N_5339,N_2235,N_3033);
and U5340 (N_5340,N_2405,N_3001);
or U5341 (N_5341,N_3233,N_3499);
and U5342 (N_5342,N_3865,N_2114);
and U5343 (N_5343,N_3748,N_3941);
nand U5344 (N_5344,N_3416,N_3826);
xor U5345 (N_5345,N_3168,N_3687);
or U5346 (N_5346,N_2514,N_3014);
nand U5347 (N_5347,N_2165,N_2255);
nor U5348 (N_5348,N_3926,N_2269);
or U5349 (N_5349,N_3452,N_3485);
and U5350 (N_5350,N_2826,N_2751);
nor U5351 (N_5351,N_3940,N_3255);
or U5352 (N_5352,N_2999,N_3979);
or U5353 (N_5353,N_3585,N_3517);
nor U5354 (N_5354,N_3734,N_3619);
or U5355 (N_5355,N_2264,N_2697);
and U5356 (N_5356,N_3156,N_3826);
or U5357 (N_5357,N_2091,N_3528);
xnor U5358 (N_5358,N_2061,N_3082);
or U5359 (N_5359,N_2477,N_2390);
nor U5360 (N_5360,N_2040,N_3502);
nand U5361 (N_5361,N_3370,N_3183);
nor U5362 (N_5362,N_3268,N_3866);
or U5363 (N_5363,N_2307,N_3121);
nand U5364 (N_5364,N_3685,N_2852);
nand U5365 (N_5365,N_3899,N_2736);
or U5366 (N_5366,N_3753,N_3696);
or U5367 (N_5367,N_2614,N_3354);
nor U5368 (N_5368,N_2374,N_3374);
nor U5369 (N_5369,N_3661,N_2078);
or U5370 (N_5370,N_3664,N_3911);
and U5371 (N_5371,N_2375,N_2631);
nor U5372 (N_5372,N_3272,N_3123);
or U5373 (N_5373,N_2215,N_3004);
and U5374 (N_5374,N_3030,N_2047);
or U5375 (N_5375,N_2179,N_2344);
nand U5376 (N_5376,N_2135,N_3152);
nand U5377 (N_5377,N_2506,N_2355);
and U5378 (N_5378,N_2977,N_2161);
xnor U5379 (N_5379,N_3993,N_3389);
xor U5380 (N_5380,N_3173,N_3696);
or U5381 (N_5381,N_2524,N_2235);
or U5382 (N_5382,N_3739,N_3978);
or U5383 (N_5383,N_3365,N_3333);
nor U5384 (N_5384,N_3045,N_2657);
or U5385 (N_5385,N_2410,N_3303);
nand U5386 (N_5386,N_3597,N_2232);
nor U5387 (N_5387,N_3273,N_2138);
nand U5388 (N_5388,N_3319,N_2003);
nor U5389 (N_5389,N_2800,N_2883);
nor U5390 (N_5390,N_3366,N_3002);
nand U5391 (N_5391,N_3792,N_2515);
nand U5392 (N_5392,N_3900,N_3161);
nand U5393 (N_5393,N_3580,N_2068);
and U5394 (N_5394,N_2125,N_3556);
nand U5395 (N_5395,N_3429,N_2710);
nor U5396 (N_5396,N_2111,N_3560);
or U5397 (N_5397,N_3803,N_3925);
or U5398 (N_5398,N_3239,N_3702);
or U5399 (N_5399,N_3810,N_3113);
nor U5400 (N_5400,N_2951,N_3797);
or U5401 (N_5401,N_2680,N_2874);
and U5402 (N_5402,N_3267,N_3705);
nor U5403 (N_5403,N_3612,N_2220);
xor U5404 (N_5404,N_2304,N_2137);
nand U5405 (N_5405,N_2664,N_2897);
nor U5406 (N_5406,N_2570,N_2707);
nand U5407 (N_5407,N_3887,N_3808);
and U5408 (N_5408,N_3297,N_2681);
or U5409 (N_5409,N_2590,N_3479);
and U5410 (N_5410,N_3429,N_3550);
nand U5411 (N_5411,N_2993,N_2663);
nand U5412 (N_5412,N_3800,N_2960);
and U5413 (N_5413,N_2435,N_2715);
xor U5414 (N_5414,N_2350,N_2143);
nand U5415 (N_5415,N_2453,N_3527);
nand U5416 (N_5416,N_2289,N_3185);
xnor U5417 (N_5417,N_2185,N_2269);
nor U5418 (N_5418,N_3449,N_3188);
or U5419 (N_5419,N_2587,N_2149);
xnor U5420 (N_5420,N_2984,N_3877);
nor U5421 (N_5421,N_2894,N_2825);
nor U5422 (N_5422,N_2188,N_2764);
nor U5423 (N_5423,N_3338,N_2134);
nor U5424 (N_5424,N_2461,N_2902);
nor U5425 (N_5425,N_2827,N_2690);
nand U5426 (N_5426,N_2293,N_2478);
and U5427 (N_5427,N_2434,N_2120);
and U5428 (N_5428,N_3464,N_3400);
nor U5429 (N_5429,N_2340,N_3055);
and U5430 (N_5430,N_2348,N_3366);
nand U5431 (N_5431,N_2108,N_2390);
and U5432 (N_5432,N_3544,N_2794);
and U5433 (N_5433,N_3012,N_2983);
or U5434 (N_5434,N_3129,N_2505);
nand U5435 (N_5435,N_2840,N_2045);
and U5436 (N_5436,N_3347,N_3122);
or U5437 (N_5437,N_3777,N_3588);
nand U5438 (N_5438,N_2665,N_2894);
nor U5439 (N_5439,N_3450,N_3135);
and U5440 (N_5440,N_3795,N_3228);
or U5441 (N_5441,N_3378,N_2197);
or U5442 (N_5442,N_3998,N_3132);
and U5443 (N_5443,N_3997,N_3925);
nand U5444 (N_5444,N_2535,N_3800);
and U5445 (N_5445,N_2895,N_3523);
xor U5446 (N_5446,N_2086,N_2650);
nand U5447 (N_5447,N_2500,N_2290);
and U5448 (N_5448,N_3152,N_2723);
or U5449 (N_5449,N_2098,N_3593);
nand U5450 (N_5450,N_2083,N_2627);
xor U5451 (N_5451,N_3883,N_2448);
or U5452 (N_5452,N_2374,N_3810);
nor U5453 (N_5453,N_2443,N_3679);
and U5454 (N_5454,N_2699,N_2480);
nor U5455 (N_5455,N_2716,N_2354);
and U5456 (N_5456,N_2719,N_2044);
or U5457 (N_5457,N_2213,N_3727);
and U5458 (N_5458,N_3887,N_2059);
nor U5459 (N_5459,N_3528,N_3694);
and U5460 (N_5460,N_3600,N_3373);
nand U5461 (N_5461,N_3223,N_2608);
nand U5462 (N_5462,N_2599,N_3933);
nand U5463 (N_5463,N_3306,N_3379);
and U5464 (N_5464,N_2571,N_2079);
or U5465 (N_5465,N_2835,N_2109);
or U5466 (N_5466,N_2425,N_3950);
or U5467 (N_5467,N_3219,N_3937);
nor U5468 (N_5468,N_2817,N_2291);
or U5469 (N_5469,N_3485,N_2702);
xor U5470 (N_5470,N_3754,N_3840);
nand U5471 (N_5471,N_2485,N_3458);
xor U5472 (N_5472,N_2474,N_3121);
or U5473 (N_5473,N_3356,N_2217);
and U5474 (N_5474,N_2419,N_2478);
nor U5475 (N_5475,N_3594,N_3647);
or U5476 (N_5476,N_3495,N_3397);
or U5477 (N_5477,N_3181,N_2779);
or U5478 (N_5478,N_3975,N_2740);
or U5479 (N_5479,N_2869,N_3573);
or U5480 (N_5480,N_2474,N_3071);
nand U5481 (N_5481,N_2846,N_3858);
nand U5482 (N_5482,N_3329,N_3218);
or U5483 (N_5483,N_3069,N_2240);
or U5484 (N_5484,N_3106,N_3248);
nand U5485 (N_5485,N_3004,N_3195);
or U5486 (N_5486,N_2564,N_3876);
nor U5487 (N_5487,N_2131,N_2814);
and U5488 (N_5488,N_3679,N_3518);
and U5489 (N_5489,N_3779,N_3918);
nor U5490 (N_5490,N_2658,N_3839);
nor U5491 (N_5491,N_2846,N_2323);
nand U5492 (N_5492,N_2695,N_3838);
or U5493 (N_5493,N_2847,N_2679);
and U5494 (N_5494,N_3264,N_2591);
or U5495 (N_5495,N_2784,N_3116);
and U5496 (N_5496,N_3573,N_2747);
or U5497 (N_5497,N_3315,N_3356);
nor U5498 (N_5498,N_2997,N_3488);
or U5499 (N_5499,N_3342,N_3574);
nor U5500 (N_5500,N_2973,N_2136);
nand U5501 (N_5501,N_3555,N_3111);
nor U5502 (N_5502,N_3881,N_2812);
and U5503 (N_5503,N_2028,N_2367);
or U5504 (N_5504,N_2013,N_3815);
nor U5505 (N_5505,N_3158,N_3214);
nor U5506 (N_5506,N_2560,N_2624);
and U5507 (N_5507,N_2536,N_2425);
nand U5508 (N_5508,N_2197,N_2120);
nand U5509 (N_5509,N_2587,N_2576);
and U5510 (N_5510,N_2277,N_3273);
xnor U5511 (N_5511,N_2667,N_2231);
nor U5512 (N_5512,N_2127,N_3075);
and U5513 (N_5513,N_3810,N_2377);
or U5514 (N_5514,N_3662,N_3218);
nor U5515 (N_5515,N_3195,N_3238);
or U5516 (N_5516,N_3608,N_3773);
nor U5517 (N_5517,N_2076,N_2154);
xnor U5518 (N_5518,N_2364,N_3927);
nor U5519 (N_5519,N_3572,N_3869);
or U5520 (N_5520,N_3074,N_2685);
and U5521 (N_5521,N_3278,N_3188);
nor U5522 (N_5522,N_2934,N_2126);
nand U5523 (N_5523,N_2888,N_2316);
or U5524 (N_5524,N_2790,N_2479);
nor U5525 (N_5525,N_2327,N_3598);
nor U5526 (N_5526,N_2449,N_2771);
or U5527 (N_5527,N_2744,N_2480);
and U5528 (N_5528,N_2515,N_2378);
xnor U5529 (N_5529,N_3787,N_3302);
or U5530 (N_5530,N_2937,N_3120);
and U5531 (N_5531,N_2223,N_2945);
and U5532 (N_5532,N_3992,N_3404);
nor U5533 (N_5533,N_3537,N_3019);
nor U5534 (N_5534,N_2211,N_2149);
nand U5535 (N_5535,N_2328,N_2456);
nand U5536 (N_5536,N_2324,N_3063);
nor U5537 (N_5537,N_3856,N_3905);
or U5538 (N_5538,N_3002,N_2841);
and U5539 (N_5539,N_3213,N_2646);
or U5540 (N_5540,N_3222,N_2010);
nand U5541 (N_5541,N_3949,N_3979);
or U5542 (N_5542,N_2346,N_2458);
and U5543 (N_5543,N_3157,N_2516);
and U5544 (N_5544,N_2242,N_2728);
and U5545 (N_5545,N_2120,N_3246);
and U5546 (N_5546,N_2342,N_2443);
nor U5547 (N_5547,N_2035,N_3254);
nor U5548 (N_5548,N_3113,N_2698);
and U5549 (N_5549,N_3939,N_3283);
nor U5550 (N_5550,N_2473,N_3874);
nor U5551 (N_5551,N_3302,N_3738);
or U5552 (N_5552,N_2868,N_2695);
or U5553 (N_5553,N_2789,N_3741);
or U5554 (N_5554,N_2310,N_3023);
or U5555 (N_5555,N_2524,N_2231);
or U5556 (N_5556,N_3610,N_2609);
nand U5557 (N_5557,N_2185,N_3444);
nand U5558 (N_5558,N_2046,N_2019);
or U5559 (N_5559,N_2900,N_3823);
xor U5560 (N_5560,N_3101,N_2402);
xnor U5561 (N_5561,N_3884,N_3406);
or U5562 (N_5562,N_2396,N_2153);
xnor U5563 (N_5563,N_3755,N_3169);
nand U5564 (N_5564,N_3519,N_3212);
and U5565 (N_5565,N_3613,N_3943);
xnor U5566 (N_5566,N_3542,N_3749);
nor U5567 (N_5567,N_3602,N_3304);
nor U5568 (N_5568,N_2163,N_2409);
or U5569 (N_5569,N_2896,N_3815);
and U5570 (N_5570,N_3435,N_3268);
nor U5571 (N_5571,N_3420,N_3418);
and U5572 (N_5572,N_3512,N_3850);
or U5573 (N_5573,N_2941,N_3633);
xnor U5574 (N_5574,N_2094,N_3820);
and U5575 (N_5575,N_3067,N_2369);
and U5576 (N_5576,N_2612,N_2140);
nand U5577 (N_5577,N_3561,N_3138);
nor U5578 (N_5578,N_2139,N_3904);
nor U5579 (N_5579,N_2196,N_3486);
or U5580 (N_5580,N_3203,N_2803);
and U5581 (N_5581,N_3476,N_3065);
or U5582 (N_5582,N_3392,N_2628);
nand U5583 (N_5583,N_2296,N_3239);
nand U5584 (N_5584,N_3330,N_3200);
nor U5585 (N_5585,N_3368,N_3947);
nand U5586 (N_5586,N_2827,N_2398);
nor U5587 (N_5587,N_2052,N_2059);
and U5588 (N_5588,N_2623,N_3840);
or U5589 (N_5589,N_2307,N_3463);
xnor U5590 (N_5590,N_2515,N_2757);
and U5591 (N_5591,N_3515,N_2650);
nand U5592 (N_5592,N_3587,N_2273);
and U5593 (N_5593,N_3882,N_3306);
nand U5594 (N_5594,N_2940,N_3439);
nand U5595 (N_5595,N_2797,N_2839);
xor U5596 (N_5596,N_2964,N_3935);
and U5597 (N_5597,N_3468,N_2588);
and U5598 (N_5598,N_3729,N_2091);
nand U5599 (N_5599,N_3758,N_3401);
or U5600 (N_5600,N_3275,N_2386);
nand U5601 (N_5601,N_2178,N_2081);
and U5602 (N_5602,N_2655,N_2345);
nand U5603 (N_5603,N_2500,N_3161);
nand U5604 (N_5604,N_2611,N_2612);
nand U5605 (N_5605,N_2731,N_2947);
and U5606 (N_5606,N_2114,N_2382);
xor U5607 (N_5607,N_3826,N_3351);
or U5608 (N_5608,N_3363,N_3004);
and U5609 (N_5609,N_3456,N_3128);
or U5610 (N_5610,N_3568,N_3681);
and U5611 (N_5611,N_2699,N_3874);
and U5612 (N_5612,N_3042,N_2946);
and U5613 (N_5613,N_2008,N_3954);
nor U5614 (N_5614,N_3152,N_2789);
and U5615 (N_5615,N_3412,N_2493);
or U5616 (N_5616,N_3162,N_2770);
and U5617 (N_5617,N_3435,N_2483);
nand U5618 (N_5618,N_3354,N_2060);
and U5619 (N_5619,N_2238,N_3957);
and U5620 (N_5620,N_3947,N_2474);
or U5621 (N_5621,N_2463,N_2807);
nand U5622 (N_5622,N_2278,N_3674);
xnor U5623 (N_5623,N_2524,N_2534);
or U5624 (N_5624,N_2145,N_3630);
nand U5625 (N_5625,N_3112,N_2765);
or U5626 (N_5626,N_2863,N_3923);
or U5627 (N_5627,N_3516,N_3092);
nand U5628 (N_5628,N_3625,N_3555);
nand U5629 (N_5629,N_2645,N_3854);
xor U5630 (N_5630,N_2820,N_2434);
and U5631 (N_5631,N_2904,N_2901);
or U5632 (N_5632,N_2023,N_2811);
xnor U5633 (N_5633,N_2048,N_2171);
xor U5634 (N_5634,N_2428,N_3305);
nor U5635 (N_5635,N_3513,N_2202);
or U5636 (N_5636,N_2510,N_3770);
and U5637 (N_5637,N_2039,N_2811);
nor U5638 (N_5638,N_2098,N_3017);
nor U5639 (N_5639,N_3707,N_3786);
xor U5640 (N_5640,N_3363,N_2315);
and U5641 (N_5641,N_3959,N_3960);
nor U5642 (N_5642,N_3656,N_3840);
xor U5643 (N_5643,N_2423,N_2340);
or U5644 (N_5644,N_2852,N_3640);
nor U5645 (N_5645,N_2050,N_3520);
or U5646 (N_5646,N_2446,N_3553);
xor U5647 (N_5647,N_3235,N_2053);
nor U5648 (N_5648,N_2870,N_2015);
and U5649 (N_5649,N_2067,N_3616);
and U5650 (N_5650,N_2512,N_2307);
and U5651 (N_5651,N_2233,N_3729);
nor U5652 (N_5652,N_2397,N_3820);
or U5653 (N_5653,N_3780,N_2163);
nor U5654 (N_5654,N_2563,N_3208);
nor U5655 (N_5655,N_3528,N_2320);
and U5656 (N_5656,N_2513,N_3009);
xnor U5657 (N_5657,N_3640,N_3600);
xnor U5658 (N_5658,N_3628,N_2715);
nand U5659 (N_5659,N_3638,N_2912);
or U5660 (N_5660,N_2731,N_2323);
or U5661 (N_5661,N_3441,N_2507);
nor U5662 (N_5662,N_2626,N_2704);
nand U5663 (N_5663,N_3316,N_2309);
nor U5664 (N_5664,N_3505,N_3103);
xnor U5665 (N_5665,N_2021,N_2635);
and U5666 (N_5666,N_3588,N_3736);
nand U5667 (N_5667,N_2136,N_2690);
nor U5668 (N_5668,N_3945,N_3631);
nor U5669 (N_5669,N_3898,N_2697);
nor U5670 (N_5670,N_2957,N_2466);
xnor U5671 (N_5671,N_2051,N_2377);
and U5672 (N_5672,N_3530,N_3543);
and U5673 (N_5673,N_2304,N_2757);
nor U5674 (N_5674,N_2776,N_2123);
and U5675 (N_5675,N_2217,N_3895);
xor U5676 (N_5676,N_3567,N_2088);
nor U5677 (N_5677,N_3995,N_2519);
and U5678 (N_5678,N_2966,N_2907);
or U5679 (N_5679,N_2348,N_2840);
nor U5680 (N_5680,N_3757,N_2198);
and U5681 (N_5681,N_2407,N_3423);
or U5682 (N_5682,N_3256,N_2549);
nor U5683 (N_5683,N_2334,N_2479);
xnor U5684 (N_5684,N_3965,N_3126);
nand U5685 (N_5685,N_3632,N_3813);
and U5686 (N_5686,N_3489,N_3881);
nor U5687 (N_5687,N_3457,N_2512);
or U5688 (N_5688,N_3834,N_3087);
or U5689 (N_5689,N_2592,N_2123);
or U5690 (N_5690,N_3652,N_2403);
nor U5691 (N_5691,N_2707,N_2553);
and U5692 (N_5692,N_3867,N_2959);
xnor U5693 (N_5693,N_3562,N_3121);
or U5694 (N_5694,N_3070,N_3122);
or U5695 (N_5695,N_2703,N_2407);
and U5696 (N_5696,N_3560,N_2698);
or U5697 (N_5697,N_2279,N_3759);
xnor U5698 (N_5698,N_2545,N_2941);
nor U5699 (N_5699,N_3392,N_2396);
nor U5700 (N_5700,N_3624,N_2463);
xnor U5701 (N_5701,N_2919,N_2927);
nand U5702 (N_5702,N_3390,N_3252);
or U5703 (N_5703,N_2266,N_3730);
and U5704 (N_5704,N_2209,N_2464);
nor U5705 (N_5705,N_2977,N_3404);
nor U5706 (N_5706,N_3640,N_3756);
xnor U5707 (N_5707,N_3428,N_2754);
nand U5708 (N_5708,N_3866,N_3651);
xnor U5709 (N_5709,N_2236,N_3406);
nor U5710 (N_5710,N_3869,N_2294);
or U5711 (N_5711,N_2319,N_2183);
nand U5712 (N_5712,N_2946,N_2366);
nor U5713 (N_5713,N_2661,N_3449);
nor U5714 (N_5714,N_2421,N_2023);
or U5715 (N_5715,N_2882,N_3895);
and U5716 (N_5716,N_2721,N_3649);
and U5717 (N_5717,N_3884,N_3017);
or U5718 (N_5718,N_2180,N_2850);
and U5719 (N_5719,N_3845,N_2745);
nor U5720 (N_5720,N_3801,N_3009);
or U5721 (N_5721,N_2369,N_3935);
and U5722 (N_5722,N_2727,N_3905);
nor U5723 (N_5723,N_3242,N_3118);
and U5724 (N_5724,N_3362,N_2990);
or U5725 (N_5725,N_2624,N_2335);
nor U5726 (N_5726,N_2656,N_2246);
nor U5727 (N_5727,N_3694,N_2173);
nor U5728 (N_5728,N_3231,N_2777);
xnor U5729 (N_5729,N_3528,N_3867);
or U5730 (N_5730,N_2564,N_2716);
xnor U5731 (N_5731,N_2770,N_2036);
or U5732 (N_5732,N_2365,N_3373);
and U5733 (N_5733,N_3448,N_3262);
nand U5734 (N_5734,N_2972,N_2111);
nor U5735 (N_5735,N_2930,N_2493);
nand U5736 (N_5736,N_3099,N_3988);
nor U5737 (N_5737,N_2390,N_2100);
or U5738 (N_5738,N_3133,N_3013);
nand U5739 (N_5739,N_3997,N_2227);
nor U5740 (N_5740,N_3437,N_3873);
or U5741 (N_5741,N_2021,N_2546);
nor U5742 (N_5742,N_2455,N_3588);
or U5743 (N_5743,N_3188,N_2832);
xnor U5744 (N_5744,N_2067,N_2832);
nor U5745 (N_5745,N_2283,N_2787);
or U5746 (N_5746,N_2102,N_2417);
nand U5747 (N_5747,N_3062,N_3807);
and U5748 (N_5748,N_3693,N_2806);
and U5749 (N_5749,N_2245,N_3872);
and U5750 (N_5750,N_3489,N_3814);
or U5751 (N_5751,N_2523,N_2070);
or U5752 (N_5752,N_3138,N_2259);
xor U5753 (N_5753,N_2845,N_3796);
xnor U5754 (N_5754,N_3582,N_2831);
nor U5755 (N_5755,N_2717,N_2648);
and U5756 (N_5756,N_2557,N_3788);
or U5757 (N_5757,N_3651,N_3698);
nor U5758 (N_5758,N_2891,N_2352);
nand U5759 (N_5759,N_3192,N_3722);
or U5760 (N_5760,N_3447,N_3196);
nand U5761 (N_5761,N_2429,N_3133);
nor U5762 (N_5762,N_3973,N_2367);
nand U5763 (N_5763,N_2192,N_3323);
or U5764 (N_5764,N_2536,N_3046);
nor U5765 (N_5765,N_2241,N_3311);
and U5766 (N_5766,N_3880,N_2840);
nor U5767 (N_5767,N_2619,N_2669);
and U5768 (N_5768,N_3941,N_2815);
or U5769 (N_5769,N_2587,N_2070);
nor U5770 (N_5770,N_2482,N_3417);
nand U5771 (N_5771,N_2071,N_3531);
and U5772 (N_5772,N_3414,N_2833);
or U5773 (N_5773,N_2654,N_2252);
or U5774 (N_5774,N_2298,N_2840);
or U5775 (N_5775,N_3634,N_2294);
xnor U5776 (N_5776,N_3296,N_2811);
nand U5777 (N_5777,N_3420,N_3665);
nand U5778 (N_5778,N_3777,N_2301);
xor U5779 (N_5779,N_2384,N_2922);
nor U5780 (N_5780,N_2303,N_3603);
or U5781 (N_5781,N_2538,N_3026);
nand U5782 (N_5782,N_2795,N_3269);
and U5783 (N_5783,N_3492,N_2767);
and U5784 (N_5784,N_3630,N_3803);
nor U5785 (N_5785,N_2408,N_3584);
or U5786 (N_5786,N_2723,N_2408);
nor U5787 (N_5787,N_2964,N_2832);
and U5788 (N_5788,N_3596,N_3368);
nor U5789 (N_5789,N_2151,N_2667);
nand U5790 (N_5790,N_2428,N_2606);
xor U5791 (N_5791,N_2992,N_3664);
and U5792 (N_5792,N_3570,N_2515);
or U5793 (N_5793,N_2413,N_2944);
nand U5794 (N_5794,N_2680,N_3744);
and U5795 (N_5795,N_3323,N_2735);
nor U5796 (N_5796,N_2334,N_3636);
nand U5797 (N_5797,N_2190,N_2330);
xnor U5798 (N_5798,N_2464,N_2752);
and U5799 (N_5799,N_3357,N_2878);
nand U5800 (N_5800,N_3334,N_2407);
nor U5801 (N_5801,N_2952,N_3245);
nand U5802 (N_5802,N_2071,N_3365);
and U5803 (N_5803,N_2076,N_2320);
and U5804 (N_5804,N_2900,N_2739);
nor U5805 (N_5805,N_3142,N_3342);
nand U5806 (N_5806,N_3969,N_3966);
xor U5807 (N_5807,N_2351,N_2014);
nor U5808 (N_5808,N_2069,N_3144);
nand U5809 (N_5809,N_2822,N_3399);
nor U5810 (N_5810,N_3990,N_3548);
nand U5811 (N_5811,N_3014,N_3448);
nor U5812 (N_5812,N_3309,N_2192);
xor U5813 (N_5813,N_3488,N_2798);
nand U5814 (N_5814,N_2028,N_2334);
and U5815 (N_5815,N_2516,N_2304);
nor U5816 (N_5816,N_3633,N_3481);
and U5817 (N_5817,N_3521,N_2582);
nand U5818 (N_5818,N_2716,N_2503);
and U5819 (N_5819,N_2272,N_2113);
nand U5820 (N_5820,N_3541,N_3797);
or U5821 (N_5821,N_2024,N_2012);
xor U5822 (N_5822,N_3253,N_2292);
or U5823 (N_5823,N_3177,N_3271);
nor U5824 (N_5824,N_2923,N_2298);
nor U5825 (N_5825,N_2273,N_3075);
nor U5826 (N_5826,N_3283,N_3431);
or U5827 (N_5827,N_3025,N_2090);
nand U5828 (N_5828,N_2530,N_3549);
nor U5829 (N_5829,N_3721,N_3378);
or U5830 (N_5830,N_2194,N_3250);
nor U5831 (N_5831,N_3971,N_2310);
or U5832 (N_5832,N_2182,N_2230);
nor U5833 (N_5833,N_3512,N_2920);
or U5834 (N_5834,N_3106,N_2858);
and U5835 (N_5835,N_3002,N_3296);
or U5836 (N_5836,N_2820,N_3843);
or U5837 (N_5837,N_3694,N_2663);
and U5838 (N_5838,N_2290,N_3299);
and U5839 (N_5839,N_2037,N_3038);
and U5840 (N_5840,N_2814,N_2930);
nand U5841 (N_5841,N_2034,N_2706);
or U5842 (N_5842,N_2045,N_2788);
nand U5843 (N_5843,N_3366,N_2353);
nand U5844 (N_5844,N_2479,N_2252);
nand U5845 (N_5845,N_2992,N_2364);
xnor U5846 (N_5846,N_3913,N_3093);
nor U5847 (N_5847,N_3737,N_3294);
xnor U5848 (N_5848,N_2686,N_3839);
or U5849 (N_5849,N_2565,N_3849);
nand U5850 (N_5850,N_3624,N_2436);
and U5851 (N_5851,N_2540,N_2687);
nand U5852 (N_5852,N_2023,N_3040);
or U5853 (N_5853,N_3201,N_2209);
or U5854 (N_5854,N_2587,N_2912);
or U5855 (N_5855,N_2975,N_2816);
nand U5856 (N_5856,N_2011,N_3893);
nor U5857 (N_5857,N_2527,N_2962);
nor U5858 (N_5858,N_2106,N_2069);
xnor U5859 (N_5859,N_2422,N_3515);
nand U5860 (N_5860,N_2013,N_2741);
nor U5861 (N_5861,N_2398,N_2253);
nor U5862 (N_5862,N_2045,N_3930);
xnor U5863 (N_5863,N_3052,N_3004);
and U5864 (N_5864,N_2455,N_3818);
xor U5865 (N_5865,N_2224,N_2574);
nand U5866 (N_5866,N_3486,N_3849);
or U5867 (N_5867,N_2106,N_3025);
xnor U5868 (N_5868,N_2342,N_2058);
or U5869 (N_5869,N_3136,N_3926);
nor U5870 (N_5870,N_2129,N_3168);
nor U5871 (N_5871,N_2133,N_3902);
and U5872 (N_5872,N_3166,N_2793);
and U5873 (N_5873,N_2362,N_3959);
and U5874 (N_5874,N_2786,N_2544);
and U5875 (N_5875,N_2632,N_3913);
and U5876 (N_5876,N_3969,N_2511);
nand U5877 (N_5877,N_2156,N_2387);
xor U5878 (N_5878,N_3300,N_2242);
xor U5879 (N_5879,N_3555,N_2235);
xor U5880 (N_5880,N_3452,N_2240);
and U5881 (N_5881,N_2776,N_3938);
nand U5882 (N_5882,N_3940,N_2385);
and U5883 (N_5883,N_3530,N_2657);
and U5884 (N_5884,N_3963,N_2506);
nor U5885 (N_5885,N_2319,N_2505);
nor U5886 (N_5886,N_2058,N_2685);
nor U5887 (N_5887,N_3826,N_3638);
or U5888 (N_5888,N_2114,N_2057);
nor U5889 (N_5889,N_3655,N_3104);
nand U5890 (N_5890,N_2833,N_2723);
nor U5891 (N_5891,N_2474,N_2993);
and U5892 (N_5892,N_2208,N_2608);
xor U5893 (N_5893,N_2960,N_3049);
and U5894 (N_5894,N_3430,N_2509);
nor U5895 (N_5895,N_3944,N_3120);
and U5896 (N_5896,N_3993,N_2028);
nor U5897 (N_5897,N_2114,N_3910);
xnor U5898 (N_5898,N_3097,N_2288);
and U5899 (N_5899,N_2918,N_2517);
nor U5900 (N_5900,N_3412,N_2260);
nand U5901 (N_5901,N_3217,N_3890);
and U5902 (N_5902,N_2319,N_2880);
and U5903 (N_5903,N_2788,N_3260);
or U5904 (N_5904,N_2755,N_3789);
and U5905 (N_5905,N_3962,N_2264);
nand U5906 (N_5906,N_2500,N_3932);
and U5907 (N_5907,N_3256,N_3173);
or U5908 (N_5908,N_3230,N_3308);
and U5909 (N_5909,N_3138,N_2146);
nand U5910 (N_5910,N_3087,N_2676);
xnor U5911 (N_5911,N_3740,N_2703);
nand U5912 (N_5912,N_3087,N_3816);
or U5913 (N_5913,N_3131,N_3250);
and U5914 (N_5914,N_2064,N_2885);
or U5915 (N_5915,N_2512,N_3938);
nor U5916 (N_5916,N_2750,N_3583);
and U5917 (N_5917,N_2031,N_2873);
or U5918 (N_5918,N_2947,N_3920);
nand U5919 (N_5919,N_3764,N_3237);
nor U5920 (N_5920,N_2433,N_2158);
xnor U5921 (N_5921,N_2080,N_2152);
or U5922 (N_5922,N_2201,N_2871);
and U5923 (N_5923,N_3096,N_2896);
nand U5924 (N_5924,N_3844,N_3933);
or U5925 (N_5925,N_2832,N_3498);
nor U5926 (N_5926,N_3630,N_2899);
and U5927 (N_5927,N_3955,N_2739);
nand U5928 (N_5928,N_2501,N_3482);
nor U5929 (N_5929,N_2885,N_2475);
nand U5930 (N_5930,N_3045,N_2972);
or U5931 (N_5931,N_3766,N_3900);
xor U5932 (N_5932,N_2763,N_2246);
nand U5933 (N_5933,N_2063,N_2770);
and U5934 (N_5934,N_3869,N_2731);
nand U5935 (N_5935,N_3133,N_3694);
or U5936 (N_5936,N_2515,N_2593);
nor U5937 (N_5937,N_3695,N_2657);
nor U5938 (N_5938,N_3997,N_2007);
nor U5939 (N_5939,N_2937,N_2868);
xor U5940 (N_5940,N_2267,N_2365);
or U5941 (N_5941,N_3643,N_2303);
and U5942 (N_5942,N_2166,N_2440);
nor U5943 (N_5943,N_3345,N_2054);
nor U5944 (N_5944,N_2860,N_2115);
nand U5945 (N_5945,N_3397,N_2506);
nand U5946 (N_5946,N_2718,N_3185);
or U5947 (N_5947,N_3913,N_3229);
and U5948 (N_5948,N_2529,N_3999);
nor U5949 (N_5949,N_3565,N_2359);
or U5950 (N_5950,N_2952,N_2851);
xnor U5951 (N_5951,N_2795,N_3986);
nor U5952 (N_5952,N_2075,N_2468);
and U5953 (N_5953,N_2958,N_3697);
nand U5954 (N_5954,N_3691,N_2004);
and U5955 (N_5955,N_2067,N_3679);
or U5956 (N_5956,N_2520,N_3715);
nand U5957 (N_5957,N_2351,N_2198);
nor U5958 (N_5958,N_3998,N_2939);
xor U5959 (N_5959,N_3720,N_3951);
nand U5960 (N_5960,N_2022,N_3982);
or U5961 (N_5961,N_2264,N_2816);
nor U5962 (N_5962,N_3038,N_2415);
nand U5963 (N_5963,N_2560,N_2153);
nor U5964 (N_5964,N_3975,N_2242);
nor U5965 (N_5965,N_2035,N_2163);
or U5966 (N_5966,N_2620,N_2768);
nor U5967 (N_5967,N_3673,N_3204);
and U5968 (N_5968,N_3179,N_3241);
xor U5969 (N_5969,N_2396,N_3904);
and U5970 (N_5970,N_2834,N_3196);
and U5971 (N_5971,N_3940,N_3493);
and U5972 (N_5972,N_3205,N_3033);
or U5973 (N_5973,N_3162,N_2864);
or U5974 (N_5974,N_2162,N_2608);
nand U5975 (N_5975,N_3639,N_2165);
nor U5976 (N_5976,N_3362,N_3305);
xnor U5977 (N_5977,N_3342,N_3101);
nand U5978 (N_5978,N_2242,N_3919);
and U5979 (N_5979,N_2811,N_3056);
and U5980 (N_5980,N_2675,N_3335);
or U5981 (N_5981,N_2416,N_3675);
nand U5982 (N_5982,N_2887,N_3442);
xor U5983 (N_5983,N_3510,N_3220);
nor U5984 (N_5984,N_3348,N_3817);
xnor U5985 (N_5985,N_2834,N_2245);
xor U5986 (N_5986,N_3236,N_3661);
and U5987 (N_5987,N_3676,N_3142);
nand U5988 (N_5988,N_2589,N_2167);
nor U5989 (N_5989,N_3261,N_3859);
nor U5990 (N_5990,N_3065,N_2767);
or U5991 (N_5991,N_2797,N_3402);
or U5992 (N_5992,N_2736,N_2654);
nand U5993 (N_5993,N_2004,N_2653);
and U5994 (N_5994,N_2567,N_2041);
xor U5995 (N_5995,N_2623,N_3428);
nor U5996 (N_5996,N_3618,N_2376);
xnor U5997 (N_5997,N_3149,N_2580);
xor U5998 (N_5998,N_3821,N_3438);
or U5999 (N_5999,N_3428,N_2083);
and U6000 (N_6000,N_5510,N_5551);
or U6001 (N_6001,N_5140,N_5371);
nand U6002 (N_6002,N_4924,N_4521);
and U6003 (N_6003,N_4442,N_4239);
nand U6004 (N_6004,N_4447,N_5192);
nor U6005 (N_6005,N_4934,N_5154);
or U6006 (N_6006,N_5022,N_5642);
nor U6007 (N_6007,N_4629,N_5345);
and U6008 (N_6008,N_4203,N_5983);
nand U6009 (N_6009,N_5786,N_4036);
nor U6010 (N_6010,N_4328,N_5383);
nand U6011 (N_6011,N_4723,N_5266);
xnor U6012 (N_6012,N_5655,N_5379);
nand U6013 (N_6013,N_5248,N_4769);
or U6014 (N_6014,N_5390,N_5298);
nor U6015 (N_6015,N_4621,N_5305);
and U6016 (N_6016,N_5450,N_4309);
or U6017 (N_6017,N_4334,N_4816);
and U6018 (N_6018,N_4730,N_4979);
nor U6019 (N_6019,N_4454,N_5168);
nor U6020 (N_6020,N_5189,N_5744);
and U6021 (N_6021,N_4133,N_5948);
nor U6022 (N_6022,N_4500,N_5087);
xnor U6023 (N_6023,N_4079,N_4834);
nand U6024 (N_6024,N_4619,N_5414);
or U6025 (N_6025,N_5497,N_4918);
and U6026 (N_6026,N_4611,N_4717);
nor U6027 (N_6027,N_4245,N_5963);
or U6028 (N_6028,N_5541,N_4909);
xnor U6029 (N_6029,N_4364,N_5552);
nor U6030 (N_6030,N_5892,N_4960);
nor U6031 (N_6031,N_5943,N_4242);
xnor U6032 (N_6032,N_4803,N_4917);
and U6033 (N_6033,N_5748,N_4468);
and U6034 (N_6034,N_4708,N_5994);
nand U6035 (N_6035,N_4870,N_5188);
and U6036 (N_6036,N_5091,N_5002);
nand U6037 (N_6037,N_4138,N_5712);
nor U6038 (N_6038,N_5187,N_5324);
or U6039 (N_6039,N_5025,N_5727);
and U6040 (N_6040,N_5207,N_5129);
or U6041 (N_6041,N_5709,N_4487);
nor U6042 (N_6042,N_4386,N_5098);
and U6043 (N_6043,N_4658,N_4096);
and U6044 (N_6044,N_4008,N_5708);
or U6045 (N_6045,N_5054,N_5910);
nor U6046 (N_6046,N_4162,N_5469);
nor U6047 (N_6047,N_4434,N_5805);
nor U6048 (N_6048,N_4012,N_4617);
and U6049 (N_6049,N_5279,N_4380);
and U6050 (N_6050,N_4940,N_5592);
nand U6051 (N_6051,N_4076,N_4910);
nor U6052 (N_6052,N_4888,N_4033);
nand U6053 (N_6053,N_5840,N_4171);
nand U6054 (N_6054,N_5882,N_4831);
nor U6055 (N_6055,N_5156,N_4892);
nor U6056 (N_6056,N_4954,N_5215);
or U6057 (N_6057,N_5494,N_5504);
and U6058 (N_6058,N_5619,N_4211);
nor U6059 (N_6059,N_5594,N_5825);
nand U6060 (N_6060,N_4990,N_4928);
or U6061 (N_6061,N_5981,N_4484);
xnor U6062 (N_6062,N_5785,N_4665);
xnor U6063 (N_6063,N_4431,N_4516);
nand U6064 (N_6064,N_5901,N_5011);
nand U6065 (N_6065,N_4677,N_5564);
xnor U6066 (N_6066,N_5627,N_5496);
or U6067 (N_6067,N_4369,N_4119);
nor U6068 (N_6068,N_4457,N_4824);
and U6069 (N_6069,N_4382,N_4958);
nand U6070 (N_6070,N_4913,N_4968);
nand U6071 (N_6071,N_5665,N_4950);
xnor U6072 (N_6072,N_5881,N_4525);
nand U6073 (N_6073,N_4664,N_5615);
or U6074 (N_6074,N_4361,N_4575);
nor U6075 (N_6075,N_4017,N_5687);
and U6076 (N_6076,N_5257,N_5718);
or U6077 (N_6077,N_4517,N_4202);
or U6078 (N_6078,N_4949,N_4763);
xor U6079 (N_6079,N_4337,N_5788);
nor U6080 (N_6080,N_4214,N_4276);
xnor U6081 (N_6081,N_5449,N_4438);
nand U6082 (N_6082,N_4445,N_5139);
nand U6083 (N_6083,N_4105,N_4261);
nor U6084 (N_6084,N_4603,N_5124);
xnor U6085 (N_6085,N_4626,N_4196);
or U6086 (N_6086,N_5406,N_5155);
or U6087 (N_6087,N_5194,N_4741);
or U6088 (N_6088,N_5782,N_4493);
nor U6089 (N_6089,N_4240,N_5427);
nor U6090 (N_6090,N_5766,N_4994);
and U6091 (N_6091,N_4419,N_4078);
nand U6092 (N_6092,N_5136,N_4997);
nor U6093 (N_6093,N_4344,N_5268);
nand U6094 (N_6094,N_5763,N_5164);
and U6095 (N_6095,N_5012,N_5259);
xnor U6096 (N_6096,N_4121,N_5440);
and U6097 (N_6097,N_5070,N_4872);
nor U6098 (N_6098,N_5149,N_4800);
xor U6099 (N_6099,N_4103,N_5082);
or U6100 (N_6100,N_5921,N_5031);
and U6101 (N_6101,N_5680,N_5018);
xor U6102 (N_6102,N_5009,N_4312);
nand U6103 (N_6103,N_4537,N_4955);
nor U6104 (N_6104,N_5442,N_5620);
nor U6105 (N_6105,N_5354,N_5797);
or U6106 (N_6106,N_4244,N_4785);
xnor U6107 (N_6107,N_4869,N_5833);
and U6108 (N_6108,N_5728,N_4791);
or U6109 (N_6109,N_4554,N_5784);
nand U6110 (N_6110,N_4031,N_5213);
nor U6111 (N_6111,N_5545,N_4465);
and U6112 (N_6112,N_5978,N_5696);
nor U6113 (N_6113,N_4993,N_4897);
and U6114 (N_6114,N_4404,N_5090);
and U6115 (N_6115,N_5692,N_4336);
or U6116 (N_6116,N_5099,N_4023);
nand U6117 (N_6117,N_5411,N_4674);
and U6118 (N_6118,N_5720,N_5398);
nand U6119 (N_6119,N_4106,N_5919);
or U6120 (N_6120,N_5794,N_5618);
xor U6121 (N_6121,N_4426,N_5484);
nor U6122 (N_6122,N_5446,N_4347);
or U6123 (N_6123,N_5804,N_5894);
and U6124 (N_6124,N_5451,N_4945);
nor U6125 (N_6125,N_4594,N_5181);
and U6126 (N_6126,N_4698,N_4802);
and U6127 (N_6127,N_5830,N_4020);
xnor U6128 (N_6128,N_5509,N_4855);
nor U6129 (N_6129,N_5348,N_5483);
or U6130 (N_6130,N_4004,N_4243);
nand U6131 (N_6131,N_4375,N_4030);
xor U6132 (N_6132,N_5112,N_5227);
and U6133 (N_6133,N_4123,N_4736);
nor U6134 (N_6134,N_4670,N_4961);
nand U6135 (N_6135,N_4641,N_4164);
and U6136 (N_6136,N_5308,N_5900);
or U6137 (N_6137,N_4492,N_4673);
nand U6138 (N_6138,N_4444,N_4652);
nand U6139 (N_6139,N_4546,N_5972);
or U6140 (N_6140,N_4387,N_4970);
and U6141 (N_6141,N_4255,N_5359);
and U6142 (N_6142,N_5238,N_4901);
nand U6143 (N_6143,N_5808,N_4238);
nor U6144 (N_6144,N_4274,N_5322);
nor U6145 (N_6145,N_4304,N_4829);
and U6146 (N_6146,N_4141,N_4067);
nand U6147 (N_6147,N_5278,N_4331);
and U6148 (N_6148,N_5679,N_5838);
xor U6149 (N_6149,N_4217,N_5613);
and U6150 (N_6150,N_4174,N_5580);
and U6151 (N_6151,N_4654,N_4275);
or U6152 (N_6152,N_5740,N_4185);
or U6153 (N_6153,N_4110,N_4354);
or U6154 (N_6154,N_4421,N_5292);
or U6155 (N_6155,N_5988,N_4620);
xor U6156 (N_6156,N_5848,N_5657);
nor U6157 (N_6157,N_4727,N_4732);
nor U6158 (N_6158,N_4657,N_5173);
xor U6159 (N_6159,N_4667,N_5318);
nor U6160 (N_6160,N_4066,N_5256);
nand U6161 (N_6161,N_4204,N_4581);
and U6162 (N_6162,N_4597,N_4108);
nor U6163 (N_6163,N_5108,N_4549);
and U6164 (N_6164,N_5950,N_5057);
or U6165 (N_6165,N_5205,N_4193);
xor U6166 (N_6166,N_4942,N_4416);
xnor U6167 (N_6167,N_4571,N_5050);
nand U6168 (N_6168,N_4854,N_5745);
nand U6169 (N_6169,N_4181,N_4087);
nand U6170 (N_6170,N_5211,N_5478);
xnor U6171 (N_6171,N_5143,N_5242);
xnor U6172 (N_6172,N_5073,N_4704);
nor U6173 (N_6173,N_5210,N_5826);
nand U6174 (N_6174,N_5653,N_5179);
nor U6175 (N_6175,N_5733,N_5621);
nand U6176 (N_6176,N_5837,N_5485);
or U6177 (N_6177,N_4482,N_5925);
xnor U6178 (N_6178,N_4071,N_4653);
and U6179 (N_6179,N_4884,N_4291);
nand U6180 (N_6180,N_5384,N_4346);
and U6181 (N_6181,N_5762,N_4359);
and U6182 (N_6182,N_5066,N_4455);
or U6183 (N_6183,N_4919,N_5223);
or U6184 (N_6184,N_5357,N_5479);
nand U6185 (N_6185,N_4634,N_4021);
or U6186 (N_6186,N_5000,N_4314);
nand U6187 (N_6187,N_5967,N_4467);
nand U6188 (N_6188,N_5832,N_5218);
and U6189 (N_6189,N_5103,N_4535);
nor U6190 (N_6190,N_4464,N_4946);
and U6191 (N_6191,N_5602,N_5421);
xor U6192 (N_6192,N_4515,N_4098);
nand U6193 (N_6193,N_5037,N_5304);
and U6194 (N_6194,N_4767,N_5120);
nor U6195 (N_6195,N_4703,N_4709);
or U6196 (N_6196,N_4499,N_4906);
xnor U6197 (N_6197,N_4338,N_4750);
xnor U6198 (N_6198,N_5104,N_5917);
and U6199 (N_6199,N_4687,N_4205);
and U6200 (N_6200,N_5321,N_4357);
nand U6201 (N_6201,N_4923,N_5755);
and U6202 (N_6202,N_4018,N_5235);
nand U6203 (N_6203,N_5676,N_4230);
and U6204 (N_6204,N_5431,N_5522);
nand U6205 (N_6205,N_5019,N_5866);
and U6206 (N_6206,N_5639,N_4567);
or U6207 (N_6207,N_4456,N_4959);
or U6208 (N_6208,N_4661,N_4795);
nand U6209 (N_6209,N_4258,N_4577);
or U6210 (N_6210,N_5128,N_4413);
nand U6211 (N_6211,N_5868,N_5918);
and U6212 (N_6212,N_4887,N_4403);
nor U6213 (N_6213,N_5113,N_4579);
nand U6214 (N_6214,N_4734,N_5550);
and U6215 (N_6215,N_5577,N_4154);
nor U6216 (N_6216,N_4083,N_5058);
and U6217 (N_6217,N_4534,N_4388);
nor U6218 (N_6218,N_5625,N_5052);
nor U6219 (N_6219,N_5616,N_5284);
or U6220 (N_6220,N_4398,N_5400);
or U6221 (N_6221,N_5820,N_4084);
nand U6222 (N_6222,N_5335,N_5372);
nand U6223 (N_6223,N_4859,N_5407);
nor U6224 (N_6224,N_5971,N_5824);
nand U6225 (N_6225,N_5117,N_5003);
or U6226 (N_6226,N_4995,N_4695);
nor U6227 (N_6227,N_4893,N_4144);
or U6228 (N_6228,N_5387,N_4801);
or U6229 (N_6229,N_4013,N_4784);
and U6230 (N_6230,N_4998,N_5017);
or U6231 (N_6231,N_4541,N_4596);
nand U6232 (N_6232,N_4074,N_5628);
xor U6233 (N_6233,N_5691,N_4749);
and U6234 (N_6234,N_5929,N_5204);
or U6235 (N_6235,N_5638,N_4268);
and U6236 (N_6236,N_4390,N_4035);
nor U6237 (N_6237,N_4285,N_5699);
nor U6238 (N_6238,N_5893,N_5317);
or U6239 (N_6239,N_5883,N_5700);
or U6240 (N_6240,N_5968,N_5723);
and U6241 (N_6241,N_5264,N_4095);
nor U6242 (N_6242,N_4234,N_4927);
or U6243 (N_6243,N_4809,N_5077);
nor U6244 (N_6244,N_4980,N_5314);
and U6245 (N_6245,N_4117,N_4552);
and U6246 (N_6246,N_4757,N_4322);
or U6247 (N_6247,N_5481,N_5942);
and U6248 (N_6248,N_5729,N_4853);
and U6249 (N_6249,N_4780,N_4828);
nor U6250 (N_6250,N_4418,N_5144);
nor U6251 (N_6251,N_4006,N_5675);
or U6252 (N_6252,N_4570,N_4000);
nand U6253 (N_6253,N_4401,N_4064);
nor U6254 (N_6254,N_4218,N_4574);
xor U6255 (N_6255,N_5222,N_4297);
xnor U6256 (N_6256,N_4608,N_4964);
xnor U6257 (N_6257,N_5206,N_4489);
or U6258 (N_6258,N_4175,N_5374);
nor U6259 (N_6259,N_5548,N_5589);
or U6260 (N_6260,N_4700,N_4632);
nand U6261 (N_6261,N_5876,N_5896);
and U6262 (N_6262,N_5097,N_4811);
nand U6263 (N_6263,N_4206,N_4545);
nor U6264 (N_6264,N_4102,N_5578);
nor U6265 (N_6265,N_4935,N_4520);
nand U6266 (N_6266,N_5319,N_4472);
nand U6267 (N_6267,N_4786,N_4441);
and U6268 (N_6268,N_4151,N_4225);
nor U6269 (N_6269,N_5587,N_4410);
nor U6270 (N_6270,N_5734,N_5851);
nor U6271 (N_6271,N_4057,N_4663);
and U6272 (N_6272,N_4335,N_4782);
xnor U6273 (N_6273,N_5637,N_4055);
and U6274 (N_6274,N_5342,N_5899);
nor U6275 (N_6275,N_5915,N_4560);
nor U6276 (N_6276,N_4898,N_5669);
or U6277 (N_6277,N_5475,N_5062);
nand U6278 (N_6278,N_4481,N_4015);
nor U6279 (N_6279,N_5861,N_4622);
or U6280 (N_6280,N_5287,N_5874);
nor U6281 (N_6281,N_4048,N_4425);
and U6282 (N_6282,N_5521,N_5579);
or U6283 (N_6283,N_5375,N_5448);
nand U6284 (N_6284,N_5422,N_4556);
or U6285 (N_6285,N_5373,N_4179);
nand U6286 (N_6286,N_5034,N_4792);
nand U6287 (N_6287,N_4407,N_4944);
nor U6288 (N_6288,N_4975,N_5749);
or U6289 (N_6289,N_5518,N_4682);
or U6290 (N_6290,N_4436,N_4532);
xnor U6291 (N_6291,N_5500,N_4394);
and U6292 (N_6292,N_5366,N_4042);
nor U6293 (N_6293,N_5531,N_4298);
nor U6294 (N_6294,N_5631,N_5358);
nand U6295 (N_6295,N_4109,N_5739);
nor U6296 (N_6296,N_5429,N_4005);
xnor U6297 (N_6297,N_5081,N_5460);
xnor U6298 (N_6298,N_4273,N_5936);
nand U6299 (N_6299,N_5307,N_4903);
nand U6300 (N_6300,N_4424,N_5228);
xnor U6301 (N_6301,N_5269,N_4733);
or U6302 (N_6302,N_5557,N_5293);
xnor U6303 (N_6303,N_5080,N_4348);
and U6304 (N_6304,N_4406,N_5309);
nand U6305 (N_6305,N_4982,N_5150);
xor U6306 (N_6306,N_4999,N_5320);
xnor U6307 (N_6307,N_5562,N_5757);
or U6308 (N_6308,N_4702,N_4894);
nand U6309 (N_6309,N_4576,N_5132);
and U6310 (N_6310,N_4987,N_4052);
or U6311 (N_6311,N_4862,N_5474);
nand U6312 (N_6312,N_5495,N_4877);
and U6313 (N_6313,N_4415,N_5667);
and U6314 (N_6314,N_5355,N_5294);
or U6315 (N_6315,N_5076,N_5525);
nor U6316 (N_6316,N_4967,N_5068);
and U6317 (N_6317,N_5296,N_5672);
and U6318 (N_6318,N_4253,N_4091);
or U6319 (N_6319,N_5890,N_5368);
nor U6320 (N_6320,N_5116,N_4192);
nor U6321 (N_6321,N_5905,N_5554);
and U6322 (N_6322,N_4743,N_4397);
nand U6323 (N_6323,N_5928,N_4186);
and U6324 (N_6324,N_5549,N_4029);
or U6325 (N_6325,N_4644,N_4257);
and U6326 (N_6326,N_5581,N_4317);
nor U6327 (N_6327,N_4219,N_4966);
nor U6328 (N_6328,N_5724,N_5752);
or U6329 (N_6329,N_4799,N_5225);
nor U6330 (N_6330,N_5865,N_5172);
nand U6331 (N_6331,N_4272,N_4662);
and U6332 (N_6332,N_4776,N_4878);
nand U6333 (N_6333,N_5529,N_4080);
xnor U6334 (N_6334,N_4719,N_4453);
nand U6335 (N_6335,N_5538,N_5847);
nand U6336 (N_6336,N_4396,N_4473);
nand U6337 (N_6337,N_4319,N_5347);
or U6338 (N_6338,N_5499,N_5490);
nand U6339 (N_6339,N_5349,N_4435);
nor U6340 (N_6340,N_5770,N_5078);
nor U6341 (N_6341,N_5853,N_4639);
nand U6342 (N_6342,N_5491,N_5392);
nor U6343 (N_6343,N_4922,N_5167);
and U6344 (N_6344,N_5244,N_5245);
or U6345 (N_6345,N_5059,N_5710);
or U6346 (N_6346,N_5773,N_4235);
and U6347 (N_6347,N_4778,N_4058);
nand U6348 (N_6348,N_5523,N_4921);
nor U6349 (N_6349,N_4583,N_5362);
xor U6350 (N_6350,N_5378,N_4810);
nand U6351 (N_6351,N_5444,N_4953);
and U6352 (N_6352,N_4787,N_5630);
nor U6353 (N_6353,N_4460,N_5004);
and U6354 (N_6354,N_4139,N_4718);
nand U6355 (N_6355,N_5998,N_4490);
or U6356 (N_6356,N_5817,N_5644);
and U6357 (N_6357,N_4104,N_5870);
nand U6358 (N_6358,N_4405,N_4009);
nand U6359 (N_6359,N_5771,N_5191);
nor U6360 (N_6360,N_5193,N_4548);
nor U6361 (N_6361,N_4610,N_4303);
nor U6362 (N_6362,N_5835,N_4601);
and U6363 (N_6363,N_5024,N_4260);
and U6364 (N_6364,N_4937,N_5743);
nor U6365 (N_6365,N_5323,N_4201);
or U6366 (N_6366,N_5722,N_4773);
xor U6367 (N_6367,N_4153,N_5694);
and U6368 (N_6368,N_5015,N_5419);
nor U6369 (N_6369,N_5420,N_4378);
and U6370 (N_6370,N_5243,N_4737);
or U6371 (N_6371,N_5877,N_5666);
nand U6372 (N_6372,N_5711,N_4696);
nor U6373 (N_6373,N_5588,N_5836);
nand U6374 (N_6374,N_4222,N_5965);
and U6375 (N_6375,N_5732,N_4002);
nand U6376 (N_6376,N_4759,N_4485);
or U6377 (N_6377,N_4930,N_4886);
nor U6378 (N_6378,N_4805,N_5267);
or U6379 (N_6379,N_4650,N_4614);
nor U6380 (N_6380,N_5539,N_4666);
nand U6381 (N_6381,N_4318,N_5986);
and U6382 (N_6382,N_5604,N_5127);
nor U6383 (N_6383,N_5337,N_5783);
nand U6384 (N_6384,N_5707,N_4631);
nor U6385 (N_6385,N_4858,N_5585);
nand U6386 (N_6386,N_5612,N_4299);
or U6387 (N_6387,N_5084,N_5693);
and U6388 (N_6388,N_5964,N_5470);
nand U6389 (N_6389,N_4561,N_5923);
and U6390 (N_6390,N_4353,N_5535);
nand U6391 (N_6391,N_4478,N_4362);
and U6392 (N_6392,N_5831,N_5537);
nand U6393 (N_6393,N_5394,N_4228);
nand U6394 (N_6394,N_4073,N_4059);
nor U6395 (N_6395,N_4963,N_4511);
nor U6396 (N_6396,N_5110,N_5561);
and U6397 (N_6397,N_4598,N_5746);
and U6398 (N_6398,N_4093,N_5975);
xor U6399 (N_6399,N_5106,N_5717);
xor U6400 (N_6400,N_5131,N_5775);
xnor U6401 (N_6401,N_4606,N_4086);
or U6402 (N_6402,N_5041,N_4705);
xnor U6403 (N_6403,N_4374,N_5403);
and U6404 (N_6404,N_4132,N_4324);
or U6405 (N_6405,N_5032,N_5536);
and U6406 (N_6406,N_5895,N_5731);
nand U6407 (N_6407,N_5114,N_4783);
nand U6408 (N_6408,N_5089,N_4756);
nor U6409 (N_6409,N_5290,N_5258);
or U6410 (N_6410,N_5043,N_4728);
and U6411 (N_6411,N_5512,N_4250);
nor U6412 (N_6412,N_4145,N_4840);
or U6413 (N_6413,N_4259,N_4300);
nor U6414 (N_6414,N_5195,N_4136);
nand U6415 (N_6415,N_5532,N_5741);
nor U6416 (N_6416,N_5811,N_4720);
or U6417 (N_6417,N_4724,N_5385);
xor U6418 (N_6418,N_5789,N_4069);
or U6419 (N_6419,N_4879,N_5664);
nand U6420 (N_6420,N_5813,N_4962);
nand U6421 (N_6421,N_4830,N_4936);
or U6422 (N_6422,N_4645,N_4707);
nor U6423 (N_6423,N_5199,N_4758);
nand U6424 (N_6424,N_5802,N_4533);
xnor U6425 (N_6425,N_4981,N_5563);
and U6426 (N_6426,N_4871,N_4262);
nor U6427 (N_6427,N_4867,N_5586);
nand U6428 (N_6428,N_5064,N_5315);
and U6429 (N_6429,N_4458,N_5683);
xor U6430 (N_6430,N_4412,N_4107);
and U6431 (N_6431,N_5288,N_5916);
nand U6432 (N_6432,N_5095,N_5914);
or U6433 (N_6433,N_4061,N_4060);
or U6434 (N_6434,N_4494,N_5331);
xnor U6435 (N_6435,N_4125,N_5458);
nor U6436 (N_6436,N_4555,N_4739);
nand U6437 (N_6437,N_5996,N_5856);
and U6438 (N_6438,N_5568,N_5013);
or U6439 (N_6439,N_4292,N_4340);
nor U6440 (N_6440,N_5884,N_4627);
or U6441 (N_6441,N_4127,N_4835);
and U6442 (N_6442,N_5208,N_4774);
and U6443 (N_6443,N_4325,N_5935);
or U6444 (N_6444,N_5338,N_5505);
xor U6445 (N_6445,N_5626,N_5945);
nor U6446 (N_6446,N_5750,N_5949);
nand U6447 (N_6447,N_4408,N_5955);
xnor U6448 (N_6448,N_4316,N_4540);
or U6449 (N_6449,N_4129,N_4607);
and U6450 (N_6450,N_4158,N_4089);
xor U6451 (N_6451,N_4553,N_5410);
nand U6452 (N_6452,N_4355,N_5133);
nand U6453 (N_6453,N_4563,N_4251);
nor U6454 (N_6454,N_5938,N_5854);
xnor U6455 (N_6455,N_5363,N_4342);
nand U6456 (N_6456,N_5897,N_4475);
nor U6457 (N_6457,N_4715,N_5931);
and U6458 (N_6458,N_5169,N_4600);
nand U6459 (N_6459,N_5688,N_4011);
xnor U6460 (N_6460,N_4024,N_5190);
xnor U6461 (N_6461,N_4523,N_4648);
nor U6462 (N_6462,N_5163,N_5962);
or U6463 (N_6463,N_5697,N_4822);
or U6464 (N_6464,N_4655,N_5203);
nor U6465 (N_6465,N_4689,N_5767);
nor U6466 (N_6466,N_4081,N_5200);
nand U6467 (N_6467,N_5232,N_5682);
nor U6468 (N_6468,N_4977,N_4122);
or U6469 (N_6469,N_4860,N_5467);
xnor U6470 (N_6470,N_4832,N_5333);
nor U6471 (N_6471,N_4628,N_5969);
and U6472 (N_6472,N_5647,N_4678);
xor U6473 (N_6473,N_5624,N_5889);
nand U6474 (N_6474,N_5715,N_5486);
or U6475 (N_6475,N_5888,N_5170);
nand U6476 (N_6476,N_4462,N_5085);
or U6477 (N_6477,N_4088,N_5800);
nor U6478 (N_6478,N_4047,N_5803);
nor U6479 (N_6479,N_4040,N_4184);
xnor U6480 (N_6480,N_4593,N_5932);
and U6481 (N_6481,N_4680,N_5607);
or U6482 (N_6482,N_5216,N_4165);
and U6483 (N_6483,N_5596,N_5356);
and U6484 (N_6484,N_5381,N_4310);
and U6485 (N_6485,N_5472,N_5301);
nand U6486 (N_6486,N_5844,N_5247);
and U6487 (N_6487,N_5903,N_5241);
or U6488 (N_6488,N_4167,N_4505);
nand U6489 (N_6489,N_4735,N_4159);
and U6490 (N_6490,N_5273,N_5121);
xor U6491 (N_6491,N_4085,N_4908);
or U6492 (N_6492,N_4329,N_4544);
xnor U6493 (N_6493,N_4818,N_5751);
and U6494 (N_6494,N_5343,N_5941);
and U6495 (N_6495,N_4745,N_4497);
xnor U6496 (N_6496,N_4714,N_4542);
and U6497 (N_6497,N_4320,N_4573);
or U6498 (N_6498,N_5622,N_5134);
and U6499 (N_6499,N_5435,N_4740);
xnor U6500 (N_6500,N_4941,N_5524);
or U6501 (N_6501,N_4512,N_4459);
or U6502 (N_6502,N_5482,N_5262);
and U6503 (N_6503,N_4543,N_5777);
or U6504 (N_6504,N_4932,N_5790);
nand U6505 (N_6505,N_4446,N_4417);
or U6506 (N_6506,N_4246,N_5927);
or U6507 (N_6507,N_4014,N_4651);
and U6508 (N_6508,N_5061,N_5507);
nand U6509 (N_6509,N_5437,N_4989);
or U6510 (N_6510,N_5001,N_5135);
xnor U6511 (N_6511,N_5702,N_4178);
and U6512 (N_6512,N_4269,N_4643);
and U6513 (N_6513,N_5401,N_5265);
or U6514 (N_6514,N_4926,N_5648);
or U6515 (N_6515,N_4642,N_4207);
nand U6516 (N_6516,N_5142,N_4001);
and U6517 (N_6517,N_4220,N_5416);
nor U6518 (N_6518,N_5300,N_5516);
nand U6519 (N_6519,N_5547,N_5063);
nor U6520 (N_6520,N_5633,N_4028);
xor U6521 (N_6521,N_4191,N_5328);
or U6522 (N_6522,N_5159,N_4474);
or U6523 (N_6523,N_5380,N_5040);
nand U6524 (N_6524,N_4812,N_4393);
and U6525 (N_6525,N_4823,N_4983);
nor U6526 (N_6526,N_4504,N_4615);
nand U6527 (N_6527,N_4659,N_4278);
or U6528 (N_6528,N_5270,N_5461);
and U6529 (N_6529,N_4379,N_4227);
nor U6530 (N_6530,N_4041,N_4889);
and U6531 (N_6531,N_4176,N_5438);
xor U6532 (N_6532,N_4612,N_5556);
nand U6533 (N_6533,N_5958,N_4430);
nand U6534 (N_6534,N_4368,N_5489);
xnor U6535 (N_6535,N_4558,N_4180);
nand U6536 (N_6536,N_4470,N_5845);
and U6537 (N_6537,N_5542,N_5249);
or U6538 (N_6538,N_4916,N_4056);
xor U6539 (N_6539,N_4358,N_5879);
or U6540 (N_6540,N_4851,N_4383);
and U6541 (N_6541,N_4849,N_4264);
nand U6542 (N_6542,N_5850,N_5346);
or U6543 (N_6543,N_5071,N_5649);
or U6544 (N_6544,N_4559,N_4978);
or U6545 (N_6545,N_4522,N_4315);
or U6546 (N_6546,N_5079,N_5201);
or U6547 (N_6547,N_5020,N_5055);
nand U6548 (N_6548,N_5344,N_5493);
nor U6549 (N_6549,N_5984,N_4026);
and U6550 (N_6550,N_5023,N_5911);
or U6551 (N_6551,N_5862,N_4697);
and U6552 (N_6552,N_5251,N_4210);
or U6553 (N_6553,N_5441,N_4586);
xnor U6554 (N_6554,N_4531,N_5576);
nand U6555 (N_6555,N_5382,N_5202);
and U6556 (N_6556,N_5157,N_4868);
xnor U6557 (N_6557,N_5424,N_4752);
nand U6558 (N_6558,N_4373,N_5118);
or U6559 (N_6559,N_4399,N_4755);
xnor U6560 (N_6560,N_4585,N_4114);
xor U6561 (N_6561,N_4766,N_5546);
nor U6562 (N_6562,N_4433,N_4507);
and U6563 (N_6563,N_5185,N_5402);
and U6564 (N_6564,N_4863,N_4688);
nand U6565 (N_6565,N_4241,N_4635);
or U6566 (N_6566,N_4838,N_5353);
nand U6567 (N_6567,N_4701,N_5898);
nand U6568 (N_6568,N_4022,N_4671);
nand U6569 (N_6569,N_5432,N_5455);
nor U6570 (N_6570,N_4118,N_5166);
nor U6571 (N_6571,N_4848,N_5409);
or U6572 (N_6572,N_4365,N_4046);
nor U6573 (N_6573,N_4725,N_4911);
nand U6574 (N_6574,N_4395,N_4686);
or U6575 (N_6575,N_5027,N_5977);
nand U6576 (N_6576,N_5180,N_4588);
nand U6577 (N_6577,N_5920,N_4039);
nand U6578 (N_6578,N_4536,N_5428);
nand U6579 (N_6579,N_5747,N_5703);
nand U6580 (N_6580,N_5130,N_5250);
and U6581 (N_6581,N_5841,N_4813);
and U6582 (N_6582,N_5255,N_5922);
and U6583 (N_6583,N_4672,N_4270);
or U6584 (N_6584,N_4744,N_5261);
nand U6585 (N_6585,N_4305,N_5812);
or U6586 (N_6586,N_4742,N_4738);
or U6587 (N_6587,N_4895,N_4873);
or U6588 (N_6588,N_5051,N_5361);
nand U6589 (N_6589,N_4592,N_5852);
and U6590 (N_6590,N_5119,N_4905);
nor U6591 (N_6591,N_5498,N_5849);
nor U6592 (N_6592,N_4307,N_5982);
or U6593 (N_6593,N_5815,N_5859);
and U6594 (N_6594,N_5765,N_5325);
nor U6595 (N_6595,N_4508,N_4969);
or U6596 (N_6596,N_4524,N_4618);
nand U6597 (N_6597,N_5086,N_4281);
or U6598 (N_6598,N_5705,N_5719);
or U6599 (N_6599,N_5555,N_5253);
nand U6600 (N_6600,N_5875,N_4070);
nor U6601 (N_6601,N_5123,N_5176);
or U6602 (N_6602,N_4350,N_5600);
or U6603 (N_6603,N_5109,N_4748);
nor U6604 (N_6604,N_4488,N_5282);
nand U6605 (N_6605,N_4360,N_4160);
nor U6606 (N_6606,N_4630,N_5219);
nand U6607 (N_6607,N_5105,N_4694);
nand U6608 (N_6608,N_5787,N_5147);
nor U6609 (N_6609,N_5014,N_4267);
nand U6610 (N_6610,N_4351,N_4526);
nand U6611 (N_6611,N_5035,N_5280);
and U6612 (N_6612,N_5514,N_5044);
nand U6613 (N_6613,N_5721,N_4142);
and U6614 (N_6614,N_4771,N_5067);
nor U6615 (N_6615,N_4126,N_5217);
xor U6616 (N_6616,N_4874,N_5761);
or U6617 (N_6617,N_5822,N_5685);
nand U6618 (N_6618,N_5138,N_4155);
nand U6619 (N_6619,N_4134,N_5939);
nand U6620 (N_6620,N_5635,N_5569);
and U6621 (N_6621,N_4925,N_5671);
nor U6622 (N_6622,N_5178,N_5567);
or U6623 (N_6623,N_5540,N_4075);
or U6624 (N_6624,N_5033,N_4034);
nand U6625 (N_6625,N_5908,N_4506);
xor U6626 (N_6626,N_4120,N_5230);
nand U6627 (N_6627,N_5453,N_4163);
nor U6628 (N_6628,N_4301,N_4381);
and U6629 (N_6629,N_5425,N_5992);
xor U6630 (N_6630,N_4595,N_5395);
nor U6631 (N_6631,N_5303,N_4437);
and U6632 (N_6632,N_5617,N_5603);
nor U6633 (N_6633,N_5662,N_4843);
and U6634 (N_6634,N_4229,N_4483);
or U6635 (N_6635,N_4288,N_5926);
nand U6636 (N_6636,N_4770,N_4775);
nor U6637 (N_6637,N_4820,N_5674);
or U6638 (N_6638,N_4777,N_4223);
xnor U6639 (N_6639,N_5686,N_4882);
and U6640 (N_6640,N_5553,N_4194);
and U6641 (N_6641,N_4476,N_5819);
or U6642 (N_6642,N_4519,N_4152);
and U6643 (N_6643,N_4833,N_4616);
and U6644 (N_6644,N_4352,N_4450);
nor U6645 (N_6645,N_5668,N_4625);
and U6646 (N_6646,N_4876,N_4856);
nand U6647 (N_6647,N_5559,N_5756);
nor U6648 (N_6648,N_5177,N_5330);
nor U6649 (N_6649,N_4043,N_5436);
xnor U6650 (N_6650,N_5184,N_5423);
and U6651 (N_6651,N_4691,N_4166);
or U6652 (N_6652,N_5957,N_5198);
nand U6653 (N_6653,N_5220,N_5995);
or U6654 (N_6654,N_5405,N_4547);
nand U6655 (N_6655,N_4432,N_5313);
nor U6656 (N_6656,N_4951,N_4938);
nand U6657 (N_6657,N_5806,N_4638);
nand U6658 (N_6658,N_4790,N_4182);
nand U6659 (N_6659,N_4112,N_5005);
or U6660 (N_6660,N_4609,N_4195);
nor U6661 (N_6661,N_5778,N_4866);
xnor U6662 (N_6662,N_4602,N_4295);
or U6663 (N_6663,N_4568,N_5291);
nand U6664 (N_6664,N_4332,N_5158);
xor U6665 (N_6665,N_4815,N_5768);
or U6666 (N_6666,N_4692,N_4414);
and U6667 (N_6667,N_4027,N_4880);
or U6668 (N_6668,N_4495,N_4865);
nand U6669 (N_6669,N_4429,N_4146);
nor U6670 (N_6670,N_4569,N_5934);
nor U6671 (N_6671,N_4647,N_5465);
nor U6672 (N_6672,N_5092,N_5060);
and U6673 (N_6673,N_4051,N_4130);
or U6674 (N_6674,N_4471,N_5316);
and U6675 (N_6675,N_5560,N_4806);
and U6676 (N_6676,N_5974,N_4754);
nand U6677 (N_6677,N_5793,N_4690);
nand U6678 (N_6678,N_4308,N_4847);
nor U6679 (N_6679,N_5565,N_4761);
and U6680 (N_6680,N_4209,N_5681);
nor U6681 (N_6681,N_5443,N_5774);
nor U6682 (N_6682,N_4054,N_5678);
nor U6683 (N_6683,N_5713,N_4323);
and U6684 (N_6684,N_5006,N_5239);
and U6685 (N_6685,N_4781,N_4965);
and U6686 (N_6686,N_5759,N_4890);
or U6687 (N_6687,N_5885,N_5397);
nor U6688 (N_6688,N_4929,N_4503);
nor U6689 (N_6689,N_5519,N_4557);
xor U6690 (N_6690,N_4236,N_5389);
nor U6691 (N_6691,N_5940,N_4660);
nand U6692 (N_6692,N_4529,N_4277);
or U6693 (N_6693,N_5985,N_4252);
and U6694 (N_6694,N_5781,N_4972);
nor U6695 (N_6695,N_5947,N_4326);
and U6696 (N_6696,N_5834,N_4807);
nor U6697 (N_6697,N_4172,N_4675);
and U6698 (N_6698,N_4306,N_5503);
nand U6699 (N_6699,N_4279,N_5049);
nand U6700 (N_6700,N_4513,N_4128);
xor U6701 (N_6701,N_4566,N_5396);
nand U6702 (N_6702,N_5433,N_4996);
and U6703 (N_6703,N_5695,N_5867);
and U6704 (N_6704,N_4794,N_5661);
and U6705 (N_6705,N_5233,N_5038);
and U6706 (N_6706,N_5350,N_4168);
nor U6707 (N_6707,N_4007,N_5386);
nor U6708 (N_6708,N_4212,N_5999);
or U6709 (N_6709,N_5843,N_5575);
nand U6710 (N_6710,N_5341,N_5197);
or U6711 (N_6711,N_5311,N_5182);
xor U6712 (N_6712,N_5285,N_5663);
nor U6713 (N_6713,N_5094,N_5021);
and U6714 (N_6714,N_4656,N_4501);
or U6715 (N_6715,N_5152,N_5096);
nor U6716 (N_6716,N_5772,N_5439);
and U6717 (N_6717,N_5100,N_4452);
nand U6718 (N_6718,N_5598,N_4985);
nor U6719 (N_6719,N_5827,N_4423);
nor U6720 (N_6720,N_4343,N_4713);
nor U6721 (N_6721,N_4837,N_4590);
and U6722 (N_6722,N_5434,N_4402);
nand U6723 (N_6723,N_4914,N_5016);
and U6724 (N_6724,N_4233,N_4502);
or U6725 (N_6725,N_5376,N_5953);
or U6726 (N_6726,N_4992,N_5590);
nor U6727 (N_6727,N_5795,N_4428);
and U6728 (N_6728,N_4065,N_4912);
and U6729 (N_6729,N_5462,N_4247);
nand U6730 (N_6730,N_4885,N_5214);
or U6731 (N_6731,N_5582,N_5487);
nor U6732 (N_6732,N_5930,N_5792);
and U6733 (N_6733,N_4904,N_4844);
or U6734 (N_6734,N_5609,N_4366);
nor U6735 (N_6735,N_5809,N_4842);
xor U6736 (N_6736,N_4090,N_5370);
or U6737 (N_6737,N_4891,N_5165);
nand U6738 (N_6738,N_5818,N_4097);
nor U6739 (N_6739,N_5231,N_4551);
nor U6740 (N_6740,N_4256,N_4762);
nor U6741 (N_6741,N_5426,N_4371);
and U6742 (N_6742,N_4864,N_4845);
or U6743 (N_6743,N_5997,N_4716);
or U6744 (N_6744,N_5543,N_4480);
nor U6745 (N_6745,N_4271,N_4572);
nor U6746 (N_6746,N_4044,N_5673);
nor U6747 (N_6747,N_4124,N_5871);
and U6748 (N_6748,N_5605,N_4190);
or U6749 (N_6749,N_4943,N_4208);
nand U6750 (N_6750,N_5821,N_4550);
nor U6751 (N_6751,N_5430,N_5829);
nand U6752 (N_6752,N_5454,N_5367);
nand U6753 (N_6753,N_5334,N_5393);
nor U6754 (N_6754,N_4311,N_4839);
xor U6755 (N_6755,N_5946,N_5042);
xor U6756 (N_6756,N_5980,N_5053);
or U6757 (N_6757,N_5069,N_4356);
xnor U6758 (N_6758,N_5629,N_5212);
and U6759 (N_6759,N_5418,N_5174);
nor U6760 (N_6760,N_5858,N_5175);
nand U6761 (N_6761,N_4440,N_5074);
or U6762 (N_6762,N_4765,N_4788);
nor U6763 (N_6763,N_4900,N_5656);
xnor U6764 (N_6764,N_4384,N_4793);
nor U6765 (N_6765,N_5297,N_5026);
and U6766 (N_6766,N_4956,N_4881);
nand U6767 (N_6767,N_4248,N_4798);
nand U6768 (N_6768,N_5591,N_4731);
and U6769 (N_6769,N_5399,N_5336);
nand U6770 (N_6770,N_5891,N_5839);
nand U6771 (N_6771,N_4016,N_4293);
nor U6772 (N_6772,N_5764,N_5171);
nor U6773 (N_6773,N_4400,N_4604);
nor U6774 (N_6774,N_4746,N_5036);
nand U6775 (N_6775,N_5445,N_4150);
nor U6776 (N_6776,N_5913,N_4768);
and U6777 (N_6777,N_5987,N_4116);
xor U6778 (N_6778,N_4376,N_4156);
and U6779 (N_6779,N_5584,N_4804);
or U6780 (N_6780,N_4565,N_4539);
or U6781 (N_6781,N_4498,N_4683);
xor U6782 (N_6782,N_5327,N_4789);
nor U6783 (N_6783,N_5102,N_5463);
or U6784 (N_6784,N_4971,N_4050);
or U6785 (N_6785,N_5162,N_4915);
nor U6786 (N_6786,N_4289,N_5634);
and U6787 (N_6787,N_4819,N_4092);
xnor U6788 (N_6788,N_5909,N_5501);
and U6789 (N_6789,N_4341,N_5991);
or U6790 (N_6790,N_4286,N_4391);
nor U6791 (N_6791,N_5528,N_5646);
nand U6792 (N_6792,N_5544,N_4282);
or U6793 (N_6793,N_4582,N_5115);
nand U6794 (N_6794,N_4427,N_4466);
nand U6795 (N_6795,N_5791,N_5970);
nand U6796 (N_6796,N_4826,N_5339);
nand U6797 (N_6797,N_4283,N_5606);
or U6798 (N_6798,N_5183,N_5122);
nand U6799 (N_6799,N_5153,N_5065);
xnor U6800 (N_6800,N_5326,N_5141);
nand U6801 (N_6801,N_4367,N_4045);
and U6802 (N_6802,N_5944,N_5126);
nor U6803 (N_6803,N_5276,N_4063);
and U6804 (N_6804,N_5735,N_5760);
nand U6805 (N_6805,N_5902,N_5417);
nand U6806 (N_6806,N_4449,N_4200);
or U6807 (N_6807,N_5221,N_4294);
and U6808 (N_6808,N_5145,N_5310);
or U6809 (N_6809,N_4562,N_4287);
and U6810 (N_6810,N_5736,N_5597);
and U6811 (N_6811,N_5570,N_5779);
or U6812 (N_6812,N_5048,N_4613);
xor U6813 (N_6813,N_4100,N_4711);
and U6814 (N_6814,N_5872,N_4947);
nor U6815 (N_6815,N_5912,N_4772);
or U6816 (N_6816,N_5107,N_5229);
and U6817 (N_6817,N_5906,N_5039);
nand U6818 (N_6818,N_4148,N_5388);
and U6819 (N_6819,N_5690,N_4976);
or U6820 (N_6820,N_5028,N_4231);
and U6821 (N_6821,N_4988,N_4385);
or U6822 (N_6822,N_5801,N_5306);
or U6823 (N_6823,N_4875,N_5976);
or U6824 (N_6824,N_4443,N_5937);
nor U6825 (N_6825,N_4514,N_5860);
nand U6826 (N_6826,N_4345,N_4263);
and U6827 (N_6827,N_4496,N_4149);
xor U6828 (N_6828,N_5471,N_4451);
or U6829 (N_6829,N_5530,N_4113);
nor U6830 (N_6830,N_4712,N_4685);
and U6831 (N_6831,N_5517,N_4491);
and U6832 (N_6832,N_5623,N_4509);
or U6833 (N_6833,N_5295,N_4439);
nor U6834 (N_6834,N_4668,N_5855);
nand U6835 (N_6835,N_5148,N_5956);
xor U6836 (N_6836,N_4479,N_4933);
nand U6837 (N_6837,N_5506,N_5904);
and U6838 (N_6838,N_4170,N_5954);
or U6839 (N_6839,N_4729,N_4215);
or U6840 (N_6840,N_4857,N_5236);
nor U6841 (N_6841,N_4313,N_5857);
and U6842 (N_6842,N_4722,N_5271);
and U6843 (N_6843,N_4684,N_4907);
or U6844 (N_6844,N_4032,N_4846);
and U6845 (N_6845,N_5526,N_5513);
and U6846 (N_6846,N_4984,N_4605);
nor U6847 (N_6847,N_5101,N_5742);
nor U6848 (N_6848,N_4902,N_5601);
nor U6849 (N_6849,N_4448,N_5404);
nor U6850 (N_6850,N_5186,N_4706);
nor U6851 (N_6851,N_5056,N_4249);
nor U6852 (N_6852,N_5726,N_5614);
nand U6853 (N_6853,N_5088,N_4189);
or U6854 (N_6854,N_5075,N_4899);
nor U6855 (N_6855,N_5636,N_5979);
nor U6856 (N_6856,N_4161,N_5706);
or U6857 (N_6857,N_4580,N_5047);
or U6858 (N_6858,N_4841,N_5533);
and U6859 (N_6859,N_5234,N_5008);
nor U6860 (N_6860,N_5030,N_5758);
nor U6861 (N_6861,N_5332,N_4131);
and U6862 (N_6862,N_4486,N_5593);
nor U6863 (N_6863,N_4721,N_4633);
xnor U6864 (N_6864,N_5640,N_5873);
and U6865 (N_6865,N_5754,N_4099);
and U6866 (N_6866,N_5274,N_4564);
or U6867 (N_6867,N_5072,N_5611);
and U6868 (N_6868,N_4290,N_5846);
nand U6869 (N_6869,N_5160,N_5302);
and U6870 (N_6870,N_4062,N_5237);
nor U6871 (N_6871,N_5670,N_4623);
nor U6872 (N_6872,N_4053,N_5352);
or U6873 (N_6873,N_5990,N_5226);
or U6874 (N_6874,N_4330,N_5689);
and U6875 (N_6875,N_4699,N_4991);
nor U6876 (N_6876,N_4469,N_5887);
nor U6877 (N_6877,N_5010,N_5457);
nand U6878 (N_6878,N_5796,N_5289);
nor U6879 (N_6879,N_5572,N_4349);
or U6880 (N_6880,N_5260,N_5459);
nand U6881 (N_6881,N_5869,N_5093);
nand U6882 (N_6882,N_5029,N_4157);
or U6883 (N_6883,N_4169,N_5224);
xnor U6884 (N_6884,N_5769,N_5704);
nand U6885 (N_6885,N_5973,N_4646);
or U6886 (N_6886,N_5574,N_4254);
nand U6887 (N_6887,N_4747,N_5701);
nor U6888 (N_6888,N_5146,N_5959);
and U6889 (N_6889,N_4077,N_4836);
nand U6890 (N_6890,N_4038,N_5254);
and U6891 (N_6891,N_5412,N_5878);
nand U6892 (N_6892,N_5595,N_4363);
and U6893 (N_6893,N_4764,N_5466);
or U6894 (N_6894,N_4094,N_5814);
or U6895 (N_6895,N_5828,N_5492);
nand U6896 (N_6896,N_4321,N_5798);
nand U6897 (N_6897,N_4422,N_4681);
nand U6898 (N_6898,N_4808,N_5365);
nor U6899 (N_6899,N_4072,N_5960);
xnor U6900 (N_6900,N_5810,N_5283);
nand U6901 (N_6901,N_4137,N_5456);
or U6902 (N_6902,N_4213,N_4518);
and U6903 (N_6903,N_5520,N_4852);
nand U6904 (N_6904,N_4710,N_4389);
and U6905 (N_6905,N_5473,N_4327);
xnor U6906 (N_6906,N_4477,N_4183);
and U6907 (N_6907,N_4010,N_4284);
and U6908 (N_6908,N_5477,N_5658);
nand U6909 (N_6909,N_5151,N_5933);
nor U6910 (N_6910,N_4232,N_4226);
and U6911 (N_6911,N_5468,N_5608);
nor U6912 (N_6912,N_5573,N_4751);
nor U6913 (N_6913,N_4224,N_5111);
nor U6914 (N_6914,N_4797,N_4530);
or U6915 (N_6915,N_4896,N_4624);
nor U6916 (N_6916,N_5391,N_4825);
and U6917 (N_6917,N_4377,N_5738);
or U6918 (N_6918,N_5907,N_4726);
and U6919 (N_6919,N_5447,N_5725);
and U6920 (N_6920,N_5508,N_5240);
nand U6921 (N_6921,N_5286,N_5677);
or U6922 (N_6922,N_5415,N_4221);
or U6923 (N_6923,N_5209,N_4392);
xnor U6924 (N_6924,N_4461,N_4669);
and U6925 (N_6925,N_5645,N_5880);
and U6926 (N_6926,N_4587,N_5566);
and U6927 (N_6927,N_4237,N_5272);
nor U6928 (N_6928,N_5476,N_5464);
or U6929 (N_6929,N_4037,N_4409);
nand U6930 (N_6930,N_5966,N_4420);
nand U6931 (N_6931,N_5641,N_4101);
and U6932 (N_6932,N_4527,N_4296);
nor U6933 (N_6933,N_5583,N_5571);
nor U6934 (N_6934,N_5488,N_5511);
nor U6935 (N_6935,N_4463,N_4003);
nand U6936 (N_6936,N_4796,N_4111);
and U6937 (N_6937,N_4115,N_4199);
nor U6938 (N_6938,N_4584,N_5799);
nor U6939 (N_6939,N_4636,N_5698);
xor U6940 (N_6940,N_4177,N_4578);
xor U6941 (N_6941,N_5340,N_4779);
or U6942 (N_6942,N_4173,N_5863);
xnor U6943 (N_6943,N_4025,N_4187);
nand U6944 (N_6944,N_4952,N_5137);
and U6945 (N_6945,N_5807,N_5652);
nor U6946 (N_6946,N_4339,N_5312);
nand U6947 (N_6947,N_5599,N_4931);
nand U6948 (N_6948,N_4266,N_4589);
and U6949 (N_6949,N_5377,N_5816);
nand U6950 (N_6950,N_5369,N_4974);
nor U6951 (N_6951,N_5780,N_4850);
nand U6952 (N_6952,N_5527,N_4939);
xor U6953 (N_6953,N_4591,N_5842);
xor U6954 (N_6954,N_5659,N_5281);
nor U6955 (N_6955,N_5951,N_5083);
nand U6956 (N_6956,N_4827,N_4821);
nor U6957 (N_6957,N_5886,N_4649);
xnor U6958 (N_6958,N_5246,N_5737);
and U6959 (N_6959,N_5753,N_4510);
nand U6960 (N_6960,N_5632,N_5558);
or U6961 (N_6961,N_5864,N_4147);
nor U6962 (N_6962,N_5989,N_5502);
xor U6963 (N_6963,N_4973,N_4920);
or U6964 (N_6964,N_5408,N_5924);
and U6965 (N_6965,N_5277,N_5351);
xor U6966 (N_6966,N_5515,N_4198);
nor U6967 (N_6967,N_4528,N_4370);
or U6968 (N_6968,N_4948,N_4019);
nor U6969 (N_6969,N_5360,N_4693);
and U6970 (N_6970,N_4637,N_4135);
nor U6971 (N_6971,N_4049,N_4640);
or U6972 (N_6972,N_4817,N_4333);
nand U6973 (N_6973,N_5480,N_4411);
nand U6974 (N_6974,N_4197,N_5196);
or U6975 (N_6975,N_4216,N_4188);
nor U6976 (N_6976,N_5961,N_4760);
and U6977 (N_6977,N_5823,N_4302);
and U6978 (N_6978,N_5046,N_4883);
and U6979 (N_6979,N_4280,N_5730);
xor U6980 (N_6980,N_5660,N_5007);
nor U6981 (N_6981,N_5263,N_5643);
and U6982 (N_6982,N_5952,N_5364);
or U6983 (N_6983,N_4676,N_5452);
xnor U6984 (N_6984,N_4957,N_5716);
and U6985 (N_6985,N_4599,N_4265);
and U6986 (N_6986,N_4814,N_5776);
or U6987 (N_6987,N_5252,N_4143);
or U6988 (N_6988,N_5714,N_4753);
and U6989 (N_6989,N_4082,N_4679);
xor U6990 (N_6990,N_4068,N_5684);
nor U6991 (N_6991,N_5610,N_5125);
xnor U6992 (N_6992,N_5299,N_4140);
or U6993 (N_6993,N_4861,N_5651);
nor U6994 (N_6994,N_5650,N_5161);
nor U6995 (N_6995,N_5534,N_5654);
or U6996 (N_6996,N_5275,N_4986);
nor U6997 (N_6997,N_5993,N_5329);
nor U6998 (N_6998,N_4372,N_5045);
nand U6999 (N_6999,N_4538,N_5413);
nor U7000 (N_7000,N_4267,N_4319);
nor U7001 (N_7001,N_4546,N_4706);
or U7002 (N_7002,N_5907,N_4887);
or U7003 (N_7003,N_4205,N_5782);
or U7004 (N_7004,N_5998,N_5825);
and U7005 (N_7005,N_4804,N_5188);
nor U7006 (N_7006,N_4993,N_5539);
and U7007 (N_7007,N_5982,N_5892);
nand U7008 (N_7008,N_4278,N_5409);
nand U7009 (N_7009,N_4682,N_5392);
xnor U7010 (N_7010,N_5241,N_4963);
nand U7011 (N_7011,N_4226,N_5192);
or U7012 (N_7012,N_5208,N_4695);
or U7013 (N_7013,N_4142,N_4693);
or U7014 (N_7014,N_5080,N_5267);
or U7015 (N_7015,N_4939,N_5972);
and U7016 (N_7016,N_5277,N_4189);
or U7017 (N_7017,N_4571,N_5151);
nand U7018 (N_7018,N_4450,N_5150);
and U7019 (N_7019,N_4709,N_5760);
and U7020 (N_7020,N_4049,N_4898);
nor U7021 (N_7021,N_5330,N_5174);
nand U7022 (N_7022,N_5255,N_4428);
nor U7023 (N_7023,N_5408,N_4366);
and U7024 (N_7024,N_5715,N_5240);
and U7025 (N_7025,N_4306,N_4585);
or U7026 (N_7026,N_4210,N_4929);
nand U7027 (N_7027,N_4063,N_4732);
nor U7028 (N_7028,N_5889,N_5565);
nor U7029 (N_7029,N_5947,N_4395);
and U7030 (N_7030,N_5071,N_5937);
and U7031 (N_7031,N_5738,N_5929);
and U7032 (N_7032,N_4013,N_4400);
nand U7033 (N_7033,N_4348,N_4848);
xor U7034 (N_7034,N_5227,N_5289);
nand U7035 (N_7035,N_4245,N_5164);
xor U7036 (N_7036,N_5356,N_5749);
nand U7037 (N_7037,N_4806,N_4263);
and U7038 (N_7038,N_5387,N_4741);
and U7039 (N_7039,N_4560,N_5233);
nand U7040 (N_7040,N_4836,N_5941);
nand U7041 (N_7041,N_4522,N_5301);
or U7042 (N_7042,N_4513,N_4721);
and U7043 (N_7043,N_4468,N_4517);
or U7044 (N_7044,N_5336,N_4433);
nand U7045 (N_7045,N_4166,N_5458);
and U7046 (N_7046,N_4800,N_5815);
or U7047 (N_7047,N_5423,N_5361);
xnor U7048 (N_7048,N_5451,N_5687);
or U7049 (N_7049,N_4915,N_4102);
or U7050 (N_7050,N_5495,N_4408);
nand U7051 (N_7051,N_4797,N_5324);
or U7052 (N_7052,N_5831,N_5405);
and U7053 (N_7053,N_4383,N_5072);
nor U7054 (N_7054,N_5403,N_4545);
and U7055 (N_7055,N_5155,N_4355);
or U7056 (N_7056,N_5996,N_4934);
or U7057 (N_7057,N_4473,N_4006);
nand U7058 (N_7058,N_4320,N_5084);
nor U7059 (N_7059,N_4719,N_4301);
or U7060 (N_7060,N_4420,N_5071);
and U7061 (N_7061,N_5154,N_4581);
xor U7062 (N_7062,N_5506,N_5708);
nand U7063 (N_7063,N_4189,N_5300);
nand U7064 (N_7064,N_5238,N_4017);
xor U7065 (N_7065,N_4097,N_4341);
and U7066 (N_7066,N_4427,N_4311);
nor U7067 (N_7067,N_4393,N_4861);
and U7068 (N_7068,N_4446,N_5846);
xor U7069 (N_7069,N_4288,N_5597);
and U7070 (N_7070,N_4951,N_4536);
and U7071 (N_7071,N_4940,N_4200);
nor U7072 (N_7072,N_5209,N_4175);
or U7073 (N_7073,N_4726,N_4428);
nor U7074 (N_7074,N_4662,N_5309);
nor U7075 (N_7075,N_5512,N_5744);
nor U7076 (N_7076,N_5091,N_5896);
nand U7077 (N_7077,N_5460,N_5562);
and U7078 (N_7078,N_5236,N_5720);
xnor U7079 (N_7079,N_4375,N_4388);
nor U7080 (N_7080,N_5751,N_4468);
nor U7081 (N_7081,N_5795,N_4091);
or U7082 (N_7082,N_4179,N_4918);
nor U7083 (N_7083,N_5023,N_4603);
nand U7084 (N_7084,N_5847,N_4821);
nor U7085 (N_7085,N_4932,N_5458);
nand U7086 (N_7086,N_5963,N_5110);
or U7087 (N_7087,N_5663,N_5872);
or U7088 (N_7088,N_5088,N_5634);
xnor U7089 (N_7089,N_4213,N_5931);
or U7090 (N_7090,N_5676,N_4636);
or U7091 (N_7091,N_4180,N_5821);
or U7092 (N_7092,N_4929,N_5810);
or U7093 (N_7093,N_5321,N_5305);
nor U7094 (N_7094,N_5864,N_5928);
or U7095 (N_7095,N_4332,N_5925);
or U7096 (N_7096,N_4879,N_4697);
or U7097 (N_7097,N_4314,N_4344);
and U7098 (N_7098,N_5847,N_4069);
xor U7099 (N_7099,N_4909,N_4408);
nor U7100 (N_7100,N_4025,N_5140);
or U7101 (N_7101,N_5465,N_4262);
and U7102 (N_7102,N_4766,N_4537);
and U7103 (N_7103,N_4414,N_4746);
nor U7104 (N_7104,N_5795,N_5223);
nand U7105 (N_7105,N_5702,N_5418);
nor U7106 (N_7106,N_5256,N_4076);
nor U7107 (N_7107,N_5977,N_4883);
and U7108 (N_7108,N_4138,N_4741);
and U7109 (N_7109,N_5700,N_4074);
nand U7110 (N_7110,N_4179,N_5513);
nand U7111 (N_7111,N_5591,N_4441);
and U7112 (N_7112,N_4942,N_5180);
nand U7113 (N_7113,N_4439,N_4682);
or U7114 (N_7114,N_4646,N_5187);
and U7115 (N_7115,N_5999,N_4997);
or U7116 (N_7116,N_4583,N_4616);
and U7117 (N_7117,N_5810,N_4403);
or U7118 (N_7118,N_5022,N_5267);
or U7119 (N_7119,N_4489,N_4547);
nor U7120 (N_7120,N_5744,N_5979);
or U7121 (N_7121,N_5729,N_4574);
nor U7122 (N_7122,N_4493,N_5697);
and U7123 (N_7123,N_4691,N_5405);
nor U7124 (N_7124,N_4536,N_4189);
nand U7125 (N_7125,N_5658,N_5317);
or U7126 (N_7126,N_5681,N_5057);
nor U7127 (N_7127,N_4723,N_5352);
nor U7128 (N_7128,N_5646,N_4293);
nor U7129 (N_7129,N_5352,N_5339);
or U7130 (N_7130,N_5412,N_5259);
nand U7131 (N_7131,N_5475,N_4403);
nor U7132 (N_7132,N_4836,N_4809);
nor U7133 (N_7133,N_5167,N_5049);
xor U7134 (N_7134,N_4203,N_4621);
xnor U7135 (N_7135,N_4899,N_4170);
nor U7136 (N_7136,N_4620,N_4263);
or U7137 (N_7137,N_4810,N_4872);
and U7138 (N_7138,N_5551,N_5291);
or U7139 (N_7139,N_5952,N_5037);
nand U7140 (N_7140,N_4878,N_4825);
and U7141 (N_7141,N_5393,N_4755);
nor U7142 (N_7142,N_4256,N_4189);
xnor U7143 (N_7143,N_4883,N_5028);
or U7144 (N_7144,N_4307,N_5096);
or U7145 (N_7145,N_5006,N_5181);
xnor U7146 (N_7146,N_5624,N_5236);
xor U7147 (N_7147,N_4538,N_5221);
and U7148 (N_7148,N_4139,N_5424);
and U7149 (N_7149,N_4564,N_4272);
nor U7150 (N_7150,N_4095,N_5326);
or U7151 (N_7151,N_5029,N_5965);
and U7152 (N_7152,N_4047,N_5888);
nand U7153 (N_7153,N_4087,N_4931);
nand U7154 (N_7154,N_5458,N_4673);
nand U7155 (N_7155,N_4162,N_4543);
and U7156 (N_7156,N_5344,N_5227);
or U7157 (N_7157,N_4741,N_4988);
and U7158 (N_7158,N_5453,N_5961);
or U7159 (N_7159,N_5043,N_4201);
nor U7160 (N_7160,N_4011,N_5917);
or U7161 (N_7161,N_4367,N_5134);
and U7162 (N_7162,N_4531,N_5646);
nand U7163 (N_7163,N_5470,N_4150);
nand U7164 (N_7164,N_5316,N_5756);
nand U7165 (N_7165,N_4573,N_5314);
and U7166 (N_7166,N_4796,N_4241);
or U7167 (N_7167,N_5240,N_4320);
or U7168 (N_7168,N_4413,N_4471);
xnor U7169 (N_7169,N_4047,N_5844);
nor U7170 (N_7170,N_5419,N_4634);
and U7171 (N_7171,N_5385,N_5798);
nand U7172 (N_7172,N_4105,N_4089);
or U7173 (N_7173,N_4207,N_4041);
or U7174 (N_7174,N_5900,N_5442);
or U7175 (N_7175,N_4748,N_4884);
or U7176 (N_7176,N_5209,N_4601);
or U7177 (N_7177,N_4872,N_5633);
nand U7178 (N_7178,N_4387,N_4842);
nand U7179 (N_7179,N_5812,N_4173);
or U7180 (N_7180,N_5716,N_4768);
nand U7181 (N_7181,N_4747,N_4215);
nor U7182 (N_7182,N_4795,N_5110);
nor U7183 (N_7183,N_4667,N_4499);
nand U7184 (N_7184,N_4223,N_4383);
or U7185 (N_7185,N_5518,N_4472);
nor U7186 (N_7186,N_5783,N_4479);
or U7187 (N_7187,N_5599,N_5410);
and U7188 (N_7188,N_4557,N_5874);
or U7189 (N_7189,N_4906,N_4559);
or U7190 (N_7190,N_4495,N_4695);
nand U7191 (N_7191,N_5320,N_5398);
nand U7192 (N_7192,N_4909,N_5120);
and U7193 (N_7193,N_4928,N_5268);
or U7194 (N_7194,N_4649,N_5088);
nand U7195 (N_7195,N_4488,N_5625);
or U7196 (N_7196,N_4092,N_4016);
and U7197 (N_7197,N_5467,N_4271);
nand U7198 (N_7198,N_4714,N_4329);
nor U7199 (N_7199,N_5377,N_4527);
nand U7200 (N_7200,N_5898,N_5009);
and U7201 (N_7201,N_4770,N_5008);
xnor U7202 (N_7202,N_5249,N_4985);
and U7203 (N_7203,N_4409,N_4904);
xor U7204 (N_7204,N_5244,N_4883);
nand U7205 (N_7205,N_5486,N_4920);
nor U7206 (N_7206,N_5479,N_4847);
nand U7207 (N_7207,N_5621,N_4744);
nor U7208 (N_7208,N_5441,N_4975);
nand U7209 (N_7209,N_4219,N_4757);
or U7210 (N_7210,N_5076,N_4676);
or U7211 (N_7211,N_4964,N_4018);
nand U7212 (N_7212,N_5495,N_4371);
or U7213 (N_7213,N_4172,N_4442);
or U7214 (N_7214,N_4349,N_4008);
and U7215 (N_7215,N_4157,N_4718);
nor U7216 (N_7216,N_5431,N_5785);
nand U7217 (N_7217,N_4540,N_5570);
nand U7218 (N_7218,N_4634,N_4875);
and U7219 (N_7219,N_5621,N_4010);
and U7220 (N_7220,N_5824,N_4477);
and U7221 (N_7221,N_4192,N_4671);
nor U7222 (N_7222,N_4175,N_4679);
or U7223 (N_7223,N_4377,N_5397);
nor U7224 (N_7224,N_5707,N_5089);
or U7225 (N_7225,N_5482,N_4794);
nand U7226 (N_7226,N_5283,N_5930);
nand U7227 (N_7227,N_5850,N_5118);
or U7228 (N_7228,N_5666,N_4522);
and U7229 (N_7229,N_4252,N_5707);
xnor U7230 (N_7230,N_5032,N_5216);
or U7231 (N_7231,N_5122,N_4717);
nor U7232 (N_7232,N_5604,N_4351);
nand U7233 (N_7233,N_4994,N_4634);
and U7234 (N_7234,N_5044,N_4064);
nor U7235 (N_7235,N_5241,N_4813);
nand U7236 (N_7236,N_4688,N_5836);
and U7237 (N_7237,N_5684,N_4673);
nand U7238 (N_7238,N_5243,N_5237);
and U7239 (N_7239,N_5658,N_5379);
nor U7240 (N_7240,N_5439,N_5173);
nand U7241 (N_7241,N_4248,N_4624);
and U7242 (N_7242,N_5253,N_5967);
nand U7243 (N_7243,N_4248,N_5738);
xor U7244 (N_7244,N_4752,N_5386);
and U7245 (N_7245,N_5565,N_4075);
nor U7246 (N_7246,N_5314,N_4097);
or U7247 (N_7247,N_5680,N_5940);
nand U7248 (N_7248,N_5584,N_5706);
and U7249 (N_7249,N_5975,N_5481);
nand U7250 (N_7250,N_5014,N_5687);
xor U7251 (N_7251,N_5264,N_5050);
xnor U7252 (N_7252,N_5053,N_5581);
and U7253 (N_7253,N_5372,N_5737);
xor U7254 (N_7254,N_4759,N_5918);
nor U7255 (N_7255,N_5652,N_4947);
nand U7256 (N_7256,N_5933,N_5315);
or U7257 (N_7257,N_5011,N_4088);
or U7258 (N_7258,N_5388,N_4181);
nand U7259 (N_7259,N_4589,N_5337);
xor U7260 (N_7260,N_5936,N_4381);
and U7261 (N_7261,N_5598,N_5089);
and U7262 (N_7262,N_4314,N_5935);
xnor U7263 (N_7263,N_4498,N_5200);
and U7264 (N_7264,N_4412,N_5359);
and U7265 (N_7265,N_4364,N_4818);
or U7266 (N_7266,N_5173,N_4789);
and U7267 (N_7267,N_5892,N_5516);
nand U7268 (N_7268,N_4996,N_5804);
or U7269 (N_7269,N_4734,N_5460);
and U7270 (N_7270,N_5724,N_4550);
or U7271 (N_7271,N_4563,N_5221);
and U7272 (N_7272,N_4416,N_5900);
or U7273 (N_7273,N_4384,N_5319);
or U7274 (N_7274,N_5441,N_4727);
xor U7275 (N_7275,N_4612,N_5563);
nand U7276 (N_7276,N_5895,N_4831);
xnor U7277 (N_7277,N_4660,N_4950);
nand U7278 (N_7278,N_4401,N_5386);
nor U7279 (N_7279,N_5490,N_5065);
nand U7280 (N_7280,N_4503,N_4572);
nand U7281 (N_7281,N_4529,N_5151);
or U7282 (N_7282,N_5685,N_4241);
and U7283 (N_7283,N_4873,N_4496);
or U7284 (N_7284,N_4435,N_5204);
and U7285 (N_7285,N_5241,N_5912);
or U7286 (N_7286,N_5077,N_5727);
and U7287 (N_7287,N_5010,N_4253);
or U7288 (N_7288,N_5670,N_4114);
nor U7289 (N_7289,N_4191,N_4959);
nor U7290 (N_7290,N_5516,N_4870);
and U7291 (N_7291,N_5549,N_5209);
xnor U7292 (N_7292,N_4903,N_5809);
or U7293 (N_7293,N_4154,N_4562);
nor U7294 (N_7294,N_5641,N_5130);
or U7295 (N_7295,N_5754,N_5369);
or U7296 (N_7296,N_5342,N_5402);
nand U7297 (N_7297,N_4465,N_4135);
or U7298 (N_7298,N_4656,N_4830);
or U7299 (N_7299,N_4248,N_5487);
and U7300 (N_7300,N_5264,N_5535);
nand U7301 (N_7301,N_4428,N_4345);
and U7302 (N_7302,N_4875,N_4580);
and U7303 (N_7303,N_4550,N_5876);
nand U7304 (N_7304,N_5519,N_4297);
xnor U7305 (N_7305,N_4274,N_4191);
and U7306 (N_7306,N_4442,N_4230);
xor U7307 (N_7307,N_4840,N_5776);
nand U7308 (N_7308,N_5690,N_5704);
and U7309 (N_7309,N_5166,N_4666);
or U7310 (N_7310,N_5951,N_4217);
and U7311 (N_7311,N_5069,N_5915);
nor U7312 (N_7312,N_5517,N_4610);
and U7313 (N_7313,N_4266,N_5666);
nor U7314 (N_7314,N_4486,N_5278);
and U7315 (N_7315,N_4740,N_5913);
or U7316 (N_7316,N_4187,N_4091);
or U7317 (N_7317,N_4057,N_5372);
xor U7318 (N_7318,N_5208,N_4713);
and U7319 (N_7319,N_5468,N_5550);
xor U7320 (N_7320,N_4630,N_5422);
nand U7321 (N_7321,N_5914,N_5793);
or U7322 (N_7322,N_5611,N_4763);
nand U7323 (N_7323,N_4801,N_5174);
nor U7324 (N_7324,N_5719,N_4436);
nand U7325 (N_7325,N_4693,N_5994);
nor U7326 (N_7326,N_5797,N_5178);
nand U7327 (N_7327,N_4260,N_5236);
nand U7328 (N_7328,N_4603,N_5777);
and U7329 (N_7329,N_4938,N_4684);
nor U7330 (N_7330,N_4402,N_4971);
or U7331 (N_7331,N_4519,N_4045);
or U7332 (N_7332,N_4625,N_4950);
nand U7333 (N_7333,N_5291,N_5924);
or U7334 (N_7334,N_5568,N_4140);
nor U7335 (N_7335,N_4444,N_4092);
or U7336 (N_7336,N_4707,N_5536);
nand U7337 (N_7337,N_5414,N_5062);
or U7338 (N_7338,N_5956,N_4352);
and U7339 (N_7339,N_5731,N_4052);
or U7340 (N_7340,N_5627,N_4572);
and U7341 (N_7341,N_4210,N_5535);
or U7342 (N_7342,N_4219,N_5681);
and U7343 (N_7343,N_4933,N_4866);
or U7344 (N_7344,N_4727,N_4186);
nor U7345 (N_7345,N_5498,N_4946);
or U7346 (N_7346,N_4601,N_4985);
nand U7347 (N_7347,N_4085,N_4461);
nand U7348 (N_7348,N_5851,N_4457);
nor U7349 (N_7349,N_5773,N_5893);
nand U7350 (N_7350,N_5704,N_5694);
nand U7351 (N_7351,N_5385,N_4819);
nand U7352 (N_7352,N_5955,N_4748);
nand U7353 (N_7353,N_5073,N_4908);
nor U7354 (N_7354,N_5060,N_4071);
nor U7355 (N_7355,N_5491,N_4231);
or U7356 (N_7356,N_5288,N_4763);
nor U7357 (N_7357,N_5626,N_4819);
or U7358 (N_7358,N_4584,N_5678);
or U7359 (N_7359,N_5662,N_5698);
nand U7360 (N_7360,N_5307,N_5739);
nor U7361 (N_7361,N_5633,N_4127);
nor U7362 (N_7362,N_5563,N_4044);
or U7363 (N_7363,N_5542,N_5474);
or U7364 (N_7364,N_4949,N_4908);
or U7365 (N_7365,N_5210,N_4178);
and U7366 (N_7366,N_4701,N_5350);
nand U7367 (N_7367,N_5021,N_5334);
and U7368 (N_7368,N_4427,N_4081);
and U7369 (N_7369,N_5799,N_4859);
nor U7370 (N_7370,N_5909,N_4420);
or U7371 (N_7371,N_5756,N_4881);
or U7372 (N_7372,N_4167,N_4937);
nor U7373 (N_7373,N_4032,N_4099);
xor U7374 (N_7374,N_4775,N_4573);
nor U7375 (N_7375,N_4551,N_5326);
nand U7376 (N_7376,N_5788,N_4408);
or U7377 (N_7377,N_5222,N_5684);
nand U7378 (N_7378,N_5579,N_5216);
xnor U7379 (N_7379,N_5411,N_4020);
nor U7380 (N_7380,N_4048,N_5948);
xnor U7381 (N_7381,N_5379,N_4921);
nand U7382 (N_7382,N_4329,N_5392);
nand U7383 (N_7383,N_5369,N_4571);
xnor U7384 (N_7384,N_4002,N_5917);
nand U7385 (N_7385,N_4482,N_5305);
or U7386 (N_7386,N_5391,N_5670);
nor U7387 (N_7387,N_5335,N_4327);
nand U7388 (N_7388,N_5627,N_5308);
xor U7389 (N_7389,N_4661,N_5793);
nor U7390 (N_7390,N_5608,N_5950);
nor U7391 (N_7391,N_4839,N_4141);
nand U7392 (N_7392,N_5710,N_5270);
and U7393 (N_7393,N_4823,N_5261);
nand U7394 (N_7394,N_4150,N_5140);
nor U7395 (N_7395,N_5267,N_4258);
nor U7396 (N_7396,N_4817,N_4424);
or U7397 (N_7397,N_4238,N_5181);
and U7398 (N_7398,N_5689,N_5680);
and U7399 (N_7399,N_5244,N_5885);
or U7400 (N_7400,N_4705,N_4858);
and U7401 (N_7401,N_4476,N_5388);
xnor U7402 (N_7402,N_5163,N_4381);
or U7403 (N_7403,N_4528,N_5231);
and U7404 (N_7404,N_5591,N_5964);
nand U7405 (N_7405,N_4979,N_4943);
nor U7406 (N_7406,N_4634,N_5007);
nand U7407 (N_7407,N_4515,N_4455);
nor U7408 (N_7408,N_5492,N_4908);
and U7409 (N_7409,N_4842,N_4872);
and U7410 (N_7410,N_4802,N_4176);
or U7411 (N_7411,N_4360,N_4244);
and U7412 (N_7412,N_5328,N_4366);
xnor U7413 (N_7413,N_5582,N_4369);
xnor U7414 (N_7414,N_4047,N_5353);
nand U7415 (N_7415,N_4533,N_4521);
and U7416 (N_7416,N_4024,N_5961);
or U7417 (N_7417,N_5976,N_5281);
and U7418 (N_7418,N_4627,N_4211);
and U7419 (N_7419,N_4972,N_4922);
or U7420 (N_7420,N_4151,N_4059);
and U7421 (N_7421,N_5076,N_4289);
or U7422 (N_7422,N_4109,N_5112);
nor U7423 (N_7423,N_5344,N_4503);
xnor U7424 (N_7424,N_4083,N_5392);
nand U7425 (N_7425,N_5876,N_5941);
and U7426 (N_7426,N_4290,N_5243);
nand U7427 (N_7427,N_5902,N_5169);
nand U7428 (N_7428,N_4365,N_4368);
nand U7429 (N_7429,N_4459,N_4077);
nor U7430 (N_7430,N_5595,N_5242);
nand U7431 (N_7431,N_4886,N_5231);
xor U7432 (N_7432,N_4048,N_5552);
nand U7433 (N_7433,N_4491,N_4189);
nor U7434 (N_7434,N_4823,N_4513);
nor U7435 (N_7435,N_5871,N_5510);
and U7436 (N_7436,N_4529,N_4207);
or U7437 (N_7437,N_4786,N_4281);
or U7438 (N_7438,N_5079,N_5052);
or U7439 (N_7439,N_4281,N_4171);
nor U7440 (N_7440,N_4421,N_4254);
nand U7441 (N_7441,N_4676,N_5475);
xnor U7442 (N_7442,N_5576,N_5443);
nor U7443 (N_7443,N_5379,N_5667);
nor U7444 (N_7444,N_4359,N_4910);
nand U7445 (N_7445,N_5649,N_5056);
and U7446 (N_7446,N_4584,N_5483);
or U7447 (N_7447,N_5475,N_5309);
and U7448 (N_7448,N_4939,N_5698);
nand U7449 (N_7449,N_5518,N_4333);
xnor U7450 (N_7450,N_5940,N_5704);
and U7451 (N_7451,N_5848,N_4187);
or U7452 (N_7452,N_5429,N_5631);
and U7453 (N_7453,N_4233,N_4914);
nand U7454 (N_7454,N_4444,N_5340);
nand U7455 (N_7455,N_4806,N_4915);
or U7456 (N_7456,N_4038,N_4305);
nand U7457 (N_7457,N_4281,N_5085);
and U7458 (N_7458,N_4132,N_4629);
nand U7459 (N_7459,N_5848,N_4794);
nand U7460 (N_7460,N_5500,N_5493);
xor U7461 (N_7461,N_5121,N_4972);
and U7462 (N_7462,N_5352,N_5405);
nand U7463 (N_7463,N_5197,N_5514);
and U7464 (N_7464,N_5155,N_5916);
and U7465 (N_7465,N_4297,N_5097);
or U7466 (N_7466,N_4477,N_4884);
nand U7467 (N_7467,N_4222,N_5225);
or U7468 (N_7468,N_4265,N_4232);
xnor U7469 (N_7469,N_4220,N_5437);
or U7470 (N_7470,N_4848,N_5969);
and U7471 (N_7471,N_5982,N_5661);
nor U7472 (N_7472,N_5491,N_5419);
and U7473 (N_7473,N_5504,N_5224);
nand U7474 (N_7474,N_5362,N_4839);
xnor U7475 (N_7475,N_5489,N_4169);
or U7476 (N_7476,N_4847,N_4618);
xor U7477 (N_7477,N_5506,N_5547);
or U7478 (N_7478,N_4702,N_5426);
nand U7479 (N_7479,N_4864,N_4567);
or U7480 (N_7480,N_5189,N_4878);
and U7481 (N_7481,N_4527,N_5634);
and U7482 (N_7482,N_4082,N_5150);
xor U7483 (N_7483,N_4522,N_4373);
and U7484 (N_7484,N_5877,N_4031);
nand U7485 (N_7485,N_5457,N_4104);
or U7486 (N_7486,N_5218,N_5589);
or U7487 (N_7487,N_5050,N_5103);
and U7488 (N_7488,N_5343,N_5320);
nor U7489 (N_7489,N_5618,N_4860);
nand U7490 (N_7490,N_4209,N_5715);
and U7491 (N_7491,N_5733,N_4689);
nor U7492 (N_7492,N_4811,N_5798);
xor U7493 (N_7493,N_5462,N_5750);
nand U7494 (N_7494,N_5614,N_4430);
nand U7495 (N_7495,N_5311,N_4422);
nand U7496 (N_7496,N_4115,N_5444);
nand U7497 (N_7497,N_5996,N_5128);
or U7498 (N_7498,N_5911,N_5798);
xor U7499 (N_7499,N_4100,N_5475);
nor U7500 (N_7500,N_5794,N_4822);
or U7501 (N_7501,N_5630,N_4755);
and U7502 (N_7502,N_5844,N_4012);
or U7503 (N_7503,N_5964,N_4283);
nor U7504 (N_7504,N_5684,N_5463);
nand U7505 (N_7505,N_4007,N_4218);
nand U7506 (N_7506,N_5433,N_5407);
nand U7507 (N_7507,N_4775,N_4057);
or U7508 (N_7508,N_4300,N_4251);
nand U7509 (N_7509,N_4396,N_5941);
nand U7510 (N_7510,N_4275,N_4460);
nand U7511 (N_7511,N_4064,N_4508);
nand U7512 (N_7512,N_5781,N_5681);
nand U7513 (N_7513,N_5168,N_5067);
and U7514 (N_7514,N_4713,N_4819);
or U7515 (N_7515,N_5079,N_5978);
or U7516 (N_7516,N_4198,N_5084);
and U7517 (N_7517,N_4265,N_5037);
and U7518 (N_7518,N_5800,N_5711);
nand U7519 (N_7519,N_5896,N_4463);
nor U7520 (N_7520,N_5614,N_5909);
and U7521 (N_7521,N_5739,N_4748);
nor U7522 (N_7522,N_5048,N_4937);
and U7523 (N_7523,N_5769,N_4811);
nand U7524 (N_7524,N_4429,N_4073);
nand U7525 (N_7525,N_5463,N_5326);
nand U7526 (N_7526,N_5333,N_5516);
or U7527 (N_7527,N_4142,N_5227);
nor U7528 (N_7528,N_4003,N_4176);
nand U7529 (N_7529,N_4211,N_4143);
xnor U7530 (N_7530,N_5147,N_5749);
or U7531 (N_7531,N_4790,N_4395);
nand U7532 (N_7532,N_4375,N_4343);
or U7533 (N_7533,N_4413,N_5101);
or U7534 (N_7534,N_4235,N_5453);
xor U7535 (N_7535,N_5348,N_4806);
and U7536 (N_7536,N_4485,N_4327);
or U7537 (N_7537,N_4006,N_5063);
or U7538 (N_7538,N_5593,N_5044);
and U7539 (N_7539,N_4555,N_5937);
nand U7540 (N_7540,N_4334,N_5798);
nand U7541 (N_7541,N_4484,N_5688);
nand U7542 (N_7542,N_4784,N_5661);
or U7543 (N_7543,N_4981,N_4911);
nor U7544 (N_7544,N_4868,N_5241);
and U7545 (N_7545,N_5414,N_5107);
nand U7546 (N_7546,N_5521,N_5547);
nor U7547 (N_7547,N_4047,N_5250);
or U7548 (N_7548,N_5854,N_5538);
nand U7549 (N_7549,N_5126,N_5723);
and U7550 (N_7550,N_5117,N_4303);
and U7551 (N_7551,N_4364,N_5267);
nand U7552 (N_7552,N_4185,N_5824);
nor U7553 (N_7553,N_5427,N_5078);
nand U7554 (N_7554,N_4306,N_4805);
or U7555 (N_7555,N_5754,N_4034);
and U7556 (N_7556,N_4907,N_4156);
or U7557 (N_7557,N_4490,N_4683);
nand U7558 (N_7558,N_4639,N_4525);
nor U7559 (N_7559,N_5765,N_4277);
nor U7560 (N_7560,N_4163,N_5074);
xnor U7561 (N_7561,N_4335,N_5737);
and U7562 (N_7562,N_4849,N_5749);
nand U7563 (N_7563,N_4819,N_5261);
or U7564 (N_7564,N_4635,N_5838);
nand U7565 (N_7565,N_5901,N_5817);
nor U7566 (N_7566,N_4776,N_5648);
nor U7567 (N_7567,N_5802,N_4358);
xnor U7568 (N_7568,N_4124,N_4544);
or U7569 (N_7569,N_5839,N_5169);
or U7570 (N_7570,N_5889,N_5324);
nand U7571 (N_7571,N_4096,N_5987);
and U7572 (N_7572,N_5262,N_5347);
nor U7573 (N_7573,N_4848,N_4733);
or U7574 (N_7574,N_5484,N_4475);
nor U7575 (N_7575,N_4711,N_5630);
nor U7576 (N_7576,N_4299,N_5549);
or U7577 (N_7577,N_4040,N_4344);
nand U7578 (N_7578,N_5910,N_4505);
xor U7579 (N_7579,N_5924,N_5152);
or U7580 (N_7580,N_4927,N_5483);
nand U7581 (N_7581,N_4978,N_5328);
or U7582 (N_7582,N_5522,N_4585);
nand U7583 (N_7583,N_4567,N_4145);
and U7584 (N_7584,N_5911,N_5535);
or U7585 (N_7585,N_5948,N_4551);
and U7586 (N_7586,N_4014,N_5485);
xnor U7587 (N_7587,N_5118,N_5121);
xnor U7588 (N_7588,N_4399,N_4814);
or U7589 (N_7589,N_5751,N_5333);
or U7590 (N_7590,N_5487,N_4919);
and U7591 (N_7591,N_5345,N_4434);
nand U7592 (N_7592,N_4877,N_5894);
or U7593 (N_7593,N_4362,N_5022);
or U7594 (N_7594,N_5661,N_5777);
and U7595 (N_7595,N_5907,N_5839);
nand U7596 (N_7596,N_4734,N_5420);
and U7597 (N_7597,N_4238,N_4268);
or U7598 (N_7598,N_5138,N_4435);
and U7599 (N_7599,N_4965,N_4660);
and U7600 (N_7600,N_5390,N_4369);
and U7601 (N_7601,N_4947,N_5374);
nor U7602 (N_7602,N_5040,N_4528);
and U7603 (N_7603,N_4690,N_4573);
or U7604 (N_7604,N_4513,N_4285);
xnor U7605 (N_7605,N_5165,N_5070);
nand U7606 (N_7606,N_4743,N_5993);
and U7607 (N_7607,N_5834,N_4283);
and U7608 (N_7608,N_5342,N_5910);
nand U7609 (N_7609,N_5543,N_5320);
and U7610 (N_7610,N_4685,N_5901);
nor U7611 (N_7611,N_5464,N_5650);
nor U7612 (N_7612,N_5387,N_5051);
and U7613 (N_7613,N_4746,N_5628);
nor U7614 (N_7614,N_5211,N_4188);
and U7615 (N_7615,N_4822,N_4952);
and U7616 (N_7616,N_4296,N_5592);
or U7617 (N_7617,N_5962,N_4830);
or U7618 (N_7618,N_5974,N_5920);
or U7619 (N_7619,N_4442,N_5054);
or U7620 (N_7620,N_4981,N_4791);
nor U7621 (N_7621,N_4220,N_4809);
and U7622 (N_7622,N_4937,N_5255);
nor U7623 (N_7623,N_5746,N_4767);
nand U7624 (N_7624,N_4728,N_5467);
or U7625 (N_7625,N_4419,N_4094);
nor U7626 (N_7626,N_4561,N_4587);
or U7627 (N_7627,N_5383,N_4829);
nand U7628 (N_7628,N_4293,N_5972);
nor U7629 (N_7629,N_4514,N_4770);
or U7630 (N_7630,N_4270,N_4785);
nor U7631 (N_7631,N_5098,N_4176);
nand U7632 (N_7632,N_4330,N_5394);
or U7633 (N_7633,N_4416,N_4761);
nand U7634 (N_7634,N_4795,N_5398);
and U7635 (N_7635,N_4573,N_5127);
and U7636 (N_7636,N_4382,N_4622);
or U7637 (N_7637,N_4621,N_4324);
xor U7638 (N_7638,N_4028,N_4338);
and U7639 (N_7639,N_4804,N_4200);
or U7640 (N_7640,N_5869,N_5992);
and U7641 (N_7641,N_5245,N_4135);
xor U7642 (N_7642,N_5764,N_5988);
nor U7643 (N_7643,N_4200,N_5231);
nand U7644 (N_7644,N_5684,N_5440);
nor U7645 (N_7645,N_4577,N_4918);
nor U7646 (N_7646,N_5365,N_4549);
and U7647 (N_7647,N_4711,N_5979);
nor U7648 (N_7648,N_4806,N_4672);
nor U7649 (N_7649,N_5079,N_4744);
or U7650 (N_7650,N_4100,N_4471);
or U7651 (N_7651,N_5737,N_4863);
and U7652 (N_7652,N_5520,N_5911);
and U7653 (N_7653,N_4030,N_5716);
nor U7654 (N_7654,N_5584,N_4100);
or U7655 (N_7655,N_5320,N_5820);
or U7656 (N_7656,N_4111,N_5059);
xor U7657 (N_7657,N_5784,N_4155);
nand U7658 (N_7658,N_4149,N_4065);
or U7659 (N_7659,N_5364,N_5184);
xnor U7660 (N_7660,N_5326,N_4242);
xor U7661 (N_7661,N_5422,N_5763);
or U7662 (N_7662,N_4249,N_5517);
or U7663 (N_7663,N_5490,N_5685);
or U7664 (N_7664,N_5856,N_5359);
and U7665 (N_7665,N_4950,N_4273);
and U7666 (N_7666,N_4782,N_5344);
and U7667 (N_7667,N_4446,N_5272);
or U7668 (N_7668,N_5556,N_5900);
nor U7669 (N_7669,N_5264,N_4769);
nand U7670 (N_7670,N_4119,N_5265);
and U7671 (N_7671,N_5833,N_4406);
nand U7672 (N_7672,N_4073,N_5061);
and U7673 (N_7673,N_4565,N_5187);
nand U7674 (N_7674,N_4547,N_5964);
or U7675 (N_7675,N_4992,N_4781);
and U7676 (N_7676,N_5777,N_5601);
nor U7677 (N_7677,N_5538,N_5660);
nand U7678 (N_7678,N_4819,N_4135);
xor U7679 (N_7679,N_4615,N_5173);
nor U7680 (N_7680,N_4353,N_4504);
nor U7681 (N_7681,N_5446,N_5427);
and U7682 (N_7682,N_5623,N_4595);
or U7683 (N_7683,N_5241,N_5051);
nand U7684 (N_7684,N_4112,N_5069);
nand U7685 (N_7685,N_5963,N_4107);
and U7686 (N_7686,N_5643,N_4803);
nand U7687 (N_7687,N_4086,N_4473);
and U7688 (N_7688,N_5992,N_5055);
nand U7689 (N_7689,N_4449,N_5805);
nor U7690 (N_7690,N_5317,N_5884);
or U7691 (N_7691,N_5449,N_4732);
nor U7692 (N_7692,N_4348,N_5822);
or U7693 (N_7693,N_5722,N_5859);
nand U7694 (N_7694,N_5191,N_5350);
xor U7695 (N_7695,N_5472,N_4448);
and U7696 (N_7696,N_4112,N_4634);
or U7697 (N_7697,N_5677,N_4139);
nand U7698 (N_7698,N_5204,N_5489);
nor U7699 (N_7699,N_5456,N_5724);
or U7700 (N_7700,N_5976,N_5844);
xnor U7701 (N_7701,N_4804,N_4363);
nand U7702 (N_7702,N_4768,N_4420);
nor U7703 (N_7703,N_5514,N_4451);
and U7704 (N_7704,N_5441,N_5534);
and U7705 (N_7705,N_4913,N_5229);
nand U7706 (N_7706,N_5751,N_4395);
or U7707 (N_7707,N_4328,N_5451);
or U7708 (N_7708,N_5095,N_4750);
nand U7709 (N_7709,N_5845,N_4285);
nand U7710 (N_7710,N_5689,N_5611);
xor U7711 (N_7711,N_5115,N_5366);
and U7712 (N_7712,N_5061,N_5828);
and U7713 (N_7713,N_5416,N_5897);
and U7714 (N_7714,N_5980,N_4830);
or U7715 (N_7715,N_5114,N_4167);
or U7716 (N_7716,N_4256,N_5264);
nor U7717 (N_7717,N_4932,N_5250);
nand U7718 (N_7718,N_5118,N_5475);
nand U7719 (N_7719,N_4023,N_5689);
nor U7720 (N_7720,N_5606,N_5907);
xnor U7721 (N_7721,N_4844,N_5303);
xor U7722 (N_7722,N_5866,N_4277);
and U7723 (N_7723,N_4992,N_5774);
and U7724 (N_7724,N_4554,N_5832);
nor U7725 (N_7725,N_5678,N_4045);
or U7726 (N_7726,N_4236,N_4651);
nand U7727 (N_7727,N_5335,N_5802);
or U7728 (N_7728,N_4052,N_5289);
nand U7729 (N_7729,N_5945,N_5532);
or U7730 (N_7730,N_4843,N_5906);
and U7731 (N_7731,N_5786,N_5997);
or U7732 (N_7732,N_4120,N_5625);
nor U7733 (N_7733,N_5913,N_4876);
or U7734 (N_7734,N_4287,N_5538);
nand U7735 (N_7735,N_4703,N_4533);
and U7736 (N_7736,N_4346,N_4666);
nand U7737 (N_7737,N_5337,N_4603);
nor U7738 (N_7738,N_5263,N_5566);
nand U7739 (N_7739,N_4372,N_4716);
and U7740 (N_7740,N_5426,N_4108);
or U7741 (N_7741,N_5502,N_5723);
nor U7742 (N_7742,N_5819,N_4790);
nor U7743 (N_7743,N_4528,N_5198);
xnor U7744 (N_7744,N_4207,N_4353);
and U7745 (N_7745,N_4212,N_4518);
nand U7746 (N_7746,N_5770,N_5970);
and U7747 (N_7747,N_5252,N_4672);
nand U7748 (N_7748,N_4442,N_4736);
xnor U7749 (N_7749,N_4006,N_4255);
nor U7750 (N_7750,N_5719,N_4456);
or U7751 (N_7751,N_5122,N_4422);
and U7752 (N_7752,N_4684,N_5278);
or U7753 (N_7753,N_5774,N_5554);
and U7754 (N_7754,N_5821,N_4197);
or U7755 (N_7755,N_4756,N_5907);
nand U7756 (N_7756,N_4147,N_5768);
or U7757 (N_7757,N_5408,N_4427);
and U7758 (N_7758,N_4274,N_4965);
nand U7759 (N_7759,N_5444,N_4129);
nand U7760 (N_7760,N_4182,N_5976);
nand U7761 (N_7761,N_5923,N_4406);
nor U7762 (N_7762,N_5525,N_5711);
and U7763 (N_7763,N_5647,N_5555);
nor U7764 (N_7764,N_4272,N_4549);
nand U7765 (N_7765,N_4308,N_4965);
xor U7766 (N_7766,N_5277,N_4848);
nor U7767 (N_7767,N_5215,N_5490);
nand U7768 (N_7768,N_4728,N_4501);
nand U7769 (N_7769,N_4714,N_5673);
nand U7770 (N_7770,N_5702,N_5242);
nor U7771 (N_7771,N_5326,N_4430);
and U7772 (N_7772,N_5317,N_5987);
or U7773 (N_7773,N_5919,N_5803);
or U7774 (N_7774,N_5843,N_5506);
nor U7775 (N_7775,N_5358,N_4745);
nand U7776 (N_7776,N_4566,N_5225);
nor U7777 (N_7777,N_4907,N_5591);
nand U7778 (N_7778,N_5657,N_5921);
nor U7779 (N_7779,N_4874,N_5966);
xnor U7780 (N_7780,N_4530,N_5566);
nor U7781 (N_7781,N_5626,N_4135);
nand U7782 (N_7782,N_5741,N_5229);
nand U7783 (N_7783,N_5484,N_4962);
nor U7784 (N_7784,N_5944,N_5792);
nor U7785 (N_7785,N_5013,N_5449);
xor U7786 (N_7786,N_5989,N_4261);
nor U7787 (N_7787,N_4488,N_5185);
nand U7788 (N_7788,N_5666,N_5770);
and U7789 (N_7789,N_5072,N_5427);
xnor U7790 (N_7790,N_4793,N_4612);
or U7791 (N_7791,N_5715,N_4862);
xor U7792 (N_7792,N_4164,N_4127);
xor U7793 (N_7793,N_4037,N_5932);
nand U7794 (N_7794,N_5862,N_5150);
nand U7795 (N_7795,N_5079,N_5481);
or U7796 (N_7796,N_5846,N_4976);
and U7797 (N_7797,N_4231,N_5818);
nand U7798 (N_7798,N_4621,N_5286);
nand U7799 (N_7799,N_4730,N_5107);
nand U7800 (N_7800,N_4318,N_5697);
nand U7801 (N_7801,N_4925,N_5251);
xor U7802 (N_7802,N_4137,N_4772);
xnor U7803 (N_7803,N_4247,N_5203);
nor U7804 (N_7804,N_4033,N_5854);
nand U7805 (N_7805,N_5342,N_5822);
nand U7806 (N_7806,N_4625,N_5589);
nor U7807 (N_7807,N_5439,N_5144);
nand U7808 (N_7808,N_5158,N_5157);
or U7809 (N_7809,N_5097,N_4501);
or U7810 (N_7810,N_5156,N_5693);
and U7811 (N_7811,N_5310,N_4295);
nor U7812 (N_7812,N_4059,N_5039);
and U7813 (N_7813,N_4241,N_4778);
xnor U7814 (N_7814,N_5965,N_4740);
or U7815 (N_7815,N_4959,N_4645);
xnor U7816 (N_7816,N_5231,N_5942);
nor U7817 (N_7817,N_5786,N_5868);
and U7818 (N_7818,N_5454,N_4816);
and U7819 (N_7819,N_5849,N_4046);
nor U7820 (N_7820,N_5664,N_4853);
nand U7821 (N_7821,N_5532,N_4919);
nor U7822 (N_7822,N_5581,N_4406);
and U7823 (N_7823,N_5578,N_5527);
nor U7824 (N_7824,N_4683,N_5661);
nand U7825 (N_7825,N_5204,N_5415);
and U7826 (N_7826,N_5504,N_4845);
or U7827 (N_7827,N_5644,N_5373);
or U7828 (N_7828,N_5379,N_4118);
nand U7829 (N_7829,N_4905,N_5321);
or U7830 (N_7830,N_5022,N_5281);
or U7831 (N_7831,N_5387,N_4283);
nor U7832 (N_7832,N_5875,N_5424);
or U7833 (N_7833,N_4966,N_4202);
nand U7834 (N_7834,N_5210,N_5050);
or U7835 (N_7835,N_4785,N_4023);
or U7836 (N_7836,N_4866,N_5702);
or U7837 (N_7837,N_5761,N_5894);
xnor U7838 (N_7838,N_4197,N_4851);
and U7839 (N_7839,N_5141,N_5445);
or U7840 (N_7840,N_4249,N_4275);
nor U7841 (N_7841,N_4854,N_5185);
or U7842 (N_7842,N_5385,N_4280);
nand U7843 (N_7843,N_4085,N_4347);
and U7844 (N_7844,N_5672,N_4059);
xnor U7845 (N_7845,N_4210,N_5675);
nor U7846 (N_7846,N_5628,N_5981);
nor U7847 (N_7847,N_4381,N_5654);
and U7848 (N_7848,N_5570,N_5500);
nor U7849 (N_7849,N_4896,N_4830);
or U7850 (N_7850,N_4786,N_4013);
or U7851 (N_7851,N_5740,N_4804);
and U7852 (N_7852,N_4964,N_4835);
nand U7853 (N_7853,N_4663,N_4788);
nor U7854 (N_7854,N_4448,N_4598);
or U7855 (N_7855,N_5231,N_5570);
nor U7856 (N_7856,N_4694,N_5457);
nand U7857 (N_7857,N_5291,N_4691);
nand U7858 (N_7858,N_5255,N_4011);
nor U7859 (N_7859,N_4556,N_4583);
xnor U7860 (N_7860,N_5118,N_5082);
xor U7861 (N_7861,N_4905,N_4460);
and U7862 (N_7862,N_5279,N_4049);
nor U7863 (N_7863,N_4345,N_4584);
and U7864 (N_7864,N_5288,N_4637);
and U7865 (N_7865,N_4091,N_4785);
nand U7866 (N_7866,N_4412,N_5793);
nand U7867 (N_7867,N_5872,N_4976);
and U7868 (N_7868,N_4309,N_5272);
or U7869 (N_7869,N_5385,N_4182);
nor U7870 (N_7870,N_5468,N_4000);
nand U7871 (N_7871,N_4697,N_5358);
and U7872 (N_7872,N_5545,N_5247);
nor U7873 (N_7873,N_4354,N_4207);
nand U7874 (N_7874,N_4678,N_5948);
nor U7875 (N_7875,N_5861,N_4713);
nand U7876 (N_7876,N_5872,N_4896);
or U7877 (N_7877,N_5279,N_4383);
nand U7878 (N_7878,N_5192,N_4381);
nor U7879 (N_7879,N_5105,N_4563);
nor U7880 (N_7880,N_4466,N_4007);
nand U7881 (N_7881,N_4168,N_5283);
or U7882 (N_7882,N_5983,N_5720);
or U7883 (N_7883,N_5637,N_5881);
or U7884 (N_7884,N_5857,N_4131);
nor U7885 (N_7885,N_4251,N_5408);
nor U7886 (N_7886,N_4648,N_5277);
nand U7887 (N_7887,N_5705,N_5941);
or U7888 (N_7888,N_5335,N_4229);
nor U7889 (N_7889,N_4836,N_5070);
nand U7890 (N_7890,N_5253,N_5260);
nand U7891 (N_7891,N_5404,N_4390);
and U7892 (N_7892,N_5477,N_4299);
nor U7893 (N_7893,N_4773,N_5956);
nor U7894 (N_7894,N_4484,N_4547);
or U7895 (N_7895,N_4245,N_5349);
nand U7896 (N_7896,N_5831,N_4233);
nor U7897 (N_7897,N_4308,N_5794);
nand U7898 (N_7898,N_4349,N_5256);
nand U7899 (N_7899,N_5992,N_4792);
and U7900 (N_7900,N_4454,N_4363);
and U7901 (N_7901,N_4619,N_5221);
nor U7902 (N_7902,N_4980,N_5867);
nand U7903 (N_7903,N_5561,N_4124);
xnor U7904 (N_7904,N_5567,N_4453);
or U7905 (N_7905,N_4255,N_5186);
xor U7906 (N_7906,N_4666,N_4188);
or U7907 (N_7907,N_4747,N_5923);
or U7908 (N_7908,N_4395,N_4988);
and U7909 (N_7909,N_4823,N_4069);
or U7910 (N_7910,N_5946,N_4244);
and U7911 (N_7911,N_5792,N_4385);
or U7912 (N_7912,N_4193,N_4392);
xnor U7913 (N_7913,N_5210,N_5545);
nor U7914 (N_7914,N_5453,N_4645);
nand U7915 (N_7915,N_5559,N_5829);
and U7916 (N_7916,N_5583,N_4190);
and U7917 (N_7917,N_4047,N_4290);
or U7918 (N_7918,N_4930,N_4202);
nor U7919 (N_7919,N_5149,N_4949);
nor U7920 (N_7920,N_4239,N_5290);
xnor U7921 (N_7921,N_4153,N_5030);
nor U7922 (N_7922,N_5877,N_5298);
and U7923 (N_7923,N_5522,N_4492);
and U7924 (N_7924,N_4154,N_4443);
and U7925 (N_7925,N_5816,N_5098);
and U7926 (N_7926,N_5917,N_4825);
and U7927 (N_7927,N_4385,N_4614);
and U7928 (N_7928,N_4592,N_4651);
and U7929 (N_7929,N_4171,N_5240);
or U7930 (N_7930,N_5224,N_4418);
nor U7931 (N_7931,N_5143,N_4433);
nand U7932 (N_7932,N_5185,N_5990);
xnor U7933 (N_7933,N_5014,N_4574);
nand U7934 (N_7934,N_5767,N_5668);
and U7935 (N_7935,N_4402,N_4009);
or U7936 (N_7936,N_4681,N_5884);
nor U7937 (N_7937,N_4142,N_4840);
or U7938 (N_7938,N_4229,N_5710);
nor U7939 (N_7939,N_5984,N_5572);
and U7940 (N_7940,N_5020,N_5969);
xor U7941 (N_7941,N_4178,N_4554);
xnor U7942 (N_7942,N_4318,N_4090);
xnor U7943 (N_7943,N_4702,N_4013);
nor U7944 (N_7944,N_4614,N_5704);
nand U7945 (N_7945,N_5184,N_4236);
or U7946 (N_7946,N_4758,N_4070);
nor U7947 (N_7947,N_5773,N_5192);
or U7948 (N_7948,N_5940,N_5097);
and U7949 (N_7949,N_4906,N_5506);
nor U7950 (N_7950,N_5425,N_5600);
nand U7951 (N_7951,N_5022,N_5473);
and U7952 (N_7952,N_4990,N_4794);
or U7953 (N_7953,N_4426,N_5790);
nor U7954 (N_7954,N_5061,N_5871);
nand U7955 (N_7955,N_5250,N_4064);
and U7956 (N_7956,N_4751,N_4357);
nor U7957 (N_7957,N_4649,N_4896);
nand U7958 (N_7958,N_4404,N_5548);
or U7959 (N_7959,N_4093,N_5650);
or U7960 (N_7960,N_4007,N_4533);
xor U7961 (N_7961,N_5011,N_4564);
or U7962 (N_7962,N_5863,N_5445);
nand U7963 (N_7963,N_5021,N_4280);
nor U7964 (N_7964,N_4785,N_4071);
nor U7965 (N_7965,N_4525,N_4932);
xor U7966 (N_7966,N_5979,N_4179);
nor U7967 (N_7967,N_5404,N_4478);
nor U7968 (N_7968,N_5268,N_5922);
nor U7969 (N_7969,N_5615,N_5651);
nor U7970 (N_7970,N_5886,N_5709);
nand U7971 (N_7971,N_4109,N_4332);
nand U7972 (N_7972,N_4161,N_5136);
nand U7973 (N_7973,N_5146,N_4344);
nor U7974 (N_7974,N_4157,N_5126);
nor U7975 (N_7975,N_4546,N_5438);
xnor U7976 (N_7976,N_5606,N_5091);
nor U7977 (N_7977,N_5421,N_4861);
nor U7978 (N_7978,N_5570,N_5071);
nor U7979 (N_7979,N_5424,N_5874);
nor U7980 (N_7980,N_5231,N_5014);
and U7981 (N_7981,N_5869,N_4497);
or U7982 (N_7982,N_5479,N_5308);
xor U7983 (N_7983,N_4678,N_5223);
or U7984 (N_7984,N_5820,N_5489);
or U7985 (N_7985,N_4860,N_5323);
and U7986 (N_7986,N_5837,N_5600);
xnor U7987 (N_7987,N_5316,N_4208);
nor U7988 (N_7988,N_5276,N_5197);
or U7989 (N_7989,N_4186,N_4482);
or U7990 (N_7990,N_4864,N_4225);
xnor U7991 (N_7991,N_5049,N_5960);
nand U7992 (N_7992,N_4032,N_5824);
xnor U7993 (N_7993,N_5663,N_5804);
nor U7994 (N_7994,N_4258,N_4593);
nor U7995 (N_7995,N_5049,N_4409);
nand U7996 (N_7996,N_5616,N_5569);
nor U7997 (N_7997,N_5756,N_4011);
or U7998 (N_7998,N_4892,N_5058);
or U7999 (N_7999,N_4468,N_5326);
or U8000 (N_8000,N_6668,N_7153);
nand U8001 (N_8001,N_6113,N_7550);
or U8002 (N_8002,N_7509,N_6003);
and U8003 (N_8003,N_7312,N_6059);
xor U8004 (N_8004,N_7492,N_6166);
nand U8005 (N_8005,N_7752,N_6007);
nand U8006 (N_8006,N_7464,N_6527);
or U8007 (N_8007,N_6469,N_6689);
and U8008 (N_8008,N_7174,N_7883);
nand U8009 (N_8009,N_7080,N_6897);
nor U8010 (N_8010,N_7846,N_6094);
or U8011 (N_8011,N_6795,N_6684);
or U8012 (N_8012,N_7479,N_7706);
xnor U8013 (N_8013,N_7860,N_6018);
or U8014 (N_8014,N_6393,N_6972);
nand U8015 (N_8015,N_7244,N_6522);
nor U8016 (N_8016,N_7100,N_6847);
and U8017 (N_8017,N_6429,N_6600);
and U8018 (N_8018,N_7903,N_7489);
xor U8019 (N_8019,N_7210,N_7146);
or U8020 (N_8020,N_6692,N_7291);
nand U8021 (N_8021,N_7305,N_6362);
nand U8022 (N_8022,N_7577,N_7920);
nand U8023 (N_8023,N_6125,N_7086);
and U8024 (N_8024,N_6793,N_7680);
or U8025 (N_8025,N_6559,N_7350);
nand U8026 (N_8026,N_7738,N_6501);
and U8027 (N_8027,N_6072,N_6833);
or U8028 (N_8028,N_7670,N_6004);
and U8029 (N_8029,N_6303,N_7557);
or U8030 (N_8030,N_6866,N_7946);
and U8031 (N_8031,N_7500,N_7295);
and U8032 (N_8032,N_7833,N_7837);
or U8033 (N_8033,N_6761,N_6807);
xnor U8034 (N_8034,N_7673,N_7540);
and U8035 (N_8035,N_7396,N_6152);
nand U8036 (N_8036,N_6546,N_6949);
or U8037 (N_8037,N_6767,N_7923);
nor U8038 (N_8038,N_7053,N_6870);
or U8039 (N_8039,N_6970,N_7416);
or U8040 (N_8040,N_7434,N_6090);
or U8041 (N_8041,N_7804,N_6998);
xnor U8042 (N_8042,N_6197,N_7071);
nand U8043 (N_8043,N_7525,N_6411);
or U8044 (N_8044,N_6046,N_6984);
or U8045 (N_8045,N_6109,N_7611);
xor U8046 (N_8046,N_7809,N_7668);
xnor U8047 (N_8047,N_7058,N_7303);
nand U8048 (N_8048,N_7934,N_6587);
or U8049 (N_8049,N_7152,N_7382);
nor U8050 (N_8050,N_6036,N_6466);
and U8051 (N_8051,N_7967,N_6500);
nand U8052 (N_8052,N_7590,N_7366);
nor U8053 (N_8053,N_6121,N_6687);
and U8054 (N_8054,N_7499,N_7377);
nor U8055 (N_8055,N_6718,N_7294);
and U8056 (N_8056,N_6924,N_7609);
and U8057 (N_8057,N_7678,N_6406);
nand U8058 (N_8058,N_7186,N_7085);
nor U8059 (N_8059,N_7290,N_6184);
and U8060 (N_8060,N_7064,N_7635);
nor U8061 (N_8061,N_7496,N_7665);
nand U8062 (N_8062,N_7664,N_7947);
and U8063 (N_8063,N_7299,N_7616);
nor U8064 (N_8064,N_7987,N_7686);
or U8065 (N_8065,N_6209,N_7584);
and U8066 (N_8066,N_6569,N_7183);
or U8067 (N_8067,N_6182,N_6159);
nand U8068 (N_8068,N_6788,N_7040);
and U8069 (N_8069,N_6370,N_7891);
and U8070 (N_8070,N_6991,N_6029);
and U8071 (N_8071,N_7547,N_6048);
and U8072 (N_8072,N_7015,N_6274);
nor U8073 (N_8073,N_7850,N_7483);
or U8074 (N_8074,N_7108,N_7684);
nand U8075 (N_8075,N_7650,N_7930);
or U8076 (N_8076,N_7451,N_6082);
and U8077 (N_8077,N_6234,N_6921);
xnor U8078 (N_8078,N_7088,N_6455);
or U8079 (N_8079,N_7750,N_6800);
and U8080 (N_8080,N_6882,N_6851);
nor U8081 (N_8081,N_6487,N_6893);
and U8082 (N_8082,N_6262,N_7359);
or U8083 (N_8083,N_7897,N_7632);
nor U8084 (N_8084,N_7954,N_6706);
nand U8085 (N_8085,N_6665,N_7010);
or U8086 (N_8086,N_7193,N_7252);
nand U8087 (N_8087,N_6315,N_7126);
or U8088 (N_8088,N_6553,N_6867);
nand U8089 (N_8089,N_6644,N_6052);
nand U8090 (N_8090,N_7983,N_7485);
nor U8091 (N_8091,N_6222,N_6281);
nor U8092 (N_8092,N_6461,N_6954);
nand U8093 (N_8093,N_6819,N_7131);
or U8094 (N_8094,N_7976,N_7534);
or U8095 (N_8095,N_7127,N_6751);
nand U8096 (N_8096,N_6936,N_7968);
and U8097 (N_8097,N_7739,N_7503);
or U8098 (N_8098,N_6865,N_7598);
nand U8099 (N_8099,N_7640,N_7212);
or U8100 (N_8100,N_7570,N_7360);
and U8101 (N_8101,N_7426,N_7147);
and U8102 (N_8102,N_6062,N_7877);
and U8103 (N_8103,N_6721,N_7567);
or U8104 (N_8104,N_7321,N_7220);
nand U8105 (N_8105,N_7807,N_6210);
xnor U8106 (N_8106,N_6280,N_7066);
nand U8107 (N_8107,N_6570,N_7263);
and U8108 (N_8108,N_7918,N_7823);
or U8109 (N_8109,N_7862,N_6131);
and U8110 (N_8110,N_6146,N_6774);
or U8111 (N_8111,N_6595,N_6314);
or U8112 (N_8112,N_7999,N_6196);
and U8113 (N_8113,N_6463,N_7710);
or U8114 (N_8114,N_6666,N_6071);
and U8115 (N_8115,N_6551,N_7472);
or U8116 (N_8116,N_6801,N_6104);
nor U8117 (N_8117,N_7356,N_6065);
or U8118 (N_8118,N_6496,N_7630);
or U8119 (N_8119,N_6444,N_6951);
and U8120 (N_8120,N_6043,N_7585);
nor U8121 (N_8121,N_7161,N_6192);
and U8122 (N_8122,N_7952,N_6535);
xor U8123 (N_8123,N_7247,N_6050);
nand U8124 (N_8124,N_6670,N_6685);
and U8125 (N_8125,N_7856,N_6763);
or U8126 (N_8126,N_6957,N_7042);
xnor U8127 (N_8127,N_6092,N_6618);
xnor U8128 (N_8128,N_7960,N_7757);
nor U8129 (N_8129,N_7746,N_6344);
nand U8130 (N_8130,N_7781,N_6704);
and U8131 (N_8131,N_7505,N_7660);
or U8132 (N_8132,N_6888,N_6662);
or U8133 (N_8133,N_7300,N_6250);
nand U8134 (N_8134,N_6517,N_6326);
and U8135 (N_8135,N_6224,N_6711);
and U8136 (N_8136,N_7620,N_7307);
or U8137 (N_8137,N_7838,N_7001);
nand U8138 (N_8138,N_7732,N_7103);
and U8139 (N_8139,N_6816,N_6433);
nand U8140 (N_8140,N_6288,N_7711);
or U8141 (N_8141,N_7339,N_7608);
and U8142 (N_8142,N_6735,N_7964);
or U8143 (N_8143,N_6329,N_6371);
nand U8144 (N_8144,N_7308,N_7970);
or U8145 (N_8145,N_7342,N_6486);
and U8146 (N_8146,N_7115,N_6724);
and U8147 (N_8147,N_6324,N_6952);
xor U8148 (N_8148,N_7043,N_7661);
or U8149 (N_8149,N_6133,N_7336);
nand U8150 (N_8150,N_6264,N_7771);
nand U8151 (N_8151,N_6843,N_6502);
nand U8152 (N_8152,N_7454,N_7248);
nor U8153 (N_8153,N_6028,N_7973);
nand U8154 (N_8154,N_7910,N_6384);
or U8155 (N_8155,N_6325,N_7888);
or U8156 (N_8156,N_6140,N_6102);
nor U8157 (N_8157,N_7148,N_6100);
or U8158 (N_8158,N_6533,N_6826);
or U8159 (N_8159,N_7639,N_7216);
and U8160 (N_8160,N_7648,N_6992);
and U8161 (N_8161,N_6039,N_6188);
and U8162 (N_8162,N_6821,N_6034);
or U8163 (N_8163,N_7438,N_6220);
or U8164 (N_8164,N_7084,N_6010);
nor U8165 (N_8165,N_7206,N_6380);
nor U8166 (N_8166,N_6478,N_7866);
or U8167 (N_8167,N_7041,N_6309);
nand U8168 (N_8168,N_6790,N_6562);
nor U8169 (N_8169,N_6943,N_7618);
or U8170 (N_8170,N_6006,N_7722);
nor U8171 (N_8171,N_7494,N_6624);
xor U8172 (N_8172,N_7676,N_7372);
or U8173 (N_8173,N_6521,N_6169);
or U8174 (N_8174,N_6253,N_7121);
or U8175 (N_8175,N_7574,N_6616);
nand U8176 (N_8176,N_7865,N_6120);
nand U8177 (N_8177,N_7328,N_6026);
or U8178 (N_8178,N_7150,N_6881);
nor U8179 (N_8179,N_7749,N_6530);
nand U8180 (N_8180,N_6519,N_7754);
or U8181 (N_8181,N_6080,N_6771);
nor U8182 (N_8182,N_6753,N_6467);
nand U8183 (N_8183,N_7994,N_7030);
nand U8184 (N_8184,N_7700,N_7013);
nor U8185 (N_8185,N_7433,N_6910);
and U8186 (N_8186,N_6555,N_7530);
or U8187 (N_8187,N_6628,N_6938);
and U8188 (N_8188,N_7319,N_6231);
or U8189 (N_8189,N_6740,N_6437);
xor U8190 (N_8190,N_6417,N_6300);
nor U8191 (N_8191,N_6000,N_6791);
or U8192 (N_8192,N_7515,N_6838);
and U8193 (N_8193,N_6889,N_7784);
nand U8194 (N_8194,N_6869,N_6173);
nand U8195 (N_8195,N_7587,N_7853);
xor U8196 (N_8196,N_7289,N_7687);
nor U8197 (N_8197,N_7997,N_6223);
nor U8198 (N_8198,N_6686,N_7021);
nor U8199 (N_8199,N_6337,N_6664);
xnor U8200 (N_8200,N_7487,N_6975);
and U8201 (N_8201,N_7471,N_6185);
nor U8202 (N_8202,N_6633,N_6859);
nand U8203 (N_8203,N_7926,N_6336);
or U8204 (N_8204,N_6585,N_7376);
nor U8205 (N_8205,N_7099,N_6515);
nand U8206 (N_8206,N_6345,N_7219);
nor U8207 (N_8207,N_7179,N_6558);
or U8208 (N_8208,N_6126,N_6232);
and U8209 (N_8209,N_7898,N_6901);
or U8210 (N_8210,N_6895,N_6009);
xor U8211 (N_8211,N_7544,N_6758);
nor U8212 (N_8212,N_7170,N_7698);
nand U8213 (N_8213,N_7518,N_6374);
xor U8214 (N_8214,N_6450,N_7681);
xnor U8215 (N_8215,N_7626,N_7832);
and U8216 (N_8216,N_7380,N_7929);
or U8217 (N_8217,N_6967,N_6612);
and U8218 (N_8218,N_7404,N_7755);
and U8219 (N_8219,N_6073,N_7800);
nor U8220 (N_8220,N_6831,N_7065);
and U8221 (N_8221,N_7940,N_7304);
or U8222 (N_8222,N_6506,N_7458);
or U8223 (N_8223,N_7427,N_7572);
xor U8224 (N_8224,N_7741,N_7641);
and U8225 (N_8225,N_6246,N_7354);
or U8226 (N_8226,N_6900,N_6702);
nand U8227 (N_8227,N_6839,N_6498);
xor U8228 (N_8228,N_7605,N_7816);
xor U8229 (N_8229,N_6592,N_7306);
or U8230 (N_8230,N_7264,N_7812);
and U8231 (N_8231,N_7774,N_6755);
and U8232 (N_8232,N_6066,N_7532);
nand U8233 (N_8233,N_7966,N_6750);
and U8234 (N_8234,N_7191,N_6454);
nor U8235 (N_8235,N_7155,N_6797);
and U8236 (N_8236,N_6135,N_7818);
nand U8237 (N_8237,N_7791,N_6708);
and U8238 (N_8238,N_7441,N_7797);
nand U8239 (N_8239,N_7675,N_6387);
or U8240 (N_8240,N_6239,N_7158);
and U8241 (N_8241,N_7344,N_7694);
nand U8242 (N_8242,N_6934,N_7275);
xor U8243 (N_8243,N_7367,N_7390);
and U8244 (N_8244,N_6923,N_6001);
and U8245 (N_8245,N_7470,N_6822);
nor U8246 (N_8246,N_7569,N_6757);
xnor U8247 (N_8247,N_7527,N_6637);
and U8248 (N_8248,N_7346,N_6574);
nand U8249 (N_8249,N_6853,N_6605);
xor U8250 (N_8250,N_7600,N_7392);
and U8251 (N_8251,N_6037,N_6656);
xnor U8252 (N_8252,N_7075,N_6557);
nand U8253 (N_8253,N_6382,N_7950);
nand U8254 (N_8254,N_6508,N_6347);
and U8255 (N_8255,N_7081,N_7703);
nor U8256 (N_8256,N_7364,N_7798);
or U8257 (N_8257,N_7627,N_6064);
or U8258 (N_8258,N_7060,N_7284);
nand U8259 (N_8259,N_7347,N_7915);
nor U8260 (N_8260,N_7769,N_6691);
nand U8261 (N_8261,N_6582,N_6658);
and U8262 (N_8262,N_7629,N_7551);
nor U8263 (N_8263,N_7421,N_6195);
nand U8264 (N_8264,N_7516,N_7748);
nor U8265 (N_8265,N_7241,N_6683);
or U8266 (N_8266,N_6805,N_7524);
or U8267 (N_8267,N_6688,N_6305);
xor U8268 (N_8268,N_7666,N_6471);
and U8269 (N_8269,N_6412,N_6678);
and U8270 (N_8270,N_6306,N_7819);
and U8271 (N_8271,N_6200,N_6842);
and U8272 (N_8272,N_7061,N_7536);
nand U8273 (N_8273,N_6675,N_6268);
or U8274 (N_8274,N_7162,N_6060);
nor U8275 (N_8275,N_6673,N_7815);
and U8276 (N_8276,N_6377,N_6573);
nand U8277 (N_8277,N_6491,N_7902);
and U8278 (N_8278,N_7900,N_7658);
or U8279 (N_8279,N_6067,N_7314);
and U8280 (N_8280,N_7413,N_6172);
nor U8281 (N_8281,N_6602,N_6410);
or U8282 (N_8282,N_6855,N_6554);
nor U8283 (N_8283,N_7669,N_7334);
or U8284 (N_8284,N_6360,N_6032);
nand U8285 (N_8285,N_6151,N_7189);
and U8286 (N_8286,N_7285,N_6969);
or U8287 (N_8287,N_7096,N_7149);
nor U8288 (N_8288,N_6453,N_6890);
or U8289 (N_8289,N_6768,N_6581);
nor U8290 (N_8290,N_6144,N_7302);
and U8291 (N_8291,N_7005,N_7282);
nand U8292 (N_8292,N_7599,N_6654);
and U8293 (N_8293,N_7274,N_6321);
nand U8294 (N_8294,N_6677,N_6627);
nand U8295 (N_8295,N_6162,N_7269);
nor U8296 (N_8296,N_7895,N_6982);
nand U8297 (N_8297,N_7337,N_6114);
nand U8298 (N_8298,N_7208,N_6055);
nor U8299 (N_8299,N_6512,N_6424);
nor U8300 (N_8300,N_6441,N_6002);
and U8301 (N_8301,N_6566,N_6995);
nor U8302 (N_8302,N_7979,N_7117);
nand U8303 (N_8303,N_7844,N_7603);
or U8304 (N_8304,N_7697,N_7178);
and U8305 (N_8305,N_7692,N_6875);
and U8306 (N_8306,N_6917,N_7429);
nor U8307 (N_8307,N_7169,N_7343);
nand U8308 (N_8308,N_6922,N_7019);
xor U8309 (N_8309,N_7459,N_6976);
or U8310 (N_8310,N_6017,N_7371);
nand U8311 (N_8311,N_7036,N_7104);
nor U8312 (N_8312,N_6525,N_7672);
and U8313 (N_8313,N_6935,N_7882);
nor U8314 (N_8314,N_7827,N_6507);
or U8315 (N_8315,N_6204,N_6304);
nand U8316 (N_8316,N_6705,N_6235);
nand U8317 (N_8317,N_7949,N_6024);
xor U8318 (N_8318,N_6458,N_6898);
or U8319 (N_8319,N_6667,N_7649);
or U8320 (N_8320,N_7932,N_6490);
and U8321 (N_8321,N_6733,N_6813);
xnor U8322 (N_8322,N_7777,N_6275);
nor U8323 (N_8323,N_7820,N_6649);
nor U8324 (N_8324,N_6416,N_7277);
nand U8325 (N_8325,N_7958,N_7631);
and U8326 (N_8326,N_7504,N_6054);
xnor U8327 (N_8327,N_7192,N_7794);
xnor U8328 (N_8328,N_6245,N_7276);
nand U8329 (N_8329,N_7773,N_7971);
or U8330 (N_8330,N_6872,N_6395);
or U8331 (N_8331,N_7792,N_6840);
or U8332 (N_8332,N_6989,N_6479);
nand U8333 (N_8333,N_7457,N_7093);
or U8334 (N_8334,N_7137,N_7028);
xor U8335 (N_8335,N_7226,N_7468);
nand U8336 (N_8336,N_6937,N_7645);
or U8337 (N_8337,N_6156,N_6459);
and U8338 (N_8338,N_6056,N_7035);
or U8339 (N_8339,N_7288,N_6023);
nor U8340 (N_8340,N_7016,N_7581);
xnor U8341 (N_8341,N_6657,N_6780);
and U8342 (N_8342,N_7431,N_6607);
nand U8343 (N_8343,N_6550,N_6744);
and U8344 (N_8344,N_7545,N_6825);
nand U8345 (N_8345,N_6348,N_6390);
nor U8346 (N_8346,N_6342,N_7154);
nor U8347 (N_8347,N_7243,N_6516);
or U8348 (N_8348,N_7232,N_6447);
nand U8349 (N_8349,N_6308,N_6332);
xnor U8350 (N_8350,N_6105,N_6394);
or U8351 (N_8351,N_6423,N_6762);
nand U8352 (N_8352,N_7576,N_6241);
and U8353 (N_8353,N_6671,N_7984);
or U8354 (N_8354,N_6697,N_7801);
and U8355 (N_8355,N_6138,N_7136);
xnor U8356 (N_8356,N_6505,N_7716);
nand U8357 (N_8357,N_7842,N_6208);
or U8358 (N_8358,N_6913,N_6426);
nor U8359 (N_8359,N_7111,N_7240);
and U8360 (N_8360,N_7786,N_7606);
xnor U8361 (N_8361,N_7062,N_6401);
nand U8362 (N_8362,N_7802,N_6715);
nor U8363 (N_8363,N_7465,N_6086);
or U8364 (N_8364,N_7765,N_7180);
nand U8365 (N_8365,N_6008,N_7486);
nand U8366 (N_8366,N_7292,N_7410);
or U8367 (N_8367,N_7133,N_6534);
or U8368 (N_8368,N_7481,N_7009);
nand U8369 (N_8369,N_7623,N_7411);
nand U8370 (N_8370,N_6057,N_7448);
nor U8371 (N_8371,N_6481,N_6645);
nand U8372 (N_8372,N_6802,N_7922);
nor U8373 (N_8373,N_7824,N_6739);
xor U8374 (N_8374,N_7480,N_6148);
nand U8375 (N_8375,N_7405,N_7267);
and U8376 (N_8376,N_6069,N_7553);
and U8377 (N_8377,N_6472,N_7869);
xnor U8378 (N_8378,N_7756,N_6389);
or U8379 (N_8379,N_7859,N_6863);
and U8380 (N_8380,N_7353,N_6396);
or U8381 (N_8381,N_7097,N_6299);
nand U8382 (N_8382,N_6742,N_6583);
nand U8383 (N_8383,N_6405,N_6812);
and U8384 (N_8384,N_7143,N_7682);
or U8385 (N_8385,N_7221,N_6435);
and U8386 (N_8386,N_7333,N_6263);
nand U8387 (N_8387,N_6544,N_6323);
or U8388 (N_8388,N_7596,N_6227);
xor U8389 (N_8389,N_7841,N_6591);
nor U8390 (N_8390,N_7981,N_7830);
and U8391 (N_8391,N_6916,N_6407);
or U8392 (N_8392,N_6122,N_6784);
nand U8393 (N_8393,N_6852,N_6119);
and U8394 (N_8394,N_7621,N_6074);
nand U8395 (N_8395,N_7293,N_7879);
and U8396 (N_8396,N_7455,N_6388);
nand U8397 (N_8397,N_7957,N_6385);
or U8398 (N_8398,N_6787,N_6880);
and U8399 (N_8399,N_7959,N_6252);
or U8400 (N_8400,N_6256,N_7597);
and U8401 (N_8401,N_7038,N_7961);
nor U8402 (N_8402,N_7988,N_6707);
and U8403 (N_8403,N_6340,N_7691);
and U8404 (N_8404,N_6904,N_7951);
and U8405 (N_8405,N_7298,N_7083);
or U8406 (N_8406,N_6249,N_7962);
and U8407 (N_8407,N_7956,N_7159);
nor U8408 (N_8408,N_7591,N_7644);
and U8409 (N_8409,N_7592,N_7510);
and U8410 (N_8410,N_6524,N_7745);
nand U8411 (N_8411,N_6351,N_7482);
or U8412 (N_8412,N_7217,N_6694);
nor U8413 (N_8413,N_7407,N_7790);
or U8414 (N_8414,N_6457,N_6640);
and U8415 (N_8415,N_6878,N_6015);
or U8416 (N_8416,N_7320,N_6700);
nor U8417 (N_8417,N_6903,N_6358);
nand U8418 (N_8418,N_7890,N_6484);
nand U8419 (N_8419,N_6817,N_7871);
and U8420 (N_8420,N_6476,N_7892);
nand U8421 (N_8421,N_6862,N_7129);
nor U8422 (N_8422,N_7449,N_6848);
nand U8423 (N_8423,N_6599,N_7759);
nor U8424 (N_8424,N_7456,N_7012);
or U8425 (N_8425,N_7370,N_7329);
and U8426 (N_8426,N_6286,N_7513);
nor U8427 (N_8427,N_7375,N_6183);
xor U8428 (N_8428,N_7017,N_6415);
nand U8429 (N_8429,N_6679,N_7727);
nor U8430 (N_8430,N_6291,N_6118);
nand U8431 (N_8431,N_6829,N_7870);
xnor U8432 (N_8432,N_6729,N_7876);
nand U8433 (N_8433,N_6690,N_7989);
nand U8434 (N_8434,N_7230,N_7717);
nor U8435 (N_8435,N_7141,N_7963);
xor U8436 (N_8436,N_6567,N_7695);
nor U8437 (N_8437,N_7995,N_7693);
and U8438 (N_8438,N_7070,N_7224);
nand U8439 (N_8439,N_7848,N_7927);
and U8440 (N_8440,N_6531,N_6451);
or U8441 (N_8441,N_6925,N_6011);
xnor U8442 (N_8442,N_7175,N_7785);
xnor U8443 (N_8443,N_6150,N_6902);
nand U8444 (N_8444,N_6199,N_7817);
nor U8445 (N_8445,N_6095,N_6808);
xnor U8446 (N_8446,N_7779,N_7165);
and U8447 (N_8447,N_7027,N_6301);
and U8448 (N_8448,N_7047,N_6497);
nand U8449 (N_8449,N_7437,N_7942);
nor U8450 (N_8450,N_7297,N_7414);
or U8451 (N_8451,N_6198,N_7140);
xnor U8452 (N_8452,N_6907,N_6021);
or U8453 (N_8453,N_6597,N_6373);
and U8454 (N_8454,N_7560,N_7533);
nor U8455 (N_8455,N_7254,N_6386);
nand U8456 (N_8456,N_7054,N_6101);
nor U8457 (N_8457,N_7938,N_6626);
nand U8458 (N_8458,N_6364,N_6214);
nor U8459 (N_8459,N_6868,N_6058);
or U8460 (N_8460,N_7562,N_7561);
nor U8461 (N_8461,N_7260,N_7102);
nand U8462 (N_8462,N_6560,N_7690);
nor U8463 (N_8463,N_6950,N_7280);
or U8464 (N_8464,N_7229,N_6155);
nand U8465 (N_8465,N_6611,N_7315);
xor U8466 (N_8466,N_7056,N_6620);
and U8467 (N_8467,N_6294,N_7969);
and U8468 (N_8468,N_6282,N_6603);
and U8469 (N_8469,N_7633,N_6652);
or U8470 (N_8470,N_6335,N_7747);
nor U8471 (N_8471,N_7855,N_7461);
nor U8472 (N_8472,N_7120,N_6089);
nand U8473 (N_8473,N_7685,N_6876);
nand U8474 (N_8474,N_7937,N_6537);
or U8475 (N_8475,N_7829,N_7993);
nor U8476 (N_8476,N_6190,N_7875);
nor U8477 (N_8477,N_7702,N_7255);
or U8478 (N_8478,N_7612,N_6614);
nand U8479 (N_8479,N_7619,N_7157);
and U8480 (N_8480,N_6322,N_6087);
nor U8481 (N_8481,N_6258,N_6350);
or U8482 (N_8482,N_6432,N_6928);
or U8483 (N_8483,N_7008,N_7132);
nor U8484 (N_8484,N_6804,N_7273);
nor U8485 (N_8485,N_7068,N_6097);
and U8486 (N_8486,N_6617,N_6170);
nor U8487 (N_8487,N_7167,N_6063);
and U8488 (N_8488,N_6355,N_6956);
nor U8489 (N_8489,N_6810,N_7018);
nand U8490 (N_8490,N_7144,N_7326);
nand U8491 (N_8491,N_6418,N_7207);
nand U8492 (N_8492,N_6356,N_6579);
or U8493 (N_8493,N_7982,N_6098);
nand U8494 (N_8494,N_6287,N_7889);
and U8495 (N_8495,N_6110,N_6661);
and U8496 (N_8496,N_7283,N_6996);
and U8497 (N_8497,N_7110,N_7874);
and U8498 (N_8498,N_7907,N_7044);
nand U8499 (N_8499,N_7767,N_6462);
or U8500 (N_8500,N_6911,N_7535);
or U8501 (N_8501,N_7974,N_7594);
nor U8502 (N_8502,N_6964,N_6716);
and U8503 (N_8503,N_7031,N_6760);
or U8504 (N_8504,N_7944,N_7839);
nand U8505 (N_8505,N_6796,N_7190);
nand U8506 (N_8506,N_7138,N_7135);
or U8507 (N_8507,N_6130,N_6206);
nand U8508 (N_8508,N_6427,N_7338);
nand U8509 (N_8509,N_6885,N_6777);
and U8510 (N_8510,N_6022,N_7601);
or U8511 (N_8511,N_7313,N_7119);
nor U8512 (N_8512,N_7721,N_7409);
or U8513 (N_8513,N_6663,N_6642);
or U8514 (N_8514,N_7520,N_6085);
nand U8515 (N_8515,N_6334,N_6720);
nor U8516 (N_8516,N_7128,N_6403);
and U8517 (N_8517,N_6365,N_7397);
nand U8518 (N_8518,N_6259,N_6277);
nand U8519 (N_8519,N_7439,N_6619);
or U8520 (N_8520,N_6174,N_7107);
nand U8521 (N_8521,N_6236,N_6307);
and U8522 (N_8522,N_7160,N_6726);
nor U8523 (N_8523,N_6465,N_7498);
nand U8524 (N_8524,N_6586,N_6932);
nor U8525 (N_8525,N_6549,N_6737);
and U8526 (N_8526,N_7381,N_7814);
nor U8527 (N_8527,N_6297,N_7556);
nand U8528 (N_8528,N_6128,N_7011);
and U8529 (N_8529,N_6674,N_7734);
and U8530 (N_8530,N_7432,N_6783);
nor U8531 (N_8531,N_7604,N_7835);
nor U8532 (N_8532,N_7378,N_7497);
nand U8533 (N_8533,N_7625,N_7256);
nand U8534 (N_8534,N_7921,N_6419);
nor U8535 (N_8535,N_6798,N_7705);
nand U8536 (N_8536,N_6404,N_7324);
nor U8537 (N_8537,N_7512,N_7425);
nor U8538 (N_8538,N_7782,N_6948);
and U8539 (N_8539,N_6955,N_6613);
and U8540 (N_8540,N_7076,N_7836);
xnor U8541 (N_8541,N_7740,N_6132);
nor U8542 (N_8542,N_7783,N_7223);
xor U8543 (N_8543,N_7125,N_7589);
and U8544 (N_8544,N_6096,N_6127);
xor U8545 (N_8545,N_6330,N_6676);
nor U8546 (N_8546,N_7873,N_6841);
and U8547 (N_8547,N_6285,N_7225);
nor U8548 (N_8548,N_7541,N_7365);
xor U8549 (N_8549,N_7887,N_7310);
nand U8550 (N_8550,N_6794,N_7444);
or U8551 (N_8551,N_6139,N_6891);
xnor U8552 (N_8552,N_6369,N_6408);
and U8553 (N_8553,N_7373,N_7399);
or U8554 (N_8554,N_6752,N_7872);
nand U8555 (N_8555,N_6042,N_7091);
or U8556 (N_8556,N_6565,N_6799);
or U8557 (N_8557,N_6070,N_7511);
nand U8558 (N_8558,N_7270,N_6115);
and U8559 (N_8559,N_6205,N_6033);
nor U8560 (N_8560,N_6860,N_7265);
or U8561 (N_8561,N_6653,N_6710);
nor U8562 (N_8562,N_7286,N_7822);
and U8563 (N_8563,N_6267,N_7696);
or U8564 (N_8564,N_7713,N_6240);
nor U8565 (N_8565,N_7116,N_7369);
or U8566 (N_8566,N_7233,N_6779);
nor U8567 (N_8567,N_7787,N_7528);
nand U8568 (N_8568,N_6584,N_7134);
and U8569 (N_8569,N_6448,N_6266);
xnor U8570 (N_8570,N_6167,N_6495);
nand U8571 (N_8571,N_7845,N_7847);
xnor U8572 (N_8572,N_7977,N_6693);
xnor U8573 (N_8573,N_6228,N_6207);
or U8574 (N_8574,N_6747,N_7123);
or U8575 (N_8575,N_7657,N_7588);
nand U8576 (N_8576,N_6473,N_7945);
and U8577 (N_8577,N_6093,N_7724);
or U8578 (N_8578,N_6594,N_7006);
xnor U8579 (N_8579,N_7151,N_7082);
nand U8580 (N_8580,N_7330,N_6164);
xnor U8581 (N_8581,N_6879,N_7435);
nor U8582 (N_8582,N_7522,N_6255);
or U8583 (N_8583,N_6545,N_6999);
and U8584 (N_8584,N_6328,N_6571);
nor U8585 (N_8585,N_7849,N_6823);
nand U8586 (N_8586,N_6449,N_7403);
or U8587 (N_8587,N_7936,N_6012);
xor U8588 (N_8588,N_6368,N_6939);
and U8589 (N_8589,N_6510,N_7523);
nor U8590 (N_8590,N_7908,N_6076);
nand U8591 (N_8591,N_7729,N_6563);
nand U8592 (N_8592,N_6078,N_7048);
and U8593 (N_8593,N_6047,N_6327);
and U8594 (N_8594,N_7362,N_7317);
and U8595 (N_8595,N_6899,N_6953);
nor U8596 (N_8596,N_6357,N_6504);
and U8597 (N_8597,N_7646,N_6141);
or U8598 (N_8598,N_6372,N_6886);
nand U8599 (N_8599,N_6414,N_7446);
and U8600 (N_8600,N_6180,N_6038);
and U8601 (N_8601,N_7316,N_7580);
and U8602 (N_8602,N_6979,N_6123);
and U8603 (N_8603,N_6019,N_7501);
and U8604 (N_8604,N_6422,N_7566);
nand U8605 (N_8605,N_6129,N_6201);
and U8606 (N_8606,N_7667,N_6470);
or U8607 (N_8607,N_6944,N_7415);
nand U8608 (N_8608,N_7358,N_7730);
nand U8609 (N_8609,N_6927,N_7939);
nand U8610 (N_8610,N_6213,N_6493);
nand U8611 (N_8611,N_7164,N_7768);
or U8612 (N_8612,N_6856,N_6143);
and U8613 (N_8613,N_7772,N_6858);
nor U8614 (N_8614,N_6920,N_6990);
or U8615 (N_8615,N_6745,N_6543);
nand U8616 (N_8616,N_6425,N_6993);
nand U8617 (N_8617,N_6828,N_7758);
or U8618 (N_8618,N_6077,N_7361);
nand U8619 (N_8619,N_7436,N_6117);
and U8620 (N_8620,N_7707,N_6806);
and U8621 (N_8621,N_6242,N_7197);
nand U8622 (N_8622,N_7831,N_6741);
or U8623 (N_8623,N_7039,N_6177);
xor U8624 (N_8624,N_7257,N_7948);
and U8625 (N_8625,N_7477,N_6257);
xnor U8626 (N_8626,N_6165,N_6346);
nor U8627 (N_8627,N_7231,N_7778);
or U8628 (N_8628,N_6238,N_6743);
and U8629 (N_8629,N_6271,N_6874);
xor U8630 (N_8630,N_7340,N_7033);
nand U8631 (N_8631,N_6809,N_7506);
or U8632 (N_8632,N_7266,N_6588);
or U8633 (N_8633,N_7901,N_6636);
and U8634 (N_8634,N_7187,N_6233);
and U8635 (N_8635,N_6727,N_7022);
nand U8636 (N_8636,N_6814,N_6379);
nand U8637 (N_8637,N_6873,N_6339);
nand U8638 (N_8638,N_6980,N_7325);
or U8639 (N_8639,N_7194,N_7301);
nor U8640 (N_8640,N_7507,N_6298);
nand U8641 (N_8641,N_7607,N_7045);
and U8642 (N_8642,N_6216,N_6699);
or U8643 (N_8643,N_6589,N_7163);
or U8644 (N_8644,N_7385,N_6475);
and U8645 (N_8645,N_6013,N_6766);
and U8646 (N_8646,N_6598,N_7218);
or U8647 (N_8647,N_6181,N_6154);
nor U8648 (N_8648,N_7215,N_6157);
xnor U8649 (N_8649,N_7508,N_7258);
nand U8650 (N_8650,N_7858,N_7546);
nand U8651 (N_8651,N_7914,N_7880);
nor U8652 (N_8652,N_7251,N_6333);
or U8653 (N_8653,N_7796,N_7460);
nand U8654 (N_8654,N_6698,N_7805);
or U8655 (N_8655,N_7014,N_6027);
and U8656 (N_8656,N_6835,N_7909);
nor U8657 (N_8657,N_6079,N_6134);
nand U8658 (N_8658,N_7762,N_6538);
xnor U8659 (N_8659,N_7057,N_6725);
nor U8660 (N_8660,N_7029,N_6520);
nor U8661 (N_8661,N_6773,N_6316);
and U8662 (N_8662,N_6445,N_7204);
or U8663 (N_8663,N_7558,N_6436);
xnor U8664 (N_8664,N_6446,N_7007);
and U8665 (N_8665,N_7857,N_7854);
nand U8666 (N_8666,N_7037,N_7234);
xnor U8667 (N_8667,N_7237,N_6575);
nor U8668 (N_8668,N_7462,N_6248);
nand U8669 (N_8669,N_7139,N_7475);
or U8670 (N_8670,N_7402,N_7495);
nand U8671 (N_8671,N_7975,N_7428);
and U8672 (N_8672,N_6542,N_7905);
or U8673 (N_8673,N_6225,N_7418);
nand U8674 (N_8674,N_6523,N_7000);
nor U8675 (N_8675,N_7327,N_6985);
and U8676 (N_8676,N_7985,N_6965);
and U8677 (N_8677,N_6049,N_6561);
or U8678 (N_8678,N_6428,N_7173);
nand U8679 (N_8679,N_6353,N_7195);
or U8680 (N_8680,N_6986,N_7529);
nor U8681 (N_8681,N_6030,N_7885);
and U8682 (N_8682,N_7202,N_7357);
and U8683 (N_8683,N_6361,N_7555);
nand U8684 (N_8684,N_6053,N_6474);
nand U8685 (N_8685,N_7978,N_6947);
nor U8686 (N_8686,N_6945,N_7704);
and U8687 (N_8687,N_7049,N_7742);
and U8688 (N_8688,N_6149,N_6005);
xor U8689 (N_8689,N_6265,N_7662);
or U8690 (N_8690,N_7559,N_6051);
nand U8691 (N_8691,N_6646,N_7184);
and U8692 (N_8692,N_6349,N_6983);
nand U8693 (N_8693,N_6732,N_6576);
nand U8694 (N_8694,N_6541,N_6811);
nor U8695 (N_8695,N_6959,N_7249);
and U8696 (N_8696,N_7253,N_7450);
or U8697 (N_8697,N_7775,N_6175);
and U8698 (N_8698,N_6375,N_7077);
nand U8699 (N_8699,N_7002,N_7737);
nor U8700 (N_8700,N_7919,N_6962);
or U8701 (N_8701,N_7568,N_6318);
or U8702 (N_8702,N_6020,N_7236);
or U8703 (N_8703,N_6713,N_6359);
nand U8704 (N_8704,N_6958,N_7677);
nor U8705 (N_8705,N_6930,N_6338);
nor U8706 (N_8706,N_6040,N_6509);
or U8707 (N_8707,N_6723,N_6278);
xor U8708 (N_8708,N_7636,N_6136);
nand U8709 (N_8709,N_7825,N_7105);
and U8710 (N_8710,N_6397,N_6734);
nor U8711 (N_8711,N_7023,N_6187);
and U8712 (N_8712,N_7332,N_6494);
nand U8713 (N_8713,N_7112,N_7986);
or U8714 (N_8714,N_6764,N_7311);
and U8715 (N_8715,N_7996,N_7751);
and U8716 (N_8716,N_6191,N_6946);
nand U8717 (N_8717,N_7679,N_7653);
nand U8718 (N_8718,N_7072,N_7776);
or U8719 (N_8719,N_7851,N_7924);
and U8720 (N_8720,N_6041,N_6528);
or U8721 (N_8721,N_7025,N_6489);
and U8722 (N_8722,N_7542,N_7764);
nor U8723 (N_8723,N_6730,N_6221);
and U8724 (N_8724,N_7795,N_6785);
or U8725 (N_8725,N_7412,N_6341);
or U8726 (N_8726,N_6914,N_7055);
and U8727 (N_8727,N_7199,N_6014);
or U8728 (N_8728,N_6601,N_6354);
xor U8729 (N_8729,N_7476,N_6756);
or U8730 (N_8730,N_6781,N_6593);
and U8731 (N_8731,N_6978,N_7205);
nand U8732 (N_8732,N_7322,N_7965);
nor U8733 (N_8733,N_6974,N_6929);
nand U8734 (N_8734,N_7181,N_6650);
or U8735 (N_8735,N_7613,N_7069);
nor U8736 (N_8736,N_7098,N_6091);
or U8737 (N_8737,N_6400,N_6638);
nor U8738 (N_8738,N_7736,N_7423);
or U8739 (N_8739,N_6896,N_6084);
xnor U8740 (N_8740,N_6492,N_7004);
nor U8741 (N_8741,N_7538,N_6572);
nor U8742 (N_8742,N_6310,N_7517);
nor U8743 (N_8743,N_7113,N_6857);
and U8744 (N_8744,N_6827,N_7388);
or U8745 (N_8745,N_7452,N_7287);
nor U8746 (N_8746,N_7656,N_7688);
nor U8747 (N_8747,N_7728,N_7122);
nand U8748 (N_8748,N_7539,N_6171);
nor U8749 (N_8749,N_7352,N_6243);
or U8750 (N_8750,N_6460,N_6391);
nand U8751 (N_8751,N_6775,N_6931);
or U8752 (N_8752,N_6477,N_6083);
xor U8753 (N_8753,N_6088,N_6776);
nand U8754 (N_8754,N_7861,N_6887);
xor U8755 (N_8755,N_7387,N_6630);
nor U8756 (N_8756,N_7593,N_7172);
and U8757 (N_8757,N_6464,N_7469);
nor U8758 (N_8758,N_7543,N_7203);
or U8759 (N_8759,N_7761,N_7899);
nand U8760 (N_8760,N_6283,N_7046);
nand U8761 (N_8761,N_6112,N_6295);
nand U8762 (N_8762,N_6655,N_6786);
nand U8763 (N_8763,N_7166,N_6376);
xor U8764 (N_8764,N_6434,N_7808);
or U8765 (N_8765,N_6844,N_6556);
or U8766 (N_8766,N_6919,N_6540);
or U8767 (N_8767,N_7374,N_6160);
or U8768 (N_8768,N_6203,N_6261);
and U8769 (N_8769,N_7200,N_7348);
xnor U8770 (N_8770,N_6648,N_6635);
or U8771 (N_8771,N_7753,N_6963);
and U8772 (N_8772,N_6398,N_7622);
and U8773 (N_8773,N_6145,N_6413);
nor U8774 (N_8774,N_6158,N_6547);
and U8775 (N_8775,N_7788,N_7349);
or U8776 (N_8776,N_7020,N_7261);
nand U8777 (N_8777,N_6659,N_7526);
xnor U8778 (N_8778,N_6580,N_7463);
nor U8779 (N_8779,N_7595,N_6442);
and U8780 (N_8780,N_7052,N_6778);
and U8781 (N_8781,N_7789,N_7770);
and U8782 (N_8782,N_7826,N_6719);
nor U8783 (N_8783,N_7925,N_6837);
nand U8784 (N_8784,N_7799,N_7318);
nor U8785 (N_8785,N_7490,N_6302);
and U8786 (N_8786,N_6099,N_6273);
or U8787 (N_8787,N_6443,N_6179);
nand U8788 (N_8788,N_7351,N_6420);
or U8789 (N_8789,N_6971,N_7916);
nand U8790 (N_8790,N_7579,N_7442);
nand U8791 (N_8791,N_6421,N_6045);
xnor U8792 (N_8792,N_7565,N_7806);
and U8793 (N_8793,N_7478,N_7554);
or U8794 (N_8794,N_6789,N_7168);
and U8795 (N_8795,N_6908,N_7643);
or U8796 (N_8796,N_6439,N_6229);
nor U8797 (N_8797,N_6623,N_6942);
nor U8798 (N_8798,N_6142,N_7473);
or U8799 (N_8799,N_6643,N_6106);
nor U8800 (N_8800,N_7514,N_6883);
or U8801 (N_8801,N_6284,N_6941);
nor U8802 (N_8802,N_7735,N_7893);
nor U8803 (N_8803,N_7709,N_6961);
nand U8804 (N_8804,N_7474,N_6513);
and U8805 (N_8805,N_6933,N_6871);
and U8806 (N_8806,N_7145,N_7445);
or U8807 (N_8807,N_7917,N_7654);
xor U8808 (N_8808,N_7674,N_7493);
or U8809 (N_8809,N_6834,N_7447);
or U8810 (N_8810,N_6312,N_6168);
nand U8811 (N_8811,N_6035,N_7272);
or U8812 (N_8812,N_7793,N_7467);
and U8813 (N_8813,N_6279,N_6854);
nor U8814 (N_8814,N_7440,N_7689);
nand U8815 (N_8815,N_7094,N_7106);
nand U8816 (N_8816,N_7384,N_6367);
nor U8817 (N_8817,N_7699,N_7156);
nand U8818 (N_8818,N_7840,N_7395);
nor U8819 (N_8819,N_7718,N_7624);
nand U8820 (N_8820,N_7419,N_6153);
or U8821 (N_8821,N_7683,N_6219);
nand U8822 (N_8822,N_7079,N_6606);
nor U8823 (N_8823,N_7953,N_7990);
nand U8824 (N_8824,N_7491,N_7443);
nand U8825 (N_8825,N_6803,N_7171);
nor U8826 (N_8826,N_7095,N_7537);
or U8827 (N_8827,N_6260,N_7034);
nand U8828 (N_8828,N_7864,N_6940);
and U8829 (N_8829,N_7637,N_7863);
and U8830 (N_8830,N_6202,N_7386);
xor U8831 (N_8831,N_6392,N_7214);
nor U8832 (N_8832,N_6244,N_6604);
or U8833 (N_8833,N_7634,N_7904);
nor U8834 (N_8834,N_6107,N_6343);
nand U8835 (N_8835,N_6681,N_7780);
nor U8836 (N_8836,N_6552,N_6877);
nor U8837 (N_8837,N_7430,N_7089);
nand U8838 (N_8838,N_6894,N_6615);
and U8839 (N_8839,N_7763,N_7379);
xnor U8840 (N_8840,N_7733,N_6824);
nor U8841 (N_8841,N_7130,N_7884);
or U8842 (N_8842,N_7063,N_6850);
or U8843 (N_8843,N_7262,N_6193);
and U8844 (N_8844,N_6217,N_6609);
and U8845 (N_8845,N_7182,N_7933);
or U8846 (N_8846,N_7578,N_7394);
and U8847 (N_8847,N_7114,N_6973);
nor U8848 (N_8848,N_7400,N_7803);
nor U8849 (N_8849,N_7331,N_6081);
nand U8850 (N_8850,N_7972,N_7843);
nor U8851 (N_8851,N_7355,N_6701);
xnor U8852 (N_8852,N_6163,N_6254);
or U8853 (N_8853,N_7810,N_6075);
and U8854 (N_8854,N_7059,N_7488);
nand U8855 (N_8855,N_6276,N_7309);
nand U8856 (N_8856,N_7575,N_7913);
or U8857 (N_8857,N_7886,N_6503);
nand U8858 (N_8858,N_7615,N_7101);
or U8859 (N_8859,N_6578,N_6468);
and U8860 (N_8860,N_6176,N_6861);
nand U8861 (N_8861,N_6717,N_7868);
and U8862 (N_8862,N_7335,N_6480);
nor U8863 (N_8863,N_7955,N_6499);
nor U8864 (N_8864,N_6782,N_7701);
xor U8865 (N_8865,N_6915,N_6968);
and U8866 (N_8866,N_6044,N_6641);
nor U8867 (N_8867,N_7196,N_7571);
nor U8868 (N_8868,N_7731,N_6313);
nand U8869 (N_8869,N_7185,N_7715);
nand U8870 (N_8870,N_6590,N_6818);
nor U8871 (N_8871,N_6320,N_6511);
xor U8872 (N_8872,N_6452,N_6987);
and U8873 (N_8873,N_7424,N_6608);
nand U8874 (N_8874,N_6680,N_6892);
nand U8875 (N_8875,N_6482,N_6864);
or U8876 (N_8876,N_7417,N_6378);
and U8877 (N_8877,N_7484,N_7296);
or U8878 (N_8878,N_6629,N_6189);
nor U8879 (N_8879,N_6714,N_7867);
or U8880 (N_8880,N_7828,N_6728);
and U8881 (N_8881,N_6269,N_7881);
nor U8882 (N_8882,N_7766,N_7714);
xor U8883 (N_8883,N_6634,N_7552);
nor U8884 (N_8884,N_6438,N_7222);
or U8885 (N_8885,N_7250,N_6296);
or U8886 (N_8886,N_6912,N_6621);
and U8887 (N_8887,N_7235,N_7651);
and U8888 (N_8888,N_6926,N_6536);
nand U8889 (N_8889,N_6988,N_7198);
nor U8890 (N_8890,N_6548,N_7073);
and U8891 (N_8891,N_6568,N_7928);
nor U8892 (N_8892,N_6247,N_7614);
nand U8893 (N_8893,N_7032,N_6366);
or U8894 (N_8894,N_7092,N_6485);
xnor U8895 (N_8895,N_7176,N_7177);
nor U8896 (N_8896,N_7401,N_6994);
nand U8897 (N_8897,N_7211,N_6529);
and U8898 (N_8898,N_6352,N_6381);
and U8899 (N_8899,N_7453,N_7744);
nand U8900 (N_8900,N_7671,N_7896);
nor U8901 (N_8901,N_6696,N_6749);
nand U8902 (N_8902,N_7617,N_7398);
and U8903 (N_8903,N_7708,N_6909);
or U8904 (N_8904,N_7209,N_7638);
nor U8905 (N_8905,N_6108,N_7894);
xnor U8906 (N_8906,N_6639,N_6748);
or U8907 (N_8907,N_6712,N_6695);
nor U8908 (N_8908,N_7992,N_7563);
or U8909 (N_8909,N_7647,N_6754);
nand U8910 (N_8910,N_6025,N_6632);
nand U8911 (N_8911,N_6722,N_6016);
xnor U8912 (N_8912,N_7259,N_6409);
or U8913 (N_8913,N_6564,N_7834);
or U8914 (N_8914,N_6226,N_7980);
nor U8915 (N_8915,N_7239,N_6815);
nor U8916 (N_8916,N_7090,N_7074);
or U8917 (N_8917,N_7719,N_7124);
or U8918 (N_8918,N_6610,N_7531);
xor U8919 (N_8919,N_6383,N_7642);
xor U8920 (N_8920,N_7201,N_6845);
or U8921 (N_8921,N_7821,N_6765);
nor U8922 (N_8922,N_7628,N_6532);
and U8923 (N_8923,N_7050,N_6622);
nand U8924 (N_8924,N_6905,N_7935);
or U8925 (N_8925,N_7586,N_7271);
and U8926 (N_8926,N_6596,N_7281);
and U8927 (N_8927,N_6215,N_6137);
nor U8928 (N_8928,N_6212,N_7991);
nor U8929 (N_8929,N_7268,N_6846);
nand U8930 (N_8930,N_6331,N_6849);
or U8931 (N_8931,N_7502,N_6709);
nor U8932 (N_8932,N_7943,N_6293);
nand U8933 (N_8933,N_7998,N_7519);
or U8934 (N_8934,N_7712,N_6736);
and U8935 (N_8935,N_7228,N_6997);
nor U8936 (N_8936,N_7564,N_6317);
nand U8937 (N_8937,N_6430,N_7878);
or U8938 (N_8938,N_6669,N_6832);
and U8939 (N_8939,N_6836,N_6211);
nor U8940 (N_8940,N_7024,N_6672);
nor U8941 (N_8941,N_7549,N_6431);
nand U8942 (N_8942,N_6906,N_6147);
and U8943 (N_8943,N_6178,N_7078);
and U8944 (N_8944,N_6960,N_6272);
and U8945 (N_8945,N_6194,N_6625);
or U8946 (N_8946,N_6270,N_7368);
and U8947 (N_8947,N_6363,N_6186);
and U8948 (N_8948,N_7213,N_6647);
nor U8949 (N_8949,N_7743,N_7246);
nand U8950 (N_8950,N_7323,N_7941);
and U8951 (N_8951,N_7279,N_6703);
and U8952 (N_8952,N_6068,N_7852);
or U8953 (N_8953,N_7087,N_6061);
nand U8954 (N_8954,N_6440,N_6103);
nand U8955 (N_8955,N_6539,N_7813);
nand U8956 (N_8956,N_7363,N_6488);
nor U8957 (N_8957,N_7602,N_6237);
and U8958 (N_8958,N_6251,N_6738);
nand U8959 (N_8959,N_7466,N_7720);
nand U8960 (N_8960,N_6770,N_6631);
xor U8961 (N_8961,N_6218,N_6518);
or U8962 (N_8962,N_7573,N_6746);
nand U8963 (N_8963,N_6161,N_7245);
or U8964 (N_8964,N_6111,N_6830);
nor U8965 (N_8965,N_6759,N_6966);
nor U8966 (N_8966,N_6116,N_7655);
nand U8967 (N_8967,N_7383,N_7242);
nor U8968 (N_8968,N_6731,N_7663);
nand U8969 (N_8969,N_7238,N_7408);
or U8970 (N_8970,N_7726,N_7911);
nand U8971 (N_8971,N_7912,N_7051);
nor U8972 (N_8972,N_6660,N_7723);
nand U8973 (N_8973,N_7582,N_7142);
or U8974 (N_8974,N_7906,N_6772);
nand U8975 (N_8975,N_7118,N_7389);
nor U8976 (N_8976,N_7422,N_6292);
nand U8977 (N_8977,N_6682,N_6311);
nor U8978 (N_8978,N_7227,N_7548);
xnor U8979 (N_8979,N_7760,N_7521);
nand U8980 (N_8980,N_7026,N_6820);
nor U8981 (N_8981,N_7931,N_6884);
and U8982 (N_8982,N_7278,N_6289);
or U8983 (N_8983,N_7109,N_7652);
nand U8984 (N_8984,N_6651,N_6918);
nor U8985 (N_8985,N_7188,N_6399);
or U8986 (N_8986,N_6402,N_7003);
and U8987 (N_8987,N_7067,N_6124);
or U8988 (N_8988,N_7725,N_6769);
and U8989 (N_8989,N_7420,N_7610);
nand U8990 (N_8990,N_6031,N_6981);
or U8991 (N_8991,N_6526,N_6977);
xor U8992 (N_8992,N_7391,N_7811);
nor U8993 (N_8993,N_6577,N_6792);
nor U8994 (N_8994,N_7345,N_7583);
and U8995 (N_8995,N_7659,N_7341);
or U8996 (N_8996,N_6290,N_6319);
or U8997 (N_8997,N_7406,N_6230);
or U8998 (N_8998,N_6456,N_6483);
nand U8999 (N_8999,N_7393,N_6514);
nand U9000 (N_9000,N_7165,N_6491);
nor U9001 (N_9001,N_6972,N_6599);
and U9002 (N_9002,N_7709,N_7190);
nand U9003 (N_9003,N_7833,N_6083);
and U9004 (N_9004,N_6044,N_7759);
or U9005 (N_9005,N_6505,N_7727);
or U9006 (N_9006,N_6626,N_6086);
or U9007 (N_9007,N_7444,N_6320);
nor U9008 (N_9008,N_6207,N_7200);
or U9009 (N_9009,N_6302,N_6581);
nand U9010 (N_9010,N_7105,N_7525);
nand U9011 (N_9011,N_7902,N_7520);
nor U9012 (N_9012,N_7838,N_7554);
nand U9013 (N_9013,N_6041,N_7778);
nand U9014 (N_9014,N_6828,N_7963);
and U9015 (N_9015,N_7310,N_6450);
nand U9016 (N_9016,N_7253,N_7960);
or U9017 (N_9017,N_7020,N_6016);
or U9018 (N_9018,N_7988,N_6480);
or U9019 (N_9019,N_6244,N_6732);
nand U9020 (N_9020,N_6798,N_6901);
nand U9021 (N_9021,N_6624,N_6101);
nand U9022 (N_9022,N_6463,N_6685);
or U9023 (N_9023,N_6318,N_6406);
xnor U9024 (N_9024,N_7144,N_7552);
or U9025 (N_9025,N_7643,N_7411);
nand U9026 (N_9026,N_7931,N_6385);
xor U9027 (N_9027,N_6659,N_7575);
nand U9028 (N_9028,N_6971,N_7413);
nor U9029 (N_9029,N_6772,N_6895);
and U9030 (N_9030,N_7699,N_6656);
or U9031 (N_9031,N_6406,N_6015);
xnor U9032 (N_9032,N_7767,N_6855);
and U9033 (N_9033,N_6271,N_7042);
nand U9034 (N_9034,N_6912,N_6587);
and U9035 (N_9035,N_6091,N_7851);
nor U9036 (N_9036,N_6660,N_6352);
and U9037 (N_9037,N_7014,N_6923);
and U9038 (N_9038,N_6246,N_6124);
nor U9039 (N_9039,N_7147,N_7825);
and U9040 (N_9040,N_6051,N_6443);
or U9041 (N_9041,N_6380,N_7281);
nand U9042 (N_9042,N_6714,N_6874);
and U9043 (N_9043,N_7597,N_7149);
nor U9044 (N_9044,N_6678,N_6363);
or U9045 (N_9045,N_6519,N_6465);
nand U9046 (N_9046,N_6369,N_6844);
nor U9047 (N_9047,N_6755,N_7183);
nor U9048 (N_9048,N_7290,N_6183);
nor U9049 (N_9049,N_7936,N_6385);
xnor U9050 (N_9050,N_6963,N_6974);
nand U9051 (N_9051,N_6737,N_7768);
and U9052 (N_9052,N_6165,N_7122);
or U9053 (N_9053,N_6628,N_6143);
and U9054 (N_9054,N_6985,N_7995);
xor U9055 (N_9055,N_6015,N_7100);
and U9056 (N_9056,N_6693,N_6979);
nand U9057 (N_9057,N_6575,N_6149);
nand U9058 (N_9058,N_6316,N_6334);
nand U9059 (N_9059,N_7865,N_7323);
and U9060 (N_9060,N_7446,N_7878);
and U9061 (N_9061,N_7438,N_7252);
nor U9062 (N_9062,N_6129,N_6199);
or U9063 (N_9063,N_7865,N_6307);
nand U9064 (N_9064,N_6728,N_6919);
nand U9065 (N_9065,N_6971,N_7452);
and U9066 (N_9066,N_6584,N_7451);
or U9067 (N_9067,N_6098,N_6555);
nor U9068 (N_9068,N_6071,N_6730);
or U9069 (N_9069,N_6606,N_7921);
and U9070 (N_9070,N_7140,N_7520);
nor U9071 (N_9071,N_6942,N_7454);
nand U9072 (N_9072,N_7852,N_7653);
or U9073 (N_9073,N_6894,N_7258);
xor U9074 (N_9074,N_6088,N_7760);
nor U9075 (N_9075,N_7506,N_7973);
nand U9076 (N_9076,N_6375,N_6042);
xnor U9077 (N_9077,N_7711,N_6284);
nand U9078 (N_9078,N_6807,N_6961);
or U9079 (N_9079,N_7856,N_6609);
nor U9080 (N_9080,N_7125,N_6000);
and U9081 (N_9081,N_7877,N_6111);
nor U9082 (N_9082,N_6836,N_7084);
nor U9083 (N_9083,N_6110,N_6937);
nand U9084 (N_9084,N_6567,N_6172);
or U9085 (N_9085,N_7073,N_7551);
or U9086 (N_9086,N_6746,N_6370);
nor U9087 (N_9087,N_6297,N_6473);
or U9088 (N_9088,N_7959,N_7567);
nor U9089 (N_9089,N_6669,N_7694);
or U9090 (N_9090,N_7877,N_6373);
nor U9091 (N_9091,N_6438,N_7797);
nor U9092 (N_9092,N_7342,N_6610);
nand U9093 (N_9093,N_6348,N_7855);
xnor U9094 (N_9094,N_6273,N_6267);
xor U9095 (N_9095,N_6551,N_7450);
nand U9096 (N_9096,N_7852,N_7351);
nand U9097 (N_9097,N_7247,N_7784);
xnor U9098 (N_9098,N_7769,N_7701);
nand U9099 (N_9099,N_6758,N_7285);
xnor U9100 (N_9100,N_6985,N_7624);
nand U9101 (N_9101,N_6431,N_7268);
or U9102 (N_9102,N_6700,N_7702);
and U9103 (N_9103,N_6246,N_6920);
xnor U9104 (N_9104,N_6839,N_7054);
xnor U9105 (N_9105,N_7952,N_7250);
nor U9106 (N_9106,N_6648,N_6662);
and U9107 (N_9107,N_7967,N_7953);
nor U9108 (N_9108,N_6194,N_6530);
nor U9109 (N_9109,N_7468,N_7363);
xor U9110 (N_9110,N_7925,N_6872);
and U9111 (N_9111,N_7514,N_6806);
nor U9112 (N_9112,N_7184,N_6748);
and U9113 (N_9113,N_7208,N_7906);
nand U9114 (N_9114,N_7673,N_6556);
nor U9115 (N_9115,N_6189,N_7843);
nor U9116 (N_9116,N_6622,N_6595);
nand U9117 (N_9117,N_7934,N_7178);
or U9118 (N_9118,N_7106,N_6138);
and U9119 (N_9119,N_6893,N_6056);
and U9120 (N_9120,N_6205,N_7852);
nand U9121 (N_9121,N_7351,N_6807);
nand U9122 (N_9122,N_7581,N_6455);
nand U9123 (N_9123,N_7444,N_7327);
and U9124 (N_9124,N_6545,N_7524);
or U9125 (N_9125,N_7813,N_7599);
nand U9126 (N_9126,N_7596,N_7378);
nand U9127 (N_9127,N_6596,N_7447);
nor U9128 (N_9128,N_7967,N_7386);
nand U9129 (N_9129,N_6176,N_6932);
nor U9130 (N_9130,N_7622,N_6360);
and U9131 (N_9131,N_6477,N_7174);
or U9132 (N_9132,N_7559,N_6725);
and U9133 (N_9133,N_6218,N_7842);
nor U9134 (N_9134,N_7241,N_7327);
or U9135 (N_9135,N_6156,N_7235);
and U9136 (N_9136,N_6679,N_6949);
nand U9137 (N_9137,N_7085,N_7542);
nor U9138 (N_9138,N_6100,N_6463);
or U9139 (N_9139,N_6512,N_7602);
nor U9140 (N_9140,N_7137,N_7031);
nor U9141 (N_9141,N_7843,N_6783);
nand U9142 (N_9142,N_7444,N_6975);
nand U9143 (N_9143,N_6766,N_7879);
or U9144 (N_9144,N_7606,N_6898);
or U9145 (N_9145,N_7944,N_6102);
and U9146 (N_9146,N_6215,N_7967);
nand U9147 (N_9147,N_7591,N_6280);
and U9148 (N_9148,N_6215,N_7442);
and U9149 (N_9149,N_7340,N_7597);
and U9150 (N_9150,N_7362,N_7509);
nor U9151 (N_9151,N_6885,N_6677);
nand U9152 (N_9152,N_7447,N_6212);
nor U9153 (N_9153,N_6873,N_6230);
and U9154 (N_9154,N_6811,N_7369);
or U9155 (N_9155,N_6931,N_6125);
and U9156 (N_9156,N_7721,N_7500);
nand U9157 (N_9157,N_7059,N_6485);
xor U9158 (N_9158,N_7448,N_6926);
or U9159 (N_9159,N_7284,N_6461);
nand U9160 (N_9160,N_7512,N_7672);
or U9161 (N_9161,N_7156,N_6568);
nand U9162 (N_9162,N_7780,N_6718);
or U9163 (N_9163,N_7062,N_7641);
nand U9164 (N_9164,N_7281,N_6953);
nand U9165 (N_9165,N_7893,N_7386);
and U9166 (N_9166,N_6618,N_7299);
nor U9167 (N_9167,N_7464,N_7256);
nor U9168 (N_9168,N_6694,N_7745);
xnor U9169 (N_9169,N_7977,N_7998);
xor U9170 (N_9170,N_6922,N_7287);
or U9171 (N_9171,N_7060,N_7105);
nor U9172 (N_9172,N_6150,N_7455);
nand U9173 (N_9173,N_6669,N_7535);
nand U9174 (N_9174,N_7565,N_7287);
nand U9175 (N_9175,N_6452,N_6666);
or U9176 (N_9176,N_7416,N_6889);
xnor U9177 (N_9177,N_7762,N_6492);
nor U9178 (N_9178,N_7138,N_7754);
xor U9179 (N_9179,N_7772,N_7785);
and U9180 (N_9180,N_7247,N_7118);
and U9181 (N_9181,N_7996,N_6386);
and U9182 (N_9182,N_7994,N_6954);
or U9183 (N_9183,N_7992,N_6076);
xnor U9184 (N_9184,N_6854,N_6412);
and U9185 (N_9185,N_6889,N_7480);
xnor U9186 (N_9186,N_7874,N_6512);
nand U9187 (N_9187,N_6440,N_7738);
nand U9188 (N_9188,N_6608,N_6172);
nand U9189 (N_9189,N_6120,N_7849);
nand U9190 (N_9190,N_6951,N_6002);
and U9191 (N_9191,N_7536,N_7790);
nand U9192 (N_9192,N_6469,N_7222);
and U9193 (N_9193,N_6763,N_6621);
or U9194 (N_9194,N_7948,N_7558);
and U9195 (N_9195,N_6164,N_7649);
nor U9196 (N_9196,N_6567,N_7626);
nand U9197 (N_9197,N_6004,N_6808);
or U9198 (N_9198,N_6498,N_7844);
or U9199 (N_9199,N_6962,N_6185);
or U9200 (N_9200,N_6190,N_7069);
xnor U9201 (N_9201,N_7886,N_6807);
or U9202 (N_9202,N_7843,N_6813);
or U9203 (N_9203,N_7213,N_7797);
nand U9204 (N_9204,N_6215,N_7928);
or U9205 (N_9205,N_6399,N_6652);
xor U9206 (N_9206,N_6909,N_6744);
or U9207 (N_9207,N_6158,N_7066);
xor U9208 (N_9208,N_6736,N_6708);
and U9209 (N_9209,N_6236,N_6800);
or U9210 (N_9210,N_6827,N_6534);
and U9211 (N_9211,N_6342,N_6391);
nor U9212 (N_9212,N_6284,N_7582);
and U9213 (N_9213,N_7517,N_7631);
nor U9214 (N_9214,N_6581,N_7357);
or U9215 (N_9215,N_6214,N_7564);
or U9216 (N_9216,N_7650,N_7644);
and U9217 (N_9217,N_7214,N_6788);
and U9218 (N_9218,N_7654,N_7162);
or U9219 (N_9219,N_6165,N_6347);
nor U9220 (N_9220,N_7428,N_7055);
nor U9221 (N_9221,N_6108,N_6962);
nor U9222 (N_9222,N_6342,N_6810);
and U9223 (N_9223,N_6523,N_7992);
nand U9224 (N_9224,N_6214,N_7185);
or U9225 (N_9225,N_6189,N_6457);
nand U9226 (N_9226,N_7624,N_7782);
nand U9227 (N_9227,N_7581,N_7914);
and U9228 (N_9228,N_6961,N_6247);
xor U9229 (N_9229,N_7003,N_6181);
nor U9230 (N_9230,N_6649,N_6282);
nand U9231 (N_9231,N_6203,N_7277);
or U9232 (N_9232,N_7708,N_6364);
xor U9233 (N_9233,N_7469,N_6748);
and U9234 (N_9234,N_6791,N_6181);
nand U9235 (N_9235,N_6965,N_7154);
or U9236 (N_9236,N_6024,N_6176);
nor U9237 (N_9237,N_7232,N_7709);
and U9238 (N_9238,N_6499,N_6582);
and U9239 (N_9239,N_7590,N_7796);
nor U9240 (N_9240,N_6053,N_7042);
and U9241 (N_9241,N_6253,N_7404);
xnor U9242 (N_9242,N_7423,N_7500);
nor U9243 (N_9243,N_6792,N_7310);
nor U9244 (N_9244,N_7952,N_7983);
nand U9245 (N_9245,N_6863,N_6443);
and U9246 (N_9246,N_7251,N_6910);
xnor U9247 (N_9247,N_6642,N_6162);
or U9248 (N_9248,N_6500,N_7007);
nor U9249 (N_9249,N_6043,N_7587);
nor U9250 (N_9250,N_6270,N_6098);
nor U9251 (N_9251,N_7341,N_7934);
xnor U9252 (N_9252,N_6902,N_6586);
and U9253 (N_9253,N_6377,N_7746);
nor U9254 (N_9254,N_6575,N_7841);
and U9255 (N_9255,N_7228,N_6334);
or U9256 (N_9256,N_6512,N_6638);
or U9257 (N_9257,N_7194,N_7886);
nor U9258 (N_9258,N_6502,N_7426);
nand U9259 (N_9259,N_7768,N_6149);
or U9260 (N_9260,N_7939,N_7843);
and U9261 (N_9261,N_7281,N_6268);
nand U9262 (N_9262,N_6698,N_7475);
or U9263 (N_9263,N_7759,N_7242);
or U9264 (N_9264,N_7893,N_7784);
and U9265 (N_9265,N_6302,N_7326);
nand U9266 (N_9266,N_6670,N_7405);
or U9267 (N_9267,N_6933,N_6238);
nor U9268 (N_9268,N_7892,N_7350);
xor U9269 (N_9269,N_6777,N_7592);
nor U9270 (N_9270,N_6284,N_7586);
or U9271 (N_9271,N_6211,N_7497);
nor U9272 (N_9272,N_6451,N_6730);
nor U9273 (N_9273,N_6972,N_7212);
nor U9274 (N_9274,N_7842,N_7386);
nand U9275 (N_9275,N_7421,N_7643);
or U9276 (N_9276,N_7153,N_7138);
nand U9277 (N_9277,N_6842,N_7662);
and U9278 (N_9278,N_6256,N_7269);
and U9279 (N_9279,N_7608,N_6979);
or U9280 (N_9280,N_7331,N_7120);
nor U9281 (N_9281,N_7268,N_6816);
and U9282 (N_9282,N_6754,N_7920);
nand U9283 (N_9283,N_6061,N_7561);
nand U9284 (N_9284,N_6784,N_6686);
or U9285 (N_9285,N_6251,N_6061);
and U9286 (N_9286,N_7189,N_7856);
and U9287 (N_9287,N_6477,N_6869);
or U9288 (N_9288,N_7497,N_7612);
and U9289 (N_9289,N_7871,N_6755);
nor U9290 (N_9290,N_7859,N_6076);
xnor U9291 (N_9291,N_6588,N_6571);
nor U9292 (N_9292,N_7868,N_6806);
and U9293 (N_9293,N_7685,N_7983);
nor U9294 (N_9294,N_7504,N_7170);
nor U9295 (N_9295,N_6858,N_6017);
nand U9296 (N_9296,N_7062,N_7818);
or U9297 (N_9297,N_6322,N_7318);
nand U9298 (N_9298,N_7633,N_7883);
nor U9299 (N_9299,N_6107,N_7719);
and U9300 (N_9300,N_7338,N_7453);
and U9301 (N_9301,N_7921,N_7935);
or U9302 (N_9302,N_6399,N_6486);
xor U9303 (N_9303,N_7251,N_6276);
and U9304 (N_9304,N_6013,N_6635);
and U9305 (N_9305,N_6979,N_6881);
nand U9306 (N_9306,N_7451,N_6063);
or U9307 (N_9307,N_7407,N_7171);
and U9308 (N_9308,N_7085,N_7114);
and U9309 (N_9309,N_6515,N_7562);
xnor U9310 (N_9310,N_6483,N_6272);
and U9311 (N_9311,N_7283,N_6436);
and U9312 (N_9312,N_6793,N_6160);
and U9313 (N_9313,N_6003,N_7638);
nand U9314 (N_9314,N_6487,N_6004);
and U9315 (N_9315,N_6064,N_6279);
and U9316 (N_9316,N_6452,N_6075);
and U9317 (N_9317,N_6743,N_6891);
nor U9318 (N_9318,N_7450,N_7694);
nand U9319 (N_9319,N_6660,N_7883);
and U9320 (N_9320,N_7175,N_7375);
nand U9321 (N_9321,N_6089,N_6505);
nand U9322 (N_9322,N_6209,N_7493);
nor U9323 (N_9323,N_7228,N_6356);
nor U9324 (N_9324,N_7061,N_7322);
and U9325 (N_9325,N_6554,N_6897);
nand U9326 (N_9326,N_7934,N_7413);
nor U9327 (N_9327,N_7615,N_6581);
nor U9328 (N_9328,N_7837,N_6343);
nor U9329 (N_9329,N_7658,N_6076);
nand U9330 (N_9330,N_6617,N_7395);
nor U9331 (N_9331,N_7820,N_7656);
or U9332 (N_9332,N_7952,N_7676);
nor U9333 (N_9333,N_6343,N_7834);
nand U9334 (N_9334,N_6225,N_7316);
nor U9335 (N_9335,N_7194,N_7005);
and U9336 (N_9336,N_6473,N_7599);
or U9337 (N_9337,N_7447,N_7504);
or U9338 (N_9338,N_7042,N_7394);
or U9339 (N_9339,N_7036,N_6270);
nand U9340 (N_9340,N_6787,N_7402);
nand U9341 (N_9341,N_6085,N_7907);
or U9342 (N_9342,N_6677,N_7296);
and U9343 (N_9343,N_7805,N_7603);
and U9344 (N_9344,N_7299,N_7912);
or U9345 (N_9345,N_6818,N_7094);
and U9346 (N_9346,N_6565,N_7817);
or U9347 (N_9347,N_7083,N_7653);
nor U9348 (N_9348,N_7919,N_7604);
nand U9349 (N_9349,N_6873,N_6483);
nand U9350 (N_9350,N_7521,N_7234);
nor U9351 (N_9351,N_7524,N_6217);
or U9352 (N_9352,N_6180,N_7745);
and U9353 (N_9353,N_6333,N_6567);
nor U9354 (N_9354,N_7992,N_7903);
nor U9355 (N_9355,N_6919,N_6851);
xnor U9356 (N_9356,N_6892,N_6071);
nand U9357 (N_9357,N_7712,N_6023);
nand U9358 (N_9358,N_6920,N_6458);
nand U9359 (N_9359,N_6659,N_7516);
and U9360 (N_9360,N_6457,N_6844);
or U9361 (N_9361,N_7696,N_7197);
nor U9362 (N_9362,N_7474,N_6021);
nor U9363 (N_9363,N_7423,N_6661);
nand U9364 (N_9364,N_6495,N_7411);
nand U9365 (N_9365,N_6050,N_6645);
xnor U9366 (N_9366,N_7021,N_7653);
nand U9367 (N_9367,N_6975,N_7537);
nand U9368 (N_9368,N_6499,N_7135);
and U9369 (N_9369,N_7732,N_7038);
or U9370 (N_9370,N_6748,N_6605);
xnor U9371 (N_9371,N_7707,N_7533);
and U9372 (N_9372,N_7733,N_7326);
or U9373 (N_9373,N_7205,N_7947);
nor U9374 (N_9374,N_7637,N_7527);
nor U9375 (N_9375,N_7624,N_7628);
or U9376 (N_9376,N_7089,N_6841);
xor U9377 (N_9377,N_6187,N_7626);
or U9378 (N_9378,N_7224,N_6337);
and U9379 (N_9379,N_7413,N_7788);
nand U9380 (N_9380,N_6586,N_6920);
nand U9381 (N_9381,N_6365,N_6217);
and U9382 (N_9382,N_7916,N_7572);
nor U9383 (N_9383,N_7064,N_7285);
nor U9384 (N_9384,N_6063,N_6217);
nand U9385 (N_9385,N_6245,N_6213);
nand U9386 (N_9386,N_6850,N_6270);
nand U9387 (N_9387,N_6160,N_6025);
nor U9388 (N_9388,N_6082,N_7032);
and U9389 (N_9389,N_7304,N_6257);
nand U9390 (N_9390,N_6842,N_7206);
nand U9391 (N_9391,N_7152,N_6068);
nand U9392 (N_9392,N_7941,N_6782);
or U9393 (N_9393,N_6499,N_7545);
nor U9394 (N_9394,N_6486,N_6697);
and U9395 (N_9395,N_6813,N_7994);
or U9396 (N_9396,N_6650,N_6792);
and U9397 (N_9397,N_7697,N_6237);
and U9398 (N_9398,N_6123,N_7797);
and U9399 (N_9399,N_6886,N_7104);
nor U9400 (N_9400,N_7467,N_6795);
nand U9401 (N_9401,N_6397,N_6402);
or U9402 (N_9402,N_6666,N_6945);
and U9403 (N_9403,N_6001,N_6280);
or U9404 (N_9404,N_7704,N_6949);
or U9405 (N_9405,N_6514,N_7594);
nand U9406 (N_9406,N_7525,N_6459);
and U9407 (N_9407,N_7969,N_7455);
or U9408 (N_9408,N_6641,N_7724);
xnor U9409 (N_9409,N_6820,N_6044);
nand U9410 (N_9410,N_6870,N_7333);
or U9411 (N_9411,N_7296,N_7794);
and U9412 (N_9412,N_7414,N_6765);
and U9413 (N_9413,N_6744,N_6179);
nand U9414 (N_9414,N_6148,N_6248);
or U9415 (N_9415,N_7963,N_7016);
nor U9416 (N_9416,N_7131,N_6929);
and U9417 (N_9417,N_6107,N_6158);
nand U9418 (N_9418,N_6238,N_6534);
or U9419 (N_9419,N_6910,N_6833);
nand U9420 (N_9420,N_6099,N_6385);
nor U9421 (N_9421,N_7591,N_7771);
nor U9422 (N_9422,N_6195,N_7740);
nand U9423 (N_9423,N_7484,N_6435);
or U9424 (N_9424,N_6116,N_6337);
nor U9425 (N_9425,N_6062,N_6192);
nor U9426 (N_9426,N_7953,N_7470);
nor U9427 (N_9427,N_7885,N_6745);
xnor U9428 (N_9428,N_7086,N_6231);
nor U9429 (N_9429,N_7672,N_7666);
nand U9430 (N_9430,N_6062,N_6462);
and U9431 (N_9431,N_6380,N_7107);
and U9432 (N_9432,N_7261,N_7855);
nand U9433 (N_9433,N_7205,N_6010);
nand U9434 (N_9434,N_6092,N_7775);
and U9435 (N_9435,N_6635,N_7083);
and U9436 (N_9436,N_7390,N_6742);
nor U9437 (N_9437,N_6980,N_6927);
and U9438 (N_9438,N_7023,N_7923);
or U9439 (N_9439,N_6376,N_6559);
nand U9440 (N_9440,N_7869,N_7053);
nand U9441 (N_9441,N_7352,N_7784);
nand U9442 (N_9442,N_6687,N_7010);
nor U9443 (N_9443,N_7631,N_7085);
or U9444 (N_9444,N_7314,N_7084);
nor U9445 (N_9445,N_6501,N_7389);
or U9446 (N_9446,N_7307,N_7741);
and U9447 (N_9447,N_7711,N_7626);
or U9448 (N_9448,N_7913,N_7336);
nand U9449 (N_9449,N_7895,N_6841);
and U9450 (N_9450,N_6071,N_6704);
nand U9451 (N_9451,N_7851,N_6299);
or U9452 (N_9452,N_7192,N_7616);
nand U9453 (N_9453,N_6920,N_7132);
or U9454 (N_9454,N_6867,N_6423);
nor U9455 (N_9455,N_7952,N_6339);
nand U9456 (N_9456,N_6077,N_6132);
or U9457 (N_9457,N_6160,N_6135);
nor U9458 (N_9458,N_6238,N_6758);
nor U9459 (N_9459,N_7752,N_6766);
or U9460 (N_9460,N_7203,N_6473);
or U9461 (N_9461,N_7676,N_7941);
nor U9462 (N_9462,N_6641,N_7230);
nor U9463 (N_9463,N_7375,N_7692);
or U9464 (N_9464,N_6562,N_6800);
nor U9465 (N_9465,N_7489,N_7949);
or U9466 (N_9466,N_7702,N_6998);
nor U9467 (N_9467,N_7338,N_7968);
nand U9468 (N_9468,N_7930,N_7789);
nor U9469 (N_9469,N_6869,N_6703);
or U9470 (N_9470,N_6854,N_7516);
nand U9471 (N_9471,N_7347,N_7920);
nor U9472 (N_9472,N_7086,N_7274);
nand U9473 (N_9473,N_7391,N_6560);
or U9474 (N_9474,N_7424,N_7175);
and U9475 (N_9475,N_6433,N_6611);
nand U9476 (N_9476,N_7738,N_7206);
and U9477 (N_9477,N_6503,N_7343);
xor U9478 (N_9478,N_7313,N_6014);
or U9479 (N_9479,N_6915,N_6630);
nand U9480 (N_9480,N_7555,N_7991);
nand U9481 (N_9481,N_7064,N_7423);
or U9482 (N_9482,N_6428,N_6078);
nor U9483 (N_9483,N_7393,N_7985);
and U9484 (N_9484,N_6967,N_7595);
or U9485 (N_9485,N_6694,N_7726);
nor U9486 (N_9486,N_7654,N_6012);
or U9487 (N_9487,N_7540,N_7745);
or U9488 (N_9488,N_7463,N_6050);
nand U9489 (N_9489,N_6924,N_7869);
or U9490 (N_9490,N_7590,N_7205);
and U9491 (N_9491,N_6716,N_6232);
xor U9492 (N_9492,N_6746,N_6683);
xnor U9493 (N_9493,N_7850,N_7434);
and U9494 (N_9494,N_7407,N_6962);
nand U9495 (N_9495,N_7259,N_6384);
nor U9496 (N_9496,N_6234,N_6412);
xor U9497 (N_9497,N_7240,N_6857);
nor U9498 (N_9498,N_6478,N_6608);
and U9499 (N_9499,N_7503,N_7733);
nor U9500 (N_9500,N_6892,N_6869);
nand U9501 (N_9501,N_7757,N_7983);
and U9502 (N_9502,N_6206,N_6476);
nor U9503 (N_9503,N_7256,N_7303);
xor U9504 (N_9504,N_7319,N_6299);
and U9505 (N_9505,N_6241,N_7334);
xnor U9506 (N_9506,N_6002,N_6388);
nand U9507 (N_9507,N_7448,N_6537);
nand U9508 (N_9508,N_7706,N_7070);
and U9509 (N_9509,N_6759,N_7984);
and U9510 (N_9510,N_7115,N_7272);
and U9511 (N_9511,N_6812,N_6727);
nor U9512 (N_9512,N_6662,N_7133);
nor U9513 (N_9513,N_7120,N_7713);
or U9514 (N_9514,N_6656,N_6338);
nor U9515 (N_9515,N_7355,N_6174);
nand U9516 (N_9516,N_6013,N_7390);
nor U9517 (N_9517,N_6825,N_7607);
nand U9518 (N_9518,N_7205,N_7868);
nor U9519 (N_9519,N_7990,N_7835);
nor U9520 (N_9520,N_7926,N_7500);
nand U9521 (N_9521,N_6678,N_6661);
nand U9522 (N_9522,N_7797,N_7464);
nand U9523 (N_9523,N_7578,N_7355);
xnor U9524 (N_9524,N_7605,N_7121);
and U9525 (N_9525,N_6270,N_6147);
or U9526 (N_9526,N_6448,N_6879);
nand U9527 (N_9527,N_7256,N_6025);
nor U9528 (N_9528,N_7483,N_7612);
xor U9529 (N_9529,N_6694,N_7938);
nand U9530 (N_9530,N_7071,N_6005);
and U9531 (N_9531,N_6692,N_7226);
and U9532 (N_9532,N_7320,N_7605);
or U9533 (N_9533,N_6608,N_6906);
nor U9534 (N_9534,N_6291,N_7377);
and U9535 (N_9535,N_7813,N_7066);
nor U9536 (N_9536,N_6296,N_6993);
and U9537 (N_9537,N_6185,N_7611);
nand U9538 (N_9538,N_7472,N_7568);
or U9539 (N_9539,N_6883,N_6875);
nand U9540 (N_9540,N_6279,N_7105);
nand U9541 (N_9541,N_6953,N_6124);
and U9542 (N_9542,N_6209,N_7821);
and U9543 (N_9543,N_6945,N_7231);
or U9544 (N_9544,N_6283,N_6690);
nand U9545 (N_9545,N_6589,N_7265);
or U9546 (N_9546,N_7445,N_7671);
nand U9547 (N_9547,N_7510,N_7420);
and U9548 (N_9548,N_7158,N_7665);
and U9549 (N_9549,N_7060,N_7628);
nor U9550 (N_9550,N_7379,N_6414);
and U9551 (N_9551,N_7578,N_7761);
and U9552 (N_9552,N_6748,N_7854);
xor U9553 (N_9553,N_7896,N_7119);
nand U9554 (N_9554,N_6108,N_6223);
nor U9555 (N_9555,N_7645,N_6025);
nor U9556 (N_9556,N_6572,N_6073);
or U9557 (N_9557,N_6749,N_7967);
nand U9558 (N_9558,N_6156,N_7309);
nand U9559 (N_9559,N_6742,N_6687);
and U9560 (N_9560,N_6319,N_6926);
and U9561 (N_9561,N_7973,N_6520);
and U9562 (N_9562,N_7053,N_6577);
nor U9563 (N_9563,N_7757,N_6237);
or U9564 (N_9564,N_6671,N_6299);
or U9565 (N_9565,N_6711,N_6528);
nand U9566 (N_9566,N_7392,N_7123);
xnor U9567 (N_9567,N_7719,N_6619);
nor U9568 (N_9568,N_6217,N_6985);
or U9569 (N_9569,N_7129,N_6741);
nor U9570 (N_9570,N_7012,N_7339);
nor U9571 (N_9571,N_6770,N_7267);
nand U9572 (N_9572,N_7163,N_6222);
nor U9573 (N_9573,N_6342,N_6302);
nor U9574 (N_9574,N_7409,N_7290);
nor U9575 (N_9575,N_7304,N_6463);
or U9576 (N_9576,N_6912,N_6301);
xnor U9577 (N_9577,N_6927,N_6623);
and U9578 (N_9578,N_7147,N_7685);
xnor U9579 (N_9579,N_6051,N_7978);
xnor U9580 (N_9580,N_6409,N_7502);
or U9581 (N_9581,N_7920,N_6256);
nor U9582 (N_9582,N_6820,N_7438);
and U9583 (N_9583,N_6128,N_7010);
nand U9584 (N_9584,N_7911,N_7202);
or U9585 (N_9585,N_7018,N_6831);
nor U9586 (N_9586,N_7624,N_7755);
and U9587 (N_9587,N_7295,N_6481);
nand U9588 (N_9588,N_7889,N_7075);
or U9589 (N_9589,N_6298,N_7351);
or U9590 (N_9590,N_6830,N_7815);
and U9591 (N_9591,N_7744,N_6336);
nor U9592 (N_9592,N_6180,N_7715);
or U9593 (N_9593,N_7548,N_7833);
nand U9594 (N_9594,N_6145,N_6425);
nor U9595 (N_9595,N_6031,N_6257);
nor U9596 (N_9596,N_7275,N_7804);
and U9597 (N_9597,N_7561,N_6908);
and U9598 (N_9598,N_6963,N_7905);
and U9599 (N_9599,N_6924,N_6656);
nor U9600 (N_9600,N_7642,N_6798);
nor U9601 (N_9601,N_7505,N_6678);
nor U9602 (N_9602,N_6674,N_6594);
nor U9603 (N_9603,N_6030,N_6914);
and U9604 (N_9604,N_6725,N_7306);
and U9605 (N_9605,N_6849,N_7056);
or U9606 (N_9606,N_7688,N_7677);
nand U9607 (N_9607,N_7235,N_7574);
xor U9608 (N_9608,N_6099,N_6072);
nor U9609 (N_9609,N_7845,N_6071);
and U9610 (N_9610,N_7193,N_7272);
xor U9611 (N_9611,N_6095,N_6716);
and U9612 (N_9612,N_6579,N_7571);
or U9613 (N_9613,N_7866,N_7449);
xnor U9614 (N_9614,N_7578,N_6408);
nand U9615 (N_9615,N_7339,N_6163);
nand U9616 (N_9616,N_6606,N_6779);
or U9617 (N_9617,N_7518,N_6942);
nor U9618 (N_9618,N_7612,N_6793);
xnor U9619 (N_9619,N_7389,N_6293);
or U9620 (N_9620,N_7099,N_7121);
and U9621 (N_9621,N_7497,N_7026);
nand U9622 (N_9622,N_6370,N_6055);
or U9623 (N_9623,N_7313,N_6777);
or U9624 (N_9624,N_6445,N_6419);
or U9625 (N_9625,N_7060,N_6853);
nor U9626 (N_9626,N_7868,N_7915);
and U9627 (N_9627,N_6383,N_6437);
nor U9628 (N_9628,N_7361,N_6119);
and U9629 (N_9629,N_7687,N_6829);
or U9630 (N_9630,N_6102,N_6707);
nand U9631 (N_9631,N_6643,N_7814);
or U9632 (N_9632,N_7432,N_7848);
xor U9633 (N_9633,N_7645,N_7401);
and U9634 (N_9634,N_6881,N_7590);
nor U9635 (N_9635,N_6641,N_6229);
nor U9636 (N_9636,N_7637,N_6573);
or U9637 (N_9637,N_6878,N_7378);
nor U9638 (N_9638,N_7995,N_7817);
or U9639 (N_9639,N_7006,N_6839);
or U9640 (N_9640,N_6425,N_6174);
xnor U9641 (N_9641,N_7198,N_7329);
and U9642 (N_9642,N_7114,N_7340);
nand U9643 (N_9643,N_7214,N_6722);
nor U9644 (N_9644,N_7309,N_7630);
or U9645 (N_9645,N_6776,N_6484);
nand U9646 (N_9646,N_6476,N_7977);
nand U9647 (N_9647,N_7891,N_7068);
nor U9648 (N_9648,N_7261,N_7223);
or U9649 (N_9649,N_7420,N_7551);
and U9650 (N_9650,N_7626,N_6048);
and U9651 (N_9651,N_7316,N_7927);
or U9652 (N_9652,N_7183,N_6599);
and U9653 (N_9653,N_7278,N_6661);
or U9654 (N_9654,N_6011,N_6954);
xnor U9655 (N_9655,N_7181,N_6971);
and U9656 (N_9656,N_7331,N_6945);
nor U9657 (N_9657,N_7078,N_7085);
nor U9658 (N_9658,N_6269,N_7829);
xor U9659 (N_9659,N_6831,N_7632);
nor U9660 (N_9660,N_7680,N_6661);
or U9661 (N_9661,N_7182,N_7380);
or U9662 (N_9662,N_7338,N_7643);
and U9663 (N_9663,N_6845,N_7254);
or U9664 (N_9664,N_7391,N_6532);
nand U9665 (N_9665,N_6296,N_7407);
xnor U9666 (N_9666,N_6964,N_6118);
and U9667 (N_9667,N_6564,N_6489);
and U9668 (N_9668,N_6921,N_6380);
nor U9669 (N_9669,N_6772,N_7815);
nand U9670 (N_9670,N_7185,N_7030);
nand U9671 (N_9671,N_7931,N_6715);
and U9672 (N_9672,N_6245,N_6352);
xor U9673 (N_9673,N_7644,N_6737);
nor U9674 (N_9674,N_6124,N_7636);
xnor U9675 (N_9675,N_7148,N_7184);
nand U9676 (N_9676,N_6059,N_7017);
nand U9677 (N_9677,N_7300,N_6918);
and U9678 (N_9678,N_6352,N_6896);
nor U9679 (N_9679,N_6034,N_7544);
or U9680 (N_9680,N_7850,N_7069);
or U9681 (N_9681,N_7448,N_7095);
or U9682 (N_9682,N_6247,N_6919);
or U9683 (N_9683,N_6761,N_7633);
or U9684 (N_9684,N_6567,N_7265);
nor U9685 (N_9685,N_7331,N_7351);
or U9686 (N_9686,N_7682,N_6027);
nand U9687 (N_9687,N_7917,N_7444);
nor U9688 (N_9688,N_6745,N_7656);
nand U9689 (N_9689,N_6326,N_7153);
nand U9690 (N_9690,N_6093,N_7792);
or U9691 (N_9691,N_6568,N_6192);
nor U9692 (N_9692,N_7642,N_6932);
nor U9693 (N_9693,N_6557,N_6331);
nand U9694 (N_9694,N_6974,N_6283);
nand U9695 (N_9695,N_6588,N_7480);
xnor U9696 (N_9696,N_7926,N_6177);
xnor U9697 (N_9697,N_7984,N_7061);
xor U9698 (N_9698,N_7497,N_7303);
and U9699 (N_9699,N_6302,N_7220);
or U9700 (N_9700,N_7048,N_6205);
nand U9701 (N_9701,N_7799,N_7148);
xnor U9702 (N_9702,N_7202,N_6654);
and U9703 (N_9703,N_6248,N_6225);
and U9704 (N_9704,N_7326,N_7910);
xor U9705 (N_9705,N_7095,N_7292);
and U9706 (N_9706,N_6161,N_6660);
or U9707 (N_9707,N_7036,N_6935);
nor U9708 (N_9708,N_7674,N_6192);
nor U9709 (N_9709,N_6565,N_7399);
or U9710 (N_9710,N_7493,N_6367);
and U9711 (N_9711,N_7037,N_7315);
or U9712 (N_9712,N_6414,N_7313);
nand U9713 (N_9713,N_7435,N_7387);
or U9714 (N_9714,N_6550,N_7443);
and U9715 (N_9715,N_6178,N_6866);
xnor U9716 (N_9716,N_6772,N_7933);
nand U9717 (N_9717,N_6229,N_6852);
nand U9718 (N_9718,N_7820,N_6275);
nand U9719 (N_9719,N_6163,N_6337);
xor U9720 (N_9720,N_6690,N_7330);
xor U9721 (N_9721,N_6731,N_7164);
xnor U9722 (N_9722,N_6949,N_7612);
nor U9723 (N_9723,N_6309,N_7430);
or U9724 (N_9724,N_7751,N_7827);
nand U9725 (N_9725,N_6928,N_7946);
or U9726 (N_9726,N_7556,N_6692);
or U9727 (N_9727,N_6477,N_7352);
xnor U9728 (N_9728,N_6846,N_7158);
and U9729 (N_9729,N_7855,N_6231);
and U9730 (N_9730,N_6995,N_7950);
nand U9731 (N_9731,N_6217,N_7253);
or U9732 (N_9732,N_7372,N_6322);
or U9733 (N_9733,N_7914,N_7639);
nand U9734 (N_9734,N_6475,N_7725);
nor U9735 (N_9735,N_6201,N_7017);
nor U9736 (N_9736,N_6589,N_7202);
and U9737 (N_9737,N_6941,N_7134);
and U9738 (N_9738,N_6334,N_6475);
and U9739 (N_9739,N_7209,N_7868);
nor U9740 (N_9740,N_6732,N_7259);
and U9741 (N_9741,N_6223,N_7989);
and U9742 (N_9742,N_7248,N_7851);
or U9743 (N_9743,N_6566,N_6604);
nor U9744 (N_9744,N_6630,N_7164);
xor U9745 (N_9745,N_6812,N_7998);
xnor U9746 (N_9746,N_6462,N_7496);
and U9747 (N_9747,N_6255,N_7370);
nor U9748 (N_9748,N_7599,N_6677);
xor U9749 (N_9749,N_7126,N_7006);
nor U9750 (N_9750,N_6065,N_7684);
and U9751 (N_9751,N_6304,N_7364);
or U9752 (N_9752,N_6899,N_7944);
or U9753 (N_9753,N_6282,N_6343);
nor U9754 (N_9754,N_7946,N_7481);
and U9755 (N_9755,N_6261,N_6477);
or U9756 (N_9756,N_7211,N_7789);
nor U9757 (N_9757,N_7440,N_7966);
or U9758 (N_9758,N_7122,N_7034);
nand U9759 (N_9759,N_7166,N_6374);
nand U9760 (N_9760,N_7542,N_7571);
and U9761 (N_9761,N_7247,N_6061);
or U9762 (N_9762,N_7790,N_7848);
or U9763 (N_9763,N_7188,N_7806);
and U9764 (N_9764,N_7313,N_6855);
nor U9765 (N_9765,N_6065,N_6007);
and U9766 (N_9766,N_6608,N_6274);
nand U9767 (N_9767,N_7410,N_6300);
xnor U9768 (N_9768,N_6765,N_7132);
and U9769 (N_9769,N_7560,N_6844);
nor U9770 (N_9770,N_7749,N_6629);
nor U9771 (N_9771,N_6110,N_7045);
nor U9772 (N_9772,N_7853,N_7642);
nor U9773 (N_9773,N_7937,N_6293);
or U9774 (N_9774,N_7566,N_6377);
and U9775 (N_9775,N_7505,N_6408);
or U9776 (N_9776,N_7208,N_6225);
nand U9777 (N_9777,N_6930,N_6223);
nand U9778 (N_9778,N_6794,N_7672);
nor U9779 (N_9779,N_7858,N_6677);
xor U9780 (N_9780,N_7433,N_7934);
nor U9781 (N_9781,N_6619,N_6020);
and U9782 (N_9782,N_6073,N_6224);
or U9783 (N_9783,N_7768,N_7243);
and U9784 (N_9784,N_7804,N_6806);
or U9785 (N_9785,N_6715,N_6879);
nor U9786 (N_9786,N_6660,N_6506);
nor U9787 (N_9787,N_7156,N_6756);
or U9788 (N_9788,N_7653,N_6378);
nor U9789 (N_9789,N_6004,N_7951);
and U9790 (N_9790,N_7129,N_7434);
nand U9791 (N_9791,N_6055,N_7250);
xor U9792 (N_9792,N_6351,N_7079);
and U9793 (N_9793,N_6792,N_7962);
and U9794 (N_9794,N_6959,N_6976);
nor U9795 (N_9795,N_6100,N_7267);
nor U9796 (N_9796,N_6863,N_6597);
nand U9797 (N_9797,N_7769,N_6408);
xnor U9798 (N_9798,N_7322,N_6277);
nor U9799 (N_9799,N_6543,N_6710);
or U9800 (N_9800,N_7573,N_7612);
and U9801 (N_9801,N_7051,N_7094);
or U9802 (N_9802,N_7235,N_6362);
nand U9803 (N_9803,N_7935,N_7243);
or U9804 (N_9804,N_7889,N_7203);
or U9805 (N_9805,N_7811,N_7299);
or U9806 (N_9806,N_7016,N_6359);
and U9807 (N_9807,N_6728,N_6949);
or U9808 (N_9808,N_7399,N_6439);
xor U9809 (N_9809,N_6889,N_7077);
nor U9810 (N_9810,N_7305,N_7167);
and U9811 (N_9811,N_7252,N_6359);
nand U9812 (N_9812,N_6146,N_7612);
nand U9813 (N_9813,N_7318,N_7301);
nor U9814 (N_9814,N_6975,N_6293);
or U9815 (N_9815,N_6488,N_6402);
or U9816 (N_9816,N_7132,N_7135);
nand U9817 (N_9817,N_7437,N_7673);
or U9818 (N_9818,N_7520,N_6118);
nand U9819 (N_9819,N_7288,N_6351);
nor U9820 (N_9820,N_6403,N_6981);
or U9821 (N_9821,N_6830,N_6690);
nand U9822 (N_9822,N_6494,N_7903);
nand U9823 (N_9823,N_6655,N_7786);
nor U9824 (N_9824,N_6117,N_7050);
nor U9825 (N_9825,N_6785,N_7535);
nand U9826 (N_9826,N_6849,N_6657);
and U9827 (N_9827,N_7173,N_6542);
nor U9828 (N_9828,N_6464,N_6118);
nand U9829 (N_9829,N_7176,N_7606);
and U9830 (N_9830,N_6120,N_7655);
and U9831 (N_9831,N_7889,N_7988);
and U9832 (N_9832,N_7773,N_7158);
and U9833 (N_9833,N_7103,N_7143);
nand U9834 (N_9834,N_6172,N_7364);
nand U9835 (N_9835,N_6101,N_6944);
and U9836 (N_9836,N_7697,N_7765);
or U9837 (N_9837,N_6400,N_6159);
or U9838 (N_9838,N_7187,N_7769);
or U9839 (N_9839,N_6180,N_6506);
nor U9840 (N_9840,N_7829,N_7909);
nand U9841 (N_9841,N_7329,N_7417);
nand U9842 (N_9842,N_7092,N_6843);
nor U9843 (N_9843,N_7243,N_7748);
nand U9844 (N_9844,N_7903,N_7107);
nor U9845 (N_9845,N_6590,N_7772);
nor U9846 (N_9846,N_6712,N_6197);
nor U9847 (N_9847,N_7233,N_7514);
or U9848 (N_9848,N_6490,N_7433);
nand U9849 (N_9849,N_6806,N_7734);
nor U9850 (N_9850,N_7092,N_6192);
and U9851 (N_9851,N_7627,N_6927);
nor U9852 (N_9852,N_6176,N_6468);
nand U9853 (N_9853,N_6941,N_7917);
and U9854 (N_9854,N_7221,N_7382);
or U9855 (N_9855,N_6547,N_6103);
and U9856 (N_9856,N_7725,N_7275);
nand U9857 (N_9857,N_7217,N_7336);
nor U9858 (N_9858,N_7903,N_6045);
or U9859 (N_9859,N_6434,N_7113);
xnor U9860 (N_9860,N_6995,N_6504);
nor U9861 (N_9861,N_7204,N_6723);
nand U9862 (N_9862,N_6077,N_6905);
nor U9863 (N_9863,N_7663,N_7102);
nand U9864 (N_9864,N_7984,N_7315);
and U9865 (N_9865,N_7404,N_6735);
nor U9866 (N_9866,N_7839,N_7546);
xor U9867 (N_9867,N_7343,N_6487);
nor U9868 (N_9868,N_6330,N_7516);
or U9869 (N_9869,N_6510,N_6040);
or U9870 (N_9870,N_7391,N_7196);
and U9871 (N_9871,N_7591,N_6800);
nor U9872 (N_9872,N_6299,N_7524);
nand U9873 (N_9873,N_6321,N_7549);
nor U9874 (N_9874,N_7356,N_7218);
nand U9875 (N_9875,N_6731,N_7945);
nand U9876 (N_9876,N_6363,N_6513);
nor U9877 (N_9877,N_7343,N_6623);
or U9878 (N_9878,N_6851,N_6596);
and U9879 (N_9879,N_6416,N_7839);
and U9880 (N_9880,N_7683,N_7309);
and U9881 (N_9881,N_6523,N_7090);
nor U9882 (N_9882,N_6189,N_6145);
and U9883 (N_9883,N_6093,N_7303);
and U9884 (N_9884,N_7093,N_6102);
and U9885 (N_9885,N_7865,N_6105);
nor U9886 (N_9886,N_6024,N_7139);
or U9887 (N_9887,N_7480,N_7765);
nand U9888 (N_9888,N_7351,N_6334);
nand U9889 (N_9889,N_6548,N_7918);
and U9890 (N_9890,N_6561,N_7844);
xnor U9891 (N_9891,N_7416,N_6896);
nor U9892 (N_9892,N_6319,N_6343);
or U9893 (N_9893,N_6508,N_6942);
and U9894 (N_9894,N_7516,N_7130);
nor U9895 (N_9895,N_7530,N_6932);
nor U9896 (N_9896,N_6571,N_6395);
and U9897 (N_9897,N_7191,N_6143);
nand U9898 (N_9898,N_6201,N_6279);
or U9899 (N_9899,N_7275,N_7108);
and U9900 (N_9900,N_6048,N_7522);
nand U9901 (N_9901,N_7555,N_6259);
nor U9902 (N_9902,N_7172,N_7551);
xnor U9903 (N_9903,N_6242,N_6442);
and U9904 (N_9904,N_7144,N_6975);
nor U9905 (N_9905,N_7660,N_6638);
nor U9906 (N_9906,N_7214,N_7483);
nand U9907 (N_9907,N_6045,N_6973);
and U9908 (N_9908,N_6254,N_7580);
nor U9909 (N_9909,N_6420,N_6435);
nor U9910 (N_9910,N_6149,N_6486);
nand U9911 (N_9911,N_6534,N_6090);
xnor U9912 (N_9912,N_6193,N_6305);
nor U9913 (N_9913,N_6709,N_7315);
nor U9914 (N_9914,N_7541,N_6473);
or U9915 (N_9915,N_6435,N_7522);
nand U9916 (N_9916,N_6395,N_7851);
and U9917 (N_9917,N_6490,N_6700);
nor U9918 (N_9918,N_6931,N_7755);
nor U9919 (N_9919,N_7584,N_6110);
nand U9920 (N_9920,N_7237,N_6233);
xor U9921 (N_9921,N_6740,N_7792);
nor U9922 (N_9922,N_6159,N_7274);
and U9923 (N_9923,N_7475,N_6491);
nor U9924 (N_9924,N_6584,N_7997);
and U9925 (N_9925,N_6862,N_6335);
nand U9926 (N_9926,N_6732,N_6937);
nand U9927 (N_9927,N_6982,N_6338);
and U9928 (N_9928,N_6384,N_6483);
and U9929 (N_9929,N_6536,N_6109);
or U9930 (N_9930,N_6710,N_6821);
nor U9931 (N_9931,N_7252,N_7146);
nor U9932 (N_9932,N_7360,N_7387);
or U9933 (N_9933,N_6686,N_6608);
and U9934 (N_9934,N_7085,N_6653);
xor U9935 (N_9935,N_6020,N_7206);
or U9936 (N_9936,N_7382,N_7406);
and U9937 (N_9937,N_7167,N_6455);
and U9938 (N_9938,N_6896,N_6035);
nand U9939 (N_9939,N_7653,N_7581);
nor U9940 (N_9940,N_7037,N_6018);
nand U9941 (N_9941,N_6583,N_6143);
xnor U9942 (N_9942,N_6941,N_6467);
xor U9943 (N_9943,N_6939,N_6100);
nand U9944 (N_9944,N_7695,N_6197);
and U9945 (N_9945,N_6419,N_7382);
nand U9946 (N_9946,N_6138,N_7051);
or U9947 (N_9947,N_7756,N_7301);
or U9948 (N_9948,N_7813,N_6571);
nand U9949 (N_9949,N_6426,N_6000);
and U9950 (N_9950,N_6083,N_6680);
or U9951 (N_9951,N_6994,N_6300);
nand U9952 (N_9952,N_6861,N_6715);
or U9953 (N_9953,N_6129,N_6963);
and U9954 (N_9954,N_7124,N_7958);
xnor U9955 (N_9955,N_6017,N_7434);
nand U9956 (N_9956,N_6780,N_7080);
nor U9957 (N_9957,N_7021,N_7562);
nor U9958 (N_9958,N_6238,N_7014);
and U9959 (N_9959,N_6536,N_7596);
nand U9960 (N_9960,N_7639,N_7276);
nand U9961 (N_9961,N_7554,N_6699);
xnor U9962 (N_9962,N_6177,N_7575);
nor U9963 (N_9963,N_7458,N_6578);
nand U9964 (N_9964,N_7711,N_7024);
xnor U9965 (N_9965,N_7897,N_6048);
nor U9966 (N_9966,N_6570,N_6566);
or U9967 (N_9967,N_7719,N_6964);
nand U9968 (N_9968,N_6688,N_6174);
nor U9969 (N_9969,N_6518,N_6210);
and U9970 (N_9970,N_6264,N_6718);
nor U9971 (N_9971,N_6707,N_6572);
xor U9972 (N_9972,N_6507,N_7740);
nor U9973 (N_9973,N_7422,N_6822);
nor U9974 (N_9974,N_7225,N_6408);
and U9975 (N_9975,N_7651,N_6647);
nand U9976 (N_9976,N_7006,N_7691);
nand U9977 (N_9977,N_6132,N_7122);
or U9978 (N_9978,N_7886,N_6770);
and U9979 (N_9979,N_7250,N_6843);
or U9980 (N_9980,N_7984,N_7998);
nor U9981 (N_9981,N_7761,N_7323);
and U9982 (N_9982,N_7264,N_7436);
and U9983 (N_9983,N_6596,N_7357);
nand U9984 (N_9984,N_6667,N_6853);
xnor U9985 (N_9985,N_7843,N_7856);
and U9986 (N_9986,N_7381,N_6323);
or U9987 (N_9987,N_7006,N_6815);
nand U9988 (N_9988,N_6893,N_7630);
or U9989 (N_9989,N_7138,N_6454);
nor U9990 (N_9990,N_7438,N_6037);
and U9991 (N_9991,N_7768,N_6761);
or U9992 (N_9992,N_6952,N_7000);
nand U9993 (N_9993,N_7227,N_6304);
nor U9994 (N_9994,N_6527,N_7535);
nor U9995 (N_9995,N_7199,N_7260);
nor U9996 (N_9996,N_6557,N_7427);
or U9997 (N_9997,N_6147,N_7781);
or U9998 (N_9998,N_7517,N_6835);
or U9999 (N_9999,N_6000,N_6950);
and UO_0 (O_0,N_9004,N_8268);
nand UO_1 (O_1,N_8596,N_9808);
nand UO_2 (O_2,N_9500,N_8141);
or UO_3 (O_3,N_8790,N_8104);
and UO_4 (O_4,N_9086,N_9692);
and UO_5 (O_5,N_8575,N_8623);
nand UO_6 (O_6,N_8282,N_9947);
or UO_7 (O_7,N_9543,N_9851);
nand UO_8 (O_8,N_9852,N_9108);
or UO_9 (O_9,N_9363,N_8209);
nor UO_10 (O_10,N_8186,N_9073);
nand UO_11 (O_11,N_9617,N_8284);
or UO_12 (O_12,N_8181,N_9737);
and UO_13 (O_13,N_9044,N_8749);
nor UO_14 (O_14,N_9504,N_8479);
or UO_15 (O_15,N_9857,N_9270);
and UO_16 (O_16,N_8836,N_9919);
nor UO_17 (O_17,N_8890,N_9755);
and UO_18 (O_18,N_9869,N_8056);
nand UO_19 (O_19,N_9656,N_8151);
and UO_20 (O_20,N_8738,N_8292);
nor UO_21 (O_21,N_9630,N_9439);
and UO_22 (O_22,N_8614,N_9578);
or UO_23 (O_23,N_9182,N_9315);
nor UO_24 (O_24,N_8742,N_9918);
nand UO_25 (O_25,N_9462,N_9001);
and UO_26 (O_26,N_8079,N_8083);
nand UO_27 (O_27,N_8859,N_8605);
nand UO_28 (O_28,N_9832,N_9533);
and UO_29 (O_29,N_9139,N_8378);
nand UO_30 (O_30,N_9340,N_9822);
and UO_31 (O_31,N_9140,N_8293);
nor UO_32 (O_32,N_9989,N_8386);
or UO_33 (O_33,N_9227,N_8794);
and UO_34 (O_34,N_8529,N_8886);
nor UO_35 (O_35,N_9278,N_8059);
and UO_36 (O_36,N_8204,N_8536);
nand UO_37 (O_37,N_8789,N_8939);
and UO_38 (O_38,N_9289,N_9901);
nand UO_39 (O_39,N_9017,N_8152);
and UO_40 (O_40,N_9539,N_8361);
nor UO_41 (O_41,N_8571,N_8868);
and UO_42 (O_42,N_9749,N_8923);
nor UO_43 (O_43,N_8520,N_8804);
and UO_44 (O_44,N_9951,N_9896);
xnor UO_45 (O_45,N_9770,N_8046);
nand UO_46 (O_46,N_8356,N_8107);
and UO_47 (O_47,N_9676,N_8705);
and UO_48 (O_48,N_9193,N_8611);
and UO_49 (O_49,N_9373,N_8171);
or UO_50 (O_50,N_9341,N_9029);
nand UO_51 (O_51,N_8864,N_8467);
nor UO_52 (O_52,N_9293,N_8768);
xor UO_53 (O_53,N_9837,N_9326);
and UO_54 (O_54,N_8678,N_8475);
nor UO_55 (O_55,N_9476,N_8949);
nand UO_56 (O_56,N_9332,N_8134);
nor UO_57 (O_57,N_8600,N_9246);
and UO_58 (O_58,N_8887,N_8343);
nand UO_59 (O_59,N_9413,N_8711);
nand UO_60 (O_60,N_9350,N_9575);
nor UO_61 (O_61,N_8621,N_9337);
nor UO_62 (O_62,N_8556,N_8454);
xor UO_63 (O_63,N_9746,N_8979);
nand UO_64 (O_64,N_9936,N_9667);
nand UO_65 (O_65,N_8910,N_9817);
and UO_66 (O_66,N_9074,N_8359);
or UO_67 (O_67,N_9060,N_9813);
xnor UO_68 (O_68,N_9566,N_8233);
or UO_69 (O_69,N_9727,N_8207);
and UO_70 (O_70,N_8324,N_8000);
nor UO_71 (O_71,N_9381,N_8875);
nand UO_72 (O_72,N_8068,N_8512);
and UO_73 (O_73,N_8214,N_9957);
or UO_74 (O_74,N_8136,N_8116);
or UO_75 (O_75,N_8322,N_8052);
nand UO_76 (O_76,N_8763,N_9952);
nor UO_77 (O_77,N_8954,N_9306);
nand UO_78 (O_78,N_9626,N_8930);
xor UO_79 (O_79,N_8936,N_9716);
and UO_80 (O_80,N_8929,N_9873);
nand UO_81 (O_81,N_8096,N_8674);
nor UO_82 (O_82,N_9101,N_8710);
or UO_83 (O_83,N_8246,N_9999);
nand UO_84 (O_84,N_9591,N_8993);
nand UO_85 (O_85,N_9927,N_9829);
or UO_86 (O_86,N_9760,N_8249);
and UO_87 (O_87,N_9549,N_8992);
nor UO_88 (O_88,N_8762,N_9427);
nand UO_89 (O_89,N_9112,N_8021);
xor UO_90 (O_90,N_9625,N_8848);
nand UO_91 (O_91,N_9877,N_8053);
and UO_92 (O_92,N_9607,N_8419);
xor UO_93 (O_93,N_8702,N_9600);
and UO_94 (O_94,N_9091,N_8659);
and UO_95 (O_95,N_8121,N_8591);
nand UO_96 (O_96,N_8128,N_8631);
nor UO_97 (O_97,N_9898,N_8552);
and UO_98 (O_98,N_8244,N_9369);
nor UO_99 (O_99,N_9364,N_8224);
nor UO_100 (O_100,N_9592,N_8471);
xnor UO_101 (O_101,N_8839,N_9700);
nand UO_102 (O_102,N_8477,N_8100);
and UO_103 (O_103,N_9587,N_8443);
nand UO_104 (O_104,N_9062,N_9257);
and UO_105 (O_105,N_8216,N_8953);
or UO_106 (O_106,N_9166,N_9122);
or UO_107 (O_107,N_8852,N_8904);
or UO_108 (O_108,N_8031,N_9342);
and UO_109 (O_109,N_8810,N_8997);
and UO_110 (O_110,N_9641,N_8262);
or UO_111 (O_111,N_9775,N_9406);
nor UO_112 (O_112,N_8338,N_8905);
or UO_113 (O_113,N_9691,N_9374);
nor UO_114 (O_114,N_9432,N_9102);
xor UO_115 (O_115,N_8668,N_9594);
nor UO_116 (O_116,N_8458,N_9751);
or UO_117 (O_117,N_8429,N_8955);
nor UO_118 (O_118,N_8109,N_9766);
nand UO_119 (O_119,N_9963,N_8387);
nand UO_120 (O_120,N_8455,N_8072);
or UO_121 (O_121,N_8959,N_8320);
or UO_122 (O_122,N_9493,N_9932);
or UO_123 (O_123,N_8285,N_8392);
nand UO_124 (O_124,N_8557,N_9411);
or UO_125 (O_125,N_9950,N_9779);
and UO_126 (O_126,N_9567,N_8604);
nor UO_127 (O_127,N_9557,N_9858);
or UO_128 (O_128,N_9097,N_8194);
nand UO_129 (O_129,N_9842,N_8202);
or UO_130 (O_130,N_9747,N_9554);
nor UO_131 (O_131,N_8987,N_8472);
xnor UO_132 (O_132,N_9684,N_8924);
nand UO_133 (O_133,N_9161,N_9865);
and UO_134 (O_134,N_8307,N_8418);
nand UO_135 (O_135,N_9731,N_8594);
nand UO_136 (O_136,N_9614,N_9258);
nand UO_137 (O_137,N_8002,N_8017);
nor UO_138 (O_138,N_8670,N_8490);
or UO_139 (O_139,N_9368,N_8970);
and UO_140 (O_140,N_8874,N_9276);
or UO_141 (O_141,N_9696,N_8309);
nand UO_142 (O_142,N_9299,N_9473);
nor UO_143 (O_143,N_8634,N_9995);
nor UO_144 (O_144,N_9359,N_9911);
nor UO_145 (O_145,N_8044,N_9114);
nor UO_146 (O_146,N_9593,N_8516);
nand UO_147 (O_147,N_9224,N_9163);
nor UO_148 (O_148,N_8425,N_9965);
nor UO_149 (O_149,N_8311,N_8519);
and UO_150 (O_150,N_9909,N_8819);
nand UO_151 (O_151,N_8135,N_9616);
nand UO_152 (O_152,N_8199,N_8532);
nand UO_153 (O_153,N_8900,N_8858);
nor UO_154 (O_154,N_8952,N_9718);
or UO_155 (O_155,N_9148,N_9467);
nand UO_156 (O_156,N_8138,N_9035);
nor UO_157 (O_157,N_8514,N_8704);
nand UO_158 (O_158,N_8357,N_9574);
nand UO_159 (O_159,N_9244,N_8669);
or UO_160 (O_160,N_9241,N_9855);
and UO_161 (O_161,N_8218,N_8741);
and UO_162 (O_162,N_9078,N_8036);
and UO_163 (O_163,N_9484,N_8753);
nor UO_164 (O_164,N_8857,N_8275);
and UO_165 (O_165,N_9084,N_8278);
or UO_166 (O_166,N_9470,N_9343);
or UO_167 (O_167,N_9392,N_8349);
or UO_168 (O_168,N_8525,N_9890);
and UO_169 (O_169,N_9092,N_8408);
and UO_170 (O_170,N_9978,N_8950);
or UO_171 (O_171,N_8767,N_9294);
and UO_172 (O_172,N_9631,N_9756);
nor UO_173 (O_173,N_9303,N_9797);
and UO_174 (O_174,N_8372,N_9531);
xor UO_175 (O_175,N_9524,N_8912);
and UO_176 (O_176,N_8572,N_9327);
and UO_177 (O_177,N_8049,N_8783);
xnor UO_178 (O_178,N_9320,N_8590);
or UO_179 (O_179,N_9164,N_8113);
or UO_180 (O_180,N_8433,N_8317);
nor UO_181 (O_181,N_9693,N_9191);
and UO_182 (O_182,N_8716,N_8251);
xnor UO_183 (O_183,N_9627,N_8290);
xor UO_184 (O_184,N_8916,N_9206);
nand UO_185 (O_185,N_9992,N_9425);
and UO_186 (O_186,N_9324,N_8757);
xor UO_187 (O_187,N_8326,N_9827);
and UO_188 (O_188,N_9125,N_9534);
nand UO_189 (O_189,N_9542,N_8791);
or UO_190 (O_190,N_9935,N_8827);
nor UO_191 (O_191,N_8974,N_8076);
nor UO_192 (O_192,N_8379,N_8942);
nor UO_193 (O_193,N_8022,N_8033);
nand UO_194 (O_194,N_9420,N_9649);
or UO_195 (O_195,N_9902,N_9668);
or UO_196 (O_196,N_9576,N_9260);
and UO_197 (O_197,N_9555,N_8144);
nand UO_198 (O_198,N_8094,N_9233);
nand UO_199 (O_199,N_8189,N_8491);
and UO_200 (O_200,N_9540,N_8560);
nand UO_201 (O_201,N_8315,N_9507);
nor UO_202 (O_202,N_8370,N_8747);
xnor UO_203 (O_203,N_9069,N_8506);
nor UO_204 (O_204,N_9885,N_9110);
xor UO_205 (O_205,N_8700,N_8940);
xor UO_206 (O_206,N_9866,N_8756);
and UO_207 (O_207,N_9606,N_8947);
or UO_208 (O_208,N_9232,N_8358);
nor UO_209 (O_209,N_8341,N_9513);
or UO_210 (O_210,N_9223,N_9882);
nor UO_211 (O_211,N_8337,N_9784);
xor UO_212 (O_212,N_8035,N_9514);
and UO_213 (O_213,N_9854,N_9177);
nor UO_214 (O_214,N_8815,N_9003);
nor UO_215 (O_215,N_8192,N_9940);
or UO_216 (O_216,N_9344,N_8761);
nand UO_217 (O_217,N_9011,N_9323);
nand UO_218 (O_218,N_8499,N_9734);
or UO_219 (O_219,N_8665,N_9188);
nand UO_220 (O_220,N_8696,N_9054);
or UO_221 (O_221,N_8126,N_9585);
nand UO_222 (O_222,N_9942,N_9875);
nand UO_223 (O_223,N_9868,N_8143);
or UO_224 (O_224,N_9584,N_8843);
nand UO_225 (O_225,N_9917,N_9652);
or UO_226 (O_226,N_9980,N_8650);
and UO_227 (O_227,N_9430,N_9419);
nor UO_228 (O_228,N_9759,N_9948);
or UO_229 (O_229,N_9900,N_9505);
nor UO_230 (O_230,N_8648,N_9710);
or UO_231 (O_231,N_8087,N_8325);
and UO_232 (O_232,N_9930,N_8080);
or UO_233 (O_233,N_9445,N_8377);
xnor UO_234 (O_234,N_8225,N_8606);
nor UO_235 (O_235,N_9711,N_9568);
nor UO_236 (O_236,N_8838,N_8101);
xor UO_237 (O_237,N_8402,N_9796);
nand UO_238 (O_238,N_8255,N_8920);
or UO_239 (O_239,N_8925,N_9480);
nand UO_240 (O_240,N_8666,N_8457);
nand UO_241 (O_241,N_8242,N_9535);
and UO_242 (O_242,N_9515,N_9519);
nand UO_243 (O_243,N_8381,N_9450);
and UO_244 (O_244,N_8303,N_8088);
xnor UO_245 (O_245,N_8567,N_8717);
nand UO_246 (O_246,N_9789,N_8375);
or UO_247 (O_247,N_8177,N_9302);
or UO_248 (O_248,N_9946,N_9672);
or UO_249 (O_249,N_9442,N_9081);
and UO_250 (O_250,N_9564,N_9118);
and UO_251 (O_251,N_9708,N_9704);
and UO_252 (O_252,N_9803,N_9521);
nand UO_253 (O_253,N_9698,N_9570);
nand UO_254 (O_254,N_9754,N_8847);
nor UO_255 (O_255,N_9903,N_9831);
xor UO_256 (O_256,N_8174,N_8941);
nor UO_257 (O_257,N_8011,N_9530);
and UO_258 (O_258,N_8740,N_8889);
or UO_259 (O_259,N_8016,N_9296);
or UO_260 (O_260,N_8420,N_8748);
nand UO_261 (O_261,N_8191,N_8680);
or UO_262 (O_262,N_9072,N_8731);
nor UO_263 (O_263,N_8619,N_9262);
and UO_264 (O_264,N_8254,N_9622);
and UO_265 (O_265,N_8095,N_9213);
nand UO_266 (O_266,N_9860,N_8279);
nor UO_267 (O_267,N_9249,N_9483);
and UO_268 (O_268,N_8462,N_9912);
and UO_269 (O_269,N_9446,N_8622);
or UO_270 (O_270,N_9853,N_9651);
or UO_271 (O_271,N_8672,N_9964);
and UO_272 (O_272,N_8423,N_9522);
nand UO_273 (O_273,N_8347,N_9428);
and UO_274 (O_274,N_8719,N_9933);
or UO_275 (O_275,N_9615,N_9207);
or UO_276 (O_276,N_8030,N_8210);
nor UO_277 (O_277,N_9977,N_8273);
or UO_278 (O_278,N_8060,N_9132);
xor UO_279 (O_279,N_8335,N_8077);
or UO_280 (O_280,N_8176,N_8978);
nand UO_281 (O_281,N_8971,N_9660);
nand UO_282 (O_282,N_8656,N_9469);
nand UO_283 (O_283,N_9157,N_8494);
or UO_284 (O_284,N_9298,N_9409);
nor UO_285 (O_285,N_9498,N_8421);
nand UO_286 (O_286,N_8996,N_9399);
nor UO_287 (O_287,N_9028,N_8917);
or UO_288 (O_288,N_9353,N_9330);
nand UO_289 (O_289,N_9713,N_8693);
nand UO_290 (O_290,N_9620,N_9601);
or UO_291 (O_291,N_9438,N_8588);
and UO_292 (O_292,N_9745,N_8260);
nand UO_293 (O_293,N_8632,N_9150);
and UO_294 (O_294,N_8872,N_8714);
nand UO_295 (O_295,N_9007,N_8793);
and UO_296 (O_296,N_9468,N_8243);
or UO_297 (O_297,N_8091,N_9846);
and UO_298 (O_298,N_9321,N_8305);
or UO_299 (O_299,N_9881,N_9448);
nand UO_300 (O_300,N_8133,N_9809);
xnor UO_301 (O_301,N_9098,N_8610);
xor UO_302 (O_302,N_9795,N_8286);
xnor UO_303 (O_303,N_9801,N_8554);
or UO_304 (O_304,N_8334,N_9407);
xnor UO_305 (O_305,N_8231,N_9629);
nor UO_306 (O_306,N_8163,N_9386);
nor UO_307 (O_307,N_9595,N_9818);
nand UO_308 (O_308,N_9429,N_9758);
or UO_309 (O_309,N_9123,N_9943);
and UO_310 (O_310,N_9002,N_8609);
nand UO_311 (O_311,N_8682,N_8637);
nand UO_312 (O_312,N_8745,N_8730);
nor UO_313 (O_313,N_9136,N_8915);
xnor UO_314 (O_314,N_8496,N_9788);
and UO_315 (O_315,N_9173,N_8266);
or UO_316 (O_316,N_9836,N_8746);
and UO_317 (O_317,N_9355,N_9352);
nor UO_318 (O_318,N_8913,N_9669);
or UO_319 (O_319,N_8898,N_8306);
and UO_320 (O_320,N_8366,N_9501);
nor UO_321 (O_321,N_8431,N_8057);
and UO_322 (O_322,N_8193,N_9435);
or UO_323 (O_323,N_9322,N_9891);
or UO_324 (O_324,N_8201,N_9970);
nor UO_325 (O_325,N_8412,N_8488);
nand UO_326 (O_326,N_8371,N_8426);
or UO_327 (O_327,N_8269,N_8099);
and UO_328 (O_328,N_8406,N_9200);
or UO_329 (O_329,N_9109,N_8019);
and UO_330 (O_330,N_8345,N_9384);
or UO_331 (O_331,N_8851,N_8690);
nand UO_332 (O_332,N_8907,N_9899);
nand UO_333 (O_333,N_9709,N_8130);
or UO_334 (O_334,N_9495,N_9408);
or UO_335 (O_335,N_8511,N_8755);
or UO_336 (O_336,N_8247,N_9644);
nand UO_337 (O_337,N_9776,N_9134);
nand UO_338 (O_338,N_9738,N_9443);
nand UO_339 (O_339,N_8617,N_9375);
nand UO_340 (O_340,N_8071,N_8627);
nand UO_341 (O_341,N_9765,N_8168);
or UO_342 (O_342,N_8543,N_8401);
nor UO_343 (O_343,N_9619,N_9723);
xnor UO_344 (O_344,N_8620,N_9781);
or UO_345 (O_345,N_9162,N_8241);
nand UO_346 (O_346,N_8879,N_9849);
xor UO_347 (O_347,N_8958,N_8432);
and UO_348 (O_348,N_9523,N_9520);
xor UO_349 (O_349,N_8041,N_8932);
xor UO_350 (O_350,N_8283,N_9966);
nand UO_351 (O_351,N_8698,N_9329);
and UO_352 (O_352,N_8544,N_9126);
or UO_353 (O_353,N_8661,N_9197);
nand UO_354 (O_354,N_9929,N_8112);
or UO_355 (O_355,N_9168,N_9843);
nand UO_356 (O_356,N_8500,N_9596);
and UO_357 (O_357,N_9488,N_9577);
or UO_358 (O_358,N_8565,N_8155);
or UO_359 (O_359,N_9671,N_8281);
or UO_360 (O_360,N_8222,N_9226);
and UO_361 (O_361,N_8183,N_8507);
nand UO_362 (O_362,N_8015,N_8641);
nand UO_363 (O_363,N_9297,N_9722);
nand UO_364 (O_364,N_9300,N_8346);
nor UO_365 (O_365,N_8502,N_8023);
or UO_366 (O_366,N_8593,N_9985);
and UO_367 (O_367,N_9958,N_9333);
xnor UO_368 (O_368,N_9389,N_8644);
xor UO_369 (O_369,N_9367,N_8237);
nand UO_370 (O_370,N_8125,N_8981);
nand UO_371 (O_371,N_9339,N_9119);
or UO_372 (O_372,N_9283,N_9886);
nor UO_373 (O_373,N_9844,N_8901);
nor UO_374 (O_374,N_8788,N_8550);
nor UO_375 (O_375,N_9867,N_9444);
nor UO_376 (O_376,N_9221,N_9472);
nor UO_377 (O_377,N_8589,N_8265);
and UO_378 (O_378,N_8545,N_9356);
nand UO_379 (O_379,N_8580,N_9021);
or UO_380 (O_380,N_8014,N_8909);
nor UO_381 (O_381,N_9705,N_9563);
nand UO_382 (O_382,N_9724,N_9458);
nand UO_383 (O_383,N_9847,N_8535);
or UO_384 (O_384,N_9214,N_8652);
and UO_385 (O_385,N_9861,N_9220);
nor UO_386 (O_386,N_9925,N_8029);
xnor UO_387 (O_387,N_9525,N_9440);
xnor UO_388 (O_388,N_8451,N_9683);
and UO_389 (O_389,N_8070,N_9962);
and UO_390 (O_390,N_9494,N_8951);
and UO_391 (O_391,N_8291,N_9403);
or UO_392 (O_392,N_8208,N_8131);
nor UO_393 (O_393,N_9208,N_8820);
nand UO_394 (O_394,N_8624,N_8537);
and UO_395 (O_395,N_8640,N_9067);
or UO_396 (O_396,N_9983,N_9526);
and UO_397 (O_397,N_9871,N_9894);
xor UO_398 (O_398,N_8166,N_9763);
or UO_399 (O_399,N_9055,N_9179);
and UO_400 (O_400,N_8758,N_8078);
and UO_401 (O_401,N_8582,N_8010);
and UO_402 (O_402,N_8328,N_9133);
and UO_403 (O_403,N_8159,N_8800);
nand UO_404 (O_404,N_9036,N_8750);
nand UO_405 (O_405,N_9639,N_8086);
nor UO_406 (O_406,N_9015,N_9018);
or UO_407 (O_407,N_8446,N_8646);
or UO_408 (O_408,N_9895,N_8196);
nor UO_409 (O_409,N_8482,N_9553);
nand UO_410 (O_410,N_8428,N_8417);
nor UO_411 (O_411,N_8775,N_9828);
nor UO_412 (O_412,N_9987,N_9441);
xnor UO_413 (O_413,N_9412,N_9635);
and UO_414 (O_414,N_8769,N_9014);
nor UO_415 (O_415,N_8221,N_9152);
nor UO_416 (O_416,N_9235,N_8132);
nor UO_417 (O_417,N_9532,N_9915);
or UO_418 (O_418,N_8528,N_8413);
nor UO_419 (O_419,N_9510,N_8256);
nor UO_420 (O_420,N_9305,N_9310);
nand UO_421 (O_421,N_9107,N_8779);
nor UO_422 (O_422,N_9024,N_9490);
nand UO_423 (O_423,N_8009,N_9741);
xor UO_424 (O_424,N_8142,N_9988);
nor UO_425 (O_425,N_8389,N_9121);
or UO_426 (O_426,N_9979,N_8764);
xor UO_427 (O_427,N_8493,N_8351);
nand UO_428 (O_428,N_8117,N_8770);
nor UO_429 (O_429,N_8300,N_8069);
xnor UO_430 (O_430,N_8054,N_8470);
nor UO_431 (O_431,N_9415,N_9464);
nand UO_432 (O_432,N_8484,N_9461);
nand UO_433 (O_433,N_9938,N_9217);
nor UO_434 (O_434,N_9556,N_9994);
nor UO_435 (O_435,N_8445,N_8759);
or UO_436 (O_436,N_8106,N_9729);
nor UO_437 (O_437,N_8965,N_9537);
nand UO_438 (O_438,N_8424,N_8312);
or UO_439 (O_439,N_8368,N_9991);
nor UO_440 (O_440,N_9334,N_9180);
xnor UO_441 (O_441,N_8220,N_8013);
nor UO_442 (O_442,N_8893,N_9046);
and UO_443 (O_443,N_9956,N_9880);
nor UO_444 (O_444,N_8835,N_8988);
or UO_445 (O_445,N_8956,N_9437);
or UO_446 (O_446,N_8729,N_8896);
nor UO_447 (O_447,N_8883,N_9888);
and UO_448 (O_448,N_8304,N_9453);
nand UO_449 (O_449,N_9878,N_9295);
or UO_450 (O_450,N_9536,N_9145);
and UO_451 (O_451,N_8739,N_9089);
xor UO_452 (O_452,N_8399,N_8382);
and UO_453 (O_453,N_9820,N_9345);
xnor UO_454 (O_454,N_8274,N_9382);
nor UO_455 (O_455,N_8055,N_9026);
nor UO_456 (O_456,N_8878,N_8983);
nor UO_457 (O_457,N_8235,N_8715);
or UO_458 (O_458,N_9783,N_8569);
nor UO_459 (O_459,N_9699,N_8466);
and UO_460 (O_460,N_9189,N_8198);
nand UO_461 (O_461,N_8206,N_8803);
nor UO_462 (O_462,N_9715,N_9138);
nor UO_463 (O_463,N_9456,N_8564);
or UO_464 (O_464,N_9893,N_9612);
xnor UO_465 (O_465,N_8105,N_9043);
or UO_466 (O_466,N_9931,N_8853);
and UO_467 (O_467,N_9551,N_9391);
nand UO_468 (O_468,N_9008,N_8720);
nand UO_469 (O_469,N_9434,N_8103);
and UO_470 (O_470,N_8568,N_8263);
nor UO_471 (O_471,N_8276,N_8436);
xor UO_472 (O_472,N_8869,N_9174);
nand UO_473 (O_473,N_8989,N_9559);
or UO_474 (O_474,N_9016,N_8679);
xnor UO_475 (O_475,N_8613,N_9400);
xor UO_476 (O_476,N_9821,N_8327);
or UO_477 (O_477,N_8919,N_9219);
nand UO_478 (O_478,N_9840,N_8531);
nor UO_479 (O_479,N_9998,N_8635);
nor UO_480 (O_480,N_9259,N_8933);
and UO_481 (O_481,N_8870,N_8694);
nand UO_482 (O_482,N_8081,N_8782);
xor UO_483 (O_483,N_9856,N_8972);
or UO_484 (O_484,N_8295,N_9056);
nor UO_485 (O_485,N_9990,N_8523);
and UO_486 (O_486,N_9204,N_8430);
or UO_487 (O_487,N_8625,N_9071);
nor UO_488 (O_488,N_9506,N_9632);
nand UO_489 (O_489,N_9274,N_9786);
and UO_490 (O_490,N_9277,N_8626);
nor UO_491 (O_491,N_8170,N_8964);
and UO_492 (O_492,N_8007,N_8754);
nand UO_493 (O_493,N_9366,N_9726);
and UO_494 (O_494,N_8108,N_8185);
and UO_495 (O_495,N_8167,N_8863);
or UO_496 (O_496,N_9194,N_8164);
and UO_497 (O_497,N_8448,N_8452);
or UO_498 (O_498,N_8442,N_9176);
or UO_499 (O_499,N_8675,N_8323);
nand UO_500 (O_500,N_8985,N_9613);
or UO_501 (O_501,N_9012,N_8365);
and UO_502 (O_502,N_8724,N_9421);
and UO_503 (O_503,N_9266,N_8510);
nand UO_504 (O_504,N_9094,N_9769);
or UO_505 (O_505,N_8146,N_9679);
and UO_506 (O_506,N_8584,N_9588);
and UO_507 (O_507,N_9792,N_9143);
nand UO_508 (O_508,N_9785,N_8288);
nand UO_509 (O_509,N_9597,N_8513);
or UO_510 (O_510,N_9969,N_9216);
or UO_511 (O_511,N_8277,N_9242);
nor UO_512 (O_512,N_8718,N_9538);
or UO_513 (O_513,N_9128,N_8837);
and UO_514 (O_514,N_8969,N_8469);
and UO_515 (O_515,N_8703,N_8409);
xnor UO_516 (O_516,N_9034,N_9778);
or UO_517 (O_517,N_8150,N_9058);
xnor UO_518 (O_518,N_8027,N_8906);
nand UO_519 (O_519,N_8050,N_9088);
xor UO_520 (O_520,N_9675,N_8828);
nand UO_521 (O_521,N_9155,N_9928);
nor UO_522 (O_522,N_9240,N_8630);
nor UO_523 (O_523,N_8555,N_8405);
and UO_524 (O_524,N_8633,N_9290);
nor UO_525 (O_525,N_8228,N_8808);
or UO_526 (O_526,N_8172,N_8829);
nor UO_527 (O_527,N_9376,N_8092);
xnor UO_528 (O_528,N_9405,N_9192);
and UO_529 (O_529,N_8977,N_9976);
nand UO_530 (O_530,N_8139,N_9961);
or UO_531 (O_531,N_8492,N_9986);
nand UO_532 (O_532,N_9486,N_9328);
nand UO_533 (O_533,N_9830,N_8809);
and UO_534 (O_534,N_9032,N_9395);
xnor UO_535 (O_535,N_9256,N_8067);
nand UO_536 (O_536,N_9512,N_8561);
nor UO_537 (O_537,N_8213,N_8197);
and UO_538 (O_538,N_9452,N_8695);
and UO_539 (O_539,N_9131,N_9984);
xor UO_540 (O_540,N_9239,N_9497);
nand UO_541 (O_541,N_9664,N_8319);
and UO_542 (O_542,N_9127,N_9025);
nand UO_543 (O_543,N_8336,N_9752);
and UO_544 (O_544,N_9268,N_9541);
nor UO_545 (O_545,N_8114,N_9061);
and UO_546 (O_546,N_9433,N_9645);
nand UO_547 (O_547,N_8570,N_8881);
nor UO_548 (O_548,N_8085,N_8227);
nand UO_549 (O_549,N_9037,N_9782);
and UO_550 (O_550,N_8712,N_9059);
nor UO_551 (O_551,N_9397,N_8169);
nand UO_552 (O_552,N_9172,N_8995);
or UO_553 (O_553,N_9317,N_9689);
nand UO_554 (O_554,N_9780,N_9806);
nor UO_555 (O_555,N_9624,N_8781);
or UO_556 (O_556,N_9316,N_9006);
and UO_557 (O_557,N_8871,N_8539);
and UO_558 (O_558,N_9424,N_8692);
xnor UO_559 (O_559,N_8824,N_9757);
nor UO_560 (O_560,N_8481,N_8342);
nor UO_561 (O_561,N_9859,N_9142);
nor UO_562 (O_562,N_8025,N_8841);
nand UO_563 (O_563,N_8505,N_8005);
and UO_564 (O_564,N_9748,N_8332);
or UO_565 (O_565,N_8573,N_9422);
nand UO_566 (O_566,N_8726,N_8708);
or UO_567 (O_567,N_8410,N_8004);
and UO_568 (O_568,N_8642,N_9973);
nor UO_569 (O_569,N_8821,N_9154);
nand UO_570 (O_570,N_9167,N_9149);
or UO_571 (O_571,N_8270,N_8396);
nor UO_572 (O_572,N_8330,N_8236);
or UO_573 (O_573,N_9706,N_8434);
or UO_574 (O_574,N_9099,N_9657);
nor UO_575 (O_575,N_8533,N_9273);
nor UO_576 (O_576,N_8774,N_8968);
nand UO_577 (O_577,N_9804,N_9934);
nand UO_578 (O_578,N_8252,N_8184);
or UO_579 (O_579,N_9038,N_9975);
and UO_580 (O_580,N_9862,N_9662);
and UO_581 (O_581,N_8040,N_8240);
and UO_582 (O_582,N_9377,N_9431);
nand UO_583 (O_583,N_8161,N_9685);
and UO_584 (O_584,N_9460,N_8707);
or UO_585 (O_585,N_9802,N_8360);
nand UO_586 (O_586,N_8527,N_9835);
or UO_587 (O_587,N_8245,N_9009);
or UO_588 (O_588,N_9816,N_9372);
nand UO_589 (O_589,N_9518,N_8006);
nor UO_590 (O_590,N_9491,N_8160);
or UO_591 (O_591,N_9231,N_8230);
or UO_592 (O_592,N_9733,N_9005);
nor UO_593 (O_593,N_8540,N_8485);
xor UO_594 (O_594,N_8615,N_9762);
xnor UO_595 (O_595,N_9186,N_8662);
or UO_596 (O_596,N_8538,N_9451);
and UO_597 (O_597,N_9253,N_9907);
or UO_598 (O_598,N_9041,N_9311);
xnor UO_599 (O_599,N_9361,N_9807);
nor UO_600 (O_600,N_9826,N_8508);
and UO_601 (O_601,N_9454,N_9347);
nor UO_602 (O_602,N_9271,N_9920);
and UO_603 (O_603,N_8549,N_8599);
xnor UO_604 (O_604,N_8706,N_9677);
nand UO_605 (O_605,N_9637,N_9687);
nor UO_606 (O_606,N_9371,N_8148);
nand UO_607 (O_607,N_9545,N_9457);
nor UO_608 (O_608,N_9565,N_9065);
and UO_609 (O_609,N_9688,N_9654);
or UO_610 (O_610,N_9459,N_9288);
and UO_611 (O_611,N_8990,N_8784);
xor UO_612 (O_612,N_8153,N_9414);
nor UO_613 (O_613,N_8946,N_8744);
or UO_614 (O_614,N_8047,N_8850);
and UO_615 (O_615,N_8563,N_9730);
nor UO_616 (O_616,N_9573,N_9237);
nor UO_617 (O_617,N_8450,N_8894);
xor UO_618 (O_618,N_8647,N_9714);
or UO_619 (O_619,N_9336,N_8474);
or UO_620 (O_620,N_8558,N_8797);
or UO_621 (O_621,N_9279,N_8699);
or UO_622 (O_622,N_9618,N_8760);
nand UO_623 (O_623,N_8587,N_8713);
nor UO_624 (O_624,N_9517,N_8728);
and UO_625 (O_625,N_8331,N_9819);
nor UO_626 (O_626,N_8817,N_9261);
nand UO_627 (O_627,N_8975,N_9198);
and UO_628 (O_628,N_8127,N_9768);
nand UO_629 (O_629,N_8562,N_9650);
or UO_630 (O_630,N_8813,N_8145);
nand UO_631 (O_631,N_9904,N_9590);
nand UO_632 (O_632,N_9883,N_9743);
or UO_633 (O_633,N_8638,N_9222);
nor UO_634 (O_634,N_8380,N_9215);
nand UO_635 (O_635,N_9338,N_9922);
nor UO_636 (O_636,N_8301,N_8945);
nand UO_637 (O_637,N_9048,N_9401);
or UO_638 (O_638,N_8862,N_9609);
and UO_639 (O_639,N_9075,N_9736);
and UO_640 (O_640,N_9833,N_8217);
and UO_641 (O_641,N_8012,N_9087);
nor UO_642 (O_642,N_9636,N_8115);
or UO_643 (O_643,N_8374,N_8001);
and UO_644 (O_644,N_9250,N_9661);
or UO_645 (O_645,N_8903,N_9423);
nand UO_646 (O_646,N_9362,N_9982);
nand UO_647 (O_647,N_9959,N_8807);
nor UO_648 (O_648,N_8676,N_9941);
or UO_649 (O_649,N_8447,N_9905);
nor UO_650 (O_650,N_9053,N_9314);
and UO_651 (O_651,N_9953,N_8823);
or UO_652 (O_652,N_9640,N_9798);
and UO_653 (O_653,N_9471,N_9187);
nor UO_654 (O_654,N_9230,N_8643);
and UO_655 (O_655,N_8308,N_8123);
nand UO_656 (O_656,N_8891,N_9199);
or UO_657 (O_657,N_8607,N_8232);
and UO_658 (O_658,N_9774,N_9552);
or UO_659 (O_659,N_9052,N_9309);
or UO_660 (O_660,N_9023,N_9019);
and UO_661 (O_661,N_9418,N_9580);
or UO_662 (O_662,N_8734,N_8542);
or UO_663 (O_663,N_8895,N_8806);
and UO_664 (O_664,N_8119,N_9740);
nand UO_665 (O_665,N_8685,N_9117);
nor UO_666 (O_666,N_9633,N_9558);
or UO_667 (O_667,N_9586,N_9105);
nor UO_668 (O_668,N_8773,N_8489);
and UO_669 (O_669,N_9203,N_8310);
and UO_670 (O_670,N_8037,N_8344);
xor UO_671 (O_671,N_9010,N_8058);
nand UO_672 (O_672,N_8785,N_8464);
nor UO_673 (O_673,N_9870,N_8664);
nand UO_674 (O_674,N_8928,N_8073);
nand UO_675 (O_675,N_9380,N_8786);
or UO_676 (O_676,N_9913,N_8960);
and UO_677 (O_677,N_8921,N_9416);
and UO_678 (O_678,N_9598,N_8752);
xor UO_679 (O_679,N_8093,N_8725);
and UO_680 (O_680,N_9908,N_9079);
or UO_681 (O_681,N_9202,N_9690);
or UO_682 (O_682,N_9178,N_9923);
and UO_683 (O_683,N_9255,N_8032);
nand UO_684 (O_684,N_9971,N_9064);
xnor UO_685 (O_685,N_9974,N_8833);
nor UO_686 (O_686,N_8253,N_9209);
nand UO_687 (O_687,N_8667,N_9864);
nand UO_688 (O_688,N_9031,N_8885);
nor UO_689 (O_689,N_9236,N_8373);
nand UO_690 (O_690,N_9546,N_8422);
or UO_691 (O_691,N_8175,N_8854);
and UO_692 (O_692,N_8534,N_8602);
nand UO_693 (O_693,N_8427,N_9926);
or UO_694 (O_694,N_8158,N_9378);
xnor UO_695 (O_695,N_8855,N_8149);
and UO_696 (O_696,N_9605,N_8998);
and UO_697 (O_697,N_9665,N_8877);
xnor UO_698 (O_698,N_9799,N_8501);
or UO_699 (O_699,N_8691,N_9892);
and UO_700 (O_700,N_8805,N_9090);
and UO_701 (O_701,N_8856,N_8234);
nor UO_702 (O_702,N_8483,N_9529);
and UO_703 (O_703,N_8400,N_8601);
or UO_704 (O_704,N_9686,N_8280);
and UO_705 (O_705,N_9147,N_8264);
nand UO_706 (O_706,N_8961,N_8618);
nor UO_707 (O_707,N_8830,N_8261);
nand UO_708 (O_708,N_8911,N_9354);
and UO_709 (O_709,N_8937,N_9287);
xor UO_710 (O_710,N_9659,N_8018);
and UO_711 (O_711,N_9447,N_8476);
nand UO_712 (O_712,N_8355,N_8849);
and UO_713 (O_713,N_9682,N_8456);
nor UO_714 (O_714,N_9582,N_9169);
or UO_715 (O_715,N_8962,N_8861);
xnor UO_716 (O_716,N_8390,N_9516);
and UO_717 (O_717,N_8271,N_9393);
nor UO_718 (O_718,N_9889,N_8162);
and UO_719 (O_719,N_8751,N_8831);
nor UO_720 (O_720,N_9475,N_9544);
nor UO_721 (O_721,N_9360,N_9390);
and UO_722 (O_722,N_9863,N_8795);
or UO_723 (O_723,N_8089,N_9761);
and UO_724 (O_724,N_9937,N_9589);
nand UO_725 (O_725,N_9394,N_9077);
and UO_726 (O_726,N_9603,N_9739);
or UO_727 (O_727,N_9485,N_9417);
and UO_728 (O_728,N_9884,N_9402);
nand UO_729 (O_729,N_9212,N_9181);
and UO_730 (O_730,N_9095,N_8984);
and UO_731 (O_731,N_9284,N_8840);
xnor UO_732 (O_732,N_8415,N_9604);
nand UO_733 (O_733,N_8948,N_8697);
nor UO_734 (O_734,N_8350,N_8551);
or UO_735 (O_735,N_8340,N_9621);
nor UO_736 (O_736,N_9717,N_8042);
or UO_737 (O_737,N_9027,N_8780);
xor UO_738 (O_738,N_9120,N_8066);
nor UO_739 (O_739,N_9810,N_8369);
nand UO_740 (O_740,N_8926,N_8553);
or UO_741 (O_741,N_8802,N_8860);
or UO_742 (O_742,N_8651,N_8395);
nand UO_743 (O_743,N_8028,N_9703);
or UO_744 (O_744,N_8986,N_9653);
and UO_745 (O_745,N_9642,N_8503);
xor UO_746 (O_746,N_8842,N_8299);
nand UO_747 (O_747,N_9104,N_8865);
nor UO_748 (O_748,N_9477,N_8737);
or UO_749 (O_749,N_9436,N_8385);
or UO_750 (O_750,N_9286,N_8701);
or UO_751 (O_751,N_8616,N_8297);
nand UO_752 (O_752,N_9106,N_9171);
and UO_753 (O_753,N_8521,N_8137);
nand UO_754 (O_754,N_8934,N_8229);
nor UO_755 (O_755,N_8684,N_8526);
or UO_756 (O_756,N_9030,N_8219);
or UO_757 (O_757,N_8043,N_9547);
or UO_758 (O_758,N_8832,N_9272);
or UO_759 (O_759,N_8663,N_9201);
or UO_760 (O_760,N_8732,N_9379);
or UO_761 (O_761,N_9238,N_9251);
and UO_762 (O_762,N_8321,N_9972);
or UO_763 (O_763,N_9872,N_9144);
xnor UO_764 (O_764,N_9426,N_9914);
nand UO_765 (O_765,N_9292,N_9548);
and UO_766 (O_766,N_8478,N_9385);
xnor UO_767 (O_767,N_9815,N_9502);
or UO_768 (O_768,N_9465,N_9674);
nor UO_769 (O_769,N_9839,N_9658);
xnor UO_770 (O_770,N_9033,N_9346);
and UO_771 (O_771,N_9897,N_8449);
and UO_772 (O_772,N_8689,N_8504);
xnor UO_773 (O_773,N_8205,N_8683);
nand UO_774 (O_774,N_9628,N_8658);
nor UO_775 (O_775,N_8074,N_8353);
and UO_776 (O_776,N_8329,N_8075);
or UO_777 (O_777,N_8259,N_9042);
nor UO_778 (O_778,N_8814,N_9185);
nand UO_779 (O_779,N_9319,N_8178);
nand UO_780 (O_780,N_9050,N_9285);
nor UO_781 (O_781,N_8258,N_8497);
nand UO_782 (O_782,N_9634,N_8364);
nand UO_783 (O_783,N_9981,N_8628);
nand UO_784 (O_784,N_8173,N_8884);
nor UO_785 (O_785,N_8778,N_8008);
and UO_786 (O_786,N_8579,N_8914);
xor UO_787 (O_787,N_8629,N_9910);
nand UO_788 (O_788,N_8899,N_9949);
and UO_789 (O_789,N_9115,N_8608);
or UO_790 (O_790,N_9481,N_9838);
and UO_791 (O_791,N_8367,N_9057);
and UO_792 (O_792,N_8129,N_8825);
or UO_793 (O_793,N_8026,N_9100);
and UO_794 (O_794,N_8190,N_8776);
nor UO_795 (O_795,N_8444,N_9744);
xnor UO_796 (O_796,N_9370,N_9254);
nand UO_797 (O_797,N_9945,N_8727);
nand UO_798 (O_798,N_8062,N_9924);
or UO_799 (O_799,N_9753,N_9794);
and UO_800 (O_800,N_9267,N_9511);
or UO_801 (O_801,N_9489,N_8180);
or UO_802 (O_802,N_9499,N_9404);
nand UO_803 (O_803,N_8302,N_9313);
and UO_804 (O_804,N_9335,N_9697);
nor UO_805 (O_805,N_8226,N_8082);
or UO_806 (O_806,N_9921,N_9165);
and UO_807 (O_807,N_9474,N_8812);
nand UO_808 (O_808,N_9349,N_8294);
nand UO_809 (O_809,N_8203,N_8407);
nor UO_810 (O_810,N_8287,N_8723);
or UO_811 (O_811,N_9280,N_8772);
or UO_812 (O_812,N_9195,N_9196);
nand UO_813 (O_813,N_8826,N_9655);
or UO_814 (O_814,N_9387,N_9479);
or UO_815 (O_815,N_8388,N_8384);
and UO_816 (O_816,N_8465,N_9263);
or UO_817 (O_817,N_9022,N_8963);
xnor UO_818 (O_818,N_8065,N_9076);
nand UO_819 (O_819,N_8140,N_9996);
nor UO_820 (O_820,N_8179,N_9608);
nand UO_821 (O_821,N_9960,N_9967);
nor UO_822 (O_822,N_9772,N_8733);
nor UO_823 (O_823,N_9720,N_8063);
or UO_824 (O_824,N_8165,N_9771);
xnor UO_825 (O_825,N_9040,N_9850);
nand UO_826 (O_826,N_8515,N_8250);
or UO_827 (O_827,N_8118,N_9825);
and UO_828 (O_828,N_8541,N_9712);
or UO_829 (O_829,N_8239,N_8238);
xnor UO_830 (O_830,N_9824,N_8333);
xnor UO_831 (O_831,N_8468,N_9906);
and UO_832 (O_832,N_8518,N_9678);
xor UO_833 (O_833,N_8416,N_9135);
and UO_834 (O_834,N_8846,N_9252);
nand UO_835 (O_835,N_8098,N_8020);
xnor UO_836 (O_836,N_9845,N_9673);
xnor UO_837 (O_837,N_9129,N_8257);
and UO_838 (O_838,N_8048,N_8980);
nand UO_839 (O_839,N_9777,N_9045);
nor UO_840 (O_840,N_8313,N_8938);
nor UO_841 (O_841,N_8024,N_8147);
nor UO_842 (O_842,N_9800,N_9275);
xor UO_843 (O_843,N_8463,N_8156);
and UO_844 (O_844,N_8660,N_9834);
or UO_845 (O_845,N_8397,N_8064);
xor UO_846 (O_846,N_9066,N_9623);
and UO_847 (O_847,N_9304,N_9175);
and UO_848 (O_848,N_9728,N_9666);
and UO_849 (O_849,N_8792,N_8480);
nand UO_850 (O_850,N_9670,N_9611);
nand UO_851 (O_851,N_9082,N_9647);
nand UO_852 (O_852,N_9301,N_9153);
or UO_853 (O_853,N_9610,N_8973);
nand UO_854 (O_854,N_8154,N_9093);
and UO_855 (O_855,N_8211,N_9348);
and UO_856 (O_856,N_8393,N_9049);
and UO_857 (O_857,N_8559,N_8765);
or UO_858 (O_858,N_8460,N_9331);
and UO_859 (O_859,N_8867,N_9787);
or UO_860 (O_860,N_8439,N_9130);
nor UO_861 (O_861,N_8935,N_9725);
or UO_862 (O_862,N_9218,N_9572);
or UO_863 (O_863,N_8362,N_9993);
nor UO_864 (O_864,N_8888,N_8931);
nor UO_865 (O_865,N_9811,N_9225);
or UO_866 (O_866,N_9137,N_8267);
and UO_867 (O_867,N_8383,N_8391);
or UO_868 (O_868,N_9205,N_9643);
nor UO_869 (O_869,N_9646,N_8876);
nand UO_870 (O_870,N_8403,N_9308);
and UO_871 (O_871,N_8524,N_9281);
or UO_872 (O_872,N_9269,N_9767);
nor UO_873 (O_873,N_9496,N_9013);
nand UO_874 (O_874,N_9968,N_8289);
or UO_875 (O_875,N_8576,N_8818);
nor UO_876 (O_876,N_8777,N_9325);
and UO_877 (O_877,N_9158,N_9228);
and UO_878 (O_878,N_9790,N_9245);
xor UO_879 (O_879,N_9184,N_8376);
and UO_880 (O_880,N_8084,N_9719);
nand UO_881 (O_881,N_8673,N_8038);
and UO_882 (O_882,N_9569,N_8517);
xor UO_883 (O_883,N_8999,N_9562);
and UO_884 (O_884,N_9211,N_8943);
nand UO_885 (O_885,N_9156,N_9528);
nand UO_886 (O_886,N_8441,N_8722);
or UO_887 (O_887,N_9916,N_9243);
nor UO_888 (O_888,N_9051,N_8188);
and UO_889 (O_889,N_9000,N_8051);
or UO_890 (O_890,N_8411,N_9887);
nand UO_891 (O_891,N_8735,N_9550);
nor UO_892 (O_892,N_9351,N_9160);
or UO_893 (O_893,N_9732,N_8438);
or UO_894 (O_894,N_8314,N_9248);
or UO_895 (O_895,N_8966,N_8157);
nand UO_896 (O_896,N_8944,N_8195);
nand UO_897 (O_897,N_8709,N_9111);
or UO_898 (O_898,N_9410,N_9742);
or UO_899 (O_899,N_8394,N_9701);
or UO_900 (O_900,N_9509,N_9229);
nand UO_901 (O_901,N_9365,N_8486);
and UO_902 (O_902,N_8866,N_9265);
nand UO_903 (O_903,N_9997,N_8547);
nand UO_904 (O_904,N_8994,N_8339);
nand UO_905 (O_905,N_8298,N_9141);
or UO_906 (O_906,N_8771,N_9190);
and UO_907 (O_907,N_9879,N_9020);
or UO_908 (O_908,N_9773,N_9848);
or UO_909 (O_909,N_9939,N_8902);
nor UO_910 (O_910,N_8548,N_8721);
nand UO_911 (O_911,N_9039,N_9210);
and UO_912 (O_912,N_9581,N_8034);
nand UO_913 (O_913,N_9388,N_8461);
nand UO_914 (O_914,N_9478,N_8348);
and UO_915 (O_915,N_9508,N_9695);
and UO_916 (O_916,N_8435,N_8509);
nand UO_917 (O_917,N_9561,N_8918);
nor UO_918 (O_918,N_9113,N_9047);
xor UO_919 (O_919,N_9602,N_8102);
nand UO_920 (O_920,N_9247,N_8459);
nand UO_921 (O_921,N_9103,N_8354);
and UO_922 (O_922,N_8546,N_9648);
xnor UO_923 (O_923,N_8845,N_8487);
or UO_924 (O_924,N_9312,N_9791);
nor UO_925 (O_925,N_8440,N_9096);
and UO_926 (O_926,N_8316,N_8967);
nand UO_927 (O_927,N_9487,N_9579);
and UO_928 (O_928,N_8223,N_9070);
or UO_929 (O_929,N_8414,N_8811);
and UO_930 (O_930,N_8473,N_8039);
and UO_931 (O_931,N_8636,N_8882);
xor UO_932 (O_932,N_8586,N_9793);
nand UO_933 (O_933,N_9358,N_9702);
xnor UO_934 (O_934,N_8111,N_9318);
or UO_935 (O_935,N_9812,N_9841);
and UO_936 (O_936,N_8612,N_9449);
nor UO_937 (O_937,N_9307,N_8681);
and UO_938 (O_938,N_8530,N_8003);
nor UO_939 (O_939,N_8578,N_8577);
or UO_940 (O_940,N_8522,N_8880);
nand UO_941 (O_941,N_8120,N_9146);
nand UO_942 (O_942,N_8982,N_9735);
or UO_943 (O_943,N_9398,N_8090);
nor UO_944 (O_944,N_9264,N_9068);
and UO_945 (O_945,N_8677,N_8200);
nand UO_946 (O_946,N_8122,N_9492);
and UO_947 (O_947,N_8822,N_9080);
or UO_948 (O_948,N_8603,N_8649);
xor UO_949 (O_949,N_8639,N_8927);
xnor UO_950 (O_950,N_8743,N_9599);
nor UO_951 (O_951,N_9638,N_9282);
nand UO_952 (O_952,N_8498,N_8766);
nand UO_953 (O_953,N_8957,N_8655);
or UO_954 (O_954,N_9063,N_9085);
xor UO_955 (O_955,N_9291,N_8110);
or UO_956 (O_956,N_8892,N_8736);
or UO_957 (O_957,N_8296,N_8495);
or UO_958 (O_958,N_8097,N_9874);
nor UO_959 (O_959,N_8398,N_8124);
nand UO_960 (O_960,N_8873,N_8061);
nor UO_961 (O_961,N_8844,N_9183);
nor UO_962 (O_962,N_8363,N_9764);
nor UO_963 (O_963,N_8976,N_9116);
nor UO_964 (O_964,N_8045,N_9455);
and UO_965 (O_965,N_9560,N_8248);
xnor UO_966 (O_966,N_9680,N_8688);
or UO_967 (O_967,N_9583,N_8318);
and UO_968 (O_968,N_8686,N_8657);
nand UO_969 (O_969,N_9466,N_8574);
or UO_970 (O_970,N_9954,N_8215);
xor UO_971 (O_971,N_8991,N_8585);
nand UO_972 (O_972,N_9234,N_9396);
or UO_973 (O_973,N_8592,N_8437);
and UO_974 (O_974,N_9527,N_8187);
or UO_975 (O_975,N_9571,N_9707);
nor UO_976 (O_976,N_9503,N_8272);
nand UO_977 (O_977,N_8908,N_9357);
or UO_978 (O_978,N_8352,N_9681);
xnor UO_979 (O_979,N_8654,N_8212);
nor UO_980 (O_980,N_8404,N_8798);
nand UO_981 (O_981,N_9876,N_8566);
nor UO_982 (O_982,N_9151,N_8653);
nand UO_983 (O_983,N_8583,N_8671);
nand UO_984 (O_984,N_9805,N_9721);
nor UO_985 (O_985,N_8796,N_9124);
nand UO_986 (O_986,N_8897,N_8597);
nand UO_987 (O_987,N_8816,N_9694);
or UO_988 (O_988,N_9955,N_8799);
nand UO_989 (O_989,N_9170,N_9463);
nor UO_990 (O_990,N_8645,N_8922);
nor UO_991 (O_991,N_8801,N_9083);
nor UO_992 (O_992,N_9159,N_9482);
and UO_993 (O_993,N_9823,N_8182);
and UO_994 (O_994,N_8453,N_9944);
and UO_995 (O_995,N_8787,N_8581);
and UO_996 (O_996,N_9663,N_8595);
and UO_997 (O_997,N_9814,N_9750);
and UO_998 (O_998,N_8834,N_8687);
nand UO_999 (O_999,N_8598,N_9383);
or UO_1000 (O_1000,N_9699,N_9358);
xor UO_1001 (O_1001,N_9033,N_8366);
and UO_1002 (O_1002,N_8612,N_8683);
or UO_1003 (O_1003,N_9591,N_9041);
xor UO_1004 (O_1004,N_8404,N_9477);
and UO_1005 (O_1005,N_8733,N_9126);
or UO_1006 (O_1006,N_9722,N_8463);
or UO_1007 (O_1007,N_8026,N_8272);
nor UO_1008 (O_1008,N_8804,N_8612);
xor UO_1009 (O_1009,N_8164,N_8141);
nand UO_1010 (O_1010,N_9257,N_9770);
xnor UO_1011 (O_1011,N_9634,N_8060);
and UO_1012 (O_1012,N_9002,N_8764);
and UO_1013 (O_1013,N_9469,N_9420);
nor UO_1014 (O_1014,N_8200,N_8342);
or UO_1015 (O_1015,N_8764,N_8347);
xnor UO_1016 (O_1016,N_9517,N_9518);
nor UO_1017 (O_1017,N_8545,N_9583);
and UO_1018 (O_1018,N_9749,N_9375);
nand UO_1019 (O_1019,N_9056,N_9260);
nand UO_1020 (O_1020,N_9264,N_8850);
xor UO_1021 (O_1021,N_9051,N_9043);
nand UO_1022 (O_1022,N_8408,N_8804);
xnor UO_1023 (O_1023,N_8258,N_9821);
nand UO_1024 (O_1024,N_9934,N_8622);
nand UO_1025 (O_1025,N_8237,N_9330);
nor UO_1026 (O_1026,N_9411,N_8562);
nand UO_1027 (O_1027,N_8900,N_9205);
nand UO_1028 (O_1028,N_8028,N_9896);
or UO_1029 (O_1029,N_9634,N_8011);
or UO_1030 (O_1030,N_9993,N_8653);
and UO_1031 (O_1031,N_9020,N_8279);
and UO_1032 (O_1032,N_8701,N_8309);
xor UO_1033 (O_1033,N_8818,N_9535);
nor UO_1034 (O_1034,N_8529,N_8332);
nand UO_1035 (O_1035,N_9662,N_9457);
xor UO_1036 (O_1036,N_9115,N_8437);
or UO_1037 (O_1037,N_9402,N_8042);
or UO_1038 (O_1038,N_9651,N_9633);
xnor UO_1039 (O_1039,N_8635,N_9407);
or UO_1040 (O_1040,N_8528,N_9292);
nand UO_1041 (O_1041,N_8071,N_8724);
xor UO_1042 (O_1042,N_8473,N_8175);
or UO_1043 (O_1043,N_9270,N_8301);
nor UO_1044 (O_1044,N_9074,N_8174);
nor UO_1045 (O_1045,N_9319,N_9356);
nand UO_1046 (O_1046,N_8555,N_8988);
and UO_1047 (O_1047,N_9704,N_8837);
xor UO_1048 (O_1048,N_9467,N_8014);
or UO_1049 (O_1049,N_9043,N_9934);
nand UO_1050 (O_1050,N_9287,N_9572);
and UO_1051 (O_1051,N_8477,N_9657);
or UO_1052 (O_1052,N_8897,N_9454);
or UO_1053 (O_1053,N_8169,N_8157);
nor UO_1054 (O_1054,N_9648,N_9733);
nand UO_1055 (O_1055,N_9040,N_8924);
or UO_1056 (O_1056,N_8164,N_8429);
nand UO_1057 (O_1057,N_9390,N_9372);
nor UO_1058 (O_1058,N_8005,N_8346);
xnor UO_1059 (O_1059,N_9541,N_8771);
nand UO_1060 (O_1060,N_8295,N_8757);
and UO_1061 (O_1061,N_9123,N_9649);
and UO_1062 (O_1062,N_8661,N_8119);
and UO_1063 (O_1063,N_9265,N_9535);
or UO_1064 (O_1064,N_8072,N_8691);
or UO_1065 (O_1065,N_8160,N_8629);
nand UO_1066 (O_1066,N_9971,N_9353);
nor UO_1067 (O_1067,N_8218,N_9103);
nor UO_1068 (O_1068,N_9584,N_8788);
nand UO_1069 (O_1069,N_9626,N_8162);
and UO_1070 (O_1070,N_9833,N_9847);
and UO_1071 (O_1071,N_9499,N_9939);
and UO_1072 (O_1072,N_8600,N_9193);
xor UO_1073 (O_1073,N_8040,N_9881);
or UO_1074 (O_1074,N_9699,N_9543);
nor UO_1075 (O_1075,N_9288,N_9561);
and UO_1076 (O_1076,N_8356,N_9883);
or UO_1077 (O_1077,N_9876,N_9718);
or UO_1078 (O_1078,N_9087,N_9659);
or UO_1079 (O_1079,N_9037,N_8052);
or UO_1080 (O_1080,N_8582,N_8473);
and UO_1081 (O_1081,N_9138,N_8534);
nor UO_1082 (O_1082,N_8000,N_9208);
and UO_1083 (O_1083,N_9774,N_9730);
xor UO_1084 (O_1084,N_9842,N_8478);
and UO_1085 (O_1085,N_9828,N_9882);
nor UO_1086 (O_1086,N_9708,N_8256);
xnor UO_1087 (O_1087,N_9010,N_9115);
or UO_1088 (O_1088,N_9042,N_9483);
nor UO_1089 (O_1089,N_9958,N_8181);
nor UO_1090 (O_1090,N_8839,N_8851);
and UO_1091 (O_1091,N_9937,N_8679);
and UO_1092 (O_1092,N_8286,N_8136);
and UO_1093 (O_1093,N_9724,N_9964);
nor UO_1094 (O_1094,N_8397,N_9525);
and UO_1095 (O_1095,N_9965,N_9444);
nand UO_1096 (O_1096,N_9382,N_8649);
xnor UO_1097 (O_1097,N_9422,N_9680);
nor UO_1098 (O_1098,N_9104,N_8754);
nand UO_1099 (O_1099,N_9408,N_9601);
and UO_1100 (O_1100,N_8354,N_9459);
nand UO_1101 (O_1101,N_9936,N_8961);
xnor UO_1102 (O_1102,N_8930,N_9026);
or UO_1103 (O_1103,N_8083,N_8858);
and UO_1104 (O_1104,N_8326,N_9627);
or UO_1105 (O_1105,N_9521,N_8234);
or UO_1106 (O_1106,N_9141,N_9999);
nor UO_1107 (O_1107,N_9779,N_9496);
nand UO_1108 (O_1108,N_9932,N_8816);
nor UO_1109 (O_1109,N_8087,N_9091);
and UO_1110 (O_1110,N_9462,N_8320);
nor UO_1111 (O_1111,N_9800,N_9134);
nor UO_1112 (O_1112,N_8435,N_9937);
nand UO_1113 (O_1113,N_9136,N_8793);
or UO_1114 (O_1114,N_8569,N_8245);
xor UO_1115 (O_1115,N_8485,N_8138);
nand UO_1116 (O_1116,N_9522,N_9380);
nor UO_1117 (O_1117,N_9850,N_8382);
nor UO_1118 (O_1118,N_9540,N_9809);
xnor UO_1119 (O_1119,N_8434,N_9163);
xnor UO_1120 (O_1120,N_8184,N_8901);
nand UO_1121 (O_1121,N_9388,N_9380);
or UO_1122 (O_1122,N_9865,N_8972);
nor UO_1123 (O_1123,N_8476,N_8196);
and UO_1124 (O_1124,N_8760,N_8354);
or UO_1125 (O_1125,N_8950,N_9180);
or UO_1126 (O_1126,N_9277,N_9275);
nor UO_1127 (O_1127,N_8665,N_8484);
or UO_1128 (O_1128,N_9073,N_9267);
and UO_1129 (O_1129,N_9466,N_9149);
nor UO_1130 (O_1130,N_9927,N_9582);
nor UO_1131 (O_1131,N_8770,N_8245);
nor UO_1132 (O_1132,N_9875,N_9080);
nand UO_1133 (O_1133,N_9505,N_8153);
and UO_1134 (O_1134,N_9534,N_9337);
nand UO_1135 (O_1135,N_9422,N_8965);
or UO_1136 (O_1136,N_9307,N_8120);
and UO_1137 (O_1137,N_8176,N_9205);
nor UO_1138 (O_1138,N_9022,N_8965);
nor UO_1139 (O_1139,N_8766,N_9222);
nand UO_1140 (O_1140,N_9496,N_8059);
and UO_1141 (O_1141,N_8510,N_8552);
and UO_1142 (O_1142,N_8998,N_9373);
and UO_1143 (O_1143,N_8966,N_8459);
nand UO_1144 (O_1144,N_8735,N_8274);
xor UO_1145 (O_1145,N_9465,N_8739);
nor UO_1146 (O_1146,N_8722,N_9349);
nor UO_1147 (O_1147,N_9085,N_8561);
and UO_1148 (O_1148,N_8111,N_8405);
or UO_1149 (O_1149,N_9464,N_8197);
and UO_1150 (O_1150,N_8615,N_9088);
and UO_1151 (O_1151,N_8859,N_9983);
or UO_1152 (O_1152,N_8101,N_8100);
nand UO_1153 (O_1153,N_9033,N_8857);
nor UO_1154 (O_1154,N_9367,N_9161);
nor UO_1155 (O_1155,N_9442,N_9650);
and UO_1156 (O_1156,N_9905,N_8160);
xor UO_1157 (O_1157,N_9522,N_9397);
nand UO_1158 (O_1158,N_9452,N_8193);
or UO_1159 (O_1159,N_9630,N_9602);
nand UO_1160 (O_1160,N_9411,N_8703);
and UO_1161 (O_1161,N_8856,N_9092);
nand UO_1162 (O_1162,N_8436,N_9531);
nand UO_1163 (O_1163,N_9921,N_8304);
nand UO_1164 (O_1164,N_9154,N_9414);
or UO_1165 (O_1165,N_8688,N_8916);
nor UO_1166 (O_1166,N_9306,N_9145);
or UO_1167 (O_1167,N_8070,N_9848);
nor UO_1168 (O_1168,N_9466,N_8083);
and UO_1169 (O_1169,N_9412,N_9194);
and UO_1170 (O_1170,N_8506,N_9987);
nand UO_1171 (O_1171,N_8364,N_8890);
nor UO_1172 (O_1172,N_9169,N_8988);
or UO_1173 (O_1173,N_9849,N_9012);
nand UO_1174 (O_1174,N_8583,N_8189);
or UO_1175 (O_1175,N_8620,N_8595);
xor UO_1176 (O_1176,N_8757,N_8494);
or UO_1177 (O_1177,N_8964,N_8919);
nand UO_1178 (O_1178,N_8144,N_8803);
nand UO_1179 (O_1179,N_8164,N_8937);
or UO_1180 (O_1180,N_9533,N_8372);
nand UO_1181 (O_1181,N_8923,N_9141);
nand UO_1182 (O_1182,N_8206,N_9507);
and UO_1183 (O_1183,N_8968,N_8893);
nand UO_1184 (O_1184,N_9762,N_8384);
nor UO_1185 (O_1185,N_9046,N_8611);
nor UO_1186 (O_1186,N_9309,N_9382);
or UO_1187 (O_1187,N_9354,N_8933);
or UO_1188 (O_1188,N_8722,N_8819);
nand UO_1189 (O_1189,N_8448,N_9341);
nor UO_1190 (O_1190,N_8331,N_9783);
nor UO_1191 (O_1191,N_9834,N_8522);
nor UO_1192 (O_1192,N_8782,N_9901);
nor UO_1193 (O_1193,N_9054,N_8342);
and UO_1194 (O_1194,N_9780,N_9575);
nand UO_1195 (O_1195,N_8271,N_9071);
and UO_1196 (O_1196,N_8582,N_9969);
or UO_1197 (O_1197,N_9479,N_9821);
nor UO_1198 (O_1198,N_8944,N_8601);
and UO_1199 (O_1199,N_8204,N_8060);
nand UO_1200 (O_1200,N_8619,N_8614);
nor UO_1201 (O_1201,N_9724,N_9217);
xor UO_1202 (O_1202,N_9136,N_9980);
xnor UO_1203 (O_1203,N_8688,N_8096);
nor UO_1204 (O_1204,N_8368,N_8721);
nand UO_1205 (O_1205,N_8165,N_9676);
nor UO_1206 (O_1206,N_8221,N_9305);
nand UO_1207 (O_1207,N_8043,N_9065);
and UO_1208 (O_1208,N_8092,N_9100);
or UO_1209 (O_1209,N_9377,N_8563);
nand UO_1210 (O_1210,N_9497,N_8337);
or UO_1211 (O_1211,N_8617,N_8334);
and UO_1212 (O_1212,N_9024,N_8145);
nor UO_1213 (O_1213,N_9431,N_9666);
nand UO_1214 (O_1214,N_8759,N_9044);
or UO_1215 (O_1215,N_9136,N_8397);
or UO_1216 (O_1216,N_9051,N_9057);
nand UO_1217 (O_1217,N_8522,N_8127);
nand UO_1218 (O_1218,N_9253,N_8920);
or UO_1219 (O_1219,N_8948,N_9203);
and UO_1220 (O_1220,N_9575,N_9676);
nand UO_1221 (O_1221,N_9624,N_8144);
nand UO_1222 (O_1222,N_8843,N_8769);
and UO_1223 (O_1223,N_9610,N_9702);
or UO_1224 (O_1224,N_9729,N_8401);
nor UO_1225 (O_1225,N_9347,N_8183);
xnor UO_1226 (O_1226,N_9080,N_9168);
nor UO_1227 (O_1227,N_8940,N_9067);
nor UO_1228 (O_1228,N_9258,N_9461);
and UO_1229 (O_1229,N_9746,N_9652);
xnor UO_1230 (O_1230,N_9323,N_9939);
nand UO_1231 (O_1231,N_8804,N_9492);
xor UO_1232 (O_1232,N_8949,N_9138);
xnor UO_1233 (O_1233,N_9951,N_9845);
nor UO_1234 (O_1234,N_8562,N_9418);
nand UO_1235 (O_1235,N_9235,N_8724);
and UO_1236 (O_1236,N_9318,N_8484);
nor UO_1237 (O_1237,N_8230,N_8846);
or UO_1238 (O_1238,N_8673,N_8646);
or UO_1239 (O_1239,N_9922,N_9251);
and UO_1240 (O_1240,N_8017,N_9350);
and UO_1241 (O_1241,N_8369,N_9096);
or UO_1242 (O_1242,N_8970,N_8888);
nand UO_1243 (O_1243,N_9687,N_9321);
or UO_1244 (O_1244,N_8897,N_8201);
or UO_1245 (O_1245,N_8540,N_8182);
nand UO_1246 (O_1246,N_9041,N_9936);
and UO_1247 (O_1247,N_8535,N_9758);
nand UO_1248 (O_1248,N_9999,N_9269);
or UO_1249 (O_1249,N_9193,N_8287);
xor UO_1250 (O_1250,N_8750,N_9992);
nor UO_1251 (O_1251,N_8851,N_8156);
nand UO_1252 (O_1252,N_8551,N_9815);
or UO_1253 (O_1253,N_9368,N_8060);
nor UO_1254 (O_1254,N_9522,N_8725);
nor UO_1255 (O_1255,N_9342,N_8615);
and UO_1256 (O_1256,N_8953,N_9708);
nand UO_1257 (O_1257,N_8415,N_8414);
and UO_1258 (O_1258,N_8398,N_8585);
or UO_1259 (O_1259,N_8770,N_8072);
nor UO_1260 (O_1260,N_9744,N_8902);
and UO_1261 (O_1261,N_8685,N_8352);
nand UO_1262 (O_1262,N_9887,N_8934);
nor UO_1263 (O_1263,N_9101,N_8540);
and UO_1264 (O_1264,N_8521,N_8888);
nand UO_1265 (O_1265,N_8943,N_9208);
nor UO_1266 (O_1266,N_8668,N_9117);
or UO_1267 (O_1267,N_9876,N_9312);
and UO_1268 (O_1268,N_9184,N_8842);
or UO_1269 (O_1269,N_9534,N_9640);
nor UO_1270 (O_1270,N_9485,N_9892);
and UO_1271 (O_1271,N_9548,N_9841);
nand UO_1272 (O_1272,N_8458,N_8836);
nand UO_1273 (O_1273,N_9733,N_9947);
and UO_1274 (O_1274,N_8019,N_9144);
and UO_1275 (O_1275,N_9936,N_8634);
nand UO_1276 (O_1276,N_9995,N_8520);
nand UO_1277 (O_1277,N_8483,N_9632);
and UO_1278 (O_1278,N_9491,N_8261);
nand UO_1279 (O_1279,N_8828,N_9883);
and UO_1280 (O_1280,N_9155,N_9087);
or UO_1281 (O_1281,N_9541,N_8752);
and UO_1282 (O_1282,N_8077,N_8000);
nand UO_1283 (O_1283,N_8391,N_8800);
nand UO_1284 (O_1284,N_8335,N_9566);
and UO_1285 (O_1285,N_9551,N_8425);
or UO_1286 (O_1286,N_8779,N_8103);
or UO_1287 (O_1287,N_9544,N_9324);
nand UO_1288 (O_1288,N_8133,N_9624);
nand UO_1289 (O_1289,N_9665,N_9893);
xnor UO_1290 (O_1290,N_9526,N_9673);
nand UO_1291 (O_1291,N_9756,N_9582);
or UO_1292 (O_1292,N_9989,N_9043);
nor UO_1293 (O_1293,N_8041,N_8623);
and UO_1294 (O_1294,N_9258,N_9941);
nand UO_1295 (O_1295,N_9994,N_9169);
and UO_1296 (O_1296,N_8993,N_9154);
nor UO_1297 (O_1297,N_9845,N_9624);
nor UO_1298 (O_1298,N_9360,N_8531);
nor UO_1299 (O_1299,N_8245,N_8051);
nor UO_1300 (O_1300,N_9953,N_9696);
nand UO_1301 (O_1301,N_9098,N_8890);
or UO_1302 (O_1302,N_9329,N_9271);
and UO_1303 (O_1303,N_8748,N_9204);
nand UO_1304 (O_1304,N_9451,N_8732);
or UO_1305 (O_1305,N_8334,N_9633);
nand UO_1306 (O_1306,N_8801,N_8068);
and UO_1307 (O_1307,N_9578,N_9863);
or UO_1308 (O_1308,N_8811,N_8695);
or UO_1309 (O_1309,N_9536,N_9628);
and UO_1310 (O_1310,N_9887,N_8368);
nand UO_1311 (O_1311,N_9531,N_9823);
nand UO_1312 (O_1312,N_8817,N_8151);
and UO_1313 (O_1313,N_9998,N_9803);
or UO_1314 (O_1314,N_8421,N_9289);
nand UO_1315 (O_1315,N_9494,N_9955);
nand UO_1316 (O_1316,N_9386,N_8736);
xor UO_1317 (O_1317,N_8960,N_9510);
and UO_1318 (O_1318,N_8195,N_9380);
and UO_1319 (O_1319,N_9640,N_8613);
nor UO_1320 (O_1320,N_9748,N_8306);
nand UO_1321 (O_1321,N_8972,N_8574);
and UO_1322 (O_1322,N_9057,N_8569);
nor UO_1323 (O_1323,N_9915,N_9259);
or UO_1324 (O_1324,N_9065,N_8811);
and UO_1325 (O_1325,N_8927,N_8146);
or UO_1326 (O_1326,N_8858,N_8143);
or UO_1327 (O_1327,N_8604,N_9314);
or UO_1328 (O_1328,N_8327,N_9665);
nor UO_1329 (O_1329,N_9505,N_9676);
and UO_1330 (O_1330,N_8112,N_9867);
nand UO_1331 (O_1331,N_9318,N_8279);
and UO_1332 (O_1332,N_9504,N_9404);
nand UO_1333 (O_1333,N_8708,N_9157);
and UO_1334 (O_1334,N_9191,N_8054);
nor UO_1335 (O_1335,N_9753,N_9718);
and UO_1336 (O_1336,N_9918,N_8352);
or UO_1337 (O_1337,N_9759,N_8072);
nor UO_1338 (O_1338,N_9576,N_9259);
nand UO_1339 (O_1339,N_8900,N_8125);
nor UO_1340 (O_1340,N_9803,N_9046);
or UO_1341 (O_1341,N_8216,N_9519);
nand UO_1342 (O_1342,N_9616,N_9208);
or UO_1343 (O_1343,N_9879,N_9083);
nor UO_1344 (O_1344,N_8104,N_9996);
nor UO_1345 (O_1345,N_9420,N_8143);
and UO_1346 (O_1346,N_9187,N_9350);
nand UO_1347 (O_1347,N_9100,N_8044);
nor UO_1348 (O_1348,N_9287,N_8615);
nor UO_1349 (O_1349,N_8308,N_9141);
nor UO_1350 (O_1350,N_8851,N_9850);
and UO_1351 (O_1351,N_9436,N_8069);
nor UO_1352 (O_1352,N_8339,N_8633);
nor UO_1353 (O_1353,N_9522,N_9961);
and UO_1354 (O_1354,N_8827,N_9522);
nand UO_1355 (O_1355,N_8124,N_8267);
nand UO_1356 (O_1356,N_8967,N_9900);
nor UO_1357 (O_1357,N_8798,N_8496);
nor UO_1358 (O_1358,N_8952,N_9548);
or UO_1359 (O_1359,N_8894,N_9858);
and UO_1360 (O_1360,N_9406,N_9090);
nand UO_1361 (O_1361,N_8972,N_9316);
nor UO_1362 (O_1362,N_8308,N_9824);
nand UO_1363 (O_1363,N_8200,N_8934);
and UO_1364 (O_1364,N_9561,N_9606);
or UO_1365 (O_1365,N_8687,N_8640);
or UO_1366 (O_1366,N_8093,N_9996);
or UO_1367 (O_1367,N_8842,N_9244);
xnor UO_1368 (O_1368,N_8437,N_9655);
and UO_1369 (O_1369,N_9493,N_8750);
nand UO_1370 (O_1370,N_9504,N_8055);
or UO_1371 (O_1371,N_9464,N_8038);
nand UO_1372 (O_1372,N_8855,N_9090);
or UO_1373 (O_1373,N_8722,N_8750);
nor UO_1374 (O_1374,N_8749,N_9625);
or UO_1375 (O_1375,N_8745,N_9252);
nand UO_1376 (O_1376,N_8419,N_9566);
and UO_1377 (O_1377,N_9351,N_9511);
and UO_1378 (O_1378,N_9294,N_9881);
nand UO_1379 (O_1379,N_9107,N_8528);
xor UO_1380 (O_1380,N_9199,N_8628);
or UO_1381 (O_1381,N_9628,N_9630);
nor UO_1382 (O_1382,N_9373,N_8658);
and UO_1383 (O_1383,N_9306,N_8243);
nor UO_1384 (O_1384,N_8071,N_9134);
and UO_1385 (O_1385,N_8936,N_9015);
xnor UO_1386 (O_1386,N_9075,N_9745);
nor UO_1387 (O_1387,N_8588,N_9659);
nand UO_1388 (O_1388,N_9351,N_8327);
nor UO_1389 (O_1389,N_8053,N_8210);
or UO_1390 (O_1390,N_9517,N_9662);
nand UO_1391 (O_1391,N_9609,N_9177);
nand UO_1392 (O_1392,N_9863,N_8862);
nor UO_1393 (O_1393,N_9309,N_8451);
and UO_1394 (O_1394,N_9456,N_9284);
nand UO_1395 (O_1395,N_8380,N_8953);
or UO_1396 (O_1396,N_8028,N_9060);
nor UO_1397 (O_1397,N_9426,N_8029);
nor UO_1398 (O_1398,N_8702,N_8521);
and UO_1399 (O_1399,N_9447,N_9502);
nand UO_1400 (O_1400,N_8343,N_8657);
and UO_1401 (O_1401,N_8017,N_8773);
or UO_1402 (O_1402,N_9224,N_9014);
xor UO_1403 (O_1403,N_8045,N_9004);
or UO_1404 (O_1404,N_9362,N_9795);
or UO_1405 (O_1405,N_8921,N_8730);
or UO_1406 (O_1406,N_8732,N_8672);
xor UO_1407 (O_1407,N_8094,N_9285);
xnor UO_1408 (O_1408,N_9660,N_8148);
and UO_1409 (O_1409,N_9005,N_9457);
nand UO_1410 (O_1410,N_8328,N_8078);
or UO_1411 (O_1411,N_8112,N_9011);
nor UO_1412 (O_1412,N_8585,N_9383);
or UO_1413 (O_1413,N_8149,N_8551);
xnor UO_1414 (O_1414,N_8745,N_8687);
nor UO_1415 (O_1415,N_9653,N_8903);
nor UO_1416 (O_1416,N_9305,N_8108);
nor UO_1417 (O_1417,N_9896,N_9768);
xnor UO_1418 (O_1418,N_8555,N_9842);
or UO_1419 (O_1419,N_8026,N_8979);
and UO_1420 (O_1420,N_9283,N_8680);
or UO_1421 (O_1421,N_8089,N_8146);
or UO_1422 (O_1422,N_8862,N_8428);
xor UO_1423 (O_1423,N_9050,N_9202);
or UO_1424 (O_1424,N_8588,N_8763);
and UO_1425 (O_1425,N_9237,N_9101);
nor UO_1426 (O_1426,N_9052,N_9237);
nor UO_1427 (O_1427,N_8647,N_9991);
or UO_1428 (O_1428,N_9423,N_8199);
or UO_1429 (O_1429,N_8893,N_9183);
nor UO_1430 (O_1430,N_8655,N_9500);
nand UO_1431 (O_1431,N_8981,N_9266);
or UO_1432 (O_1432,N_8975,N_9813);
nand UO_1433 (O_1433,N_8030,N_8293);
nor UO_1434 (O_1434,N_9212,N_8388);
and UO_1435 (O_1435,N_8290,N_8710);
nor UO_1436 (O_1436,N_8580,N_9282);
nand UO_1437 (O_1437,N_8107,N_9639);
nor UO_1438 (O_1438,N_8978,N_9963);
nor UO_1439 (O_1439,N_8646,N_8194);
and UO_1440 (O_1440,N_9641,N_9941);
nand UO_1441 (O_1441,N_8709,N_9624);
or UO_1442 (O_1442,N_9341,N_9234);
and UO_1443 (O_1443,N_9647,N_9038);
or UO_1444 (O_1444,N_9599,N_9191);
nand UO_1445 (O_1445,N_8717,N_9318);
nand UO_1446 (O_1446,N_8699,N_8087);
and UO_1447 (O_1447,N_8260,N_8866);
nand UO_1448 (O_1448,N_9050,N_8564);
or UO_1449 (O_1449,N_8151,N_8603);
nand UO_1450 (O_1450,N_8772,N_8029);
and UO_1451 (O_1451,N_8843,N_8614);
nor UO_1452 (O_1452,N_9010,N_8665);
nor UO_1453 (O_1453,N_8659,N_9690);
nor UO_1454 (O_1454,N_9079,N_8862);
xor UO_1455 (O_1455,N_8208,N_8254);
nor UO_1456 (O_1456,N_9073,N_8040);
and UO_1457 (O_1457,N_9432,N_9833);
nand UO_1458 (O_1458,N_8984,N_9734);
xnor UO_1459 (O_1459,N_9758,N_8175);
and UO_1460 (O_1460,N_9154,N_9311);
nor UO_1461 (O_1461,N_8689,N_9436);
nand UO_1462 (O_1462,N_9380,N_8346);
or UO_1463 (O_1463,N_8271,N_9160);
nor UO_1464 (O_1464,N_9098,N_8306);
nor UO_1465 (O_1465,N_9955,N_9571);
xor UO_1466 (O_1466,N_8042,N_9561);
nand UO_1467 (O_1467,N_9887,N_8608);
and UO_1468 (O_1468,N_8033,N_8623);
nand UO_1469 (O_1469,N_8648,N_9872);
or UO_1470 (O_1470,N_8404,N_8823);
or UO_1471 (O_1471,N_8733,N_9460);
and UO_1472 (O_1472,N_8878,N_8599);
or UO_1473 (O_1473,N_9496,N_8162);
or UO_1474 (O_1474,N_9666,N_9612);
and UO_1475 (O_1475,N_8578,N_9234);
or UO_1476 (O_1476,N_9107,N_8488);
or UO_1477 (O_1477,N_8424,N_9637);
and UO_1478 (O_1478,N_9884,N_8066);
and UO_1479 (O_1479,N_8372,N_9713);
or UO_1480 (O_1480,N_8255,N_8337);
and UO_1481 (O_1481,N_9065,N_8150);
nand UO_1482 (O_1482,N_8831,N_8559);
nand UO_1483 (O_1483,N_9817,N_9130);
nor UO_1484 (O_1484,N_8694,N_8368);
nor UO_1485 (O_1485,N_9867,N_9705);
or UO_1486 (O_1486,N_9083,N_9244);
and UO_1487 (O_1487,N_9856,N_8258);
nand UO_1488 (O_1488,N_9033,N_9340);
or UO_1489 (O_1489,N_8535,N_9601);
or UO_1490 (O_1490,N_9228,N_9923);
nor UO_1491 (O_1491,N_9188,N_8387);
and UO_1492 (O_1492,N_9980,N_8454);
nor UO_1493 (O_1493,N_9012,N_8995);
and UO_1494 (O_1494,N_8113,N_8884);
nand UO_1495 (O_1495,N_8862,N_8601);
nor UO_1496 (O_1496,N_9695,N_8496);
nor UO_1497 (O_1497,N_8177,N_9997);
or UO_1498 (O_1498,N_8570,N_8562);
and UO_1499 (O_1499,N_8561,N_9327);
endmodule