module basic_1500_15000_2000_20_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_727,In_1494);
nand U1 (N_1,In_772,In_672);
nand U2 (N_2,In_1478,In_685);
nor U3 (N_3,In_124,In_68);
and U4 (N_4,In_1171,In_1033);
or U5 (N_5,In_638,In_984);
or U6 (N_6,In_1022,In_405);
nand U7 (N_7,In_504,In_283);
nor U8 (N_8,In_600,In_397);
and U9 (N_9,In_636,In_307);
or U10 (N_10,In_565,In_35);
xor U11 (N_11,In_438,In_666);
and U12 (N_12,In_905,In_325);
nand U13 (N_13,In_312,In_48);
nand U14 (N_14,In_778,In_590);
or U15 (N_15,In_191,In_1416);
and U16 (N_16,In_308,In_616);
nand U17 (N_17,In_228,In_701);
nor U18 (N_18,In_1,In_844);
nand U19 (N_19,In_907,In_737);
nand U20 (N_20,In_761,In_225);
xor U21 (N_21,In_40,In_1231);
xnor U22 (N_22,In_1151,In_474);
nor U23 (N_23,In_917,In_708);
or U24 (N_24,In_190,In_525);
and U25 (N_25,In_1343,In_835);
nor U26 (N_26,In_1107,In_1496);
nand U27 (N_27,In_1443,In_112);
and U28 (N_28,In_1346,In_1261);
nand U29 (N_29,In_1075,In_482);
nor U30 (N_30,In_533,In_650);
nor U31 (N_31,In_94,In_161);
and U32 (N_32,In_1334,In_285);
nor U33 (N_33,In_986,In_87);
nor U34 (N_34,In_802,In_207);
and U35 (N_35,In_412,In_997);
nor U36 (N_36,In_1299,In_1275);
or U37 (N_37,In_1253,In_764);
nor U38 (N_38,In_807,In_1193);
or U39 (N_39,In_377,In_1441);
and U40 (N_40,In_88,In_828);
and U41 (N_41,In_169,In_732);
nand U42 (N_42,In_555,In_1139);
nor U43 (N_43,In_1276,In_1135);
nor U44 (N_44,In_860,In_54);
xor U45 (N_45,In_181,In_479);
nand U46 (N_46,In_469,In_591);
and U47 (N_47,In_619,In_795);
nor U48 (N_48,In_1472,In_463);
nand U49 (N_49,In_970,In_961);
nand U50 (N_50,In_951,In_382);
or U51 (N_51,In_1322,In_402);
or U52 (N_52,In_1485,In_959);
or U53 (N_53,In_1398,In_938);
nor U54 (N_54,In_343,In_461);
or U55 (N_55,In_73,In_639);
nand U56 (N_56,In_233,In_1024);
nand U57 (N_57,In_769,In_282);
nor U58 (N_58,In_1187,In_381);
nand U59 (N_59,In_787,In_925);
or U60 (N_60,In_42,In_695);
or U61 (N_61,In_768,In_1399);
nor U62 (N_62,In_1116,In_1094);
or U63 (N_63,In_257,In_184);
and U64 (N_64,In_738,In_155);
or U65 (N_65,In_836,In_369);
nand U66 (N_66,In_515,In_483);
and U67 (N_67,In_934,In_566);
nor U68 (N_68,In_739,In_306);
or U69 (N_69,In_1360,In_110);
or U70 (N_70,In_1464,In_9);
nand U71 (N_71,In_1270,In_539);
nand U72 (N_72,In_60,In_1384);
nor U73 (N_73,In_960,In_1450);
or U74 (N_74,In_454,In_676);
nand U75 (N_75,In_256,In_1380);
or U76 (N_76,In_661,In_1027);
and U77 (N_77,In_1148,In_770);
nor U78 (N_78,In_1310,In_1195);
xnor U79 (N_79,In_76,In_1141);
nand U80 (N_80,In_611,In_99);
nor U81 (N_81,In_909,In_355);
nor U82 (N_82,In_602,In_678);
or U83 (N_83,In_940,In_77);
nand U84 (N_84,In_126,In_1348);
nor U85 (N_85,In_850,In_1045);
xor U86 (N_86,In_1272,In_496);
nor U87 (N_87,In_1475,In_1216);
xnor U88 (N_88,In_36,In_598);
and U89 (N_89,In_982,In_927);
nor U90 (N_90,In_1482,In_398);
nor U91 (N_91,In_432,In_908);
or U92 (N_92,In_544,In_197);
nand U93 (N_93,In_958,In_164);
or U94 (N_94,In_100,In_1223);
nand U95 (N_95,In_689,In_945);
or U96 (N_96,In_728,In_129);
nand U97 (N_97,In_581,In_471);
nand U98 (N_98,In_631,In_1147);
xor U99 (N_99,In_1473,In_304);
nor U100 (N_100,In_509,In_1286);
or U101 (N_101,In_1397,In_535);
nor U102 (N_102,In_1489,In_131);
or U103 (N_103,In_104,In_105);
or U104 (N_104,In_706,In_275);
and U105 (N_105,In_675,In_1121);
xor U106 (N_106,In_599,In_31);
nand U107 (N_107,In_3,In_1209);
or U108 (N_108,In_752,In_683);
or U109 (N_109,In_627,In_289);
and U110 (N_110,In_107,In_258);
nor U111 (N_111,In_594,In_1156);
nand U112 (N_112,In_1032,In_1467);
or U113 (N_113,In_799,In_116);
nor U114 (N_114,In_429,In_362);
xor U115 (N_115,In_295,In_348);
nor U116 (N_116,In_710,In_1492);
and U117 (N_117,In_494,In_530);
and U118 (N_118,In_1145,In_1059);
nor U119 (N_119,In_58,In_1378);
nand U120 (N_120,In_878,In_447);
nor U121 (N_121,In_1211,In_735);
nor U122 (N_122,In_121,In_936);
nand U123 (N_123,In_19,In_97);
and U124 (N_124,In_895,In_1428);
nand U125 (N_125,In_1029,In_929);
nor U126 (N_126,In_726,In_839);
nand U127 (N_127,In_1290,In_711);
nand U128 (N_128,In_404,In_317);
nor U129 (N_129,In_1285,In_941);
or U130 (N_130,In_21,In_705);
or U131 (N_131,In_490,In_903);
nand U132 (N_132,In_550,In_871);
nor U133 (N_133,In_990,In_645);
xnor U134 (N_134,In_491,In_1407);
nor U135 (N_135,In_204,In_1037);
nand U136 (N_136,In_758,In_250);
and U137 (N_137,In_1008,In_406);
nor U138 (N_138,In_1184,In_441);
or U139 (N_139,In_6,In_1048);
nor U140 (N_140,In_367,In_712);
nand U141 (N_141,In_1414,In_1143);
or U142 (N_142,In_1257,In_648);
and U143 (N_143,In_1000,In_651);
or U144 (N_144,In_538,In_460);
nand U145 (N_145,In_98,In_1199);
nor U146 (N_146,In_75,In_588);
and U147 (N_147,In_324,In_1132);
and U148 (N_148,In_840,In_623);
or U149 (N_149,In_380,In_760);
nor U150 (N_150,In_403,In_1434);
and U151 (N_151,In_1134,In_937);
and U152 (N_152,In_239,In_1046);
or U153 (N_153,In_1375,In_407);
and U154 (N_154,In_477,In_580);
and U155 (N_155,In_597,In_755);
nor U156 (N_156,In_1152,In_1198);
xnor U157 (N_157,In_1393,In_891);
nor U158 (N_158,In_1294,In_847);
or U159 (N_159,In_1469,In_459);
and U160 (N_160,In_357,In_794);
nor U161 (N_161,In_323,In_366);
and U162 (N_162,In_1004,In_352);
nor U163 (N_163,In_514,In_302);
xor U164 (N_164,In_1210,In_526);
xnor U165 (N_165,In_1074,In_1459);
and U166 (N_166,In_618,In_299);
and U167 (N_167,In_427,In_488);
or U168 (N_168,In_417,In_863);
nor U169 (N_169,In_291,In_866);
nor U170 (N_170,In_1361,In_249);
nor U171 (N_171,In_390,In_342);
xnor U172 (N_172,In_1355,In_1205);
nand U173 (N_173,In_767,In_521);
nor U174 (N_174,In_27,In_1268);
and U175 (N_175,In_1206,In_1288);
or U176 (N_176,In_1405,In_1289);
and U177 (N_177,In_893,In_884);
and U178 (N_178,In_1096,In_1076);
nand U179 (N_179,In_101,In_862);
or U180 (N_180,In_243,In_842);
xor U181 (N_181,In_215,In_911);
nand U182 (N_182,In_1435,In_644);
or U183 (N_183,In_217,In_1153);
nand U184 (N_184,In_805,In_1243);
nor U185 (N_185,In_41,In_725);
nor U186 (N_186,In_1367,In_480);
or U187 (N_187,In_1326,In_797);
or U188 (N_188,In_487,In_1300);
nor U189 (N_189,In_1460,In_817);
nor U190 (N_190,In_679,In_913);
nor U191 (N_191,In_1126,In_139);
nor U192 (N_192,In_1189,In_1035);
or U193 (N_193,In_1279,In_142);
and U194 (N_194,In_1425,In_1330);
and U195 (N_195,In_775,In_1474);
nor U196 (N_196,In_790,In_232);
nor U197 (N_197,In_1018,In_271);
and U198 (N_198,In_125,In_159);
and U199 (N_199,In_437,In_1258);
and U200 (N_200,In_720,In_694);
or U201 (N_201,In_151,In_95);
nand U202 (N_202,In_700,In_974);
and U203 (N_203,In_507,In_1431);
nand U204 (N_204,In_655,In_292);
nor U205 (N_205,In_50,In_33);
nor U206 (N_206,In_821,In_85);
nor U207 (N_207,In_1142,In_1287);
nor U208 (N_208,In_495,In_829);
nor U209 (N_209,In_1341,In_1255);
nand U210 (N_210,In_212,In_1138);
or U211 (N_211,In_1026,In_718);
nand U212 (N_212,In_1201,In_358);
and U213 (N_213,In_1240,In_1207);
or U214 (N_214,In_1127,In_1117);
or U215 (N_215,In_187,In_90);
or U216 (N_216,In_854,In_691);
or U217 (N_217,In_1386,In_920);
nand U218 (N_218,In_313,In_742);
or U219 (N_219,In_1063,In_183);
nor U220 (N_220,In_696,In_11);
and U221 (N_221,In_702,In_1477);
nand U222 (N_222,In_1222,In_57);
and U223 (N_223,In_133,In_815);
and U224 (N_224,In_26,In_1146);
nand U225 (N_225,In_994,In_527);
nand U226 (N_226,In_579,In_176);
or U227 (N_227,In_1486,In_1248);
nand U228 (N_228,In_944,In_420);
nand U229 (N_229,In_1093,In_154);
or U230 (N_230,In_965,In_269);
nand U231 (N_231,In_901,In_1200);
xor U232 (N_232,In_692,In_1254);
or U233 (N_233,In_595,In_1365);
and U234 (N_234,In_793,In_740);
xor U235 (N_235,In_8,In_556);
or U236 (N_236,In_956,In_673);
nand U237 (N_237,In_1252,In_368);
or U238 (N_238,In_475,In_1172);
and U239 (N_239,In_1364,In_52);
nand U240 (N_240,In_567,In_1323);
xor U241 (N_241,In_1176,In_1418);
and U242 (N_242,In_1455,In_410);
and U243 (N_243,In_470,In_175);
nand U244 (N_244,In_1087,In_1149);
nor U245 (N_245,In_660,In_723);
nor U246 (N_246,In_346,In_559);
and U247 (N_247,In_721,In_1266);
or U248 (N_248,In_468,In_549);
nor U249 (N_249,In_677,In_806);
and U250 (N_250,In_259,In_456);
nor U251 (N_251,In_1065,In_684);
and U252 (N_252,In_422,In_583);
nand U253 (N_253,In_1180,In_800);
or U254 (N_254,In_857,In_1498);
or U255 (N_255,In_798,In_1395);
or U256 (N_256,In_569,In_1133);
nor U257 (N_257,In_1379,In_1389);
xnor U258 (N_258,In_1280,In_536);
and U259 (N_259,In_516,In_1235);
and U260 (N_260,In_1366,In_56);
nand U261 (N_261,In_1442,In_1354);
nand U262 (N_262,In_66,In_61);
and U263 (N_263,In_180,In_848);
nand U264 (N_264,In_37,In_1043);
nor U265 (N_265,In_1462,In_545);
and U266 (N_266,In_1369,In_411);
and U267 (N_267,In_344,In_1137);
nand U268 (N_268,In_140,In_869);
nor U269 (N_269,In_1017,In_868);
nand U270 (N_270,In_122,In_251);
nor U271 (N_271,In_179,In_17);
xnor U272 (N_272,In_1150,In_141);
or U273 (N_273,In_575,In_1256);
nor U274 (N_274,In_1038,In_703);
nor U275 (N_275,In_788,In_394);
and U276 (N_276,In_267,In_642);
nand U277 (N_277,In_156,In_260);
nand U278 (N_278,In_1073,In_209);
and U279 (N_279,In_478,In_13);
nor U280 (N_280,In_1100,In_1362);
nand U281 (N_281,In_316,In_238);
nand U282 (N_282,In_326,In_656);
nand U283 (N_283,In_1174,In_1005);
or U284 (N_284,In_808,In_1274);
and U285 (N_285,In_263,In_255);
nand U286 (N_286,In_601,In_1480);
and U287 (N_287,In_174,In_1404);
nor U288 (N_288,In_995,In_949);
or U289 (N_289,In_34,In_446);
or U290 (N_290,In_32,In_1356);
nand U291 (N_291,In_1284,In_28);
or U292 (N_292,In_379,In_560);
nand U293 (N_293,In_485,In_1490);
and U294 (N_294,In_1324,In_1186);
xnor U295 (N_295,In_51,In_1120);
nand U296 (N_296,In_520,In_1451);
xor U297 (N_297,In_301,In_46);
nand U298 (N_298,In_864,In_1337);
and U299 (N_299,In_149,In_551);
and U300 (N_300,In_1164,In_473);
or U301 (N_301,In_278,In_168);
nand U302 (N_302,In_1122,In_1085);
and U303 (N_303,In_1304,In_219);
xor U304 (N_304,In_1099,In_210);
and U305 (N_305,In_522,In_1055);
nand U306 (N_306,In_421,In_1196);
nor U307 (N_307,In_12,In_596);
xnor U308 (N_308,In_436,In_153);
xor U309 (N_309,In_1316,In_464);
nor U310 (N_310,In_236,In_1039);
xor U311 (N_311,In_237,In_1488);
or U312 (N_312,In_814,In_163);
nor U313 (N_313,In_783,In_782);
nand U314 (N_314,In_363,In_1106);
nor U315 (N_315,In_640,In_288);
nor U316 (N_316,In_1463,In_743);
or U317 (N_317,In_719,In_1349);
or U318 (N_318,In_1173,In_199);
and U319 (N_319,In_1471,In_1079);
nor U320 (N_320,In_628,In_1333);
and U321 (N_321,In_1111,In_115);
and U322 (N_322,In_353,In_1358);
nor U323 (N_323,In_201,In_1371);
xnor U324 (N_324,In_218,In_1052);
nor U325 (N_325,In_582,In_717);
nor U326 (N_326,In_883,In_327);
and U327 (N_327,In_966,In_264);
xnor U328 (N_328,In_423,In_562);
nand U329 (N_329,In_1329,In_546);
xnor U330 (N_330,In_593,In_753);
nor U331 (N_331,In_1381,In_1229);
and U332 (N_332,In_383,In_855);
nand U333 (N_333,In_500,In_192);
and U334 (N_334,In_1188,In_334);
and U335 (N_335,In_1320,In_1204);
xor U336 (N_336,In_501,In_347);
and U337 (N_337,In_426,In_189);
and U338 (N_338,In_178,In_1491);
or U339 (N_339,In_273,In_846);
or U340 (N_340,In_502,In_221);
and U341 (N_341,In_823,In_1102);
and U342 (N_342,In_682,In_333);
and U343 (N_343,In_1015,In_1128);
and U344 (N_344,In_613,In_1160);
nand U345 (N_345,In_607,In_413);
nand U346 (N_346,In_853,In_1267);
or U347 (N_347,In_1430,In_796);
or U348 (N_348,In_177,In_942);
and U349 (N_349,In_513,In_103);
and U350 (N_350,In_1031,In_1377);
nand U351 (N_351,In_472,In_923);
or U352 (N_352,In_592,In_950);
or U353 (N_353,In_572,In_418);
nor U354 (N_354,In_455,In_335);
or U355 (N_355,In_1466,In_1495);
nand U356 (N_356,In_584,In_939);
and U357 (N_357,In_999,In_667);
and U358 (N_358,In_64,In_1309);
nor U359 (N_359,In_336,In_298);
nor U360 (N_360,In_1129,In_303);
or U361 (N_361,In_43,In_1056);
nand U362 (N_362,In_898,In_963);
nor U363 (N_363,In_157,In_230);
nand U364 (N_364,In_216,In_89);
and U365 (N_365,In_1327,In_763);
nor U366 (N_366,In_268,In_320);
and U367 (N_367,In_1387,In_635);
or U368 (N_368,In_211,In_453);
and U369 (N_369,In_561,In_130);
nand U370 (N_370,In_1400,In_1244);
nor U371 (N_371,In_246,In_486);
or U372 (N_372,In_29,In_374);
or U373 (N_373,In_874,In_1057);
xnor U374 (N_374,In_1006,In_1020);
and U375 (N_375,In_1083,In_765);
or U376 (N_376,In_1417,In_1090);
or U377 (N_377,In_892,In_387);
nand U378 (N_378,In_146,In_1250);
and U379 (N_379,In_467,In_851);
or U380 (N_380,In_1307,In_573);
nor U381 (N_381,In_305,In_1166);
xnor U382 (N_382,In_617,In_1476);
and U383 (N_383,In_1202,In_499);
nand U384 (N_384,In_693,In_756);
nor U385 (N_385,In_558,In_1217);
nor U386 (N_386,In_71,In_1060);
and U387 (N_387,In_332,In_870);
nand U388 (N_388,In_1383,In_1112);
or U389 (N_389,In_1318,In_1497);
nand U390 (N_390,In_668,In_1155);
and U391 (N_391,In_1260,In_395);
nor U392 (N_392,In_372,In_449);
nand U393 (N_393,In_1419,In_1273);
and U394 (N_394,In_193,In_136);
xor U395 (N_395,In_605,In_881);
xnor U396 (N_396,In_396,In_906);
nand U397 (N_397,In_910,In_1242);
nor U398 (N_398,In_5,In_896);
nand U399 (N_399,In_445,In_1344);
and U400 (N_400,In_1277,In_1221);
nor U401 (N_401,In_1426,In_262);
xnor U402 (N_402,In_370,In_248);
nor U403 (N_403,In_329,In_816);
and U404 (N_404,In_1282,In_652);
xor U405 (N_405,In_1078,In_277);
and U406 (N_406,In_505,In_875);
nor U407 (N_407,In_813,In_1119);
nand U408 (N_408,In_80,In_206);
xnor U409 (N_409,In_1336,In_663);
nand U410 (N_410,In_14,In_967);
nand U411 (N_411,In_1203,In_63);
nor U412 (N_412,In_1224,In_160);
or U413 (N_413,In_977,In_820);
nand U414 (N_414,In_1044,In_55);
nand U415 (N_415,In_1278,In_785);
nor U416 (N_416,In_843,In_120);
nand U417 (N_417,In_894,In_953);
and U418 (N_418,In_284,In_451);
or U419 (N_419,In_279,In_531);
nor U420 (N_420,In_1013,In_1408);
and U421 (N_421,In_1302,In_62);
nand U422 (N_422,In_637,In_356);
or U423 (N_423,In_1457,In_457);
nor U424 (N_424,In_933,In_812);
or U425 (N_425,In_1179,In_385);
or U426 (N_426,In_414,In_900);
xnor U427 (N_427,In_1089,In_1036);
nand U428 (N_428,In_1479,In_1338);
or U429 (N_429,In_235,In_1016);
nand U430 (N_430,In_1319,In_662);
and U431 (N_431,In_1051,In_388);
and U432 (N_432,In_730,In_552);
nor U433 (N_433,In_902,In_916);
nor U434 (N_434,In_1245,In_1439);
nor U435 (N_435,In_213,In_1410);
and U436 (N_436,In_253,In_946);
and U437 (N_437,In_106,In_810);
or U438 (N_438,In_1177,In_571);
nand U439 (N_439,In_882,In_506);
nor U440 (N_440,In_361,In_1025);
nor U441 (N_441,In_983,In_444);
nand U442 (N_442,In_1424,In_621);
nand U443 (N_443,In_1220,In_1352);
and U444 (N_444,In_1181,In_1454);
nor U445 (N_445,In_524,In_542);
xor U446 (N_446,In_23,In_744);
xnor U447 (N_447,In_254,In_762);
and U448 (N_448,In_1458,In_1009);
xor U449 (N_449,In_1236,In_604);
nand U450 (N_450,In_976,In_1070);
nand U451 (N_451,In_1317,In_614);
nand U452 (N_452,In_608,In_1350);
xnor U453 (N_453,In_1170,In_328);
and U454 (N_454,In_38,In_1230);
nor U455 (N_455,In_1413,In_972);
nand U456 (N_456,In_1305,In_553);
and U457 (N_457,In_364,In_1215);
nand U458 (N_458,In_484,In_78);
and U459 (N_459,In_1340,In_1308);
nor U460 (N_460,In_975,In_265);
and U461 (N_461,In_143,In_170);
and U462 (N_462,In_2,In_989);
nor U463 (N_463,In_59,In_1234);
or U464 (N_464,In_957,In_624);
and U465 (N_465,In_754,In_1314);
and U466 (N_466,In_96,In_18);
nand U467 (N_467,In_1144,In_928);
and U468 (N_468,In_714,In_987);
nor U469 (N_469,In_713,In_1264);
nor U470 (N_470,In_1328,In_1429);
or U471 (N_471,In_158,In_1301);
and U472 (N_472,In_24,In_399);
and U473 (N_473,In_947,In_1238);
and U474 (N_474,In_386,In_557);
or U475 (N_475,In_401,In_102);
and U476 (N_476,In_276,In_1023);
nand U477 (N_477,In_606,In_922);
or U478 (N_478,In_879,In_620);
xnor U479 (N_479,In_709,In_296);
nand U480 (N_480,In_899,In_1483);
nand U481 (N_481,In_1312,In_832);
or U482 (N_482,In_150,In_921);
xnor U483 (N_483,In_234,In_564);
and U484 (N_484,In_10,In_1335);
xnor U485 (N_485,In_971,In_819);
nand U486 (N_486,In_135,In_350);
and U487 (N_487,In_1040,In_1159);
nand U488 (N_488,In_433,In_1071);
or U489 (N_489,In_261,In_885);
nor U490 (N_490,In_224,In_969);
and U491 (N_491,In_634,In_771);
or U492 (N_492,In_280,In_82);
nand U493 (N_493,In_1091,In_781);
and U494 (N_494,In_1140,In_1001);
and U495 (N_495,In_1219,In_931);
or U496 (N_496,In_1239,In_365);
nor U497 (N_497,In_904,In_632);
or U498 (N_498,In_200,In_1098);
nor U499 (N_499,In_1086,In_511);
nor U500 (N_500,In_1370,In_543);
and U501 (N_501,In_1014,In_162);
nand U502 (N_502,In_389,In_930);
nand U503 (N_503,In_450,In_1194);
nor U504 (N_504,In_890,In_1342);
or U505 (N_505,In_202,In_1053);
nand U506 (N_506,In_1420,In_804);
nor U507 (N_507,In_1103,In_998);
nor U508 (N_508,In_1226,In_801);
nand U509 (N_509,In_784,In_1163);
or U510 (N_510,In_980,In_1283);
or U511 (N_511,In_1092,In_290);
nand U512 (N_512,In_39,In_241);
and U513 (N_513,In_337,In_952);
nor U514 (N_514,In_1192,In_1481);
nand U515 (N_515,In_186,In_699);
nor U516 (N_516,In_670,In_603);
nor U517 (N_517,In_45,In_272);
nand U518 (N_518,In_452,In_119);
nand U519 (N_519,In_1225,In_1259);
and U520 (N_520,In_226,In_1213);
and U521 (N_521,In_880,In_74);
xnor U522 (N_522,In_127,In_0);
nor U523 (N_523,In_1049,In_858);
nor U524 (N_524,In_722,In_988);
or U525 (N_525,In_1262,In_1263);
nor U526 (N_526,In_194,In_751);
or U527 (N_527,In_973,In_465);
xnor U528 (N_528,In_1162,In_789);
nand U529 (N_529,In_49,In_1157);
or U530 (N_530,In_540,In_220);
xor U531 (N_531,In_1321,In_425);
nor U532 (N_532,In_1315,In_1402);
and U533 (N_533,In_1391,In_1372);
nand U534 (N_534,In_270,In_1465);
xnor U535 (N_535,In_887,In_319);
nand U536 (N_536,In_132,In_1110);
xor U537 (N_537,In_79,In_943);
and U538 (N_538,In_1281,In_1376);
or U539 (N_539,In_736,In_697);
and U540 (N_540,In_1109,In_803);
or U541 (N_541,In_1453,In_574);
and U542 (N_542,In_440,In_750);
or U543 (N_543,In_926,In_979);
nand U544 (N_544,In_1452,In_1123);
nand U545 (N_545,In_1058,In_227);
nand U546 (N_546,In_1191,In_654);
or U547 (N_547,In_1347,In_442);
xor U548 (N_548,In_69,In_834);
xnor U549 (N_549,In_371,In_659);
and U550 (N_550,In_1249,In_91);
and U551 (N_551,In_1412,In_822);
nand U552 (N_552,In_746,In_665);
and U553 (N_553,In_827,In_757);
and U554 (N_554,In_825,In_182);
or U555 (N_555,In_378,In_297);
nor U556 (N_556,In_865,In_166);
or U557 (N_557,In_391,In_1105);
and U558 (N_558,In_1118,In_15);
nand U559 (N_559,In_510,In_1228);
nor U560 (N_560,In_172,In_741);
nand U561 (N_561,In_1440,In_83);
and U562 (N_562,In_81,In_698);
nor U563 (N_563,In_1449,In_924);
nand U564 (N_564,In_1108,In_568);
or U565 (N_565,In_435,In_114);
nand U566 (N_566,In_1406,In_1197);
or U567 (N_567,In_476,In_991);
nor U568 (N_568,In_489,In_914);
xor U569 (N_569,In_294,In_1295);
or U570 (N_570,In_1168,In_1247);
xnor U571 (N_571,In_1182,In_1487);
nand U572 (N_572,In_349,In_1351);
nor U573 (N_573,In_647,In_338);
and U574 (N_574,In_876,In_955);
and U575 (N_575,In_144,In_1169);
nand U576 (N_576,In_570,In_1421);
and U577 (N_577,In_643,In_1214);
nor U578 (N_578,In_872,In_503);
and U579 (N_579,In_376,In_1437);
nor U580 (N_580,In_393,In_247);
nand U581 (N_581,In_252,In_311);
nor U582 (N_582,In_354,In_462);
nor U583 (N_583,In_830,In_118);
nor U584 (N_584,In_629,In_1461);
and U585 (N_585,In_1002,In_113);
nor U586 (N_586,In_1227,In_646);
xnor U587 (N_587,In_321,In_408);
xor U588 (N_588,In_792,In_1422);
nand U589 (N_589,In_1332,In_384);
nand U590 (N_590,In_244,In_985);
and U591 (N_591,In_633,In_1010);
and U592 (N_592,In_466,In_415);
and U593 (N_593,In_1432,In_147);
and U594 (N_594,In_996,In_1084);
nand U595 (N_595,In_766,In_1161);
and U596 (N_596,In_1265,In_1136);
or U597 (N_597,In_1095,In_1493);
xnor U598 (N_598,In_826,In_1499);
nor U599 (N_599,In_1382,In_109);
and U600 (N_600,In_4,In_877);
nor U601 (N_601,In_537,In_962);
nand U602 (N_602,In_704,In_777);
nand U603 (N_603,In_1021,In_286);
nor U604 (N_604,In_1241,In_1298);
nor U605 (N_605,In_1396,In_300);
nand U606 (N_606,In_1411,In_993);
nor U607 (N_607,In_716,In_203);
nand U608 (N_608,In_108,In_86);
nor U609 (N_609,In_345,In_1047);
nand U610 (N_610,In_724,In_888);
or U611 (N_611,In_610,In_1339);
and U612 (N_612,In_563,In_1445);
and U613 (N_613,In_1011,In_1403);
or U614 (N_614,In_134,In_167);
nor U615 (N_615,In_330,In_481);
nand U616 (N_616,In_554,In_25);
nand U617 (N_617,In_748,In_439);
or U618 (N_618,In_715,In_548);
nand U619 (N_619,In_424,In_231);
nor U620 (N_620,In_44,In_1373);
xnor U621 (N_621,In_171,In_1271);
xor U622 (N_622,In_859,In_1028);
or U623 (N_623,In_1246,In_1415);
and U624 (N_624,In_534,In_1007);
and U625 (N_625,In_630,In_431);
nor U626 (N_626,In_20,In_811);
and U627 (N_627,In_242,In_978);
nor U628 (N_628,In_1232,In_745);
or U629 (N_629,In_1353,In_615);
and U630 (N_630,In_519,In_1468);
and U631 (N_631,In_458,In_293);
nand U632 (N_632,In_123,In_609);
and U633 (N_633,In_359,In_310);
or U634 (N_634,In_1124,In_1313);
nor U635 (N_635,In_392,In_1212);
nor U636 (N_636,In_314,In_223);
nand U637 (N_637,In_749,In_214);
and U638 (N_638,In_707,In_649);
nor U639 (N_639,In_776,In_84);
nand U640 (N_640,In_315,In_1293);
or U641 (N_641,In_626,In_681);
and U642 (N_642,In_1030,In_1167);
and U643 (N_643,In_589,In_1061);
and U644 (N_644,In_690,In_508);
or U645 (N_645,In_1388,In_448);
and U646 (N_646,In_245,In_873);
nor U647 (N_647,In_1456,In_287);
nor U648 (N_648,In_443,In_915);
nor U649 (N_649,In_196,In_1385);
nand U650 (N_650,In_222,In_831);
nand U651 (N_651,In_1292,In_968);
and U652 (N_652,In_1392,In_849);
and U653 (N_653,In_964,In_493);
or U654 (N_654,In_779,In_1374);
or U655 (N_655,In_92,In_932);
nand U656 (N_656,In_1054,In_400);
and U657 (N_657,In_1251,In_773);
or U658 (N_658,In_1218,In_1068);
nand U659 (N_659,In_281,In_375);
xnor U660 (N_660,In_1066,In_1034);
or U661 (N_661,In_1131,In_1067);
or U662 (N_662,In_430,In_1345);
nand U663 (N_663,In_173,In_318);
nor U664 (N_664,In_165,In_824);
and U665 (N_665,In_1470,In_852);
and U666 (N_666,In_1125,In_838);
nand U667 (N_667,In_1233,In_1113);
nand U668 (N_668,In_687,In_188);
nand U669 (N_669,In_528,In_1325);
or U670 (N_670,In_774,In_351);
and U671 (N_671,In_492,In_992);
nor U672 (N_672,In_532,In_67);
and U673 (N_673,In_1041,In_1269);
nand U674 (N_674,In_1359,In_1115);
or U675 (N_675,In_517,In_1446);
and U676 (N_676,In_529,In_1448);
nor U677 (N_677,In_674,In_340);
nor U678 (N_678,In_185,In_1165);
nor U679 (N_679,In_117,In_198);
xor U680 (N_680,In_1394,In_1363);
nor U681 (N_681,In_791,In_780);
nand U682 (N_682,In_416,In_1438);
nand U683 (N_683,In_65,In_409);
and U684 (N_684,In_954,In_148);
and U685 (N_685,In_845,In_578);
xor U686 (N_686,In_981,In_841);
nand U687 (N_687,In_1427,In_686);
or U688 (N_688,In_912,In_1311);
and U689 (N_689,In_30,In_1368);
or U690 (N_690,In_1183,In_733);
xor U691 (N_691,In_759,In_1077);
nand U692 (N_692,In_47,In_53);
nand U693 (N_693,In_72,In_1080);
nand U694 (N_694,In_889,In_1401);
nor U695 (N_695,In_518,In_1114);
xor U696 (N_696,In_657,In_1130);
nand U697 (N_697,In_625,In_419);
xor U698 (N_698,In_111,In_137);
nor U699 (N_699,In_586,In_734);
or U700 (N_700,In_1297,In_208);
and U701 (N_701,In_935,In_274);
nor U702 (N_702,In_809,In_1101);
or U703 (N_703,In_145,In_1436);
nor U704 (N_704,In_152,In_428);
nand U705 (N_705,In_434,In_1158);
and U706 (N_706,In_612,In_498);
and U707 (N_707,In_1291,In_1081);
and U708 (N_708,In_1296,In_731);
and U709 (N_709,In_1185,In_497);
nand U710 (N_710,In_1444,In_919);
nor U711 (N_711,In_266,In_1237);
nand U712 (N_712,In_1088,In_1303);
nand U713 (N_713,In_1178,In_818);
nand U714 (N_714,In_1097,In_1104);
nand U715 (N_715,In_1390,In_587);
nor U716 (N_716,In_1447,In_541);
nor U717 (N_717,In_1175,In_341);
and U718 (N_718,In_322,In_1082);
or U719 (N_719,In_7,In_93);
and U720 (N_720,In_1190,In_856);
nand U721 (N_721,In_669,In_861);
or U722 (N_722,In_22,In_918);
or U723 (N_723,In_729,In_897);
and U724 (N_724,In_339,In_195);
xor U725 (N_725,In_658,In_1069);
or U726 (N_726,In_680,In_1062);
nand U727 (N_727,In_1154,In_653);
nand U728 (N_728,In_1423,In_837);
nand U729 (N_729,In_1433,In_128);
or U730 (N_730,In_240,In_1306);
and U731 (N_731,In_622,In_577);
or U732 (N_732,In_1064,In_1072);
nor U733 (N_733,In_70,In_948);
xor U734 (N_734,In_1409,In_833);
nand U735 (N_735,In_688,In_1012);
and U736 (N_736,In_360,In_1484);
xnor U737 (N_737,In_1357,In_523);
nand U738 (N_738,In_1042,In_1019);
nor U739 (N_739,In_229,In_547);
or U740 (N_740,In_138,In_786);
or U741 (N_741,In_585,In_641);
or U742 (N_742,In_576,In_664);
nor U743 (N_743,In_512,In_16);
and U744 (N_744,In_331,In_1050);
and U745 (N_745,In_886,In_671);
and U746 (N_746,In_867,In_1208);
nor U747 (N_747,In_1331,In_1003);
nor U748 (N_748,In_747,In_309);
nor U749 (N_749,In_373,In_205);
and U750 (N_750,N_319,N_596);
nand U751 (N_751,N_720,N_456);
nand U752 (N_752,N_45,N_725);
or U753 (N_753,N_369,N_736);
nor U754 (N_754,N_461,N_642);
or U755 (N_755,N_395,N_215);
nor U756 (N_756,N_411,N_353);
nor U757 (N_757,N_171,N_93);
or U758 (N_758,N_740,N_714);
nand U759 (N_759,N_376,N_143);
nand U760 (N_760,N_123,N_420);
nand U761 (N_761,N_646,N_57);
nand U762 (N_762,N_622,N_8);
and U763 (N_763,N_523,N_28);
or U764 (N_764,N_298,N_721);
nor U765 (N_765,N_628,N_127);
or U766 (N_766,N_405,N_426);
or U767 (N_767,N_675,N_626);
xor U768 (N_768,N_739,N_193);
nand U769 (N_769,N_368,N_149);
nor U770 (N_770,N_67,N_110);
or U771 (N_771,N_292,N_272);
or U772 (N_772,N_727,N_643);
nand U773 (N_773,N_489,N_185);
nand U774 (N_774,N_683,N_423);
nor U775 (N_775,N_65,N_109);
or U776 (N_776,N_696,N_301);
nor U777 (N_777,N_283,N_222);
nor U778 (N_778,N_705,N_55);
and U779 (N_779,N_595,N_354);
and U780 (N_780,N_158,N_464);
nand U781 (N_781,N_673,N_713);
and U782 (N_782,N_364,N_553);
and U783 (N_783,N_620,N_113);
and U784 (N_784,N_180,N_413);
and U785 (N_785,N_446,N_733);
and U786 (N_786,N_359,N_470);
and U787 (N_787,N_666,N_617);
nor U788 (N_788,N_314,N_267);
and U789 (N_789,N_308,N_73);
nor U790 (N_790,N_380,N_138);
nor U791 (N_791,N_178,N_650);
nor U792 (N_792,N_521,N_281);
nor U793 (N_793,N_150,N_517);
and U794 (N_794,N_414,N_291);
nor U795 (N_795,N_707,N_384);
nand U796 (N_796,N_391,N_716);
nand U797 (N_797,N_657,N_124);
and U798 (N_798,N_318,N_460);
and U799 (N_799,N_410,N_174);
nor U800 (N_800,N_102,N_355);
and U801 (N_801,N_88,N_35);
nor U802 (N_802,N_40,N_605);
and U803 (N_803,N_552,N_522);
or U804 (N_804,N_94,N_60);
and U805 (N_805,N_285,N_336);
or U806 (N_806,N_609,N_462);
and U807 (N_807,N_545,N_579);
nor U808 (N_808,N_341,N_220);
xor U809 (N_809,N_76,N_170);
nand U810 (N_810,N_307,N_234);
nor U811 (N_811,N_106,N_10);
nand U812 (N_812,N_404,N_156);
xor U813 (N_813,N_242,N_483);
or U814 (N_814,N_197,N_644);
nand U815 (N_815,N_566,N_616);
and U816 (N_816,N_477,N_358);
nand U817 (N_817,N_23,N_257);
or U818 (N_818,N_655,N_131);
and U819 (N_819,N_322,N_196);
nor U820 (N_820,N_256,N_735);
or U821 (N_821,N_70,N_402);
nand U822 (N_822,N_651,N_61);
nand U823 (N_823,N_310,N_16);
xnor U824 (N_824,N_636,N_79);
nor U825 (N_825,N_603,N_315);
and U826 (N_826,N_611,N_352);
nand U827 (N_827,N_224,N_181);
xor U828 (N_828,N_134,N_248);
nor U829 (N_829,N_87,N_249);
or U830 (N_830,N_250,N_290);
and U831 (N_831,N_621,N_253);
nor U832 (N_832,N_370,N_530);
and U833 (N_833,N_533,N_348);
or U834 (N_834,N_154,N_419);
nand U835 (N_835,N_279,N_639);
or U836 (N_836,N_678,N_31);
or U837 (N_837,N_345,N_371);
and U838 (N_838,N_120,N_610);
nor U839 (N_839,N_490,N_440);
and U840 (N_840,N_510,N_367);
or U841 (N_841,N_518,N_274);
and U842 (N_842,N_12,N_471);
nor U843 (N_843,N_38,N_670);
or U844 (N_844,N_11,N_209);
nor U845 (N_845,N_577,N_416);
xnor U846 (N_846,N_656,N_407);
or U847 (N_847,N_722,N_165);
or U848 (N_848,N_488,N_64);
nor U849 (N_849,N_732,N_571);
nor U850 (N_850,N_211,N_9);
or U851 (N_851,N_572,N_326);
nor U852 (N_852,N_205,N_637);
or U853 (N_853,N_737,N_155);
or U854 (N_854,N_235,N_241);
or U855 (N_855,N_260,N_288);
nor U856 (N_856,N_647,N_560);
or U857 (N_857,N_382,N_32);
or U858 (N_858,N_672,N_115);
nand U859 (N_859,N_406,N_700);
nand U860 (N_860,N_112,N_748);
and U861 (N_861,N_467,N_17);
or U862 (N_862,N_468,N_728);
and U863 (N_863,N_543,N_432);
and U864 (N_864,N_693,N_484);
xor U865 (N_865,N_339,N_633);
or U866 (N_866,N_320,N_41);
and U867 (N_867,N_428,N_598);
nor U868 (N_868,N_259,N_195);
nor U869 (N_869,N_337,N_689);
nand U870 (N_870,N_625,N_329);
nand U871 (N_871,N_738,N_50);
or U872 (N_872,N_328,N_677);
nand U873 (N_873,N_627,N_581);
nor U874 (N_874,N_590,N_424);
or U875 (N_875,N_648,N_239);
nand U876 (N_876,N_258,N_383);
or U877 (N_877,N_442,N_140);
and U878 (N_878,N_303,N_293);
or U879 (N_879,N_679,N_100);
or U880 (N_880,N_139,N_47);
xnor U881 (N_881,N_589,N_487);
nor U882 (N_882,N_569,N_389);
nand U883 (N_883,N_187,N_379);
or U884 (N_884,N_403,N_494);
or U885 (N_885,N_172,N_325);
xnor U886 (N_886,N_731,N_434);
or U887 (N_887,N_63,N_323);
and U888 (N_888,N_27,N_481);
nor U889 (N_889,N_708,N_438);
nor U890 (N_890,N_210,N_575);
or U891 (N_891,N_694,N_82);
or U892 (N_892,N_527,N_444);
nor U893 (N_893,N_271,N_166);
or U894 (N_894,N_128,N_742);
nand U895 (N_895,N_299,N_218);
nand U896 (N_896,N_486,N_321);
or U897 (N_897,N_167,N_624);
xor U898 (N_898,N_231,N_591);
xnor U899 (N_899,N_316,N_48);
nor U900 (N_900,N_294,N_556);
nor U901 (N_901,N_480,N_671);
nand U902 (N_902,N_709,N_13);
nor U903 (N_903,N_711,N_300);
nand U904 (N_904,N_664,N_525);
or U905 (N_905,N_573,N_85);
xor U906 (N_906,N_629,N_511);
nor U907 (N_907,N_287,N_587);
or U908 (N_908,N_344,N_472);
xnor U909 (N_909,N_394,N_365);
and U910 (N_910,N_302,N_743);
xor U911 (N_911,N_493,N_619);
and U912 (N_912,N_505,N_561);
and U913 (N_913,N_295,N_546);
nor U914 (N_914,N_531,N_331);
nor U915 (N_915,N_284,N_529);
nor U916 (N_916,N_179,N_532);
or U917 (N_917,N_544,N_396);
and U918 (N_918,N_99,N_356);
nand U919 (N_919,N_238,N_507);
or U920 (N_920,N_135,N_433);
nand U921 (N_921,N_450,N_385);
and U922 (N_922,N_191,N_14);
nand U923 (N_923,N_439,N_96);
xor U924 (N_924,N_551,N_91);
nand U925 (N_925,N_681,N_72);
or U926 (N_926,N_608,N_719);
nor U927 (N_927,N_309,N_746);
nand U928 (N_928,N_363,N_496);
and U929 (N_929,N_607,N_111);
and U930 (N_930,N_421,N_216);
nand U931 (N_931,N_597,N_482);
nor U932 (N_932,N_706,N_223);
nor U933 (N_933,N_126,N_334);
nand U934 (N_934,N_540,N_116);
and U935 (N_935,N_199,N_710);
nor U936 (N_936,N_520,N_19);
or U937 (N_937,N_661,N_66);
or U938 (N_938,N_554,N_375);
nand U939 (N_939,N_244,N_233);
xnor U940 (N_940,N_262,N_152);
or U941 (N_941,N_567,N_588);
nand U942 (N_942,N_297,N_212);
nor U943 (N_943,N_21,N_491);
or U944 (N_944,N_125,N_599);
nor U945 (N_945,N_278,N_631);
and U946 (N_946,N_660,N_270);
xor U947 (N_947,N_208,N_43);
and U948 (N_948,N_680,N_362);
nor U949 (N_949,N_600,N_687);
nand U950 (N_950,N_653,N_665);
or U951 (N_951,N_3,N_228);
or U952 (N_952,N_652,N_275);
xor U953 (N_953,N_243,N_397);
and U954 (N_954,N_0,N_401);
nand U955 (N_955,N_347,N_269);
nor U956 (N_956,N_221,N_534);
nor U957 (N_957,N_519,N_332);
or U958 (N_958,N_632,N_236);
and U959 (N_959,N_24,N_176);
nor U960 (N_960,N_726,N_500);
or U961 (N_961,N_549,N_718);
xnor U962 (N_962,N_141,N_667);
nor U963 (N_963,N_747,N_701);
and U964 (N_964,N_557,N_312);
nand U965 (N_965,N_18,N_92);
or U966 (N_966,N_502,N_695);
or U967 (N_967,N_219,N_492);
nand U968 (N_968,N_475,N_53);
nand U969 (N_969,N_559,N_251);
nor U970 (N_970,N_390,N_463);
and U971 (N_971,N_654,N_688);
nor U972 (N_972,N_90,N_340);
nand U973 (N_973,N_697,N_684);
nand U974 (N_974,N_184,N_422);
nand U975 (N_975,N_466,N_430);
and U976 (N_976,N_506,N_604);
or U977 (N_977,N_311,N_36);
nor U978 (N_978,N_641,N_451);
nand U979 (N_979,N_198,N_441);
or U980 (N_980,N_137,N_330);
or U981 (N_981,N_144,N_59);
or U982 (N_982,N_49,N_454);
nand U983 (N_983,N_161,N_202);
or U984 (N_984,N_188,N_204);
xnor U985 (N_985,N_246,N_22);
nand U986 (N_986,N_415,N_190);
or U987 (N_987,N_514,N_564);
nand U988 (N_988,N_459,N_634);
nand U989 (N_989,N_495,N_485);
nor U990 (N_990,N_458,N_75);
nor U991 (N_991,N_372,N_240);
nand U992 (N_992,N_717,N_277);
nor U993 (N_993,N_412,N_227);
nand U994 (N_994,N_431,N_437);
or U995 (N_995,N_592,N_305);
nor U996 (N_996,N_715,N_338);
nor U997 (N_997,N_6,N_175);
xor U998 (N_998,N_162,N_173);
nor U999 (N_999,N_255,N_163);
nor U1000 (N_1000,N_547,N_498);
xor U1001 (N_1001,N_584,N_663);
nand U1002 (N_1002,N_388,N_427);
xor U1003 (N_1003,N_669,N_445);
and U1004 (N_1004,N_712,N_1);
and U1005 (N_1005,N_89,N_145);
xor U1006 (N_1006,N_304,N_563);
or U1007 (N_1007,N_261,N_606);
and U1008 (N_1008,N_528,N_474);
or U1009 (N_1009,N_457,N_536);
nor U1010 (N_1010,N_465,N_214);
or U1011 (N_1011,N_392,N_5);
or U1012 (N_1012,N_30,N_130);
nand U1013 (N_1013,N_381,N_132);
or U1014 (N_1014,N_15,N_576);
and U1015 (N_1015,N_108,N_263);
and U1016 (N_1016,N_698,N_133);
or U1017 (N_1017,N_105,N_95);
and U1018 (N_1018,N_515,N_741);
or U1019 (N_1019,N_393,N_366);
xor U1020 (N_1020,N_585,N_668);
nor U1021 (N_1021,N_229,N_62);
nand U1022 (N_1022,N_51,N_296);
nand U1023 (N_1023,N_97,N_455);
and U1024 (N_1024,N_418,N_729);
nor U1025 (N_1025,N_582,N_586);
nor U1026 (N_1026,N_453,N_583);
nand U1027 (N_1027,N_26,N_226);
or U1028 (N_1028,N_542,N_476);
nor U1029 (N_1029,N_509,N_74);
nor U1030 (N_1030,N_33,N_730);
nand U1031 (N_1031,N_245,N_452);
or U1032 (N_1032,N_645,N_623);
or U1033 (N_1033,N_317,N_266);
and U1034 (N_1034,N_479,N_101);
and U1035 (N_1035,N_435,N_734);
nand U1036 (N_1036,N_699,N_377);
xor U1037 (N_1037,N_192,N_146);
nor U1038 (N_1038,N_56,N_703);
nand U1039 (N_1039,N_268,N_638);
or U1040 (N_1040,N_225,N_58);
nor U1041 (N_1041,N_54,N_335);
and U1042 (N_1042,N_409,N_548);
nor U1043 (N_1043,N_98,N_103);
nor U1044 (N_1044,N_513,N_449);
and U1045 (N_1045,N_7,N_114);
nor U1046 (N_1046,N_568,N_447);
and U1047 (N_1047,N_349,N_230);
nand U1048 (N_1048,N_203,N_524);
nand U1049 (N_1049,N_682,N_39);
or U1050 (N_1050,N_52,N_252);
and U1051 (N_1051,N_723,N_237);
or U1052 (N_1052,N_744,N_538);
nor U1053 (N_1053,N_136,N_151);
nor U1054 (N_1054,N_286,N_118);
nor U1055 (N_1055,N_207,N_399);
or U1056 (N_1056,N_280,N_408);
nand U1057 (N_1057,N_189,N_350);
nand U1058 (N_1058,N_34,N_749);
xor U1059 (N_1059,N_386,N_541);
nand U1060 (N_1060,N_473,N_273);
and U1061 (N_1061,N_232,N_550);
nand U1062 (N_1062,N_374,N_247);
nand U1063 (N_1063,N_46,N_69);
and U1064 (N_1064,N_289,N_429);
xor U1065 (N_1065,N_276,N_122);
xor U1066 (N_1066,N_20,N_612);
xnor U1067 (N_1067,N_360,N_177);
xnor U1068 (N_1068,N_674,N_614);
or U1069 (N_1069,N_640,N_618);
xnor U1070 (N_1070,N_142,N_745);
or U1071 (N_1071,N_2,N_44);
nor U1072 (N_1072,N_217,N_690);
nor U1073 (N_1073,N_685,N_168);
nand U1074 (N_1074,N_508,N_264);
xor U1075 (N_1075,N_265,N_686);
or U1076 (N_1076,N_539,N_164);
or U1077 (N_1077,N_148,N_562);
and U1078 (N_1078,N_565,N_121);
and U1079 (N_1079,N_346,N_201);
nand U1080 (N_1080,N_448,N_558);
and U1081 (N_1081,N_37,N_324);
or U1082 (N_1082,N_516,N_83);
or U1083 (N_1083,N_692,N_29);
nor U1084 (N_1084,N_501,N_206);
nand U1085 (N_1085,N_186,N_81);
or U1086 (N_1086,N_659,N_400);
or U1087 (N_1087,N_436,N_361);
and U1088 (N_1088,N_662,N_306);
or U1089 (N_1089,N_387,N_25);
nor U1090 (N_1090,N_613,N_594);
nand U1091 (N_1091,N_71,N_84);
nand U1092 (N_1092,N_537,N_555);
or U1093 (N_1093,N_4,N_649);
and U1094 (N_1094,N_159,N_602);
xor U1095 (N_1095,N_342,N_443);
or U1096 (N_1096,N_601,N_119);
xor U1097 (N_1097,N_77,N_213);
or U1098 (N_1098,N_504,N_351);
nand U1099 (N_1099,N_86,N_478);
and U1100 (N_1100,N_704,N_147);
and U1101 (N_1101,N_499,N_182);
nor U1102 (N_1102,N_107,N_658);
nor U1103 (N_1103,N_157,N_570);
or U1104 (N_1104,N_635,N_327);
and U1105 (N_1105,N_282,N_68);
or U1106 (N_1106,N_343,N_357);
or U1107 (N_1107,N_702,N_169);
xnor U1108 (N_1108,N_42,N_160);
or U1109 (N_1109,N_526,N_615);
nor U1110 (N_1110,N_200,N_512);
nand U1111 (N_1111,N_574,N_593);
and U1112 (N_1112,N_183,N_497);
or U1113 (N_1113,N_630,N_80);
and U1114 (N_1114,N_580,N_104);
nand U1115 (N_1115,N_333,N_724);
nor U1116 (N_1116,N_469,N_373);
or U1117 (N_1117,N_378,N_535);
or U1118 (N_1118,N_117,N_425);
nand U1119 (N_1119,N_676,N_398);
nor U1120 (N_1120,N_503,N_691);
or U1121 (N_1121,N_153,N_129);
or U1122 (N_1122,N_78,N_254);
nand U1123 (N_1123,N_417,N_313);
nor U1124 (N_1124,N_194,N_578);
and U1125 (N_1125,N_709,N_745);
nand U1126 (N_1126,N_602,N_469);
and U1127 (N_1127,N_209,N_724);
xnor U1128 (N_1128,N_588,N_658);
and U1129 (N_1129,N_58,N_150);
and U1130 (N_1130,N_191,N_264);
nand U1131 (N_1131,N_331,N_728);
or U1132 (N_1132,N_386,N_517);
nor U1133 (N_1133,N_701,N_115);
nor U1134 (N_1134,N_125,N_78);
nor U1135 (N_1135,N_148,N_388);
nand U1136 (N_1136,N_68,N_338);
or U1137 (N_1137,N_142,N_42);
nand U1138 (N_1138,N_79,N_577);
or U1139 (N_1139,N_597,N_413);
nand U1140 (N_1140,N_742,N_255);
nand U1141 (N_1141,N_35,N_292);
and U1142 (N_1142,N_443,N_23);
or U1143 (N_1143,N_404,N_407);
xor U1144 (N_1144,N_235,N_93);
nor U1145 (N_1145,N_410,N_396);
xor U1146 (N_1146,N_571,N_299);
nand U1147 (N_1147,N_160,N_556);
nand U1148 (N_1148,N_416,N_546);
nand U1149 (N_1149,N_439,N_654);
xor U1150 (N_1150,N_221,N_306);
or U1151 (N_1151,N_656,N_273);
or U1152 (N_1152,N_16,N_34);
and U1153 (N_1153,N_111,N_4);
nor U1154 (N_1154,N_536,N_520);
and U1155 (N_1155,N_561,N_6);
and U1156 (N_1156,N_72,N_707);
and U1157 (N_1157,N_332,N_382);
or U1158 (N_1158,N_362,N_692);
and U1159 (N_1159,N_720,N_53);
xnor U1160 (N_1160,N_454,N_307);
or U1161 (N_1161,N_109,N_192);
and U1162 (N_1162,N_153,N_120);
and U1163 (N_1163,N_325,N_622);
and U1164 (N_1164,N_397,N_407);
xnor U1165 (N_1165,N_741,N_43);
nand U1166 (N_1166,N_110,N_631);
nor U1167 (N_1167,N_229,N_379);
nand U1168 (N_1168,N_325,N_304);
and U1169 (N_1169,N_17,N_18);
or U1170 (N_1170,N_8,N_435);
and U1171 (N_1171,N_384,N_256);
or U1172 (N_1172,N_536,N_260);
and U1173 (N_1173,N_631,N_630);
nand U1174 (N_1174,N_500,N_57);
or U1175 (N_1175,N_143,N_429);
nand U1176 (N_1176,N_247,N_19);
and U1177 (N_1177,N_172,N_171);
nand U1178 (N_1178,N_34,N_215);
nor U1179 (N_1179,N_104,N_36);
nand U1180 (N_1180,N_636,N_65);
nor U1181 (N_1181,N_716,N_184);
and U1182 (N_1182,N_15,N_218);
or U1183 (N_1183,N_414,N_250);
nand U1184 (N_1184,N_620,N_572);
nand U1185 (N_1185,N_740,N_539);
xnor U1186 (N_1186,N_248,N_51);
nand U1187 (N_1187,N_254,N_696);
nor U1188 (N_1188,N_601,N_484);
xor U1189 (N_1189,N_51,N_397);
nor U1190 (N_1190,N_540,N_276);
or U1191 (N_1191,N_165,N_135);
or U1192 (N_1192,N_493,N_288);
nand U1193 (N_1193,N_123,N_528);
xnor U1194 (N_1194,N_588,N_93);
nor U1195 (N_1195,N_58,N_153);
or U1196 (N_1196,N_202,N_731);
or U1197 (N_1197,N_19,N_673);
nor U1198 (N_1198,N_173,N_688);
nor U1199 (N_1199,N_692,N_89);
or U1200 (N_1200,N_671,N_212);
nand U1201 (N_1201,N_399,N_480);
and U1202 (N_1202,N_130,N_224);
xnor U1203 (N_1203,N_362,N_621);
nor U1204 (N_1204,N_14,N_110);
xor U1205 (N_1205,N_629,N_710);
or U1206 (N_1206,N_352,N_439);
nand U1207 (N_1207,N_603,N_566);
nand U1208 (N_1208,N_404,N_706);
nand U1209 (N_1209,N_391,N_362);
nor U1210 (N_1210,N_621,N_104);
or U1211 (N_1211,N_514,N_130);
nor U1212 (N_1212,N_428,N_527);
nand U1213 (N_1213,N_1,N_742);
nand U1214 (N_1214,N_662,N_243);
and U1215 (N_1215,N_484,N_26);
nor U1216 (N_1216,N_586,N_436);
nand U1217 (N_1217,N_730,N_550);
nor U1218 (N_1218,N_37,N_70);
nand U1219 (N_1219,N_457,N_648);
xnor U1220 (N_1220,N_200,N_10);
xor U1221 (N_1221,N_447,N_567);
nand U1222 (N_1222,N_180,N_743);
nand U1223 (N_1223,N_32,N_217);
or U1224 (N_1224,N_187,N_274);
xor U1225 (N_1225,N_434,N_9);
and U1226 (N_1226,N_279,N_135);
nand U1227 (N_1227,N_239,N_300);
or U1228 (N_1228,N_252,N_333);
nand U1229 (N_1229,N_529,N_589);
xnor U1230 (N_1230,N_100,N_720);
or U1231 (N_1231,N_617,N_747);
and U1232 (N_1232,N_114,N_110);
xnor U1233 (N_1233,N_216,N_618);
nand U1234 (N_1234,N_292,N_480);
nor U1235 (N_1235,N_56,N_683);
and U1236 (N_1236,N_726,N_74);
nor U1237 (N_1237,N_220,N_264);
nor U1238 (N_1238,N_398,N_456);
or U1239 (N_1239,N_574,N_33);
nand U1240 (N_1240,N_578,N_34);
nand U1241 (N_1241,N_578,N_172);
nor U1242 (N_1242,N_175,N_243);
nand U1243 (N_1243,N_167,N_397);
or U1244 (N_1244,N_31,N_511);
nand U1245 (N_1245,N_705,N_296);
or U1246 (N_1246,N_83,N_71);
nor U1247 (N_1247,N_137,N_295);
and U1248 (N_1248,N_561,N_583);
or U1249 (N_1249,N_60,N_208);
nand U1250 (N_1250,N_743,N_22);
nand U1251 (N_1251,N_170,N_421);
nor U1252 (N_1252,N_221,N_497);
and U1253 (N_1253,N_641,N_437);
nand U1254 (N_1254,N_273,N_727);
or U1255 (N_1255,N_510,N_362);
xnor U1256 (N_1256,N_702,N_67);
and U1257 (N_1257,N_417,N_335);
nor U1258 (N_1258,N_632,N_54);
nor U1259 (N_1259,N_524,N_448);
or U1260 (N_1260,N_555,N_67);
nor U1261 (N_1261,N_226,N_494);
and U1262 (N_1262,N_372,N_478);
or U1263 (N_1263,N_487,N_306);
nor U1264 (N_1264,N_360,N_359);
nor U1265 (N_1265,N_129,N_455);
or U1266 (N_1266,N_259,N_112);
nor U1267 (N_1267,N_508,N_588);
nand U1268 (N_1268,N_612,N_115);
nand U1269 (N_1269,N_83,N_119);
or U1270 (N_1270,N_276,N_434);
nor U1271 (N_1271,N_104,N_164);
nor U1272 (N_1272,N_317,N_596);
xnor U1273 (N_1273,N_452,N_550);
nor U1274 (N_1274,N_491,N_323);
or U1275 (N_1275,N_370,N_68);
nand U1276 (N_1276,N_533,N_747);
xor U1277 (N_1277,N_292,N_712);
nor U1278 (N_1278,N_202,N_64);
or U1279 (N_1279,N_127,N_183);
and U1280 (N_1280,N_36,N_715);
and U1281 (N_1281,N_551,N_514);
nand U1282 (N_1282,N_369,N_258);
nand U1283 (N_1283,N_698,N_101);
or U1284 (N_1284,N_429,N_540);
or U1285 (N_1285,N_555,N_433);
nor U1286 (N_1286,N_10,N_118);
or U1287 (N_1287,N_476,N_748);
nand U1288 (N_1288,N_596,N_249);
and U1289 (N_1289,N_484,N_582);
nor U1290 (N_1290,N_187,N_233);
and U1291 (N_1291,N_534,N_186);
nor U1292 (N_1292,N_374,N_664);
nor U1293 (N_1293,N_646,N_727);
or U1294 (N_1294,N_648,N_406);
nor U1295 (N_1295,N_721,N_576);
nand U1296 (N_1296,N_425,N_662);
or U1297 (N_1297,N_165,N_665);
and U1298 (N_1298,N_146,N_116);
and U1299 (N_1299,N_343,N_233);
or U1300 (N_1300,N_41,N_473);
nand U1301 (N_1301,N_106,N_40);
or U1302 (N_1302,N_356,N_273);
nand U1303 (N_1303,N_597,N_587);
nor U1304 (N_1304,N_698,N_272);
nor U1305 (N_1305,N_455,N_607);
and U1306 (N_1306,N_498,N_83);
and U1307 (N_1307,N_321,N_154);
nand U1308 (N_1308,N_576,N_401);
nand U1309 (N_1309,N_279,N_133);
and U1310 (N_1310,N_179,N_126);
nand U1311 (N_1311,N_476,N_694);
nor U1312 (N_1312,N_446,N_188);
and U1313 (N_1313,N_122,N_329);
nor U1314 (N_1314,N_679,N_241);
nand U1315 (N_1315,N_137,N_718);
nor U1316 (N_1316,N_110,N_188);
xor U1317 (N_1317,N_659,N_540);
or U1318 (N_1318,N_657,N_222);
and U1319 (N_1319,N_486,N_481);
nor U1320 (N_1320,N_597,N_107);
nor U1321 (N_1321,N_48,N_77);
nor U1322 (N_1322,N_356,N_678);
and U1323 (N_1323,N_252,N_150);
and U1324 (N_1324,N_686,N_491);
xor U1325 (N_1325,N_249,N_587);
nor U1326 (N_1326,N_416,N_11);
nand U1327 (N_1327,N_299,N_626);
and U1328 (N_1328,N_664,N_282);
and U1329 (N_1329,N_478,N_235);
and U1330 (N_1330,N_296,N_20);
or U1331 (N_1331,N_502,N_202);
nor U1332 (N_1332,N_294,N_161);
and U1333 (N_1333,N_720,N_79);
xnor U1334 (N_1334,N_283,N_594);
nand U1335 (N_1335,N_106,N_270);
nand U1336 (N_1336,N_229,N_49);
nor U1337 (N_1337,N_537,N_319);
and U1338 (N_1338,N_597,N_671);
nor U1339 (N_1339,N_238,N_690);
xnor U1340 (N_1340,N_730,N_198);
nand U1341 (N_1341,N_134,N_426);
and U1342 (N_1342,N_255,N_117);
or U1343 (N_1343,N_589,N_97);
nand U1344 (N_1344,N_493,N_10);
and U1345 (N_1345,N_707,N_393);
nor U1346 (N_1346,N_559,N_188);
nand U1347 (N_1347,N_547,N_308);
or U1348 (N_1348,N_200,N_360);
or U1349 (N_1349,N_592,N_69);
and U1350 (N_1350,N_289,N_651);
nand U1351 (N_1351,N_150,N_402);
or U1352 (N_1352,N_708,N_576);
nand U1353 (N_1353,N_678,N_270);
nand U1354 (N_1354,N_616,N_14);
and U1355 (N_1355,N_234,N_441);
nand U1356 (N_1356,N_739,N_205);
nand U1357 (N_1357,N_521,N_275);
nor U1358 (N_1358,N_604,N_550);
nor U1359 (N_1359,N_340,N_358);
nand U1360 (N_1360,N_749,N_462);
xor U1361 (N_1361,N_33,N_98);
xnor U1362 (N_1362,N_621,N_698);
nor U1363 (N_1363,N_740,N_147);
xnor U1364 (N_1364,N_56,N_636);
or U1365 (N_1365,N_305,N_746);
nor U1366 (N_1366,N_83,N_352);
or U1367 (N_1367,N_106,N_218);
or U1368 (N_1368,N_715,N_215);
or U1369 (N_1369,N_671,N_567);
or U1370 (N_1370,N_311,N_579);
or U1371 (N_1371,N_594,N_590);
nand U1372 (N_1372,N_70,N_626);
or U1373 (N_1373,N_124,N_625);
nor U1374 (N_1374,N_732,N_606);
nand U1375 (N_1375,N_5,N_662);
or U1376 (N_1376,N_736,N_558);
or U1377 (N_1377,N_30,N_133);
nand U1378 (N_1378,N_222,N_458);
or U1379 (N_1379,N_657,N_204);
or U1380 (N_1380,N_423,N_206);
and U1381 (N_1381,N_654,N_195);
xnor U1382 (N_1382,N_369,N_30);
and U1383 (N_1383,N_612,N_1);
nor U1384 (N_1384,N_685,N_329);
or U1385 (N_1385,N_450,N_506);
and U1386 (N_1386,N_674,N_542);
nor U1387 (N_1387,N_176,N_382);
and U1388 (N_1388,N_590,N_22);
and U1389 (N_1389,N_549,N_289);
nand U1390 (N_1390,N_259,N_534);
nor U1391 (N_1391,N_69,N_317);
and U1392 (N_1392,N_237,N_536);
and U1393 (N_1393,N_535,N_373);
nand U1394 (N_1394,N_550,N_493);
and U1395 (N_1395,N_65,N_56);
or U1396 (N_1396,N_491,N_409);
nand U1397 (N_1397,N_634,N_340);
xor U1398 (N_1398,N_619,N_674);
nor U1399 (N_1399,N_687,N_241);
or U1400 (N_1400,N_605,N_633);
nand U1401 (N_1401,N_573,N_684);
and U1402 (N_1402,N_199,N_444);
and U1403 (N_1403,N_399,N_388);
and U1404 (N_1404,N_666,N_713);
nor U1405 (N_1405,N_417,N_99);
xnor U1406 (N_1406,N_516,N_386);
nor U1407 (N_1407,N_315,N_4);
nor U1408 (N_1408,N_196,N_164);
and U1409 (N_1409,N_223,N_595);
or U1410 (N_1410,N_601,N_668);
or U1411 (N_1411,N_685,N_689);
nand U1412 (N_1412,N_206,N_301);
or U1413 (N_1413,N_624,N_137);
or U1414 (N_1414,N_648,N_35);
nand U1415 (N_1415,N_447,N_570);
nand U1416 (N_1416,N_49,N_704);
nand U1417 (N_1417,N_457,N_720);
nand U1418 (N_1418,N_574,N_592);
and U1419 (N_1419,N_728,N_549);
and U1420 (N_1420,N_110,N_392);
and U1421 (N_1421,N_409,N_505);
and U1422 (N_1422,N_678,N_486);
or U1423 (N_1423,N_661,N_214);
nand U1424 (N_1424,N_307,N_551);
and U1425 (N_1425,N_388,N_248);
nand U1426 (N_1426,N_368,N_43);
or U1427 (N_1427,N_264,N_307);
xor U1428 (N_1428,N_732,N_616);
and U1429 (N_1429,N_460,N_217);
xor U1430 (N_1430,N_53,N_91);
or U1431 (N_1431,N_473,N_594);
nand U1432 (N_1432,N_702,N_604);
xor U1433 (N_1433,N_316,N_287);
and U1434 (N_1434,N_604,N_575);
and U1435 (N_1435,N_642,N_551);
or U1436 (N_1436,N_335,N_207);
nor U1437 (N_1437,N_685,N_546);
or U1438 (N_1438,N_623,N_173);
or U1439 (N_1439,N_677,N_535);
and U1440 (N_1440,N_407,N_376);
nand U1441 (N_1441,N_182,N_527);
nor U1442 (N_1442,N_91,N_106);
nand U1443 (N_1443,N_505,N_520);
nor U1444 (N_1444,N_601,N_319);
and U1445 (N_1445,N_457,N_364);
nand U1446 (N_1446,N_95,N_102);
or U1447 (N_1447,N_744,N_195);
nand U1448 (N_1448,N_495,N_330);
nand U1449 (N_1449,N_485,N_606);
xnor U1450 (N_1450,N_281,N_5);
nand U1451 (N_1451,N_362,N_199);
nor U1452 (N_1452,N_387,N_86);
and U1453 (N_1453,N_306,N_713);
nand U1454 (N_1454,N_213,N_453);
or U1455 (N_1455,N_629,N_516);
or U1456 (N_1456,N_423,N_585);
nor U1457 (N_1457,N_702,N_355);
nor U1458 (N_1458,N_62,N_294);
nand U1459 (N_1459,N_18,N_87);
and U1460 (N_1460,N_454,N_46);
xnor U1461 (N_1461,N_5,N_291);
nor U1462 (N_1462,N_142,N_151);
and U1463 (N_1463,N_468,N_49);
or U1464 (N_1464,N_461,N_229);
nor U1465 (N_1465,N_604,N_602);
and U1466 (N_1466,N_147,N_198);
or U1467 (N_1467,N_229,N_343);
xnor U1468 (N_1468,N_88,N_276);
xnor U1469 (N_1469,N_483,N_633);
and U1470 (N_1470,N_128,N_400);
nor U1471 (N_1471,N_465,N_675);
nand U1472 (N_1472,N_87,N_95);
and U1473 (N_1473,N_284,N_438);
and U1474 (N_1474,N_72,N_557);
and U1475 (N_1475,N_229,N_20);
and U1476 (N_1476,N_575,N_151);
nor U1477 (N_1477,N_51,N_418);
or U1478 (N_1478,N_418,N_294);
and U1479 (N_1479,N_480,N_13);
nor U1480 (N_1480,N_668,N_545);
or U1481 (N_1481,N_214,N_191);
nor U1482 (N_1482,N_113,N_216);
or U1483 (N_1483,N_133,N_453);
nand U1484 (N_1484,N_60,N_51);
and U1485 (N_1485,N_486,N_129);
and U1486 (N_1486,N_576,N_709);
and U1487 (N_1487,N_342,N_146);
and U1488 (N_1488,N_702,N_662);
or U1489 (N_1489,N_593,N_101);
nor U1490 (N_1490,N_503,N_536);
nor U1491 (N_1491,N_222,N_169);
and U1492 (N_1492,N_665,N_109);
nor U1493 (N_1493,N_321,N_479);
xor U1494 (N_1494,N_255,N_339);
nand U1495 (N_1495,N_120,N_198);
nand U1496 (N_1496,N_109,N_721);
and U1497 (N_1497,N_270,N_519);
nand U1498 (N_1498,N_206,N_240);
or U1499 (N_1499,N_265,N_715);
and U1500 (N_1500,N_1152,N_993);
xor U1501 (N_1501,N_1024,N_780);
xor U1502 (N_1502,N_1224,N_1198);
xor U1503 (N_1503,N_1197,N_871);
nand U1504 (N_1504,N_791,N_1269);
or U1505 (N_1505,N_963,N_1079);
and U1506 (N_1506,N_992,N_1442);
and U1507 (N_1507,N_1389,N_1359);
or U1508 (N_1508,N_889,N_1218);
nand U1509 (N_1509,N_1363,N_950);
nor U1510 (N_1510,N_999,N_769);
or U1511 (N_1511,N_1025,N_1291);
nand U1512 (N_1512,N_1346,N_1320);
xor U1513 (N_1513,N_1114,N_899);
or U1514 (N_1514,N_954,N_1028);
and U1515 (N_1515,N_1158,N_1265);
nor U1516 (N_1516,N_1378,N_1102);
and U1517 (N_1517,N_1138,N_767);
or U1518 (N_1518,N_904,N_1487);
and U1519 (N_1519,N_805,N_924);
nor U1520 (N_1520,N_1264,N_1143);
and U1521 (N_1521,N_1271,N_1117);
and U1522 (N_1522,N_1154,N_1493);
and U1523 (N_1523,N_1282,N_1292);
nor U1524 (N_1524,N_1093,N_1407);
xnor U1525 (N_1525,N_1465,N_1182);
nand U1526 (N_1526,N_1202,N_1082);
nand U1527 (N_1527,N_793,N_1210);
nand U1528 (N_1528,N_857,N_1468);
nor U1529 (N_1529,N_1180,N_1009);
and U1530 (N_1530,N_1149,N_1023);
or U1531 (N_1531,N_808,N_1496);
or U1532 (N_1532,N_1075,N_949);
or U1533 (N_1533,N_1452,N_1344);
nor U1534 (N_1534,N_1020,N_1122);
or U1535 (N_1535,N_812,N_810);
nor U1536 (N_1536,N_896,N_1308);
or U1537 (N_1537,N_920,N_1053);
nand U1538 (N_1538,N_923,N_1206);
xor U1539 (N_1539,N_1064,N_1033);
xnor U1540 (N_1540,N_1228,N_875);
or U1541 (N_1541,N_1433,N_977);
and U1542 (N_1542,N_1425,N_960);
and U1543 (N_1543,N_1119,N_1044);
nand U1544 (N_1544,N_1034,N_955);
or U1545 (N_1545,N_909,N_1427);
and U1546 (N_1546,N_1065,N_1259);
xor U1547 (N_1547,N_1406,N_1343);
or U1548 (N_1548,N_1306,N_1051);
xor U1549 (N_1549,N_1032,N_1485);
nand U1550 (N_1550,N_892,N_1013);
nand U1551 (N_1551,N_1091,N_983);
xor U1552 (N_1552,N_801,N_1455);
nand U1553 (N_1553,N_1055,N_1109);
or U1554 (N_1554,N_1410,N_1043);
nor U1555 (N_1555,N_1123,N_1412);
nand U1556 (N_1556,N_1103,N_1021);
or U1557 (N_1557,N_879,N_1453);
and U1558 (N_1558,N_1225,N_1379);
nand U1559 (N_1559,N_867,N_1466);
xnor U1560 (N_1560,N_1337,N_1164);
or U1561 (N_1561,N_902,N_976);
xor U1562 (N_1562,N_989,N_1219);
and U1563 (N_1563,N_1071,N_1004);
and U1564 (N_1564,N_886,N_1112);
and U1565 (N_1565,N_1294,N_1173);
or U1566 (N_1566,N_1090,N_1480);
and U1567 (N_1567,N_1041,N_1003);
xor U1568 (N_1568,N_802,N_952);
xor U1569 (N_1569,N_1106,N_1200);
and U1570 (N_1570,N_1131,N_1335);
and U1571 (N_1571,N_1230,N_1481);
or U1572 (N_1572,N_1416,N_1369);
and U1573 (N_1573,N_1147,N_1247);
nand U1574 (N_1574,N_958,N_1145);
and U1575 (N_1575,N_1100,N_1423);
and U1576 (N_1576,N_990,N_1397);
nand U1577 (N_1577,N_824,N_794);
or U1578 (N_1578,N_1178,N_1139);
xor U1579 (N_1579,N_1323,N_1205);
xor U1580 (N_1580,N_1047,N_809);
nor U1581 (N_1581,N_1284,N_850);
and U1582 (N_1582,N_913,N_1495);
nand U1583 (N_1583,N_1234,N_760);
nor U1584 (N_1584,N_863,N_1263);
and U1585 (N_1585,N_1413,N_1017);
and U1586 (N_1586,N_1299,N_1007);
nand U1587 (N_1587,N_1048,N_1411);
nor U1588 (N_1588,N_925,N_798);
nand U1589 (N_1589,N_1362,N_1050);
and U1590 (N_1590,N_1080,N_1318);
or U1591 (N_1591,N_837,N_986);
nor U1592 (N_1592,N_1421,N_891);
and U1593 (N_1593,N_897,N_1222);
xor U1594 (N_1594,N_1054,N_817);
and U1595 (N_1595,N_1437,N_1087);
nand U1596 (N_1596,N_934,N_1332);
or U1597 (N_1597,N_1317,N_907);
nor U1598 (N_1598,N_1488,N_931);
and U1599 (N_1599,N_1078,N_1297);
xnor U1600 (N_1600,N_1108,N_1461);
nand U1601 (N_1601,N_750,N_1486);
xnor U1602 (N_1602,N_1333,N_1267);
or U1603 (N_1603,N_985,N_1430);
and U1604 (N_1604,N_1467,N_1236);
and U1605 (N_1605,N_888,N_1160);
nor U1606 (N_1606,N_858,N_1400);
nand U1607 (N_1607,N_1209,N_978);
xor U1608 (N_1608,N_1336,N_831);
and U1609 (N_1609,N_1376,N_1321);
and U1610 (N_1610,N_1287,N_1331);
xor U1611 (N_1611,N_1029,N_1185);
nor U1612 (N_1612,N_1440,N_796);
nor U1613 (N_1613,N_906,N_1128);
or U1614 (N_1614,N_773,N_1245);
and U1615 (N_1615,N_894,N_1240);
nor U1616 (N_1616,N_1310,N_938);
and U1617 (N_1617,N_765,N_1166);
or U1618 (N_1618,N_1221,N_1327);
nand U1619 (N_1619,N_1489,N_1303);
or U1620 (N_1620,N_1450,N_1449);
nand U1621 (N_1621,N_1364,N_865);
and U1622 (N_1622,N_1130,N_1268);
xor U1623 (N_1623,N_905,N_1010);
nor U1624 (N_1624,N_806,N_1027);
nor U1625 (N_1625,N_1001,N_1146);
and U1626 (N_1626,N_1329,N_1148);
nor U1627 (N_1627,N_873,N_1172);
nor U1628 (N_1628,N_820,N_755);
nand U1629 (N_1629,N_844,N_829);
or U1630 (N_1630,N_1005,N_1373);
or U1631 (N_1631,N_1115,N_1340);
and U1632 (N_1632,N_1042,N_1213);
or U1633 (N_1633,N_1249,N_1476);
nor U1634 (N_1634,N_1235,N_1127);
nor U1635 (N_1635,N_1399,N_1479);
nand U1636 (N_1636,N_1081,N_1351);
nand U1637 (N_1637,N_1260,N_1132);
and U1638 (N_1638,N_860,N_1133);
and U1639 (N_1639,N_1251,N_1286);
or U1640 (N_1640,N_781,N_1325);
nor U1641 (N_1641,N_987,N_1422);
nand U1642 (N_1642,N_821,N_1420);
nand U1643 (N_1643,N_935,N_1324);
or U1644 (N_1644,N_1285,N_1229);
and U1645 (N_1645,N_1445,N_1328);
nor U1646 (N_1646,N_1076,N_1295);
xnor U1647 (N_1647,N_1298,N_957);
and U1648 (N_1648,N_1176,N_1339);
nor U1649 (N_1649,N_973,N_1342);
xnor U1650 (N_1650,N_996,N_951);
or U1651 (N_1651,N_968,N_1444);
nor U1652 (N_1652,N_1434,N_834);
and U1653 (N_1653,N_1068,N_937);
nor U1654 (N_1654,N_842,N_1414);
or U1655 (N_1655,N_883,N_1107);
nor U1656 (N_1656,N_784,N_1385);
xnor U1657 (N_1657,N_1405,N_1223);
nor U1658 (N_1658,N_1375,N_1037);
and U1659 (N_1659,N_1384,N_856);
nand U1660 (N_1660,N_1409,N_1458);
nand U1661 (N_1661,N_1456,N_1426);
nor U1662 (N_1662,N_1401,N_882);
or U1663 (N_1663,N_1490,N_855);
and U1664 (N_1664,N_754,N_1239);
nor U1665 (N_1665,N_1367,N_921);
and U1666 (N_1666,N_1256,N_1386);
and U1667 (N_1667,N_1111,N_1261);
and U1668 (N_1668,N_911,N_1159);
or U1669 (N_1669,N_1242,N_1110);
nor U1670 (N_1670,N_1475,N_1377);
or U1671 (N_1671,N_1366,N_1454);
nand U1672 (N_1672,N_1214,N_1136);
nand U1673 (N_1673,N_1408,N_1459);
nand U1674 (N_1674,N_861,N_1276);
nand U1675 (N_1675,N_1305,N_940);
or U1676 (N_1676,N_851,N_1253);
nand U1677 (N_1677,N_1163,N_1365);
or U1678 (N_1678,N_1290,N_918);
or U1679 (N_1679,N_1443,N_759);
nand U1680 (N_1680,N_1330,N_1015);
nand U1681 (N_1681,N_964,N_1431);
xnor U1682 (N_1682,N_1415,N_971);
or U1683 (N_1683,N_1322,N_752);
nand U1684 (N_1684,N_947,N_1275);
nand U1685 (N_1685,N_982,N_1266);
nand U1686 (N_1686,N_1189,N_862);
and U1687 (N_1687,N_1302,N_1220);
nand U1688 (N_1688,N_1125,N_933);
nor U1689 (N_1689,N_1368,N_1199);
nand U1690 (N_1690,N_1462,N_941);
nand U1691 (N_1691,N_816,N_1313);
and U1692 (N_1692,N_1392,N_1135);
or U1693 (N_1693,N_1057,N_942);
and U1694 (N_1694,N_1066,N_813);
nand U1695 (N_1695,N_1341,N_811);
and U1696 (N_1696,N_870,N_853);
or U1697 (N_1697,N_1436,N_1097);
xor U1698 (N_1698,N_1073,N_803);
xor U1699 (N_1699,N_1250,N_1393);
nor U1700 (N_1700,N_1194,N_1049);
and U1701 (N_1701,N_770,N_1304);
and U1702 (N_1702,N_901,N_1204);
xor U1703 (N_1703,N_1216,N_1428);
or U1704 (N_1704,N_763,N_772);
and U1705 (N_1705,N_1226,N_916);
nor U1706 (N_1706,N_1498,N_864);
or U1707 (N_1707,N_1022,N_1390);
nor U1708 (N_1708,N_936,N_1244);
nor U1709 (N_1709,N_927,N_1432);
nand U1710 (N_1710,N_1491,N_764);
xnor U1711 (N_1711,N_1447,N_797);
and U1712 (N_1712,N_838,N_1274);
or U1713 (N_1713,N_1056,N_782);
and U1714 (N_1714,N_959,N_1012);
or U1715 (N_1715,N_1283,N_1246);
and U1716 (N_1716,N_1315,N_1120);
and U1717 (N_1717,N_1096,N_1312);
nor U1718 (N_1718,N_1077,N_975);
xnor U1719 (N_1719,N_1070,N_1035);
nand U1720 (N_1720,N_1060,N_756);
nor U1721 (N_1721,N_966,N_946);
xor U1722 (N_1722,N_1195,N_1349);
or U1723 (N_1723,N_1484,N_1497);
and U1724 (N_1724,N_910,N_1464);
or U1725 (N_1725,N_1374,N_914);
or U1726 (N_1726,N_827,N_1063);
and U1727 (N_1727,N_1179,N_1227);
or U1728 (N_1728,N_1355,N_1463);
xor U1729 (N_1729,N_792,N_859);
nor U1730 (N_1730,N_1208,N_1477);
nand U1731 (N_1731,N_1352,N_1254);
and U1732 (N_1732,N_790,N_1046);
xor U1733 (N_1733,N_783,N_893);
nor U1734 (N_1734,N_1086,N_1238);
and U1735 (N_1735,N_1347,N_945);
and U1736 (N_1736,N_1121,N_1356);
nand U1737 (N_1737,N_1045,N_1262);
nand U1738 (N_1738,N_930,N_1278);
and U1739 (N_1739,N_994,N_1277);
nand U1740 (N_1740,N_1129,N_1190);
xor U1741 (N_1741,N_1174,N_819);
or U1742 (N_1742,N_1289,N_887);
or U1743 (N_1743,N_1067,N_836);
and U1744 (N_1744,N_997,N_1248);
xnor U1745 (N_1745,N_1357,N_751);
and U1746 (N_1746,N_1191,N_854);
nor U1747 (N_1747,N_1232,N_1137);
and U1748 (N_1748,N_1473,N_1470);
or U1749 (N_1749,N_974,N_962);
nor U1750 (N_1750,N_1217,N_1417);
and U1751 (N_1751,N_1358,N_1101);
and U1752 (N_1752,N_1014,N_1175);
or U1753 (N_1753,N_815,N_972);
nor U1754 (N_1754,N_852,N_1058);
xnor U1755 (N_1755,N_1439,N_1059);
or U1756 (N_1756,N_1438,N_1288);
or U1757 (N_1757,N_1293,N_1441);
nor U1758 (N_1758,N_1429,N_1052);
or U1759 (N_1759,N_1492,N_1372);
nor U1760 (N_1760,N_1469,N_984);
nand U1761 (N_1761,N_1201,N_1168);
xnor U1762 (N_1762,N_1134,N_1124);
nand U1763 (N_1763,N_1074,N_1457);
nand U1764 (N_1764,N_832,N_1451);
xnor U1765 (N_1765,N_1167,N_762);
nand U1766 (N_1766,N_1171,N_1471);
xnor U1767 (N_1767,N_1231,N_915);
or U1768 (N_1768,N_1085,N_779);
xnor U1769 (N_1769,N_1169,N_1170);
xor U1770 (N_1770,N_1279,N_1398);
and U1771 (N_1771,N_1151,N_758);
or U1772 (N_1772,N_1088,N_768);
nand U1773 (N_1773,N_1104,N_1241);
and U1774 (N_1774,N_912,N_1006);
nand U1775 (N_1775,N_979,N_1144);
nor U1776 (N_1776,N_1150,N_1309);
nor U1777 (N_1777,N_1387,N_908);
and U1778 (N_1778,N_1403,N_1326);
or U1779 (N_1779,N_967,N_1162);
and U1780 (N_1780,N_1113,N_1192);
or U1781 (N_1781,N_866,N_1301);
nand U1782 (N_1782,N_1094,N_1038);
nand U1783 (N_1783,N_847,N_998);
or U1784 (N_1784,N_868,N_1370);
nand U1785 (N_1785,N_789,N_953);
nor U1786 (N_1786,N_1116,N_1435);
xor U1787 (N_1787,N_799,N_991);
nor U1788 (N_1788,N_1019,N_775);
and U1789 (N_1789,N_939,N_823);
and U1790 (N_1790,N_919,N_980);
nand U1791 (N_1791,N_818,N_771);
nand U1792 (N_1792,N_766,N_1062);
nor U1793 (N_1793,N_1040,N_1272);
or U1794 (N_1794,N_849,N_1098);
nor U1795 (N_1795,N_1396,N_1237);
nor U1796 (N_1796,N_878,N_1207);
nor U1797 (N_1797,N_1311,N_1345);
xor U1798 (N_1798,N_1193,N_988);
nor U1799 (N_1799,N_922,N_965);
nor U1800 (N_1800,N_1002,N_970);
nand U1801 (N_1801,N_903,N_1233);
nor U1802 (N_1802,N_1354,N_1196);
or U1803 (N_1803,N_1319,N_848);
and U1804 (N_1804,N_1008,N_877);
nor U1805 (N_1805,N_841,N_814);
nand U1806 (N_1806,N_1203,N_1424);
nand U1807 (N_1807,N_1156,N_885);
nor U1808 (N_1808,N_1140,N_761);
nor U1809 (N_1809,N_840,N_872);
nor U1810 (N_1810,N_1281,N_788);
and U1811 (N_1811,N_1338,N_777);
and U1812 (N_1812,N_926,N_1141);
nor U1813 (N_1813,N_1165,N_1212);
or U1814 (N_1814,N_1155,N_1280);
and U1815 (N_1815,N_1383,N_835);
and U1816 (N_1816,N_1069,N_1446);
or U1817 (N_1817,N_1419,N_1030);
and U1818 (N_1818,N_1000,N_1348);
and U1819 (N_1819,N_1036,N_876);
and U1820 (N_1820,N_757,N_776);
or U1821 (N_1821,N_932,N_948);
or U1822 (N_1822,N_869,N_1460);
xnor U1823 (N_1823,N_1395,N_1494);
and U1824 (N_1824,N_826,N_1270);
nand U1825 (N_1825,N_1381,N_1211);
or U1826 (N_1826,N_1072,N_1105);
nand U1827 (N_1827,N_1483,N_1361);
nand U1828 (N_1828,N_753,N_833);
xor U1829 (N_1829,N_874,N_917);
nand U1830 (N_1830,N_778,N_944);
or U1831 (N_1831,N_1255,N_1157);
xor U1832 (N_1832,N_1404,N_943);
nor U1833 (N_1833,N_1448,N_961);
nor U1834 (N_1834,N_1118,N_1126);
or U1835 (N_1835,N_881,N_1187);
xor U1836 (N_1836,N_1084,N_807);
and U1837 (N_1837,N_1382,N_1095);
nor U1838 (N_1838,N_995,N_822);
xor U1839 (N_1839,N_1394,N_884);
or U1840 (N_1840,N_969,N_1258);
xor U1841 (N_1841,N_1257,N_1418);
and U1842 (N_1842,N_1161,N_830);
and U1843 (N_1843,N_785,N_1391);
nand U1844 (N_1844,N_1089,N_804);
or U1845 (N_1845,N_1153,N_1402);
nor U1846 (N_1846,N_1016,N_1188);
and U1847 (N_1847,N_1371,N_1083);
or U1848 (N_1848,N_1388,N_929);
or U1849 (N_1849,N_1472,N_900);
and U1850 (N_1850,N_1252,N_1215);
or U1851 (N_1851,N_1474,N_774);
or U1852 (N_1852,N_1177,N_1350);
and U1853 (N_1853,N_1353,N_1092);
nand U1854 (N_1854,N_1099,N_981);
nand U1855 (N_1855,N_1186,N_825);
nor U1856 (N_1856,N_1026,N_1273);
and U1857 (N_1857,N_1018,N_1031);
nand U1858 (N_1858,N_787,N_1316);
and U1859 (N_1859,N_845,N_1296);
and U1860 (N_1860,N_1184,N_1314);
xnor U1861 (N_1861,N_1380,N_786);
nor U1862 (N_1862,N_1478,N_898);
nor U1863 (N_1863,N_1300,N_1061);
nand U1864 (N_1864,N_839,N_1011);
xnor U1865 (N_1865,N_1482,N_828);
and U1866 (N_1866,N_1307,N_846);
xnor U1867 (N_1867,N_1334,N_843);
nor U1868 (N_1868,N_895,N_795);
nand U1869 (N_1869,N_800,N_956);
nand U1870 (N_1870,N_1243,N_1039);
nand U1871 (N_1871,N_1183,N_1499);
nor U1872 (N_1872,N_928,N_1142);
nor U1873 (N_1873,N_1360,N_890);
and U1874 (N_1874,N_880,N_1181);
nand U1875 (N_1875,N_1337,N_790);
nor U1876 (N_1876,N_1128,N_1444);
nand U1877 (N_1877,N_845,N_1129);
nand U1878 (N_1878,N_824,N_765);
nand U1879 (N_1879,N_915,N_1489);
nor U1880 (N_1880,N_824,N_868);
nand U1881 (N_1881,N_998,N_1204);
and U1882 (N_1882,N_935,N_1249);
and U1883 (N_1883,N_922,N_1146);
or U1884 (N_1884,N_893,N_1092);
or U1885 (N_1885,N_959,N_1194);
or U1886 (N_1886,N_1452,N_1238);
and U1887 (N_1887,N_1235,N_1243);
or U1888 (N_1888,N_1467,N_822);
and U1889 (N_1889,N_1408,N_776);
xor U1890 (N_1890,N_1376,N_1048);
nor U1891 (N_1891,N_1280,N_861);
and U1892 (N_1892,N_759,N_875);
nand U1893 (N_1893,N_1413,N_1411);
xor U1894 (N_1894,N_825,N_1465);
and U1895 (N_1895,N_903,N_764);
nand U1896 (N_1896,N_1366,N_847);
nor U1897 (N_1897,N_1326,N_1386);
nor U1898 (N_1898,N_979,N_817);
nor U1899 (N_1899,N_1468,N_1167);
nor U1900 (N_1900,N_1443,N_1020);
nor U1901 (N_1901,N_1396,N_753);
nor U1902 (N_1902,N_1089,N_1115);
xor U1903 (N_1903,N_1217,N_1033);
or U1904 (N_1904,N_1449,N_1074);
nor U1905 (N_1905,N_1141,N_1447);
nand U1906 (N_1906,N_758,N_1128);
and U1907 (N_1907,N_1493,N_1237);
and U1908 (N_1908,N_1018,N_1332);
and U1909 (N_1909,N_995,N_1402);
and U1910 (N_1910,N_1366,N_1409);
and U1911 (N_1911,N_1109,N_1129);
nand U1912 (N_1912,N_882,N_972);
nor U1913 (N_1913,N_1398,N_1114);
and U1914 (N_1914,N_929,N_1209);
nor U1915 (N_1915,N_1270,N_896);
nand U1916 (N_1916,N_941,N_1031);
nand U1917 (N_1917,N_974,N_1152);
and U1918 (N_1918,N_1489,N_1337);
xnor U1919 (N_1919,N_1379,N_808);
nand U1920 (N_1920,N_1213,N_918);
nor U1921 (N_1921,N_1247,N_1092);
nor U1922 (N_1922,N_1181,N_1406);
or U1923 (N_1923,N_1103,N_1433);
nor U1924 (N_1924,N_915,N_1083);
xnor U1925 (N_1925,N_920,N_1259);
or U1926 (N_1926,N_1152,N_1415);
nor U1927 (N_1927,N_921,N_767);
and U1928 (N_1928,N_835,N_1047);
and U1929 (N_1929,N_925,N_1279);
xnor U1930 (N_1930,N_818,N_996);
nand U1931 (N_1931,N_1060,N_1446);
or U1932 (N_1932,N_1229,N_993);
xor U1933 (N_1933,N_884,N_1184);
and U1934 (N_1934,N_1270,N_1075);
nor U1935 (N_1935,N_1003,N_1186);
nand U1936 (N_1936,N_965,N_1223);
nor U1937 (N_1937,N_1193,N_891);
nor U1938 (N_1938,N_917,N_1427);
nand U1939 (N_1939,N_1376,N_953);
and U1940 (N_1940,N_1381,N_804);
nor U1941 (N_1941,N_1364,N_963);
and U1942 (N_1942,N_1486,N_954);
and U1943 (N_1943,N_1043,N_936);
nor U1944 (N_1944,N_855,N_954);
and U1945 (N_1945,N_769,N_1267);
nor U1946 (N_1946,N_1229,N_900);
nor U1947 (N_1947,N_1053,N_1253);
or U1948 (N_1948,N_950,N_1456);
nor U1949 (N_1949,N_1171,N_1113);
and U1950 (N_1950,N_1021,N_1459);
or U1951 (N_1951,N_1075,N_834);
nor U1952 (N_1952,N_825,N_767);
nand U1953 (N_1953,N_1373,N_1338);
nor U1954 (N_1954,N_1479,N_1045);
and U1955 (N_1955,N_880,N_1058);
nand U1956 (N_1956,N_935,N_1334);
and U1957 (N_1957,N_1132,N_1190);
nand U1958 (N_1958,N_1202,N_1138);
and U1959 (N_1959,N_877,N_841);
nor U1960 (N_1960,N_875,N_1241);
and U1961 (N_1961,N_1378,N_1237);
or U1962 (N_1962,N_1006,N_790);
nor U1963 (N_1963,N_889,N_1140);
nor U1964 (N_1964,N_1114,N_834);
or U1965 (N_1965,N_1253,N_1340);
or U1966 (N_1966,N_950,N_1179);
or U1967 (N_1967,N_1248,N_1243);
or U1968 (N_1968,N_973,N_763);
or U1969 (N_1969,N_1301,N_903);
and U1970 (N_1970,N_1325,N_1170);
and U1971 (N_1971,N_1136,N_1404);
nand U1972 (N_1972,N_1132,N_1312);
nor U1973 (N_1973,N_1079,N_1129);
nor U1974 (N_1974,N_1469,N_1096);
and U1975 (N_1975,N_1300,N_1271);
nor U1976 (N_1976,N_984,N_1470);
and U1977 (N_1977,N_1466,N_1355);
nor U1978 (N_1978,N_984,N_1147);
xnor U1979 (N_1979,N_1311,N_888);
nand U1980 (N_1980,N_1412,N_1342);
nand U1981 (N_1981,N_1184,N_756);
and U1982 (N_1982,N_1483,N_1294);
nand U1983 (N_1983,N_1280,N_920);
and U1984 (N_1984,N_754,N_766);
and U1985 (N_1985,N_861,N_975);
or U1986 (N_1986,N_1407,N_1161);
nand U1987 (N_1987,N_781,N_1457);
and U1988 (N_1988,N_1379,N_1047);
and U1989 (N_1989,N_1243,N_1339);
nor U1990 (N_1990,N_1447,N_1348);
and U1991 (N_1991,N_941,N_969);
and U1992 (N_1992,N_1024,N_1349);
or U1993 (N_1993,N_1335,N_1328);
nor U1994 (N_1994,N_1074,N_962);
nand U1995 (N_1995,N_792,N_1204);
and U1996 (N_1996,N_1476,N_1136);
or U1997 (N_1997,N_1305,N_792);
and U1998 (N_1998,N_1456,N_1351);
and U1999 (N_1999,N_971,N_1142);
nand U2000 (N_2000,N_1486,N_994);
nand U2001 (N_2001,N_1048,N_861);
nor U2002 (N_2002,N_1275,N_854);
and U2003 (N_2003,N_1189,N_1437);
or U2004 (N_2004,N_1063,N_1464);
and U2005 (N_2005,N_1191,N_1152);
xnor U2006 (N_2006,N_825,N_770);
nand U2007 (N_2007,N_1237,N_783);
nand U2008 (N_2008,N_1328,N_764);
nand U2009 (N_2009,N_1469,N_1205);
and U2010 (N_2010,N_1138,N_819);
nor U2011 (N_2011,N_766,N_1171);
nor U2012 (N_2012,N_1169,N_1005);
or U2013 (N_2013,N_1138,N_1397);
nand U2014 (N_2014,N_1358,N_1267);
and U2015 (N_2015,N_975,N_1394);
or U2016 (N_2016,N_1226,N_1392);
and U2017 (N_2017,N_878,N_839);
and U2018 (N_2018,N_1300,N_1337);
nand U2019 (N_2019,N_1423,N_1040);
nor U2020 (N_2020,N_1110,N_1432);
or U2021 (N_2021,N_840,N_1455);
nor U2022 (N_2022,N_903,N_1076);
nand U2023 (N_2023,N_846,N_1249);
nor U2024 (N_2024,N_1231,N_1014);
nand U2025 (N_2025,N_1495,N_1441);
nor U2026 (N_2026,N_1400,N_851);
or U2027 (N_2027,N_1491,N_1395);
or U2028 (N_2028,N_774,N_1118);
nand U2029 (N_2029,N_1390,N_886);
or U2030 (N_2030,N_1023,N_1274);
or U2031 (N_2031,N_1317,N_1267);
nand U2032 (N_2032,N_1263,N_1189);
or U2033 (N_2033,N_1224,N_1077);
or U2034 (N_2034,N_1084,N_1251);
nor U2035 (N_2035,N_1064,N_1316);
or U2036 (N_2036,N_1114,N_941);
and U2037 (N_2037,N_1361,N_1093);
nand U2038 (N_2038,N_1224,N_1300);
nand U2039 (N_2039,N_865,N_1087);
and U2040 (N_2040,N_1455,N_1365);
nand U2041 (N_2041,N_790,N_1095);
nand U2042 (N_2042,N_991,N_1117);
xor U2043 (N_2043,N_928,N_1322);
or U2044 (N_2044,N_1153,N_1484);
nand U2045 (N_2045,N_1209,N_1279);
nor U2046 (N_2046,N_1484,N_1166);
nand U2047 (N_2047,N_1189,N_1422);
nand U2048 (N_2048,N_1236,N_889);
xor U2049 (N_2049,N_1302,N_1056);
nor U2050 (N_2050,N_1348,N_796);
nand U2051 (N_2051,N_997,N_1229);
xor U2052 (N_2052,N_1301,N_1236);
xor U2053 (N_2053,N_1277,N_1367);
and U2054 (N_2054,N_992,N_820);
nor U2055 (N_2055,N_777,N_1107);
or U2056 (N_2056,N_1284,N_1494);
nor U2057 (N_2057,N_1432,N_858);
and U2058 (N_2058,N_996,N_1188);
nand U2059 (N_2059,N_1123,N_908);
nand U2060 (N_2060,N_1364,N_827);
nor U2061 (N_2061,N_1421,N_1463);
nand U2062 (N_2062,N_835,N_1136);
or U2063 (N_2063,N_1403,N_1390);
and U2064 (N_2064,N_1034,N_1439);
or U2065 (N_2065,N_898,N_784);
nor U2066 (N_2066,N_1370,N_1199);
or U2067 (N_2067,N_1130,N_1100);
or U2068 (N_2068,N_885,N_798);
nor U2069 (N_2069,N_1121,N_1074);
nor U2070 (N_2070,N_785,N_1440);
nor U2071 (N_2071,N_865,N_1115);
nand U2072 (N_2072,N_770,N_1187);
or U2073 (N_2073,N_1160,N_902);
nand U2074 (N_2074,N_1394,N_1181);
xnor U2075 (N_2075,N_1452,N_979);
and U2076 (N_2076,N_811,N_1082);
or U2077 (N_2077,N_1329,N_914);
and U2078 (N_2078,N_1106,N_1251);
or U2079 (N_2079,N_1306,N_1289);
and U2080 (N_2080,N_1485,N_1103);
and U2081 (N_2081,N_1036,N_1194);
xnor U2082 (N_2082,N_887,N_1245);
and U2083 (N_2083,N_932,N_1414);
and U2084 (N_2084,N_986,N_1422);
or U2085 (N_2085,N_1150,N_1434);
nor U2086 (N_2086,N_945,N_764);
nand U2087 (N_2087,N_1067,N_1287);
and U2088 (N_2088,N_1434,N_1390);
or U2089 (N_2089,N_1093,N_767);
nor U2090 (N_2090,N_1432,N_977);
xnor U2091 (N_2091,N_1079,N_1429);
xor U2092 (N_2092,N_927,N_801);
xor U2093 (N_2093,N_1046,N_1333);
nand U2094 (N_2094,N_1375,N_1196);
or U2095 (N_2095,N_1458,N_788);
nand U2096 (N_2096,N_1056,N_775);
nand U2097 (N_2097,N_1000,N_1261);
or U2098 (N_2098,N_797,N_753);
nand U2099 (N_2099,N_786,N_835);
nand U2100 (N_2100,N_1082,N_1384);
or U2101 (N_2101,N_1319,N_892);
or U2102 (N_2102,N_1012,N_992);
nor U2103 (N_2103,N_936,N_1447);
or U2104 (N_2104,N_1112,N_1487);
nand U2105 (N_2105,N_1462,N_756);
xnor U2106 (N_2106,N_1208,N_1162);
nor U2107 (N_2107,N_1042,N_1361);
or U2108 (N_2108,N_1026,N_870);
or U2109 (N_2109,N_829,N_1070);
nor U2110 (N_2110,N_1053,N_1427);
nor U2111 (N_2111,N_880,N_902);
nand U2112 (N_2112,N_882,N_945);
or U2113 (N_2113,N_1052,N_1169);
nand U2114 (N_2114,N_1402,N_1013);
nor U2115 (N_2115,N_975,N_1285);
nand U2116 (N_2116,N_794,N_1338);
nor U2117 (N_2117,N_1477,N_1295);
nand U2118 (N_2118,N_960,N_920);
nand U2119 (N_2119,N_1447,N_807);
nand U2120 (N_2120,N_996,N_1267);
nor U2121 (N_2121,N_942,N_916);
nor U2122 (N_2122,N_950,N_1289);
or U2123 (N_2123,N_807,N_786);
nand U2124 (N_2124,N_959,N_1067);
nand U2125 (N_2125,N_1372,N_1316);
xnor U2126 (N_2126,N_809,N_1295);
and U2127 (N_2127,N_1140,N_1155);
nand U2128 (N_2128,N_812,N_1309);
nand U2129 (N_2129,N_1253,N_1276);
and U2130 (N_2130,N_1211,N_807);
xor U2131 (N_2131,N_866,N_984);
nand U2132 (N_2132,N_1082,N_1026);
and U2133 (N_2133,N_1081,N_1219);
or U2134 (N_2134,N_901,N_1247);
nand U2135 (N_2135,N_1284,N_1262);
nand U2136 (N_2136,N_916,N_859);
and U2137 (N_2137,N_895,N_956);
xor U2138 (N_2138,N_1033,N_835);
or U2139 (N_2139,N_983,N_1220);
and U2140 (N_2140,N_1354,N_1409);
xor U2141 (N_2141,N_972,N_1181);
and U2142 (N_2142,N_1040,N_1331);
nand U2143 (N_2143,N_1050,N_958);
nand U2144 (N_2144,N_1474,N_815);
nand U2145 (N_2145,N_1094,N_1049);
and U2146 (N_2146,N_951,N_906);
or U2147 (N_2147,N_859,N_1321);
nand U2148 (N_2148,N_793,N_1242);
nand U2149 (N_2149,N_900,N_783);
or U2150 (N_2150,N_1184,N_1334);
nand U2151 (N_2151,N_1001,N_818);
nor U2152 (N_2152,N_999,N_1477);
or U2153 (N_2153,N_965,N_905);
nor U2154 (N_2154,N_1171,N_1155);
and U2155 (N_2155,N_1433,N_1184);
xor U2156 (N_2156,N_1067,N_1249);
nand U2157 (N_2157,N_1177,N_1130);
nand U2158 (N_2158,N_902,N_1108);
and U2159 (N_2159,N_953,N_1417);
and U2160 (N_2160,N_878,N_1308);
or U2161 (N_2161,N_1259,N_1473);
nor U2162 (N_2162,N_907,N_1102);
nand U2163 (N_2163,N_1027,N_832);
and U2164 (N_2164,N_1152,N_1198);
or U2165 (N_2165,N_1252,N_1209);
and U2166 (N_2166,N_1341,N_1173);
nand U2167 (N_2167,N_1016,N_998);
nand U2168 (N_2168,N_915,N_1021);
nor U2169 (N_2169,N_1158,N_754);
nand U2170 (N_2170,N_1406,N_929);
xor U2171 (N_2171,N_898,N_806);
nand U2172 (N_2172,N_1087,N_1445);
nand U2173 (N_2173,N_959,N_1243);
or U2174 (N_2174,N_959,N_1451);
xnor U2175 (N_2175,N_1321,N_1257);
nor U2176 (N_2176,N_1300,N_868);
and U2177 (N_2177,N_766,N_1309);
nor U2178 (N_2178,N_1201,N_1383);
and U2179 (N_2179,N_886,N_1126);
nor U2180 (N_2180,N_1095,N_1094);
nand U2181 (N_2181,N_1399,N_905);
xnor U2182 (N_2182,N_1263,N_1050);
and U2183 (N_2183,N_1297,N_845);
nor U2184 (N_2184,N_898,N_1325);
or U2185 (N_2185,N_913,N_941);
nand U2186 (N_2186,N_1214,N_1302);
nand U2187 (N_2187,N_995,N_775);
nand U2188 (N_2188,N_817,N_1420);
nand U2189 (N_2189,N_1058,N_1374);
or U2190 (N_2190,N_1457,N_869);
nand U2191 (N_2191,N_1143,N_775);
nand U2192 (N_2192,N_1297,N_1216);
or U2193 (N_2193,N_990,N_1161);
and U2194 (N_2194,N_1429,N_1414);
nor U2195 (N_2195,N_1180,N_1077);
xor U2196 (N_2196,N_901,N_1463);
or U2197 (N_2197,N_835,N_1097);
xor U2198 (N_2198,N_1428,N_1073);
or U2199 (N_2199,N_1381,N_1437);
and U2200 (N_2200,N_1203,N_1477);
and U2201 (N_2201,N_1113,N_1269);
nor U2202 (N_2202,N_1229,N_1088);
nor U2203 (N_2203,N_894,N_1441);
and U2204 (N_2204,N_1250,N_929);
nand U2205 (N_2205,N_1492,N_1138);
or U2206 (N_2206,N_1427,N_1243);
or U2207 (N_2207,N_956,N_902);
xor U2208 (N_2208,N_1358,N_877);
xor U2209 (N_2209,N_1245,N_1269);
xor U2210 (N_2210,N_792,N_1447);
nor U2211 (N_2211,N_1097,N_1030);
or U2212 (N_2212,N_1063,N_1225);
nand U2213 (N_2213,N_1232,N_990);
or U2214 (N_2214,N_890,N_1411);
nor U2215 (N_2215,N_1373,N_1366);
xor U2216 (N_2216,N_894,N_1200);
and U2217 (N_2217,N_1464,N_1438);
nor U2218 (N_2218,N_1325,N_1099);
and U2219 (N_2219,N_1197,N_1496);
xor U2220 (N_2220,N_1417,N_958);
and U2221 (N_2221,N_1395,N_923);
and U2222 (N_2222,N_854,N_801);
nor U2223 (N_2223,N_802,N_1220);
nor U2224 (N_2224,N_1186,N_1384);
xor U2225 (N_2225,N_1308,N_1301);
or U2226 (N_2226,N_873,N_1231);
nand U2227 (N_2227,N_1465,N_947);
nand U2228 (N_2228,N_959,N_1486);
nor U2229 (N_2229,N_1007,N_1225);
nand U2230 (N_2230,N_1336,N_844);
or U2231 (N_2231,N_1056,N_1438);
xor U2232 (N_2232,N_901,N_902);
nand U2233 (N_2233,N_1429,N_1241);
xor U2234 (N_2234,N_974,N_852);
nand U2235 (N_2235,N_1088,N_1405);
and U2236 (N_2236,N_826,N_1081);
or U2237 (N_2237,N_1317,N_1266);
nand U2238 (N_2238,N_977,N_796);
or U2239 (N_2239,N_1238,N_838);
nand U2240 (N_2240,N_883,N_1254);
or U2241 (N_2241,N_1499,N_1179);
or U2242 (N_2242,N_1264,N_862);
nor U2243 (N_2243,N_1071,N_1293);
nor U2244 (N_2244,N_940,N_1485);
and U2245 (N_2245,N_988,N_1221);
xor U2246 (N_2246,N_884,N_919);
nor U2247 (N_2247,N_1340,N_806);
and U2248 (N_2248,N_871,N_1274);
nand U2249 (N_2249,N_1388,N_1129);
or U2250 (N_2250,N_1509,N_1597);
nand U2251 (N_2251,N_1561,N_2193);
or U2252 (N_2252,N_2005,N_1841);
xor U2253 (N_2253,N_2006,N_1556);
nor U2254 (N_2254,N_2054,N_1697);
nor U2255 (N_2255,N_2019,N_1536);
nand U2256 (N_2256,N_1600,N_1892);
nor U2257 (N_2257,N_2033,N_1682);
nor U2258 (N_2258,N_2173,N_1636);
and U2259 (N_2259,N_1696,N_1854);
and U2260 (N_2260,N_1555,N_1825);
or U2261 (N_2261,N_2246,N_2237);
or U2262 (N_2262,N_1716,N_1727);
or U2263 (N_2263,N_2013,N_1686);
or U2264 (N_2264,N_2231,N_2039);
and U2265 (N_2265,N_1544,N_1874);
nor U2266 (N_2266,N_2205,N_2027);
nor U2267 (N_2267,N_1670,N_2144);
nand U2268 (N_2268,N_1647,N_2131);
nand U2269 (N_2269,N_2097,N_2084);
nand U2270 (N_2270,N_1777,N_1606);
nor U2271 (N_2271,N_1560,N_2004);
nor U2272 (N_2272,N_1602,N_1804);
and U2273 (N_2273,N_1963,N_2244);
and U2274 (N_2274,N_1713,N_2143);
or U2275 (N_2275,N_1968,N_1537);
nor U2276 (N_2276,N_2122,N_1843);
nand U2277 (N_2277,N_2216,N_1876);
nor U2278 (N_2278,N_1778,N_1562);
nand U2279 (N_2279,N_2111,N_2167);
or U2280 (N_2280,N_2243,N_1699);
nor U2281 (N_2281,N_2140,N_1956);
nor U2282 (N_2282,N_1770,N_1848);
or U2283 (N_2283,N_1621,N_2209);
xor U2284 (N_2284,N_2032,N_2046);
or U2285 (N_2285,N_2170,N_1741);
nand U2286 (N_2286,N_2057,N_1888);
or U2287 (N_2287,N_1932,N_2211);
or U2288 (N_2288,N_1835,N_1588);
nand U2289 (N_2289,N_2227,N_1813);
and U2290 (N_2290,N_1583,N_2195);
or U2291 (N_2291,N_1726,N_1883);
nor U2292 (N_2292,N_1873,N_1833);
nand U2293 (N_2293,N_1782,N_2048);
xnor U2294 (N_2294,N_1720,N_2015);
nor U2295 (N_2295,N_1812,N_1750);
nor U2296 (N_2296,N_1521,N_1623);
or U2297 (N_2297,N_1648,N_1516);
nor U2298 (N_2298,N_1771,N_1965);
or U2299 (N_2299,N_2150,N_1901);
nand U2300 (N_2300,N_2207,N_1858);
nand U2301 (N_2301,N_1882,N_1659);
or U2302 (N_2302,N_2029,N_1590);
or U2303 (N_2303,N_2105,N_1959);
or U2304 (N_2304,N_1625,N_1717);
or U2305 (N_2305,N_2003,N_1802);
nor U2306 (N_2306,N_1893,N_1995);
or U2307 (N_2307,N_2183,N_1649);
xnor U2308 (N_2308,N_1994,N_1834);
or U2309 (N_2309,N_1880,N_1706);
nor U2310 (N_2310,N_2241,N_1530);
or U2311 (N_2311,N_1891,N_1755);
nor U2312 (N_2312,N_1567,N_1928);
and U2313 (N_2313,N_2191,N_1573);
and U2314 (N_2314,N_1635,N_1950);
and U2315 (N_2315,N_1576,N_1526);
and U2316 (N_2316,N_1681,N_1952);
nor U2317 (N_2317,N_1768,N_1695);
or U2318 (N_2318,N_2229,N_1594);
or U2319 (N_2319,N_2206,N_1667);
and U2320 (N_2320,N_1679,N_1759);
or U2321 (N_2321,N_1933,N_2001);
nor U2322 (N_2322,N_1515,N_1924);
or U2323 (N_2323,N_2014,N_1601);
or U2324 (N_2324,N_2182,N_1735);
xnor U2325 (N_2325,N_2224,N_2116);
nand U2326 (N_2326,N_2129,N_1700);
or U2327 (N_2327,N_2093,N_1661);
or U2328 (N_2328,N_1578,N_1748);
or U2329 (N_2329,N_1957,N_1614);
nand U2330 (N_2330,N_1714,N_1853);
and U2331 (N_2331,N_2215,N_1624);
or U2332 (N_2332,N_1511,N_1524);
xor U2333 (N_2333,N_1532,N_1973);
and U2334 (N_2334,N_1751,N_1514);
xnor U2335 (N_2335,N_2175,N_2024);
and U2336 (N_2336,N_1620,N_1784);
and U2337 (N_2337,N_2007,N_1707);
xor U2338 (N_2338,N_1722,N_1809);
nand U2339 (N_2339,N_1508,N_2091);
nor U2340 (N_2340,N_2010,N_2164);
nand U2341 (N_2341,N_1541,N_1799);
and U2342 (N_2342,N_2184,N_1864);
nand U2343 (N_2343,N_1830,N_1810);
xor U2344 (N_2344,N_1910,N_1746);
xnor U2345 (N_2345,N_1862,N_1985);
nor U2346 (N_2346,N_1840,N_2133);
nand U2347 (N_2347,N_1917,N_1897);
or U2348 (N_2348,N_1775,N_1628);
xnor U2349 (N_2349,N_1905,N_1806);
nor U2350 (N_2350,N_1797,N_2149);
nor U2351 (N_2351,N_1736,N_1603);
nor U2352 (N_2352,N_1629,N_2221);
or U2353 (N_2353,N_1923,N_2192);
nor U2354 (N_2354,N_2198,N_1640);
nor U2355 (N_2355,N_2147,N_1946);
nor U2356 (N_2356,N_2132,N_1823);
or U2357 (N_2357,N_2135,N_1839);
or U2358 (N_2358,N_1633,N_1749);
nand U2359 (N_2359,N_1643,N_2063);
xnor U2360 (N_2360,N_1572,N_2159);
or U2361 (N_2361,N_1738,N_2138);
or U2362 (N_2362,N_1915,N_2061);
and U2363 (N_2363,N_2125,N_1800);
xnor U2364 (N_2364,N_1570,N_1691);
nand U2365 (N_2365,N_1523,N_1550);
nor U2366 (N_2366,N_1980,N_2021);
nand U2367 (N_2367,N_2194,N_2062);
or U2368 (N_2368,N_2071,N_1737);
nand U2369 (N_2369,N_1710,N_1857);
and U2370 (N_2370,N_2233,N_2226);
or U2371 (N_2371,N_1983,N_1894);
and U2372 (N_2372,N_1676,N_2079);
and U2373 (N_2373,N_2176,N_1916);
nor U2374 (N_2374,N_2179,N_1861);
nand U2375 (N_2375,N_1796,N_1967);
xnor U2376 (N_2376,N_1575,N_2165);
and U2377 (N_2377,N_2174,N_1920);
or U2378 (N_2378,N_2186,N_2108);
or U2379 (N_2379,N_1757,N_1531);
and U2380 (N_2380,N_1780,N_2092);
nand U2381 (N_2381,N_1731,N_1569);
xnor U2382 (N_2382,N_1961,N_1831);
nor U2383 (N_2383,N_1551,N_1564);
and U2384 (N_2384,N_2080,N_1964);
or U2385 (N_2385,N_1520,N_2100);
nor U2386 (N_2386,N_1895,N_1673);
nor U2387 (N_2387,N_1984,N_1711);
nand U2388 (N_2388,N_1728,N_1535);
nor U2389 (N_2389,N_2230,N_1921);
nand U2390 (N_2390,N_2248,N_1558);
or U2391 (N_2391,N_1553,N_1791);
nand U2392 (N_2392,N_1918,N_2234);
nor U2393 (N_2393,N_2118,N_2223);
and U2394 (N_2394,N_1886,N_1906);
xor U2395 (N_2395,N_2225,N_1653);
or U2396 (N_2396,N_1846,N_2085);
and U2397 (N_2397,N_1552,N_1721);
or U2398 (N_2398,N_1817,N_2086);
nand U2399 (N_2399,N_1724,N_1715);
or U2400 (N_2400,N_1815,N_1926);
or U2401 (N_2401,N_1518,N_1881);
or U2402 (N_2402,N_1505,N_1546);
nor U2403 (N_2403,N_2200,N_2065);
and U2404 (N_2404,N_2107,N_1589);
or U2405 (N_2405,N_1938,N_1912);
and U2406 (N_2406,N_2247,N_1645);
nor U2407 (N_2407,N_2128,N_1855);
and U2408 (N_2408,N_1534,N_1794);
nor U2409 (N_2409,N_1739,N_2012);
nand U2410 (N_2410,N_1798,N_2037);
and U2411 (N_2411,N_1903,N_1887);
and U2412 (N_2412,N_1890,N_1745);
or U2413 (N_2413,N_2096,N_1754);
nand U2414 (N_2414,N_1540,N_1847);
xnor U2415 (N_2415,N_2017,N_1948);
nand U2416 (N_2416,N_1610,N_1944);
nand U2417 (N_2417,N_1677,N_1851);
or U2418 (N_2418,N_1599,N_1548);
and U2419 (N_2419,N_1925,N_1683);
or U2420 (N_2420,N_1631,N_2090);
or U2421 (N_2421,N_1877,N_1818);
nand U2422 (N_2422,N_1816,N_1609);
nor U2423 (N_2423,N_1704,N_2011);
nor U2424 (N_2424,N_1795,N_1662);
nand U2425 (N_2425,N_1842,N_1725);
and U2426 (N_2426,N_2047,N_1752);
and U2427 (N_2427,N_2002,N_2172);
nor U2428 (N_2428,N_1978,N_2056);
and U2429 (N_2429,N_1668,N_1652);
and U2430 (N_2430,N_1593,N_1740);
nor U2431 (N_2431,N_1630,N_1547);
xor U2432 (N_2432,N_2127,N_2137);
xor U2433 (N_2433,N_1519,N_2213);
nand U2434 (N_2434,N_1580,N_1940);
and U2435 (N_2435,N_2232,N_1618);
nor U2436 (N_2436,N_1859,N_2134);
and U2437 (N_2437,N_2074,N_1774);
nor U2438 (N_2438,N_1539,N_1969);
nand U2439 (N_2439,N_1522,N_1612);
or U2440 (N_2440,N_1875,N_1646);
and U2441 (N_2441,N_1786,N_1783);
nand U2442 (N_2442,N_1733,N_1581);
or U2443 (N_2443,N_1878,N_1598);
and U2444 (N_2444,N_1658,N_1885);
nor U2445 (N_2445,N_1904,N_1650);
nor U2446 (N_2446,N_1970,N_2113);
nor U2447 (N_2447,N_1793,N_2154);
and U2448 (N_2448,N_1512,N_1849);
xnor U2449 (N_2449,N_1604,N_1587);
and U2450 (N_2450,N_2210,N_1690);
or U2451 (N_2451,N_2228,N_1909);
xnor U2452 (N_2452,N_1586,N_2066);
nor U2453 (N_2453,N_2058,N_1987);
nand U2454 (N_2454,N_2160,N_2123);
nor U2455 (N_2455,N_2030,N_2064);
nand U2456 (N_2456,N_2031,N_1898);
nand U2457 (N_2457,N_1563,N_1951);
nand U2458 (N_2458,N_1712,N_1922);
and U2459 (N_2459,N_2162,N_1568);
or U2460 (N_2460,N_2052,N_1701);
and U2461 (N_2461,N_2217,N_1977);
nor U2462 (N_2462,N_1822,N_1545);
nor U2463 (N_2463,N_1732,N_1958);
nand U2464 (N_2464,N_2189,N_1960);
or U2465 (N_2465,N_2009,N_1582);
and U2466 (N_2466,N_1884,N_2095);
xor U2467 (N_2467,N_2023,N_1503);
nand U2468 (N_2468,N_1989,N_1900);
and U2469 (N_2469,N_1819,N_1975);
and U2470 (N_2470,N_1845,N_1743);
xnor U2471 (N_2471,N_1642,N_1947);
nand U2472 (N_2472,N_2078,N_1927);
nand U2473 (N_2473,N_2060,N_1979);
xnor U2474 (N_2474,N_1651,N_2117);
xnor U2475 (N_2475,N_1929,N_1765);
nor U2476 (N_2476,N_1756,N_2124);
nand U2477 (N_2477,N_1773,N_2073);
xor U2478 (N_2478,N_1914,N_2051);
and U2479 (N_2479,N_1982,N_1501);
or U2480 (N_2480,N_2059,N_1675);
nor U2481 (N_2481,N_1634,N_1709);
or U2482 (N_2482,N_2098,N_1592);
nor U2483 (N_2483,N_1513,N_1502);
and U2484 (N_2484,N_2103,N_1571);
xor U2485 (N_2485,N_1870,N_2161);
nand U2486 (N_2486,N_2219,N_1767);
nor U2487 (N_2487,N_1872,N_1674);
or U2488 (N_2488,N_1981,N_1814);
or U2489 (N_2489,N_1931,N_2049);
nand U2490 (N_2490,N_1654,N_2136);
nand U2491 (N_2491,N_2145,N_1821);
and U2492 (N_2492,N_2045,N_1787);
and U2493 (N_2493,N_1678,N_1708);
nand U2494 (N_2494,N_2163,N_1533);
nand U2495 (N_2495,N_1828,N_2034);
and U2496 (N_2496,N_1999,N_1663);
and U2497 (N_2497,N_1865,N_1992);
nor U2498 (N_2498,N_1954,N_2028);
and U2499 (N_2499,N_2110,N_1638);
and U2500 (N_2500,N_1693,N_1500);
nand U2501 (N_2501,N_2155,N_2130);
nand U2502 (N_2502,N_2242,N_2181);
or U2503 (N_2503,N_1998,N_1769);
nand U2504 (N_2504,N_2177,N_1908);
and U2505 (N_2505,N_1829,N_1669);
and U2506 (N_2506,N_2044,N_1781);
and U2507 (N_2507,N_1761,N_1507);
or U2508 (N_2508,N_2099,N_1703);
nor U2509 (N_2509,N_1808,N_1805);
or U2510 (N_2510,N_1694,N_1807);
or U2511 (N_2511,N_1692,N_1758);
and U2512 (N_2512,N_1939,N_2249);
nand U2513 (N_2513,N_1632,N_1837);
nor U2514 (N_2514,N_1510,N_1949);
nor U2515 (N_2515,N_1579,N_1962);
or U2516 (N_2516,N_1907,N_1988);
xor U2517 (N_2517,N_1689,N_1971);
nand U2518 (N_2518,N_1655,N_2083);
or U2519 (N_2519,N_2082,N_2196);
and U2520 (N_2520,N_1820,N_1911);
or U2521 (N_2521,N_2094,N_1584);
xor U2522 (N_2522,N_2141,N_1826);
nor U2523 (N_2523,N_1574,N_2114);
nand U2524 (N_2524,N_1542,N_1672);
or U2525 (N_2525,N_1665,N_1976);
and U2526 (N_2526,N_1698,N_1607);
or U2527 (N_2527,N_2120,N_1811);
nand U2528 (N_2528,N_2235,N_1827);
nand U2529 (N_2529,N_1986,N_2158);
or U2530 (N_2530,N_2101,N_2070);
nor U2531 (N_2531,N_2199,N_1559);
and U2532 (N_2532,N_1566,N_1702);
or U2533 (N_2533,N_1506,N_1760);
and U2534 (N_2534,N_1896,N_2166);
nor U2535 (N_2535,N_1991,N_2240);
and U2536 (N_2536,N_1644,N_2043);
and U2537 (N_2537,N_1863,N_2236);
and U2538 (N_2538,N_1687,N_1776);
nand U2539 (N_2539,N_1930,N_2000);
nor U2540 (N_2540,N_1788,N_1657);
xor U2541 (N_2541,N_2201,N_2239);
xnor U2542 (N_2542,N_1844,N_2026);
and U2543 (N_2543,N_1742,N_2168);
xnor U2544 (N_2544,N_2053,N_2121);
nand U2545 (N_2545,N_1527,N_2050);
xor U2546 (N_2546,N_1943,N_2157);
or U2547 (N_2547,N_2180,N_1608);
nand U2548 (N_2548,N_1622,N_2112);
nand U2549 (N_2549,N_1639,N_2055);
xor U2550 (N_2550,N_1718,N_1688);
nor U2551 (N_2551,N_2202,N_1744);
or U2552 (N_2552,N_2020,N_2212);
nor U2553 (N_2553,N_2178,N_1705);
and U2554 (N_2554,N_2220,N_2075);
nor U2555 (N_2555,N_1615,N_1902);
nand U2556 (N_2556,N_2142,N_1504);
nand U2557 (N_2557,N_1641,N_1966);
xnor U2558 (N_2558,N_2077,N_1763);
or U2559 (N_2559,N_1734,N_1684);
and U2560 (N_2560,N_1942,N_1529);
nor U2561 (N_2561,N_2156,N_1517);
nand U2562 (N_2562,N_1866,N_2018);
or U2563 (N_2563,N_2067,N_1790);
or U2564 (N_2564,N_1990,N_1792);
nand U2565 (N_2565,N_2126,N_2008);
nand U2566 (N_2566,N_2088,N_2115);
and U2567 (N_2567,N_2089,N_2188);
xnor U2568 (N_2568,N_1730,N_2204);
nor U2569 (N_2569,N_2102,N_2016);
nand U2570 (N_2570,N_1656,N_1785);
or U2571 (N_2571,N_1596,N_1953);
nand U2572 (N_2572,N_1549,N_1753);
nand U2573 (N_2573,N_1850,N_2081);
nand U2574 (N_2574,N_1936,N_1637);
xor U2575 (N_2575,N_2146,N_1605);
and U2576 (N_2576,N_1838,N_1762);
nand U2577 (N_2577,N_2035,N_1803);
xor U2578 (N_2578,N_1772,N_2152);
and U2579 (N_2579,N_2025,N_1801);
nand U2580 (N_2580,N_2069,N_1627);
and U2581 (N_2581,N_1889,N_2076);
or U2582 (N_2582,N_2041,N_1913);
nor U2583 (N_2583,N_1955,N_2245);
nor U2584 (N_2584,N_1935,N_1836);
or U2585 (N_2585,N_1729,N_1613);
nor U2586 (N_2586,N_2185,N_2038);
and U2587 (N_2587,N_1554,N_1993);
nand U2588 (N_2588,N_2169,N_1577);
xor U2589 (N_2589,N_1779,N_1671);
or U2590 (N_2590,N_1871,N_2208);
and U2591 (N_2591,N_1766,N_1868);
or U2592 (N_2592,N_1660,N_2106);
nor U2593 (N_2593,N_2171,N_2109);
nand U2594 (N_2594,N_2203,N_2104);
nand U2595 (N_2595,N_1997,N_2139);
nor U2596 (N_2596,N_1972,N_1941);
or U2597 (N_2597,N_2040,N_1565);
and U2598 (N_2598,N_2072,N_2036);
or U2599 (N_2599,N_1832,N_1723);
nand U2600 (N_2600,N_2190,N_1945);
or U2601 (N_2601,N_2238,N_1626);
nand U2602 (N_2602,N_2151,N_1824);
nor U2603 (N_2603,N_2153,N_1617);
nor U2604 (N_2604,N_1680,N_1719);
and U2605 (N_2605,N_1869,N_1856);
or U2606 (N_2606,N_1611,N_1860);
xor U2607 (N_2607,N_2214,N_1974);
nand U2608 (N_2608,N_1619,N_1879);
nor U2609 (N_2609,N_2218,N_2042);
nor U2610 (N_2610,N_2087,N_1538);
nand U2611 (N_2611,N_2197,N_2022);
nor U2612 (N_2612,N_1528,N_1996);
nand U2613 (N_2613,N_2119,N_1591);
and U2614 (N_2614,N_1525,N_1747);
nor U2615 (N_2615,N_1867,N_1685);
nor U2616 (N_2616,N_1585,N_1919);
and U2617 (N_2617,N_1666,N_2222);
or U2618 (N_2618,N_1934,N_1616);
nand U2619 (N_2619,N_2148,N_1664);
nor U2620 (N_2620,N_1789,N_2068);
or U2621 (N_2621,N_1899,N_1764);
nor U2622 (N_2622,N_1557,N_1543);
xor U2623 (N_2623,N_1852,N_1937);
xnor U2624 (N_2624,N_2187,N_1595);
nor U2625 (N_2625,N_1623,N_1790);
nor U2626 (N_2626,N_2030,N_1733);
nand U2627 (N_2627,N_1777,N_2015);
or U2628 (N_2628,N_1788,N_1517);
and U2629 (N_2629,N_2195,N_2213);
nor U2630 (N_2630,N_1568,N_1867);
nor U2631 (N_2631,N_1950,N_1801);
nand U2632 (N_2632,N_2234,N_1972);
nand U2633 (N_2633,N_1631,N_1519);
and U2634 (N_2634,N_1761,N_1595);
and U2635 (N_2635,N_1829,N_1507);
xor U2636 (N_2636,N_2016,N_2180);
or U2637 (N_2637,N_2053,N_2143);
and U2638 (N_2638,N_1634,N_1532);
nor U2639 (N_2639,N_1990,N_2007);
nor U2640 (N_2640,N_2199,N_2059);
nor U2641 (N_2641,N_2129,N_1870);
nor U2642 (N_2642,N_1962,N_1530);
or U2643 (N_2643,N_2196,N_2028);
and U2644 (N_2644,N_1981,N_1572);
nand U2645 (N_2645,N_1564,N_2151);
nand U2646 (N_2646,N_1564,N_1876);
and U2647 (N_2647,N_2029,N_1943);
nor U2648 (N_2648,N_2104,N_1748);
or U2649 (N_2649,N_1642,N_1504);
xnor U2650 (N_2650,N_1666,N_1699);
nand U2651 (N_2651,N_1928,N_1852);
and U2652 (N_2652,N_1668,N_1902);
xnor U2653 (N_2653,N_1614,N_2249);
nand U2654 (N_2654,N_1555,N_2014);
and U2655 (N_2655,N_1907,N_2016);
or U2656 (N_2656,N_2132,N_1652);
or U2657 (N_2657,N_2205,N_1765);
or U2658 (N_2658,N_2027,N_1962);
and U2659 (N_2659,N_2209,N_1568);
nand U2660 (N_2660,N_1918,N_1805);
and U2661 (N_2661,N_1673,N_1509);
nand U2662 (N_2662,N_1740,N_1909);
xnor U2663 (N_2663,N_1993,N_2004);
xor U2664 (N_2664,N_2130,N_2038);
or U2665 (N_2665,N_2248,N_1617);
nor U2666 (N_2666,N_1800,N_1619);
nor U2667 (N_2667,N_2089,N_1509);
nor U2668 (N_2668,N_1532,N_1869);
or U2669 (N_2669,N_1748,N_2065);
nor U2670 (N_2670,N_2125,N_2074);
or U2671 (N_2671,N_2004,N_1765);
nor U2672 (N_2672,N_1889,N_1715);
or U2673 (N_2673,N_1682,N_2165);
nand U2674 (N_2674,N_2179,N_1561);
xnor U2675 (N_2675,N_1623,N_2021);
nor U2676 (N_2676,N_2069,N_1935);
xor U2677 (N_2677,N_1629,N_2020);
nand U2678 (N_2678,N_1714,N_1737);
nor U2679 (N_2679,N_1738,N_1684);
or U2680 (N_2680,N_2068,N_2103);
nor U2681 (N_2681,N_1590,N_2035);
or U2682 (N_2682,N_2199,N_1861);
or U2683 (N_2683,N_1802,N_1991);
and U2684 (N_2684,N_2075,N_1729);
nand U2685 (N_2685,N_1919,N_1742);
xnor U2686 (N_2686,N_1669,N_2213);
xor U2687 (N_2687,N_2215,N_2062);
or U2688 (N_2688,N_2006,N_2158);
nor U2689 (N_2689,N_1568,N_2164);
and U2690 (N_2690,N_2057,N_1927);
nand U2691 (N_2691,N_2110,N_1847);
nor U2692 (N_2692,N_2074,N_1761);
nand U2693 (N_2693,N_2078,N_1937);
nand U2694 (N_2694,N_2161,N_2190);
or U2695 (N_2695,N_2117,N_1994);
nor U2696 (N_2696,N_1867,N_1974);
xor U2697 (N_2697,N_2080,N_1833);
nor U2698 (N_2698,N_1968,N_2006);
xnor U2699 (N_2699,N_1509,N_1865);
nor U2700 (N_2700,N_1509,N_1706);
and U2701 (N_2701,N_1870,N_2079);
nor U2702 (N_2702,N_1699,N_2163);
and U2703 (N_2703,N_2210,N_2241);
nor U2704 (N_2704,N_1992,N_1820);
nand U2705 (N_2705,N_1906,N_2101);
nand U2706 (N_2706,N_1705,N_1757);
or U2707 (N_2707,N_1982,N_1589);
nand U2708 (N_2708,N_1583,N_2228);
nor U2709 (N_2709,N_1547,N_1926);
or U2710 (N_2710,N_2159,N_1609);
nor U2711 (N_2711,N_2112,N_1744);
or U2712 (N_2712,N_1808,N_2190);
or U2713 (N_2713,N_2111,N_1775);
or U2714 (N_2714,N_2078,N_1914);
nand U2715 (N_2715,N_1937,N_2141);
nand U2716 (N_2716,N_2020,N_1909);
or U2717 (N_2717,N_2100,N_1529);
or U2718 (N_2718,N_1707,N_2135);
and U2719 (N_2719,N_1764,N_1742);
and U2720 (N_2720,N_1886,N_1664);
and U2721 (N_2721,N_1886,N_1761);
or U2722 (N_2722,N_1957,N_1952);
nand U2723 (N_2723,N_2059,N_2187);
nor U2724 (N_2724,N_1721,N_2098);
or U2725 (N_2725,N_1646,N_1899);
or U2726 (N_2726,N_1838,N_2204);
nor U2727 (N_2727,N_2195,N_1722);
and U2728 (N_2728,N_1830,N_2245);
and U2729 (N_2729,N_1813,N_2023);
nand U2730 (N_2730,N_2077,N_1681);
xnor U2731 (N_2731,N_1895,N_1737);
nand U2732 (N_2732,N_1870,N_1608);
xor U2733 (N_2733,N_1895,N_2195);
nand U2734 (N_2734,N_2221,N_1657);
nand U2735 (N_2735,N_1809,N_1522);
and U2736 (N_2736,N_2049,N_2227);
nand U2737 (N_2737,N_1620,N_1933);
nand U2738 (N_2738,N_1513,N_1562);
nor U2739 (N_2739,N_1949,N_1969);
and U2740 (N_2740,N_1802,N_1511);
xor U2741 (N_2741,N_2080,N_2206);
and U2742 (N_2742,N_1971,N_2155);
nor U2743 (N_2743,N_1753,N_1776);
nor U2744 (N_2744,N_1735,N_2230);
nor U2745 (N_2745,N_2075,N_2242);
and U2746 (N_2746,N_1880,N_1733);
and U2747 (N_2747,N_1819,N_2043);
or U2748 (N_2748,N_1542,N_1903);
and U2749 (N_2749,N_1880,N_1943);
or U2750 (N_2750,N_1661,N_1510);
or U2751 (N_2751,N_1954,N_1996);
nand U2752 (N_2752,N_2157,N_1668);
and U2753 (N_2753,N_1738,N_1503);
nand U2754 (N_2754,N_1791,N_1623);
nand U2755 (N_2755,N_1548,N_1848);
and U2756 (N_2756,N_2005,N_1802);
and U2757 (N_2757,N_1593,N_1699);
nor U2758 (N_2758,N_2061,N_2144);
or U2759 (N_2759,N_1990,N_1549);
nor U2760 (N_2760,N_1882,N_1817);
and U2761 (N_2761,N_1540,N_2213);
nand U2762 (N_2762,N_1796,N_1912);
or U2763 (N_2763,N_1793,N_1542);
or U2764 (N_2764,N_1958,N_1795);
or U2765 (N_2765,N_1844,N_2004);
and U2766 (N_2766,N_1557,N_2247);
or U2767 (N_2767,N_2152,N_1507);
and U2768 (N_2768,N_1968,N_1853);
nor U2769 (N_2769,N_2205,N_1976);
and U2770 (N_2770,N_1596,N_2022);
nand U2771 (N_2771,N_1875,N_1890);
nand U2772 (N_2772,N_1731,N_1502);
nor U2773 (N_2773,N_1628,N_1536);
nor U2774 (N_2774,N_2067,N_2025);
nor U2775 (N_2775,N_1608,N_1860);
nor U2776 (N_2776,N_2090,N_1677);
nor U2777 (N_2777,N_2217,N_1844);
or U2778 (N_2778,N_2231,N_1935);
and U2779 (N_2779,N_1613,N_1636);
or U2780 (N_2780,N_1978,N_1609);
xnor U2781 (N_2781,N_1840,N_1516);
xor U2782 (N_2782,N_2162,N_1730);
nand U2783 (N_2783,N_2212,N_2206);
nand U2784 (N_2784,N_1825,N_2149);
and U2785 (N_2785,N_2004,N_2214);
nor U2786 (N_2786,N_2242,N_2188);
nor U2787 (N_2787,N_2236,N_1593);
nor U2788 (N_2788,N_1835,N_1516);
xnor U2789 (N_2789,N_1841,N_1858);
nand U2790 (N_2790,N_1615,N_1505);
xor U2791 (N_2791,N_1977,N_2212);
nand U2792 (N_2792,N_1998,N_1690);
nor U2793 (N_2793,N_1773,N_1822);
and U2794 (N_2794,N_1939,N_1966);
or U2795 (N_2795,N_2105,N_1949);
and U2796 (N_2796,N_1897,N_1821);
or U2797 (N_2797,N_1885,N_2113);
or U2798 (N_2798,N_1892,N_1802);
nand U2799 (N_2799,N_2014,N_2038);
and U2800 (N_2800,N_1975,N_1556);
and U2801 (N_2801,N_1566,N_1997);
and U2802 (N_2802,N_2178,N_1839);
nand U2803 (N_2803,N_1542,N_1981);
nor U2804 (N_2804,N_1907,N_1937);
and U2805 (N_2805,N_2191,N_1545);
or U2806 (N_2806,N_2239,N_1911);
xnor U2807 (N_2807,N_1718,N_1974);
nand U2808 (N_2808,N_2099,N_2035);
xor U2809 (N_2809,N_2211,N_1996);
and U2810 (N_2810,N_1969,N_1509);
and U2811 (N_2811,N_1565,N_1683);
nor U2812 (N_2812,N_1928,N_2076);
nand U2813 (N_2813,N_2182,N_2207);
nand U2814 (N_2814,N_2034,N_1902);
or U2815 (N_2815,N_1748,N_1560);
nand U2816 (N_2816,N_1613,N_1677);
nand U2817 (N_2817,N_1794,N_2019);
nor U2818 (N_2818,N_1569,N_2225);
nand U2819 (N_2819,N_1810,N_2076);
and U2820 (N_2820,N_1736,N_1925);
xor U2821 (N_2821,N_1668,N_1892);
or U2822 (N_2822,N_1514,N_1543);
and U2823 (N_2823,N_2003,N_2072);
or U2824 (N_2824,N_1792,N_1885);
nand U2825 (N_2825,N_2238,N_1961);
and U2826 (N_2826,N_1783,N_2205);
and U2827 (N_2827,N_1946,N_1813);
nand U2828 (N_2828,N_1606,N_2140);
nor U2829 (N_2829,N_2123,N_1501);
or U2830 (N_2830,N_1675,N_1833);
nand U2831 (N_2831,N_1992,N_1787);
and U2832 (N_2832,N_1964,N_2109);
and U2833 (N_2833,N_1658,N_1592);
nor U2834 (N_2834,N_1682,N_1685);
nand U2835 (N_2835,N_2096,N_1516);
or U2836 (N_2836,N_2186,N_1853);
nand U2837 (N_2837,N_1864,N_1794);
nand U2838 (N_2838,N_2217,N_1639);
nor U2839 (N_2839,N_1731,N_1896);
and U2840 (N_2840,N_1969,N_1809);
or U2841 (N_2841,N_1506,N_2202);
nor U2842 (N_2842,N_2127,N_2145);
or U2843 (N_2843,N_1731,N_1779);
nor U2844 (N_2844,N_1825,N_1929);
or U2845 (N_2845,N_1966,N_1510);
or U2846 (N_2846,N_1958,N_1998);
nand U2847 (N_2847,N_1668,N_1882);
or U2848 (N_2848,N_2004,N_2187);
xnor U2849 (N_2849,N_1526,N_1524);
nand U2850 (N_2850,N_1888,N_2041);
or U2851 (N_2851,N_2121,N_2187);
nand U2852 (N_2852,N_1727,N_2158);
and U2853 (N_2853,N_2205,N_1748);
and U2854 (N_2854,N_1919,N_1642);
nand U2855 (N_2855,N_2170,N_1657);
nor U2856 (N_2856,N_1937,N_2064);
and U2857 (N_2857,N_1798,N_1751);
or U2858 (N_2858,N_1965,N_1642);
and U2859 (N_2859,N_1538,N_1941);
or U2860 (N_2860,N_1576,N_1951);
nor U2861 (N_2861,N_2031,N_1836);
nor U2862 (N_2862,N_1981,N_1916);
nand U2863 (N_2863,N_2022,N_1893);
nand U2864 (N_2864,N_2010,N_1922);
nand U2865 (N_2865,N_2095,N_1569);
nand U2866 (N_2866,N_1780,N_1790);
and U2867 (N_2867,N_1863,N_2023);
or U2868 (N_2868,N_1867,N_1631);
nand U2869 (N_2869,N_1963,N_2044);
nor U2870 (N_2870,N_1816,N_1894);
or U2871 (N_2871,N_1870,N_2242);
nand U2872 (N_2872,N_2094,N_1801);
and U2873 (N_2873,N_1978,N_1998);
nor U2874 (N_2874,N_2225,N_1719);
nor U2875 (N_2875,N_1937,N_1966);
xor U2876 (N_2876,N_2098,N_1736);
or U2877 (N_2877,N_2101,N_2121);
and U2878 (N_2878,N_1889,N_2199);
and U2879 (N_2879,N_2101,N_1655);
nor U2880 (N_2880,N_1854,N_1795);
and U2881 (N_2881,N_1564,N_1581);
nor U2882 (N_2882,N_1632,N_1649);
xor U2883 (N_2883,N_2232,N_1930);
nand U2884 (N_2884,N_1870,N_1857);
and U2885 (N_2885,N_1933,N_2080);
xnor U2886 (N_2886,N_2017,N_1620);
or U2887 (N_2887,N_1841,N_1871);
or U2888 (N_2888,N_1955,N_1592);
nor U2889 (N_2889,N_1930,N_1791);
or U2890 (N_2890,N_1670,N_2068);
and U2891 (N_2891,N_1504,N_1875);
and U2892 (N_2892,N_1803,N_1822);
nand U2893 (N_2893,N_1762,N_1858);
or U2894 (N_2894,N_1573,N_2155);
and U2895 (N_2895,N_1667,N_1639);
and U2896 (N_2896,N_1722,N_1563);
and U2897 (N_2897,N_2169,N_2071);
and U2898 (N_2898,N_1713,N_1884);
xor U2899 (N_2899,N_2102,N_1970);
xnor U2900 (N_2900,N_1908,N_2236);
nor U2901 (N_2901,N_1837,N_2230);
or U2902 (N_2902,N_1896,N_2017);
and U2903 (N_2903,N_2247,N_1696);
xnor U2904 (N_2904,N_2074,N_2159);
nand U2905 (N_2905,N_1919,N_1574);
nand U2906 (N_2906,N_2107,N_1984);
nand U2907 (N_2907,N_2019,N_1795);
xnor U2908 (N_2908,N_1864,N_1672);
or U2909 (N_2909,N_1844,N_1508);
nand U2910 (N_2910,N_1924,N_1721);
xnor U2911 (N_2911,N_1946,N_1801);
nand U2912 (N_2912,N_1885,N_1508);
and U2913 (N_2913,N_1557,N_1538);
nand U2914 (N_2914,N_1648,N_2096);
and U2915 (N_2915,N_1720,N_1901);
nand U2916 (N_2916,N_2002,N_2241);
nor U2917 (N_2917,N_1717,N_2032);
or U2918 (N_2918,N_1668,N_2247);
nand U2919 (N_2919,N_2015,N_1759);
or U2920 (N_2920,N_2159,N_1748);
or U2921 (N_2921,N_1617,N_1579);
nand U2922 (N_2922,N_1637,N_1713);
nand U2923 (N_2923,N_2175,N_1693);
and U2924 (N_2924,N_1650,N_2095);
and U2925 (N_2925,N_1685,N_1681);
or U2926 (N_2926,N_2227,N_1862);
xor U2927 (N_2927,N_1744,N_2071);
xnor U2928 (N_2928,N_1887,N_1955);
and U2929 (N_2929,N_2087,N_2065);
nor U2930 (N_2930,N_1649,N_1781);
and U2931 (N_2931,N_2009,N_1655);
nor U2932 (N_2932,N_2159,N_1777);
nor U2933 (N_2933,N_1716,N_1867);
nand U2934 (N_2934,N_2149,N_2012);
nand U2935 (N_2935,N_2162,N_2198);
nor U2936 (N_2936,N_1900,N_1771);
nor U2937 (N_2937,N_1572,N_1641);
and U2938 (N_2938,N_1717,N_1841);
or U2939 (N_2939,N_1568,N_1889);
or U2940 (N_2940,N_1885,N_1604);
and U2941 (N_2941,N_2114,N_1668);
xor U2942 (N_2942,N_2168,N_2042);
nand U2943 (N_2943,N_1703,N_1637);
and U2944 (N_2944,N_2030,N_2014);
or U2945 (N_2945,N_2231,N_2196);
nor U2946 (N_2946,N_1505,N_2152);
nor U2947 (N_2947,N_1753,N_1858);
nand U2948 (N_2948,N_1796,N_2087);
nand U2949 (N_2949,N_1875,N_1567);
nand U2950 (N_2950,N_1644,N_2215);
and U2951 (N_2951,N_1669,N_2137);
and U2952 (N_2952,N_2098,N_1975);
xor U2953 (N_2953,N_1889,N_1934);
nand U2954 (N_2954,N_1546,N_1678);
and U2955 (N_2955,N_1575,N_1972);
nor U2956 (N_2956,N_1789,N_1656);
xnor U2957 (N_2957,N_1887,N_2161);
nand U2958 (N_2958,N_1939,N_2001);
and U2959 (N_2959,N_1958,N_1685);
nand U2960 (N_2960,N_2018,N_1861);
and U2961 (N_2961,N_1784,N_1519);
or U2962 (N_2962,N_1876,N_1671);
nand U2963 (N_2963,N_1961,N_1599);
nand U2964 (N_2964,N_1990,N_1649);
or U2965 (N_2965,N_1508,N_1769);
or U2966 (N_2966,N_2105,N_1827);
nand U2967 (N_2967,N_2187,N_2098);
or U2968 (N_2968,N_1971,N_2010);
or U2969 (N_2969,N_2046,N_1740);
nand U2970 (N_2970,N_1626,N_2070);
nor U2971 (N_2971,N_1581,N_2207);
xnor U2972 (N_2972,N_1716,N_1615);
nor U2973 (N_2973,N_1709,N_1984);
or U2974 (N_2974,N_1849,N_1589);
nor U2975 (N_2975,N_1786,N_1969);
xnor U2976 (N_2976,N_1542,N_1640);
nand U2977 (N_2977,N_1521,N_2189);
or U2978 (N_2978,N_1796,N_2244);
and U2979 (N_2979,N_1531,N_2057);
and U2980 (N_2980,N_1990,N_1639);
nand U2981 (N_2981,N_2114,N_1749);
and U2982 (N_2982,N_1985,N_2032);
and U2983 (N_2983,N_1781,N_1601);
nor U2984 (N_2984,N_2043,N_2113);
or U2985 (N_2985,N_1508,N_2130);
and U2986 (N_2986,N_1955,N_2043);
nand U2987 (N_2987,N_2222,N_1691);
or U2988 (N_2988,N_2023,N_2198);
nor U2989 (N_2989,N_1964,N_1790);
and U2990 (N_2990,N_2194,N_1745);
or U2991 (N_2991,N_1767,N_2016);
nand U2992 (N_2992,N_2153,N_2170);
nand U2993 (N_2993,N_2090,N_1867);
nor U2994 (N_2994,N_1895,N_1970);
and U2995 (N_2995,N_1833,N_2082);
or U2996 (N_2996,N_1727,N_2106);
or U2997 (N_2997,N_2113,N_1525);
xor U2998 (N_2998,N_1778,N_1800);
nand U2999 (N_2999,N_1504,N_1910);
nor U3000 (N_3000,N_2851,N_2373);
xnor U3001 (N_3001,N_2385,N_2926);
and U3002 (N_3002,N_2308,N_2407);
and U3003 (N_3003,N_2590,N_2299);
and U3004 (N_3004,N_2670,N_2597);
nor U3005 (N_3005,N_2493,N_2434);
or U3006 (N_3006,N_2560,N_2591);
nor U3007 (N_3007,N_2883,N_2819);
nand U3008 (N_3008,N_2963,N_2980);
and U3009 (N_3009,N_2947,N_2262);
nor U3010 (N_3010,N_2632,N_2577);
nand U3011 (N_3011,N_2619,N_2635);
xnor U3012 (N_3012,N_2456,N_2664);
and U3013 (N_3013,N_2368,N_2302);
nor U3014 (N_3014,N_2773,N_2985);
nand U3015 (N_3015,N_2854,N_2379);
or U3016 (N_3016,N_2486,N_2604);
and U3017 (N_3017,N_2370,N_2537);
xnor U3018 (N_3018,N_2827,N_2957);
nand U3019 (N_3019,N_2720,N_2575);
xor U3020 (N_3020,N_2975,N_2551);
nor U3021 (N_3021,N_2607,N_2718);
or U3022 (N_3022,N_2406,N_2991);
nor U3023 (N_3023,N_2319,N_2504);
nand U3024 (N_3024,N_2335,N_2918);
or U3025 (N_3025,N_2982,N_2450);
nor U3026 (N_3026,N_2367,N_2789);
nand U3027 (N_3027,N_2608,N_2453);
or U3028 (N_3028,N_2275,N_2512);
and U3029 (N_3029,N_2655,N_2998);
nand U3030 (N_3030,N_2618,N_2436);
and U3031 (N_3031,N_2557,N_2993);
nand U3032 (N_3032,N_2818,N_2855);
or U3033 (N_3033,N_2836,N_2609);
xor U3034 (N_3034,N_2476,N_2558);
or U3035 (N_3035,N_2904,N_2555);
and U3036 (N_3036,N_2972,N_2936);
nor U3037 (N_3037,N_2938,N_2573);
or U3038 (N_3038,N_2441,N_2853);
and U3039 (N_3039,N_2790,N_2509);
or U3040 (N_3040,N_2382,N_2674);
or U3041 (N_3041,N_2268,N_2584);
nor U3042 (N_3042,N_2812,N_2890);
or U3043 (N_3043,N_2580,N_2873);
and U3044 (N_3044,N_2876,N_2333);
and U3045 (N_3045,N_2704,N_2317);
or U3046 (N_3046,N_2990,N_2857);
nand U3047 (N_3047,N_2538,N_2387);
or U3048 (N_3048,N_2606,N_2878);
nand U3049 (N_3049,N_2426,N_2347);
and U3050 (N_3050,N_2359,N_2399);
nand U3051 (N_3051,N_2658,N_2971);
nor U3052 (N_3052,N_2381,N_2907);
nor U3053 (N_3053,N_2893,N_2772);
nand U3054 (N_3054,N_2973,N_2517);
nor U3055 (N_3055,N_2711,N_2432);
nand U3056 (N_3056,N_2375,N_2523);
nand U3057 (N_3057,N_2542,N_2826);
or U3058 (N_3058,N_2532,N_2384);
or U3059 (N_3059,N_2657,N_2752);
or U3060 (N_3060,N_2461,N_2395);
or U3061 (N_3061,N_2277,N_2933);
xnor U3062 (N_3062,N_2910,N_2321);
or U3063 (N_3063,N_2847,N_2294);
and U3064 (N_3064,N_2948,N_2968);
nand U3065 (N_3065,N_2688,N_2997);
xor U3066 (N_3066,N_2912,N_2735);
and U3067 (N_3067,N_2462,N_2895);
nand U3068 (N_3068,N_2874,N_2653);
or U3069 (N_3069,N_2411,N_2334);
or U3070 (N_3070,N_2499,N_2686);
nor U3071 (N_3071,N_2964,N_2842);
nand U3072 (N_3072,N_2626,N_2760);
or U3073 (N_3073,N_2543,N_2640);
nand U3074 (N_3074,N_2502,N_2482);
nand U3075 (N_3075,N_2516,N_2297);
or U3076 (N_3076,N_2679,N_2746);
nor U3077 (N_3077,N_2736,N_2872);
nor U3078 (N_3078,N_2738,N_2312);
nor U3079 (N_3079,N_2977,N_2780);
nor U3080 (N_3080,N_2505,N_2937);
nand U3081 (N_3081,N_2293,N_2860);
xnor U3082 (N_3082,N_2298,N_2729);
or U3083 (N_3083,N_2917,N_2324);
nor U3084 (N_3084,N_2898,N_2353);
nand U3085 (N_3085,N_2750,N_2545);
or U3086 (N_3086,N_2452,N_2583);
or U3087 (N_3087,N_2613,N_2371);
nand U3088 (N_3088,N_2341,N_2565);
and U3089 (N_3089,N_2496,N_2338);
nand U3090 (N_3090,N_2749,N_2783);
and U3091 (N_3091,N_2322,N_2465);
nand U3092 (N_3092,N_2392,N_2848);
nand U3093 (N_3093,N_2548,N_2942);
and U3094 (N_3094,N_2721,N_2634);
nand U3095 (N_3095,N_2908,N_2582);
nand U3096 (N_3096,N_2377,N_2472);
and U3097 (N_3097,N_2801,N_2984);
nand U3098 (N_3098,N_2571,N_2497);
nor U3099 (N_3099,N_2285,N_2253);
nand U3100 (N_3100,N_2800,N_2273);
and U3101 (N_3101,N_2956,N_2845);
and U3102 (N_3102,N_2650,N_2739);
nand U3103 (N_3103,N_2405,N_2612);
or U3104 (N_3104,N_2627,N_2888);
and U3105 (N_3105,N_2727,N_2578);
and U3106 (N_3106,N_2471,N_2394);
xnor U3107 (N_3107,N_2306,N_2362);
and U3108 (N_3108,N_2336,N_2445);
or U3109 (N_3109,N_2420,N_2741);
and U3110 (N_3110,N_2447,N_2556);
and U3111 (N_3111,N_2771,N_2320);
nand U3112 (N_3112,N_2266,N_2871);
or U3113 (N_3113,N_2702,N_2289);
nand U3114 (N_3114,N_2553,N_2965);
nand U3115 (N_3115,N_2389,N_2717);
and U3116 (N_3116,N_2858,N_2882);
or U3117 (N_3117,N_2398,N_2979);
xnor U3118 (N_3118,N_2255,N_2962);
and U3119 (N_3119,N_2498,N_2519);
xnor U3120 (N_3120,N_2552,N_2374);
nor U3121 (N_3121,N_2707,N_2564);
or U3122 (N_3122,N_2680,N_2601);
nor U3123 (N_3123,N_2383,N_2403);
or U3124 (N_3124,N_2342,N_2929);
nor U3125 (N_3125,N_2615,N_2326);
nor U3126 (N_3126,N_2649,N_2391);
nand U3127 (N_3127,N_2891,N_2574);
nand U3128 (N_3128,N_2410,N_2969);
xor U3129 (N_3129,N_2678,N_2660);
nand U3130 (N_3130,N_2559,N_2814);
and U3131 (N_3131,N_2799,N_2927);
and U3132 (N_3132,N_2614,N_2313);
xor U3133 (N_3133,N_2838,N_2753);
xor U3134 (N_3134,N_2837,N_2596);
and U3135 (N_3135,N_2828,N_2880);
xnor U3136 (N_3136,N_2911,N_2251);
or U3137 (N_3137,N_2380,N_2639);
xor U3138 (N_3138,N_2781,N_2572);
nand U3139 (N_3139,N_2585,N_2343);
and U3140 (N_3140,N_2784,N_2340);
nand U3141 (N_3141,N_2446,N_2743);
nor U3142 (N_3142,N_2633,N_2843);
nor U3143 (N_3143,N_2501,N_2526);
or U3144 (N_3144,N_2386,N_2284);
or U3145 (N_3145,N_2327,N_2355);
nand U3146 (N_3146,N_2346,N_2349);
and U3147 (N_3147,N_2372,N_2654);
and U3148 (N_3148,N_2744,N_2408);
and U3149 (N_3149,N_2598,N_2357);
nor U3150 (N_3150,N_2835,N_2464);
xor U3151 (N_3151,N_2805,N_2413);
xor U3152 (N_3152,N_2409,N_2731);
and U3153 (N_3153,N_2282,N_2943);
xnor U3154 (N_3154,N_2989,N_2666);
or U3155 (N_3155,N_2323,N_2378);
nand U3156 (N_3156,N_2494,N_2762);
and U3157 (N_3157,N_2265,N_2276);
or U3158 (N_3158,N_2622,N_2659);
nor U3159 (N_3159,N_2288,N_2491);
nor U3160 (N_3160,N_2316,N_2777);
and U3161 (N_3161,N_2473,N_2528);
xnor U3162 (N_3162,N_2388,N_2460);
nand U3163 (N_3163,N_2468,N_2899);
xor U3164 (N_3164,N_2694,N_2987);
and U3165 (N_3165,N_2879,N_2850);
nor U3166 (N_3166,N_2280,N_2624);
and U3167 (N_3167,N_2592,N_2539);
and U3168 (N_3168,N_2719,N_2797);
nand U3169 (N_3169,N_2529,N_2258);
nor U3170 (N_3170,N_2867,N_2648);
and U3171 (N_3171,N_2747,N_2569);
nor U3172 (N_3172,N_2424,N_2810);
nor U3173 (N_3173,N_2617,N_2562);
and U3174 (N_3174,N_2960,N_2546);
nor U3175 (N_3175,N_2830,N_2300);
or U3176 (N_3176,N_2934,N_2687);
and U3177 (N_3177,N_2806,N_2976);
nand U3178 (N_3178,N_2820,N_2250);
nor U3179 (N_3179,N_2438,N_2791);
xor U3180 (N_3180,N_2514,N_2671);
nor U3181 (N_3181,N_2390,N_2522);
and U3182 (N_3182,N_2602,N_2595);
xor U3183 (N_3183,N_2787,N_2412);
nand U3184 (N_3184,N_2986,N_2260);
and U3185 (N_3185,N_2682,N_2715);
or U3186 (N_3186,N_2629,N_2396);
and U3187 (N_3187,N_2541,N_2896);
nor U3188 (N_3188,N_2701,N_2520);
nand U3189 (N_3189,N_2647,N_2939);
nor U3190 (N_3190,N_2621,N_2315);
nor U3191 (N_3191,N_2710,N_2841);
and U3192 (N_3192,N_2903,N_2885);
or U3193 (N_3193,N_2568,N_2834);
and U3194 (N_3194,N_2822,N_2274);
nor U3195 (N_3195,N_2970,N_2278);
or U3196 (N_3196,N_2469,N_2605);
nor U3197 (N_3197,N_2946,N_2974);
or U3198 (N_3198,N_2511,N_2803);
nor U3199 (N_3199,N_2515,N_2570);
and U3200 (N_3200,N_2713,N_2492);
xnor U3201 (N_3201,N_2796,N_2625);
or U3202 (N_3202,N_2485,N_2610);
xnor U3203 (N_3203,N_2536,N_2795);
and U3204 (N_3204,N_2429,N_2863);
nor U3205 (N_3205,N_2906,N_2350);
nor U3206 (N_3206,N_2292,N_2466);
and U3207 (N_3207,N_2716,N_2695);
nand U3208 (N_3208,N_2839,N_2593);
and U3209 (N_3209,N_2667,N_2495);
nor U3210 (N_3210,N_2478,N_2951);
nand U3211 (N_3211,N_2920,N_2527);
nor U3212 (N_3212,N_2698,N_2270);
nand U3213 (N_3213,N_2281,N_2488);
xnor U3214 (N_3214,N_2978,N_2700);
or U3215 (N_3215,N_2849,N_2474);
or U3216 (N_3216,N_2475,N_2755);
xnor U3217 (N_3217,N_2547,N_2561);
or U3218 (N_3218,N_2508,N_2661);
or U3219 (N_3219,N_2865,N_2269);
and U3220 (N_3220,N_2706,N_2430);
nand U3221 (N_3221,N_2870,N_2534);
and U3222 (N_3222,N_2919,N_2480);
xor U3223 (N_3223,N_2877,N_2345);
nand U3224 (N_3224,N_2643,N_2483);
nor U3225 (N_3225,N_2490,N_2628);
nand U3226 (N_3226,N_2369,N_2813);
and U3227 (N_3227,N_2959,N_2677);
and U3228 (N_3228,N_2665,N_2914);
nor U3229 (N_3229,N_2309,N_2256);
and U3230 (N_3230,N_2301,N_2623);
or U3231 (N_3231,N_2861,N_2786);
or U3232 (N_3232,N_2354,N_2524);
and U3233 (N_3233,N_2785,N_2272);
nor U3234 (N_3234,N_2815,N_2846);
and U3235 (N_3235,N_2563,N_2449);
or U3236 (N_3236,N_2440,N_2988);
or U3237 (N_3237,N_2435,N_2763);
xor U3238 (N_3238,N_2756,N_2966);
nand U3239 (N_3239,N_2588,N_2332);
or U3240 (N_3240,N_2689,N_2905);
and U3241 (N_3241,N_2533,N_2808);
nor U3242 (N_3242,N_2685,N_2360);
or U3243 (N_3243,N_2467,N_2458);
or U3244 (N_3244,N_2656,N_2587);
xnor U3245 (N_3245,N_2669,N_2824);
and U3246 (N_3246,N_2931,N_2924);
nand U3247 (N_3247,N_2454,N_2544);
nand U3248 (N_3248,N_2376,N_2697);
xnor U3249 (N_3249,N_2699,N_2645);
and U3250 (N_3250,N_2287,N_2603);
nand U3251 (N_3251,N_2804,N_2922);
and U3252 (N_3252,N_2792,N_2404);
nor U3253 (N_3253,N_2616,N_2897);
xnor U3254 (N_3254,N_2310,N_2887);
xor U3255 (N_3255,N_2952,N_2489);
nand U3256 (N_3256,N_2257,N_2337);
and U3257 (N_3257,N_2642,N_2503);
nor U3258 (N_3258,N_2894,N_2892);
or U3259 (N_3259,N_2477,N_2881);
nand U3260 (N_3260,N_2550,N_2766);
nand U3261 (N_3261,N_2733,N_2296);
nor U3262 (N_3262,N_2856,N_2869);
nand U3263 (N_3263,N_2611,N_2705);
nor U3264 (N_3264,N_2983,N_2295);
or U3265 (N_3265,N_2829,N_2330);
xor U3266 (N_3266,N_2339,N_2932);
and U3267 (N_3267,N_2646,N_2428);
and U3268 (N_3268,N_2443,N_2751);
nand U3269 (N_3269,N_2402,N_2651);
or U3270 (N_3270,N_2817,N_2431);
nand U3271 (N_3271,N_2261,N_2949);
and U3272 (N_3272,N_2442,N_2459);
or U3273 (N_3273,N_2364,N_2684);
or U3274 (N_3274,N_2400,N_2290);
or U3275 (N_3275,N_2994,N_2305);
nand U3276 (N_3276,N_2708,N_2866);
nor U3277 (N_3277,N_2513,N_2271);
xor U3278 (N_3278,N_2692,N_2567);
nor U3279 (N_3279,N_2637,N_2311);
xor U3280 (N_3280,N_2267,N_2254);
and U3281 (N_3281,N_2525,N_2868);
or U3282 (N_3282,N_2900,N_2955);
and U3283 (N_3283,N_2945,N_2832);
or U3284 (N_3284,N_2728,N_2793);
nor U3285 (N_3285,N_2652,N_2352);
or U3286 (N_3286,N_2967,N_2314);
and U3287 (N_3287,N_2875,N_2416);
or U3288 (N_3288,N_2725,N_2630);
nand U3289 (N_3289,N_2506,N_2307);
and U3290 (N_3290,N_2500,N_2530);
and U3291 (N_3291,N_2798,N_2864);
and U3292 (N_3292,N_2916,N_2852);
and U3293 (N_3293,N_2775,N_2930);
nor U3294 (N_3294,N_2999,N_2778);
nor U3295 (N_3295,N_2414,N_2809);
nand U3296 (N_3296,N_2745,N_2724);
or U3297 (N_3297,N_2693,N_2318);
nor U3298 (N_3298,N_2779,N_2279);
xnor U3299 (N_3299,N_2363,N_2953);
and U3300 (N_3300,N_2992,N_2662);
nor U3301 (N_3301,N_2726,N_2788);
nand U3302 (N_3302,N_2833,N_2366);
xnor U3303 (N_3303,N_2549,N_2954);
or U3304 (N_3304,N_2831,N_2862);
nor U3305 (N_3305,N_2518,N_2393);
nor U3306 (N_3306,N_2740,N_2764);
xnor U3307 (N_3307,N_2510,N_2487);
nor U3308 (N_3308,N_2397,N_2770);
and U3309 (N_3309,N_2884,N_2676);
nand U3310 (N_3310,N_2263,N_2419);
and U3311 (N_3311,N_2507,N_2748);
nand U3312 (N_3312,N_2811,N_2673);
and U3313 (N_3313,N_2644,N_2737);
xor U3314 (N_3314,N_2958,N_2641);
and U3315 (N_3315,N_2636,N_2423);
nand U3316 (N_3316,N_2291,N_2540);
nor U3317 (N_3317,N_2925,N_2754);
or U3318 (N_3318,N_2928,N_2995);
nor U3319 (N_3319,N_2709,N_2821);
and U3320 (N_3320,N_2663,N_2586);
nand U3321 (N_3321,N_2767,N_2734);
and U3322 (N_3322,N_2470,N_2825);
and U3323 (N_3323,N_2361,N_2921);
nand U3324 (N_3324,N_2631,N_2768);
or U3325 (N_3325,N_2742,N_2283);
nor U3326 (N_3326,N_2807,N_2448);
nand U3327 (N_3327,N_2484,N_2913);
xor U3328 (N_3328,N_2433,N_2981);
nand U3329 (N_3329,N_2421,N_2479);
xor U3330 (N_3330,N_2759,N_2437);
or U3331 (N_3331,N_2422,N_2840);
and U3332 (N_3332,N_2286,N_2365);
nor U3333 (N_3333,N_2451,N_2304);
nor U3334 (N_3334,N_2769,N_2535);
xor U3335 (N_3335,N_2901,N_2599);
nand U3336 (N_3336,N_2259,N_2455);
and U3337 (N_3337,N_2329,N_2765);
xor U3338 (N_3338,N_2696,N_2417);
nand U3339 (N_3339,N_2776,N_2774);
xor U3340 (N_3340,N_2579,N_2427);
nor U3341 (N_3341,N_2802,N_2714);
and U3342 (N_3342,N_2344,N_2672);
nor U3343 (N_3343,N_2909,N_2521);
nand U3344 (N_3344,N_2668,N_2600);
and U3345 (N_3345,N_2566,N_2844);
or U3346 (N_3346,N_2594,N_2794);
nand U3347 (N_3347,N_2620,N_2444);
nand U3348 (N_3348,N_2358,N_2439);
nand U3349 (N_3349,N_2712,N_2418);
and U3350 (N_3350,N_2859,N_2425);
nand U3351 (N_3351,N_2457,N_2531);
nor U3352 (N_3352,N_2356,N_2481);
nand U3353 (N_3353,N_2940,N_2554);
nand U3354 (N_3354,N_2691,N_2681);
xnor U3355 (N_3355,N_2703,N_2328);
nor U3356 (N_3356,N_2252,N_2816);
nor U3357 (N_3357,N_2732,N_2675);
and U3358 (N_3358,N_2941,N_2722);
xor U3359 (N_3359,N_2758,N_2638);
or U3360 (N_3360,N_2576,N_2923);
nand U3361 (N_3361,N_2348,N_2902);
or U3362 (N_3362,N_2823,N_2723);
nor U3363 (N_3363,N_2730,N_2690);
xnor U3364 (N_3364,N_2961,N_2401);
nand U3365 (N_3365,N_2683,N_2331);
xor U3366 (N_3366,N_2303,N_2351);
nand U3367 (N_3367,N_2589,N_2950);
nand U3368 (N_3368,N_2889,N_2935);
and U3369 (N_3369,N_2782,N_2325);
or U3370 (N_3370,N_2996,N_2757);
nor U3371 (N_3371,N_2944,N_2415);
nor U3372 (N_3372,N_2886,N_2264);
and U3373 (N_3373,N_2915,N_2463);
xnor U3374 (N_3374,N_2581,N_2761);
nand U3375 (N_3375,N_2566,N_2717);
xor U3376 (N_3376,N_2699,N_2443);
or U3377 (N_3377,N_2717,N_2333);
nor U3378 (N_3378,N_2965,N_2895);
nand U3379 (N_3379,N_2687,N_2355);
xnor U3380 (N_3380,N_2341,N_2949);
xnor U3381 (N_3381,N_2582,N_2750);
or U3382 (N_3382,N_2599,N_2771);
xnor U3383 (N_3383,N_2285,N_2801);
xnor U3384 (N_3384,N_2999,N_2885);
or U3385 (N_3385,N_2787,N_2256);
or U3386 (N_3386,N_2918,N_2396);
xnor U3387 (N_3387,N_2406,N_2949);
or U3388 (N_3388,N_2443,N_2400);
nand U3389 (N_3389,N_2997,N_2947);
nand U3390 (N_3390,N_2438,N_2849);
nor U3391 (N_3391,N_2961,N_2708);
or U3392 (N_3392,N_2440,N_2975);
nand U3393 (N_3393,N_2272,N_2424);
and U3394 (N_3394,N_2540,N_2633);
or U3395 (N_3395,N_2312,N_2411);
nand U3396 (N_3396,N_2949,N_2304);
nand U3397 (N_3397,N_2469,N_2993);
nor U3398 (N_3398,N_2461,N_2317);
nor U3399 (N_3399,N_2499,N_2393);
and U3400 (N_3400,N_2557,N_2380);
nor U3401 (N_3401,N_2406,N_2681);
nand U3402 (N_3402,N_2424,N_2283);
nor U3403 (N_3403,N_2284,N_2845);
nand U3404 (N_3404,N_2844,N_2416);
or U3405 (N_3405,N_2316,N_2611);
or U3406 (N_3406,N_2310,N_2272);
nor U3407 (N_3407,N_2673,N_2774);
and U3408 (N_3408,N_2961,N_2853);
or U3409 (N_3409,N_2648,N_2984);
xnor U3410 (N_3410,N_2641,N_2832);
nor U3411 (N_3411,N_2305,N_2838);
xor U3412 (N_3412,N_2626,N_2676);
or U3413 (N_3413,N_2560,N_2644);
nor U3414 (N_3414,N_2446,N_2536);
xnor U3415 (N_3415,N_2521,N_2687);
and U3416 (N_3416,N_2491,N_2321);
nor U3417 (N_3417,N_2316,N_2292);
and U3418 (N_3418,N_2929,N_2595);
and U3419 (N_3419,N_2540,N_2759);
nand U3420 (N_3420,N_2699,N_2639);
nor U3421 (N_3421,N_2352,N_2275);
or U3422 (N_3422,N_2409,N_2919);
and U3423 (N_3423,N_2976,N_2698);
nand U3424 (N_3424,N_2485,N_2891);
or U3425 (N_3425,N_2554,N_2776);
xnor U3426 (N_3426,N_2312,N_2340);
and U3427 (N_3427,N_2571,N_2446);
nor U3428 (N_3428,N_2369,N_2525);
and U3429 (N_3429,N_2748,N_2772);
or U3430 (N_3430,N_2476,N_2657);
nor U3431 (N_3431,N_2863,N_2978);
nor U3432 (N_3432,N_2330,N_2519);
nor U3433 (N_3433,N_2531,N_2704);
and U3434 (N_3434,N_2711,N_2809);
or U3435 (N_3435,N_2570,N_2824);
xor U3436 (N_3436,N_2535,N_2523);
nand U3437 (N_3437,N_2902,N_2598);
nand U3438 (N_3438,N_2628,N_2336);
or U3439 (N_3439,N_2376,N_2367);
nand U3440 (N_3440,N_2799,N_2560);
nor U3441 (N_3441,N_2671,N_2462);
or U3442 (N_3442,N_2767,N_2800);
and U3443 (N_3443,N_2481,N_2899);
nor U3444 (N_3444,N_2704,N_2963);
nor U3445 (N_3445,N_2382,N_2566);
xnor U3446 (N_3446,N_2676,N_2353);
and U3447 (N_3447,N_2485,N_2704);
nand U3448 (N_3448,N_2905,N_2398);
nor U3449 (N_3449,N_2615,N_2985);
xnor U3450 (N_3450,N_2455,N_2891);
xor U3451 (N_3451,N_2404,N_2857);
or U3452 (N_3452,N_2831,N_2586);
nand U3453 (N_3453,N_2716,N_2916);
nor U3454 (N_3454,N_2764,N_2613);
nand U3455 (N_3455,N_2698,N_2881);
nand U3456 (N_3456,N_2674,N_2412);
and U3457 (N_3457,N_2698,N_2906);
nor U3458 (N_3458,N_2841,N_2265);
nand U3459 (N_3459,N_2976,N_2476);
or U3460 (N_3460,N_2297,N_2920);
nand U3461 (N_3461,N_2748,N_2639);
nand U3462 (N_3462,N_2401,N_2742);
xor U3463 (N_3463,N_2756,N_2450);
and U3464 (N_3464,N_2362,N_2998);
xnor U3465 (N_3465,N_2297,N_2401);
nand U3466 (N_3466,N_2658,N_2462);
and U3467 (N_3467,N_2353,N_2762);
and U3468 (N_3468,N_2743,N_2853);
nand U3469 (N_3469,N_2656,N_2299);
nor U3470 (N_3470,N_2934,N_2935);
nor U3471 (N_3471,N_2996,N_2699);
nor U3472 (N_3472,N_2358,N_2816);
xnor U3473 (N_3473,N_2899,N_2367);
nand U3474 (N_3474,N_2255,N_2809);
and U3475 (N_3475,N_2570,N_2309);
nor U3476 (N_3476,N_2501,N_2872);
and U3477 (N_3477,N_2742,N_2333);
and U3478 (N_3478,N_2913,N_2312);
xor U3479 (N_3479,N_2930,N_2881);
or U3480 (N_3480,N_2518,N_2964);
and U3481 (N_3481,N_2546,N_2793);
nor U3482 (N_3482,N_2639,N_2989);
and U3483 (N_3483,N_2420,N_2788);
nand U3484 (N_3484,N_2389,N_2998);
or U3485 (N_3485,N_2937,N_2673);
and U3486 (N_3486,N_2785,N_2400);
or U3487 (N_3487,N_2525,N_2636);
nor U3488 (N_3488,N_2635,N_2599);
and U3489 (N_3489,N_2336,N_2666);
nand U3490 (N_3490,N_2993,N_2446);
and U3491 (N_3491,N_2809,N_2518);
and U3492 (N_3492,N_2679,N_2955);
and U3493 (N_3493,N_2674,N_2337);
and U3494 (N_3494,N_2275,N_2932);
and U3495 (N_3495,N_2490,N_2955);
and U3496 (N_3496,N_2914,N_2667);
nand U3497 (N_3497,N_2794,N_2258);
or U3498 (N_3498,N_2302,N_2422);
or U3499 (N_3499,N_2599,N_2909);
and U3500 (N_3500,N_2847,N_2990);
nand U3501 (N_3501,N_2266,N_2631);
nor U3502 (N_3502,N_2352,N_2860);
and U3503 (N_3503,N_2383,N_2935);
nor U3504 (N_3504,N_2370,N_2831);
xnor U3505 (N_3505,N_2417,N_2700);
xor U3506 (N_3506,N_2623,N_2456);
nand U3507 (N_3507,N_2310,N_2796);
nand U3508 (N_3508,N_2939,N_2710);
and U3509 (N_3509,N_2353,N_2855);
nand U3510 (N_3510,N_2695,N_2631);
xor U3511 (N_3511,N_2528,N_2974);
or U3512 (N_3512,N_2668,N_2972);
or U3513 (N_3513,N_2597,N_2312);
nor U3514 (N_3514,N_2891,N_2851);
or U3515 (N_3515,N_2396,N_2946);
nand U3516 (N_3516,N_2668,N_2625);
nor U3517 (N_3517,N_2402,N_2656);
or U3518 (N_3518,N_2724,N_2520);
nand U3519 (N_3519,N_2693,N_2310);
xnor U3520 (N_3520,N_2910,N_2622);
nand U3521 (N_3521,N_2916,N_2531);
or U3522 (N_3522,N_2447,N_2713);
or U3523 (N_3523,N_2367,N_2874);
nor U3524 (N_3524,N_2659,N_2439);
or U3525 (N_3525,N_2744,N_2706);
nor U3526 (N_3526,N_2866,N_2578);
nand U3527 (N_3527,N_2487,N_2746);
xor U3528 (N_3528,N_2402,N_2771);
xor U3529 (N_3529,N_2373,N_2539);
and U3530 (N_3530,N_2570,N_2819);
nor U3531 (N_3531,N_2320,N_2268);
nor U3532 (N_3532,N_2911,N_2694);
or U3533 (N_3533,N_2947,N_2541);
and U3534 (N_3534,N_2275,N_2782);
or U3535 (N_3535,N_2985,N_2797);
and U3536 (N_3536,N_2468,N_2949);
and U3537 (N_3537,N_2263,N_2554);
xor U3538 (N_3538,N_2868,N_2848);
and U3539 (N_3539,N_2991,N_2420);
and U3540 (N_3540,N_2695,N_2333);
and U3541 (N_3541,N_2578,N_2371);
and U3542 (N_3542,N_2811,N_2828);
nor U3543 (N_3543,N_2988,N_2853);
and U3544 (N_3544,N_2397,N_2301);
nand U3545 (N_3545,N_2278,N_2418);
and U3546 (N_3546,N_2262,N_2364);
nand U3547 (N_3547,N_2892,N_2521);
nand U3548 (N_3548,N_2441,N_2769);
or U3549 (N_3549,N_2273,N_2986);
nor U3550 (N_3550,N_2510,N_2404);
and U3551 (N_3551,N_2340,N_2298);
xor U3552 (N_3552,N_2677,N_2341);
nand U3553 (N_3553,N_2994,N_2292);
nand U3554 (N_3554,N_2578,N_2609);
and U3555 (N_3555,N_2849,N_2492);
xor U3556 (N_3556,N_2497,N_2333);
nand U3557 (N_3557,N_2539,N_2897);
or U3558 (N_3558,N_2440,N_2545);
and U3559 (N_3559,N_2536,N_2975);
and U3560 (N_3560,N_2979,N_2550);
or U3561 (N_3561,N_2530,N_2681);
or U3562 (N_3562,N_2882,N_2735);
nand U3563 (N_3563,N_2320,N_2636);
nor U3564 (N_3564,N_2819,N_2641);
or U3565 (N_3565,N_2594,N_2974);
and U3566 (N_3566,N_2804,N_2681);
xor U3567 (N_3567,N_2682,N_2845);
and U3568 (N_3568,N_2586,N_2253);
or U3569 (N_3569,N_2998,N_2489);
xor U3570 (N_3570,N_2835,N_2605);
nor U3571 (N_3571,N_2372,N_2256);
nor U3572 (N_3572,N_2861,N_2477);
or U3573 (N_3573,N_2361,N_2706);
or U3574 (N_3574,N_2294,N_2554);
and U3575 (N_3575,N_2316,N_2790);
and U3576 (N_3576,N_2921,N_2536);
or U3577 (N_3577,N_2927,N_2305);
and U3578 (N_3578,N_2957,N_2554);
nand U3579 (N_3579,N_2825,N_2393);
xnor U3580 (N_3580,N_2391,N_2714);
and U3581 (N_3581,N_2490,N_2878);
and U3582 (N_3582,N_2546,N_2370);
nand U3583 (N_3583,N_2252,N_2671);
xor U3584 (N_3584,N_2669,N_2980);
xnor U3585 (N_3585,N_2779,N_2687);
nor U3586 (N_3586,N_2748,N_2320);
or U3587 (N_3587,N_2598,N_2291);
and U3588 (N_3588,N_2963,N_2356);
nor U3589 (N_3589,N_2656,N_2917);
nand U3590 (N_3590,N_2403,N_2454);
nand U3591 (N_3591,N_2603,N_2283);
or U3592 (N_3592,N_2739,N_2789);
and U3593 (N_3593,N_2391,N_2690);
xor U3594 (N_3594,N_2888,N_2621);
nor U3595 (N_3595,N_2500,N_2712);
nand U3596 (N_3596,N_2957,N_2531);
and U3597 (N_3597,N_2818,N_2275);
and U3598 (N_3598,N_2462,N_2624);
xnor U3599 (N_3599,N_2693,N_2759);
nor U3600 (N_3600,N_2390,N_2994);
nor U3601 (N_3601,N_2819,N_2330);
nand U3602 (N_3602,N_2864,N_2292);
nor U3603 (N_3603,N_2827,N_2790);
nor U3604 (N_3604,N_2271,N_2610);
nor U3605 (N_3605,N_2422,N_2623);
and U3606 (N_3606,N_2456,N_2977);
nor U3607 (N_3607,N_2657,N_2887);
and U3608 (N_3608,N_2480,N_2651);
nand U3609 (N_3609,N_2791,N_2503);
nand U3610 (N_3610,N_2433,N_2692);
or U3611 (N_3611,N_2929,N_2748);
and U3612 (N_3612,N_2328,N_2831);
or U3613 (N_3613,N_2390,N_2440);
and U3614 (N_3614,N_2273,N_2500);
nor U3615 (N_3615,N_2895,N_2589);
or U3616 (N_3616,N_2272,N_2452);
nand U3617 (N_3617,N_2515,N_2961);
nor U3618 (N_3618,N_2653,N_2782);
nand U3619 (N_3619,N_2668,N_2936);
and U3620 (N_3620,N_2770,N_2805);
xnor U3621 (N_3621,N_2647,N_2294);
and U3622 (N_3622,N_2377,N_2872);
nor U3623 (N_3623,N_2971,N_2818);
nor U3624 (N_3624,N_2730,N_2986);
nand U3625 (N_3625,N_2686,N_2894);
or U3626 (N_3626,N_2650,N_2756);
or U3627 (N_3627,N_2488,N_2654);
nor U3628 (N_3628,N_2617,N_2525);
xnor U3629 (N_3629,N_2832,N_2433);
xor U3630 (N_3630,N_2516,N_2508);
or U3631 (N_3631,N_2395,N_2894);
or U3632 (N_3632,N_2498,N_2998);
nand U3633 (N_3633,N_2882,N_2964);
nor U3634 (N_3634,N_2338,N_2783);
and U3635 (N_3635,N_2264,N_2937);
nor U3636 (N_3636,N_2434,N_2251);
nand U3637 (N_3637,N_2802,N_2341);
nor U3638 (N_3638,N_2849,N_2581);
nand U3639 (N_3639,N_2584,N_2579);
nor U3640 (N_3640,N_2575,N_2822);
xnor U3641 (N_3641,N_2350,N_2964);
nor U3642 (N_3642,N_2381,N_2706);
nand U3643 (N_3643,N_2496,N_2441);
nand U3644 (N_3644,N_2763,N_2387);
or U3645 (N_3645,N_2878,N_2846);
or U3646 (N_3646,N_2584,N_2415);
or U3647 (N_3647,N_2986,N_2493);
and U3648 (N_3648,N_2969,N_2659);
nor U3649 (N_3649,N_2527,N_2882);
and U3650 (N_3650,N_2741,N_2512);
and U3651 (N_3651,N_2508,N_2260);
xor U3652 (N_3652,N_2782,N_2453);
or U3653 (N_3653,N_2271,N_2492);
xnor U3654 (N_3654,N_2841,N_2307);
or U3655 (N_3655,N_2804,N_2910);
and U3656 (N_3656,N_2563,N_2826);
and U3657 (N_3657,N_2601,N_2941);
nand U3658 (N_3658,N_2949,N_2771);
nand U3659 (N_3659,N_2786,N_2783);
and U3660 (N_3660,N_2567,N_2294);
nor U3661 (N_3661,N_2825,N_2998);
or U3662 (N_3662,N_2552,N_2715);
nor U3663 (N_3663,N_2483,N_2256);
xor U3664 (N_3664,N_2696,N_2423);
or U3665 (N_3665,N_2750,N_2993);
nor U3666 (N_3666,N_2918,N_2904);
or U3667 (N_3667,N_2930,N_2931);
and U3668 (N_3668,N_2730,N_2773);
nor U3669 (N_3669,N_2304,N_2823);
and U3670 (N_3670,N_2440,N_2345);
or U3671 (N_3671,N_2357,N_2610);
and U3672 (N_3672,N_2736,N_2799);
nand U3673 (N_3673,N_2550,N_2359);
and U3674 (N_3674,N_2349,N_2751);
nand U3675 (N_3675,N_2511,N_2979);
nand U3676 (N_3676,N_2565,N_2544);
and U3677 (N_3677,N_2996,N_2504);
xor U3678 (N_3678,N_2968,N_2280);
nand U3679 (N_3679,N_2969,N_2884);
or U3680 (N_3680,N_2950,N_2793);
nor U3681 (N_3681,N_2594,N_2775);
or U3682 (N_3682,N_2523,N_2851);
or U3683 (N_3683,N_2552,N_2795);
nand U3684 (N_3684,N_2317,N_2520);
nand U3685 (N_3685,N_2985,N_2277);
and U3686 (N_3686,N_2966,N_2510);
or U3687 (N_3687,N_2252,N_2595);
nand U3688 (N_3688,N_2433,N_2616);
nor U3689 (N_3689,N_2624,N_2475);
or U3690 (N_3690,N_2899,N_2838);
nand U3691 (N_3691,N_2678,N_2437);
and U3692 (N_3692,N_2329,N_2429);
nand U3693 (N_3693,N_2760,N_2975);
nor U3694 (N_3694,N_2843,N_2659);
and U3695 (N_3695,N_2359,N_2619);
or U3696 (N_3696,N_2890,N_2565);
or U3697 (N_3697,N_2382,N_2273);
nor U3698 (N_3698,N_2937,N_2759);
and U3699 (N_3699,N_2793,N_2305);
nor U3700 (N_3700,N_2888,N_2880);
and U3701 (N_3701,N_2956,N_2448);
and U3702 (N_3702,N_2305,N_2567);
and U3703 (N_3703,N_2884,N_2888);
xor U3704 (N_3704,N_2624,N_2391);
or U3705 (N_3705,N_2356,N_2700);
or U3706 (N_3706,N_2434,N_2809);
nor U3707 (N_3707,N_2691,N_2793);
and U3708 (N_3708,N_2511,N_2332);
nor U3709 (N_3709,N_2410,N_2765);
or U3710 (N_3710,N_2546,N_2523);
and U3711 (N_3711,N_2851,N_2423);
and U3712 (N_3712,N_2651,N_2440);
nand U3713 (N_3713,N_2932,N_2689);
or U3714 (N_3714,N_2378,N_2400);
nand U3715 (N_3715,N_2266,N_2427);
nand U3716 (N_3716,N_2981,N_2849);
or U3717 (N_3717,N_2482,N_2963);
or U3718 (N_3718,N_2555,N_2621);
and U3719 (N_3719,N_2561,N_2809);
nand U3720 (N_3720,N_2766,N_2447);
nand U3721 (N_3721,N_2881,N_2492);
xor U3722 (N_3722,N_2853,N_2608);
and U3723 (N_3723,N_2516,N_2997);
nor U3724 (N_3724,N_2898,N_2770);
nor U3725 (N_3725,N_2652,N_2709);
or U3726 (N_3726,N_2838,N_2971);
nand U3727 (N_3727,N_2379,N_2464);
nor U3728 (N_3728,N_2761,N_2338);
nor U3729 (N_3729,N_2956,N_2351);
nand U3730 (N_3730,N_2662,N_2976);
and U3731 (N_3731,N_2997,N_2305);
and U3732 (N_3732,N_2357,N_2288);
and U3733 (N_3733,N_2433,N_2867);
nand U3734 (N_3734,N_2830,N_2841);
and U3735 (N_3735,N_2925,N_2978);
or U3736 (N_3736,N_2922,N_2796);
nand U3737 (N_3737,N_2916,N_2501);
nand U3738 (N_3738,N_2579,N_2453);
nand U3739 (N_3739,N_2859,N_2306);
nand U3740 (N_3740,N_2802,N_2579);
or U3741 (N_3741,N_2915,N_2527);
or U3742 (N_3742,N_2678,N_2369);
nand U3743 (N_3743,N_2292,N_2974);
or U3744 (N_3744,N_2442,N_2731);
nand U3745 (N_3745,N_2602,N_2729);
and U3746 (N_3746,N_2283,N_2922);
or U3747 (N_3747,N_2371,N_2476);
or U3748 (N_3748,N_2569,N_2301);
nor U3749 (N_3749,N_2767,N_2343);
nor U3750 (N_3750,N_3438,N_3598);
and U3751 (N_3751,N_3114,N_3188);
or U3752 (N_3752,N_3467,N_3148);
or U3753 (N_3753,N_3245,N_3400);
and U3754 (N_3754,N_3265,N_3544);
nand U3755 (N_3755,N_3257,N_3374);
xnor U3756 (N_3756,N_3299,N_3701);
or U3757 (N_3757,N_3558,N_3127);
or U3758 (N_3758,N_3517,N_3235);
or U3759 (N_3759,N_3232,N_3738);
nor U3760 (N_3760,N_3206,N_3056);
nand U3761 (N_3761,N_3640,N_3332);
nor U3762 (N_3762,N_3227,N_3673);
nor U3763 (N_3763,N_3748,N_3717);
nand U3764 (N_3764,N_3100,N_3158);
or U3765 (N_3765,N_3182,N_3381);
or U3766 (N_3766,N_3122,N_3401);
and U3767 (N_3767,N_3493,N_3347);
and U3768 (N_3768,N_3111,N_3157);
and U3769 (N_3769,N_3631,N_3274);
and U3770 (N_3770,N_3041,N_3471);
or U3771 (N_3771,N_3339,N_3358);
and U3772 (N_3772,N_3003,N_3051);
and U3773 (N_3773,N_3349,N_3448);
nor U3774 (N_3774,N_3585,N_3474);
xnor U3775 (N_3775,N_3125,N_3675);
and U3776 (N_3776,N_3676,N_3175);
nand U3777 (N_3777,N_3123,N_3000);
nor U3778 (N_3778,N_3340,N_3120);
nor U3779 (N_3779,N_3407,N_3033);
or U3780 (N_3780,N_3511,N_3117);
or U3781 (N_3781,N_3069,N_3691);
and U3782 (N_3782,N_3255,N_3537);
and U3783 (N_3783,N_3472,N_3485);
or U3784 (N_3784,N_3654,N_3508);
nor U3785 (N_3785,N_3398,N_3744);
and U3786 (N_3786,N_3626,N_3115);
nand U3787 (N_3787,N_3080,N_3151);
xnor U3788 (N_3788,N_3382,N_3217);
nor U3789 (N_3789,N_3361,N_3663);
nor U3790 (N_3790,N_3499,N_3124);
nor U3791 (N_3791,N_3700,N_3501);
or U3792 (N_3792,N_3276,N_3666);
and U3793 (N_3793,N_3498,N_3481);
or U3794 (N_3794,N_3713,N_3062);
or U3795 (N_3795,N_3319,N_3475);
nor U3796 (N_3796,N_3538,N_3521);
xor U3797 (N_3797,N_3327,N_3311);
or U3798 (N_3798,N_3615,N_3518);
nor U3799 (N_3799,N_3006,N_3684);
and U3800 (N_3800,N_3431,N_3489);
nor U3801 (N_3801,N_3196,N_3366);
or U3802 (N_3802,N_3015,N_3238);
nor U3803 (N_3803,N_3243,N_3293);
nand U3804 (N_3804,N_3163,N_3030);
or U3805 (N_3805,N_3420,N_3424);
nor U3806 (N_3806,N_3283,N_3466);
nor U3807 (N_3807,N_3270,N_3009);
nor U3808 (N_3808,N_3688,N_3669);
and U3809 (N_3809,N_3025,N_3614);
or U3810 (N_3810,N_3742,N_3433);
xnor U3811 (N_3811,N_3601,N_3556);
nand U3812 (N_3812,N_3596,N_3272);
nand U3813 (N_3813,N_3342,N_3568);
nand U3814 (N_3814,N_3533,N_3636);
or U3815 (N_3815,N_3098,N_3239);
or U3816 (N_3816,N_3309,N_3279);
or U3817 (N_3817,N_3152,N_3018);
or U3818 (N_3818,N_3099,N_3021);
nand U3819 (N_3819,N_3324,N_3728);
nor U3820 (N_3820,N_3269,N_3638);
nor U3821 (N_3821,N_3065,N_3328);
or U3822 (N_3822,N_3144,N_3121);
nand U3823 (N_3823,N_3330,N_3579);
nor U3824 (N_3824,N_3621,N_3622);
nor U3825 (N_3825,N_3256,N_3671);
nor U3826 (N_3826,N_3735,N_3116);
and U3827 (N_3827,N_3209,N_3378);
and U3828 (N_3828,N_3672,N_3668);
xor U3829 (N_3829,N_3600,N_3402);
nor U3830 (N_3830,N_3641,N_3444);
or U3831 (N_3831,N_3428,N_3457);
nand U3832 (N_3832,N_3250,N_3179);
nor U3833 (N_3833,N_3388,N_3126);
nor U3834 (N_3834,N_3734,N_3649);
nand U3835 (N_3835,N_3618,N_3722);
nor U3836 (N_3836,N_3743,N_3530);
and U3837 (N_3837,N_3494,N_3060);
nand U3838 (N_3838,N_3220,N_3718);
or U3839 (N_3839,N_3632,N_3681);
nor U3840 (N_3840,N_3200,N_3139);
and U3841 (N_3841,N_3561,N_3307);
or U3842 (N_3842,N_3159,N_3244);
nor U3843 (N_3843,N_3298,N_3635);
xnor U3844 (N_3844,N_3383,N_3067);
or U3845 (N_3845,N_3746,N_3507);
or U3846 (N_3846,N_3189,N_3606);
nor U3847 (N_3847,N_3091,N_3130);
nor U3848 (N_3848,N_3287,N_3429);
xnor U3849 (N_3849,N_3054,N_3617);
nand U3850 (N_3850,N_3716,N_3252);
or U3851 (N_3851,N_3173,N_3459);
nand U3852 (N_3852,N_3704,N_3500);
nand U3853 (N_3853,N_3384,N_3164);
nand U3854 (N_3854,N_3645,N_3451);
and U3855 (N_3855,N_3741,N_3480);
or U3856 (N_3856,N_3247,N_3028);
nand U3857 (N_3857,N_3277,N_3723);
or U3858 (N_3858,N_3204,N_3412);
and U3859 (N_3859,N_3532,N_3588);
or U3860 (N_3860,N_3246,N_3107);
nand U3861 (N_3861,N_3195,N_3369);
or U3862 (N_3862,N_3035,N_3686);
and U3863 (N_3863,N_3652,N_3039);
xor U3864 (N_3864,N_3304,N_3219);
xor U3865 (N_3865,N_3371,N_3657);
nor U3866 (N_3866,N_3233,N_3578);
nand U3867 (N_3867,N_3357,N_3540);
nand U3868 (N_3868,N_3291,N_3013);
nand U3869 (N_3869,N_3613,N_3551);
nand U3870 (N_3870,N_3553,N_3446);
xor U3871 (N_3871,N_3418,N_3720);
nor U3872 (N_3872,N_3002,N_3300);
or U3873 (N_3873,N_3329,N_3104);
nor U3874 (N_3874,N_3354,N_3180);
or U3875 (N_3875,N_3226,N_3083);
or U3876 (N_3876,N_3222,N_3043);
nor U3877 (N_3877,N_3515,N_3207);
nand U3878 (N_3878,N_3172,N_3519);
xnor U3879 (N_3879,N_3674,N_3655);
and U3880 (N_3880,N_3040,N_3468);
or U3881 (N_3881,N_3086,N_3085);
or U3882 (N_3882,N_3557,N_3203);
nor U3883 (N_3883,N_3084,N_3461);
nand U3884 (N_3884,N_3453,N_3186);
or U3885 (N_3885,N_3310,N_3387);
nand U3886 (N_3886,N_3590,N_3516);
and U3887 (N_3887,N_3278,N_3047);
and U3888 (N_3888,N_3731,N_3647);
nor U3889 (N_3889,N_3736,N_3706);
or U3890 (N_3890,N_3667,N_3425);
and U3891 (N_3891,N_3503,N_3696);
nand U3892 (N_3892,N_3237,N_3592);
or U3893 (N_3893,N_3112,N_3583);
nor U3894 (N_3894,N_3405,N_3464);
nand U3895 (N_3895,N_3137,N_3413);
nand U3896 (N_3896,N_3423,N_3092);
and U3897 (N_3897,N_3184,N_3094);
or U3898 (N_3898,N_3619,N_3694);
nor U3899 (N_3899,N_3665,N_3303);
nor U3900 (N_3900,N_3271,N_3629);
nor U3901 (N_3901,N_3611,N_3462);
and U3902 (N_3902,N_3333,N_3174);
nor U3903 (N_3903,N_3660,N_3465);
or U3904 (N_3904,N_3078,N_3531);
nand U3905 (N_3905,N_3076,N_3221);
nand U3906 (N_3906,N_3261,N_3662);
or U3907 (N_3907,N_3698,N_3230);
and U3908 (N_3908,N_3612,N_3029);
nor U3909 (N_3909,N_3389,N_3241);
or U3910 (N_3910,N_3609,N_3460);
nand U3911 (N_3911,N_3156,N_3452);
or U3912 (N_3912,N_3703,N_3058);
nor U3913 (N_3913,N_3089,N_3725);
and U3914 (N_3914,N_3208,N_3143);
and U3915 (N_3915,N_3059,N_3005);
nor U3916 (N_3916,N_3042,N_3314);
nand U3917 (N_3917,N_3229,N_3570);
nand U3918 (N_3918,N_3527,N_3749);
nor U3919 (N_3919,N_3607,N_3105);
nor U3920 (N_3920,N_3334,N_3093);
nor U3921 (N_3921,N_3740,N_3392);
or U3922 (N_3922,N_3012,N_3138);
nand U3923 (N_3923,N_3224,N_3305);
nor U3924 (N_3924,N_3032,N_3267);
nor U3925 (N_3925,N_3348,N_3170);
and U3926 (N_3926,N_3068,N_3693);
nand U3927 (N_3927,N_3399,N_3658);
or U3928 (N_3928,N_3439,N_3166);
and U3929 (N_3929,N_3323,N_3386);
and U3930 (N_3930,N_3677,N_3132);
or U3931 (N_3931,N_3604,N_3571);
nor U3932 (N_3932,N_3223,N_3726);
nand U3933 (N_3933,N_3633,N_3258);
nand U3934 (N_3934,N_3251,N_3705);
nor U3935 (N_3935,N_3338,N_3010);
nor U3936 (N_3936,N_3211,N_3729);
xor U3937 (N_3937,N_3721,N_3397);
nand U3938 (N_3938,N_3316,N_3072);
nor U3939 (N_3939,N_3712,N_3739);
xnor U3940 (N_3940,N_3280,N_3315);
and U3941 (N_3941,N_3441,N_3052);
nor U3942 (N_3942,N_3595,N_3391);
nor U3943 (N_3943,N_3212,N_3552);
and U3944 (N_3944,N_3525,N_3414);
nor U3945 (N_3945,N_3496,N_3482);
or U3946 (N_3946,N_3470,N_3373);
or U3947 (N_3947,N_3565,N_3699);
and U3948 (N_3948,N_3682,N_3101);
or U3949 (N_3949,N_3345,N_3313);
nor U3950 (N_3950,N_3536,N_3341);
or U3951 (N_3951,N_3259,N_3526);
nand U3952 (N_3952,N_3097,N_3591);
xor U3953 (N_3953,N_3231,N_3082);
and U3954 (N_3954,N_3434,N_3487);
nand U3955 (N_3955,N_3048,N_3432);
or U3956 (N_3956,N_3061,N_3199);
and U3957 (N_3957,N_3071,N_3484);
nor U3958 (N_3958,N_3119,N_3106);
nand U3959 (N_3959,N_3075,N_3447);
or U3960 (N_3960,N_3034,N_3559);
or U3961 (N_3961,N_3201,N_3608);
nand U3962 (N_3962,N_3630,N_3282);
nor U3963 (N_3963,N_3073,N_3449);
nor U3964 (N_3964,N_3213,N_3528);
and U3965 (N_3965,N_3050,N_3288);
nand U3966 (N_3966,N_3587,N_3134);
or U3967 (N_3967,N_3478,N_3090);
and U3968 (N_3968,N_3594,N_3602);
or U3969 (N_3969,N_3053,N_3197);
and U3970 (N_3970,N_3648,N_3437);
nand U3971 (N_3971,N_3483,N_3422);
and U3972 (N_3972,N_3236,N_3194);
and U3973 (N_3973,N_3351,N_3308);
and U3974 (N_3974,N_3379,N_3008);
nand U3975 (N_3975,N_3367,N_3644);
or U3976 (N_3976,N_3455,N_3190);
nand U3977 (N_3977,N_3262,N_3365);
or U3978 (N_3978,N_3593,N_3435);
nand U3979 (N_3979,N_3142,N_3491);
nand U3980 (N_3980,N_3171,N_3046);
or U3981 (N_3981,N_3337,N_3504);
nor U3982 (N_3982,N_3456,N_3192);
nor U3983 (N_3983,N_3469,N_3589);
xor U3984 (N_3984,N_3599,N_3294);
nor U3985 (N_3985,N_3113,N_3577);
or U3986 (N_3986,N_3024,N_3572);
or U3987 (N_3987,N_3044,N_3545);
nand U3988 (N_3988,N_3178,N_3234);
nor U3989 (N_3989,N_3352,N_3637);
and U3990 (N_3990,N_3268,N_3031);
or U3991 (N_3991,N_3359,N_3249);
or U3992 (N_3992,N_3240,N_3715);
nand U3993 (N_3993,N_3548,N_3266);
xnor U3994 (N_3994,N_3620,N_3616);
or U3995 (N_3995,N_3543,N_3576);
nor U3996 (N_3996,N_3318,N_3542);
or U3997 (N_3997,N_3653,N_3580);
or U3998 (N_3998,N_3146,N_3473);
and U3999 (N_3999,N_3479,N_3403);
nor U4000 (N_4000,N_3218,N_3356);
and U4001 (N_4001,N_3719,N_3198);
or U4002 (N_4002,N_3575,N_3514);
xor U4003 (N_4003,N_3045,N_3443);
nand U4004 (N_4004,N_3295,N_3177);
and U4005 (N_4005,N_3642,N_3529);
nand U4006 (N_4006,N_3087,N_3074);
nand U4007 (N_4007,N_3605,N_3225);
nor U4008 (N_4008,N_3560,N_3037);
and U4009 (N_4009,N_3363,N_3296);
xor U4010 (N_4010,N_3128,N_3393);
xnor U4011 (N_4011,N_3183,N_3541);
and U4012 (N_4012,N_3440,N_3070);
and U4013 (N_4013,N_3664,N_3331);
nand U4014 (N_4014,N_3522,N_3375);
nor U4015 (N_4015,N_3185,N_3297);
or U4016 (N_4016,N_3108,N_3205);
xnor U4017 (N_4017,N_3490,N_3697);
or U4018 (N_4018,N_3510,N_3004);
xnor U4019 (N_4019,N_3563,N_3584);
and U4020 (N_4020,N_3216,N_3289);
xor U4021 (N_4021,N_3714,N_3057);
and U4022 (N_4022,N_3546,N_3110);
xnor U4023 (N_4023,N_3215,N_3547);
nor U4024 (N_4024,N_3370,N_3505);
nor U4025 (N_4025,N_3509,N_3372);
or U4026 (N_4026,N_3165,N_3396);
or U4027 (N_4027,N_3680,N_3394);
nor U4028 (N_4028,N_3495,N_3564);
and U4029 (N_4029,N_3670,N_3646);
nor U4030 (N_4030,N_3079,N_3709);
nand U4031 (N_4031,N_3155,N_3254);
nand U4032 (N_4032,N_3659,N_3077);
and U4033 (N_4033,N_3695,N_3285);
and U4034 (N_4034,N_3610,N_3325);
xor U4035 (N_4035,N_3454,N_3368);
xnor U4036 (N_4036,N_3477,N_3430);
or U4037 (N_4037,N_3566,N_3118);
xor U4038 (N_4038,N_3150,N_3678);
and U4039 (N_4039,N_3095,N_3707);
xor U4040 (N_4040,N_3063,N_3160);
or U4041 (N_4041,N_3539,N_3355);
or U4042 (N_4042,N_3103,N_3362);
nor U4043 (N_4043,N_3214,N_3248);
nor U4044 (N_4044,N_3162,N_3747);
and U4045 (N_4045,N_3275,N_3395);
or U4046 (N_4046,N_3281,N_3016);
nor U4047 (N_4047,N_3286,N_3421);
nand U4048 (N_4048,N_3569,N_3623);
nand U4049 (N_4049,N_3711,N_3426);
or U4050 (N_4050,N_3458,N_3129);
and U4051 (N_4051,N_3167,N_3102);
and U4052 (N_4052,N_3140,N_3520);
nor U4053 (N_4053,N_3136,N_3161);
or U4054 (N_4054,N_3055,N_3502);
nand U4055 (N_4055,N_3679,N_3476);
or U4056 (N_4056,N_3022,N_3168);
and U4057 (N_4057,N_3036,N_3326);
nand U4058 (N_4058,N_3650,N_3390);
and U4059 (N_4059,N_3683,N_3169);
or U4060 (N_4060,N_3141,N_3581);
or U4061 (N_4061,N_3450,N_3643);
nand U4062 (N_4062,N_3336,N_3523);
nand U4063 (N_4063,N_3317,N_3512);
and U4064 (N_4064,N_3692,N_3135);
nor U4065 (N_4065,N_3154,N_3625);
and U4066 (N_4066,N_3210,N_3639);
nor U4067 (N_4067,N_3263,N_3320);
and U4068 (N_4068,N_3550,N_3346);
xor U4069 (N_4069,N_3627,N_3687);
and U4070 (N_4070,N_3685,N_3409);
or U4071 (N_4071,N_3582,N_3586);
nor U4072 (N_4072,N_3385,N_3377);
nand U4073 (N_4073,N_3153,N_3436);
and U4074 (N_4074,N_3109,N_3181);
nand U4075 (N_4075,N_3322,N_3253);
nor U4076 (N_4076,N_3360,N_3284);
and U4077 (N_4077,N_3689,N_3064);
nand U4078 (N_4078,N_3191,N_3007);
or U4079 (N_4079,N_3406,N_3131);
nor U4080 (N_4080,N_3023,N_3096);
xnor U4081 (N_4081,N_3497,N_3260);
nand U4082 (N_4082,N_3488,N_3081);
and U4083 (N_4083,N_3302,N_3442);
or U4084 (N_4084,N_3187,N_3702);
or U4085 (N_4085,N_3014,N_3149);
xor U4086 (N_4086,N_3486,N_3321);
and U4087 (N_4087,N_3710,N_3535);
nor U4088 (N_4088,N_3343,N_3376);
nand U4089 (N_4089,N_3634,N_3410);
nor U4090 (N_4090,N_3088,N_3353);
nor U4091 (N_4091,N_3651,N_3417);
nand U4092 (N_4092,N_3408,N_3427);
nor U4093 (N_4093,N_3554,N_3573);
nand U4094 (N_4094,N_3027,N_3020);
nor U4095 (N_4095,N_3290,N_3524);
nand U4096 (N_4096,N_3549,N_3292);
nand U4097 (N_4097,N_3555,N_3350);
nand U4098 (N_4098,N_3737,N_3597);
and U4099 (N_4099,N_3411,N_3574);
and U4100 (N_4100,N_3492,N_3306);
nand U4101 (N_4101,N_3017,N_3176);
nand U4102 (N_4102,N_3415,N_3628);
or U4103 (N_4103,N_3732,N_3445);
and U4104 (N_4104,N_3011,N_3242);
or U4105 (N_4105,N_3567,N_3724);
xor U4106 (N_4106,N_3416,N_3133);
nor U4107 (N_4107,N_3335,N_3049);
or U4108 (N_4108,N_3228,N_3603);
nor U4109 (N_4109,N_3202,N_3730);
or U4110 (N_4110,N_3301,N_3419);
nor U4111 (N_4111,N_3404,N_3463);
nor U4112 (N_4112,N_3312,N_3364);
nand U4113 (N_4113,N_3193,N_3624);
nor U4114 (N_4114,N_3066,N_3344);
xor U4115 (N_4115,N_3727,N_3145);
nor U4116 (N_4116,N_3733,N_3745);
nand U4117 (N_4117,N_3661,N_3026);
nand U4118 (N_4118,N_3038,N_3019);
and U4119 (N_4119,N_3562,N_3147);
and U4120 (N_4120,N_3690,N_3708);
and U4121 (N_4121,N_3264,N_3273);
nor U4122 (N_4122,N_3380,N_3506);
nor U4123 (N_4123,N_3656,N_3001);
nor U4124 (N_4124,N_3534,N_3513);
nor U4125 (N_4125,N_3281,N_3514);
and U4126 (N_4126,N_3394,N_3589);
xor U4127 (N_4127,N_3603,N_3626);
nand U4128 (N_4128,N_3685,N_3222);
or U4129 (N_4129,N_3377,N_3252);
or U4130 (N_4130,N_3674,N_3261);
nor U4131 (N_4131,N_3508,N_3385);
nor U4132 (N_4132,N_3240,N_3008);
nand U4133 (N_4133,N_3516,N_3465);
and U4134 (N_4134,N_3149,N_3225);
nor U4135 (N_4135,N_3450,N_3330);
nor U4136 (N_4136,N_3685,N_3547);
nor U4137 (N_4137,N_3150,N_3366);
nand U4138 (N_4138,N_3294,N_3649);
nand U4139 (N_4139,N_3021,N_3512);
and U4140 (N_4140,N_3474,N_3475);
and U4141 (N_4141,N_3290,N_3091);
nor U4142 (N_4142,N_3728,N_3057);
and U4143 (N_4143,N_3693,N_3116);
nand U4144 (N_4144,N_3307,N_3550);
nand U4145 (N_4145,N_3098,N_3003);
and U4146 (N_4146,N_3607,N_3534);
or U4147 (N_4147,N_3494,N_3707);
and U4148 (N_4148,N_3068,N_3085);
nor U4149 (N_4149,N_3644,N_3035);
nor U4150 (N_4150,N_3563,N_3327);
nor U4151 (N_4151,N_3385,N_3574);
or U4152 (N_4152,N_3200,N_3637);
and U4153 (N_4153,N_3005,N_3748);
and U4154 (N_4154,N_3552,N_3508);
and U4155 (N_4155,N_3085,N_3184);
xor U4156 (N_4156,N_3303,N_3649);
or U4157 (N_4157,N_3052,N_3020);
or U4158 (N_4158,N_3331,N_3305);
nor U4159 (N_4159,N_3050,N_3739);
nor U4160 (N_4160,N_3458,N_3288);
nor U4161 (N_4161,N_3402,N_3450);
or U4162 (N_4162,N_3359,N_3267);
nand U4163 (N_4163,N_3440,N_3414);
nor U4164 (N_4164,N_3691,N_3461);
nand U4165 (N_4165,N_3147,N_3341);
and U4166 (N_4166,N_3137,N_3363);
and U4167 (N_4167,N_3605,N_3402);
nand U4168 (N_4168,N_3097,N_3064);
and U4169 (N_4169,N_3414,N_3054);
nand U4170 (N_4170,N_3502,N_3254);
nand U4171 (N_4171,N_3372,N_3610);
and U4172 (N_4172,N_3706,N_3556);
nor U4173 (N_4173,N_3185,N_3542);
or U4174 (N_4174,N_3693,N_3010);
nand U4175 (N_4175,N_3149,N_3306);
nor U4176 (N_4176,N_3291,N_3246);
nand U4177 (N_4177,N_3109,N_3539);
or U4178 (N_4178,N_3590,N_3196);
or U4179 (N_4179,N_3469,N_3426);
nor U4180 (N_4180,N_3043,N_3629);
nand U4181 (N_4181,N_3231,N_3583);
and U4182 (N_4182,N_3424,N_3674);
nand U4183 (N_4183,N_3364,N_3640);
nor U4184 (N_4184,N_3012,N_3528);
or U4185 (N_4185,N_3031,N_3359);
or U4186 (N_4186,N_3228,N_3243);
or U4187 (N_4187,N_3547,N_3213);
and U4188 (N_4188,N_3688,N_3034);
xnor U4189 (N_4189,N_3422,N_3366);
nor U4190 (N_4190,N_3120,N_3513);
or U4191 (N_4191,N_3036,N_3494);
or U4192 (N_4192,N_3498,N_3596);
nor U4193 (N_4193,N_3687,N_3464);
nor U4194 (N_4194,N_3412,N_3541);
nor U4195 (N_4195,N_3639,N_3066);
or U4196 (N_4196,N_3502,N_3217);
nand U4197 (N_4197,N_3419,N_3201);
nor U4198 (N_4198,N_3682,N_3040);
nand U4199 (N_4199,N_3198,N_3180);
and U4200 (N_4200,N_3735,N_3547);
or U4201 (N_4201,N_3342,N_3182);
nor U4202 (N_4202,N_3098,N_3362);
nor U4203 (N_4203,N_3400,N_3262);
nand U4204 (N_4204,N_3097,N_3243);
or U4205 (N_4205,N_3278,N_3034);
nor U4206 (N_4206,N_3250,N_3621);
nand U4207 (N_4207,N_3630,N_3409);
nand U4208 (N_4208,N_3496,N_3376);
and U4209 (N_4209,N_3316,N_3055);
nor U4210 (N_4210,N_3092,N_3070);
or U4211 (N_4211,N_3130,N_3032);
and U4212 (N_4212,N_3237,N_3571);
nor U4213 (N_4213,N_3282,N_3413);
and U4214 (N_4214,N_3737,N_3005);
nor U4215 (N_4215,N_3554,N_3480);
nand U4216 (N_4216,N_3117,N_3587);
nand U4217 (N_4217,N_3529,N_3414);
nand U4218 (N_4218,N_3170,N_3033);
nor U4219 (N_4219,N_3411,N_3036);
xor U4220 (N_4220,N_3493,N_3559);
nand U4221 (N_4221,N_3510,N_3544);
nand U4222 (N_4222,N_3320,N_3211);
nor U4223 (N_4223,N_3741,N_3552);
nand U4224 (N_4224,N_3470,N_3107);
xnor U4225 (N_4225,N_3313,N_3460);
nand U4226 (N_4226,N_3746,N_3728);
nand U4227 (N_4227,N_3398,N_3017);
or U4228 (N_4228,N_3385,N_3032);
and U4229 (N_4229,N_3280,N_3427);
nand U4230 (N_4230,N_3618,N_3027);
nor U4231 (N_4231,N_3421,N_3236);
nor U4232 (N_4232,N_3613,N_3454);
xor U4233 (N_4233,N_3192,N_3601);
nand U4234 (N_4234,N_3116,N_3076);
or U4235 (N_4235,N_3018,N_3441);
and U4236 (N_4236,N_3176,N_3512);
nor U4237 (N_4237,N_3415,N_3486);
or U4238 (N_4238,N_3443,N_3308);
and U4239 (N_4239,N_3523,N_3512);
nand U4240 (N_4240,N_3287,N_3175);
or U4241 (N_4241,N_3258,N_3689);
or U4242 (N_4242,N_3186,N_3343);
and U4243 (N_4243,N_3677,N_3673);
nand U4244 (N_4244,N_3153,N_3483);
or U4245 (N_4245,N_3188,N_3546);
nand U4246 (N_4246,N_3447,N_3503);
nand U4247 (N_4247,N_3349,N_3290);
and U4248 (N_4248,N_3519,N_3688);
nor U4249 (N_4249,N_3079,N_3517);
and U4250 (N_4250,N_3200,N_3075);
nand U4251 (N_4251,N_3640,N_3005);
or U4252 (N_4252,N_3116,N_3212);
nor U4253 (N_4253,N_3679,N_3576);
xnor U4254 (N_4254,N_3479,N_3284);
nor U4255 (N_4255,N_3474,N_3021);
nand U4256 (N_4256,N_3374,N_3377);
nor U4257 (N_4257,N_3593,N_3135);
and U4258 (N_4258,N_3605,N_3115);
and U4259 (N_4259,N_3017,N_3518);
or U4260 (N_4260,N_3622,N_3037);
nand U4261 (N_4261,N_3391,N_3375);
or U4262 (N_4262,N_3477,N_3647);
and U4263 (N_4263,N_3247,N_3727);
xnor U4264 (N_4264,N_3643,N_3501);
and U4265 (N_4265,N_3687,N_3209);
nor U4266 (N_4266,N_3242,N_3643);
and U4267 (N_4267,N_3493,N_3520);
nand U4268 (N_4268,N_3038,N_3429);
nand U4269 (N_4269,N_3672,N_3351);
and U4270 (N_4270,N_3748,N_3460);
and U4271 (N_4271,N_3582,N_3511);
nand U4272 (N_4272,N_3009,N_3106);
or U4273 (N_4273,N_3374,N_3201);
nor U4274 (N_4274,N_3009,N_3199);
or U4275 (N_4275,N_3572,N_3090);
xor U4276 (N_4276,N_3580,N_3684);
and U4277 (N_4277,N_3600,N_3470);
or U4278 (N_4278,N_3681,N_3389);
and U4279 (N_4279,N_3460,N_3560);
nand U4280 (N_4280,N_3280,N_3317);
or U4281 (N_4281,N_3009,N_3300);
or U4282 (N_4282,N_3432,N_3308);
nand U4283 (N_4283,N_3304,N_3681);
nor U4284 (N_4284,N_3249,N_3440);
nor U4285 (N_4285,N_3638,N_3557);
nand U4286 (N_4286,N_3222,N_3354);
and U4287 (N_4287,N_3345,N_3398);
and U4288 (N_4288,N_3273,N_3476);
and U4289 (N_4289,N_3743,N_3662);
nor U4290 (N_4290,N_3035,N_3373);
and U4291 (N_4291,N_3266,N_3667);
nand U4292 (N_4292,N_3696,N_3071);
nor U4293 (N_4293,N_3451,N_3295);
nor U4294 (N_4294,N_3667,N_3017);
or U4295 (N_4295,N_3613,N_3306);
or U4296 (N_4296,N_3453,N_3391);
and U4297 (N_4297,N_3678,N_3673);
nor U4298 (N_4298,N_3039,N_3710);
nand U4299 (N_4299,N_3359,N_3195);
and U4300 (N_4300,N_3664,N_3366);
nor U4301 (N_4301,N_3704,N_3553);
nor U4302 (N_4302,N_3497,N_3044);
xor U4303 (N_4303,N_3224,N_3265);
and U4304 (N_4304,N_3123,N_3032);
or U4305 (N_4305,N_3302,N_3635);
or U4306 (N_4306,N_3626,N_3204);
nor U4307 (N_4307,N_3003,N_3250);
and U4308 (N_4308,N_3618,N_3007);
nor U4309 (N_4309,N_3518,N_3551);
and U4310 (N_4310,N_3006,N_3594);
and U4311 (N_4311,N_3610,N_3518);
and U4312 (N_4312,N_3229,N_3267);
nor U4313 (N_4313,N_3004,N_3435);
and U4314 (N_4314,N_3160,N_3245);
or U4315 (N_4315,N_3589,N_3324);
or U4316 (N_4316,N_3047,N_3079);
nand U4317 (N_4317,N_3299,N_3630);
and U4318 (N_4318,N_3401,N_3546);
or U4319 (N_4319,N_3068,N_3580);
nand U4320 (N_4320,N_3039,N_3318);
or U4321 (N_4321,N_3357,N_3031);
nor U4322 (N_4322,N_3662,N_3046);
or U4323 (N_4323,N_3135,N_3577);
nor U4324 (N_4324,N_3708,N_3299);
and U4325 (N_4325,N_3533,N_3482);
and U4326 (N_4326,N_3287,N_3668);
or U4327 (N_4327,N_3485,N_3717);
and U4328 (N_4328,N_3186,N_3251);
xor U4329 (N_4329,N_3488,N_3012);
nand U4330 (N_4330,N_3041,N_3331);
nor U4331 (N_4331,N_3146,N_3274);
nand U4332 (N_4332,N_3611,N_3440);
or U4333 (N_4333,N_3446,N_3020);
nor U4334 (N_4334,N_3018,N_3256);
nor U4335 (N_4335,N_3524,N_3002);
and U4336 (N_4336,N_3725,N_3457);
xor U4337 (N_4337,N_3484,N_3268);
nor U4338 (N_4338,N_3407,N_3373);
and U4339 (N_4339,N_3079,N_3350);
xor U4340 (N_4340,N_3192,N_3271);
and U4341 (N_4341,N_3063,N_3552);
nand U4342 (N_4342,N_3316,N_3503);
nand U4343 (N_4343,N_3707,N_3659);
nor U4344 (N_4344,N_3087,N_3423);
and U4345 (N_4345,N_3354,N_3445);
nand U4346 (N_4346,N_3028,N_3588);
xnor U4347 (N_4347,N_3129,N_3041);
and U4348 (N_4348,N_3737,N_3114);
and U4349 (N_4349,N_3168,N_3586);
or U4350 (N_4350,N_3233,N_3241);
nor U4351 (N_4351,N_3480,N_3072);
nand U4352 (N_4352,N_3534,N_3526);
nor U4353 (N_4353,N_3236,N_3630);
nor U4354 (N_4354,N_3654,N_3258);
nand U4355 (N_4355,N_3462,N_3425);
nand U4356 (N_4356,N_3465,N_3035);
nor U4357 (N_4357,N_3064,N_3377);
nor U4358 (N_4358,N_3266,N_3287);
and U4359 (N_4359,N_3246,N_3364);
and U4360 (N_4360,N_3637,N_3411);
nor U4361 (N_4361,N_3223,N_3113);
or U4362 (N_4362,N_3569,N_3083);
and U4363 (N_4363,N_3720,N_3056);
nor U4364 (N_4364,N_3459,N_3067);
nand U4365 (N_4365,N_3311,N_3354);
and U4366 (N_4366,N_3546,N_3107);
nand U4367 (N_4367,N_3735,N_3132);
and U4368 (N_4368,N_3042,N_3355);
nand U4369 (N_4369,N_3340,N_3565);
nand U4370 (N_4370,N_3339,N_3226);
and U4371 (N_4371,N_3248,N_3412);
and U4372 (N_4372,N_3401,N_3564);
and U4373 (N_4373,N_3217,N_3017);
nor U4374 (N_4374,N_3414,N_3181);
nor U4375 (N_4375,N_3059,N_3030);
xnor U4376 (N_4376,N_3731,N_3187);
or U4377 (N_4377,N_3726,N_3334);
or U4378 (N_4378,N_3687,N_3192);
and U4379 (N_4379,N_3280,N_3110);
nor U4380 (N_4380,N_3075,N_3011);
and U4381 (N_4381,N_3239,N_3500);
and U4382 (N_4382,N_3329,N_3413);
or U4383 (N_4383,N_3324,N_3479);
xnor U4384 (N_4384,N_3735,N_3138);
nor U4385 (N_4385,N_3312,N_3035);
or U4386 (N_4386,N_3610,N_3649);
and U4387 (N_4387,N_3683,N_3470);
or U4388 (N_4388,N_3571,N_3350);
nand U4389 (N_4389,N_3505,N_3029);
and U4390 (N_4390,N_3282,N_3067);
nor U4391 (N_4391,N_3280,N_3140);
or U4392 (N_4392,N_3009,N_3435);
nor U4393 (N_4393,N_3521,N_3023);
and U4394 (N_4394,N_3734,N_3035);
nor U4395 (N_4395,N_3323,N_3028);
or U4396 (N_4396,N_3288,N_3443);
xnor U4397 (N_4397,N_3027,N_3219);
and U4398 (N_4398,N_3676,N_3713);
or U4399 (N_4399,N_3665,N_3028);
nor U4400 (N_4400,N_3271,N_3716);
nand U4401 (N_4401,N_3660,N_3379);
and U4402 (N_4402,N_3225,N_3400);
xnor U4403 (N_4403,N_3449,N_3026);
xor U4404 (N_4404,N_3204,N_3705);
nand U4405 (N_4405,N_3284,N_3615);
and U4406 (N_4406,N_3686,N_3715);
or U4407 (N_4407,N_3183,N_3098);
nor U4408 (N_4408,N_3296,N_3234);
and U4409 (N_4409,N_3696,N_3544);
nor U4410 (N_4410,N_3738,N_3061);
nand U4411 (N_4411,N_3105,N_3095);
or U4412 (N_4412,N_3262,N_3555);
or U4413 (N_4413,N_3279,N_3200);
or U4414 (N_4414,N_3744,N_3499);
and U4415 (N_4415,N_3530,N_3418);
xnor U4416 (N_4416,N_3299,N_3176);
nand U4417 (N_4417,N_3593,N_3080);
nor U4418 (N_4418,N_3122,N_3667);
nor U4419 (N_4419,N_3594,N_3097);
nor U4420 (N_4420,N_3359,N_3055);
nand U4421 (N_4421,N_3138,N_3540);
nor U4422 (N_4422,N_3351,N_3526);
nand U4423 (N_4423,N_3687,N_3321);
nor U4424 (N_4424,N_3608,N_3046);
or U4425 (N_4425,N_3580,N_3646);
or U4426 (N_4426,N_3159,N_3362);
nor U4427 (N_4427,N_3731,N_3403);
xnor U4428 (N_4428,N_3446,N_3362);
nor U4429 (N_4429,N_3283,N_3220);
or U4430 (N_4430,N_3329,N_3027);
nand U4431 (N_4431,N_3555,N_3007);
or U4432 (N_4432,N_3265,N_3288);
or U4433 (N_4433,N_3230,N_3693);
and U4434 (N_4434,N_3350,N_3367);
or U4435 (N_4435,N_3524,N_3399);
and U4436 (N_4436,N_3555,N_3322);
and U4437 (N_4437,N_3400,N_3317);
nand U4438 (N_4438,N_3230,N_3395);
nor U4439 (N_4439,N_3707,N_3575);
nor U4440 (N_4440,N_3516,N_3215);
nor U4441 (N_4441,N_3368,N_3372);
xnor U4442 (N_4442,N_3564,N_3719);
or U4443 (N_4443,N_3175,N_3650);
nand U4444 (N_4444,N_3079,N_3381);
nor U4445 (N_4445,N_3661,N_3115);
nand U4446 (N_4446,N_3606,N_3239);
and U4447 (N_4447,N_3534,N_3476);
nor U4448 (N_4448,N_3217,N_3583);
nand U4449 (N_4449,N_3710,N_3746);
and U4450 (N_4450,N_3177,N_3537);
and U4451 (N_4451,N_3457,N_3421);
or U4452 (N_4452,N_3696,N_3016);
nand U4453 (N_4453,N_3353,N_3402);
or U4454 (N_4454,N_3242,N_3346);
nand U4455 (N_4455,N_3070,N_3163);
nand U4456 (N_4456,N_3220,N_3192);
or U4457 (N_4457,N_3138,N_3508);
nor U4458 (N_4458,N_3534,N_3079);
and U4459 (N_4459,N_3515,N_3333);
nor U4460 (N_4460,N_3473,N_3396);
nand U4461 (N_4461,N_3463,N_3653);
and U4462 (N_4462,N_3064,N_3161);
xor U4463 (N_4463,N_3131,N_3663);
nand U4464 (N_4464,N_3166,N_3593);
or U4465 (N_4465,N_3360,N_3427);
nand U4466 (N_4466,N_3628,N_3645);
nand U4467 (N_4467,N_3699,N_3270);
nor U4468 (N_4468,N_3263,N_3496);
nor U4469 (N_4469,N_3181,N_3705);
xnor U4470 (N_4470,N_3432,N_3182);
nor U4471 (N_4471,N_3577,N_3294);
nor U4472 (N_4472,N_3430,N_3286);
and U4473 (N_4473,N_3564,N_3069);
and U4474 (N_4474,N_3204,N_3408);
or U4475 (N_4475,N_3596,N_3633);
or U4476 (N_4476,N_3093,N_3219);
nand U4477 (N_4477,N_3659,N_3529);
and U4478 (N_4478,N_3155,N_3697);
or U4479 (N_4479,N_3304,N_3107);
or U4480 (N_4480,N_3697,N_3422);
xnor U4481 (N_4481,N_3358,N_3456);
and U4482 (N_4482,N_3720,N_3020);
xor U4483 (N_4483,N_3376,N_3473);
nand U4484 (N_4484,N_3098,N_3574);
and U4485 (N_4485,N_3692,N_3489);
nor U4486 (N_4486,N_3491,N_3066);
nand U4487 (N_4487,N_3469,N_3135);
xnor U4488 (N_4488,N_3201,N_3636);
or U4489 (N_4489,N_3195,N_3573);
nand U4490 (N_4490,N_3494,N_3156);
nand U4491 (N_4491,N_3103,N_3059);
nand U4492 (N_4492,N_3255,N_3661);
or U4493 (N_4493,N_3048,N_3447);
or U4494 (N_4494,N_3682,N_3301);
xor U4495 (N_4495,N_3546,N_3331);
nand U4496 (N_4496,N_3371,N_3219);
nand U4497 (N_4497,N_3605,N_3533);
and U4498 (N_4498,N_3331,N_3218);
nor U4499 (N_4499,N_3547,N_3079);
or U4500 (N_4500,N_4133,N_4378);
and U4501 (N_4501,N_4037,N_4495);
nand U4502 (N_4502,N_4362,N_3917);
nand U4503 (N_4503,N_4425,N_4075);
nand U4504 (N_4504,N_3872,N_3892);
or U4505 (N_4505,N_3891,N_4089);
nor U4506 (N_4506,N_4262,N_3989);
nand U4507 (N_4507,N_4160,N_4418);
and U4508 (N_4508,N_4094,N_4124);
and U4509 (N_4509,N_4257,N_4103);
nand U4510 (N_4510,N_3995,N_3804);
nor U4511 (N_4511,N_3925,N_4175);
xor U4512 (N_4512,N_4063,N_4235);
xor U4513 (N_4513,N_4461,N_4408);
nor U4514 (N_4514,N_4048,N_4351);
nor U4515 (N_4515,N_3919,N_4392);
nor U4516 (N_4516,N_4131,N_4347);
or U4517 (N_4517,N_3902,N_4421);
nor U4518 (N_4518,N_3833,N_4014);
xor U4519 (N_4519,N_4333,N_4396);
nand U4520 (N_4520,N_3910,N_3881);
and U4521 (N_4521,N_4406,N_4422);
and U4522 (N_4522,N_4470,N_4491);
xnor U4523 (N_4523,N_4200,N_4376);
xor U4524 (N_4524,N_3807,N_4213);
and U4525 (N_4525,N_4332,N_4352);
nor U4526 (N_4526,N_4184,N_4182);
and U4527 (N_4527,N_4085,N_4442);
nor U4528 (N_4528,N_4122,N_3847);
nand U4529 (N_4529,N_4045,N_3815);
nand U4530 (N_4530,N_4278,N_3887);
nor U4531 (N_4531,N_3997,N_4210);
nand U4532 (N_4532,N_4290,N_4194);
nand U4533 (N_4533,N_3785,N_4368);
nor U4534 (N_4534,N_4449,N_3788);
xnor U4535 (N_4535,N_4393,N_4467);
or U4536 (N_4536,N_3894,N_3950);
nand U4537 (N_4537,N_4371,N_4439);
and U4538 (N_4538,N_4028,N_4060);
nor U4539 (N_4539,N_3914,N_3928);
xnor U4540 (N_4540,N_3784,N_3853);
nor U4541 (N_4541,N_4440,N_4460);
nor U4542 (N_4542,N_4321,N_4082);
nor U4543 (N_4543,N_3761,N_4212);
and U4544 (N_4544,N_3806,N_3777);
or U4545 (N_4545,N_3766,N_4125);
nor U4546 (N_4546,N_4404,N_3754);
and U4547 (N_4547,N_4030,N_4494);
nand U4548 (N_4548,N_4146,N_4346);
nor U4549 (N_4549,N_3759,N_3933);
nor U4550 (N_4550,N_4398,N_4118);
nor U4551 (N_4551,N_4019,N_4051);
or U4552 (N_4552,N_4056,N_4480);
nand U4553 (N_4553,N_4033,N_3857);
or U4554 (N_4554,N_3998,N_3852);
and U4555 (N_4555,N_4230,N_4203);
xor U4556 (N_4556,N_4098,N_3974);
and U4557 (N_4557,N_4369,N_3792);
xor U4558 (N_4558,N_4324,N_3967);
or U4559 (N_4559,N_4445,N_3948);
and U4560 (N_4560,N_4465,N_4026);
nor U4561 (N_4561,N_4229,N_4223);
and U4562 (N_4562,N_4293,N_4271);
and U4563 (N_4563,N_3913,N_4284);
nand U4564 (N_4564,N_4147,N_4226);
nand U4565 (N_4565,N_3886,N_3964);
or U4566 (N_4566,N_4297,N_4416);
or U4567 (N_4567,N_3813,N_3803);
or U4568 (N_4568,N_4486,N_3811);
nand U4569 (N_4569,N_3856,N_3757);
or U4570 (N_4570,N_4400,N_3775);
nand U4571 (N_4571,N_3812,N_4110);
xor U4572 (N_4572,N_4020,N_4473);
and U4573 (N_4573,N_4090,N_4342);
nand U4574 (N_4574,N_3888,N_4313);
nor U4575 (N_4575,N_4397,N_4143);
nand U4576 (N_4576,N_4062,N_4234);
nand U4577 (N_4577,N_4323,N_4220);
nand U4578 (N_4578,N_4101,N_4145);
nor U4579 (N_4579,N_4240,N_3973);
and U4580 (N_4580,N_4036,N_3823);
or U4581 (N_4581,N_4302,N_4214);
nor U4582 (N_4582,N_3979,N_4358);
xnor U4583 (N_4583,N_4039,N_4468);
xor U4584 (N_4584,N_4373,N_3843);
or U4585 (N_4585,N_4005,N_3970);
nor U4586 (N_4586,N_4107,N_4492);
nor U4587 (N_4587,N_3965,N_4064);
xor U4588 (N_4588,N_4413,N_4209);
or U4589 (N_4589,N_4218,N_4304);
or U4590 (N_4590,N_4247,N_3846);
nor U4591 (N_4591,N_3981,N_4242);
nor U4592 (N_4592,N_4032,N_3984);
nand U4593 (N_4593,N_3962,N_4379);
xor U4594 (N_4594,N_4169,N_3939);
or U4595 (N_4595,N_4205,N_3835);
nand U4596 (N_4596,N_4248,N_4488);
nand U4597 (N_4597,N_4289,N_4186);
nand U4598 (N_4598,N_3953,N_4104);
xor U4599 (N_4599,N_3924,N_4409);
nand U4600 (N_4600,N_4482,N_4034);
nand U4601 (N_4601,N_4010,N_3779);
or U4602 (N_4602,N_3916,N_4263);
nand U4603 (N_4603,N_4357,N_4129);
nand U4604 (N_4604,N_4306,N_4047);
nand U4605 (N_4605,N_3909,N_4399);
nor U4606 (N_4606,N_3845,N_3848);
nor U4607 (N_4607,N_3922,N_4275);
nor U4608 (N_4608,N_3960,N_4188);
or U4609 (N_4609,N_4299,N_4432);
xor U4610 (N_4610,N_3935,N_3762);
and U4611 (N_4611,N_4250,N_4419);
and U4612 (N_4612,N_4384,N_3946);
nor U4613 (N_4613,N_4068,N_4088);
xnor U4614 (N_4614,N_4154,N_4174);
xnor U4615 (N_4615,N_4374,N_4336);
and U4616 (N_4616,N_4080,N_3800);
nor U4617 (N_4617,N_4287,N_4448);
nand U4618 (N_4618,N_4318,N_4023);
and U4619 (N_4619,N_4149,N_3771);
and U4620 (N_4620,N_3791,N_3863);
nand U4621 (N_4621,N_3927,N_4029);
nor U4622 (N_4622,N_4076,N_4164);
nand U4623 (N_4623,N_4338,N_4326);
and U4624 (N_4624,N_3824,N_4121);
and U4625 (N_4625,N_4298,N_4158);
or U4626 (N_4626,N_4215,N_4095);
nor U4627 (N_4627,N_4006,N_4241);
nor U4628 (N_4628,N_3937,N_4017);
or U4629 (N_4629,N_4363,N_4252);
nand U4630 (N_4630,N_4462,N_3987);
nand U4631 (N_4631,N_3921,N_3790);
nand U4632 (N_4632,N_3929,N_4192);
nand U4633 (N_4633,N_4222,N_4433);
nor U4634 (N_4634,N_4128,N_4083);
or U4635 (N_4635,N_4345,N_3993);
nor U4636 (N_4636,N_4196,N_4420);
and U4637 (N_4637,N_4280,N_3770);
nand U4638 (N_4638,N_3977,N_3978);
nand U4639 (N_4639,N_3963,N_4141);
or U4640 (N_4640,N_4477,N_4489);
or U4641 (N_4641,N_4475,N_4407);
nand U4642 (N_4642,N_4191,N_3947);
xor U4643 (N_4643,N_4092,N_3911);
and U4644 (N_4644,N_4097,N_4208);
or U4645 (N_4645,N_3932,N_4484);
xor U4646 (N_4646,N_4153,N_3959);
or U4647 (N_4647,N_4386,N_4190);
and U4648 (N_4648,N_4024,N_4310);
nor U4649 (N_4649,N_4071,N_4403);
nor U4650 (N_4650,N_4211,N_3855);
nand U4651 (N_4651,N_4282,N_4086);
nor U4652 (N_4652,N_4007,N_3957);
nor U4653 (N_4653,N_3873,N_4243);
or U4654 (N_4654,N_4108,N_4339);
nand U4655 (N_4655,N_4219,N_3840);
nand U4656 (N_4656,N_3865,N_3915);
nor U4657 (N_4657,N_4109,N_3930);
nand U4658 (N_4658,N_4319,N_3841);
xnor U4659 (N_4659,N_3849,N_4344);
xor U4660 (N_4660,N_4389,N_4277);
nor U4661 (N_4661,N_4453,N_4189);
or U4662 (N_4662,N_4452,N_4053);
nand U4663 (N_4663,N_3988,N_4159);
or U4664 (N_4664,N_4325,N_4112);
nand U4665 (N_4665,N_4443,N_4180);
xnor U4666 (N_4666,N_4308,N_4274);
or U4667 (N_4667,N_4178,N_3765);
nand U4668 (N_4668,N_4424,N_4411);
xnor U4669 (N_4669,N_4315,N_4127);
and U4670 (N_4670,N_3763,N_3837);
nand U4671 (N_4671,N_4099,N_4165);
and U4672 (N_4672,N_4138,N_4349);
and U4673 (N_4673,N_4198,N_3890);
and U4674 (N_4674,N_3870,N_3944);
and U4675 (N_4675,N_4043,N_3842);
nand U4676 (N_4676,N_4172,N_4431);
or U4677 (N_4677,N_4327,N_4073);
and U4678 (N_4678,N_3758,N_3901);
or U4679 (N_4679,N_3829,N_4052);
and U4680 (N_4680,N_4091,N_3889);
xnor U4681 (N_4681,N_4206,N_3897);
or U4682 (N_4682,N_4116,N_3864);
nor U4683 (N_4683,N_4246,N_4027);
or U4684 (N_4684,N_4444,N_4295);
and U4685 (N_4685,N_3755,N_4055);
nand U4686 (N_4686,N_3808,N_4476);
and U4687 (N_4687,N_3908,N_4354);
or U4688 (N_4688,N_4231,N_3793);
nand U4689 (N_4689,N_4311,N_3831);
nand U4690 (N_4690,N_4372,N_4312);
nand U4691 (N_4691,N_3900,N_4309);
nor U4692 (N_4692,N_3912,N_4256);
nand U4693 (N_4693,N_4058,N_3884);
nand U4694 (N_4694,N_3810,N_4464);
nand U4695 (N_4695,N_4276,N_4305);
nand U4696 (N_4696,N_4016,N_4385);
nand U4697 (N_4697,N_4337,N_4292);
nor U4698 (N_4698,N_3874,N_4152);
or U4699 (N_4699,N_3828,N_4003);
or U4700 (N_4700,N_4365,N_4340);
and U4701 (N_4701,N_4140,N_4474);
and U4702 (N_4702,N_4417,N_3976);
and U4703 (N_4703,N_4427,N_4004);
xnor U4704 (N_4704,N_3877,N_4022);
or U4705 (N_4705,N_3936,N_3839);
nor U4706 (N_4706,N_3895,N_3868);
or U4707 (N_4707,N_4496,N_4359);
or U4708 (N_4708,N_3801,N_3776);
nor U4709 (N_4709,N_4167,N_4166);
or U4710 (N_4710,N_4267,N_4197);
nor U4711 (N_4711,N_4456,N_3955);
xnor U4712 (N_4712,N_3867,N_4307);
or U4713 (N_4713,N_3869,N_4114);
xnor U4714 (N_4714,N_4258,N_3904);
nor U4715 (N_4715,N_3906,N_4283);
and U4716 (N_4716,N_3954,N_3861);
nand U4717 (N_4717,N_4078,N_3943);
nand U4718 (N_4718,N_3972,N_4438);
nand U4719 (N_4719,N_4040,N_4328);
or U4720 (N_4720,N_4430,N_3926);
xor U4721 (N_4721,N_4294,N_4130);
nand U4722 (N_4722,N_4105,N_3781);
or U4723 (N_4723,N_4296,N_4395);
nand U4724 (N_4724,N_3994,N_3885);
nor U4725 (N_4725,N_4410,N_3898);
nor U4726 (N_4726,N_3805,N_4119);
or U4727 (N_4727,N_4377,N_4054);
or U4728 (N_4728,N_4300,N_4193);
nor U4729 (N_4729,N_4483,N_3951);
and U4730 (N_4730,N_3850,N_4157);
or U4731 (N_4731,N_4111,N_3796);
or U4732 (N_4732,N_4261,N_4335);
and U4733 (N_4733,N_4434,N_4132);
nor U4734 (N_4734,N_4177,N_3787);
and U4735 (N_4735,N_3799,N_4102);
nand U4736 (N_4736,N_3756,N_3920);
nand U4737 (N_4737,N_4270,N_4100);
and U4738 (N_4738,N_4050,N_4285);
xnor U4739 (N_4739,N_4435,N_4485);
or U4740 (N_4740,N_4471,N_3764);
xnor U4741 (N_4741,N_4322,N_4142);
xnor U4742 (N_4742,N_3825,N_4459);
or U4743 (N_4743,N_4015,N_4035);
and U4744 (N_4744,N_3999,N_4254);
nor U4745 (N_4745,N_4402,N_3778);
and U4746 (N_4746,N_4446,N_3938);
and U4747 (N_4747,N_3934,N_4170);
nand U4748 (N_4748,N_3838,N_3956);
or U4749 (N_4749,N_4176,N_4331);
xnor U4750 (N_4750,N_4233,N_3883);
nand U4751 (N_4751,N_4199,N_4139);
or U4752 (N_4752,N_3918,N_3996);
or U4753 (N_4753,N_3942,N_4227);
nor U4754 (N_4754,N_4320,N_4454);
and U4755 (N_4755,N_4273,N_3751);
nor U4756 (N_4756,N_4437,N_4245);
nor U4757 (N_4757,N_4136,N_4217);
or U4758 (N_4758,N_4002,N_4096);
xnor U4759 (N_4759,N_4087,N_4441);
and U4760 (N_4760,N_3858,N_4497);
nand U4761 (N_4761,N_4093,N_4120);
and U4762 (N_4762,N_4181,N_4429);
nor U4763 (N_4763,N_4106,N_4458);
or U4764 (N_4764,N_4239,N_4260);
nand U4765 (N_4765,N_3878,N_4394);
and U4766 (N_4766,N_4498,N_4117);
nor U4767 (N_4767,N_3975,N_4388);
or U4768 (N_4768,N_4135,N_3971);
and U4769 (N_4769,N_4066,N_4038);
nand U4770 (N_4770,N_4163,N_3814);
xnor U4771 (N_4771,N_4162,N_4367);
nor U4772 (N_4772,N_4207,N_3783);
nor U4773 (N_4773,N_4046,N_3896);
nand U4774 (N_4774,N_4259,N_3931);
xnor U4775 (N_4775,N_3860,N_4356);
and U4776 (N_4776,N_4341,N_4081);
and U4777 (N_4777,N_4171,N_4405);
and U4778 (N_4778,N_3798,N_4065);
nor U4779 (N_4779,N_4353,N_4375);
nor U4780 (N_4780,N_4330,N_4021);
nor U4781 (N_4781,N_3822,N_4264);
or U4782 (N_4782,N_4202,N_3985);
or U4783 (N_4783,N_4291,N_4079);
nand U4784 (N_4784,N_4244,N_4195);
nor U4785 (N_4785,N_3820,N_4450);
nor U4786 (N_4786,N_3818,N_4478);
or U4787 (N_4787,N_4481,N_3862);
or U4788 (N_4788,N_4401,N_4070);
or U4789 (N_4789,N_4150,N_3923);
and U4790 (N_4790,N_4255,N_4072);
nor U4791 (N_4791,N_4451,N_4301);
and U4792 (N_4792,N_4382,N_3980);
or U4793 (N_4793,N_4155,N_4390);
nor U4794 (N_4794,N_3958,N_3899);
nand U4795 (N_4795,N_4348,N_3986);
xnor U4796 (N_4796,N_3871,N_3795);
nor U4797 (N_4797,N_4161,N_4134);
nor U4798 (N_4798,N_4236,N_3767);
nand U4799 (N_4799,N_4077,N_4251);
nand U4800 (N_4800,N_4185,N_3752);
xnor U4801 (N_4801,N_4115,N_4415);
nand U4802 (N_4802,N_4499,N_3830);
nand U4803 (N_4803,N_4237,N_4041);
or U4804 (N_4804,N_4355,N_3816);
nand U4805 (N_4805,N_4423,N_4216);
or U4806 (N_4806,N_4487,N_4316);
or U4807 (N_4807,N_4084,N_3827);
xnor U4808 (N_4808,N_4286,N_4472);
and U4809 (N_4809,N_4364,N_3832);
and U4810 (N_4810,N_4329,N_4069);
nor U4811 (N_4811,N_4168,N_3940);
nor U4812 (N_4812,N_4001,N_4279);
nor U4813 (N_4813,N_4387,N_3949);
and U4814 (N_4814,N_3880,N_3797);
and U4815 (N_4815,N_3769,N_4228);
nor U4816 (N_4816,N_3794,N_4018);
xor U4817 (N_4817,N_3750,N_4317);
nor U4818 (N_4818,N_4201,N_3780);
and U4819 (N_4819,N_4059,N_4426);
nand U4820 (N_4820,N_3905,N_3772);
nor U4821 (N_4821,N_4123,N_3991);
or U4822 (N_4822,N_4113,N_3893);
xor U4823 (N_4823,N_4288,N_4334);
nor U4824 (N_4824,N_4221,N_4490);
xor U4825 (N_4825,N_4187,N_4151);
xnor U4826 (N_4826,N_3859,N_3851);
and U4827 (N_4827,N_4493,N_3819);
or U4828 (N_4828,N_4391,N_3760);
nor U4829 (N_4829,N_4232,N_4225);
nand U4830 (N_4830,N_4013,N_4061);
or U4831 (N_4831,N_4381,N_4025);
or U4832 (N_4832,N_3983,N_4126);
nor U4833 (N_4833,N_3903,N_4455);
nor U4834 (N_4834,N_4303,N_3992);
nor U4835 (N_4835,N_3866,N_4224);
xor U4836 (N_4836,N_4009,N_4466);
nor U4837 (N_4837,N_4204,N_4011);
xnor U4838 (N_4838,N_4380,N_4148);
and U4839 (N_4839,N_3789,N_3836);
nand U4840 (N_4840,N_4057,N_4457);
xor U4841 (N_4841,N_3809,N_3990);
nor U4842 (N_4842,N_4067,N_3826);
nand U4843 (N_4843,N_4008,N_3968);
and U4844 (N_4844,N_4074,N_3802);
nand U4845 (N_4845,N_4272,N_4469);
nor U4846 (N_4846,N_4042,N_4436);
nor U4847 (N_4847,N_3774,N_4479);
xnor U4848 (N_4848,N_3952,N_3945);
or U4849 (N_4849,N_4414,N_4265);
or U4850 (N_4850,N_3821,N_4463);
and U4851 (N_4851,N_4350,N_4281);
nor U4852 (N_4852,N_4179,N_3941);
nor U4853 (N_4853,N_4266,N_3844);
nor U4854 (N_4854,N_3834,N_3753);
nor U4855 (N_4855,N_3773,N_4253);
and U4856 (N_4856,N_4137,N_4156);
and U4857 (N_4857,N_4049,N_3875);
nand U4858 (N_4858,N_4412,N_3961);
and U4859 (N_4859,N_4370,N_4343);
xnor U4860 (N_4860,N_3817,N_4428);
or U4861 (N_4861,N_3854,N_4360);
nand U4862 (N_4862,N_4383,N_4447);
nor U4863 (N_4863,N_4000,N_3876);
xor U4864 (N_4864,N_4031,N_3786);
or U4865 (N_4865,N_4012,N_4173);
and U4866 (N_4866,N_3768,N_3882);
xor U4867 (N_4867,N_4044,N_4238);
nand U4868 (N_4868,N_4249,N_4314);
and U4869 (N_4869,N_3982,N_4183);
or U4870 (N_4870,N_3966,N_3782);
nand U4871 (N_4871,N_4144,N_3907);
nand U4872 (N_4872,N_3879,N_4366);
xor U4873 (N_4873,N_4268,N_4269);
nor U4874 (N_4874,N_4361,N_3969);
or U4875 (N_4875,N_4033,N_4324);
nor U4876 (N_4876,N_3835,N_4224);
nor U4877 (N_4877,N_3949,N_4415);
or U4878 (N_4878,N_3989,N_4074);
or U4879 (N_4879,N_4344,N_4441);
or U4880 (N_4880,N_3892,N_4036);
or U4881 (N_4881,N_4038,N_4078);
nor U4882 (N_4882,N_4472,N_4050);
and U4883 (N_4883,N_4189,N_3991);
nor U4884 (N_4884,N_3759,N_4258);
and U4885 (N_4885,N_4164,N_4098);
nor U4886 (N_4886,N_4318,N_3766);
nand U4887 (N_4887,N_4471,N_3758);
nand U4888 (N_4888,N_3836,N_4361);
nor U4889 (N_4889,N_3946,N_4232);
or U4890 (N_4890,N_4046,N_4068);
or U4891 (N_4891,N_4428,N_4470);
xor U4892 (N_4892,N_4240,N_4209);
nor U4893 (N_4893,N_4019,N_4476);
nand U4894 (N_4894,N_3820,N_3772);
nor U4895 (N_4895,N_4266,N_3821);
or U4896 (N_4896,N_4083,N_4217);
nand U4897 (N_4897,N_4051,N_3894);
and U4898 (N_4898,N_4020,N_3976);
and U4899 (N_4899,N_3989,N_4412);
and U4900 (N_4900,N_3824,N_4290);
and U4901 (N_4901,N_4113,N_4077);
or U4902 (N_4902,N_4122,N_3795);
nand U4903 (N_4903,N_4248,N_4244);
and U4904 (N_4904,N_4444,N_4160);
nand U4905 (N_4905,N_3919,N_4248);
nand U4906 (N_4906,N_4412,N_4386);
or U4907 (N_4907,N_4218,N_4057);
and U4908 (N_4908,N_4484,N_3887);
xor U4909 (N_4909,N_4090,N_3780);
or U4910 (N_4910,N_4093,N_3912);
and U4911 (N_4911,N_3905,N_4287);
and U4912 (N_4912,N_4220,N_3811);
and U4913 (N_4913,N_4144,N_4311);
and U4914 (N_4914,N_4235,N_4303);
nor U4915 (N_4915,N_3906,N_3932);
nor U4916 (N_4916,N_3970,N_4127);
and U4917 (N_4917,N_4238,N_4338);
nor U4918 (N_4918,N_3995,N_4271);
nor U4919 (N_4919,N_4461,N_3920);
nor U4920 (N_4920,N_4379,N_4150);
nand U4921 (N_4921,N_3766,N_3995);
or U4922 (N_4922,N_4068,N_3976);
or U4923 (N_4923,N_3827,N_4261);
and U4924 (N_4924,N_4064,N_3756);
xor U4925 (N_4925,N_4441,N_4468);
nand U4926 (N_4926,N_3958,N_3901);
xnor U4927 (N_4927,N_4167,N_3990);
nor U4928 (N_4928,N_4454,N_4058);
or U4929 (N_4929,N_4026,N_3858);
or U4930 (N_4930,N_4371,N_4292);
nand U4931 (N_4931,N_4380,N_3887);
or U4932 (N_4932,N_4317,N_4215);
or U4933 (N_4933,N_3877,N_4471);
nor U4934 (N_4934,N_3912,N_4032);
xnor U4935 (N_4935,N_3851,N_3764);
and U4936 (N_4936,N_3836,N_3827);
or U4937 (N_4937,N_3910,N_4354);
xnor U4938 (N_4938,N_3791,N_3962);
nand U4939 (N_4939,N_4008,N_4175);
or U4940 (N_4940,N_3987,N_4358);
nand U4941 (N_4941,N_3825,N_4189);
nor U4942 (N_4942,N_3977,N_3960);
and U4943 (N_4943,N_4468,N_3912);
and U4944 (N_4944,N_4480,N_4406);
and U4945 (N_4945,N_4225,N_4162);
nand U4946 (N_4946,N_4120,N_3969);
nor U4947 (N_4947,N_4083,N_4050);
xor U4948 (N_4948,N_3802,N_4239);
nand U4949 (N_4949,N_4385,N_4448);
nand U4950 (N_4950,N_3969,N_4420);
or U4951 (N_4951,N_4441,N_4263);
or U4952 (N_4952,N_4459,N_4253);
nand U4953 (N_4953,N_4434,N_4024);
and U4954 (N_4954,N_4495,N_3812);
nand U4955 (N_4955,N_3788,N_4329);
nor U4956 (N_4956,N_4078,N_4483);
and U4957 (N_4957,N_4389,N_4110);
and U4958 (N_4958,N_4227,N_3980);
or U4959 (N_4959,N_4097,N_4299);
or U4960 (N_4960,N_4306,N_4409);
or U4961 (N_4961,N_4150,N_3769);
nand U4962 (N_4962,N_3775,N_3863);
nand U4963 (N_4963,N_3788,N_3896);
or U4964 (N_4964,N_3981,N_4498);
xor U4965 (N_4965,N_3981,N_4478);
and U4966 (N_4966,N_3783,N_3822);
nand U4967 (N_4967,N_3812,N_4343);
nand U4968 (N_4968,N_4056,N_4273);
nor U4969 (N_4969,N_4273,N_3972);
xnor U4970 (N_4970,N_4290,N_3845);
and U4971 (N_4971,N_4230,N_4211);
and U4972 (N_4972,N_3772,N_4065);
or U4973 (N_4973,N_3794,N_3988);
xnor U4974 (N_4974,N_4010,N_4193);
nor U4975 (N_4975,N_4107,N_3924);
xnor U4976 (N_4976,N_4297,N_3999);
and U4977 (N_4977,N_4328,N_4434);
nor U4978 (N_4978,N_3984,N_4410);
and U4979 (N_4979,N_3960,N_4027);
and U4980 (N_4980,N_4416,N_4183);
or U4981 (N_4981,N_4073,N_3843);
nand U4982 (N_4982,N_3801,N_4150);
nand U4983 (N_4983,N_4260,N_3870);
nor U4984 (N_4984,N_3950,N_4421);
or U4985 (N_4985,N_3940,N_4006);
nor U4986 (N_4986,N_3912,N_4477);
and U4987 (N_4987,N_4278,N_4032);
and U4988 (N_4988,N_4488,N_4411);
and U4989 (N_4989,N_4214,N_4146);
nand U4990 (N_4990,N_4408,N_4172);
xnor U4991 (N_4991,N_4084,N_4053);
and U4992 (N_4992,N_4462,N_3759);
or U4993 (N_4993,N_4481,N_3792);
nand U4994 (N_4994,N_4178,N_4182);
or U4995 (N_4995,N_4099,N_3955);
and U4996 (N_4996,N_3909,N_4417);
and U4997 (N_4997,N_4035,N_4183);
nor U4998 (N_4998,N_4214,N_4244);
xnor U4999 (N_4999,N_4061,N_3767);
nand U5000 (N_5000,N_3946,N_4114);
nand U5001 (N_5001,N_4409,N_4235);
xnor U5002 (N_5002,N_3922,N_4312);
nor U5003 (N_5003,N_3773,N_4096);
nor U5004 (N_5004,N_4066,N_4019);
nor U5005 (N_5005,N_3846,N_3800);
nand U5006 (N_5006,N_3764,N_3834);
and U5007 (N_5007,N_3769,N_3934);
nor U5008 (N_5008,N_4101,N_3926);
nor U5009 (N_5009,N_3849,N_4010);
and U5010 (N_5010,N_3933,N_4045);
and U5011 (N_5011,N_4236,N_4178);
and U5012 (N_5012,N_4282,N_3832);
and U5013 (N_5013,N_4313,N_4496);
xnor U5014 (N_5014,N_4030,N_3810);
and U5015 (N_5015,N_4241,N_4296);
or U5016 (N_5016,N_4431,N_4222);
nor U5017 (N_5017,N_3966,N_4102);
and U5018 (N_5018,N_4380,N_4074);
nor U5019 (N_5019,N_3894,N_3982);
nand U5020 (N_5020,N_4037,N_3835);
or U5021 (N_5021,N_3847,N_3965);
or U5022 (N_5022,N_4140,N_4081);
nor U5023 (N_5023,N_4108,N_4309);
nand U5024 (N_5024,N_3811,N_3792);
or U5025 (N_5025,N_4255,N_4174);
and U5026 (N_5026,N_3764,N_4187);
nor U5027 (N_5027,N_4266,N_3925);
nor U5028 (N_5028,N_3909,N_4478);
nor U5029 (N_5029,N_4106,N_4359);
and U5030 (N_5030,N_4286,N_3944);
nand U5031 (N_5031,N_4226,N_4411);
or U5032 (N_5032,N_3910,N_4337);
nor U5033 (N_5033,N_4496,N_4230);
or U5034 (N_5034,N_3817,N_4396);
nand U5035 (N_5035,N_3909,N_4379);
or U5036 (N_5036,N_3909,N_4346);
nor U5037 (N_5037,N_4094,N_4300);
and U5038 (N_5038,N_4272,N_4027);
xnor U5039 (N_5039,N_4184,N_4281);
xnor U5040 (N_5040,N_4025,N_4347);
and U5041 (N_5041,N_3850,N_4021);
nand U5042 (N_5042,N_4091,N_3793);
nor U5043 (N_5043,N_3903,N_3940);
xnor U5044 (N_5044,N_4342,N_4339);
or U5045 (N_5045,N_4223,N_3936);
or U5046 (N_5046,N_3797,N_4447);
nor U5047 (N_5047,N_4182,N_4132);
nand U5048 (N_5048,N_4165,N_4193);
nor U5049 (N_5049,N_3750,N_3873);
xnor U5050 (N_5050,N_4068,N_3941);
or U5051 (N_5051,N_4185,N_4090);
or U5052 (N_5052,N_4476,N_3956);
and U5053 (N_5053,N_4222,N_3952);
and U5054 (N_5054,N_3819,N_4235);
nand U5055 (N_5055,N_3871,N_3815);
or U5056 (N_5056,N_4411,N_4355);
nor U5057 (N_5057,N_4120,N_4045);
nor U5058 (N_5058,N_4417,N_4258);
nor U5059 (N_5059,N_3925,N_4359);
nand U5060 (N_5060,N_4069,N_4040);
xor U5061 (N_5061,N_4211,N_3891);
and U5062 (N_5062,N_4379,N_4054);
nand U5063 (N_5063,N_3853,N_4308);
or U5064 (N_5064,N_4075,N_4155);
and U5065 (N_5065,N_4208,N_3898);
nand U5066 (N_5066,N_3973,N_4176);
or U5067 (N_5067,N_4405,N_3963);
and U5068 (N_5068,N_4283,N_4035);
nand U5069 (N_5069,N_4213,N_4153);
and U5070 (N_5070,N_4214,N_4402);
or U5071 (N_5071,N_4370,N_4045);
xor U5072 (N_5072,N_3765,N_3920);
nor U5073 (N_5073,N_4044,N_4182);
or U5074 (N_5074,N_3816,N_4010);
nand U5075 (N_5075,N_4071,N_3841);
or U5076 (N_5076,N_4466,N_4132);
and U5077 (N_5077,N_3885,N_4052);
and U5078 (N_5078,N_3795,N_4034);
and U5079 (N_5079,N_4086,N_4038);
nor U5080 (N_5080,N_3994,N_4023);
nor U5081 (N_5081,N_4299,N_4321);
and U5082 (N_5082,N_3921,N_4367);
nor U5083 (N_5083,N_3839,N_3857);
nor U5084 (N_5084,N_4267,N_4149);
xor U5085 (N_5085,N_4392,N_4212);
or U5086 (N_5086,N_3957,N_4215);
nor U5087 (N_5087,N_3923,N_4312);
nor U5088 (N_5088,N_3833,N_3995);
or U5089 (N_5089,N_3970,N_3980);
and U5090 (N_5090,N_3788,N_4263);
nand U5091 (N_5091,N_4397,N_4077);
and U5092 (N_5092,N_4233,N_4346);
and U5093 (N_5093,N_4395,N_3777);
nor U5094 (N_5094,N_4478,N_4279);
nor U5095 (N_5095,N_4384,N_4230);
nand U5096 (N_5096,N_3901,N_4242);
and U5097 (N_5097,N_4188,N_4152);
and U5098 (N_5098,N_4256,N_4368);
nand U5099 (N_5099,N_3872,N_4145);
nand U5100 (N_5100,N_3782,N_4199);
nand U5101 (N_5101,N_4118,N_3877);
or U5102 (N_5102,N_4415,N_4116);
and U5103 (N_5103,N_4053,N_4111);
xor U5104 (N_5104,N_3918,N_4240);
and U5105 (N_5105,N_3776,N_4016);
and U5106 (N_5106,N_3914,N_4194);
and U5107 (N_5107,N_4065,N_3980);
xnor U5108 (N_5108,N_3832,N_4340);
or U5109 (N_5109,N_3912,N_4475);
nor U5110 (N_5110,N_4268,N_4319);
nor U5111 (N_5111,N_4249,N_3795);
and U5112 (N_5112,N_3945,N_4198);
nand U5113 (N_5113,N_4407,N_3797);
nand U5114 (N_5114,N_4070,N_4195);
or U5115 (N_5115,N_4210,N_4444);
nor U5116 (N_5116,N_4413,N_4472);
or U5117 (N_5117,N_4138,N_4139);
nand U5118 (N_5118,N_4186,N_3775);
and U5119 (N_5119,N_4388,N_4187);
nor U5120 (N_5120,N_4362,N_4220);
or U5121 (N_5121,N_3828,N_3944);
or U5122 (N_5122,N_3794,N_3871);
nand U5123 (N_5123,N_3763,N_3896);
and U5124 (N_5124,N_3842,N_4050);
nand U5125 (N_5125,N_4040,N_3893);
nand U5126 (N_5126,N_3797,N_4306);
xnor U5127 (N_5127,N_3764,N_3945);
nand U5128 (N_5128,N_4100,N_4127);
xnor U5129 (N_5129,N_4198,N_4111);
nor U5130 (N_5130,N_3971,N_4347);
nand U5131 (N_5131,N_4304,N_4454);
nand U5132 (N_5132,N_3973,N_4496);
nor U5133 (N_5133,N_3758,N_4392);
nand U5134 (N_5134,N_4118,N_4442);
nor U5135 (N_5135,N_4172,N_3930);
and U5136 (N_5136,N_4302,N_3829);
nand U5137 (N_5137,N_3964,N_4482);
nand U5138 (N_5138,N_4216,N_3999);
and U5139 (N_5139,N_4309,N_3790);
and U5140 (N_5140,N_4305,N_4314);
nand U5141 (N_5141,N_3980,N_4086);
or U5142 (N_5142,N_4155,N_4449);
nand U5143 (N_5143,N_3755,N_4496);
xor U5144 (N_5144,N_4290,N_3915);
nand U5145 (N_5145,N_3987,N_4111);
nand U5146 (N_5146,N_4289,N_3968);
nand U5147 (N_5147,N_3912,N_4235);
and U5148 (N_5148,N_4074,N_4110);
and U5149 (N_5149,N_4052,N_4461);
nand U5150 (N_5150,N_4087,N_4367);
nand U5151 (N_5151,N_4406,N_4424);
or U5152 (N_5152,N_4408,N_4193);
or U5153 (N_5153,N_3825,N_3962);
xor U5154 (N_5154,N_4095,N_4261);
nor U5155 (N_5155,N_3805,N_3950);
nor U5156 (N_5156,N_3772,N_4483);
nand U5157 (N_5157,N_4456,N_3753);
nor U5158 (N_5158,N_4277,N_3875);
xor U5159 (N_5159,N_4053,N_4406);
nand U5160 (N_5160,N_3830,N_4325);
and U5161 (N_5161,N_3806,N_3775);
nor U5162 (N_5162,N_3834,N_3879);
nor U5163 (N_5163,N_4148,N_4484);
nand U5164 (N_5164,N_4398,N_4203);
xnor U5165 (N_5165,N_3842,N_4347);
and U5166 (N_5166,N_4334,N_4302);
and U5167 (N_5167,N_3938,N_4499);
or U5168 (N_5168,N_4249,N_3904);
nand U5169 (N_5169,N_4177,N_4270);
nor U5170 (N_5170,N_4417,N_4103);
or U5171 (N_5171,N_4189,N_4301);
nand U5172 (N_5172,N_4484,N_4057);
nor U5173 (N_5173,N_4226,N_4128);
nor U5174 (N_5174,N_4314,N_3777);
and U5175 (N_5175,N_3943,N_4484);
and U5176 (N_5176,N_4214,N_4126);
nor U5177 (N_5177,N_4375,N_4357);
nand U5178 (N_5178,N_3932,N_4137);
nor U5179 (N_5179,N_4407,N_4200);
and U5180 (N_5180,N_4251,N_4201);
and U5181 (N_5181,N_4400,N_4192);
nand U5182 (N_5182,N_3932,N_4101);
and U5183 (N_5183,N_4127,N_3769);
nand U5184 (N_5184,N_3965,N_4126);
nor U5185 (N_5185,N_4219,N_4392);
and U5186 (N_5186,N_4281,N_4139);
or U5187 (N_5187,N_4296,N_4216);
or U5188 (N_5188,N_4095,N_4028);
and U5189 (N_5189,N_4160,N_4337);
and U5190 (N_5190,N_4160,N_4082);
and U5191 (N_5191,N_3963,N_4325);
or U5192 (N_5192,N_4379,N_4377);
or U5193 (N_5193,N_4055,N_4214);
nand U5194 (N_5194,N_3855,N_4445);
or U5195 (N_5195,N_4042,N_4393);
or U5196 (N_5196,N_3924,N_4403);
nor U5197 (N_5197,N_3994,N_3837);
nand U5198 (N_5198,N_4010,N_3844);
and U5199 (N_5199,N_3752,N_3925);
and U5200 (N_5200,N_4045,N_3849);
nand U5201 (N_5201,N_4167,N_4177);
xor U5202 (N_5202,N_3917,N_4149);
nor U5203 (N_5203,N_3797,N_4175);
nand U5204 (N_5204,N_4044,N_3851);
nor U5205 (N_5205,N_4385,N_3965);
or U5206 (N_5206,N_4347,N_4449);
nand U5207 (N_5207,N_4190,N_4282);
and U5208 (N_5208,N_4039,N_4497);
nand U5209 (N_5209,N_3789,N_4033);
and U5210 (N_5210,N_4052,N_4159);
nor U5211 (N_5211,N_4211,N_4178);
or U5212 (N_5212,N_4129,N_4221);
nor U5213 (N_5213,N_4178,N_4000);
xnor U5214 (N_5214,N_3902,N_4083);
nor U5215 (N_5215,N_3979,N_3917);
nor U5216 (N_5216,N_3843,N_4470);
nand U5217 (N_5217,N_4477,N_4171);
xor U5218 (N_5218,N_4363,N_4096);
or U5219 (N_5219,N_4146,N_3895);
nor U5220 (N_5220,N_3998,N_3911);
and U5221 (N_5221,N_4277,N_3860);
or U5222 (N_5222,N_4061,N_4106);
or U5223 (N_5223,N_4039,N_4162);
nor U5224 (N_5224,N_3960,N_4496);
and U5225 (N_5225,N_4389,N_4249);
nor U5226 (N_5226,N_4072,N_3875);
nand U5227 (N_5227,N_3869,N_3868);
nor U5228 (N_5228,N_4268,N_4286);
and U5229 (N_5229,N_4078,N_3791);
or U5230 (N_5230,N_4030,N_4140);
nor U5231 (N_5231,N_4457,N_3931);
or U5232 (N_5232,N_4354,N_4266);
and U5233 (N_5233,N_4247,N_4004);
nand U5234 (N_5234,N_4091,N_4296);
nor U5235 (N_5235,N_4405,N_4022);
or U5236 (N_5236,N_4197,N_3961);
nand U5237 (N_5237,N_3771,N_3905);
nor U5238 (N_5238,N_4142,N_3883);
nand U5239 (N_5239,N_4454,N_4461);
and U5240 (N_5240,N_3833,N_4228);
or U5241 (N_5241,N_4368,N_4196);
nor U5242 (N_5242,N_4157,N_4391);
nor U5243 (N_5243,N_4137,N_4084);
and U5244 (N_5244,N_3765,N_3799);
and U5245 (N_5245,N_3995,N_3836);
nand U5246 (N_5246,N_4256,N_4416);
nor U5247 (N_5247,N_4475,N_4351);
nor U5248 (N_5248,N_3916,N_4288);
nor U5249 (N_5249,N_3919,N_3826);
and U5250 (N_5250,N_4607,N_5121);
nor U5251 (N_5251,N_4641,N_5174);
or U5252 (N_5252,N_5203,N_5100);
nand U5253 (N_5253,N_5195,N_5166);
or U5254 (N_5254,N_4866,N_4980);
nor U5255 (N_5255,N_4803,N_5101);
or U5256 (N_5256,N_4945,N_4736);
and U5257 (N_5257,N_4507,N_4824);
nor U5258 (N_5258,N_4617,N_4990);
or U5259 (N_5259,N_5171,N_4875);
nor U5260 (N_5260,N_4602,N_5050);
or U5261 (N_5261,N_4960,N_4936);
or U5262 (N_5262,N_4531,N_4819);
nor U5263 (N_5263,N_5069,N_5149);
xnor U5264 (N_5264,N_5218,N_4884);
xnor U5265 (N_5265,N_5191,N_4744);
xor U5266 (N_5266,N_4780,N_5172);
nor U5267 (N_5267,N_4688,N_4995);
and U5268 (N_5268,N_4613,N_4991);
nand U5269 (N_5269,N_4532,N_5045);
or U5270 (N_5270,N_5041,N_4652);
or U5271 (N_5271,N_5066,N_4810);
nor U5272 (N_5272,N_5159,N_4895);
nand U5273 (N_5273,N_4592,N_5161);
nor U5274 (N_5274,N_4709,N_5020);
or U5275 (N_5275,N_4831,N_5219);
or U5276 (N_5276,N_4615,N_4983);
nor U5277 (N_5277,N_5181,N_5094);
nor U5278 (N_5278,N_4850,N_5182);
and U5279 (N_5279,N_5215,N_4857);
nand U5280 (N_5280,N_5241,N_5225);
or U5281 (N_5281,N_4612,N_5097);
nand U5282 (N_5282,N_4528,N_4878);
xor U5283 (N_5283,N_4811,N_4835);
nor U5284 (N_5284,N_4791,N_5247);
nor U5285 (N_5285,N_4674,N_4972);
and U5286 (N_5286,N_5137,N_5236);
xnor U5287 (N_5287,N_5011,N_4921);
or U5288 (N_5288,N_4651,N_4925);
nor U5289 (N_5289,N_4687,N_5115);
or U5290 (N_5290,N_4695,N_4992);
or U5291 (N_5291,N_4853,N_4816);
and U5292 (N_5292,N_4950,N_5063);
nor U5293 (N_5293,N_5070,N_5139);
nand U5294 (N_5294,N_4545,N_4978);
xnor U5295 (N_5295,N_4685,N_4920);
or U5296 (N_5296,N_4672,N_4629);
nor U5297 (N_5297,N_4970,N_4976);
nand U5298 (N_5298,N_4724,N_5224);
nand U5299 (N_5299,N_5245,N_4514);
and U5300 (N_5300,N_5013,N_4900);
nor U5301 (N_5301,N_4564,N_5228);
nor U5302 (N_5302,N_5235,N_4733);
nand U5303 (N_5303,N_5096,N_4509);
nand U5304 (N_5304,N_4745,N_4975);
and U5305 (N_5305,N_4626,N_4984);
or U5306 (N_5306,N_5176,N_5160);
nor U5307 (N_5307,N_5105,N_4817);
or U5308 (N_5308,N_5022,N_4655);
nand U5309 (N_5309,N_4735,N_4918);
nand U5310 (N_5310,N_5158,N_4877);
nor U5311 (N_5311,N_4833,N_4986);
nor U5312 (N_5312,N_4597,N_4851);
or U5313 (N_5313,N_4790,N_4845);
or U5314 (N_5314,N_4912,N_4746);
or U5315 (N_5315,N_4739,N_5221);
and U5316 (N_5316,N_5116,N_4600);
nor U5317 (N_5317,N_4549,N_4692);
or U5318 (N_5318,N_4806,N_4580);
nor U5319 (N_5319,N_5086,N_4708);
and U5320 (N_5320,N_4722,N_4561);
nand U5321 (N_5321,N_5140,N_5056);
nor U5322 (N_5322,N_4684,N_4729);
nor U5323 (N_5323,N_4516,N_5111);
and U5324 (N_5324,N_5090,N_4798);
and U5325 (N_5325,N_5244,N_4563);
nand U5326 (N_5326,N_5146,N_5223);
nand U5327 (N_5327,N_4794,N_4671);
nor U5328 (N_5328,N_5125,N_5205);
nor U5329 (N_5329,N_5145,N_4604);
nand U5330 (N_5330,N_4996,N_4732);
nor U5331 (N_5331,N_4734,N_4934);
and U5332 (N_5332,N_5000,N_5135);
or U5333 (N_5333,N_4873,N_4951);
and U5334 (N_5334,N_5201,N_5151);
or U5335 (N_5335,N_4874,N_5026);
and U5336 (N_5336,N_5134,N_4681);
or U5337 (N_5337,N_4620,N_5231);
nor U5338 (N_5338,N_5153,N_4969);
xor U5339 (N_5339,N_5027,N_4955);
and U5340 (N_5340,N_5177,N_4664);
or U5341 (N_5341,N_4616,N_4503);
or U5342 (N_5342,N_5222,N_4582);
nand U5343 (N_5343,N_5104,N_4520);
nor U5344 (N_5344,N_5242,N_4640);
or U5345 (N_5345,N_4930,N_4855);
nand U5346 (N_5346,N_5192,N_4710);
or U5347 (N_5347,N_4784,N_5129);
nor U5348 (N_5348,N_5138,N_4959);
xnor U5349 (N_5349,N_4775,N_4856);
nor U5350 (N_5350,N_4890,N_5091);
or U5351 (N_5351,N_4658,N_5190);
or U5352 (N_5352,N_4979,N_4994);
or U5353 (N_5353,N_4829,N_5187);
and U5354 (N_5354,N_4800,N_4888);
nor U5355 (N_5355,N_4630,N_4511);
xnor U5356 (N_5356,N_4909,N_4590);
nand U5357 (N_5357,N_4847,N_5233);
nor U5358 (N_5358,N_5024,N_4740);
nand U5359 (N_5359,N_4765,N_5180);
nand U5360 (N_5360,N_4501,N_4749);
nor U5361 (N_5361,N_4832,N_4727);
or U5362 (N_5362,N_5015,N_4720);
nand U5363 (N_5363,N_4965,N_5120);
and U5364 (N_5364,N_4534,N_5142);
nor U5365 (N_5365,N_5232,N_4789);
or U5366 (N_5366,N_5162,N_4715);
nand U5367 (N_5367,N_4657,N_5119);
xor U5368 (N_5368,N_5112,N_4656);
and U5369 (N_5369,N_4842,N_4881);
nand U5370 (N_5370,N_4947,N_5124);
and U5371 (N_5371,N_4578,N_4863);
nor U5372 (N_5372,N_5229,N_5189);
nor U5373 (N_5373,N_4714,N_4702);
nor U5374 (N_5374,N_5117,N_5002);
and U5375 (N_5375,N_4587,N_5183);
nand U5376 (N_5376,N_4682,N_4570);
and U5377 (N_5377,N_5230,N_4525);
xor U5378 (N_5378,N_4669,N_5110);
nand U5379 (N_5379,N_4987,N_5216);
nand U5380 (N_5380,N_4772,N_4982);
xnor U5381 (N_5381,N_5003,N_5240);
nand U5382 (N_5382,N_4974,N_4956);
or U5383 (N_5383,N_4805,N_4500);
or U5384 (N_5384,N_4823,N_4954);
and U5385 (N_5385,N_4953,N_4539);
nor U5386 (N_5386,N_5073,N_4802);
nand U5387 (N_5387,N_4773,N_5025);
xnor U5388 (N_5388,N_5239,N_4760);
nor U5389 (N_5389,N_4861,N_5102);
or U5390 (N_5390,N_4697,N_5147);
nor U5391 (N_5391,N_4860,N_4826);
nor U5392 (N_5392,N_5061,N_4968);
and U5393 (N_5393,N_4661,N_4717);
nor U5394 (N_5394,N_4521,N_4785);
or U5395 (N_5395,N_4675,N_4737);
nor U5396 (N_5396,N_4690,N_4694);
and U5397 (N_5397,N_5186,N_4914);
nand U5398 (N_5398,N_4973,N_5008);
xor U5399 (N_5399,N_4828,N_4858);
and U5400 (N_5400,N_5131,N_5021);
nand U5401 (N_5401,N_4783,N_4634);
nor U5402 (N_5402,N_4632,N_5047);
and U5403 (N_5403,N_5028,N_4927);
nor U5404 (N_5404,N_4779,N_4769);
or U5405 (N_5405,N_5023,N_4639);
or U5406 (N_5406,N_4577,N_4718);
nand U5407 (N_5407,N_4703,N_4966);
or U5408 (N_5408,N_4862,N_4840);
or U5409 (N_5409,N_4583,N_4753);
and U5410 (N_5410,N_4892,N_5234);
and U5411 (N_5411,N_4571,N_4662);
and U5412 (N_5412,N_4886,N_4971);
and U5413 (N_5413,N_4725,N_4777);
xnor U5414 (N_5414,N_4841,N_5157);
nor U5415 (N_5415,N_5141,N_4942);
nand U5416 (N_5416,N_4541,N_5082);
or U5417 (N_5417,N_4601,N_4898);
and U5418 (N_5418,N_4929,N_4876);
nand U5419 (N_5419,N_4502,N_4911);
and U5420 (N_5420,N_4807,N_4931);
and U5421 (N_5421,N_5243,N_4663);
and U5422 (N_5422,N_5164,N_5208);
xnor U5423 (N_5423,N_5109,N_4542);
nand U5424 (N_5424,N_4893,N_4887);
and U5425 (N_5425,N_4839,N_4679);
nor U5426 (N_5426,N_5006,N_4894);
or U5427 (N_5427,N_4618,N_5046);
and U5428 (N_5428,N_4820,N_4754);
or U5429 (N_5429,N_4988,N_4993);
nor U5430 (N_5430,N_4799,N_5175);
nand U5431 (N_5431,N_4774,N_5044);
nor U5432 (N_5432,N_4650,N_4701);
xor U5433 (N_5433,N_5128,N_5155);
xnor U5434 (N_5434,N_4693,N_4957);
and U5435 (N_5435,N_5207,N_4830);
and U5436 (N_5436,N_4848,N_4771);
nand U5437 (N_5437,N_5217,N_4917);
and U5438 (N_5438,N_4998,N_4882);
nor U5439 (N_5439,N_4786,N_4748);
or U5440 (N_5440,N_4854,N_5185);
xor U5441 (N_5441,N_4868,N_4522);
and U5442 (N_5442,N_4747,N_5012);
nor U5443 (N_5443,N_4599,N_5055);
or U5444 (N_5444,N_4818,N_4595);
nor U5445 (N_5445,N_4933,N_5030);
and U5446 (N_5446,N_5078,N_4506);
nor U5447 (N_5447,N_5246,N_4940);
or U5448 (N_5448,N_4598,N_4551);
and U5449 (N_5449,N_4846,N_4883);
nand U5450 (N_5450,N_5060,N_4897);
and U5451 (N_5451,N_4844,N_5103);
nor U5452 (N_5452,N_4908,N_4568);
nor U5453 (N_5453,N_4614,N_5038);
nor U5454 (N_5454,N_4644,N_5092);
nand U5455 (N_5455,N_5068,N_4548);
nor U5456 (N_5456,N_5178,N_4762);
or U5457 (N_5457,N_5052,N_4575);
and U5458 (N_5458,N_4645,N_4852);
and U5459 (N_5459,N_5076,N_5204);
nand U5460 (N_5460,N_4728,N_4670);
nor U5461 (N_5461,N_4939,N_4591);
nor U5462 (N_5462,N_4686,N_4588);
nor U5463 (N_5463,N_5214,N_4849);
nor U5464 (N_5464,N_4719,N_4924);
and U5465 (N_5465,N_4683,N_4889);
and U5466 (N_5466,N_5039,N_4543);
xor U5467 (N_5467,N_5048,N_5077);
nor U5468 (N_5468,N_5184,N_4546);
and U5469 (N_5469,N_5163,N_4812);
and U5470 (N_5470,N_4901,N_5007);
nor U5471 (N_5471,N_5065,N_4586);
nand U5472 (N_5472,N_4961,N_4822);
or U5473 (N_5473,N_4723,N_4680);
and U5474 (N_5474,N_5197,N_4837);
nor U5475 (N_5475,N_4573,N_4964);
nor U5476 (N_5476,N_4622,N_5199);
nor U5477 (N_5477,N_4836,N_5144);
nor U5478 (N_5478,N_5085,N_4946);
nor U5479 (N_5479,N_4537,N_4756);
or U5480 (N_5480,N_4554,N_4827);
nand U5481 (N_5481,N_4880,N_4606);
nor U5482 (N_5482,N_4553,N_5212);
nand U5483 (N_5483,N_4646,N_4764);
nor U5484 (N_5484,N_4903,N_5001);
and U5485 (N_5485,N_4944,N_4743);
xnor U5486 (N_5486,N_5004,N_4891);
nand U5487 (N_5487,N_5126,N_4758);
nor U5488 (N_5488,N_5080,N_4556);
nor U5489 (N_5489,N_4750,N_4547);
nand U5490 (N_5490,N_4530,N_4605);
nand U5491 (N_5491,N_4948,N_4608);
nor U5492 (N_5492,N_4631,N_5042);
nor U5493 (N_5493,N_4904,N_4711);
or U5494 (N_5494,N_5083,N_4518);
and U5495 (N_5495,N_5031,N_4544);
nor U5496 (N_5496,N_4825,N_5037);
or U5497 (N_5497,N_4768,N_4519);
or U5498 (N_5498,N_4653,N_4906);
nor U5499 (N_5499,N_5095,N_5194);
and U5500 (N_5500,N_4603,N_4654);
nand U5501 (N_5501,N_5084,N_5168);
nor U5502 (N_5502,N_5029,N_4926);
nor U5503 (N_5503,N_5054,N_4752);
or U5504 (N_5504,N_4742,N_5074);
nand U5505 (N_5505,N_4517,N_4985);
nand U5506 (N_5506,N_4668,N_4667);
nor U5507 (N_5507,N_5040,N_4566);
nor U5508 (N_5508,N_5211,N_4689);
and U5509 (N_5509,N_4943,N_4751);
nand U5510 (N_5510,N_4958,N_5079);
nand U5511 (N_5511,N_4636,N_4627);
nand U5512 (N_5512,N_5133,N_4787);
nor U5513 (N_5513,N_4967,N_4731);
or U5514 (N_5514,N_4788,N_5209);
or U5515 (N_5515,N_4997,N_5136);
nor U5516 (N_5516,N_4691,N_4567);
nand U5517 (N_5517,N_4726,N_4673);
or U5518 (N_5518,N_4624,N_4505);
or U5519 (N_5519,N_4512,N_5033);
nor U5520 (N_5520,N_5098,N_5064);
nor U5521 (N_5521,N_4952,N_5108);
nor U5522 (N_5522,N_4870,N_4907);
nor U5523 (N_5523,N_4843,N_5034);
or U5524 (N_5524,N_5202,N_4621);
nand U5525 (N_5525,N_4504,N_5248);
nand U5526 (N_5526,N_4928,N_5062);
nand U5527 (N_5527,N_4778,N_4649);
nand U5528 (N_5528,N_5173,N_4526);
nor U5529 (N_5529,N_4558,N_5058);
and U5530 (N_5530,N_5072,N_4633);
or U5531 (N_5531,N_4759,N_4796);
xnor U5532 (N_5532,N_4915,N_4707);
xnor U5533 (N_5533,N_4938,N_4919);
nand U5534 (N_5534,N_4659,N_4941);
and U5535 (N_5535,N_4741,N_4565);
nand U5536 (N_5536,N_4536,N_4913);
or U5537 (N_5537,N_4706,N_4834);
and U5538 (N_5538,N_4813,N_5127);
or U5539 (N_5539,N_4677,N_4696);
and U5540 (N_5540,N_5019,N_4515);
or U5541 (N_5541,N_4814,N_4896);
or U5542 (N_5542,N_5099,N_4916);
or U5543 (N_5543,N_4801,N_5220);
nor U5544 (N_5544,N_4795,N_5237);
nor U5545 (N_5545,N_5053,N_4619);
or U5546 (N_5546,N_5018,N_4755);
nand U5547 (N_5547,N_5122,N_4625);
and U5548 (N_5548,N_5170,N_4923);
or U5549 (N_5549,N_4574,N_5143);
and U5550 (N_5550,N_5014,N_4579);
nor U5551 (N_5551,N_4859,N_4665);
and U5552 (N_5552,N_5200,N_5088);
nand U5553 (N_5553,N_4527,N_4676);
or U5554 (N_5554,N_4838,N_4782);
nand U5555 (N_5555,N_5123,N_4738);
nand U5556 (N_5556,N_4569,N_4529);
nor U5557 (N_5557,N_5032,N_4809);
and U5558 (N_5558,N_4623,N_4648);
nand U5559 (N_5559,N_4660,N_4699);
and U5560 (N_5560,N_4510,N_4712);
or U5561 (N_5561,N_5087,N_4585);
nand U5562 (N_5562,N_4932,N_4647);
and U5563 (N_5563,N_4678,N_5010);
or U5564 (N_5564,N_4962,N_5148);
nand U5565 (N_5565,N_4638,N_4767);
nor U5566 (N_5566,N_4584,N_4865);
and U5567 (N_5567,N_4864,N_4922);
nor U5568 (N_5568,N_4637,N_4963);
nor U5569 (N_5569,N_5093,N_5005);
xor U5570 (N_5570,N_4628,N_5210);
nor U5571 (N_5571,N_4808,N_4763);
nand U5572 (N_5572,N_4523,N_4821);
or U5573 (N_5573,N_5132,N_4589);
or U5574 (N_5574,N_4730,N_5067);
nand U5575 (N_5575,N_4989,N_5213);
or U5576 (N_5576,N_5075,N_4793);
or U5577 (N_5577,N_5130,N_4879);
or U5578 (N_5578,N_5113,N_4642);
nand U5579 (N_5579,N_5118,N_4704);
or U5580 (N_5580,N_5238,N_5106);
and U5581 (N_5581,N_5193,N_4576);
nor U5582 (N_5582,N_4905,N_4776);
and U5583 (N_5583,N_5049,N_4761);
nand U5584 (N_5584,N_4937,N_4949);
xnor U5585 (N_5585,N_5156,N_4533);
or U5586 (N_5586,N_4513,N_5167);
nand U5587 (N_5587,N_4977,N_4611);
nand U5588 (N_5588,N_5043,N_4552);
and U5589 (N_5589,N_4885,N_4713);
nand U5590 (N_5590,N_4700,N_5059);
or U5591 (N_5591,N_5009,N_4902);
xor U5592 (N_5592,N_4867,N_4871);
nor U5593 (N_5593,N_4804,N_4766);
nand U5594 (N_5594,N_4562,N_4550);
nand U5595 (N_5595,N_4559,N_5188);
and U5596 (N_5596,N_4698,N_5057);
or U5597 (N_5597,N_4560,N_5071);
and U5598 (N_5598,N_4872,N_5206);
nand U5599 (N_5599,N_4635,N_4999);
nand U5600 (N_5600,N_4781,N_4935);
and U5601 (N_5601,N_5179,N_4721);
nand U5602 (N_5602,N_5036,N_4666);
xor U5603 (N_5603,N_4535,N_4643);
nor U5604 (N_5604,N_4869,N_4593);
and U5605 (N_5605,N_4716,N_4705);
nor U5606 (N_5606,N_4757,N_4899);
nor U5607 (N_5607,N_4524,N_4792);
nand U5608 (N_5608,N_4581,N_5249);
nand U5609 (N_5609,N_4540,N_5227);
and U5610 (N_5610,N_4596,N_5017);
and U5611 (N_5611,N_4610,N_4609);
xnor U5612 (N_5612,N_5154,N_4508);
nor U5613 (N_5613,N_5114,N_5196);
or U5614 (N_5614,N_5089,N_4797);
and U5615 (N_5615,N_4770,N_5107);
nand U5616 (N_5616,N_5198,N_5016);
nand U5617 (N_5617,N_5169,N_5152);
xnor U5618 (N_5618,N_4572,N_5150);
nor U5619 (N_5619,N_5081,N_4555);
xor U5620 (N_5620,N_4538,N_5051);
and U5621 (N_5621,N_4594,N_5165);
nand U5622 (N_5622,N_5226,N_5035);
nor U5623 (N_5623,N_4910,N_4981);
nand U5624 (N_5624,N_4815,N_4557);
and U5625 (N_5625,N_5086,N_4885);
and U5626 (N_5626,N_4766,N_5064);
or U5627 (N_5627,N_5208,N_4786);
and U5628 (N_5628,N_4695,N_4696);
nand U5629 (N_5629,N_4634,N_4939);
nor U5630 (N_5630,N_4657,N_4572);
nand U5631 (N_5631,N_4776,N_4635);
and U5632 (N_5632,N_4943,N_5005);
nor U5633 (N_5633,N_4956,N_4605);
or U5634 (N_5634,N_5182,N_5092);
and U5635 (N_5635,N_4889,N_4816);
or U5636 (N_5636,N_5249,N_4616);
or U5637 (N_5637,N_4739,N_4815);
xor U5638 (N_5638,N_4618,N_4546);
or U5639 (N_5639,N_5033,N_5082);
nand U5640 (N_5640,N_4778,N_4792);
nand U5641 (N_5641,N_4510,N_5058);
and U5642 (N_5642,N_4926,N_4758);
nor U5643 (N_5643,N_5178,N_4989);
nor U5644 (N_5644,N_4885,N_4909);
nor U5645 (N_5645,N_4774,N_4731);
nand U5646 (N_5646,N_4569,N_5116);
or U5647 (N_5647,N_5142,N_4503);
xnor U5648 (N_5648,N_4659,N_4689);
xor U5649 (N_5649,N_4648,N_4501);
nand U5650 (N_5650,N_5144,N_4798);
and U5651 (N_5651,N_5042,N_5085);
nor U5652 (N_5652,N_4735,N_5127);
and U5653 (N_5653,N_5083,N_5172);
or U5654 (N_5654,N_4844,N_4731);
or U5655 (N_5655,N_4996,N_4654);
or U5656 (N_5656,N_4784,N_4552);
nor U5657 (N_5657,N_5079,N_5195);
nor U5658 (N_5658,N_4810,N_5095);
and U5659 (N_5659,N_4814,N_5233);
nand U5660 (N_5660,N_5140,N_5205);
or U5661 (N_5661,N_5101,N_5211);
nand U5662 (N_5662,N_4573,N_4601);
nand U5663 (N_5663,N_4683,N_4598);
nor U5664 (N_5664,N_4948,N_4602);
and U5665 (N_5665,N_4831,N_4580);
and U5666 (N_5666,N_4928,N_4955);
and U5667 (N_5667,N_4831,N_5245);
xor U5668 (N_5668,N_5065,N_5005);
and U5669 (N_5669,N_5022,N_4565);
xor U5670 (N_5670,N_5036,N_5062);
or U5671 (N_5671,N_5011,N_4940);
and U5672 (N_5672,N_4831,N_4651);
nand U5673 (N_5673,N_4739,N_4773);
nor U5674 (N_5674,N_4664,N_5175);
nand U5675 (N_5675,N_4651,N_4662);
and U5676 (N_5676,N_5196,N_5202);
nor U5677 (N_5677,N_5103,N_5151);
nor U5678 (N_5678,N_5173,N_4675);
nor U5679 (N_5679,N_4669,N_4998);
and U5680 (N_5680,N_5248,N_4685);
or U5681 (N_5681,N_4501,N_4608);
nor U5682 (N_5682,N_4922,N_5042);
or U5683 (N_5683,N_5240,N_5236);
and U5684 (N_5684,N_4606,N_5021);
and U5685 (N_5685,N_4928,N_5169);
and U5686 (N_5686,N_4751,N_5131);
or U5687 (N_5687,N_4539,N_4759);
and U5688 (N_5688,N_4622,N_5247);
nand U5689 (N_5689,N_4607,N_5192);
or U5690 (N_5690,N_5061,N_4673);
nand U5691 (N_5691,N_4675,N_4838);
xnor U5692 (N_5692,N_4928,N_4855);
nand U5693 (N_5693,N_5030,N_4963);
xor U5694 (N_5694,N_4747,N_5043);
xor U5695 (N_5695,N_5081,N_5168);
nand U5696 (N_5696,N_4742,N_4620);
xor U5697 (N_5697,N_5106,N_5154);
nand U5698 (N_5698,N_4753,N_4696);
or U5699 (N_5699,N_4992,N_4728);
nor U5700 (N_5700,N_4700,N_4889);
and U5701 (N_5701,N_4892,N_4675);
nor U5702 (N_5702,N_4654,N_4823);
and U5703 (N_5703,N_4698,N_4555);
nand U5704 (N_5704,N_4698,N_5196);
nor U5705 (N_5705,N_5107,N_4863);
or U5706 (N_5706,N_4998,N_4880);
nand U5707 (N_5707,N_4645,N_4778);
xnor U5708 (N_5708,N_4669,N_5097);
and U5709 (N_5709,N_4947,N_5103);
or U5710 (N_5710,N_5094,N_4638);
and U5711 (N_5711,N_5030,N_4971);
nand U5712 (N_5712,N_4641,N_4864);
xor U5713 (N_5713,N_5212,N_4952);
xnor U5714 (N_5714,N_5111,N_4864);
nand U5715 (N_5715,N_4825,N_5203);
and U5716 (N_5716,N_4652,N_4589);
nand U5717 (N_5717,N_4646,N_5136);
nor U5718 (N_5718,N_5144,N_4978);
and U5719 (N_5719,N_4548,N_5124);
xnor U5720 (N_5720,N_5176,N_5133);
and U5721 (N_5721,N_4649,N_5200);
nor U5722 (N_5722,N_5227,N_5244);
or U5723 (N_5723,N_4745,N_4693);
nand U5724 (N_5724,N_5126,N_5113);
nor U5725 (N_5725,N_4749,N_4784);
and U5726 (N_5726,N_4701,N_5150);
and U5727 (N_5727,N_4876,N_4741);
nor U5728 (N_5728,N_4769,N_5016);
and U5729 (N_5729,N_4774,N_4644);
or U5730 (N_5730,N_4583,N_4908);
and U5731 (N_5731,N_5003,N_5175);
nor U5732 (N_5732,N_4983,N_4822);
or U5733 (N_5733,N_5217,N_5043);
or U5734 (N_5734,N_4822,N_4967);
and U5735 (N_5735,N_5233,N_4638);
nor U5736 (N_5736,N_4804,N_4957);
or U5737 (N_5737,N_5095,N_4606);
or U5738 (N_5738,N_4714,N_5023);
nor U5739 (N_5739,N_4570,N_4516);
nor U5740 (N_5740,N_4600,N_4599);
nand U5741 (N_5741,N_4955,N_4566);
nor U5742 (N_5742,N_4673,N_4770);
and U5743 (N_5743,N_4997,N_4904);
and U5744 (N_5744,N_4782,N_4915);
and U5745 (N_5745,N_4957,N_4985);
nor U5746 (N_5746,N_4813,N_4846);
nand U5747 (N_5747,N_4780,N_5216);
and U5748 (N_5748,N_4883,N_5241);
nand U5749 (N_5749,N_4976,N_4944);
or U5750 (N_5750,N_4976,N_5191);
nand U5751 (N_5751,N_4881,N_4901);
and U5752 (N_5752,N_4605,N_4627);
and U5753 (N_5753,N_5090,N_4741);
nand U5754 (N_5754,N_5061,N_4554);
nor U5755 (N_5755,N_4945,N_5103);
and U5756 (N_5756,N_4795,N_5154);
or U5757 (N_5757,N_4643,N_4648);
and U5758 (N_5758,N_4873,N_4980);
or U5759 (N_5759,N_4600,N_5169);
nor U5760 (N_5760,N_4951,N_5100);
and U5761 (N_5761,N_5243,N_4727);
nor U5762 (N_5762,N_4570,N_5019);
or U5763 (N_5763,N_5050,N_5238);
or U5764 (N_5764,N_4963,N_5210);
or U5765 (N_5765,N_5243,N_5185);
or U5766 (N_5766,N_5032,N_4939);
xor U5767 (N_5767,N_4508,N_4652);
or U5768 (N_5768,N_4682,N_4618);
nor U5769 (N_5769,N_4814,N_4645);
or U5770 (N_5770,N_5025,N_4998);
nand U5771 (N_5771,N_4983,N_5060);
and U5772 (N_5772,N_5088,N_5201);
nor U5773 (N_5773,N_5148,N_5074);
and U5774 (N_5774,N_5093,N_5052);
nand U5775 (N_5775,N_4793,N_5158);
or U5776 (N_5776,N_4681,N_4686);
and U5777 (N_5777,N_4800,N_4868);
or U5778 (N_5778,N_4730,N_5082);
nand U5779 (N_5779,N_5056,N_4940);
xor U5780 (N_5780,N_4580,N_4559);
nand U5781 (N_5781,N_4752,N_4523);
or U5782 (N_5782,N_4693,N_4701);
nand U5783 (N_5783,N_4611,N_4841);
nand U5784 (N_5784,N_5171,N_4982);
or U5785 (N_5785,N_4650,N_5182);
nand U5786 (N_5786,N_4751,N_4681);
nor U5787 (N_5787,N_4695,N_4993);
nor U5788 (N_5788,N_5124,N_4534);
nand U5789 (N_5789,N_5009,N_4654);
nor U5790 (N_5790,N_4801,N_4872);
nor U5791 (N_5791,N_5100,N_4501);
and U5792 (N_5792,N_4713,N_4642);
or U5793 (N_5793,N_5109,N_4758);
nor U5794 (N_5794,N_5006,N_4983);
and U5795 (N_5795,N_4937,N_4884);
and U5796 (N_5796,N_4818,N_4898);
or U5797 (N_5797,N_5154,N_4614);
or U5798 (N_5798,N_4937,N_4655);
or U5799 (N_5799,N_4512,N_5005);
and U5800 (N_5800,N_4604,N_4944);
nor U5801 (N_5801,N_4809,N_5082);
nand U5802 (N_5802,N_4845,N_4952);
or U5803 (N_5803,N_4559,N_4905);
nor U5804 (N_5804,N_5166,N_4647);
nand U5805 (N_5805,N_4711,N_5059);
nand U5806 (N_5806,N_4919,N_4992);
nand U5807 (N_5807,N_4606,N_5240);
and U5808 (N_5808,N_5200,N_5050);
nand U5809 (N_5809,N_4978,N_5062);
nand U5810 (N_5810,N_4584,N_5052);
or U5811 (N_5811,N_4933,N_5189);
xor U5812 (N_5812,N_5203,N_4508);
xor U5813 (N_5813,N_4581,N_4676);
nor U5814 (N_5814,N_4952,N_5057);
xnor U5815 (N_5815,N_4501,N_5101);
nor U5816 (N_5816,N_4817,N_4891);
xor U5817 (N_5817,N_5084,N_4613);
and U5818 (N_5818,N_4855,N_4902);
nand U5819 (N_5819,N_4620,N_4851);
nor U5820 (N_5820,N_4671,N_5236);
nor U5821 (N_5821,N_4676,N_4941);
or U5822 (N_5822,N_5228,N_4981);
or U5823 (N_5823,N_4616,N_5162);
and U5824 (N_5824,N_5096,N_5103);
nor U5825 (N_5825,N_5064,N_4800);
nand U5826 (N_5826,N_4972,N_5106);
nor U5827 (N_5827,N_4875,N_4827);
nor U5828 (N_5828,N_4689,N_4847);
and U5829 (N_5829,N_4611,N_4924);
xnor U5830 (N_5830,N_5018,N_4923);
or U5831 (N_5831,N_4959,N_4966);
and U5832 (N_5832,N_4825,N_4892);
and U5833 (N_5833,N_4807,N_4675);
and U5834 (N_5834,N_4913,N_5147);
nand U5835 (N_5835,N_4695,N_5202);
or U5836 (N_5836,N_4591,N_5140);
and U5837 (N_5837,N_4996,N_5009);
and U5838 (N_5838,N_5229,N_4628);
nand U5839 (N_5839,N_4638,N_5059);
or U5840 (N_5840,N_4814,N_5085);
nand U5841 (N_5841,N_4650,N_5206);
nor U5842 (N_5842,N_4771,N_4923);
or U5843 (N_5843,N_4560,N_4886);
nor U5844 (N_5844,N_4534,N_5211);
nor U5845 (N_5845,N_5216,N_4933);
xor U5846 (N_5846,N_5151,N_4692);
nand U5847 (N_5847,N_4705,N_4754);
and U5848 (N_5848,N_5012,N_4774);
nor U5849 (N_5849,N_5181,N_5137);
nor U5850 (N_5850,N_4664,N_4838);
nand U5851 (N_5851,N_4792,N_4601);
and U5852 (N_5852,N_4916,N_4997);
xnor U5853 (N_5853,N_5154,N_4786);
nor U5854 (N_5854,N_4549,N_4982);
nand U5855 (N_5855,N_5232,N_4921);
nand U5856 (N_5856,N_5068,N_4934);
and U5857 (N_5857,N_4608,N_4968);
xor U5858 (N_5858,N_4950,N_5197);
nor U5859 (N_5859,N_4925,N_4772);
xor U5860 (N_5860,N_4603,N_5044);
xnor U5861 (N_5861,N_5033,N_5044);
nand U5862 (N_5862,N_4755,N_4910);
nand U5863 (N_5863,N_4987,N_4738);
nand U5864 (N_5864,N_5170,N_4735);
xnor U5865 (N_5865,N_4754,N_5116);
nand U5866 (N_5866,N_4918,N_4532);
xor U5867 (N_5867,N_5200,N_4947);
nor U5868 (N_5868,N_4644,N_5070);
or U5869 (N_5869,N_4669,N_5147);
nand U5870 (N_5870,N_5032,N_4619);
and U5871 (N_5871,N_4620,N_4580);
or U5872 (N_5872,N_4588,N_5107);
and U5873 (N_5873,N_4515,N_4736);
or U5874 (N_5874,N_5227,N_4989);
or U5875 (N_5875,N_4578,N_5144);
xnor U5876 (N_5876,N_4543,N_5114);
xor U5877 (N_5877,N_4527,N_4768);
nor U5878 (N_5878,N_4782,N_4787);
xnor U5879 (N_5879,N_4547,N_4760);
nand U5880 (N_5880,N_4632,N_5109);
nor U5881 (N_5881,N_4776,N_5148);
and U5882 (N_5882,N_4934,N_5201);
nor U5883 (N_5883,N_5129,N_5178);
or U5884 (N_5884,N_4630,N_4680);
and U5885 (N_5885,N_4749,N_5072);
or U5886 (N_5886,N_4587,N_5074);
nor U5887 (N_5887,N_4656,N_5166);
and U5888 (N_5888,N_4884,N_4536);
or U5889 (N_5889,N_4803,N_4575);
or U5890 (N_5890,N_4921,N_4719);
xnor U5891 (N_5891,N_4931,N_4989);
and U5892 (N_5892,N_4555,N_4914);
or U5893 (N_5893,N_4686,N_5009);
nor U5894 (N_5894,N_5213,N_4986);
or U5895 (N_5895,N_4738,N_5200);
nand U5896 (N_5896,N_5060,N_5171);
nor U5897 (N_5897,N_4519,N_5036);
nand U5898 (N_5898,N_4681,N_4935);
nand U5899 (N_5899,N_5198,N_4727);
xnor U5900 (N_5900,N_4705,N_5077);
or U5901 (N_5901,N_4641,N_4578);
xor U5902 (N_5902,N_5069,N_5147);
nand U5903 (N_5903,N_5074,N_4680);
and U5904 (N_5904,N_5104,N_4834);
xor U5905 (N_5905,N_4815,N_4913);
and U5906 (N_5906,N_5039,N_4784);
nor U5907 (N_5907,N_4746,N_5095);
nor U5908 (N_5908,N_4613,N_4995);
nand U5909 (N_5909,N_4836,N_4706);
or U5910 (N_5910,N_4946,N_4850);
and U5911 (N_5911,N_4706,N_4845);
xor U5912 (N_5912,N_5155,N_4530);
nor U5913 (N_5913,N_5005,N_4678);
nor U5914 (N_5914,N_4742,N_4524);
or U5915 (N_5915,N_5145,N_5227);
nor U5916 (N_5916,N_5159,N_5149);
nand U5917 (N_5917,N_5243,N_4584);
nor U5918 (N_5918,N_5180,N_5176);
nor U5919 (N_5919,N_4715,N_4933);
nand U5920 (N_5920,N_4522,N_4748);
or U5921 (N_5921,N_4933,N_5196);
or U5922 (N_5922,N_4551,N_4748);
or U5923 (N_5923,N_4912,N_4986);
and U5924 (N_5924,N_4865,N_4998);
or U5925 (N_5925,N_4949,N_4581);
and U5926 (N_5926,N_4848,N_4657);
nand U5927 (N_5927,N_4774,N_4984);
and U5928 (N_5928,N_5184,N_4863);
nand U5929 (N_5929,N_4947,N_4880);
or U5930 (N_5930,N_4808,N_5144);
nor U5931 (N_5931,N_5046,N_5071);
and U5932 (N_5932,N_4512,N_5023);
nand U5933 (N_5933,N_4650,N_4544);
and U5934 (N_5934,N_5196,N_5093);
nand U5935 (N_5935,N_4592,N_4758);
nor U5936 (N_5936,N_4903,N_5234);
xnor U5937 (N_5937,N_4732,N_4513);
nor U5938 (N_5938,N_5246,N_4968);
nand U5939 (N_5939,N_4689,N_5021);
or U5940 (N_5940,N_4865,N_5162);
or U5941 (N_5941,N_5199,N_4745);
and U5942 (N_5942,N_5172,N_5055);
nor U5943 (N_5943,N_4681,N_5059);
nor U5944 (N_5944,N_4546,N_5013);
or U5945 (N_5945,N_4805,N_5160);
or U5946 (N_5946,N_4892,N_4658);
or U5947 (N_5947,N_4682,N_4510);
nand U5948 (N_5948,N_4723,N_4526);
or U5949 (N_5949,N_4688,N_4860);
or U5950 (N_5950,N_4929,N_4850);
nor U5951 (N_5951,N_4871,N_5240);
and U5952 (N_5952,N_4680,N_5142);
nand U5953 (N_5953,N_4619,N_4613);
or U5954 (N_5954,N_4761,N_5182);
nand U5955 (N_5955,N_4838,N_4656);
nor U5956 (N_5956,N_4839,N_4888);
or U5957 (N_5957,N_4617,N_5135);
and U5958 (N_5958,N_4738,N_5112);
nand U5959 (N_5959,N_4551,N_4734);
or U5960 (N_5960,N_5061,N_4602);
or U5961 (N_5961,N_4561,N_5239);
or U5962 (N_5962,N_4535,N_5028);
or U5963 (N_5963,N_4677,N_5107);
or U5964 (N_5964,N_4970,N_5081);
and U5965 (N_5965,N_4755,N_5004);
and U5966 (N_5966,N_4859,N_5181);
xor U5967 (N_5967,N_4775,N_4894);
nor U5968 (N_5968,N_4923,N_4735);
nor U5969 (N_5969,N_4664,N_5157);
nand U5970 (N_5970,N_4509,N_5109);
nand U5971 (N_5971,N_4999,N_5154);
xor U5972 (N_5972,N_5022,N_4842);
and U5973 (N_5973,N_4754,N_4775);
and U5974 (N_5974,N_5157,N_4853);
xnor U5975 (N_5975,N_4770,N_4929);
nor U5976 (N_5976,N_4889,N_5196);
and U5977 (N_5977,N_5180,N_4749);
xnor U5978 (N_5978,N_4813,N_4685);
and U5979 (N_5979,N_5211,N_4510);
nor U5980 (N_5980,N_4681,N_5008);
nor U5981 (N_5981,N_5033,N_4937);
or U5982 (N_5982,N_4702,N_4555);
or U5983 (N_5983,N_5095,N_4556);
or U5984 (N_5984,N_4625,N_4857);
and U5985 (N_5985,N_4675,N_4685);
and U5986 (N_5986,N_4557,N_5057);
and U5987 (N_5987,N_4779,N_4671);
nor U5988 (N_5988,N_4835,N_5052);
nor U5989 (N_5989,N_4897,N_4515);
nor U5990 (N_5990,N_5019,N_4628);
nand U5991 (N_5991,N_4989,N_5187);
or U5992 (N_5992,N_4706,N_4694);
or U5993 (N_5993,N_5097,N_4791);
or U5994 (N_5994,N_5074,N_4981);
nor U5995 (N_5995,N_4945,N_4835);
nand U5996 (N_5996,N_4708,N_5219);
or U5997 (N_5997,N_4924,N_4840);
and U5998 (N_5998,N_4545,N_5235);
or U5999 (N_5999,N_4819,N_4774);
nor U6000 (N_6000,N_5448,N_5361);
and U6001 (N_6001,N_5813,N_5648);
nand U6002 (N_6002,N_5451,N_5996);
nand U6003 (N_6003,N_5659,N_5786);
nor U6004 (N_6004,N_5710,N_5657);
nand U6005 (N_6005,N_5439,N_5663);
or U6006 (N_6006,N_5263,N_5740);
or U6007 (N_6007,N_5409,N_5565);
or U6008 (N_6008,N_5771,N_5310);
nand U6009 (N_6009,N_5745,N_5769);
or U6010 (N_6010,N_5727,N_5681);
xnor U6011 (N_6011,N_5684,N_5729);
nand U6012 (N_6012,N_5765,N_5287);
nand U6013 (N_6013,N_5967,N_5644);
xor U6014 (N_6014,N_5906,N_5955);
and U6015 (N_6015,N_5567,N_5416);
and U6016 (N_6016,N_5751,N_5533);
and U6017 (N_6017,N_5760,N_5469);
nand U6018 (N_6018,N_5337,N_5397);
nor U6019 (N_6019,N_5275,N_5406);
xor U6020 (N_6020,N_5608,N_5991);
or U6021 (N_6021,N_5484,N_5324);
and U6022 (N_6022,N_5258,N_5641);
and U6023 (N_6023,N_5876,N_5251);
or U6024 (N_6024,N_5798,N_5921);
nand U6025 (N_6025,N_5851,N_5800);
and U6026 (N_6026,N_5988,N_5327);
xor U6027 (N_6027,N_5985,N_5370);
nand U6028 (N_6028,N_5815,N_5366);
or U6029 (N_6029,N_5343,N_5650);
or U6030 (N_6030,N_5457,N_5829);
and U6031 (N_6031,N_5444,N_5592);
nor U6032 (N_6032,N_5643,N_5598);
or U6033 (N_6033,N_5852,N_5807);
or U6034 (N_6034,N_5630,N_5652);
xor U6035 (N_6035,N_5423,N_5868);
xnor U6036 (N_6036,N_5999,N_5562);
nand U6037 (N_6037,N_5981,N_5490);
and U6038 (N_6038,N_5520,N_5712);
xnor U6039 (N_6039,N_5892,N_5395);
or U6040 (N_6040,N_5538,N_5739);
and U6041 (N_6041,N_5979,N_5887);
nor U6042 (N_6042,N_5808,N_5855);
and U6043 (N_6043,N_5420,N_5349);
nor U6044 (N_6044,N_5314,N_5552);
or U6045 (N_6045,N_5537,N_5792);
or U6046 (N_6046,N_5722,N_5685);
xnor U6047 (N_6047,N_5894,N_5627);
and U6048 (N_6048,N_5289,N_5637);
and U6049 (N_6049,N_5672,N_5434);
nor U6050 (N_6050,N_5818,N_5619);
nand U6051 (N_6051,N_5534,N_5990);
xnor U6052 (N_6052,N_5462,N_5570);
xor U6053 (N_6053,N_5977,N_5762);
or U6054 (N_6054,N_5827,N_5593);
or U6055 (N_6055,N_5513,N_5880);
nor U6056 (N_6056,N_5297,N_5661);
xor U6057 (N_6057,N_5521,N_5847);
and U6058 (N_6058,N_5628,N_5507);
and U6059 (N_6059,N_5501,N_5526);
and U6060 (N_6060,N_5986,N_5651);
nand U6061 (N_6061,N_5972,N_5445);
nor U6062 (N_6062,N_5335,N_5560);
nand U6063 (N_6063,N_5557,N_5464);
and U6064 (N_6064,N_5857,N_5495);
nor U6065 (N_6065,N_5730,N_5353);
nor U6066 (N_6066,N_5779,N_5781);
or U6067 (N_6067,N_5806,N_5276);
nand U6068 (N_6068,N_5456,N_5290);
nand U6069 (N_6069,N_5614,N_5579);
nand U6070 (N_6070,N_5820,N_5519);
and U6071 (N_6071,N_5753,N_5328);
nand U6072 (N_6072,N_5586,N_5839);
nor U6073 (N_6073,N_5634,N_5767);
xnor U6074 (N_6074,N_5948,N_5359);
and U6075 (N_6075,N_5803,N_5399);
nand U6076 (N_6076,N_5272,N_5891);
and U6077 (N_6077,N_5723,N_5804);
xor U6078 (N_6078,N_5487,N_5429);
nor U6079 (N_6079,N_5437,N_5285);
nand U6080 (N_6080,N_5882,N_5532);
nor U6081 (N_6081,N_5400,N_5941);
nor U6082 (N_6082,N_5318,N_5449);
nand U6083 (N_6083,N_5854,N_5728);
nand U6084 (N_6084,N_5408,N_5884);
or U6085 (N_6085,N_5775,N_5711);
or U6086 (N_6086,N_5580,N_5367);
nand U6087 (N_6087,N_5571,N_5927);
nor U6088 (N_6088,N_5871,N_5415);
nand U6089 (N_6089,N_5840,N_5475);
nor U6090 (N_6090,N_5597,N_5755);
or U6091 (N_6091,N_5334,N_5443);
nor U6092 (N_6092,N_5794,N_5333);
and U6093 (N_6093,N_5486,N_5364);
and U6094 (N_6094,N_5446,N_5960);
xnor U6095 (N_6095,N_5515,N_5543);
xnor U6096 (N_6096,N_5547,N_5474);
nor U6097 (N_6097,N_5340,N_5363);
nand U6098 (N_6098,N_5494,N_5938);
nor U6099 (N_6099,N_5584,N_5724);
and U6100 (N_6100,N_5461,N_5304);
or U6101 (N_6101,N_5269,N_5431);
and U6102 (N_6102,N_5743,N_5286);
nor U6103 (N_6103,N_5528,N_5971);
and U6104 (N_6104,N_5396,N_5890);
xor U6105 (N_6105,N_5823,N_5780);
or U6106 (N_6106,N_5504,N_5961);
nor U6107 (N_6107,N_5326,N_5572);
nand U6108 (N_6108,N_5609,N_5553);
and U6109 (N_6109,N_5838,N_5670);
nor U6110 (N_6110,N_5508,N_5658);
and U6111 (N_6111,N_5788,N_5413);
or U6112 (N_6112,N_5330,N_5482);
or U6113 (N_6113,N_5789,N_5994);
nand U6114 (N_6114,N_5959,N_5913);
or U6115 (N_6115,N_5554,N_5802);
and U6116 (N_6116,N_5302,N_5678);
and U6117 (N_6117,N_5814,N_5790);
nand U6118 (N_6118,N_5261,N_5380);
nand U6119 (N_6119,N_5911,N_5489);
or U6120 (N_6120,N_5510,N_5902);
nand U6121 (N_6121,N_5516,N_5590);
nor U6122 (N_6122,N_5525,N_5517);
or U6123 (N_6123,N_5308,N_5732);
and U6124 (N_6124,N_5603,N_5773);
nor U6125 (N_6125,N_5425,N_5292);
and U6126 (N_6126,N_5686,N_5713);
nor U6127 (N_6127,N_5316,N_5312);
and U6128 (N_6128,N_5940,N_5784);
nand U6129 (N_6129,N_5345,N_5797);
xnor U6130 (N_6130,N_5618,N_5726);
nand U6131 (N_6131,N_5404,N_5379);
nand U6132 (N_6132,N_5864,N_5688);
nand U6133 (N_6133,N_5331,N_5264);
or U6134 (N_6134,N_5680,N_5358);
nor U6135 (N_6135,N_5509,N_5371);
nand U6136 (N_6136,N_5811,N_5756);
nand U6137 (N_6137,N_5410,N_5271);
nand U6138 (N_6138,N_5842,N_5468);
nand U6139 (N_6139,N_5667,N_5524);
and U6140 (N_6140,N_5717,N_5666);
nor U6141 (N_6141,N_5746,N_5752);
nand U6142 (N_6142,N_5817,N_5772);
and U6143 (N_6143,N_5934,N_5480);
xor U6144 (N_6144,N_5390,N_5859);
xor U6145 (N_6145,N_5821,N_5668);
nand U6146 (N_6146,N_5878,N_5897);
and U6147 (N_6147,N_5964,N_5427);
and U6148 (N_6148,N_5600,N_5500);
and U6149 (N_6149,N_5267,N_5856);
nand U6150 (N_6150,N_5952,N_5435);
nor U6151 (N_6151,N_5671,N_5702);
nor U6152 (N_6152,N_5968,N_5925);
or U6153 (N_6153,N_5796,N_5785);
nand U6154 (N_6154,N_5268,N_5346);
xnor U6155 (N_6155,N_5776,N_5926);
nor U6156 (N_6156,N_5873,N_5622);
or U6157 (N_6157,N_5632,N_5541);
nor U6158 (N_6158,N_5759,N_5280);
xor U6159 (N_6159,N_5253,N_5669);
and U6160 (N_6160,N_5903,N_5578);
nand U6161 (N_6161,N_5675,N_5962);
or U6162 (N_6162,N_5975,N_5270);
nand U6163 (N_6163,N_5283,N_5910);
or U6164 (N_6164,N_5633,N_5354);
nor U6165 (N_6165,N_5260,N_5692);
nor U6166 (N_6166,N_5610,N_5473);
nand U6167 (N_6167,N_5417,N_5942);
or U6168 (N_6168,N_5662,N_5492);
and U6169 (N_6169,N_5398,N_5407);
and U6170 (N_6170,N_5587,N_5376);
and U6171 (N_6171,N_5656,N_5944);
or U6172 (N_6172,N_5881,N_5714);
or U6173 (N_6173,N_5362,N_5946);
xnor U6174 (N_6174,N_5273,N_5992);
nor U6175 (N_6175,N_5378,N_5899);
and U6176 (N_6176,N_5556,N_5505);
xnor U6177 (N_6177,N_5664,N_5947);
nand U6178 (N_6178,N_5418,N_5809);
and U6179 (N_6179,N_5497,N_5577);
nor U6180 (N_6180,N_5889,N_5574);
and U6181 (N_6181,N_5825,N_5617);
nand U6182 (N_6182,N_5496,N_5665);
and U6183 (N_6183,N_5322,N_5843);
xnor U6184 (N_6184,N_5604,N_5357);
or U6185 (N_6185,N_5278,N_5502);
or U6186 (N_6186,N_5734,N_5706);
nor U6187 (N_6187,N_5383,N_5382);
or U6188 (N_6188,N_5514,N_5539);
nand U6189 (N_6189,N_5956,N_5836);
nor U6190 (N_6190,N_5687,N_5984);
or U6191 (N_6191,N_5774,N_5422);
and U6192 (N_6192,N_5682,N_5372);
nand U6193 (N_6193,N_5653,N_5965);
and U6194 (N_6194,N_5388,N_5877);
nor U6195 (N_6195,N_5471,N_5305);
and U6196 (N_6196,N_5830,N_5476);
or U6197 (N_6197,N_5731,N_5615);
nand U6198 (N_6198,N_5858,N_5834);
and U6199 (N_6199,N_5736,N_5438);
or U6200 (N_6200,N_5602,N_5920);
and U6201 (N_6201,N_5315,N_5987);
and U6202 (N_6202,N_5943,N_5875);
nor U6203 (N_6203,N_5924,N_5953);
and U6204 (N_6204,N_5606,N_5850);
nor U6205 (N_6205,N_5581,N_5932);
nor U6206 (N_6206,N_5885,N_5758);
nor U6207 (N_6207,N_5693,N_5266);
or U6208 (N_6208,N_5594,N_5320);
nor U6209 (N_6209,N_5296,N_5566);
nor U6210 (N_6210,N_5442,N_5317);
and U6211 (N_6211,N_5936,N_5582);
xor U6212 (N_6212,N_5323,N_5708);
or U6213 (N_6213,N_5801,N_5735);
and U6214 (N_6214,N_5791,N_5522);
xnor U6215 (N_6215,N_5564,N_5403);
nand U6216 (N_6216,N_5822,N_5389);
or U6217 (N_6217,N_5826,N_5623);
or U6218 (N_6218,N_5368,N_5997);
nand U6219 (N_6219,N_5683,N_5405);
or U6220 (N_6220,N_5607,N_5846);
nand U6221 (N_6221,N_5957,N_5763);
and U6222 (N_6222,N_5392,N_5419);
or U6223 (N_6223,N_5470,N_5893);
or U6224 (N_6224,N_5620,N_5585);
nand U6225 (N_6225,N_5748,N_5568);
and U6226 (N_6226,N_5591,N_5387);
nor U6227 (N_6227,N_5447,N_5540);
nor U6228 (N_6228,N_5835,N_5612);
and U6229 (N_6229,N_5799,N_5983);
or U6230 (N_6230,N_5660,N_5527);
and U6231 (N_6231,N_5795,N_5698);
nand U6232 (N_6232,N_5321,N_5970);
nor U6233 (N_6233,N_5485,N_5605);
nor U6234 (N_6234,N_5848,N_5766);
and U6235 (N_6235,N_5467,N_5428);
and U6236 (N_6236,N_5365,N_5595);
or U6237 (N_6237,N_5674,N_5336);
and U6238 (N_6238,N_5649,N_5279);
nand U6239 (N_6239,N_5872,N_5945);
nand U6240 (N_6240,N_5341,N_5549);
or U6241 (N_6241,N_5309,N_5436);
xor U6242 (N_6242,N_5908,N_5866);
nand U6243 (N_6243,N_5294,N_5655);
and U6244 (N_6244,N_5441,N_5589);
xor U6245 (N_6245,N_5596,N_5274);
xor U6246 (N_6246,N_5518,N_5548);
and U6247 (N_6247,N_5512,N_5503);
nand U6248 (N_6248,N_5647,N_5998);
or U6249 (N_6249,N_5969,N_5454);
nor U6250 (N_6250,N_5394,N_5939);
and U6251 (N_6251,N_5601,N_5298);
nand U6252 (N_6252,N_5426,N_5931);
nor U6253 (N_6253,N_5530,N_5831);
and U6254 (N_6254,N_5546,N_5883);
xor U6255 (N_6255,N_5583,N_5412);
or U6256 (N_6256,N_5332,N_5355);
and U6257 (N_6257,N_5561,N_5531);
nand U6258 (N_6258,N_5465,N_5411);
nand U6259 (N_6259,N_5923,N_5569);
or U6260 (N_6260,N_5707,N_5709);
nor U6261 (N_6261,N_5812,N_5478);
and U6262 (N_6262,N_5989,N_5414);
nor U6263 (N_6263,N_5576,N_5914);
nor U6264 (N_6264,N_5777,N_5282);
or U6265 (N_6265,N_5401,N_5973);
nor U6266 (N_6266,N_5845,N_5374);
or U6267 (N_6267,N_5816,N_5351);
and U6268 (N_6268,N_5654,N_5252);
nor U6269 (N_6269,N_5329,N_5342);
nor U6270 (N_6270,N_5645,N_5339);
and U6271 (N_6271,N_5499,N_5306);
and U6272 (N_6272,N_5313,N_5477);
xnor U6273 (N_6273,N_5385,N_5744);
nand U6274 (N_6274,N_5916,N_5348);
nor U6275 (N_6275,N_5599,N_5262);
nor U6276 (N_6276,N_5624,N_5611);
nand U6277 (N_6277,N_5917,N_5483);
or U6278 (N_6278,N_5935,N_5950);
nand U6279 (N_6279,N_5293,N_5841);
or U6280 (N_6280,N_5481,N_5742);
or U6281 (N_6281,N_5963,N_5421);
nand U6282 (N_6282,N_5819,N_5810);
or U6283 (N_6283,N_5550,N_5958);
nor U6284 (N_6284,N_5928,N_5265);
xnor U6285 (N_6285,N_5311,N_5255);
and U6286 (N_6286,N_5793,N_5951);
and U6287 (N_6287,N_5640,N_5629);
nor U6288 (N_6288,N_5886,N_5974);
nand U6289 (N_6289,N_5621,N_5778);
or U6290 (N_6290,N_5912,N_5511);
and U6291 (N_6291,N_5929,N_5460);
nand U6292 (N_6292,N_5472,N_5690);
nor U6293 (N_6293,N_5749,N_5575);
and U6294 (N_6294,N_5625,N_5277);
or U6295 (N_6295,N_5679,N_5613);
and U6296 (N_6296,N_5631,N_5555);
nand U6297 (N_6297,N_5386,N_5463);
nand U6298 (N_6298,N_5761,N_5874);
nand U6299 (N_6299,N_5704,N_5824);
or U6300 (N_6300,N_5573,N_5733);
and U6301 (N_6301,N_5867,N_5638);
nand U6302 (N_6302,N_5837,N_5291);
nand U6303 (N_6303,N_5558,N_5673);
nand U6304 (N_6304,N_5995,N_5689);
and U6305 (N_6305,N_5901,N_5430);
nor U6306 (N_6306,N_5369,N_5787);
nand U6307 (N_6307,N_5741,N_5720);
and U6308 (N_6308,N_5393,N_5699);
xor U6309 (N_6309,N_5879,N_5782);
or U6310 (N_6310,N_5319,N_5450);
or U6311 (N_6311,N_5738,N_5909);
or U6312 (N_6312,N_5506,N_5853);
nor U6313 (N_6313,N_5360,N_5978);
nand U6314 (N_6314,N_5980,N_5697);
nand U6315 (N_6315,N_5551,N_5966);
nor U6316 (N_6316,N_5373,N_5307);
nand U6317 (N_6317,N_5860,N_5694);
or U6318 (N_6318,N_5863,N_5303);
or U6319 (N_6319,N_5677,N_5545);
xnor U6320 (N_6320,N_5535,N_5256);
nand U6321 (N_6321,N_5300,N_5700);
or U6322 (N_6322,N_5844,N_5350);
nor U6323 (N_6323,N_5933,N_5384);
nand U6324 (N_6324,N_5725,N_5895);
nor U6325 (N_6325,N_5433,N_5288);
nor U6326 (N_6326,N_5301,N_5299);
and U6327 (N_6327,N_5559,N_5750);
nor U6328 (N_6328,N_5452,N_5616);
and U6329 (N_6329,N_5805,N_5783);
xnor U6330 (N_6330,N_5459,N_5754);
and U6331 (N_6331,N_5381,N_5828);
or U6332 (N_6332,N_5356,N_5402);
nand U6333 (N_6333,N_5498,N_5701);
or U6334 (N_6334,N_5695,N_5900);
xnor U6335 (N_6335,N_5455,N_5424);
and U6336 (N_6336,N_5696,N_5375);
and U6337 (N_6337,N_5715,N_5281);
xnor U6338 (N_6338,N_5466,N_5491);
nor U6339 (N_6339,N_5284,N_5544);
nand U6340 (N_6340,N_5479,N_5691);
or U6341 (N_6341,N_5377,N_5898);
and U6342 (N_6342,N_5930,N_5865);
and U6343 (N_6343,N_5703,N_5705);
nor U6344 (N_6344,N_5922,N_5737);
nand U6345 (N_6345,N_5918,N_5523);
and U6346 (N_6346,N_5250,N_5721);
and U6347 (N_6347,N_5904,N_5563);
nor U6348 (N_6348,N_5832,N_5993);
or U6349 (N_6349,N_5536,N_5888);
xnor U6350 (N_6350,N_5639,N_5982);
nand U6351 (N_6351,N_5344,N_5529);
or U6352 (N_6352,N_5768,N_5764);
and U6353 (N_6353,N_5646,N_5849);
xor U6354 (N_6354,N_5642,N_5861);
nand U6355 (N_6355,N_5352,N_5635);
and U6356 (N_6356,N_5719,N_5432);
and U6357 (N_6357,N_5295,N_5954);
and U6358 (N_6358,N_5833,N_5862);
or U6359 (N_6359,N_5347,N_5325);
xnor U6360 (N_6360,N_5949,N_5770);
or U6361 (N_6361,N_5588,N_5869);
nor U6362 (N_6362,N_5338,N_5757);
and U6363 (N_6363,N_5493,N_5542);
and U6364 (N_6364,N_5870,N_5919);
or U6365 (N_6365,N_5636,N_5907);
and U6366 (N_6366,N_5453,N_5488);
or U6367 (N_6367,N_5896,N_5626);
nand U6368 (N_6368,N_5458,N_5915);
and U6369 (N_6369,N_5254,N_5747);
and U6370 (N_6370,N_5976,N_5440);
and U6371 (N_6371,N_5259,N_5391);
xnor U6372 (N_6372,N_5937,N_5718);
nand U6373 (N_6373,N_5905,N_5676);
xnor U6374 (N_6374,N_5257,N_5716);
or U6375 (N_6375,N_5535,N_5610);
and U6376 (N_6376,N_5340,N_5766);
nand U6377 (N_6377,N_5478,N_5954);
and U6378 (N_6378,N_5610,N_5927);
and U6379 (N_6379,N_5619,N_5337);
nand U6380 (N_6380,N_5947,N_5310);
or U6381 (N_6381,N_5682,N_5884);
nor U6382 (N_6382,N_5753,N_5438);
or U6383 (N_6383,N_5888,N_5985);
or U6384 (N_6384,N_5755,N_5972);
or U6385 (N_6385,N_5272,N_5678);
or U6386 (N_6386,N_5270,N_5638);
xor U6387 (N_6387,N_5487,N_5865);
and U6388 (N_6388,N_5589,N_5832);
nand U6389 (N_6389,N_5888,N_5367);
or U6390 (N_6390,N_5925,N_5268);
or U6391 (N_6391,N_5417,N_5834);
xor U6392 (N_6392,N_5575,N_5602);
nor U6393 (N_6393,N_5578,N_5983);
nor U6394 (N_6394,N_5460,N_5250);
nor U6395 (N_6395,N_5319,N_5372);
or U6396 (N_6396,N_5277,N_5377);
or U6397 (N_6397,N_5599,N_5988);
and U6398 (N_6398,N_5456,N_5708);
nor U6399 (N_6399,N_5736,N_5672);
xnor U6400 (N_6400,N_5412,N_5897);
nand U6401 (N_6401,N_5330,N_5296);
and U6402 (N_6402,N_5631,N_5438);
or U6403 (N_6403,N_5285,N_5993);
nand U6404 (N_6404,N_5589,N_5925);
and U6405 (N_6405,N_5917,N_5584);
nor U6406 (N_6406,N_5979,N_5743);
and U6407 (N_6407,N_5902,N_5830);
or U6408 (N_6408,N_5396,N_5668);
or U6409 (N_6409,N_5515,N_5993);
and U6410 (N_6410,N_5631,N_5814);
or U6411 (N_6411,N_5610,N_5588);
or U6412 (N_6412,N_5667,N_5411);
xor U6413 (N_6413,N_5757,N_5284);
or U6414 (N_6414,N_5737,N_5772);
xor U6415 (N_6415,N_5468,N_5252);
nor U6416 (N_6416,N_5828,N_5816);
and U6417 (N_6417,N_5464,N_5697);
nor U6418 (N_6418,N_5937,N_5934);
nor U6419 (N_6419,N_5631,N_5829);
or U6420 (N_6420,N_5813,N_5403);
or U6421 (N_6421,N_5783,N_5598);
nand U6422 (N_6422,N_5913,N_5615);
or U6423 (N_6423,N_5279,N_5531);
nor U6424 (N_6424,N_5987,N_5472);
and U6425 (N_6425,N_5767,N_5366);
nand U6426 (N_6426,N_5691,N_5383);
or U6427 (N_6427,N_5564,N_5623);
and U6428 (N_6428,N_5358,N_5569);
or U6429 (N_6429,N_5640,N_5656);
and U6430 (N_6430,N_5456,N_5294);
nor U6431 (N_6431,N_5351,N_5509);
nand U6432 (N_6432,N_5845,N_5883);
nor U6433 (N_6433,N_5518,N_5507);
and U6434 (N_6434,N_5394,N_5636);
and U6435 (N_6435,N_5733,N_5572);
nand U6436 (N_6436,N_5554,N_5396);
nor U6437 (N_6437,N_5911,N_5972);
nor U6438 (N_6438,N_5723,N_5471);
nand U6439 (N_6439,N_5600,N_5403);
and U6440 (N_6440,N_5796,N_5855);
nand U6441 (N_6441,N_5356,N_5830);
and U6442 (N_6442,N_5703,N_5747);
nand U6443 (N_6443,N_5555,N_5433);
and U6444 (N_6444,N_5736,N_5297);
nand U6445 (N_6445,N_5303,N_5399);
nor U6446 (N_6446,N_5537,N_5694);
or U6447 (N_6447,N_5314,N_5571);
and U6448 (N_6448,N_5970,N_5447);
nor U6449 (N_6449,N_5961,N_5912);
or U6450 (N_6450,N_5729,N_5370);
nand U6451 (N_6451,N_5723,N_5693);
and U6452 (N_6452,N_5642,N_5349);
and U6453 (N_6453,N_5802,N_5881);
nand U6454 (N_6454,N_5620,N_5804);
and U6455 (N_6455,N_5922,N_5539);
or U6456 (N_6456,N_5290,N_5911);
nand U6457 (N_6457,N_5455,N_5753);
or U6458 (N_6458,N_5984,N_5468);
nand U6459 (N_6459,N_5640,N_5917);
nor U6460 (N_6460,N_5459,N_5634);
nor U6461 (N_6461,N_5468,N_5386);
or U6462 (N_6462,N_5502,N_5547);
nand U6463 (N_6463,N_5926,N_5612);
nor U6464 (N_6464,N_5985,N_5811);
nand U6465 (N_6465,N_5770,N_5814);
xor U6466 (N_6466,N_5339,N_5458);
xnor U6467 (N_6467,N_5553,N_5597);
nand U6468 (N_6468,N_5294,N_5732);
xor U6469 (N_6469,N_5455,N_5619);
nor U6470 (N_6470,N_5307,N_5511);
nand U6471 (N_6471,N_5925,N_5591);
and U6472 (N_6472,N_5886,N_5369);
nand U6473 (N_6473,N_5402,N_5665);
or U6474 (N_6474,N_5432,N_5713);
or U6475 (N_6475,N_5328,N_5422);
or U6476 (N_6476,N_5878,N_5674);
and U6477 (N_6477,N_5435,N_5811);
and U6478 (N_6478,N_5346,N_5761);
or U6479 (N_6479,N_5689,N_5625);
or U6480 (N_6480,N_5849,N_5715);
and U6481 (N_6481,N_5540,N_5379);
nand U6482 (N_6482,N_5627,N_5276);
nand U6483 (N_6483,N_5916,N_5722);
or U6484 (N_6484,N_5915,N_5896);
and U6485 (N_6485,N_5515,N_5535);
nand U6486 (N_6486,N_5314,N_5810);
nand U6487 (N_6487,N_5635,N_5296);
and U6488 (N_6488,N_5789,N_5404);
or U6489 (N_6489,N_5452,N_5704);
nor U6490 (N_6490,N_5666,N_5996);
nand U6491 (N_6491,N_5858,N_5357);
xnor U6492 (N_6492,N_5533,N_5346);
nand U6493 (N_6493,N_5593,N_5462);
or U6494 (N_6494,N_5860,N_5796);
nand U6495 (N_6495,N_5993,N_5683);
nor U6496 (N_6496,N_5683,N_5413);
or U6497 (N_6497,N_5615,N_5972);
nor U6498 (N_6498,N_5826,N_5665);
and U6499 (N_6499,N_5840,N_5923);
or U6500 (N_6500,N_5281,N_5497);
and U6501 (N_6501,N_5328,N_5795);
and U6502 (N_6502,N_5750,N_5628);
and U6503 (N_6503,N_5315,N_5403);
and U6504 (N_6504,N_5384,N_5251);
xnor U6505 (N_6505,N_5387,N_5941);
or U6506 (N_6506,N_5256,N_5579);
nor U6507 (N_6507,N_5290,N_5551);
nand U6508 (N_6508,N_5976,N_5284);
nor U6509 (N_6509,N_5390,N_5895);
nand U6510 (N_6510,N_5927,N_5540);
and U6511 (N_6511,N_5267,N_5750);
nand U6512 (N_6512,N_5925,N_5709);
nand U6513 (N_6513,N_5864,N_5334);
nor U6514 (N_6514,N_5409,N_5653);
nand U6515 (N_6515,N_5289,N_5910);
or U6516 (N_6516,N_5476,N_5530);
and U6517 (N_6517,N_5309,N_5431);
and U6518 (N_6518,N_5293,N_5973);
or U6519 (N_6519,N_5936,N_5853);
and U6520 (N_6520,N_5341,N_5696);
or U6521 (N_6521,N_5715,N_5378);
and U6522 (N_6522,N_5854,N_5965);
or U6523 (N_6523,N_5426,N_5995);
xor U6524 (N_6524,N_5592,N_5863);
xnor U6525 (N_6525,N_5993,N_5362);
and U6526 (N_6526,N_5876,N_5991);
nand U6527 (N_6527,N_5757,N_5422);
nor U6528 (N_6528,N_5739,N_5939);
xnor U6529 (N_6529,N_5538,N_5634);
nand U6530 (N_6530,N_5393,N_5496);
or U6531 (N_6531,N_5318,N_5859);
nand U6532 (N_6532,N_5617,N_5852);
nor U6533 (N_6533,N_5805,N_5263);
or U6534 (N_6534,N_5279,N_5893);
nor U6535 (N_6535,N_5584,N_5884);
nand U6536 (N_6536,N_5842,N_5465);
nand U6537 (N_6537,N_5954,N_5272);
nor U6538 (N_6538,N_5839,N_5267);
and U6539 (N_6539,N_5545,N_5724);
nor U6540 (N_6540,N_5526,N_5518);
nand U6541 (N_6541,N_5797,N_5437);
nor U6542 (N_6542,N_5675,N_5830);
or U6543 (N_6543,N_5476,N_5633);
or U6544 (N_6544,N_5294,N_5627);
xnor U6545 (N_6545,N_5741,N_5734);
or U6546 (N_6546,N_5858,N_5657);
nor U6547 (N_6547,N_5580,N_5907);
nand U6548 (N_6548,N_5830,N_5916);
nand U6549 (N_6549,N_5629,N_5604);
nor U6550 (N_6550,N_5379,N_5664);
nand U6551 (N_6551,N_5615,N_5404);
nor U6552 (N_6552,N_5432,N_5584);
nand U6553 (N_6553,N_5758,N_5332);
xnor U6554 (N_6554,N_5334,N_5703);
or U6555 (N_6555,N_5308,N_5698);
and U6556 (N_6556,N_5815,N_5708);
xor U6557 (N_6557,N_5470,N_5590);
nor U6558 (N_6558,N_5875,N_5710);
nor U6559 (N_6559,N_5331,N_5449);
or U6560 (N_6560,N_5770,N_5760);
nor U6561 (N_6561,N_5444,N_5294);
or U6562 (N_6562,N_5510,N_5620);
nand U6563 (N_6563,N_5461,N_5366);
nand U6564 (N_6564,N_5665,N_5706);
or U6565 (N_6565,N_5686,N_5434);
or U6566 (N_6566,N_5876,N_5269);
nor U6567 (N_6567,N_5537,N_5863);
nor U6568 (N_6568,N_5650,N_5366);
nand U6569 (N_6569,N_5287,N_5640);
or U6570 (N_6570,N_5343,N_5576);
or U6571 (N_6571,N_5595,N_5918);
nor U6572 (N_6572,N_5317,N_5815);
nand U6573 (N_6573,N_5295,N_5310);
and U6574 (N_6574,N_5910,N_5542);
nand U6575 (N_6575,N_5840,N_5335);
or U6576 (N_6576,N_5666,N_5967);
nor U6577 (N_6577,N_5596,N_5650);
or U6578 (N_6578,N_5285,N_5482);
or U6579 (N_6579,N_5388,N_5281);
or U6580 (N_6580,N_5428,N_5620);
or U6581 (N_6581,N_5435,N_5663);
and U6582 (N_6582,N_5711,N_5583);
and U6583 (N_6583,N_5968,N_5590);
and U6584 (N_6584,N_5794,N_5497);
xnor U6585 (N_6585,N_5461,N_5280);
nor U6586 (N_6586,N_5740,N_5731);
and U6587 (N_6587,N_5344,N_5897);
or U6588 (N_6588,N_5639,N_5403);
and U6589 (N_6589,N_5666,N_5607);
nor U6590 (N_6590,N_5916,N_5296);
nand U6591 (N_6591,N_5348,N_5345);
and U6592 (N_6592,N_5903,N_5587);
or U6593 (N_6593,N_5680,N_5274);
and U6594 (N_6594,N_5784,N_5954);
and U6595 (N_6595,N_5406,N_5673);
nor U6596 (N_6596,N_5579,N_5943);
nor U6597 (N_6597,N_5569,N_5568);
nand U6598 (N_6598,N_5388,N_5331);
nand U6599 (N_6599,N_5308,N_5574);
nor U6600 (N_6600,N_5336,N_5467);
nor U6601 (N_6601,N_5386,N_5917);
xor U6602 (N_6602,N_5849,N_5547);
and U6603 (N_6603,N_5671,N_5825);
nor U6604 (N_6604,N_5323,N_5627);
nand U6605 (N_6605,N_5608,N_5504);
nor U6606 (N_6606,N_5908,N_5823);
or U6607 (N_6607,N_5863,N_5582);
nor U6608 (N_6608,N_5961,N_5590);
nand U6609 (N_6609,N_5732,N_5745);
nor U6610 (N_6610,N_5575,N_5738);
and U6611 (N_6611,N_5969,N_5939);
nor U6612 (N_6612,N_5709,N_5627);
and U6613 (N_6613,N_5415,N_5614);
and U6614 (N_6614,N_5907,N_5583);
nand U6615 (N_6615,N_5830,N_5746);
nand U6616 (N_6616,N_5583,N_5699);
xor U6617 (N_6617,N_5554,N_5921);
or U6618 (N_6618,N_5809,N_5599);
and U6619 (N_6619,N_5347,N_5546);
nor U6620 (N_6620,N_5561,N_5781);
or U6621 (N_6621,N_5834,N_5583);
xnor U6622 (N_6622,N_5339,N_5495);
xnor U6623 (N_6623,N_5798,N_5953);
or U6624 (N_6624,N_5444,N_5847);
xor U6625 (N_6625,N_5934,N_5583);
and U6626 (N_6626,N_5386,N_5947);
nand U6627 (N_6627,N_5589,N_5852);
xor U6628 (N_6628,N_5288,N_5910);
or U6629 (N_6629,N_5924,N_5346);
nor U6630 (N_6630,N_5842,N_5668);
nor U6631 (N_6631,N_5765,N_5289);
or U6632 (N_6632,N_5588,N_5849);
or U6633 (N_6633,N_5300,N_5844);
or U6634 (N_6634,N_5507,N_5260);
nand U6635 (N_6635,N_5668,N_5495);
and U6636 (N_6636,N_5362,N_5937);
or U6637 (N_6637,N_5271,N_5585);
nor U6638 (N_6638,N_5437,N_5518);
and U6639 (N_6639,N_5437,N_5496);
nor U6640 (N_6640,N_5362,N_5540);
nand U6641 (N_6641,N_5416,N_5694);
nand U6642 (N_6642,N_5756,N_5683);
xor U6643 (N_6643,N_5628,N_5941);
xnor U6644 (N_6644,N_5907,N_5534);
and U6645 (N_6645,N_5957,N_5506);
and U6646 (N_6646,N_5408,N_5685);
nand U6647 (N_6647,N_5625,N_5903);
or U6648 (N_6648,N_5559,N_5912);
nand U6649 (N_6649,N_5451,N_5841);
nor U6650 (N_6650,N_5903,N_5939);
nand U6651 (N_6651,N_5289,N_5341);
nor U6652 (N_6652,N_5371,N_5462);
xnor U6653 (N_6653,N_5766,N_5350);
nand U6654 (N_6654,N_5338,N_5865);
nor U6655 (N_6655,N_5810,N_5305);
and U6656 (N_6656,N_5385,N_5513);
or U6657 (N_6657,N_5272,N_5900);
nor U6658 (N_6658,N_5922,N_5380);
or U6659 (N_6659,N_5329,N_5728);
and U6660 (N_6660,N_5308,N_5787);
and U6661 (N_6661,N_5809,N_5251);
nand U6662 (N_6662,N_5391,N_5385);
nor U6663 (N_6663,N_5952,N_5269);
or U6664 (N_6664,N_5982,N_5531);
and U6665 (N_6665,N_5770,N_5617);
nor U6666 (N_6666,N_5908,N_5555);
and U6667 (N_6667,N_5899,N_5609);
nor U6668 (N_6668,N_5316,N_5996);
and U6669 (N_6669,N_5833,N_5656);
and U6670 (N_6670,N_5751,N_5889);
nand U6671 (N_6671,N_5479,N_5423);
nand U6672 (N_6672,N_5863,N_5844);
or U6673 (N_6673,N_5755,N_5877);
nand U6674 (N_6674,N_5426,N_5724);
nand U6675 (N_6675,N_5951,N_5635);
nor U6676 (N_6676,N_5703,N_5880);
nor U6677 (N_6677,N_5615,N_5350);
or U6678 (N_6678,N_5466,N_5915);
xor U6679 (N_6679,N_5816,N_5979);
nand U6680 (N_6680,N_5748,N_5844);
and U6681 (N_6681,N_5697,N_5515);
nand U6682 (N_6682,N_5769,N_5676);
or U6683 (N_6683,N_5797,N_5837);
nor U6684 (N_6684,N_5326,N_5725);
or U6685 (N_6685,N_5332,N_5653);
nand U6686 (N_6686,N_5280,N_5398);
nand U6687 (N_6687,N_5580,N_5461);
nand U6688 (N_6688,N_5782,N_5913);
nor U6689 (N_6689,N_5924,N_5448);
and U6690 (N_6690,N_5652,N_5890);
and U6691 (N_6691,N_5996,N_5587);
nor U6692 (N_6692,N_5508,N_5779);
and U6693 (N_6693,N_5848,N_5969);
nor U6694 (N_6694,N_5606,N_5995);
and U6695 (N_6695,N_5737,N_5859);
or U6696 (N_6696,N_5950,N_5476);
and U6697 (N_6697,N_5253,N_5980);
xnor U6698 (N_6698,N_5641,N_5691);
nand U6699 (N_6699,N_5393,N_5304);
and U6700 (N_6700,N_5934,N_5275);
and U6701 (N_6701,N_5710,N_5294);
nand U6702 (N_6702,N_5796,N_5583);
xnor U6703 (N_6703,N_5739,N_5620);
or U6704 (N_6704,N_5860,N_5475);
nand U6705 (N_6705,N_5433,N_5702);
nor U6706 (N_6706,N_5467,N_5442);
and U6707 (N_6707,N_5648,N_5947);
nand U6708 (N_6708,N_5496,N_5854);
or U6709 (N_6709,N_5483,N_5798);
and U6710 (N_6710,N_5329,N_5649);
nor U6711 (N_6711,N_5818,N_5895);
or U6712 (N_6712,N_5493,N_5845);
nor U6713 (N_6713,N_5530,N_5298);
or U6714 (N_6714,N_5893,N_5463);
nor U6715 (N_6715,N_5585,N_5536);
nand U6716 (N_6716,N_5561,N_5894);
nand U6717 (N_6717,N_5891,N_5791);
nand U6718 (N_6718,N_5714,N_5679);
nor U6719 (N_6719,N_5417,N_5275);
nor U6720 (N_6720,N_5843,N_5330);
nand U6721 (N_6721,N_5325,N_5659);
xor U6722 (N_6722,N_5648,N_5975);
or U6723 (N_6723,N_5818,N_5366);
nor U6724 (N_6724,N_5907,N_5856);
nand U6725 (N_6725,N_5566,N_5647);
nor U6726 (N_6726,N_5453,N_5348);
nand U6727 (N_6727,N_5767,N_5355);
or U6728 (N_6728,N_5250,N_5684);
and U6729 (N_6729,N_5717,N_5737);
or U6730 (N_6730,N_5379,N_5353);
nand U6731 (N_6731,N_5523,N_5898);
or U6732 (N_6732,N_5498,N_5937);
xor U6733 (N_6733,N_5289,N_5350);
xnor U6734 (N_6734,N_5986,N_5325);
nor U6735 (N_6735,N_5887,N_5512);
nor U6736 (N_6736,N_5924,N_5728);
nor U6737 (N_6737,N_5298,N_5704);
nand U6738 (N_6738,N_5578,N_5441);
xnor U6739 (N_6739,N_5274,N_5351);
nor U6740 (N_6740,N_5994,N_5764);
nor U6741 (N_6741,N_5528,N_5543);
and U6742 (N_6742,N_5852,N_5933);
nand U6743 (N_6743,N_5340,N_5359);
nand U6744 (N_6744,N_5279,N_5930);
nor U6745 (N_6745,N_5838,N_5540);
nor U6746 (N_6746,N_5947,N_5555);
and U6747 (N_6747,N_5826,N_5744);
xor U6748 (N_6748,N_5478,N_5523);
xor U6749 (N_6749,N_5994,N_5767);
nand U6750 (N_6750,N_6354,N_6508);
nand U6751 (N_6751,N_6233,N_6637);
nand U6752 (N_6752,N_6633,N_6662);
or U6753 (N_6753,N_6591,N_6568);
nand U6754 (N_6754,N_6024,N_6313);
or U6755 (N_6755,N_6713,N_6470);
or U6756 (N_6756,N_6415,N_6264);
or U6757 (N_6757,N_6562,N_6465);
and U6758 (N_6758,N_6600,N_6551);
and U6759 (N_6759,N_6521,N_6715);
nor U6760 (N_6760,N_6188,N_6114);
and U6761 (N_6761,N_6646,N_6458);
nand U6762 (N_6762,N_6126,N_6216);
nor U6763 (N_6763,N_6681,N_6084);
nand U6764 (N_6764,N_6003,N_6747);
and U6765 (N_6765,N_6655,N_6207);
nand U6766 (N_6766,N_6648,N_6694);
xor U6767 (N_6767,N_6168,N_6328);
nor U6768 (N_6768,N_6193,N_6395);
or U6769 (N_6769,N_6279,N_6263);
and U6770 (N_6770,N_6295,N_6402);
and U6771 (N_6771,N_6705,N_6134);
or U6772 (N_6772,N_6350,N_6135);
and U6773 (N_6773,N_6391,N_6092);
nand U6774 (N_6774,N_6399,N_6019);
nor U6775 (N_6775,N_6013,N_6348);
nand U6776 (N_6776,N_6556,N_6507);
or U6777 (N_6777,N_6192,N_6589);
nor U6778 (N_6778,N_6386,N_6246);
and U6779 (N_6779,N_6308,N_6298);
nor U6780 (N_6780,N_6383,N_6492);
nand U6781 (N_6781,N_6529,N_6702);
and U6782 (N_6782,N_6017,N_6374);
or U6783 (N_6783,N_6527,N_6157);
nand U6784 (N_6784,N_6208,N_6620);
nand U6785 (N_6785,N_6360,N_6359);
or U6786 (N_6786,N_6397,N_6689);
or U6787 (N_6787,N_6707,N_6483);
nor U6788 (N_6788,N_6209,N_6164);
and U6789 (N_6789,N_6479,N_6115);
and U6790 (N_6790,N_6627,N_6594);
nor U6791 (N_6791,N_6212,N_6364);
nor U6792 (N_6792,N_6503,N_6042);
nor U6793 (N_6793,N_6730,N_6645);
and U6794 (N_6794,N_6224,N_6160);
nor U6795 (N_6795,N_6007,N_6446);
or U6796 (N_6796,N_6119,N_6581);
nand U6797 (N_6797,N_6588,N_6317);
or U6798 (N_6798,N_6526,N_6053);
nand U6799 (N_6799,N_6252,N_6016);
nand U6800 (N_6800,N_6618,N_6131);
and U6801 (N_6801,N_6002,N_6210);
xor U6802 (N_6802,N_6250,N_6525);
nand U6803 (N_6803,N_6401,N_6741);
nor U6804 (N_6804,N_6675,N_6404);
or U6805 (N_6805,N_6190,N_6251);
nor U6806 (N_6806,N_6276,N_6143);
nand U6807 (N_6807,N_6309,N_6561);
and U6808 (N_6808,N_6486,N_6221);
nand U6809 (N_6809,N_6191,N_6304);
and U6810 (N_6810,N_6596,N_6129);
or U6811 (N_6811,N_6287,N_6378);
or U6812 (N_6812,N_6472,N_6669);
nand U6813 (N_6813,N_6547,N_6540);
or U6814 (N_6814,N_6621,N_6430);
nor U6815 (N_6815,N_6686,N_6611);
or U6816 (N_6816,N_6709,N_6578);
and U6817 (N_6817,N_6368,N_6502);
and U6818 (N_6818,N_6375,N_6083);
nand U6819 (N_6819,N_6613,N_6008);
nand U6820 (N_6820,N_6184,N_6334);
nor U6821 (N_6821,N_6055,N_6481);
and U6822 (N_6822,N_6161,N_6282);
and U6823 (N_6823,N_6117,N_6006);
nor U6824 (N_6824,N_6087,N_6047);
or U6825 (N_6825,N_6325,N_6239);
nand U6826 (N_6826,N_6431,N_6189);
and U6827 (N_6827,N_6429,N_6450);
nand U6828 (N_6828,N_6376,N_6103);
or U6829 (N_6829,N_6064,N_6518);
nand U6830 (N_6830,N_6292,N_6330);
or U6831 (N_6831,N_6372,N_6660);
and U6832 (N_6832,N_6629,N_6068);
nor U6833 (N_6833,N_6125,N_6543);
and U6834 (N_6834,N_6601,N_6605);
and U6835 (N_6835,N_6559,N_6583);
and U6836 (N_6836,N_6738,N_6177);
nor U6837 (N_6837,N_6365,N_6461);
nor U6838 (N_6838,N_6632,N_6370);
or U6839 (N_6839,N_6418,N_6541);
xor U6840 (N_6840,N_6028,N_6333);
nor U6841 (N_6841,N_6471,N_6687);
nor U6842 (N_6842,N_6736,N_6244);
or U6843 (N_6843,N_6570,N_6535);
or U6844 (N_6844,N_6265,N_6548);
nor U6845 (N_6845,N_6155,N_6424);
nand U6846 (N_6846,N_6555,N_6717);
nand U6847 (N_6847,N_6312,N_6513);
nand U6848 (N_6848,N_6666,N_6392);
and U6849 (N_6849,N_6178,N_6703);
or U6850 (N_6850,N_6284,N_6080);
xor U6851 (N_6851,N_6145,N_6255);
xnor U6852 (N_6852,N_6170,N_6104);
nor U6853 (N_6853,N_6054,N_6094);
and U6854 (N_6854,N_6058,N_6343);
nand U6855 (N_6855,N_6511,N_6671);
or U6856 (N_6856,N_6035,N_6664);
or U6857 (N_6857,N_6065,N_6480);
and U6858 (N_6858,N_6070,N_6537);
xor U6859 (N_6859,N_6678,N_6152);
nor U6860 (N_6860,N_6714,N_6565);
nand U6861 (N_6861,N_6652,N_6531);
or U6862 (N_6862,N_6195,N_6725);
xnor U6863 (N_6863,N_6194,N_6358);
nor U6864 (N_6864,N_6593,N_6416);
xor U6865 (N_6865,N_6090,N_6744);
or U6866 (N_6866,N_6642,N_6238);
and U6867 (N_6867,N_6014,N_6258);
and U6868 (N_6868,N_6100,N_6202);
xnor U6869 (N_6869,N_6504,N_6271);
nand U6870 (N_6870,N_6356,N_6569);
nand U6871 (N_6871,N_6528,N_6732);
xnor U6872 (N_6872,N_6329,N_6641);
or U6873 (N_6873,N_6663,N_6388);
or U6874 (N_6874,N_6259,N_6727);
and U6875 (N_6875,N_6366,N_6726);
or U6876 (N_6876,N_6022,N_6708);
and U6877 (N_6877,N_6417,N_6020);
nand U6878 (N_6878,N_6640,N_6563);
and U6879 (N_6879,N_6522,N_6237);
or U6880 (N_6880,N_6724,N_6575);
nor U6881 (N_6881,N_6112,N_6536);
nor U6882 (N_6882,N_6558,N_6576);
xor U6883 (N_6883,N_6186,N_6434);
nand U6884 (N_6884,N_6398,N_6082);
and U6885 (N_6885,N_6610,N_6567);
or U6886 (N_6886,N_6665,N_6027);
or U6887 (N_6887,N_6696,N_6327);
nor U6888 (N_6888,N_6475,N_6373);
or U6889 (N_6889,N_6236,N_6420);
nor U6890 (N_6890,N_6101,N_6049);
nand U6891 (N_6891,N_6682,N_6712);
nor U6892 (N_6892,N_6181,N_6249);
and U6893 (N_6893,N_6441,N_6426);
or U6894 (N_6894,N_6196,N_6023);
and U6895 (N_6895,N_6319,N_6464);
nand U6896 (N_6896,N_6288,N_6369);
nor U6897 (N_6897,N_6011,N_6009);
and U6898 (N_6898,N_6274,N_6089);
or U6899 (N_6899,N_6113,N_6407);
or U6900 (N_6900,N_6381,N_6198);
and U6901 (N_6901,N_6139,N_6220);
nand U6902 (N_6902,N_6384,N_6661);
or U6903 (N_6903,N_6311,N_6728);
or U6904 (N_6904,N_6506,N_6411);
or U6905 (N_6905,N_6338,N_6056);
nor U6906 (N_6906,N_6602,N_6116);
nand U6907 (N_6907,N_6467,N_6076);
nor U6908 (N_6908,N_6590,N_6377);
nand U6909 (N_6909,N_6452,N_6061);
nand U6910 (N_6910,N_6608,N_6297);
or U6911 (N_6911,N_6294,N_6063);
nand U6912 (N_6912,N_6273,N_6240);
xnor U6913 (N_6913,N_6459,N_6435);
or U6914 (N_6914,N_6021,N_6519);
xnor U6915 (N_6915,N_6739,N_6630);
and U6916 (N_6916,N_6137,N_6187);
or U6917 (N_6917,N_6408,N_6302);
or U6918 (N_6918,N_6214,N_6501);
nor U6919 (N_6919,N_6124,N_6166);
nand U6920 (N_6920,N_6173,N_6720);
or U6921 (N_6921,N_6073,N_6695);
nand U6922 (N_6922,N_6731,N_6444);
nor U6923 (N_6923,N_6544,N_6676);
nor U6924 (N_6924,N_6440,N_6336);
nand U6925 (N_6925,N_6428,N_6253);
nand U6926 (N_6926,N_6644,N_6599);
or U6927 (N_6927,N_6109,N_6482);
nand U6928 (N_6928,N_6159,N_6005);
or U6929 (N_6929,N_6289,N_6619);
or U6930 (N_6930,N_6066,N_6406);
nand U6931 (N_6931,N_6534,N_6110);
and U6932 (N_6932,N_6422,N_6683);
nand U6933 (N_6933,N_6303,N_6427);
and U6934 (N_6934,N_6026,N_6517);
or U6935 (N_6935,N_6150,N_6491);
nor U6936 (N_6936,N_6339,N_6140);
or U6937 (N_6937,N_6476,N_6051);
nor U6938 (N_6938,N_6211,N_6704);
and U6939 (N_6939,N_6332,N_6275);
xnor U6940 (N_6940,N_6658,N_6097);
nand U6941 (N_6941,N_6495,N_6261);
nand U6942 (N_6942,N_6001,N_6463);
nor U6943 (N_6943,N_6291,N_6650);
nor U6944 (N_6944,N_6579,N_6489);
nor U6945 (N_6945,N_6743,N_6585);
xor U6946 (N_6946,N_6012,N_6423);
nor U6947 (N_6947,N_6635,N_6105);
and U6948 (N_6948,N_6315,N_6039);
nand U6949 (N_6949,N_6046,N_6432);
or U6950 (N_6950,N_6015,N_6691);
or U6951 (N_6951,N_6574,N_6283);
and U6952 (N_6952,N_6509,N_6118);
nand U6953 (N_6953,N_6552,N_6234);
or U6954 (N_6954,N_6530,N_6631);
and U6955 (N_6955,N_6523,N_6301);
and U6956 (N_6956,N_6074,N_6560);
or U6957 (N_6957,N_6380,N_6342);
nor U6958 (N_6958,N_6512,N_6043);
or U6959 (N_6959,N_6546,N_6050);
and U6960 (N_6960,N_6612,N_6349);
and U6961 (N_6961,N_6353,N_6673);
and U6962 (N_6962,N_6004,N_6499);
and U6963 (N_6963,N_6414,N_6044);
or U6964 (N_6964,N_6086,N_6219);
nor U6965 (N_6965,N_6093,N_6247);
and U6966 (N_6966,N_6278,N_6445);
or U6967 (N_6967,N_6542,N_6197);
nand U6968 (N_6968,N_6060,N_6394);
and U6969 (N_6969,N_6668,N_6493);
or U6970 (N_6970,N_6698,N_6151);
nor U6971 (N_6971,N_6697,N_6153);
or U6972 (N_6972,N_6607,N_6469);
and U6973 (N_6973,N_6036,N_6451);
xor U6974 (N_6974,N_6688,N_6123);
and U6975 (N_6975,N_6127,N_6742);
nand U6976 (N_6976,N_6268,N_6412);
and U6977 (N_6977,N_6107,N_6218);
nor U6978 (N_6978,N_6099,N_6515);
and U6979 (N_6979,N_6174,N_6716);
or U6980 (N_6980,N_6740,N_6566);
nor U6981 (N_6981,N_6448,N_6609);
nand U6982 (N_6982,N_6604,N_6723);
and U6983 (N_6983,N_6539,N_6443);
or U6984 (N_6984,N_6136,N_6685);
nor U6985 (N_6985,N_6037,N_6337);
nand U6986 (N_6986,N_6748,N_6180);
nor U6987 (N_6987,N_6711,N_6162);
and U6988 (N_6988,N_6222,N_6382);
nor U6989 (N_6989,N_6514,N_6355);
nor U6990 (N_6990,N_6616,N_6128);
or U6991 (N_6991,N_6000,N_6651);
and U6992 (N_6992,N_6674,N_6403);
and U6993 (N_6993,N_6700,N_6079);
nor U6994 (N_6994,N_6692,N_6231);
nand U6995 (N_6995,N_6453,N_6436);
nand U6996 (N_6996,N_6223,N_6667);
or U6997 (N_6997,N_6624,N_6679);
nand U6998 (N_6998,N_6167,N_6213);
or U6999 (N_6999,N_6324,N_6085);
nand U7000 (N_7000,N_6267,N_6179);
or U7001 (N_7001,N_6299,N_6072);
nand U7002 (N_7002,N_6735,N_6734);
nor U7003 (N_7003,N_6277,N_6321);
nand U7004 (N_7004,N_6549,N_6749);
or U7005 (N_7005,N_6318,N_6217);
nor U7006 (N_7006,N_6520,N_6307);
nor U7007 (N_7007,N_6351,N_6228);
xor U7008 (N_7008,N_6266,N_6477);
nor U7009 (N_7009,N_6389,N_6410);
nand U7010 (N_7010,N_6182,N_6462);
xor U7011 (N_7011,N_6120,N_6030);
nand U7012 (N_7012,N_6133,N_6634);
nand U7013 (N_7013,N_6572,N_6052);
and U7014 (N_7014,N_6326,N_6146);
and U7015 (N_7015,N_6710,N_6571);
nor U7016 (N_7016,N_6447,N_6286);
or U7017 (N_7017,N_6362,N_6320);
nand U7018 (N_7018,N_6488,N_6405);
and U7019 (N_7019,N_6690,N_6096);
nor U7020 (N_7020,N_6656,N_6256);
nor U7021 (N_7021,N_6516,N_6672);
and U7022 (N_7022,N_6498,N_6331);
or U7023 (N_7023,N_6699,N_6653);
and U7024 (N_7024,N_6626,N_6468);
or U7025 (N_7025,N_6154,N_6121);
nor U7026 (N_7026,N_6306,N_6729);
xor U7027 (N_7027,N_6163,N_6684);
and U7028 (N_7028,N_6737,N_6147);
and U7029 (N_7029,N_6361,N_6425);
nand U7030 (N_7030,N_6490,N_6200);
nor U7031 (N_7031,N_6484,N_6587);
nand U7032 (N_7032,N_6533,N_6067);
nor U7033 (N_7033,N_6553,N_6647);
and U7034 (N_7034,N_6346,N_6718);
or U7035 (N_7035,N_6038,N_6433);
and U7036 (N_7036,N_6657,N_6018);
and U7037 (N_7037,N_6345,N_6385);
xor U7038 (N_7038,N_6597,N_6033);
nor U7039 (N_7039,N_6029,N_6183);
xnor U7040 (N_7040,N_6454,N_6034);
nor U7041 (N_7041,N_6025,N_6230);
nand U7042 (N_7042,N_6071,N_6148);
and U7043 (N_7043,N_6138,N_6260);
and U7044 (N_7044,N_6144,N_6245);
nand U7045 (N_7045,N_6316,N_6280);
nand U7046 (N_7046,N_6693,N_6248);
and U7047 (N_7047,N_6032,N_6122);
nor U7048 (N_7048,N_6296,N_6323);
or U7049 (N_7049,N_6721,N_6095);
xnor U7050 (N_7050,N_6367,N_6040);
nand U7051 (N_7051,N_6081,N_6595);
nand U7052 (N_7052,N_6473,N_6387);
or U7053 (N_7053,N_6413,N_6111);
or U7054 (N_7054,N_6746,N_6670);
xnor U7055 (N_7055,N_6204,N_6557);
nand U7056 (N_7056,N_6466,N_6232);
nand U7057 (N_7057,N_6564,N_6442);
nor U7058 (N_7058,N_6165,N_6057);
and U7059 (N_7059,N_6171,N_6628);
and U7060 (N_7060,N_6176,N_6156);
nor U7061 (N_7061,N_6643,N_6439);
and U7062 (N_7062,N_6215,N_6106);
nand U7063 (N_7063,N_6449,N_6281);
or U7064 (N_7064,N_6241,N_6041);
nor U7065 (N_7065,N_6262,N_6305);
nor U7066 (N_7066,N_6659,N_6371);
xnor U7067 (N_7067,N_6226,N_6108);
nand U7068 (N_7068,N_6460,N_6494);
and U7069 (N_7069,N_6510,N_6206);
or U7070 (N_7070,N_6456,N_6638);
and U7071 (N_7071,N_6603,N_6701);
and U7072 (N_7072,N_6497,N_6269);
and U7073 (N_7073,N_6199,N_6098);
and U7074 (N_7074,N_6719,N_6352);
nor U7075 (N_7075,N_6500,N_6545);
or U7076 (N_7076,N_6438,N_6290);
xnor U7077 (N_7077,N_6584,N_6496);
nor U7078 (N_7078,N_6457,N_6254);
and U7079 (N_7079,N_6293,N_6062);
xor U7080 (N_7080,N_6573,N_6649);
nand U7081 (N_7081,N_6270,N_6314);
xnor U7082 (N_7082,N_6580,N_6532);
and U7083 (N_7083,N_6606,N_6598);
xnor U7084 (N_7084,N_6623,N_6745);
nor U7085 (N_7085,N_6322,N_6393);
and U7086 (N_7086,N_6615,N_6185);
nor U7087 (N_7087,N_6175,N_6243);
nor U7088 (N_7088,N_6069,N_6582);
or U7089 (N_7089,N_6091,N_6625);
nor U7090 (N_7090,N_6680,N_6614);
nor U7091 (N_7091,N_6478,N_6227);
nor U7092 (N_7092,N_6577,N_6733);
or U7093 (N_7093,N_6169,N_6088);
nand U7094 (N_7094,N_6487,N_6421);
xnor U7095 (N_7095,N_6285,N_6235);
or U7096 (N_7096,N_6078,N_6172);
nand U7097 (N_7097,N_6357,N_6257);
nor U7098 (N_7098,N_6335,N_6554);
nor U7099 (N_7099,N_6059,N_6341);
and U7100 (N_7100,N_6409,N_6344);
or U7101 (N_7101,N_6400,N_6419);
nand U7102 (N_7102,N_6031,N_6654);
or U7103 (N_7103,N_6505,N_6205);
xnor U7104 (N_7104,N_6203,N_6102);
nand U7105 (N_7105,N_6524,N_6229);
and U7106 (N_7106,N_6045,N_6132);
and U7107 (N_7107,N_6142,N_6141);
or U7108 (N_7108,N_6474,N_6485);
xor U7109 (N_7109,N_6010,N_6550);
and U7110 (N_7110,N_6722,N_6538);
nor U7111 (N_7111,N_6310,N_6617);
xnor U7112 (N_7112,N_6130,N_6390);
and U7113 (N_7113,N_6158,N_6149);
nor U7114 (N_7114,N_6636,N_6455);
and U7115 (N_7115,N_6300,N_6677);
or U7116 (N_7116,N_6077,N_6622);
or U7117 (N_7117,N_6201,N_6396);
nor U7118 (N_7118,N_6347,N_6272);
nand U7119 (N_7119,N_6586,N_6639);
nor U7120 (N_7120,N_6340,N_6706);
or U7121 (N_7121,N_6592,N_6225);
nand U7122 (N_7122,N_6363,N_6437);
nand U7123 (N_7123,N_6048,N_6379);
xor U7124 (N_7124,N_6075,N_6242);
nand U7125 (N_7125,N_6539,N_6425);
and U7126 (N_7126,N_6329,N_6210);
xnor U7127 (N_7127,N_6689,N_6287);
or U7128 (N_7128,N_6071,N_6511);
nand U7129 (N_7129,N_6423,N_6622);
or U7130 (N_7130,N_6710,N_6695);
or U7131 (N_7131,N_6590,N_6515);
nand U7132 (N_7132,N_6701,N_6642);
nor U7133 (N_7133,N_6455,N_6368);
or U7134 (N_7134,N_6542,N_6651);
nor U7135 (N_7135,N_6353,N_6658);
xnor U7136 (N_7136,N_6150,N_6031);
nor U7137 (N_7137,N_6112,N_6075);
nor U7138 (N_7138,N_6516,N_6371);
nand U7139 (N_7139,N_6096,N_6452);
nor U7140 (N_7140,N_6491,N_6420);
nand U7141 (N_7141,N_6491,N_6012);
nor U7142 (N_7142,N_6495,N_6133);
or U7143 (N_7143,N_6516,N_6416);
or U7144 (N_7144,N_6619,N_6177);
xnor U7145 (N_7145,N_6539,N_6509);
nand U7146 (N_7146,N_6442,N_6736);
xor U7147 (N_7147,N_6620,N_6338);
or U7148 (N_7148,N_6280,N_6563);
and U7149 (N_7149,N_6138,N_6433);
nor U7150 (N_7150,N_6443,N_6464);
and U7151 (N_7151,N_6364,N_6493);
and U7152 (N_7152,N_6449,N_6732);
nand U7153 (N_7153,N_6129,N_6152);
nor U7154 (N_7154,N_6374,N_6175);
or U7155 (N_7155,N_6538,N_6112);
or U7156 (N_7156,N_6229,N_6348);
nand U7157 (N_7157,N_6702,N_6488);
and U7158 (N_7158,N_6392,N_6717);
xor U7159 (N_7159,N_6345,N_6692);
and U7160 (N_7160,N_6305,N_6567);
xnor U7161 (N_7161,N_6185,N_6696);
and U7162 (N_7162,N_6132,N_6010);
nor U7163 (N_7163,N_6171,N_6681);
nor U7164 (N_7164,N_6648,N_6392);
xor U7165 (N_7165,N_6384,N_6001);
nand U7166 (N_7166,N_6186,N_6465);
nand U7167 (N_7167,N_6193,N_6477);
xor U7168 (N_7168,N_6289,N_6210);
xnor U7169 (N_7169,N_6407,N_6000);
or U7170 (N_7170,N_6198,N_6698);
nor U7171 (N_7171,N_6005,N_6465);
and U7172 (N_7172,N_6053,N_6068);
and U7173 (N_7173,N_6136,N_6515);
nand U7174 (N_7174,N_6360,N_6676);
nor U7175 (N_7175,N_6039,N_6572);
nor U7176 (N_7176,N_6394,N_6726);
or U7177 (N_7177,N_6141,N_6416);
and U7178 (N_7178,N_6156,N_6443);
and U7179 (N_7179,N_6030,N_6439);
or U7180 (N_7180,N_6042,N_6668);
xor U7181 (N_7181,N_6225,N_6607);
and U7182 (N_7182,N_6292,N_6416);
xnor U7183 (N_7183,N_6684,N_6174);
nand U7184 (N_7184,N_6268,N_6637);
nand U7185 (N_7185,N_6578,N_6037);
and U7186 (N_7186,N_6006,N_6697);
nor U7187 (N_7187,N_6276,N_6517);
nand U7188 (N_7188,N_6194,N_6089);
xor U7189 (N_7189,N_6077,N_6309);
and U7190 (N_7190,N_6118,N_6593);
nor U7191 (N_7191,N_6378,N_6320);
and U7192 (N_7192,N_6115,N_6621);
nor U7193 (N_7193,N_6180,N_6413);
nor U7194 (N_7194,N_6262,N_6198);
and U7195 (N_7195,N_6091,N_6054);
nor U7196 (N_7196,N_6669,N_6141);
nor U7197 (N_7197,N_6550,N_6279);
nand U7198 (N_7198,N_6673,N_6614);
or U7199 (N_7199,N_6674,N_6352);
nor U7200 (N_7200,N_6115,N_6091);
and U7201 (N_7201,N_6734,N_6238);
nand U7202 (N_7202,N_6582,N_6080);
xor U7203 (N_7203,N_6409,N_6135);
nor U7204 (N_7204,N_6239,N_6340);
nand U7205 (N_7205,N_6676,N_6190);
and U7206 (N_7206,N_6110,N_6457);
nand U7207 (N_7207,N_6544,N_6044);
xnor U7208 (N_7208,N_6368,N_6743);
or U7209 (N_7209,N_6373,N_6323);
nand U7210 (N_7210,N_6532,N_6689);
xor U7211 (N_7211,N_6021,N_6443);
xnor U7212 (N_7212,N_6043,N_6392);
nand U7213 (N_7213,N_6297,N_6096);
or U7214 (N_7214,N_6312,N_6535);
nor U7215 (N_7215,N_6484,N_6726);
nand U7216 (N_7216,N_6033,N_6199);
or U7217 (N_7217,N_6432,N_6505);
xnor U7218 (N_7218,N_6559,N_6494);
xor U7219 (N_7219,N_6276,N_6587);
nand U7220 (N_7220,N_6377,N_6312);
nand U7221 (N_7221,N_6167,N_6428);
nand U7222 (N_7222,N_6719,N_6375);
or U7223 (N_7223,N_6694,N_6588);
nand U7224 (N_7224,N_6270,N_6661);
and U7225 (N_7225,N_6718,N_6716);
xor U7226 (N_7226,N_6397,N_6290);
or U7227 (N_7227,N_6159,N_6349);
xor U7228 (N_7228,N_6504,N_6312);
nand U7229 (N_7229,N_6163,N_6443);
nor U7230 (N_7230,N_6148,N_6712);
and U7231 (N_7231,N_6514,N_6596);
or U7232 (N_7232,N_6299,N_6508);
nor U7233 (N_7233,N_6240,N_6039);
nor U7234 (N_7234,N_6440,N_6112);
or U7235 (N_7235,N_6050,N_6609);
nor U7236 (N_7236,N_6174,N_6064);
xor U7237 (N_7237,N_6679,N_6430);
or U7238 (N_7238,N_6238,N_6146);
nor U7239 (N_7239,N_6600,N_6432);
nor U7240 (N_7240,N_6294,N_6093);
or U7241 (N_7241,N_6640,N_6216);
and U7242 (N_7242,N_6705,N_6019);
and U7243 (N_7243,N_6632,N_6108);
nand U7244 (N_7244,N_6616,N_6424);
or U7245 (N_7245,N_6453,N_6609);
nand U7246 (N_7246,N_6721,N_6709);
nor U7247 (N_7247,N_6292,N_6401);
nand U7248 (N_7248,N_6739,N_6368);
or U7249 (N_7249,N_6155,N_6580);
or U7250 (N_7250,N_6674,N_6119);
or U7251 (N_7251,N_6468,N_6410);
nor U7252 (N_7252,N_6685,N_6651);
nor U7253 (N_7253,N_6647,N_6406);
or U7254 (N_7254,N_6073,N_6427);
and U7255 (N_7255,N_6297,N_6458);
or U7256 (N_7256,N_6002,N_6710);
or U7257 (N_7257,N_6195,N_6529);
nand U7258 (N_7258,N_6312,N_6749);
and U7259 (N_7259,N_6571,N_6023);
nor U7260 (N_7260,N_6089,N_6297);
or U7261 (N_7261,N_6670,N_6357);
nor U7262 (N_7262,N_6123,N_6191);
nor U7263 (N_7263,N_6503,N_6127);
nor U7264 (N_7264,N_6691,N_6468);
nand U7265 (N_7265,N_6563,N_6287);
nand U7266 (N_7266,N_6509,N_6367);
or U7267 (N_7267,N_6737,N_6611);
xnor U7268 (N_7268,N_6102,N_6251);
xor U7269 (N_7269,N_6579,N_6575);
and U7270 (N_7270,N_6415,N_6370);
and U7271 (N_7271,N_6503,N_6665);
nor U7272 (N_7272,N_6526,N_6533);
or U7273 (N_7273,N_6581,N_6371);
and U7274 (N_7274,N_6716,N_6440);
nand U7275 (N_7275,N_6567,N_6114);
nand U7276 (N_7276,N_6271,N_6118);
nand U7277 (N_7277,N_6476,N_6109);
and U7278 (N_7278,N_6055,N_6181);
nand U7279 (N_7279,N_6491,N_6203);
or U7280 (N_7280,N_6360,N_6155);
and U7281 (N_7281,N_6263,N_6451);
nand U7282 (N_7282,N_6398,N_6742);
nor U7283 (N_7283,N_6219,N_6646);
or U7284 (N_7284,N_6211,N_6745);
nor U7285 (N_7285,N_6553,N_6261);
nor U7286 (N_7286,N_6258,N_6484);
nor U7287 (N_7287,N_6532,N_6300);
nor U7288 (N_7288,N_6372,N_6303);
nand U7289 (N_7289,N_6595,N_6606);
nand U7290 (N_7290,N_6499,N_6474);
or U7291 (N_7291,N_6236,N_6472);
nor U7292 (N_7292,N_6340,N_6177);
and U7293 (N_7293,N_6260,N_6222);
and U7294 (N_7294,N_6511,N_6500);
nand U7295 (N_7295,N_6117,N_6547);
nand U7296 (N_7296,N_6296,N_6597);
nand U7297 (N_7297,N_6086,N_6295);
and U7298 (N_7298,N_6507,N_6322);
or U7299 (N_7299,N_6299,N_6684);
xnor U7300 (N_7300,N_6619,N_6479);
and U7301 (N_7301,N_6453,N_6015);
nand U7302 (N_7302,N_6468,N_6374);
nand U7303 (N_7303,N_6712,N_6463);
xnor U7304 (N_7304,N_6198,N_6500);
nand U7305 (N_7305,N_6026,N_6529);
and U7306 (N_7306,N_6014,N_6605);
and U7307 (N_7307,N_6627,N_6390);
nor U7308 (N_7308,N_6179,N_6313);
xor U7309 (N_7309,N_6079,N_6351);
nor U7310 (N_7310,N_6444,N_6340);
nand U7311 (N_7311,N_6371,N_6558);
and U7312 (N_7312,N_6646,N_6350);
and U7313 (N_7313,N_6093,N_6590);
nor U7314 (N_7314,N_6252,N_6149);
xor U7315 (N_7315,N_6081,N_6709);
and U7316 (N_7316,N_6421,N_6273);
or U7317 (N_7317,N_6073,N_6091);
xnor U7318 (N_7318,N_6263,N_6419);
xor U7319 (N_7319,N_6130,N_6483);
and U7320 (N_7320,N_6633,N_6664);
nand U7321 (N_7321,N_6452,N_6030);
nand U7322 (N_7322,N_6012,N_6476);
xnor U7323 (N_7323,N_6728,N_6495);
nand U7324 (N_7324,N_6559,N_6423);
xnor U7325 (N_7325,N_6287,N_6612);
or U7326 (N_7326,N_6510,N_6475);
and U7327 (N_7327,N_6178,N_6304);
nand U7328 (N_7328,N_6131,N_6366);
xor U7329 (N_7329,N_6526,N_6673);
xor U7330 (N_7330,N_6514,N_6470);
and U7331 (N_7331,N_6455,N_6447);
and U7332 (N_7332,N_6041,N_6163);
and U7333 (N_7333,N_6658,N_6047);
and U7334 (N_7334,N_6310,N_6402);
nand U7335 (N_7335,N_6385,N_6690);
or U7336 (N_7336,N_6013,N_6308);
and U7337 (N_7337,N_6210,N_6704);
or U7338 (N_7338,N_6169,N_6269);
nor U7339 (N_7339,N_6543,N_6078);
and U7340 (N_7340,N_6505,N_6249);
nor U7341 (N_7341,N_6337,N_6300);
nor U7342 (N_7342,N_6592,N_6620);
or U7343 (N_7343,N_6645,N_6557);
or U7344 (N_7344,N_6523,N_6279);
xor U7345 (N_7345,N_6472,N_6195);
or U7346 (N_7346,N_6029,N_6386);
nand U7347 (N_7347,N_6236,N_6616);
nand U7348 (N_7348,N_6483,N_6371);
or U7349 (N_7349,N_6300,N_6628);
or U7350 (N_7350,N_6674,N_6506);
nor U7351 (N_7351,N_6603,N_6236);
nor U7352 (N_7352,N_6195,N_6135);
xor U7353 (N_7353,N_6500,N_6462);
xor U7354 (N_7354,N_6151,N_6084);
or U7355 (N_7355,N_6078,N_6120);
and U7356 (N_7356,N_6353,N_6472);
xnor U7357 (N_7357,N_6596,N_6153);
and U7358 (N_7358,N_6523,N_6190);
xor U7359 (N_7359,N_6280,N_6729);
or U7360 (N_7360,N_6611,N_6570);
or U7361 (N_7361,N_6701,N_6485);
nor U7362 (N_7362,N_6162,N_6588);
and U7363 (N_7363,N_6143,N_6735);
or U7364 (N_7364,N_6175,N_6549);
nor U7365 (N_7365,N_6212,N_6376);
nand U7366 (N_7366,N_6056,N_6562);
or U7367 (N_7367,N_6595,N_6233);
nand U7368 (N_7368,N_6233,N_6372);
and U7369 (N_7369,N_6397,N_6651);
and U7370 (N_7370,N_6558,N_6397);
or U7371 (N_7371,N_6033,N_6417);
xor U7372 (N_7372,N_6086,N_6274);
nor U7373 (N_7373,N_6556,N_6152);
nor U7374 (N_7374,N_6264,N_6624);
and U7375 (N_7375,N_6566,N_6224);
or U7376 (N_7376,N_6456,N_6633);
and U7377 (N_7377,N_6275,N_6505);
nand U7378 (N_7378,N_6010,N_6740);
or U7379 (N_7379,N_6715,N_6151);
nor U7380 (N_7380,N_6654,N_6705);
xnor U7381 (N_7381,N_6698,N_6691);
nor U7382 (N_7382,N_6223,N_6310);
nor U7383 (N_7383,N_6569,N_6400);
nand U7384 (N_7384,N_6180,N_6673);
or U7385 (N_7385,N_6682,N_6342);
and U7386 (N_7386,N_6725,N_6109);
xor U7387 (N_7387,N_6474,N_6600);
nand U7388 (N_7388,N_6737,N_6094);
or U7389 (N_7389,N_6031,N_6020);
nor U7390 (N_7390,N_6186,N_6217);
or U7391 (N_7391,N_6285,N_6571);
and U7392 (N_7392,N_6410,N_6667);
or U7393 (N_7393,N_6436,N_6141);
or U7394 (N_7394,N_6689,N_6396);
nand U7395 (N_7395,N_6711,N_6085);
or U7396 (N_7396,N_6238,N_6415);
nor U7397 (N_7397,N_6553,N_6705);
and U7398 (N_7398,N_6249,N_6570);
and U7399 (N_7399,N_6095,N_6214);
nor U7400 (N_7400,N_6490,N_6377);
nor U7401 (N_7401,N_6383,N_6295);
or U7402 (N_7402,N_6270,N_6743);
nor U7403 (N_7403,N_6375,N_6104);
or U7404 (N_7404,N_6311,N_6257);
or U7405 (N_7405,N_6287,N_6613);
nand U7406 (N_7406,N_6152,N_6357);
nor U7407 (N_7407,N_6655,N_6514);
nand U7408 (N_7408,N_6351,N_6391);
xor U7409 (N_7409,N_6745,N_6226);
nor U7410 (N_7410,N_6677,N_6319);
or U7411 (N_7411,N_6656,N_6211);
nor U7412 (N_7412,N_6553,N_6655);
nand U7413 (N_7413,N_6289,N_6243);
nand U7414 (N_7414,N_6552,N_6642);
and U7415 (N_7415,N_6366,N_6343);
or U7416 (N_7416,N_6521,N_6643);
or U7417 (N_7417,N_6382,N_6705);
xnor U7418 (N_7418,N_6303,N_6087);
xor U7419 (N_7419,N_6714,N_6637);
or U7420 (N_7420,N_6603,N_6344);
nand U7421 (N_7421,N_6722,N_6002);
nor U7422 (N_7422,N_6002,N_6223);
nand U7423 (N_7423,N_6657,N_6245);
nor U7424 (N_7424,N_6472,N_6672);
or U7425 (N_7425,N_6406,N_6117);
nand U7426 (N_7426,N_6408,N_6484);
or U7427 (N_7427,N_6657,N_6670);
xnor U7428 (N_7428,N_6718,N_6373);
and U7429 (N_7429,N_6206,N_6217);
and U7430 (N_7430,N_6477,N_6665);
xor U7431 (N_7431,N_6390,N_6239);
and U7432 (N_7432,N_6128,N_6118);
xnor U7433 (N_7433,N_6140,N_6112);
and U7434 (N_7434,N_6041,N_6193);
nand U7435 (N_7435,N_6158,N_6741);
xnor U7436 (N_7436,N_6100,N_6600);
or U7437 (N_7437,N_6296,N_6088);
nor U7438 (N_7438,N_6687,N_6063);
nand U7439 (N_7439,N_6668,N_6611);
and U7440 (N_7440,N_6423,N_6516);
and U7441 (N_7441,N_6736,N_6130);
and U7442 (N_7442,N_6170,N_6166);
xnor U7443 (N_7443,N_6043,N_6351);
xor U7444 (N_7444,N_6652,N_6074);
and U7445 (N_7445,N_6359,N_6617);
nor U7446 (N_7446,N_6459,N_6218);
nand U7447 (N_7447,N_6651,N_6475);
xnor U7448 (N_7448,N_6598,N_6459);
nand U7449 (N_7449,N_6068,N_6326);
or U7450 (N_7450,N_6662,N_6418);
nand U7451 (N_7451,N_6180,N_6005);
nand U7452 (N_7452,N_6696,N_6083);
or U7453 (N_7453,N_6220,N_6603);
or U7454 (N_7454,N_6465,N_6700);
xor U7455 (N_7455,N_6327,N_6465);
nand U7456 (N_7456,N_6155,N_6725);
or U7457 (N_7457,N_6657,N_6747);
and U7458 (N_7458,N_6396,N_6001);
xnor U7459 (N_7459,N_6434,N_6085);
or U7460 (N_7460,N_6726,N_6567);
or U7461 (N_7461,N_6396,N_6239);
xor U7462 (N_7462,N_6644,N_6096);
and U7463 (N_7463,N_6536,N_6716);
and U7464 (N_7464,N_6579,N_6260);
nor U7465 (N_7465,N_6159,N_6704);
or U7466 (N_7466,N_6653,N_6644);
nor U7467 (N_7467,N_6298,N_6010);
or U7468 (N_7468,N_6386,N_6566);
nor U7469 (N_7469,N_6692,N_6589);
nor U7470 (N_7470,N_6541,N_6615);
nand U7471 (N_7471,N_6115,N_6389);
and U7472 (N_7472,N_6159,N_6679);
nand U7473 (N_7473,N_6542,N_6697);
nor U7474 (N_7474,N_6357,N_6662);
and U7475 (N_7475,N_6268,N_6505);
nand U7476 (N_7476,N_6339,N_6473);
and U7477 (N_7477,N_6398,N_6378);
nor U7478 (N_7478,N_6533,N_6516);
or U7479 (N_7479,N_6323,N_6547);
nand U7480 (N_7480,N_6199,N_6371);
or U7481 (N_7481,N_6329,N_6243);
xor U7482 (N_7482,N_6362,N_6269);
nand U7483 (N_7483,N_6184,N_6539);
and U7484 (N_7484,N_6597,N_6711);
nor U7485 (N_7485,N_6653,N_6669);
or U7486 (N_7486,N_6676,N_6512);
nor U7487 (N_7487,N_6314,N_6198);
nand U7488 (N_7488,N_6619,N_6376);
and U7489 (N_7489,N_6068,N_6218);
and U7490 (N_7490,N_6705,N_6330);
nand U7491 (N_7491,N_6689,N_6037);
or U7492 (N_7492,N_6001,N_6651);
nand U7493 (N_7493,N_6421,N_6439);
nand U7494 (N_7494,N_6326,N_6404);
and U7495 (N_7495,N_6420,N_6188);
and U7496 (N_7496,N_6255,N_6399);
nand U7497 (N_7497,N_6265,N_6493);
xor U7498 (N_7498,N_6155,N_6096);
nand U7499 (N_7499,N_6202,N_6277);
nand U7500 (N_7500,N_7109,N_7210);
nand U7501 (N_7501,N_7255,N_7405);
xor U7502 (N_7502,N_7192,N_7181);
nor U7503 (N_7503,N_7009,N_7498);
nand U7504 (N_7504,N_7486,N_6914);
or U7505 (N_7505,N_7441,N_7048);
nor U7506 (N_7506,N_7477,N_7375);
nor U7507 (N_7507,N_6927,N_7120);
xnor U7508 (N_7508,N_7424,N_7444);
nand U7509 (N_7509,N_7184,N_6824);
nor U7510 (N_7510,N_7067,N_6990);
and U7511 (N_7511,N_7202,N_7413);
xnor U7512 (N_7512,N_6835,N_7332);
or U7513 (N_7513,N_7061,N_7302);
nor U7514 (N_7514,N_7482,N_7215);
nor U7515 (N_7515,N_7133,N_7260);
and U7516 (N_7516,N_6834,N_7279);
and U7517 (N_7517,N_7071,N_6888);
nor U7518 (N_7518,N_6836,N_7068);
and U7519 (N_7519,N_7174,N_7226);
nor U7520 (N_7520,N_7420,N_6881);
nand U7521 (N_7521,N_7209,N_7101);
nor U7522 (N_7522,N_7348,N_6801);
nor U7523 (N_7523,N_6754,N_7432);
nand U7524 (N_7524,N_7337,N_7082);
and U7525 (N_7525,N_7126,N_6929);
and U7526 (N_7526,N_7100,N_7435);
nor U7527 (N_7527,N_7154,N_7195);
nand U7528 (N_7528,N_7028,N_6902);
and U7529 (N_7529,N_6892,N_7378);
or U7530 (N_7530,N_7415,N_7197);
or U7531 (N_7531,N_7236,N_7468);
nor U7532 (N_7532,N_6961,N_7496);
and U7533 (N_7533,N_7066,N_7078);
or U7534 (N_7534,N_7092,N_7326);
nand U7535 (N_7535,N_7085,N_7096);
or U7536 (N_7536,N_7024,N_7450);
xor U7537 (N_7537,N_7385,N_7227);
nand U7538 (N_7538,N_7475,N_7162);
or U7539 (N_7539,N_7060,N_7318);
nand U7540 (N_7540,N_7291,N_7178);
and U7541 (N_7541,N_7214,N_6986);
nand U7542 (N_7542,N_7419,N_7108);
and U7543 (N_7543,N_6793,N_6829);
nor U7544 (N_7544,N_6758,N_6753);
or U7545 (N_7545,N_7084,N_7252);
and U7546 (N_7546,N_7485,N_7118);
nor U7547 (N_7547,N_7299,N_6864);
xnor U7548 (N_7548,N_6890,N_6819);
xnor U7549 (N_7549,N_7220,N_7153);
nand U7550 (N_7550,N_6974,N_6932);
xnor U7551 (N_7551,N_6772,N_7171);
nand U7552 (N_7552,N_6830,N_7287);
nand U7553 (N_7553,N_6942,N_7044);
and U7554 (N_7554,N_7191,N_6878);
and U7555 (N_7555,N_7314,N_6977);
nor U7556 (N_7556,N_6783,N_6940);
and U7557 (N_7557,N_7081,N_7063);
and U7558 (N_7558,N_7165,N_7446);
xnor U7559 (N_7559,N_6782,N_6759);
and U7560 (N_7560,N_7377,N_7073);
nand U7561 (N_7561,N_7104,N_7380);
nor U7562 (N_7562,N_7203,N_7199);
nor U7563 (N_7563,N_7272,N_6963);
xor U7564 (N_7564,N_6854,N_7484);
nor U7565 (N_7565,N_6839,N_7286);
or U7566 (N_7566,N_6833,N_6761);
nand U7567 (N_7567,N_6943,N_6915);
nand U7568 (N_7568,N_7264,N_7400);
or U7569 (N_7569,N_7399,N_7059);
nand U7570 (N_7570,N_6950,N_7176);
or U7571 (N_7571,N_7459,N_7017);
or U7572 (N_7572,N_7443,N_6857);
or U7573 (N_7573,N_7295,N_6844);
and U7574 (N_7574,N_6906,N_7053);
and U7575 (N_7575,N_6838,N_6869);
and U7576 (N_7576,N_6802,N_7389);
or U7577 (N_7577,N_7004,N_7304);
or U7578 (N_7578,N_7397,N_7351);
or U7579 (N_7579,N_7107,N_7379);
and U7580 (N_7580,N_7265,N_7343);
or U7581 (N_7581,N_6922,N_7467);
and U7582 (N_7582,N_6887,N_7499);
or U7583 (N_7583,N_6889,N_7269);
or U7584 (N_7584,N_6936,N_7311);
nand U7585 (N_7585,N_6752,N_6894);
nand U7586 (N_7586,N_6945,N_7026);
and U7587 (N_7587,N_6938,N_6908);
nand U7588 (N_7588,N_7131,N_6980);
nor U7589 (N_7589,N_7452,N_7228);
and U7590 (N_7590,N_6930,N_6780);
nand U7591 (N_7591,N_7451,N_6868);
or U7592 (N_7592,N_7305,N_7079);
nor U7593 (N_7593,N_6787,N_6764);
or U7594 (N_7594,N_6918,N_6928);
or U7595 (N_7595,N_7074,N_7278);
nor U7596 (N_7596,N_7409,N_7289);
and U7597 (N_7597,N_7022,N_7157);
nor U7598 (N_7598,N_7367,N_7119);
and U7599 (N_7599,N_7117,N_6806);
nand U7600 (N_7600,N_7231,N_6852);
and U7601 (N_7601,N_7453,N_7402);
and U7602 (N_7602,N_6978,N_7350);
nor U7603 (N_7603,N_6847,N_7390);
nor U7604 (N_7604,N_6919,N_7470);
nand U7605 (N_7605,N_6882,N_6900);
and U7606 (N_7606,N_6968,N_6954);
nand U7607 (N_7607,N_7075,N_6766);
and U7608 (N_7608,N_6804,N_6840);
or U7609 (N_7609,N_6907,N_7064);
or U7610 (N_7610,N_7110,N_7325);
nand U7611 (N_7611,N_7128,N_7427);
or U7612 (N_7612,N_7247,N_7431);
nor U7613 (N_7613,N_6867,N_7448);
or U7614 (N_7614,N_6973,N_7010);
nand U7615 (N_7615,N_7412,N_6821);
nand U7616 (N_7616,N_7457,N_7015);
xnor U7617 (N_7617,N_7102,N_7455);
nor U7618 (N_7618,N_6891,N_6988);
or U7619 (N_7619,N_7246,N_7386);
or U7620 (N_7620,N_6750,N_7393);
or U7621 (N_7621,N_6760,N_6941);
or U7622 (N_7622,N_7354,N_7481);
or U7623 (N_7623,N_6858,N_6933);
or U7624 (N_7624,N_7211,N_6816);
or U7625 (N_7625,N_6874,N_6998);
and U7626 (N_7626,N_7140,N_7320);
or U7627 (N_7627,N_7275,N_7323);
or U7628 (N_7628,N_7250,N_7298);
nor U7629 (N_7629,N_7147,N_6897);
nand U7630 (N_7630,N_6755,N_7045);
nor U7631 (N_7631,N_7346,N_7168);
and U7632 (N_7632,N_7205,N_7463);
and U7633 (N_7633,N_7051,N_7098);
or U7634 (N_7634,N_6994,N_7113);
nand U7635 (N_7635,N_6850,N_6953);
xnor U7636 (N_7636,N_7033,N_7173);
nand U7637 (N_7637,N_7274,N_6967);
or U7638 (N_7638,N_7186,N_6789);
nand U7639 (N_7639,N_7458,N_6926);
nand U7640 (N_7640,N_6814,N_7035);
or U7641 (N_7641,N_7369,N_7421);
and U7642 (N_7642,N_7480,N_7471);
nand U7643 (N_7643,N_7317,N_7127);
and U7644 (N_7644,N_7262,N_7341);
or U7645 (N_7645,N_7232,N_6810);
and U7646 (N_7646,N_6939,N_6981);
nor U7647 (N_7647,N_7495,N_6831);
xor U7648 (N_7648,N_6879,N_6811);
nor U7649 (N_7649,N_7077,N_6822);
nand U7650 (N_7650,N_6898,N_6958);
or U7651 (N_7651,N_7259,N_7103);
xor U7652 (N_7652,N_7138,N_7285);
nor U7653 (N_7653,N_6866,N_6883);
or U7654 (N_7654,N_7179,N_6809);
or U7655 (N_7655,N_7404,N_7465);
and U7656 (N_7656,N_7461,N_7288);
nand U7657 (N_7657,N_7454,N_7099);
or U7658 (N_7658,N_7036,N_7093);
nand U7659 (N_7659,N_6777,N_6962);
nand U7660 (N_7660,N_7002,N_7169);
nor U7661 (N_7661,N_6856,N_7237);
nor U7662 (N_7662,N_7437,N_6855);
xor U7663 (N_7663,N_6903,N_7141);
and U7664 (N_7664,N_7356,N_6909);
nor U7665 (N_7665,N_7057,N_7216);
nand U7666 (N_7666,N_7309,N_7387);
nor U7667 (N_7667,N_7308,N_7364);
nor U7668 (N_7668,N_6959,N_6957);
nor U7669 (N_7669,N_7392,N_7408);
nand U7670 (N_7670,N_7310,N_7200);
and U7671 (N_7671,N_6946,N_7294);
or U7672 (N_7672,N_7023,N_7156);
or U7673 (N_7673,N_6796,N_7012);
nand U7674 (N_7674,N_7124,N_7058);
nor U7675 (N_7675,N_6767,N_7353);
or U7676 (N_7676,N_7426,N_7115);
nor U7677 (N_7677,N_6825,N_7358);
and U7678 (N_7678,N_7307,N_7152);
nor U7679 (N_7679,N_7204,N_6917);
and U7680 (N_7680,N_6845,N_6989);
nor U7681 (N_7681,N_7160,N_7097);
and U7682 (N_7682,N_7473,N_6899);
nand U7683 (N_7683,N_6937,N_6861);
or U7684 (N_7684,N_6965,N_7217);
and U7685 (N_7685,N_6873,N_6901);
nor U7686 (N_7686,N_7383,N_7462);
and U7687 (N_7687,N_7362,N_6944);
nor U7688 (N_7688,N_7005,N_6876);
and U7689 (N_7689,N_7031,N_7225);
or U7690 (N_7690,N_7395,N_6853);
nor U7691 (N_7691,N_7041,N_7245);
and U7692 (N_7692,N_7042,N_7145);
nand U7693 (N_7693,N_7394,N_6948);
or U7694 (N_7694,N_6773,N_7207);
nor U7695 (N_7695,N_6972,N_6762);
or U7696 (N_7696,N_7373,N_7352);
and U7697 (N_7697,N_7371,N_7436);
or U7698 (N_7698,N_6960,N_7258);
and U7699 (N_7699,N_7396,N_7251);
nor U7700 (N_7700,N_7322,N_7034);
nand U7701 (N_7701,N_6949,N_6803);
and U7702 (N_7702,N_7449,N_7105);
nand U7703 (N_7703,N_7334,N_7312);
and U7704 (N_7704,N_7229,N_7000);
nor U7705 (N_7705,N_7201,N_6871);
nor U7706 (N_7706,N_7223,N_7052);
and U7707 (N_7707,N_7280,N_6911);
or U7708 (N_7708,N_7313,N_7328);
or U7709 (N_7709,N_6790,N_6827);
nand U7710 (N_7710,N_7430,N_6983);
and U7711 (N_7711,N_7206,N_6863);
and U7712 (N_7712,N_6774,N_7170);
or U7713 (N_7713,N_7129,N_7315);
nor U7714 (N_7714,N_6984,N_7142);
xnor U7715 (N_7715,N_6828,N_7194);
nand U7716 (N_7716,N_7407,N_6784);
or U7717 (N_7717,N_7406,N_7083);
and U7718 (N_7718,N_7188,N_7384);
nor U7719 (N_7719,N_6812,N_6875);
and U7720 (N_7720,N_7253,N_6815);
nor U7721 (N_7721,N_6924,N_6860);
and U7722 (N_7722,N_7198,N_7076);
nor U7723 (N_7723,N_6995,N_6923);
or U7724 (N_7724,N_7422,N_7149);
nor U7725 (N_7725,N_7489,N_6769);
or U7726 (N_7726,N_7055,N_7072);
and U7727 (N_7727,N_7243,N_7344);
nand U7728 (N_7728,N_7347,N_6786);
xnor U7729 (N_7729,N_7277,N_6770);
and U7730 (N_7730,N_7339,N_6987);
or U7731 (N_7731,N_6935,N_7248);
nor U7732 (N_7732,N_7111,N_6993);
or U7733 (N_7733,N_7150,N_7401);
and U7734 (N_7734,N_6808,N_6997);
xnor U7735 (N_7735,N_7479,N_7433);
and U7736 (N_7736,N_6820,N_6970);
nor U7737 (N_7737,N_7418,N_7376);
and U7738 (N_7738,N_7106,N_7290);
xor U7739 (N_7739,N_7382,N_6893);
nand U7740 (N_7740,N_7398,N_6931);
xor U7741 (N_7741,N_7239,N_7218);
or U7742 (N_7742,N_6768,N_7365);
and U7743 (N_7743,N_7233,N_6934);
or U7744 (N_7744,N_7013,N_7429);
and U7745 (N_7745,N_7027,N_7439);
nand U7746 (N_7746,N_6862,N_7135);
nand U7747 (N_7747,N_7266,N_6880);
nand U7748 (N_7748,N_7366,N_7018);
or U7749 (N_7749,N_7440,N_7158);
and U7750 (N_7750,N_7086,N_7306);
and U7751 (N_7751,N_7242,N_7333);
nand U7752 (N_7752,N_7193,N_7370);
and U7753 (N_7753,N_7241,N_7182);
nor U7754 (N_7754,N_7222,N_7038);
and U7755 (N_7755,N_6921,N_7230);
and U7756 (N_7756,N_6800,N_7423);
nor U7757 (N_7757,N_6859,N_7136);
nor U7758 (N_7758,N_7144,N_7177);
nand U7759 (N_7759,N_6916,N_7282);
nor U7760 (N_7760,N_7014,N_7020);
and U7761 (N_7761,N_7008,N_7273);
and U7762 (N_7762,N_7301,N_7006);
or U7763 (N_7763,N_6964,N_6870);
nand U7764 (N_7764,N_6895,N_7442);
and U7765 (N_7765,N_6791,N_6795);
nand U7766 (N_7766,N_6877,N_6886);
and U7767 (N_7767,N_7183,N_6788);
xor U7768 (N_7768,N_7039,N_7292);
and U7769 (N_7769,N_6912,N_7281);
nor U7770 (N_7770,N_6872,N_7056);
nor U7771 (N_7771,N_7032,N_7132);
or U7772 (N_7772,N_7316,N_7335);
nor U7773 (N_7773,N_7488,N_7491);
or U7774 (N_7774,N_7125,N_7297);
or U7775 (N_7775,N_7161,N_7094);
nor U7776 (N_7776,N_7187,N_7212);
nand U7777 (N_7777,N_7293,N_7345);
or U7778 (N_7778,N_7011,N_7411);
nor U7779 (N_7779,N_7047,N_6763);
or U7780 (N_7780,N_7490,N_7062);
and U7781 (N_7781,N_7434,N_7134);
nor U7782 (N_7782,N_7021,N_6781);
or U7783 (N_7783,N_6979,N_7151);
nand U7784 (N_7784,N_7487,N_6823);
nor U7785 (N_7785,N_7166,N_7372);
or U7786 (N_7786,N_6848,N_7284);
nor U7787 (N_7787,N_7342,N_6851);
and U7788 (N_7788,N_6813,N_7175);
or U7789 (N_7789,N_7240,N_7474);
nand U7790 (N_7790,N_6996,N_7219);
and U7791 (N_7791,N_7054,N_7329);
nand U7792 (N_7792,N_7137,N_7087);
and U7793 (N_7793,N_6778,N_6841);
or U7794 (N_7794,N_7112,N_7095);
or U7795 (N_7795,N_7003,N_7007);
and U7796 (N_7796,N_7167,N_6799);
nand U7797 (N_7797,N_7019,N_7050);
xnor U7798 (N_7798,N_7464,N_7276);
or U7799 (N_7799,N_7261,N_6966);
nand U7800 (N_7800,N_7361,N_7121);
nor U7801 (N_7801,N_7249,N_7472);
and U7802 (N_7802,N_6797,N_6982);
and U7803 (N_7803,N_7257,N_7324);
xor U7804 (N_7804,N_6832,N_7234);
nand U7805 (N_7805,N_7381,N_7303);
nand U7806 (N_7806,N_7224,N_7070);
nand U7807 (N_7807,N_7460,N_7091);
nor U7808 (N_7808,N_7355,N_6849);
and U7809 (N_7809,N_7359,N_7030);
or U7810 (N_7810,N_6955,N_7368);
nand U7811 (N_7811,N_6807,N_6969);
or U7812 (N_7812,N_6756,N_7331);
nand U7813 (N_7813,N_7494,N_7116);
or U7814 (N_7814,N_7123,N_7180);
xnor U7815 (N_7815,N_6884,N_6779);
or U7816 (N_7816,N_7040,N_6751);
nor U7817 (N_7817,N_6792,N_7296);
xnor U7818 (N_7818,N_7330,N_7391);
or U7819 (N_7819,N_6826,N_7148);
or U7820 (N_7820,N_7043,N_6976);
nand U7821 (N_7821,N_7374,N_7414);
xor U7822 (N_7822,N_7256,N_7088);
or U7823 (N_7823,N_6885,N_7069);
nand U7824 (N_7824,N_7476,N_6910);
nand U7825 (N_7825,N_7235,N_7029);
or U7826 (N_7826,N_6951,N_7447);
and U7827 (N_7827,N_7155,N_7139);
nor U7828 (N_7828,N_6913,N_7037);
and U7829 (N_7829,N_7159,N_6846);
nor U7830 (N_7830,N_7172,N_7065);
or U7831 (N_7831,N_6999,N_6818);
and U7832 (N_7832,N_7089,N_7466);
nand U7833 (N_7833,N_7146,N_7221);
nand U7834 (N_7834,N_7340,N_7438);
and U7835 (N_7835,N_7270,N_7016);
and U7836 (N_7836,N_6794,N_7208);
and U7837 (N_7837,N_7164,N_6991);
nand U7838 (N_7838,N_7493,N_7271);
nand U7839 (N_7839,N_7321,N_7338);
or U7840 (N_7840,N_7163,N_7492);
and U7841 (N_7841,N_6771,N_6896);
and U7842 (N_7842,N_6985,N_7363);
nor U7843 (N_7843,N_7049,N_6776);
xnor U7844 (N_7844,N_7319,N_6817);
or U7845 (N_7845,N_7445,N_7478);
or U7846 (N_7846,N_6843,N_7001);
nor U7847 (N_7847,N_6757,N_7417);
or U7848 (N_7848,N_7143,N_7114);
or U7849 (N_7849,N_7263,N_7238);
nand U7850 (N_7850,N_6865,N_7360);
nor U7851 (N_7851,N_7410,N_6947);
xnor U7852 (N_7852,N_6925,N_6992);
or U7853 (N_7853,N_7090,N_7283);
or U7854 (N_7854,N_7300,N_7425);
or U7855 (N_7855,N_6956,N_7428);
nor U7856 (N_7856,N_6971,N_6842);
nand U7857 (N_7857,N_7483,N_7080);
or U7858 (N_7858,N_6805,N_7196);
nor U7859 (N_7859,N_7268,N_7497);
or U7860 (N_7860,N_7349,N_7388);
or U7861 (N_7861,N_6905,N_7025);
xor U7862 (N_7862,N_6952,N_7336);
nor U7863 (N_7863,N_7130,N_7327);
or U7864 (N_7864,N_7267,N_7244);
xor U7865 (N_7865,N_6785,N_7189);
nor U7866 (N_7866,N_7254,N_7416);
and U7867 (N_7867,N_7122,N_6904);
and U7868 (N_7868,N_6765,N_7046);
nand U7869 (N_7869,N_6837,N_6775);
nor U7870 (N_7870,N_6920,N_7456);
and U7871 (N_7871,N_7403,N_7469);
or U7872 (N_7872,N_7190,N_7185);
nor U7873 (N_7873,N_7213,N_7357);
or U7874 (N_7874,N_6975,N_6798);
and U7875 (N_7875,N_6781,N_7407);
xor U7876 (N_7876,N_6848,N_7071);
nor U7877 (N_7877,N_6948,N_7270);
nand U7878 (N_7878,N_7467,N_7250);
or U7879 (N_7879,N_7365,N_7309);
nor U7880 (N_7880,N_7219,N_7276);
nor U7881 (N_7881,N_7347,N_6889);
and U7882 (N_7882,N_7068,N_7428);
or U7883 (N_7883,N_7367,N_6953);
nor U7884 (N_7884,N_7214,N_7462);
xor U7885 (N_7885,N_6799,N_7335);
nor U7886 (N_7886,N_7165,N_7401);
or U7887 (N_7887,N_6909,N_7166);
and U7888 (N_7888,N_7349,N_6753);
nand U7889 (N_7889,N_6996,N_6783);
and U7890 (N_7890,N_7322,N_7177);
and U7891 (N_7891,N_6948,N_6852);
and U7892 (N_7892,N_6921,N_6768);
nor U7893 (N_7893,N_7481,N_7459);
and U7894 (N_7894,N_6951,N_7475);
or U7895 (N_7895,N_7095,N_7308);
and U7896 (N_7896,N_7315,N_7439);
or U7897 (N_7897,N_7134,N_6845);
and U7898 (N_7898,N_7302,N_7451);
or U7899 (N_7899,N_6884,N_7270);
nand U7900 (N_7900,N_7029,N_7361);
and U7901 (N_7901,N_7075,N_6811);
or U7902 (N_7902,N_7119,N_7056);
or U7903 (N_7903,N_6944,N_7183);
nand U7904 (N_7904,N_7243,N_7165);
nand U7905 (N_7905,N_7413,N_6887);
nor U7906 (N_7906,N_7013,N_7099);
nor U7907 (N_7907,N_6755,N_6926);
or U7908 (N_7908,N_7366,N_7093);
nor U7909 (N_7909,N_6776,N_6988);
or U7910 (N_7910,N_6789,N_7304);
nand U7911 (N_7911,N_7393,N_7377);
nor U7912 (N_7912,N_6923,N_7012);
or U7913 (N_7913,N_7062,N_6882);
xor U7914 (N_7914,N_7062,N_7317);
and U7915 (N_7915,N_7442,N_6791);
nand U7916 (N_7916,N_6941,N_6830);
or U7917 (N_7917,N_7303,N_6807);
and U7918 (N_7918,N_6880,N_6906);
and U7919 (N_7919,N_7112,N_6856);
or U7920 (N_7920,N_7466,N_7128);
xnor U7921 (N_7921,N_7416,N_6864);
and U7922 (N_7922,N_7320,N_7328);
xor U7923 (N_7923,N_7044,N_6898);
nand U7924 (N_7924,N_6779,N_7259);
xnor U7925 (N_7925,N_6994,N_7296);
or U7926 (N_7926,N_7127,N_6904);
or U7927 (N_7927,N_6956,N_7355);
or U7928 (N_7928,N_6942,N_7094);
or U7929 (N_7929,N_7077,N_7195);
and U7930 (N_7930,N_7072,N_7075);
nand U7931 (N_7931,N_6966,N_6841);
nand U7932 (N_7932,N_6931,N_6765);
nand U7933 (N_7933,N_6762,N_7482);
nor U7934 (N_7934,N_7241,N_7291);
or U7935 (N_7935,N_7450,N_6968);
and U7936 (N_7936,N_7032,N_6803);
or U7937 (N_7937,N_7263,N_7027);
nor U7938 (N_7938,N_7323,N_7222);
nor U7939 (N_7939,N_7456,N_6864);
and U7940 (N_7940,N_7355,N_7431);
and U7941 (N_7941,N_7423,N_7349);
or U7942 (N_7942,N_6886,N_6887);
or U7943 (N_7943,N_7262,N_6936);
nand U7944 (N_7944,N_7369,N_7144);
nand U7945 (N_7945,N_7114,N_6838);
nand U7946 (N_7946,N_6763,N_6983);
and U7947 (N_7947,N_7331,N_6963);
nand U7948 (N_7948,N_6795,N_7156);
nand U7949 (N_7949,N_6947,N_7179);
nand U7950 (N_7950,N_6834,N_6926);
nand U7951 (N_7951,N_7346,N_7395);
and U7952 (N_7952,N_7235,N_7364);
xnor U7953 (N_7953,N_7478,N_7376);
or U7954 (N_7954,N_7362,N_7345);
and U7955 (N_7955,N_6899,N_7183);
nor U7956 (N_7956,N_7330,N_7490);
xor U7957 (N_7957,N_7114,N_7026);
nand U7958 (N_7958,N_7096,N_6935);
and U7959 (N_7959,N_6864,N_7339);
or U7960 (N_7960,N_6928,N_7452);
nand U7961 (N_7961,N_7092,N_7445);
or U7962 (N_7962,N_7025,N_7019);
or U7963 (N_7963,N_7447,N_7422);
and U7964 (N_7964,N_7058,N_6875);
nor U7965 (N_7965,N_7040,N_7012);
nand U7966 (N_7966,N_7475,N_6924);
xor U7967 (N_7967,N_6778,N_7349);
xnor U7968 (N_7968,N_7142,N_7464);
nand U7969 (N_7969,N_7248,N_6981);
and U7970 (N_7970,N_6862,N_6950);
and U7971 (N_7971,N_6989,N_7321);
xnor U7972 (N_7972,N_6792,N_7474);
and U7973 (N_7973,N_7018,N_7266);
nand U7974 (N_7974,N_7144,N_6810);
or U7975 (N_7975,N_7341,N_7193);
and U7976 (N_7976,N_7001,N_6844);
or U7977 (N_7977,N_7005,N_7231);
and U7978 (N_7978,N_7142,N_7467);
nand U7979 (N_7979,N_7001,N_7182);
nor U7980 (N_7980,N_6756,N_7395);
and U7981 (N_7981,N_6825,N_6838);
xnor U7982 (N_7982,N_7121,N_7196);
xor U7983 (N_7983,N_7011,N_7472);
or U7984 (N_7984,N_7121,N_7266);
or U7985 (N_7985,N_7101,N_6972);
and U7986 (N_7986,N_7401,N_6899);
and U7987 (N_7987,N_7139,N_6907);
xnor U7988 (N_7988,N_7461,N_7092);
and U7989 (N_7989,N_7135,N_6886);
nor U7990 (N_7990,N_7026,N_6969);
or U7991 (N_7991,N_7037,N_7296);
or U7992 (N_7992,N_6915,N_6805);
or U7993 (N_7993,N_7207,N_7143);
or U7994 (N_7994,N_7367,N_7162);
or U7995 (N_7995,N_6941,N_7193);
nor U7996 (N_7996,N_7380,N_7361);
or U7997 (N_7997,N_6863,N_6966);
and U7998 (N_7998,N_7047,N_7326);
nor U7999 (N_7999,N_7417,N_7260);
nand U8000 (N_8000,N_6819,N_7455);
or U8001 (N_8001,N_7366,N_7245);
nand U8002 (N_8002,N_7106,N_7057);
nor U8003 (N_8003,N_7365,N_7249);
nand U8004 (N_8004,N_6902,N_7301);
or U8005 (N_8005,N_7167,N_7234);
or U8006 (N_8006,N_6817,N_7315);
and U8007 (N_8007,N_7066,N_6753);
and U8008 (N_8008,N_6941,N_7476);
nand U8009 (N_8009,N_7234,N_7499);
nor U8010 (N_8010,N_7222,N_6879);
and U8011 (N_8011,N_6891,N_6804);
or U8012 (N_8012,N_7217,N_7014);
or U8013 (N_8013,N_6819,N_7231);
nand U8014 (N_8014,N_7120,N_6750);
and U8015 (N_8015,N_6902,N_6815);
or U8016 (N_8016,N_6991,N_7380);
and U8017 (N_8017,N_7373,N_7366);
and U8018 (N_8018,N_6794,N_7397);
xnor U8019 (N_8019,N_7065,N_7489);
nand U8020 (N_8020,N_7488,N_6780);
nand U8021 (N_8021,N_6901,N_7197);
and U8022 (N_8022,N_6758,N_7021);
or U8023 (N_8023,N_7272,N_7096);
xnor U8024 (N_8024,N_7286,N_7142);
nand U8025 (N_8025,N_6916,N_7362);
nor U8026 (N_8026,N_7117,N_7014);
nand U8027 (N_8027,N_6885,N_7228);
nand U8028 (N_8028,N_6956,N_7498);
nand U8029 (N_8029,N_7245,N_7371);
xnor U8030 (N_8030,N_7486,N_7272);
and U8031 (N_8031,N_7206,N_6762);
or U8032 (N_8032,N_7083,N_7329);
nor U8033 (N_8033,N_7400,N_7204);
and U8034 (N_8034,N_7104,N_7078);
xnor U8035 (N_8035,N_7352,N_7353);
nand U8036 (N_8036,N_7315,N_6823);
nor U8037 (N_8037,N_7101,N_7361);
and U8038 (N_8038,N_7434,N_7450);
and U8039 (N_8039,N_7446,N_6876);
and U8040 (N_8040,N_6995,N_7224);
nand U8041 (N_8041,N_6901,N_7334);
nand U8042 (N_8042,N_7359,N_7339);
nand U8043 (N_8043,N_7428,N_7406);
nand U8044 (N_8044,N_7220,N_6965);
and U8045 (N_8045,N_7230,N_6775);
and U8046 (N_8046,N_7165,N_6903);
nor U8047 (N_8047,N_6889,N_7028);
nand U8048 (N_8048,N_6832,N_7164);
and U8049 (N_8049,N_7042,N_6934);
nor U8050 (N_8050,N_6832,N_6805);
nand U8051 (N_8051,N_7200,N_6978);
and U8052 (N_8052,N_7369,N_7215);
nand U8053 (N_8053,N_7424,N_7303);
xor U8054 (N_8054,N_7047,N_6760);
nor U8055 (N_8055,N_7180,N_6969);
and U8056 (N_8056,N_6865,N_7493);
nand U8057 (N_8057,N_7378,N_7471);
or U8058 (N_8058,N_7133,N_6793);
nand U8059 (N_8059,N_7298,N_7448);
and U8060 (N_8060,N_7406,N_7172);
nand U8061 (N_8061,N_7363,N_6801);
nand U8062 (N_8062,N_6837,N_6763);
nor U8063 (N_8063,N_7245,N_6794);
or U8064 (N_8064,N_6958,N_7191);
nor U8065 (N_8065,N_6798,N_7453);
xnor U8066 (N_8066,N_7350,N_6952);
nor U8067 (N_8067,N_7337,N_7126);
or U8068 (N_8068,N_7187,N_7481);
and U8069 (N_8069,N_6940,N_7055);
nand U8070 (N_8070,N_6883,N_7046);
xnor U8071 (N_8071,N_6803,N_7359);
xnor U8072 (N_8072,N_7400,N_6967);
nand U8073 (N_8073,N_7309,N_6902);
nand U8074 (N_8074,N_6870,N_7259);
or U8075 (N_8075,N_7378,N_6891);
and U8076 (N_8076,N_7308,N_7046);
and U8077 (N_8077,N_7498,N_6830);
xor U8078 (N_8078,N_7084,N_6885);
or U8079 (N_8079,N_6774,N_6970);
or U8080 (N_8080,N_6922,N_7274);
nor U8081 (N_8081,N_7488,N_7232);
or U8082 (N_8082,N_7169,N_7072);
and U8083 (N_8083,N_6845,N_7480);
xnor U8084 (N_8084,N_6750,N_6885);
nor U8085 (N_8085,N_6968,N_7243);
nand U8086 (N_8086,N_6793,N_7467);
or U8087 (N_8087,N_7382,N_7422);
xnor U8088 (N_8088,N_7183,N_6933);
or U8089 (N_8089,N_7162,N_6904);
and U8090 (N_8090,N_6812,N_7075);
and U8091 (N_8091,N_7201,N_7249);
and U8092 (N_8092,N_7474,N_6814);
nand U8093 (N_8093,N_7490,N_7290);
nand U8094 (N_8094,N_7076,N_7054);
or U8095 (N_8095,N_7069,N_6958);
or U8096 (N_8096,N_6957,N_7423);
nor U8097 (N_8097,N_6916,N_6929);
or U8098 (N_8098,N_7466,N_6882);
nand U8099 (N_8099,N_6828,N_7044);
and U8100 (N_8100,N_6980,N_7321);
and U8101 (N_8101,N_7429,N_7120);
or U8102 (N_8102,N_6900,N_6855);
nand U8103 (N_8103,N_7306,N_6955);
and U8104 (N_8104,N_7332,N_6864);
nand U8105 (N_8105,N_6900,N_7251);
nor U8106 (N_8106,N_7118,N_6848);
and U8107 (N_8107,N_6825,N_7238);
and U8108 (N_8108,N_7017,N_6928);
nand U8109 (N_8109,N_7481,N_6771);
and U8110 (N_8110,N_7395,N_6781);
nor U8111 (N_8111,N_7122,N_7465);
and U8112 (N_8112,N_7281,N_7397);
nand U8113 (N_8113,N_6868,N_7415);
or U8114 (N_8114,N_6799,N_6905);
xor U8115 (N_8115,N_7362,N_7390);
nor U8116 (N_8116,N_6861,N_6808);
nor U8117 (N_8117,N_7464,N_6890);
xnor U8118 (N_8118,N_7368,N_6950);
nand U8119 (N_8119,N_6801,N_6882);
xnor U8120 (N_8120,N_7307,N_7282);
xor U8121 (N_8121,N_7165,N_7308);
and U8122 (N_8122,N_6829,N_7111);
and U8123 (N_8123,N_7471,N_6756);
and U8124 (N_8124,N_7205,N_7221);
and U8125 (N_8125,N_7203,N_7406);
and U8126 (N_8126,N_6776,N_7479);
nor U8127 (N_8127,N_7188,N_7240);
nand U8128 (N_8128,N_7059,N_7054);
and U8129 (N_8129,N_6964,N_6923);
nand U8130 (N_8130,N_7160,N_7193);
nor U8131 (N_8131,N_7322,N_7284);
xor U8132 (N_8132,N_7171,N_7285);
nand U8133 (N_8133,N_7239,N_6766);
nor U8134 (N_8134,N_7457,N_6868);
or U8135 (N_8135,N_7076,N_7346);
nand U8136 (N_8136,N_6854,N_7458);
nor U8137 (N_8137,N_7360,N_6998);
nand U8138 (N_8138,N_7204,N_7061);
nand U8139 (N_8139,N_6954,N_7472);
nor U8140 (N_8140,N_7439,N_7070);
or U8141 (N_8141,N_7197,N_7078);
nand U8142 (N_8142,N_6891,N_7135);
or U8143 (N_8143,N_7398,N_6834);
nand U8144 (N_8144,N_7154,N_7160);
nor U8145 (N_8145,N_7462,N_7453);
and U8146 (N_8146,N_7453,N_6996);
xor U8147 (N_8147,N_6765,N_6808);
and U8148 (N_8148,N_6798,N_7349);
and U8149 (N_8149,N_6939,N_7157);
nor U8150 (N_8150,N_7480,N_7304);
nand U8151 (N_8151,N_7310,N_7345);
xnor U8152 (N_8152,N_6754,N_6880);
xnor U8153 (N_8153,N_6939,N_7488);
or U8154 (N_8154,N_7314,N_7167);
nand U8155 (N_8155,N_6752,N_7160);
or U8156 (N_8156,N_7249,N_7215);
xor U8157 (N_8157,N_7284,N_6842);
xnor U8158 (N_8158,N_7310,N_7478);
or U8159 (N_8159,N_7328,N_7351);
nor U8160 (N_8160,N_6763,N_6791);
xor U8161 (N_8161,N_6755,N_7219);
nor U8162 (N_8162,N_7156,N_7410);
or U8163 (N_8163,N_7475,N_7471);
nor U8164 (N_8164,N_6762,N_7159);
nand U8165 (N_8165,N_6949,N_7004);
and U8166 (N_8166,N_7256,N_7444);
or U8167 (N_8167,N_7081,N_6991);
nor U8168 (N_8168,N_7364,N_6801);
or U8169 (N_8169,N_7018,N_7053);
nor U8170 (N_8170,N_7340,N_7025);
or U8171 (N_8171,N_7414,N_7168);
or U8172 (N_8172,N_7437,N_7182);
nor U8173 (N_8173,N_7355,N_6828);
nor U8174 (N_8174,N_7096,N_7494);
or U8175 (N_8175,N_6919,N_7035);
nor U8176 (N_8176,N_7282,N_7229);
and U8177 (N_8177,N_7221,N_7428);
nand U8178 (N_8178,N_7119,N_7030);
nand U8179 (N_8179,N_6798,N_6851);
and U8180 (N_8180,N_6926,N_6859);
nand U8181 (N_8181,N_7253,N_7215);
and U8182 (N_8182,N_7458,N_7472);
and U8183 (N_8183,N_7450,N_6960);
nor U8184 (N_8184,N_7325,N_6938);
or U8185 (N_8185,N_6954,N_6950);
nor U8186 (N_8186,N_7482,N_7110);
and U8187 (N_8187,N_7061,N_7239);
nor U8188 (N_8188,N_7485,N_6907);
and U8189 (N_8189,N_7006,N_6936);
and U8190 (N_8190,N_7462,N_7008);
or U8191 (N_8191,N_7154,N_7139);
nor U8192 (N_8192,N_7175,N_7236);
nand U8193 (N_8193,N_6797,N_6987);
and U8194 (N_8194,N_7466,N_7151);
nand U8195 (N_8195,N_7201,N_6928);
nor U8196 (N_8196,N_6928,N_7004);
nand U8197 (N_8197,N_6907,N_6894);
or U8198 (N_8198,N_7004,N_7285);
and U8199 (N_8199,N_6943,N_6792);
nand U8200 (N_8200,N_7288,N_7035);
or U8201 (N_8201,N_7255,N_7460);
or U8202 (N_8202,N_7315,N_7218);
nor U8203 (N_8203,N_7226,N_7066);
and U8204 (N_8204,N_7171,N_6764);
and U8205 (N_8205,N_7058,N_6969);
nand U8206 (N_8206,N_7156,N_7359);
nor U8207 (N_8207,N_7244,N_7109);
or U8208 (N_8208,N_6985,N_7375);
nand U8209 (N_8209,N_6847,N_6887);
nand U8210 (N_8210,N_7357,N_6967);
and U8211 (N_8211,N_7295,N_6819);
nand U8212 (N_8212,N_7305,N_7307);
nor U8213 (N_8213,N_6815,N_6809);
or U8214 (N_8214,N_7207,N_7491);
nand U8215 (N_8215,N_7267,N_7090);
xor U8216 (N_8216,N_7312,N_7397);
nand U8217 (N_8217,N_7122,N_7114);
nand U8218 (N_8218,N_6966,N_7210);
nor U8219 (N_8219,N_6985,N_7181);
or U8220 (N_8220,N_6835,N_7069);
and U8221 (N_8221,N_7085,N_7446);
nand U8222 (N_8222,N_7033,N_7357);
nor U8223 (N_8223,N_7152,N_7091);
nand U8224 (N_8224,N_7073,N_7407);
or U8225 (N_8225,N_7499,N_7071);
nor U8226 (N_8226,N_7482,N_7361);
nand U8227 (N_8227,N_7382,N_7240);
nand U8228 (N_8228,N_6811,N_6780);
nand U8229 (N_8229,N_6901,N_6760);
or U8230 (N_8230,N_6889,N_7179);
and U8231 (N_8231,N_7254,N_6986);
and U8232 (N_8232,N_6814,N_7340);
nand U8233 (N_8233,N_7421,N_6831);
nor U8234 (N_8234,N_7224,N_6966);
nand U8235 (N_8235,N_7087,N_7236);
and U8236 (N_8236,N_7251,N_6962);
or U8237 (N_8237,N_6851,N_6951);
xor U8238 (N_8238,N_7182,N_6917);
or U8239 (N_8239,N_7093,N_6907);
and U8240 (N_8240,N_7234,N_7031);
and U8241 (N_8241,N_7456,N_6836);
and U8242 (N_8242,N_7291,N_6879);
nor U8243 (N_8243,N_7345,N_6994);
or U8244 (N_8244,N_7377,N_7347);
nand U8245 (N_8245,N_6847,N_7083);
nand U8246 (N_8246,N_6833,N_7418);
or U8247 (N_8247,N_7305,N_7304);
and U8248 (N_8248,N_7005,N_7319);
nor U8249 (N_8249,N_7025,N_6833);
xor U8250 (N_8250,N_7963,N_8197);
xnor U8251 (N_8251,N_7865,N_7795);
nand U8252 (N_8252,N_8102,N_7551);
or U8253 (N_8253,N_8193,N_8070);
nand U8254 (N_8254,N_8135,N_7894);
nor U8255 (N_8255,N_7992,N_8151);
nor U8256 (N_8256,N_7696,N_7820);
xnor U8257 (N_8257,N_7756,N_8202);
nor U8258 (N_8258,N_7919,N_7692);
and U8259 (N_8259,N_7760,N_7782);
and U8260 (N_8260,N_7873,N_8170);
nand U8261 (N_8261,N_7661,N_7931);
and U8262 (N_8262,N_7723,N_7883);
nand U8263 (N_8263,N_8066,N_8038);
or U8264 (N_8264,N_7535,N_7629);
or U8265 (N_8265,N_8163,N_7889);
and U8266 (N_8266,N_7749,N_7779);
or U8267 (N_8267,N_7624,N_8246);
nor U8268 (N_8268,N_8198,N_8090);
or U8269 (N_8269,N_8210,N_8003);
and U8270 (N_8270,N_7801,N_8009);
or U8271 (N_8271,N_7742,N_8116);
or U8272 (N_8272,N_8084,N_7672);
nor U8273 (N_8273,N_7840,N_7577);
nand U8274 (N_8274,N_8051,N_7519);
nor U8275 (N_8275,N_7855,N_7614);
nor U8276 (N_8276,N_7950,N_8013);
nand U8277 (N_8277,N_7677,N_7842);
and U8278 (N_8278,N_7619,N_8074);
and U8279 (N_8279,N_8027,N_7556);
xnor U8280 (N_8280,N_7606,N_7566);
nor U8281 (N_8281,N_7562,N_7632);
nand U8282 (N_8282,N_7526,N_7622);
nand U8283 (N_8283,N_7508,N_7648);
nand U8284 (N_8284,N_7985,N_7949);
xnor U8285 (N_8285,N_8219,N_7937);
nand U8286 (N_8286,N_8049,N_8120);
or U8287 (N_8287,N_7633,N_7991);
or U8288 (N_8288,N_7559,N_8212);
nor U8289 (N_8289,N_7687,N_8171);
and U8290 (N_8290,N_8002,N_7878);
nor U8291 (N_8291,N_8187,N_7858);
nand U8292 (N_8292,N_7800,N_8065);
and U8293 (N_8293,N_7954,N_7918);
or U8294 (N_8294,N_7595,N_7706);
and U8295 (N_8295,N_8149,N_7603);
or U8296 (N_8296,N_7515,N_8091);
or U8297 (N_8297,N_8112,N_7784);
or U8298 (N_8298,N_8180,N_8182);
nor U8299 (N_8299,N_7589,N_8006);
nor U8300 (N_8300,N_8078,N_7912);
and U8301 (N_8301,N_7695,N_7665);
or U8302 (N_8302,N_7882,N_7935);
and U8303 (N_8303,N_8014,N_7529);
nor U8304 (N_8304,N_7952,N_8114);
or U8305 (N_8305,N_8201,N_7591);
or U8306 (N_8306,N_7817,N_7792);
and U8307 (N_8307,N_8162,N_7793);
nor U8308 (N_8308,N_7543,N_7905);
nor U8309 (N_8309,N_8101,N_8016);
nand U8310 (N_8310,N_8008,N_8139);
nor U8311 (N_8311,N_7707,N_8123);
nand U8312 (N_8312,N_7890,N_8222);
or U8313 (N_8313,N_8045,N_7576);
nor U8314 (N_8314,N_8068,N_7548);
nand U8315 (N_8315,N_8158,N_8209);
xnor U8316 (N_8316,N_8073,N_8096);
or U8317 (N_8317,N_7970,N_8040);
or U8318 (N_8318,N_7995,N_7829);
nand U8319 (N_8319,N_7989,N_7537);
nand U8320 (N_8320,N_8143,N_7788);
or U8321 (N_8321,N_8213,N_8098);
nor U8322 (N_8322,N_8075,N_7722);
nand U8323 (N_8323,N_7976,N_8233);
nor U8324 (N_8324,N_7901,N_7521);
and U8325 (N_8325,N_8226,N_8001);
and U8326 (N_8326,N_8230,N_8062);
or U8327 (N_8327,N_7634,N_7744);
or U8328 (N_8328,N_7850,N_8224);
nor U8329 (N_8329,N_7763,N_7567);
or U8330 (N_8330,N_7520,N_8111);
nor U8331 (N_8331,N_7814,N_8020);
nand U8332 (N_8332,N_7874,N_7533);
or U8333 (N_8333,N_7859,N_8173);
nand U8334 (N_8334,N_8137,N_7982);
and U8335 (N_8335,N_8227,N_8134);
nor U8336 (N_8336,N_7825,N_7839);
or U8337 (N_8337,N_8059,N_7563);
nand U8338 (N_8338,N_8154,N_8247);
nand U8339 (N_8339,N_7538,N_7908);
nand U8340 (N_8340,N_7765,N_7694);
and U8341 (N_8341,N_8105,N_8211);
xor U8342 (N_8342,N_7539,N_7588);
or U8343 (N_8343,N_7900,N_8196);
or U8344 (N_8344,N_7510,N_8144);
nand U8345 (N_8345,N_7868,N_7586);
nand U8346 (N_8346,N_7846,N_7754);
xnor U8347 (N_8347,N_7869,N_7953);
nor U8348 (N_8348,N_7804,N_7827);
xor U8349 (N_8349,N_7778,N_7776);
or U8350 (N_8350,N_7861,N_7922);
or U8351 (N_8351,N_8189,N_7896);
nor U8352 (N_8352,N_7994,N_7546);
and U8353 (N_8353,N_7964,N_7828);
or U8354 (N_8354,N_7715,N_8086);
and U8355 (N_8355,N_7862,N_7888);
and U8356 (N_8356,N_7810,N_8136);
xor U8357 (N_8357,N_7596,N_7643);
nor U8358 (N_8358,N_8216,N_7848);
nand U8359 (N_8359,N_7913,N_7818);
nor U8360 (N_8360,N_8044,N_7892);
and U8361 (N_8361,N_7791,N_7711);
and U8362 (N_8362,N_7833,N_8005);
nor U8363 (N_8363,N_7613,N_8155);
and U8364 (N_8364,N_7960,N_8035);
nor U8365 (N_8365,N_7679,N_7772);
nand U8366 (N_8366,N_7803,N_7587);
nor U8367 (N_8367,N_7944,N_7738);
or U8368 (N_8368,N_8050,N_7977);
nor U8369 (N_8369,N_7652,N_8199);
nor U8370 (N_8370,N_8053,N_8106);
or U8371 (N_8371,N_8025,N_7719);
or U8372 (N_8372,N_8220,N_7579);
nor U8373 (N_8373,N_7518,N_7501);
nor U8374 (N_8374,N_7700,N_7623);
nor U8375 (N_8375,N_7550,N_8063);
nor U8376 (N_8376,N_8099,N_7545);
or U8377 (N_8377,N_7747,N_8019);
or U8378 (N_8378,N_7794,N_7555);
nor U8379 (N_8379,N_7815,N_7647);
or U8380 (N_8380,N_7787,N_7656);
nor U8381 (N_8381,N_7955,N_7986);
or U8382 (N_8382,N_8153,N_7993);
nor U8383 (N_8383,N_7712,N_8249);
nor U8384 (N_8384,N_7728,N_8054);
nand U8385 (N_8385,N_8110,N_7662);
nor U8386 (N_8386,N_7998,N_7832);
nand U8387 (N_8387,N_8118,N_7564);
or U8388 (N_8388,N_8089,N_8010);
and U8389 (N_8389,N_7867,N_7920);
or U8390 (N_8390,N_7798,N_8129);
and U8391 (N_8391,N_7565,N_7973);
nand U8392 (N_8392,N_8192,N_7852);
or U8393 (N_8393,N_8125,N_7940);
and U8394 (N_8394,N_7531,N_8085);
nor U8395 (N_8395,N_7724,N_8043);
or U8396 (N_8396,N_8057,N_7698);
xor U8397 (N_8397,N_7664,N_8121);
xnor U8398 (N_8398,N_7681,N_7831);
and U8399 (N_8399,N_8093,N_8113);
nor U8400 (N_8400,N_7945,N_7968);
and U8401 (N_8401,N_7758,N_7618);
or U8402 (N_8402,N_7860,N_7797);
nand U8403 (N_8403,N_7605,N_7886);
nand U8404 (N_8404,N_8244,N_8150);
nor U8405 (N_8405,N_8072,N_7513);
or U8406 (N_8406,N_7512,N_7733);
and U8407 (N_8407,N_7522,N_8164);
nor U8408 (N_8408,N_7561,N_7974);
nor U8409 (N_8409,N_7654,N_7528);
xnor U8410 (N_8410,N_7872,N_8235);
or U8411 (N_8411,N_7688,N_7957);
xnor U8412 (N_8412,N_7752,N_7607);
xor U8413 (N_8413,N_7547,N_8083);
and U8414 (N_8414,N_7708,N_7525);
xnor U8415 (N_8415,N_7777,N_7939);
nor U8416 (N_8416,N_7673,N_7731);
or U8417 (N_8417,N_7783,N_8022);
nand U8418 (N_8418,N_8061,N_7870);
nor U8419 (N_8419,N_7650,N_7796);
and U8420 (N_8420,N_8087,N_7500);
nand U8421 (N_8421,N_7927,N_7536);
or U8422 (N_8422,N_7549,N_7785);
nand U8423 (N_8423,N_7568,N_7844);
nor U8424 (N_8424,N_7903,N_7714);
or U8425 (N_8425,N_7693,N_7880);
and U8426 (N_8426,N_7612,N_7925);
and U8427 (N_8427,N_7946,N_7930);
nand U8428 (N_8428,N_7737,N_8141);
nor U8429 (N_8429,N_7646,N_7504);
nor U8430 (N_8430,N_8152,N_7864);
nand U8431 (N_8431,N_7572,N_7685);
or U8432 (N_8432,N_7990,N_7630);
nand U8433 (N_8433,N_7574,N_8168);
nor U8434 (N_8434,N_7773,N_7530);
or U8435 (N_8435,N_8228,N_7909);
and U8436 (N_8436,N_7583,N_7740);
and U8437 (N_8437,N_7759,N_8071);
xnor U8438 (N_8438,N_8131,N_8119);
nor U8439 (N_8439,N_7610,N_8145);
nor U8440 (N_8440,N_7999,N_7819);
nor U8441 (N_8441,N_8240,N_7780);
and U8442 (N_8442,N_7808,N_8148);
nand U8443 (N_8443,N_8094,N_7902);
or U8444 (N_8444,N_8109,N_8024);
nor U8445 (N_8445,N_7716,N_7769);
nor U8446 (N_8446,N_7802,N_7657);
xnor U8447 (N_8447,N_8183,N_7721);
and U8448 (N_8448,N_7812,N_8077);
nor U8449 (N_8449,N_7557,N_8241);
nand U8450 (N_8450,N_8195,N_8181);
and U8451 (N_8451,N_7996,N_7635);
xor U8452 (N_8452,N_7703,N_7626);
nand U8453 (N_8453,N_8214,N_7961);
or U8454 (N_8454,N_8076,N_7891);
nor U8455 (N_8455,N_7628,N_8052);
nor U8456 (N_8456,N_7600,N_8012);
and U8457 (N_8457,N_7604,N_7534);
nor U8458 (N_8458,N_7942,N_7581);
xor U8459 (N_8459,N_8229,N_7962);
or U8460 (N_8460,N_7933,N_7898);
and U8461 (N_8461,N_7938,N_8069);
and U8462 (N_8462,N_8004,N_7674);
or U8463 (N_8463,N_8200,N_7569);
nand U8464 (N_8464,N_8215,N_8174);
nor U8465 (N_8465,N_7746,N_8081);
nand U8466 (N_8466,N_7910,N_8048);
and U8467 (N_8467,N_7897,N_8056);
nor U8468 (N_8468,N_8232,N_7841);
nand U8469 (N_8469,N_8100,N_8021);
nand U8470 (N_8470,N_8217,N_8178);
or U8471 (N_8471,N_7699,N_7836);
or U8472 (N_8472,N_8184,N_7823);
or U8473 (N_8473,N_8218,N_8206);
or U8474 (N_8474,N_7751,N_7638);
xnor U8475 (N_8475,N_7690,N_8029);
nor U8476 (N_8476,N_8132,N_7729);
nand U8477 (N_8477,N_7834,N_7771);
and U8478 (N_8478,N_7975,N_8169);
or U8479 (N_8479,N_7697,N_7669);
nor U8480 (N_8480,N_8231,N_7851);
nor U8481 (N_8481,N_7959,N_8046);
and U8482 (N_8482,N_7762,N_8166);
or U8483 (N_8483,N_8064,N_7843);
nand U8484 (N_8484,N_7578,N_7757);
or U8485 (N_8485,N_8037,N_8140);
xor U8486 (N_8486,N_8128,N_8042);
nor U8487 (N_8487,N_7552,N_7866);
and U8488 (N_8488,N_7683,N_8221);
nand U8489 (N_8489,N_7764,N_7884);
or U8490 (N_8490,N_7593,N_7667);
xnor U8491 (N_8491,N_7824,N_8034);
and U8492 (N_8492,N_7936,N_8124);
nand U8493 (N_8493,N_7921,N_7658);
xnor U8494 (N_8494,N_7987,N_7702);
and U8495 (N_8495,N_7854,N_7725);
nor U8496 (N_8496,N_8203,N_7932);
and U8497 (N_8497,N_7570,N_7617);
or U8498 (N_8498,N_8242,N_7571);
and U8499 (N_8499,N_7666,N_7822);
and U8500 (N_8500,N_7659,N_7680);
nor U8501 (N_8501,N_7809,N_7701);
nand U8502 (N_8502,N_8165,N_7911);
and U8503 (N_8503,N_7620,N_7582);
nand U8504 (N_8504,N_7966,N_8107);
nor U8505 (N_8505,N_8234,N_7718);
nand U8506 (N_8506,N_7503,N_7806);
and U8507 (N_8507,N_7726,N_7713);
or U8508 (N_8508,N_8033,N_7653);
nor U8509 (N_8509,N_7790,N_7743);
xor U8510 (N_8510,N_7830,N_8156);
nor U8511 (N_8511,N_7736,N_7934);
nand U8512 (N_8512,N_8122,N_7660);
and U8513 (N_8513,N_7984,N_7789);
or U8514 (N_8514,N_7527,N_8138);
or U8515 (N_8515,N_7615,N_7732);
nand U8516 (N_8516,N_7691,N_8167);
or U8517 (N_8517,N_7745,N_7641);
nand U8518 (N_8518,N_7983,N_7770);
nand U8519 (N_8519,N_8194,N_7849);
and U8520 (N_8520,N_7580,N_8060);
or U8521 (N_8521,N_7906,N_7877);
nor U8522 (N_8522,N_7924,N_7717);
and U8523 (N_8523,N_7835,N_8157);
or U8524 (N_8524,N_8204,N_7923);
or U8525 (N_8525,N_7705,N_7967);
nand U8526 (N_8526,N_7649,N_8092);
nor U8527 (N_8527,N_7871,N_7767);
or U8528 (N_8528,N_8097,N_7709);
nand U8529 (N_8529,N_7904,N_8236);
nand U8530 (N_8530,N_8205,N_7948);
xor U8531 (N_8531,N_7676,N_7544);
nand U8532 (N_8532,N_8115,N_7997);
and U8533 (N_8533,N_8245,N_7826);
or U8534 (N_8534,N_7766,N_7730);
or U8535 (N_8535,N_8055,N_7926);
and U8536 (N_8536,N_7821,N_7917);
or U8537 (N_8537,N_7636,N_8047);
nand U8538 (N_8538,N_7863,N_7799);
nor U8539 (N_8539,N_8108,N_7507);
nor U8540 (N_8540,N_8179,N_7644);
or U8541 (N_8541,N_8036,N_7813);
nor U8542 (N_8542,N_8007,N_7558);
nand U8543 (N_8543,N_7502,N_8238);
nor U8544 (N_8544,N_8223,N_7958);
or U8545 (N_8545,N_8104,N_8175);
or U8546 (N_8546,N_7682,N_7811);
nor U8547 (N_8547,N_7590,N_7734);
and U8548 (N_8548,N_7592,N_7875);
xor U8549 (N_8549,N_7601,N_7585);
nand U8550 (N_8550,N_8058,N_7684);
nor U8551 (N_8551,N_8133,N_8207);
or U8552 (N_8552,N_8185,N_8082);
nand U8553 (N_8553,N_8095,N_7514);
nand U8554 (N_8554,N_8041,N_8237);
or U8555 (N_8555,N_7720,N_7663);
xor U8556 (N_8556,N_7879,N_7602);
xor U8557 (N_8557,N_7943,N_7837);
and U8558 (N_8558,N_7786,N_7838);
nor U8559 (N_8559,N_8142,N_8103);
xor U8560 (N_8560,N_7505,N_7907);
and U8561 (N_8561,N_8000,N_7542);
nand U8562 (N_8562,N_8130,N_7978);
nand U8563 (N_8563,N_7847,N_7853);
and U8564 (N_8564,N_7972,N_7775);
and U8565 (N_8565,N_7554,N_7640);
xnor U8566 (N_8566,N_8030,N_8079);
and U8567 (N_8567,N_7753,N_8015);
or U8568 (N_8568,N_8191,N_7857);
nand U8569 (N_8569,N_7980,N_7584);
xnor U8570 (N_8570,N_7748,N_7689);
or U8571 (N_8571,N_8080,N_7651);
or U8572 (N_8572,N_7807,N_8188);
or U8573 (N_8573,N_7637,N_7727);
nand U8574 (N_8574,N_8088,N_7541);
nor U8575 (N_8575,N_7941,N_7971);
xor U8576 (N_8576,N_8225,N_7928);
or U8577 (N_8577,N_7951,N_7881);
xnor U8578 (N_8578,N_7627,N_7670);
and U8579 (N_8579,N_7616,N_8039);
and U8580 (N_8580,N_7781,N_7671);
and U8581 (N_8581,N_7675,N_7540);
nand U8582 (N_8582,N_7710,N_8159);
and U8583 (N_8583,N_8023,N_8172);
or U8584 (N_8584,N_7739,N_7678);
and U8585 (N_8585,N_8208,N_7553);
nand U8586 (N_8586,N_7965,N_7741);
and U8587 (N_8587,N_8031,N_8186);
nor U8588 (N_8588,N_8147,N_7524);
xnor U8589 (N_8589,N_7845,N_7621);
or U8590 (N_8590,N_7611,N_8243);
and U8591 (N_8591,N_8127,N_7599);
nand U8592 (N_8592,N_7517,N_8026);
and U8593 (N_8593,N_7668,N_7750);
or U8594 (N_8594,N_7774,N_8177);
and U8595 (N_8595,N_7885,N_8067);
nand U8596 (N_8596,N_7704,N_8160);
nor U8597 (N_8597,N_7876,N_7893);
and U8598 (N_8598,N_7856,N_8018);
and U8599 (N_8599,N_7645,N_7915);
or U8600 (N_8600,N_7895,N_8176);
and U8601 (N_8601,N_7532,N_8126);
xor U8602 (N_8602,N_7768,N_7969);
nor U8603 (N_8603,N_7598,N_7631);
nand U8604 (N_8604,N_7686,N_7597);
xor U8605 (N_8605,N_7575,N_7979);
or U8606 (N_8606,N_7642,N_8117);
nand U8607 (N_8607,N_8032,N_7947);
or U8608 (N_8608,N_7816,N_7560);
and U8609 (N_8609,N_7761,N_7625);
nor U8610 (N_8610,N_7755,N_7608);
xnor U8611 (N_8611,N_7981,N_7916);
or U8612 (N_8612,N_7609,N_7594);
and U8613 (N_8613,N_8017,N_7573);
nand U8614 (N_8614,N_8146,N_7735);
or U8615 (N_8615,N_7956,N_7506);
and U8616 (N_8616,N_8161,N_7523);
and U8617 (N_8617,N_8239,N_7988);
nand U8618 (N_8618,N_7511,N_7516);
and U8619 (N_8619,N_7655,N_8190);
xnor U8620 (N_8620,N_7929,N_7509);
or U8621 (N_8621,N_7805,N_8248);
and U8622 (N_8622,N_7639,N_7914);
or U8623 (N_8623,N_8011,N_7899);
and U8624 (N_8624,N_7887,N_8028);
nand U8625 (N_8625,N_7971,N_7813);
or U8626 (N_8626,N_8039,N_7824);
and U8627 (N_8627,N_7711,N_8091);
nor U8628 (N_8628,N_8079,N_7889);
nand U8629 (N_8629,N_7631,N_8206);
or U8630 (N_8630,N_8042,N_7719);
nand U8631 (N_8631,N_7545,N_8182);
nor U8632 (N_8632,N_8142,N_7579);
nor U8633 (N_8633,N_8006,N_8162);
xnor U8634 (N_8634,N_7584,N_7918);
and U8635 (N_8635,N_7956,N_7662);
xor U8636 (N_8636,N_8230,N_7671);
xor U8637 (N_8637,N_8204,N_7908);
nor U8638 (N_8638,N_7622,N_8212);
or U8639 (N_8639,N_7634,N_7674);
and U8640 (N_8640,N_8144,N_7575);
nor U8641 (N_8641,N_8031,N_7641);
or U8642 (N_8642,N_7964,N_7690);
and U8643 (N_8643,N_8170,N_7560);
nand U8644 (N_8644,N_8115,N_7902);
nor U8645 (N_8645,N_8124,N_7894);
and U8646 (N_8646,N_7877,N_7903);
nor U8647 (N_8647,N_8185,N_7709);
nor U8648 (N_8648,N_7968,N_8242);
xor U8649 (N_8649,N_7500,N_7915);
or U8650 (N_8650,N_7605,N_7867);
xnor U8651 (N_8651,N_8083,N_7535);
xor U8652 (N_8652,N_8130,N_8011);
nor U8653 (N_8653,N_8077,N_7776);
or U8654 (N_8654,N_7715,N_7976);
and U8655 (N_8655,N_7548,N_7885);
nor U8656 (N_8656,N_7945,N_7569);
or U8657 (N_8657,N_7830,N_7621);
xnor U8658 (N_8658,N_7806,N_7523);
or U8659 (N_8659,N_8130,N_7688);
nand U8660 (N_8660,N_7868,N_8039);
nor U8661 (N_8661,N_8242,N_7576);
nor U8662 (N_8662,N_7599,N_7867);
nand U8663 (N_8663,N_7767,N_7595);
or U8664 (N_8664,N_7753,N_8049);
and U8665 (N_8665,N_7924,N_7730);
and U8666 (N_8666,N_7710,N_8015);
nor U8667 (N_8667,N_8029,N_7935);
xor U8668 (N_8668,N_8230,N_7568);
and U8669 (N_8669,N_7613,N_8015);
nand U8670 (N_8670,N_7665,N_8156);
xnor U8671 (N_8671,N_7848,N_8077);
or U8672 (N_8672,N_7941,N_7562);
nand U8673 (N_8673,N_7966,N_7752);
nand U8674 (N_8674,N_7838,N_7898);
and U8675 (N_8675,N_7614,N_7964);
nand U8676 (N_8676,N_8159,N_7980);
nand U8677 (N_8677,N_7820,N_7778);
nand U8678 (N_8678,N_7720,N_7582);
nand U8679 (N_8679,N_7511,N_8076);
and U8680 (N_8680,N_7547,N_7542);
xor U8681 (N_8681,N_7513,N_7944);
or U8682 (N_8682,N_8112,N_7730);
and U8683 (N_8683,N_7726,N_7589);
xnor U8684 (N_8684,N_7659,N_8188);
or U8685 (N_8685,N_7698,N_8004);
nor U8686 (N_8686,N_8163,N_8128);
and U8687 (N_8687,N_7518,N_7756);
nand U8688 (N_8688,N_8148,N_7824);
nor U8689 (N_8689,N_7721,N_8221);
nand U8690 (N_8690,N_7666,N_7975);
nor U8691 (N_8691,N_7657,N_7634);
and U8692 (N_8692,N_7833,N_7616);
nand U8693 (N_8693,N_8226,N_7726);
or U8694 (N_8694,N_7872,N_8216);
nand U8695 (N_8695,N_8174,N_7937);
or U8696 (N_8696,N_7597,N_8020);
nor U8697 (N_8697,N_7648,N_7641);
and U8698 (N_8698,N_8070,N_7611);
nand U8699 (N_8699,N_7592,N_7754);
nor U8700 (N_8700,N_7753,N_7577);
or U8701 (N_8701,N_7577,N_7872);
nand U8702 (N_8702,N_7845,N_7695);
nor U8703 (N_8703,N_7644,N_8022);
and U8704 (N_8704,N_7942,N_8012);
xor U8705 (N_8705,N_7573,N_7857);
and U8706 (N_8706,N_7628,N_7901);
nand U8707 (N_8707,N_7843,N_7794);
and U8708 (N_8708,N_7532,N_7937);
or U8709 (N_8709,N_7652,N_7530);
and U8710 (N_8710,N_7733,N_7526);
nor U8711 (N_8711,N_7776,N_8210);
or U8712 (N_8712,N_7701,N_7514);
nor U8713 (N_8713,N_8215,N_8120);
and U8714 (N_8714,N_7796,N_7941);
or U8715 (N_8715,N_7908,N_7791);
and U8716 (N_8716,N_7534,N_8024);
nand U8717 (N_8717,N_8144,N_8101);
or U8718 (N_8718,N_7751,N_7741);
nor U8719 (N_8719,N_7672,N_7654);
or U8720 (N_8720,N_7513,N_8113);
or U8721 (N_8721,N_7582,N_8155);
nor U8722 (N_8722,N_7749,N_7647);
nand U8723 (N_8723,N_7826,N_7878);
xnor U8724 (N_8724,N_7554,N_7699);
and U8725 (N_8725,N_8027,N_8147);
or U8726 (N_8726,N_8224,N_7865);
nor U8727 (N_8727,N_7692,N_7567);
xor U8728 (N_8728,N_7621,N_8053);
nand U8729 (N_8729,N_7962,N_7831);
or U8730 (N_8730,N_7738,N_7872);
nand U8731 (N_8731,N_7881,N_7821);
nor U8732 (N_8732,N_7703,N_8148);
or U8733 (N_8733,N_8197,N_7766);
and U8734 (N_8734,N_7871,N_8090);
or U8735 (N_8735,N_8036,N_7868);
or U8736 (N_8736,N_7642,N_8018);
and U8737 (N_8737,N_7501,N_7572);
nor U8738 (N_8738,N_8160,N_7962);
or U8739 (N_8739,N_8052,N_8032);
nand U8740 (N_8740,N_8235,N_7519);
or U8741 (N_8741,N_7658,N_8215);
xor U8742 (N_8742,N_7789,N_8065);
nand U8743 (N_8743,N_7817,N_7875);
and U8744 (N_8744,N_8145,N_7688);
and U8745 (N_8745,N_8233,N_7686);
or U8746 (N_8746,N_7778,N_8006);
nand U8747 (N_8747,N_7511,N_8214);
and U8748 (N_8748,N_7816,N_7826);
and U8749 (N_8749,N_7873,N_7888);
nor U8750 (N_8750,N_7915,N_7755);
nor U8751 (N_8751,N_8236,N_8111);
or U8752 (N_8752,N_7809,N_8000);
or U8753 (N_8753,N_8118,N_7750);
nor U8754 (N_8754,N_8179,N_8227);
or U8755 (N_8755,N_7951,N_7667);
and U8756 (N_8756,N_7693,N_8238);
nand U8757 (N_8757,N_7982,N_8117);
nand U8758 (N_8758,N_7534,N_8072);
xor U8759 (N_8759,N_7798,N_8060);
and U8760 (N_8760,N_8044,N_7578);
or U8761 (N_8761,N_7537,N_7611);
nor U8762 (N_8762,N_8215,N_7716);
or U8763 (N_8763,N_7569,N_7941);
nand U8764 (N_8764,N_7519,N_7751);
xor U8765 (N_8765,N_8188,N_7978);
nand U8766 (N_8766,N_7766,N_7915);
or U8767 (N_8767,N_7987,N_8209);
and U8768 (N_8768,N_7640,N_8095);
or U8769 (N_8769,N_7752,N_8197);
nand U8770 (N_8770,N_7644,N_7891);
or U8771 (N_8771,N_7999,N_7550);
nor U8772 (N_8772,N_7730,N_8165);
or U8773 (N_8773,N_7743,N_7897);
and U8774 (N_8774,N_8069,N_7944);
or U8775 (N_8775,N_7616,N_8027);
and U8776 (N_8776,N_7950,N_8222);
or U8777 (N_8777,N_8214,N_8108);
and U8778 (N_8778,N_7848,N_8231);
nand U8779 (N_8779,N_8111,N_8177);
xor U8780 (N_8780,N_7866,N_7549);
or U8781 (N_8781,N_7585,N_8049);
nand U8782 (N_8782,N_7784,N_7689);
nand U8783 (N_8783,N_8237,N_8066);
nand U8784 (N_8784,N_7650,N_8087);
nand U8785 (N_8785,N_8246,N_7914);
nand U8786 (N_8786,N_7758,N_8225);
nor U8787 (N_8787,N_7892,N_7800);
nand U8788 (N_8788,N_8225,N_8190);
nand U8789 (N_8789,N_7745,N_7818);
xnor U8790 (N_8790,N_7800,N_7926);
nor U8791 (N_8791,N_7787,N_7590);
or U8792 (N_8792,N_7862,N_7689);
and U8793 (N_8793,N_7855,N_7551);
and U8794 (N_8794,N_7845,N_8210);
or U8795 (N_8795,N_7864,N_7861);
nand U8796 (N_8796,N_8065,N_7919);
nor U8797 (N_8797,N_7979,N_7626);
and U8798 (N_8798,N_7580,N_7503);
nor U8799 (N_8799,N_7526,N_7748);
nand U8800 (N_8800,N_8123,N_7899);
and U8801 (N_8801,N_7813,N_7521);
and U8802 (N_8802,N_8117,N_7829);
and U8803 (N_8803,N_7916,N_7667);
nand U8804 (N_8804,N_7660,N_7858);
nand U8805 (N_8805,N_8057,N_7814);
nand U8806 (N_8806,N_7662,N_8044);
and U8807 (N_8807,N_8185,N_7932);
or U8808 (N_8808,N_7557,N_7879);
nor U8809 (N_8809,N_7629,N_7947);
nand U8810 (N_8810,N_7574,N_8244);
or U8811 (N_8811,N_8037,N_7943);
and U8812 (N_8812,N_8246,N_8044);
xnor U8813 (N_8813,N_7897,N_7921);
xor U8814 (N_8814,N_7763,N_8160);
nor U8815 (N_8815,N_7584,N_7810);
nor U8816 (N_8816,N_7548,N_8091);
nand U8817 (N_8817,N_7655,N_7795);
nor U8818 (N_8818,N_7938,N_8157);
nand U8819 (N_8819,N_7629,N_8241);
xor U8820 (N_8820,N_8014,N_7879);
nand U8821 (N_8821,N_8117,N_7912);
and U8822 (N_8822,N_7992,N_8050);
and U8823 (N_8823,N_7829,N_7800);
and U8824 (N_8824,N_8030,N_8031);
or U8825 (N_8825,N_8238,N_7760);
or U8826 (N_8826,N_7658,N_8126);
and U8827 (N_8827,N_7951,N_7690);
and U8828 (N_8828,N_8200,N_8004);
and U8829 (N_8829,N_7970,N_7549);
nand U8830 (N_8830,N_7911,N_7633);
nand U8831 (N_8831,N_8038,N_7722);
and U8832 (N_8832,N_7524,N_8047);
nand U8833 (N_8833,N_7919,N_7997);
and U8834 (N_8834,N_7894,N_8238);
and U8835 (N_8835,N_7676,N_7889);
nand U8836 (N_8836,N_7685,N_8025);
xnor U8837 (N_8837,N_7926,N_8132);
nor U8838 (N_8838,N_7632,N_7725);
xor U8839 (N_8839,N_8175,N_7581);
nand U8840 (N_8840,N_7952,N_7574);
and U8841 (N_8841,N_7832,N_7654);
or U8842 (N_8842,N_8036,N_7693);
nand U8843 (N_8843,N_8080,N_7836);
nor U8844 (N_8844,N_8055,N_8099);
and U8845 (N_8845,N_8166,N_7730);
nor U8846 (N_8846,N_7806,N_7899);
nand U8847 (N_8847,N_7897,N_8193);
xor U8848 (N_8848,N_8225,N_7976);
and U8849 (N_8849,N_8104,N_7678);
nand U8850 (N_8850,N_8209,N_8122);
xnor U8851 (N_8851,N_7579,N_8066);
and U8852 (N_8852,N_7980,N_7704);
nand U8853 (N_8853,N_7841,N_8078);
nand U8854 (N_8854,N_7563,N_8203);
and U8855 (N_8855,N_7582,N_7952);
nand U8856 (N_8856,N_8118,N_7588);
xnor U8857 (N_8857,N_7812,N_7796);
nor U8858 (N_8858,N_8007,N_7915);
and U8859 (N_8859,N_8198,N_7954);
or U8860 (N_8860,N_7978,N_8049);
nor U8861 (N_8861,N_7715,N_7687);
or U8862 (N_8862,N_7782,N_8182);
nand U8863 (N_8863,N_8187,N_7874);
or U8864 (N_8864,N_8244,N_7741);
nor U8865 (N_8865,N_8206,N_7705);
nor U8866 (N_8866,N_7778,N_8116);
nand U8867 (N_8867,N_7730,N_8196);
nand U8868 (N_8868,N_7535,N_7503);
or U8869 (N_8869,N_7637,N_7603);
nand U8870 (N_8870,N_7973,N_8143);
nor U8871 (N_8871,N_7553,N_7841);
nor U8872 (N_8872,N_8027,N_7971);
xor U8873 (N_8873,N_7593,N_8125);
nand U8874 (N_8874,N_7842,N_8157);
nand U8875 (N_8875,N_7924,N_7701);
or U8876 (N_8876,N_7703,N_8072);
or U8877 (N_8877,N_7970,N_7954);
nand U8878 (N_8878,N_7865,N_7571);
xnor U8879 (N_8879,N_8118,N_7551);
or U8880 (N_8880,N_7857,N_8069);
or U8881 (N_8881,N_8046,N_7800);
nand U8882 (N_8882,N_8114,N_7508);
and U8883 (N_8883,N_7952,N_7942);
xor U8884 (N_8884,N_7724,N_7716);
xnor U8885 (N_8885,N_8050,N_7779);
nand U8886 (N_8886,N_7563,N_7582);
nand U8887 (N_8887,N_7873,N_7655);
and U8888 (N_8888,N_8119,N_7937);
nor U8889 (N_8889,N_7919,N_7770);
and U8890 (N_8890,N_7555,N_8202);
nand U8891 (N_8891,N_8048,N_7538);
nor U8892 (N_8892,N_7637,N_7509);
and U8893 (N_8893,N_8049,N_7635);
nand U8894 (N_8894,N_8007,N_8137);
nand U8895 (N_8895,N_8133,N_7508);
and U8896 (N_8896,N_7818,N_8062);
nand U8897 (N_8897,N_7567,N_7722);
nand U8898 (N_8898,N_7744,N_8245);
and U8899 (N_8899,N_7549,N_8084);
and U8900 (N_8900,N_8043,N_7871);
xor U8901 (N_8901,N_7959,N_8059);
nor U8902 (N_8902,N_7822,N_7869);
or U8903 (N_8903,N_8121,N_7692);
or U8904 (N_8904,N_7882,N_8034);
nand U8905 (N_8905,N_8036,N_8156);
or U8906 (N_8906,N_7947,N_8184);
nor U8907 (N_8907,N_7919,N_7816);
nand U8908 (N_8908,N_7560,N_7540);
nor U8909 (N_8909,N_7969,N_8159);
xor U8910 (N_8910,N_7733,N_8200);
and U8911 (N_8911,N_7501,N_8233);
xor U8912 (N_8912,N_7549,N_7992);
nor U8913 (N_8913,N_7662,N_7912);
or U8914 (N_8914,N_8100,N_7608);
nor U8915 (N_8915,N_7587,N_8055);
and U8916 (N_8916,N_8072,N_8026);
nor U8917 (N_8917,N_7682,N_8104);
nand U8918 (N_8918,N_7519,N_7633);
or U8919 (N_8919,N_8131,N_7925);
or U8920 (N_8920,N_7549,N_7742);
nor U8921 (N_8921,N_7802,N_8181);
or U8922 (N_8922,N_7722,N_7612);
nor U8923 (N_8923,N_7729,N_8218);
nor U8924 (N_8924,N_8054,N_7694);
and U8925 (N_8925,N_8043,N_7814);
nor U8926 (N_8926,N_8019,N_7602);
and U8927 (N_8927,N_8209,N_7690);
xnor U8928 (N_8928,N_7748,N_7739);
nand U8929 (N_8929,N_8207,N_8140);
xor U8930 (N_8930,N_7646,N_7983);
and U8931 (N_8931,N_7982,N_7614);
nand U8932 (N_8932,N_7528,N_7776);
nand U8933 (N_8933,N_7644,N_8129);
nand U8934 (N_8934,N_7820,N_7981);
nor U8935 (N_8935,N_7913,N_7698);
nor U8936 (N_8936,N_8099,N_7542);
nor U8937 (N_8937,N_7903,N_8190);
and U8938 (N_8938,N_7695,N_8047);
or U8939 (N_8939,N_7791,N_8045);
and U8940 (N_8940,N_7930,N_7705);
nand U8941 (N_8941,N_8053,N_7633);
and U8942 (N_8942,N_7511,N_7570);
or U8943 (N_8943,N_7809,N_7527);
and U8944 (N_8944,N_8089,N_7940);
nor U8945 (N_8945,N_7919,N_7766);
or U8946 (N_8946,N_7985,N_7765);
or U8947 (N_8947,N_7874,N_7626);
and U8948 (N_8948,N_7954,N_7931);
or U8949 (N_8949,N_7851,N_7952);
and U8950 (N_8950,N_7983,N_7884);
nand U8951 (N_8951,N_7616,N_7602);
nor U8952 (N_8952,N_7719,N_8178);
nand U8953 (N_8953,N_7599,N_7934);
xnor U8954 (N_8954,N_8155,N_7817);
nor U8955 (N_8955,N_8197,N_7625);
and U8956 (N_8956,N_7673,N_7645);
nand U8957 (N_8957,N_7878,N_8193);
nor U8958 (N_8958,N_7958,N_7547);
nand U8959 (N_8959,N_7537,N_7913);
nand U8960 (N_8960,N_8236,N_8033);
or U8961 (N_8961,N_7748,N_8111);
nand U8962 (N_8962,N_8247,N_8169);
xor U8963 (N_8963,N_8131,N_8078);
nor U8964 (N_8964,N_8046,N_7536);
nand U8965 (N_8965,N_7979,N_8245);
nor U8966 (N_8966,N_7885,N_7589);
and U8967 (N_8967,N_8045,N_8153);
and U8968 (N_8968,N_7846,N_8197);
nor U8969 (N_8969,N_8040,N_8044);
and U8970 (N_8970,N_7928,N_8132);
and U8971 (N_8971,N_7981,N_7590);
and U8972 (N_8972,N_7655,N_8034);
xor U8973 (N_8973,N_8189,N_8184);
and U8974 (N_8974,N_7941,N_8198);
xor U8975 (N_8975,N_7673,N_7709);
and U8976 (N_8976,N_7809,N_8106);
or U8977 (N_8977,N_8172,N_7859);
nor U8978 (N_8978,N_8218,N_7976);
nand U8979 (N_8979,N_7856,N_8202);
or U8980 (N_8980,N_8132,N_7730);
and U8981 (N_8981,N_7643,N_7659);
and U8982 (N_8982,N_8242,N_7530);
nand U8983 (N_8983,N_8053,N_7720);
or U8984 (N_8984,N_8202,N_7779);
and U8985 (N_8985,N_8013,N_8086);
or U8986 (N_8986,N_8141,N_8129);
and U8987 (N_8987,N_7859,N_8235);
nor U8988 (N_8988,N_7679,N_7514);
nand U8989 (N_8989,N_7568,N_7840);
and U8990 (N_8990,N_7747,N_7559);
nand U8991 (N_8991,N_7991,N_8204);
nor U8992 (N_8992,N_8134,N_8241);
and U8993 (N_8993,N_7830,N_7538);
and U8994 (N_8994,N_8105,N_7570);
nor U8995 (N_8995,N_8110,N_7954);
nand U8996 (N_8996,N_8201,N_8188);
or U8997 (N_8997,N_7766,N_8218);
nor U8998 (N_8998,N_8051,N_8082);
and U8999 (N_8999,N_7962,N_7713);
nand U9000 (N_9000,N_8782,N_8351);
and U9001 (N_9001,N_8940,N_8493);
or U9002 (N_9002,N_8402,N_8676);
nor U9003 (N_9003,N_8689,N_8749);
or U9004 (N_9004,N_8721,N_8844);
nand U9005 (N_9005,N_8711,N_8411);
nor U9006 (N_9006,N_8769,N_8594);
nand U9007 (N_9007,N_8967,N_8706);
nand U9008 (N_9008,N_8751,N_8636);
nand U9009 (N_9009,N_8754,N_8976);
and U9010 (N_9010,N_8959,N_8894);
or U9011 (N_9011,N_8270,N_8687);
or U9012 (N_9012,N_8743,N_8739);
nor U9013 (N_9013,N_8622,N_8454);
xnor U9014 (N_9014,N_8436,N_8780);
nand U9015 (N_9015,N_8474,N_8898);
nor U9016 (N_9016,N_8364,N_8465);
and U9017 (N_9017,N_8934,N_8503);
and U9018 (N_9018,N_8539,N_8987);
nor U9019 (N_9019,N_8356,N_8334);
and U9020 (N_9020,N_8758,N_8651);
and U9021 (N_9021,N_8602,N_8981);
and U9022 (N_9022,N_8808,N_8870);
or U9023 (N_9023,N_8853,N_8256);
nor U9024 (N_9024,N_8813,N_8513);
and U9025 (N_9025,N_8328,N_8891);
xnor U9026 (N_9026,N_8648,N_8455);
and U9027 (N_9027,N_8771,N_8260);
xor U9028 (N_9028,N_8635,N_8292);
and U9029 (N_9029,N_8600,N_8606);
nor U9030 (N_9030,N_8816,N_8578);
nand U9031 (N_9031,N_8327,N_8984);
and U9032 (N_9032,N_8793,N_8779);
nor U9033 (N_9033,N_8387,N_8800);
and U9034 (N_9034,N_8755,N_8551);
nor U9035 (N_9035,N_8308,N_8753);
and U9036 (N_9036,N_8877,N_8737);
nor U9037 (N_9037,N_8952,N_8838);
and U9038 (N_9038,N_8437,N_8610);
or U9039 (N_9039,N_8840,N_8945);
and U9040 (N_9040,N_8629,N_8564);
and U9041 (N_9041,N_8814,N_8863);
and U9042 (N_9042,N_8943,N_8842);
or U9043 (N_9043,N_8765,N_8540);
nor U9044 (N_9044,N_8825,N_8896);
nand U9045 (N_9045,N_8382,N_8354);
or U9046 (N_9046,N_8748,N_8846);
nor U9047 (N_9047,N_8867,N_8901);
and U9048 (N_9048,N_8884,N_8484);
xnor U9049 (N_9049,N_8433,N_8831);
and U9050 (N_9050,N_8650,N_8533);
and U9051 (N_9051,N_8968,N_8611);
and U9052 (N_9052,N_8274,N_8306);
and U9053 (N_9053,N_8847,N_8851);
nand U9054 (N_9054,N_8605,N_8567);
nor U9055 (N_9055,N_8671,N_8326);
xnor U9056 (N_9056,N_8691,N_8582);
or U9057 (N_9057,N_8604,N_8584);
and U9058 (N_9058,N_8313,N_8427);
or U9059 (N_9059,N_8276,N_8441);
nand U9060 (N_9060,N_8845,N_8478);
nand U9061 (N_9061,N_8617,N_8544);
nor U9062 (N_9062,N_8268,N_8833);
and U9063 (N_9063,N_8592,N_8486);
nor U9064 (N_9064,N_8775,N_8294);
and U9065 (N_9065,N_8962,N_8649);
nor U9066 (N_9066,N_8405,N_8878);
xor U9067 (N_9067,N_8708,N_8498);
and U9068 (N_9068,N_8657,N_8798);
nor U9069 (N_9069,N_8668,N_8861);
and U9070 (N_9070,N_8709,N_8507);
and U9071 (N_9071,N_8438,N_8596);
nor U9072 (N_9072,N_8778,N_8640);
nor U9073 (N_9073,N_8581,N_8397);
xnor U9074 (N_9074,N_8911,N_8712);
nor U9075 (N_9075,N_8527,N_8757);
nor U9076 (N_9076,N_8324,N_8745);
or U9077 (N_9077,N_8783,N_8546);
nor U9078 (N_9078,N_8789,N_8407);
xor U9079 (N_9079,N_8693,N_8499);
and U9080 (N_9080,N_8419,N_8497);
nor U9081 (N_9081,N_8866,N_8740);
nor U9082 (N_9082,N_8995,N_8763);
xor U9083 (N_9083,N_8271,N_8876);
nor U9084 (N_9084,N_8543,N_8572);
xnor U9085 (N_9085,N_8509,N_8742);
and U9086 (N_9086,N_8930,N_8346);
and U9087 (N_9087,N_8929,N_8905);
nand U9088 (N_9088,N_8926,N_8342);
xnor U9089 (N_9089,N_8426,N_8983);
or U9090 (N_9090,N_8374,N_8283);
nand U9091 (N_9091,N_8439,N_8381);
and U9092 (N_9092,N_8373,N_8423);
xnor U9093 (N_9093,N_8852,N_8261);
and U9094 (N_9094,N_8817,N_8922);
nor U9095 (N_9095,N_8570,N_8915);
and U9096 (N_9096,N_8280,N_8655);
or U9097 (N_9097,N_8273,N_8704);
nand U9098 (N_9098,N_8781,N_8398);
nand U9099 (N_9099,N_8278,N_8453);
nor U9100 (N_9100,N_8723,N_8660);
and U9101 (N_9101,N_8580,N_8591);
nor U9102 (N_9102,N_8744,N_8514);
nand U9103 (N_9103,N_8836,N_8658);
nand U9104 (N_9104,N_8795,N_8377);
nand U9105 (N_9105,N_8431,N_8850);
and U9106 (N_9106,N_8625,N_8647);
nand U9107 (N_9107,N_8621,N_8803);
and U9108 (N_9108,N_8309,N_8534);
or U9109 (N_9109,N_8408,N_8291);
and U9110 (N_9110,N_8424,N_8715);
nand U9111 (N_9111,N_8978,N_8479);
xnor U9112 (N_9112,N_8832,N_8725);
nor U9113 (N_9113,N_8862,N_8906);
nor U9114 (N_9114,N_8951,N_8632);
and U9115 (N_9115,N_8400,N_8390);
and U9116 (N_9116,N_8488,N_8489);
nor U9117 (N_9117,N_8440,N_8536);
or U9118 (N_9118,N_8824,N_8675);
xnor U9119 (N_9119,N_8619,N_8756);
nor U9120 (N_9120,N_8826,N_8264);
xnor U9121 (N_9121,N_8928,N_8996);
nand U9122 (N_9122,N_8521,N_8639);
and U9123 (N_9123,N_8883,N_8975);
xnor U9124 (N_9124,N_8343,N_8993);
and U9125 (N_9125,N_8319,N_8552);
nor U9126 (N_9126,N_8760,N_8731);
nor U9127 (N_9127,N_8912,N_8307);
nor U9128 (N_9128,N_8537,N_8662);
and U9129 (N_9129,N_8827,N_8627);
and U9130 (N_9130,N_8614,N_8525);
nor U9131 (N_9131,N_8577,N_8332);
nand U9132 (N_9132,N_8900,N_8909);
and U9133 (N_9133,N_8750,N_8349);
or U9134 (N_9134,N_8821,N_8475);
nand U9135 (N_9135,N_8910,N_8561);
or U9136 (N_9136,N_8253,N_8504);
nand U9137 (N_9137,N_8683,N_8378);
and U9138 (N_9138,N_8340,N_8686);
or U9139 (N_9139,N_8776,N_8970);
nor U9140 (N_9140,N_8624,N_8696);
nor U9141 (N_9141,N_8937,N_8545);
and U9142 (N_9142,N_8288,N_8979);
or U9143 (N_9143,N_8277,N_8938);
nand U9144 (N_9144,N_8416,N_8616);
and U9145 (N_9145,N_8746,N_8576);
or U9146 (N_9146,N_8347,N_8442);
nand U9147 (N_9147,N_8257,N_8275);
nand U9148 (N_9148,N_8388,N_8366);
or U9149 (N_9149,N_8293,N_8550);
and U9150 (N_9150,N_8464,N_8738);
or U9151 (N_9151,N_8716,N_8941);
nand U9152 (N_9152,N_8532,N_8519);
nor U9153 (N_9153,N_8394,N_8384);
and U9154 (N_9154,N_8855,N_8574);
and U9155 (N_9155,N_8741,N_8659);
or U9156 (N_9156,N_8881,N_8892);
xnor U9157 (N_9157,N_8661,N_8508);
and U9158 (N_9158,N_8430,N_8589);
nand U9159 (N_9159,N_8897,N_8372);
nand U9160 (N_9160,N_8321,N_8797);
and U9161 (N_9161,N_8553,N_8457);
nor U9162 (N_9162,N_8396,N_8542);
and U9163 (N_9163,N_8429,N_8316);
nand U9164 (N_9164,N_8931,N_8980);
nand U9165 (N_9165,N_8714,N_8669);
or U9166 (N_9166,N_8871,N_8713);
nor U9167 (N_9167,N_8925,N_8972);
and U9168 (N_9168,N_8963,N_8365);
or U9169 (N_9169,N_8722,N_8494);
nor U9170 (N_9170,N_8330,N_8939);
nor U9171 (N_9171,N_8734,N_8391);
or U9172 (N_9172,N_8893,N_8302);
and U9173 (N_9173,N_8263,N_8692);
and U9174 (N_9174,N_8554,N_8946);
nor U9175 (N_9175,N_8667,N_8947);
nand U9176 (N_9176,N_8541,N_8727);
xnor U9177 (N_9177,N_8267,N_8523);
or U9178 (N_9178,N_8412,N_8485);
nor U9179 (N_9179,N_8918,N_8673);
or U9180 (N_9180,N_8456,N_8585);
and U9181 (N_9181,N_8392,N_8259);
nand U9182 (N_9182,N_8305,N_8468);
nand U9183 (N_9183,N_8341,N_8279);
xnor U9184 (N_9184,N_8875,N_8409);
or U9185 (N_9185,N_8774,N_8312);
and U9186 (N_9186,N_8435,N_8914);
nor U9187 (N_9187,N_8904,N_8467);
or U9188 (N_9188,N_8618,N_8815);
nor U9189 (N_9189,N_8530,N_8482);
or U9190 (N_9190,N_8960,N_8777);
or U9191 (N_9191,N_8566,N_8496);
nor U9192 (N_9192,N_8913,N_8811);
nand U9193 (N_9193,N_8401,N_8720);
and U9194 (N_9194,N_8282,N_8703);
and U9195 (N_9195,N_8702,N_8997);
nand U9196 (N_9196,N_8698,N_8770);
and U9197 (N_9197,N_8518,N_8690);
nor U9198 (N_9198,N_8994,N_8339);
nand U9199 (N_9199,N_8251,N_8303);
nor U9200 (N_9200,N_8590,N_8785);
and U9201 (N_9201,N_8699,N_8895);
nor U9202 (N_9202,N_8471,N_8790);
xor U9203 (N_9203,N_8563,N_8344);
nand U9204 (N_9204,N_8626,N_8950);
nor U9205 (N_9205,N_8425,N_8869);
nor U9206 (N_9206,N_8807,N_8924);
and U9207 (N_9207,N_8375,N_8656);
and U9208 (N_9208,N_8599,N_8961);
or U9209 (N_9209,N_8859,N_8643);
and U9210 (N_9210,N_8593,N_8359);
nand U9211 (N_9211,N_8501,N_8399);
nand U9212 (N_9212,N_8254,N_8357);
nand U9213 (N_9213,N_8290,N_8907);
nor U9214 (N_9214,N_8644,N_8747);
and U9215 (N_9215,N_8607,N_8973);
or U9216 (N_9216,N_8752,N_8443);
and U9217 (N_9217,N_8483,N_8571);
or U9218 (N_9218,N_8730,N_8452);
nand U9219 (N_9219,N_8965,N_8565);
or U9220 (N_9220,N_8728,N_8726);
or U9221 (N_9221,N_8410,N_8935);
or U9222 (N_9222,N_8573,N_8792);
nand U9223 (N_9223,N_8265,N_8286);
nor U9224 (N_9224,N_8879,N_8701);
nand U9225 (N_9225,N_8612,N_8255);
nor U9226 (N_9226,N_8472,N_8466);
or U9227 (N_9227,N_8562,N_8989);
and U9228 (N_9228,N_8856,N_8874);
nand U9229 (N_9229,N_8733,N_8415);
nand U9230 (N_9230,N_8393,N_8603);
and U9231 (N_9231,N_8369,N_8784);
nand U9232 (N_9232,N_8538,N_8395);
nand U9233 (N_9233,N_8956,N_8318);
and U9234 (N_9234,N_8890,N_8526);
nor U9235 (N_9235,N_8791,N_8977);
nor U9236 (N_9236,N_8331,N_8470);
and U9237 (N_9237,N_8707,N_8522);
nor U9238 (N_9238,N_8837,N_8272);
nor U9239 (N_9239,N_8487,N_8645);
or U9240 (N_9240,N_8336,N_8759);
and U9241 (N_9241,N_8587,N_8736);
nor U9242 (N_9242,N_8828,N_8506);
and U9243 (N_9243,N_8505,N_8250);
nor U9244 (N_9244,N_8413,N_8547);
nor U9245 (N_9245,N_8404,N_8732);
and U9246 (N_9246,N_8502,N_8700);
and U9247 (N_9247,N_8322,N_8964);
xnor U9248 (N_9248,N_8469,N_8969);
nor U9249 (N_9249,N_8841,N_8764);
and U9250 (N_9250,N_8462,N_8985);
and U9251 (N_9251,N_8490,N_8666);
nand U9252 (N_9252,N_8447,N_8609);
xor U9253 (N_9253,N_8857,N_8849);
nand U9254 (N_9254,N_8949,N_8588);
nor U9255 (N_9255,N_8459,N_8434);
nor U9256 (N_9256,N_8460,N_8865);
xnor U9257 (N_9257,N_8421,N_8284);
nor U9258 (N_9258,N_8524,N_8886);
nand U9259 (N_9259,N_8445,N_8310);
or U9260 (N_9260,N_8932,N_8766);
nand U9261 (N_9261,N_8717,N_8287);
nor U9262 (N_9262,N_8966,N_8812);
xor U9263 (N_9263,N_8835,N_8678);
nand U9264 (N_9264,N_8569,N_8406);
nand U9265 (N_9265,N_8642,N_8451);
or U9266 (N_9266,N_8559,N_8363);
nor U9267 (N_9267,N_8555,N_8848);
or U9268 (N_9268,N_8927,N_8768);
or U9269 (N_9269,N_8510,N_8535);
and U9270 (N_9270,N_8512,N_8586);
and U9271 (N_9271,N_8684,N_8608);
and U9272 (N_9272,N_8481,N_8988);
nor U9273 (N_9273,N_8954,N_8805);
or U9274 (N_9274,N_8549,N_8677);
and U9275 (N_9275,N_8615,N_8296);
and U9276 (N_9276,N_8773,N_8903);
and U9277 (N_9277,N_8633,N_8380);
xor U9278 (N_9278,N_8320,N_8990);
nor U9279 (N_9279,N_8473,N_8794);
or U9280 (N_9280,N_8575,N_8450);
nand U9281 (N_9281,N_8560,N_8806);
and U9282 (N_9282,N_8414,N_8799);
nand U9283 (N_9283,N_8338,N_8360);
xnor U9284 (N_9284,N_8697,N_8315);
nand U9285 (N_9285,N_8786,N_8665);
nand U9286 (N_9286,N_8323,N_8368);
or U9287 (N_9287,N_8477,N_8637);
nand U9288 (N_9288,N_8515,N_8705);
or U9289 (N_9289,N_8718,N_8352);
nand U9290 (N_9290,N_8682,N_8528);
xor U9291 (N_9291,N_8860,N_8556);
nor U9292 (N_9292,N_8834,N_8295);
nor U9293 (N_9293,N_8646,N_8719);
nand U9294 (N_9294,N_8289,N_8371);
and U9295 (N_9295,N_8921,N_8449);
nor U9296 (N_9296,N_8558,N_8819);
xor U9297 (N_9297,N_8767,N_8333);
xor U9298 (N_9298,N_8376,N_8641);
nor U9299 (N_9299,N_8818,N_8936);
nor U9300 (N_9300,N_8694,N_8325);
or U9301 (N_9301,N_8735,N_8262);
nor U9302 (N_9302,N_8680,N_8971);
and U9303 (N_9303,N_8948,N_8461);
or U9304 (N_9304,N_8919,N_8362);
nor U9305 (N_9305,N_8724,N_8269);
nor U9306 (N_9306,N_8298,N_8796);
and U9307 (N_9307,N_8548,N_8579);
nand U9308 (N_9308,N_8500,N_8998);
or U9309 (N_9309,N_8953,N_8864);
nand U9310 (N_9310,N_8557,N_8598);
nand U9311 (N_9311,N_8568,N_8999);
or U9312 (N_9312,N_8920,N_8628);
nor U9313 (N_9313,N_8710,N_8670);
nor U9314 (N_9314,N_8385,N_8531);
and U9315 (N_9315,N_8986,N_8882);
nand U9316 (N_9316,N_8788,N_8417);
nor U9317 (N_9317,N_8944,N_8448);
nand U9318 (N_9318,N_8982,N_8285);
and U9319 (N_9319,N_8762,N_8992);
nor U9320 (N_9320,N_8353,N_8420);
and U9321 (N_9321,N_8252,N_8418);
or U9322 (N_9322,N_8370,N_8383);
nor U9323 (N_9323,N_8444,N_8311);
nand U9324 (N_9324,N_8335,N_8428);
nand U9325 (N_9325,N_8787,N_8258);
nand U9326 (N_9326,N_8367,N_8495);
nand U9327 (N_9327,N_8634,N_8804);
and U9328 (N_9328,N_8653,N_8809);
and U9329 (N_9329,N_8991,N_8888);
and U9330 (N_9330,N_8297,N_8957);
xnor U9331 (N_9331,N_8317,N_8638);
and U9332 (N_9332,N_8491,N_8299);
and U9333 (N_9333,N_8595,N_8301);
xor U9334 (N_9334,N_8917,N_8652);
nand U9335 (N_9335,N_8663,N_8955);
and U9336 (N_9336,N_8422,N_8511);
xor U9337 (N_9337,N_8823,N_8873);
and U9338 (N_9338,N_8654,N_8885);
nor U9339 (N_9339,N_8872,N_8345);
or U9340 (N_9340,N_8772,N_8386);
xnor U9341 (N_9341,N_8446,N_8516);
nand U9342 (N_9342,N_8902,N_8379);
nand U9343 (N_9343,N_8520,N_8761);
nor U9344 (N_9344,N_8672,N_8880);
or U9345 (N_9345,N_8529,N_8432);
nand U9346 (N_9346,N_8300,N_8942);
nand U9347 (N_9347,N_8729,N_8854);
nand U9348 (N_9348,N_8908,N_8304);
nor U9349 (N_9349,N_8403,N_8355);
xnor U9350 (N_9350,N_8517,N_8348);
and U9351 (N_9351,N_8887,N_8281);
nor U9352 (N_9352,N_8933,N_8458);
nor U9353 (N_9353,N_8889,N_8923);
and U9354 (N_9354,N_8916,N_8695);
xor U9355 (N_9355,N_8358,N_8480);
xnor U9356 (N_9356,N_8389,N_8613);
nor U9357 (N_9357,N_8820,N_8664);
nand U9358 (N_9358,N_8858,N_8463);
nand U9359 (N_9359,N_8839,N_8958);
nor U9360 (N_9360,N_8829,N_8583);
nand U9361 (N_9361,N_8620,N_8685);
nand U9362 (N_9362,N_8899,N_8688);
nand U9363 (N_9363,N_8601,N_8597);
nor U9364 (N_9364,N_8314,N_8679);
nand U9365 (N_9365,N_8476,N_8802);
and U9366 (N_9366,N_8266,N_8623);
nor U9367 (N_9367,N_8350,N_8674);
nand U9368 (N_9368,N_8843,N_8974);
and U9369 (N_9369,N_8681,N_8810);
nand U9370 (N_9370,N_8492,N_8630);
or U9371 (N_9371,N_8361,N_8631);
or U9372 (N_9372,N_8868,N_8830);
and U9373 (N_9373,N_8329,N_8822);
nand U9374 (N_9374,N_8801,N_8337);
nand U9375 (N_9375,N_8279,N_8934);
and U9376 (N_9376,N_8699,N_8506);
or U9377 (N_9377,N_8510,N_8873);
nor U9378 (N_9378,N_8649,N_8558);
and U9379 (N_9379,N_8366,N_8988);
nand U9380 (N_9380,N_8701,N_8784);
xor U9381 (N_9381,N_8680,N_8935);
and U9382 (N_9382,N_8634,N_8950);
or U9383 (N_9383,N_8578,N_8566);
or U9384 (N_9384,N_8591,N_8946);
nand U9385 (N_9385,N_8739,N_8560);
and U9386 (N_9386,N_8460,N_8805);
and U9387 (N_9387,N_8552,N_8672);
or U9388 (N_9388,N_8441,N_8609);
and U9389 (N_9389,N_8590,N_8669);
or U9390 (N_9390,N_8268,N_8364);
and U9391 (N_9391,N_8683,N_8595);
and U9392 (N_9392,N_8423,N_8651);
nor U9393 (N_9393,N_8937,N_8958);
and U9394 (N_9394,N_8669,N_8336);
nand U9395 (N_9395,N_8574,N_8743);
nor U9396 (N_9396,N_8283,N_8901);
nand U9397 (N_9397,N_8731,N_8435);
or U9398 (N_9398,N_8821,N_8610);
and U9399 (N_9399,N_8807,N_8949);
nand U9400 (N_9400,N_8517,N_8653);
nor U9401 (N_9401,N_8616,N_8251);
and U9402 (N_9402,N_8304,N_8254);
nand U9403 (N_9403,N_8650,N_8497);
or U9404 (N_9404,N_8746,N_8420);
nand U9405 (N_9405,N_8336,N_8765);
xnor U9406 (N_9406,N_8735,N_8362);
nand U9407 (N_9407,N_8747,N_8552);
and U9408 (N_9408,N_8393,N_8327);
nor U9409 (N_9409,N_8634,N_8372);
xnor U9410 (N_9410,N_8692,N_8261);
or U9411 (N_9411,N_8526,N_8853);
nand U9412 (N_9412,N_8971,N_8779);
and U9413 (N_9413,N_8544,N_8951);
and U9414 (N_9414,N_8456,N_8251);
and U9415 (N_9415,N_8303,N_8984);
or U9416 (N_9416,N_8446,N_8513);
xor U9417 (N_9417,N_8500,N_8598);
and U9418 (N_9418,N_8768,N_8841);
nor U9419 (N_9419,N_8452,N_8692);
or U9420 (N_9420,N_8815,N_8692);
nand U9421 (N_9421,N_8455,N_8596);
nand U9422 (N_9422,N_8525,N_8658);
or U9423 (N_9423,N_8515,N_8842);
nand U9424 (N_9424,N_8616,N_8431);
nand U9425 (N_9425,N_8883,N_8800);
nor U9426 (N_9426,N_8779,N_8309);
or U9427 (N_9427,N_8686,N_8758);
and U9428 (N_9428,N_8487,N_8885);
or U9429 (N_9429,N_8729,N_8939);
or U9430 (N_9430,N_8444,N_8877);
or U9431 (N_9431,N_8925,N_8611);
nand U9432 (N_9432,N_8333,N_8906);
nor U9433 (N_9433,N_8927,N_8803);
and U9434 (N_9434,N_8335,N_8880);
nor U9435 (N_9435,N_8819,N_8697);
and U9436 (N_9436,N_8901,N_8784);
xnor U9437 (N_9437,N_8408,N_8791);
nand U9438 (N_9438,N_8865,N_8426);
and U9439 (N_9439,N_8686,N_8850);
and U9440 (N_9440,N_8689,N_8918);
and U9441 (N_9441,N_8702,N_8671);
and U9442 (N_9442,N_8444,N_8734);
or U9443 (N_9443,N_8549,N_8517);
xnor U9444 (N_9444,N_8804,N_8640);
and U9445 (N_9445,N_8785,N_8984);
nand U9446 (N_9446,N_8793,N_8297);
nand U9447 (N_9447,N_8631,N_8683);
nor U9448 (N_9448,N_8982,N_8428);
and U9449 (N_9449,N_8408,N_8565);
nor U9450 (N_9450,N_8364,N_8631);
and U9451 (N_9451,N_8474,N_8514);
nand U9452 (N_9452,N_8642,N_8424);
xor U9453 (N_9453,N_8423,N_8571);
nor U9454 (N_9454,N_8680,N_8706);
nand U9455 (N_9455,N_8884,N_8916);
nand U9456 (N_9456,N_8491,N_8979);
xnor U9457 (N_9457,N_8976,N_8693);
nand U9458 (N_9458,N_8945,N_8567);
or U9459 (N_9459,N_8951,N_8834);
nand U9460 (N_9460,N_8475,N_8836);
or U9461 (N_9461,N_8906,N_8934);
and U9462 (N_9462,N_8507,N_8508);
nand U9463 (N_9463,N_8561,N_8266);
or U9464 (N_9464,N_8867,N_8559);
nor U9465 (N_9465,N_8931,N_8383);
xnor U9466 (N_9466,N_8492,N_8607);
xnor U9467 (N_9467,N_8376,N_8595);
or U9468 (N_9468,N_8654,N_8746);
nor U9469 (N_9469,N_8686,N_8740);
and U9470 (N_9470,N_8969,N_8745);
xor U9471 (N_9471,N_8598,N_8963);
or U9472 (N_9472,N_8937,N_8872);
and U9473 (N_9473,N_8916,N_8345);
nand U9474 (N_9474,N_8513,N_8475);
or U9475 (N_9475,N_8336,N_8893);
or U9476 (N_9476,N_8833,N_8261);
nand U9477 (N_9477,N_8348,N_8793);
nand U9478 (N_9478,N_8592,N_8417);
nor U9479 (N_9479,N_8590,N_8543);
nand U9480 (N_9480,N_8301,N_8674);
or U9481 (N_9481,N_8483,N_8926);
nor U9482 (N_9482,N_8893,N_8921);
nand U9483 (N_9483,N_8418,N_8267);
or U9484 (N_9484,N_8670,N_8426);
nor U9485 (N_9485,N_8620,N_8323);
nand U9486 (N_9486,N_8397,N_8452);
and U9487 (N_9487,N_8993,N_8716);
nand U9488 (N_9488,N_8870,N_8995);
or U9489 (N_9489,N_8924,N_8856);
nor U9490 (N_9490,N_8339,N_8420);
nand U9491 (N_9491,N_8597,N_8675);
nand U9492 (N_9492,N_8942,N_8870);
xor U9493 (N_9493,N_8601,N_8556);
or U9494 (N_9494,N_8880,N_8478);
nand U9495 (N_9495,N_8939,N_8302);
or U9496 (N_9496,N_8490,N_8618);
nor U9497 (N_9497,N_8278,N_8767);
nand U9498 (N_9498,N_8921,N_8382);
nand U9499 (N_9499,N_8805,N_8337);
xor U9500 (N_9500,N_8895,N_8689);
nor U9501 (N_9501,N_8409,N_8571);
nand U9502 (N_9502,N_8801,N_8485);
nor U9503 (N_9503,N_8711,N_8581);
xor U9504 (N_9504,N_8976,N_8950);
or U9505 (N_9505,N_8726,N_8483);
or U9506 (N_9506,N_8908,N_8421);
and U9507 (N_9507,N_8277,N_8478);
or U9508 (N_9508,N_8723,N_8619);
nand U9509 (N_9509,N_8755,N_8690);
xor U9510 (N_9510,N_8842,N_8273);
nand U9511 (N_9511,N_8546,N_8667);
xnor U9512 (N_9512,N_8827,N_8749);
and U9513 (N_9513,N_8849,N_8765);
nand U9514 (N_9514,N_8941,N_8335);
and U9515 (N_9515,N_8739,N_8303);
or U9516 (N_9516,N_8564,N_8940);
and U9517 (N_9517,N_8299,N_8762);
nand U9518 (N_9518,N_8588,N_8334);
xor U9519 (N_9519,N_8660,N_8919);
nand U9520 (N_9520,N_8325,N_8278);
or U9521 (N_9521,N_8777,N_8751);
nand U9522 (N_9522,N_8444,N_8912);
xor U9523 (N_9523,N_8998,N_8580);
nand U9524 (N_9524,N_8991,N_8868);
or U9525 (N_9525,N_8709,N_8436);
and U9526 (N_9526,N_8929,N_8797);
or U9527 (N_9527,N_8866,N_8503);
and U9528 (N_9528,N_8352,N_8856);
nor U9529 (N_9529,N_8832,N_8653);
or U9530 (N_9530,N_8686,N_8370);
xnor U9531 (N_9531,N_8423,N_8548);
nor U9532 (N_9532,N_8800,N_8429);
and U9533 (N_9533,N_8338,N_8742);
nand U9534 (N_9534,N_8463,N_8326);
nand U9535 (N_9535,N_8726,N_8659);
nor U9536 (N_9536,N_8612,N_8974);
nand U9537 (N_9537,N_8912,N_8520);
and U9538 (N_9538,N_8996,N_8406);
or U9539 (N_9539,N_8754,N_8722);
or U9540 (N_9540,N_8543,N_8518);
and U9541 (N_9541,N_8736,N_8904);
nand U9542 (N_9542,N_8580,N_8701);
nor U9543 (N_9543,N_8410,N_8483);
and U9544 (N_9544,N_8396,N_8867);
xnor U9545 (N_9545,N_8340,N_8917);
or U9546 (N_9546,N_8365,N_8466);
nor U9547 (N_9547,N_8438,N_8675);
or U9548 (N_9548,N_8346,N_8372);
or U9549 (N_9549,N_8502,N_8777);
or U9550 (N_9550,N_8952,N_8358);
nor U9551 (N_9551,N_8823,N_8964);
nand U9552 (N_9552,N_8890,N_8651);
or U9553 (N_9553,N_8771,N_8504);
and U9554 (N_9554,N_8509,N_8368);
nor U9555 (N_9555,N_8367,N_8604);
or U9556 (N_9556,N_8621,N_8332);
xor U9557 (N_9557,N_8582,N_8363);
and U9558 (N_9558,N_8716,N_8718);
or U9559 (N_9559,N_8914,N_8556);
xor U9560 (N_9560,N_8587,N_8975);
or U9561 (N_9561,N_8292,N_8579);
and U9562 (N_9562,N_8813,N_8797);
nand U9563 (N_9563,N_8574,N_8792);
or U9564 (N_9564,N_8704,N_8442);
and U9565 (N_9565,N_8987,N_8293);
and U9566 (N_9566,N_8758,N_8539);
nor U9567 (N_9567,N_8505,N_8592);
nand U9568 (N_9568,N_8995,N_8472);
or U9569 (N_9569,N_8472,N_8963);
and U9570 (N_9570,N_8581,N_8843);
or U9571 (N_9571,N_8716,N_8487);
nor U9572 (N_9572,N_8550,N_8351);
nand U9573 (N_9573,N_8474,N_8972);
or U9574 (N_9574,N_8821,N_8918);
and U9575 (N_9575,N_8888,N_8526);
or U9576 (N_9576,N_8397,N_8710);
and U9577 (N_9577,N_8264,N_8904);
nor U9578 (N_9578,N_8880,N_8596);
nand U9579 (N_9579,N_8664,N_8434);
nand U9580 (N_9580,N_8694,N_8479);
or U9581 (N_9581,N_8952,N_8382);
nor U9582 (N_9582,N_8774,N_8958);
nand U9583 (N_9583,N_8592,N_8922);
or U9584 (N_9584,N_8678,N_8749);
or U9585 (N_9585,N_8387,N_8595);
nor U9586 (N_9586,N_8908,N_8856);
nor U9587 (N_9587,N_8411,N_8628);
nor U9588 (N_9588,N_8294,N_8425);
xor U9589 (N_9589,N_8399,N_8645);
and U9590 (N_9590,N_8718,N_8415);
nor U9591 (N_9591,N_8631,N_8443);
or U9592 (N_9592,N_8934,N_8667);
or U9593 (N_9593,N_8999,N_8269);
nor U9594 (N_9594,N_8290,N_8865);
nand U9595 (N_9595,N_8896,N_8680);
nor U9596 (N_9596,N_8346,N_8545);
xor U9597 (N_9597,N_8577,N_8423);
and U9598 (N_9598,N_8367,N_8369);
and U9599 (N_9599,N_8388,N_8368);
nor U9600 (N_9600,N_8617,N_8718);
or U9601 (N_9601,N_8396,N_8988);
or U9602 (N_9602,N_8822,N_8654);
nand U9603 (N_9603,N_8919,N_8987);
nor U9604 (N_9604,N_8571,N_8912);
nor U9605 (N_9605,N_8396,N_8842);
or U9606 (N_9606,N_8505,N_8282);
nor U9607 (N_9607,N_8339,N_8851);
and U9608 (N_9608,N_8839,N_8386);
or U9609 (N_9609,N_8748,N_8834);
and U9610 (N_9610,N_8696,N_8289);
and U9611 (N_9611,N_8754,N_8844);
and U9612 (N_9612,N_8529,N_8871);
nand U9613 (N_9613,N_8379,N_8787);
nand U9614 (N_9614,N_8863,N_8682);
or U9615 (N_9615,N_8756,N_8918);
and U9616 (N_9616,N_8770,N_8942);
and U9617 (N_9617,N_8859,N_8377);
nand U9618 (N_9618,N_8708,N_8286);
and U9619 (N_9619,N_8426,N_8449);
nor U9620 (N_9620,N_8937,N_8564);
or U9621 (N_9621,N_8665,N_8742);
and U9622 (N_9622,N_8740,N_8415);
nand U9623 (N_9623,N_8906,N_8978);
xor U9624 (N_9624,N_8948,N_8985);
xnor U9625 (N_9625,N_8496,N_8930);
nor U9626 (N_9626,N_8712,N_8352);
nand U9627 (N_9627,N_8578,N_8398);
or U9628 (N_9628,N_8934,N_8941);
or U9629 (N_9629,N_8560,N_8938);
nor U9630 (N_9630,N_8380,N_8928);
xor U9631 (N_9631,N_8723,N_8278);
xnor U9632 (N_9632,N_8748,N_8753);
or U9633 (N_9633,N_8552,N_8886);
nor U9634 (N_9634,N_8675,N_8761);
nor U9635 (N_9635,N_8559,N_8378);
nand U9636 (N_9636,N_8662,N_8453);
or U9637 (N_9637,N_8771,N_8798);
xnor U9638 (N_9638,N_8890,N_8250);
or U9639 (N_9639,N_8600,N_8914);
or U9640 (N_9640,N_8646,N_8419);
nand U9641 (N_9641,N_8609,N_8847);
and U9642 (N_9642,N_8988,N_8672);
or U9643 (N_9643,N_8889,N_8474);
xor U9644 (N_9644,N_8642,N_8341);
xnor U9645 (N_9645,N_8748,N_8371);
nor U9646 (N_9646,N_8992,N_8543);
nand U9647 (N_9647,N_8779,N_8949);
nand U9648 (N_9648,N_8631,N_8626);
nor U9649 (N_9649,N_8977,N_8510);
or U9650 (N_9650,N_8711,N_8871);
nand U9651 (N_9651,N_8971,N_8305);
nand U9652 (N_9652,N_8304,N_8904);
nand U9653 (N_9653,N_8428,N_8802);
nor U9654 (N_9654,N_8670,N_8564);
and U9655 (N_9655,N_8410,N_8638);
or U9656 (N_9656,N_8904,N_8657);
and U9657 (N_9657,N_8423,N_8803);
and U9658 (N_9658,N_8528,N_8718);
or U9659 (N_9659,N_8756,N_8350);
nor U9660 (N_9660,N_8368,N_8691);
nor U9661 (N_9661,N_8676,N_8489);
nor U9662 (N_9662,N_8988,N_8817);
nand U9663 (N_9663,N_8527,N_8471);
and U9664 (N_9664,N_8953,N_8603);
and U9665 (N_9665,N_8781,N_8901);
nor U9666 (N_9666,N_8811,N_8898);
nor U9667 (N_9667,N_8959,N_8895);
or U9668 (N_9668,N_8899,N_8548);
or U9669 (N_9669,N_8532,N_8418);
nand U9670 (N_9670,N_8470,N_8766);
or U9671 (N_9671,N_8870,N_8810);
nand U9672 (N_9672,N_8882,N_8983);
nand U9673 (N_9673,N_8516,N_8594);
nor U9674 (N_9674,N_8875,N_8444);
nand U9675 (N_9675,N_8573,N_8298);
nand U9676 (N_9676,N_8666,N_8255);
nor U9677 (N_9677,N_8582,N_8355);
or U9678 (N_9678,N_8511,N_8770);
nand U9679 (N_9679,N_8648,N_8906);
nor U9680 (N_9680,N_8418,N_8997);
and U9681 (N_9681,N_8278,N_8609);
and U9682 (N_9682,N_8854,N_8505);
nand U9683 (N_9683,N_8667,N_8536);
nor U9684 (N_9684,N_8678,N_8422);
or U9685 (N_9685,N_8731,N_8696);
or U9686 (N_9686,N_8812,N_8361);
and U9687 (N_9687,N_8390,N_8396);
nor U9688 (N_9688,N_8491,N_8451);
nor U9689 (N_9689,N_8473,N_8495);
and U9690 (N_9690,N_8489,N_8576);
and U9691 (N_9691,N_8387,N_8593);
nor U9692 (N_9692,N_8399,N_8744);
or U9693 (N_9693,N_8257,N_8580);
nor U9694 (N_9694,N_8251,N_8629);
nand U9695 (N_9695,N_8379,N_8933);
nand U9696 (N_9696,N_8960,N_8512);
and U9697 (N_9697,N_8703,N_8329);
nor U9698 (N_9698,N_8488,N_8594);
nand U9699 (N_9699,N_8998,N_8560);
nor U9700 (N_9700,N_8344,N_8601);
xnor U9701 (N_9701,N_8277,N_8879);
and U9702 (N_9702,N_8478,N_8488);
and U9703 (N_9703,N_8928,N_8269);
nand U9704 (N_9704,N_8980,N_8889);
xnor U9705 (N_9705,N_8453,N_8594);
or U9706 (N_9706,N_8636,N_8353);
nor U9707 (N_9707,N_8411,N_8861);
nand U9708 (N_9708,N_8922,N_8981);
xor U9709 (N_9709,N_8643,N_8825);
xnor U9710 (N_9710,N_8471,N_8273);
or U9711 (N_9711,N_8358,N_8832);
nand U9712 (N_9712,N_8431,N_8283);
or U9713 (N_9713,N_8497,N_8924);
or U9714 (N_9714,N_8472,N_8921);
nand U9715 (N_9715,N_8838,N_8805);
and U9716 (N_9716,N_8649,N_8542);
nor U9717 (N_9717,N_8273,N_8406);
xor U9718 (N_9718,N_8520,N_8906);
or U9719 (N_9719,N_8582,N_8464);
and U9720 (N_9720,N_8435,N_8382);
and U9721 (N_9721,N_8399,N_8648);
xor U9722 (N_9722,N_8911,N_8290);
nor U9723 (N_9723,N_8927,N_8287);
nand U9724 (N_9724,N_8344,N_8702);
nor U9725 (N_9725,N_8655,N_8383);
nor U9726 (N_9726,N_8995,N_8263);
and U9727 (N_9727,N_8924,N_8554);
xnor U9728 (N_9728,N_8405,N_8366);
nor U9729 (N_9729,N_8549,N_8841);
and U9730 (N_9730,N_8764,N_8292);
or U9731 (N_9731,N_8368,N_8893);
xor U9732 (N_9732,N_8756,N_8261);
nand U9733 (N_9733,N_8875,N_8348);
or U9734 (N_9734,N_8572,N_8337);
nor U9735 (N_9735,N_8824,N_8271);
nor U9736 (N_9736,N_8320,N_8817);
nand U9737 (N_9737,N_8796,N_8424);
xnor U9738 (N_9738,N_8478,N_8983);
and U9739 (N_9739,N_8999,N_8887);
nand U9740 (N_9740,N_8919,N_8720);
and U9741 (N_9741,N_8410,N_8685);
or U9742 (N_9742,N_8722,N_8624);
and U9743 (N_9743,N_8826,N_8367);
nand U9744 (N_9744,N_8967,N_8977);
nor U9745 (N_9745,N_8695,N_8452);
nand U9746 (N_9746,N_8686,N_8322);
nor U9747 (N_9747,N_8401,N_8830);
nor U9748 (N_9748,N_8403,N_8624);
nor U9749 (N_9749,N_8288,N_8738);
nor U9750 (N_9750,N_9627,N_9578);
xor U9751 (N_9751,N_9381,N_9096);
and U9752 (N_9752,N_9666,N_9515);
or U9753 (N_9753,N_9300,N_9063);
nor U9754 (N_9754,N_9620,N_9140);
nor U9755 (N_9755,N_9661,N_9614);
nand U9756 (N_9756,N_9498,N_9223);
and U9757 (N_9757,N_9095,N_9424);
or U9758 (N_9758,N_9748,N_9071);
nor U9759 (N_9759,N_9342,N_9746);
and U9760 (N_9760,N_9189,N_9728);
or U9761 (N_9761,N_9016,N_9123);
and U9762 (N_9762,N_9397,N_9744);
nor U9763 (N_9763,N_9443,N_9311);
nand U9764 (N_9764,N_9507,N_9710);
nand U9765 (N_9765,N_9359,N_9470);
nor U9766 (N_9766,N_9029,N_9668);
nand U9767 (N_9767,N_9177,N_9567);
and U9768 (N_9768,N_9678,N_9256);
nor U9769 (N_9769,N_9524,N_9345);
nor U9770 (N_9770,N_9012,N_9416);
or U9771 (N_9771,N_9482,N_9546);
nor U9772 (N_9772,N_9210,N_9303);
and U9773 (N_9773,N_9525,N_9636);
or U9774 (N_9774,N_9611,N_9164);
nand U9775 (N_9775,N_9370,N_9708);
nor U9776 (N_9776,N_9101,N_9421);
or U9777 (N_9777,N_9079,N_9669);
or U9778 (N_9778,N_9100,N_9230);
xnor U9779 (N_9779,N_9175,N_9267);
or U9780 (N_9780,N_9486,N_9640);
or U9781 (N_9781,N_9149,N_9255);
or U9782 (N_9782,N_9201,N_9682);
nor U9783 (N_9783,N_9539,N_9146);
xnor U9784 (N_9784,N_9185,N_9444);
nor U9785 (N_9785,N_9225,N_9472);
and U9786 (N_9786,N_9504,N_9377);
and U9787 (N_9787,N_9566,N_9325);
and U9788 (N_9788,N_9235,N_9160);
or U9789 (N_9789,N_9371,N_9511);
or U9790 (N_9790,N_9464,N_9270);
nand U9791 (N_9791,N_9142,N_9642);
or U9792 (N_9792,N_9112,N_9493);
nor U9793 (N_9793,N_9109,N_9473);
nand U9794 (N_9794,N_9242,N_9222);
nand U9795 (N_9795,N_9147,N_9042);
nor U9796 (N_9796,N_9332,N_9205);
or U9797 (N_9797,N_9038,N_9172);
nand U9798 (N_9798,N_9502,N_9400);
and U9799 (N_9799,N_9088,N_9239);
and U9800 (N_9800,N_9035,N_9451);
and U9801 (N_9801,N_9186,N_9036);
nand U9802 (N_9802,N_9570,N_9388);
or U9803 (N_9803,N_9415,N_9393);
or U9804 (N_9804,N_9612,N_9729);
nor U9805 (N_9805,N_9544,N_9138);
xor U9806 (N_9806,N_9010,N_9173);
xor U9807 (N_9807,N_9425,N_9298);
or U9808 (N_9808,N_9619,N_9509);
or U9809 (N_9809,N_9686,N_9580);
or U9810 (N_9810,N_9534,N_9553);
and U9811 (N_9811,N_9248,N_9412);
or U9812 (N_9812,N_9284,N_9521);
nor U9813 (N_9813,N_9059,N_9306);
and U9814 (N_9814,N_9536,N_9015);
and U9815 (N_9815,N_9389,N_9658);
and U9816 (N_9816,N_9090,N_9179);
nand U9817 (N_9817,N_9049,N_9593);
and U9818 (N_9818,N_9354,N_9572);
nor U9819 (N_9819,N_9152,N_9241);
and U9820 (N_9820,N_9556,N_9322);
xor U9821 (N_9821,N_9745,N_9081);
nand U9822 (N_9822,N_9585,N_9635);
and U9823 (N_9823,N_9691,N_9655);
nand U9824 (N_9824,N_9277,N_9613);
or U9825 (N_9825,N_9219,N_9232);
or U9826 (N_9826,N_9467,N_9356);
nor U9827 (N_9827,N_9517,N_9254);
nand U9828 (N_9828,N_9542,N_9537);
or U9829 (N_9829,N_9383,N_9192);
nor U9830 (N_9830,N_9286,N_9700);
or U9831 (N_9831,N_9725,N_9721);
or U9832 (N_9832,N_9519,N_9245);
or U9833 (N_9833,N_9044,N_9500);
nand U9834 (N_9834,N_9604,N_9183);
or U9835 (N_9835,N_9422,N_9603);
or U9836 (N_9836,N_9363,N_9233);
or U9837 (N_9837,N_9153,N_9382);
nand U9838 (N_9838,N_9471,N_9034);
xor U9839 (N_9839,N_9115,N_9633);
or U9840 (N_9840,N_9740,N_9558);
nor U9841 (N_9841,N_9538,N_9430);
nand U9842 (N_9842,N_9310,N_9176);
or U9843 (N_9843,N_9628,N_9344);
nor U9844 (N_9844,N_9391,N_9738);
and U9845 (N_9845,N_9560,N_9196);
and U9846 (N_9846,N_9261,N_9439);
or U9847 (N_9847,N_9132,N_9257);
xnor U9848 (N_9848,N_9328,N_9301);
nor U9849 (N_9849,N_9271,N_9625);
nor U9850 (N_9850,N_9663,N_9720);
or U9851 (N_9851,N_9126,N_9372);
nand U9852 (N_9852,N_9013,N_9074);
xor U9853 (N_9853,N_9073,N_9208);
and U9854 (N_9854,N_9413,N_9699);
and U9855 (N_9855,N_9212,N_9707);
nand U9856 (N_9856,N_9170,N_9343);
and U9857 (N_9857,N_9541,N_9549);
xnor U9858 (N_9858,N_9703,N_9463);
or U9859 (N_9859,N_9449,N_9357);
and U9860 (N_9860,N_9169,N_9351);
and U9861 (N_9861,N_9369,N_9436);
nand U9862 (N_9862,N_9395,N_9253);
and U9863 (N_9863,N_9227,N_9615);
or U9864 (N_9864,N_9695,N_9045);
or U9865 (N_9865,N_9522,N_9597);
xor U9866 (N_9866,N_9462,N_9319);
or U9867 (N_9867,N_9005,N_9487);
xor U9868 (N_9868,N_9419,N_9739);
nor U9869 (N_9869,N_9075,N_9122);
nor U9870 (N_9870,N_9320,N_9608);
nor U9871 (N_9871,N_9237,N_9398);
nor U9872 (N_9872,N_9428,N_9280);
nand U9873 (N_9873,N_9569,N_9204);
or U9874 (N_9874,N_9143,N_9066);
nor U9875 (N_9875,N_9070,N_9749);
nand U9876 (N_9876,N_9503,N_9292);
or U9877 (N_9877,N_9526,N_9694);
nand U9878 (N_9878,N_9052,N_9673);
and U9879 (N_9879,N_9350,N_9531);
or U9880 (N_9880,N_9043,N_9165);
and U9881 (N_9881,N_9574,N_9547);
or U9882 (N_9882,N_9730,N_9330);
and U9883 (N_9883,N_9656,N_9665);
or U9884 (N_9884,N_9732,N_9590);
nand U9885 (N_9885,N_9247,N_9483);
and U9886 (N_9886,N_9137,N_9119);
nor U9887 (N_9887,N_9394,N_9209);
and U9888 (N_9888,N_9705,N_9014);
nor U9889 (N_9889,N_9039,N_9638);
and U9890 (N_9890,N_9453,N_9402);
nor U9891 (N_9891,N_9206,N_9654);
nor U9892 (N_9892,N_9262,N_9194);
or U9893 (N_9893,N_9027,N_9226);
nor U9894 (N_9894,N_9168,N_9392);
nand U9895 (N_9895,N_9671,N_9246);
xor U9896 (N_9896,N_9452,N_9494);
nor U9897 (N_9897,N_9200,N_9698);
nor U9898 (N_9898,N_9490,N_9631);
nor U9899 (N_9899,N_9712,N_9315);
or U9900 (N_9900,N_9557,N_9065);
and U9901 (N_9901,N_9496,N_9723);
xor U9902 (N_9902,N_9459,N_9437);
nand U9903 (N_9903,N_9530,N_9337);
xor U9904 (N_9904,N_9622,N_9743);
nand U9905 (N_9905,N_9684,N_9180);
nand U9906 (N_9906,N_9327,N_9644);
nor U9907 (N_9907,N_9385,N_9680);
nor U9908 (N_9908,N_9404,N_9440);
xor U9909 (N_9909,N_9528,N_9195);
xor U9910 (N_9910,N_9064,N_9019);
nand U9911 (N_9911,N_9202,N_9069);
and U9912 (N_9912,N_9163,N_9505);
or U9913 (N_9913,N_9040,N_9150);
xnor U9914 (N_9914,N_9353,N_9349);
xor U9915 (N_9915,N_9610,N_9555);
and U9916 (N_9916,N_9217,N_9406);
or U9917 (N_9917,N_9662,N_9191);
or U9918 (N_9918,N_9594,N_9649);
nand U9919 (N_9919,N_9252,N_9347);
or U9920 (N_9920,N_9076,N_9031);
xor U9921 (N_9921,N_9719,N_9333);
nand U9922 (N_9922,N_9450,N_9057);
or U9923 (N_9923,N_9024,N_9427);
or U9924 (N_9924,N_9514,N_9533);
or U9925 (N_9925,N_9687,N_9285);
xnor U9926 (N_9926,N_9484,N_9139);
xor U9927 (N_9927,N_9659,N_9460);
and U9928 (N_9928,N_9268,N_9685);
and U9929 (N_9929,N_9561,N_9414);
and U9930 (N_9930,N_9197,N_9477);
or U9931 (N_9931,N_9532,N_9418);
and U9932 (N_9932,N_9367,N_9621);
nor U9933 (N_9933,N_9141,N_9274);
and U9934 (N_9934,N_9485,N_9410);
and U9935 (N_9935,N_9396,N_9060);
nand U9936 (N_9936,N_9488,N_9512);
xor U9937 (N_9937,N_9429,N_9214);
nor U9938 (N_9938,N_9110,N_9352);
or U9939 (N_9939,N_9058,N_9606);
and U9940 (N_9940,N_9455,N_9251);
and U9941 (N_9941,N_9228,N_9432);
nor U9942 (N_9942,N_9198,N_9596);
nand U9943 (N_9943,N_9171,N_9346);
or U9944 (N_9944,N_9617,N_9051);
and U9945 (N_9945,N_9297,N_9364);
nor U9946 (N_9946,N_9092,N_9605);
and U9947 (N_9947,N_9588,N_9305);
or U9948 (N_9948,N_9121,N_9269);
nor U9949 (N_9949,N_9704,N_9296);
nand U9950 (N_9950,N_9543,N_9366);
nand U9951 (N_9951,N_9001,N_9133);
or U9952 (N_9952,N_9696,N_9011);
and U9953 (N_9953,N_9706,N_9053);
or U9954 (N_9954,N_9408,N_9355);
nand U9955 (N_9955,N_9316,N_9334);
or U9956 (N_9956,N_9061,N_9181);
or U9957 (N_9957,N_9469,N_9067);
or U9958 (N_9958,N_9336,N_9577);
or U9959 (N_9959,N_9162,N_9586);
xnor U9960 (N_9960,N_9124,N_9637);
nor U9961 (N_9961,N_9134,N_9495);
nand U9962 (N_9962,N_9379,N_9135);
or U9963 (N_9963,N_9231,N_9144);
or U9964 (N_9964,N_9513,N_9474);
or U9965 (N_9965,N_9341,N_9098);
or U9966 (N_9966,N_9224,N_9329);
or U9967 (N_9967,N_9264,N_9527);
nand U9968 (N_9968,N_9551,N_9007);
or U9969 (N_9969,N_9082,N_9667);
nor U9970 (N_9970,N_9576,N_9672);
nor U9971 (N_9971,N_9457,N_9105);
and U9972 (N_9972,N_9697,N_9199);
nor U9973 (N_9973,N_9564,N_9326);
nor U9974 (N_9974,N_9565,N_9523);
or U9975 (N_9975,N_9461,N_9454);
nand U9976 (N_9976,N_9314,N_9358);
nor U9977 (N_9977,N_9709,N_9106);
or U9978 (N_9978,N_9289,N_9002);
nor U9979 (N_9979,N_9368,N_9188);
or U9980 (N_9980,N_9203,N_9476);
xor U9981 (N_9981,N_9003,N_9318);
nor U9982 (N_9982,N_9047,N_9041);
nor U9983 (N_9983,N_9216,N_9234);
or U9984 (N_9984,N_9161,N_9616);
or U9985 (N_9985,N_9591,N_9650);
or U9986 (N_9986,N_9579,N_9028);
and U9987 (N_9987,N_9025,N_9032);
nand U9988 (N_9988,N_9365,N_9736);
nand U9989 (N_9989,N_9290,N_9384);
or U9990 (N_9990,N_9229,N_9747);
nor U9991 (N_9991,N_9540,N_9117);
xor U9992 (N_9992,N_9131,N_9087);
and U9993 (N_9993,N_9022,N_9128);
nor U9994 (N_9994,N_9715,N_9294);
and U9995 (N_9995,N_9475,N_9714);
nor U9996 (N_9996,N_9091,N_9407);
nor U9997 (N_9997,N_9446,N_9478);
nand U9998 (N_9998,N_9033,N_9727);
and U9999 (N_9999,N_9584,N_9275);
and U10000 (N_10000,N_9545,N_9323);
nor U10001 (N_10001,N_9307,N_9273);
or U10002 (N_10002,N_9102,N_9742);
nand U10003 (N_10003,N_9211,N_9518);
and U10004 (N_10004,N_9236,N_9713);
and U10005 (N_10005,N_9660,N_9501);
nor U10006 (N_10006,N_9260,N_9624);
nor U10007 (N_10007,N_9592,N_9598);
and U10008 (N_10008,N_9120,N_9244);
or U10009 (N_10009,N_9386,N_9026);
nand U10010 (N_10010,N_9479,N_9447);
and U10011 (N_10011,N_9093,N_9568);
or U10012 (N_10012,N_9589,N_9480);
or U10013 (N_10013,N_9021,N_9481);
xor U10014 (N_10014,N_9733,N_9272);
nor U10015 (N_10015,N_9127,N_9731);
and U10016 (N_10016,N_9103,N_9664);
or U10017 (N_10017,N_9441,N_9735);
and U10018 (N_10018,N_9466,N_9068);
and U10019 (N_10019,N_9238,N_9409);
xor U10020 (N_10020,N_9159,N_9417);
xor U10021 (N_10021,N_9607,N_9240);
nor U10022 (N_10022,N_9675,N_9701);
nand U10023 (N_10023,N_9676,N_9023);
nand U10024 (N_10024,N_9104,N_9506);
nand U10025 (N_10025,N_9692,N_9420);
nand U10026 (N_10026,N_9499,N_9335);
nor U10027 (N_10027,N_9339,N_9157);
xor U10028 (N_10028,N_9259,N_9009);
nor U10029 (N_10029,N_9178,N_9581);
xor U10030 (N_10030,N_9213,N_9378);
and U10031 (N_10031,N_9250,N_9623);
or U10032 (N_10032,N_9113,N_9380);
nand U10033 (N_10033,N_9340,N_9677);
nor U10034 (N_10034,N_9702,N_9048);
xnor U10035 (N_10035,N_9174,N_9717);
and U10036 (N_10036,N_9072,N_9657);
and U10037 (N_10037,N_9037,N_9403);
nand U10038 (N_10038,N_9629,N_9489);
nor U10039 (N_10039,N_9510,N_9711);
nand U10040 (N_10040,N_9375,N_9000);
or U10041 (N_10041,N_9004,N_9182);
or U10042 (N_10042,N_9331,N_9582);
or U10043 (N_10043,N_9600,N_9626);
or U10044 (N_10044,N_9287,N_9291);
or U10045 (N_10045,N_9107,N_9046);
nand U10046 (N_10046,N_9575,N_9387);
nand U10047 (N_10047,N_9652,N_9258);
or U10048 (N_10048,N_9030,N_9554);
nor U10049 (N_10049,N_9550,N_9207);
xnor U10050 (N_10050,N_9423,N_9641);
nor U10051 (N_10051,N_9362,N_9653);
and U10052 (N_10052,N_9167,N_9215);
or U10053 (N_10053,N_9679,N_9338);
or U10054 (N_10054,N_9559,N_9151);
nand U10055 (N_10055,N_9136,N_9630);
nand U10056 (N_10056,N_9078,N_9618);
and U10057 (N_10057,N_9373,N_9639);
nor U10058 (N_10058,N_9573,N_9737);
xor U10059 (N_10059,N_9376,N_9056);
or U10060 (N_10060,N_9017,N_9348);
and U10061 (N_10061,N_9094,N_9693);
nand U10062 (N_10062,N_9166,N_9321);
xnor U10063 (N_10063,N_9187,N_9099);
or U10064 (N_10064,N_9243,N_9266);
or U10065 (N_10065,N_9020,N_9360);
nor U10066 (N_10066,N_9448,N_9516);
or U10067 (N_10067,N_9249,N_9722);
and U10068 (N_10068,N_9643,N_9426);
or U10069 (N_10069,N_9651,N_9724);
nor U10070 (N_10070,N_9263,N_9114);
and U10071 (N_10071,N_9312,N_9218);
and U10072 (N_10072,N_9190,N_9125);
and U10073 (N_10073,N_9097,N_9718);
and U10074 (N_10074,N_9609,N_9688);
nor U10075 (N_10075,N_9492,N_9265);
nor U10076 (N_10076,N_9465,N_9220);
nor U10077 (N_10077,N_9085,N_9129);
nand U10078 (N_10078,N_9062,N_9283);
and U10079 (N_10079,N_9055,N_9317);
and U10080 (N_10080,N_9390,N_9018);
and U10081 (N_10081,N_9304,N_9563);
xor U10082 (N_10082,N_9108,N_9299);
and U10083 (N_10083,N_9741,N_9158);
nand U10084 (N_10084,N_9434,N_9086);
nor U10085 (N_10085,N_9324,N_9435);
and U10086 (N_10086,N_9552,N_9497);
and U10087 (N_10087,N_9156,N_9399);
xor U10088 (N_10088,N_9084,N_9726);
nand U10089 (N_10089,N_9595,N_9083);
or U10090 (N_10090,N_9520,N_9193);
nand U10091 (N_10091,N_9008,N_9130);
or U10092 (N_10092,N_9411,N_9282);
nand U10093 (N_10093,N_9361,N_9681);
and U10094 (N_10094,N_9080,N_9689);
xnor U10095 (N_10095,N_9433,N_9508);
and U10096 (N_10096,N_9690,N_9599);
nor U10097 (N_10097,N_9154,N_9632);
nand U10098 (N_10098,N_9148,N_9313);
nand U10099 (N_10099,N_9445,N_9645);
or U10100 (N_10100,N_9221,N_9456);
or U10101 (N_10101,N_9155,N_9468);
nand U10102 (N_10102,N_9438,N_9302);
nor U10103 (N_10103,N_9683,N_9646);
nand U10104 (N_10104,N_9548,N_9648);
and U10105 (N_10105,N_9279,N_9006);
nor U10106 (N_10106,N_9431,N_9118);
or U10107 (N_10107,N_9184,N_9308);
or U10108 (N_10108,N_9281,N_9401);
nor U10109 (N_10109,N_9089,N_9571);
xnor U10110 (N_10110,N_9647,N_9734);
or U10111 (N_10111,N_9674,N_9293);
or U10112 (N_10112,N_9716,N_9145);
nand U10113 (N_10113,N_9562,N_9077);
xor U10114 (N_10114,N_9491,N_9374);
nor U10115 (N_10115,N_9583,N_9529);
nand U10116 (N_10116,N_9442,N_9288);
nor U10117 (N_10117,N_9309,N_9278);
nor U10118 (N_10118,N_9405,N_9602);
nor U10119 (N_10119,N_9601,N_9634);
and U10120 (N_10120,N_9054,N_9458);
and U10121 (N_10121,N_9276,N_9535);
nor U10122 (N_10122,N_9116,N_9587);
and U10123 (N_10123,N_9295,N_9050);
or U10124 (N_10124,N_9670,N_9111);
nor U10125 (N_10125,N_9678,N_9356);
and U10126 (N_10126,N_9367,N_9315);
nand U10127 (N_10127,N_9347,N_9293);
nand U10128 (N_10128,N_9311,N_9527);
nand U10129 (N_10129,N_9573,N_9225);
xor U10130 (N_10130,N_9047,N_9435);
nor U10131 (N_10131,N_9273,N_9597);
nor U10132 (N_10132,N_9064,N_9329);
xnor U10133 (N_10133,N_9587,N_9726);
nand U10134 (N_10134,N_9500,N_9350);
or U10135 (N_10135,N_9273,N_9563);
xor U10136 (N_10136,N_9453,N_9571);
xnor U10137 (N_10137,N_9703,N_9695);
nand U10138 (N_10138,N_9567,N_9646);
nand U10139 (N_10139,N_9195,N_9689);
and U10140 (N_10140,N_9624,N_9245);
nor U10141 (N_10141,N_9063,N_9105);
nand U10142 (N_10142,N_9262,N_9320);
nand U10143 (N_10143,N_9230,N_9618);
or U10144 (N_10144,N_9733,N_9718);
nand U10145 (N_10145,N_9651,N_9111);
and U10146 (N_10146,N_9661,N_9333);
or U10147 (N_10147,N_9524,N_9197);
xnor U10148 (N_10148,N_9282,N_9274);
nand U10149 (N_10149,N_9707,N_9288);
nand U10150 (N_10150,N_9442,N_9627);
xnor U10151 (N_10151,N_9565,N_9129);
nor U10152 (N_10152,N_9641,N_9131);
nand U10153 (N_10153,N_9372,N_9701);
and U10154 (N_10154,N_9738,N_9361);
nor U10155 (N_10155,N_9555,N_9365);
and U10156 (N_10156,N_9445,N_9580);
and U10157 (N_10157,N_9322,N_9017);
nor U10158 (N_10158,N_9555,N_9224);
nand U10159 (N_10159,N_9129,N_9260);
or U10160 (N_10160,N_9681,N_9048);
and U10161 (N_10161,N_9467,N_9261);
nand U10162 (N_10162,N_9640,N_9702);
or U10163 (N_10163,N_9472,N_9453);
or U10164 (N_10164,N_9697,N_9223);
nand U10165 (N_10165,N_9172,N_9579);
nor U10166 (N_10166,N_9010,N_9433);
and U10167 (N_10167,N_9729,N_9346);
or U10168 (N_10168,N_9729,N_9517);
and U10169 (N_10169,N_9519,N_9647);
and U10170 (N_10170,N_9461,N_9144);
nand U10171 (N_10171,N_9553,N_9043);
nor U10172 (N_10172,N_9164,N_9732);
and U10173 (N_10173,N_9238,N_9429);
nor U10174 (N_10174,N_9155,N_9534);
or U10175 (N_10175,N_9244,N_9450);
and U10176 (N_10176,N_9550,N_9614);
and U10177 (N_10177,N_9559,N_9610);
or U10178 (N_10178,N_9039,N_9260);
or U10179 (N_10179,N_9289,N_9446);
nand U10180 (N_10180,N_9575,N_9150);
nor U10181 (N_10181,N_9415,N_9372);
nand U10182 (N_10182,N_9056,N_9658);
and U10183 (N_10183,N_9406,N_9228);
nand U10184 (N_10184,N_9407,N_9295);
or U10185 (N_10185,N_9240,N_9490);
and U10186 (N_10186,N_9114,N_9565);
or U10187 (N_10187,N_9520,N_9583);
nand U10188 (N_10188,N_9604,N_9247);
nand U10189 (N_10189,N_9594,N_9278);
or U10190 (N_10190,N_9178,N_9090);
or U10191 (N_10191,N_9491,N_9240);
nand U10192 (N_10192,N_9245,N_9644);
nand U10193 (N_10193,N_9429,N_9299);
nor U10194 (N_10194,N_9369,N_9499);
and U10195 (N_10195,N_9157,N_9712);
xnor U10196 (N_10196,N_9546,N_9118);
or U10197 (N_10197,N_9528,N_9280);
and U10198 (N_10198,N_9046,N_9350);
xnor U10199 (N_10199,N_9567,N_9280);
xor U10200 (N_10200,N_9271,N_9742);
xor U10201 (N_10201,N_9651,N_9714);
xnor U10202 (N_10202,N_9740,N_9138);
nor U10203 (N_10203,N_9748,N_9124);
xor U10204 (N_10204,N_9728,N_9726);
nand U10205 (N_10205,N_9371,N_9304);
and U10206 (N_10206,N_9089,N_9508);
and U10207 (N_10207,N_9677,N_9094);
nor U10208 (N_10208,N_9588,N_9576);
and U10209 (N_10209,N_9352,N_9153);
nand U10210 (N_10210,N_9614,N_9448);
and U10211 (N_10211,N_9576,N_9547);
or U10212 (N_10212,N_9504,N_9514);
xnor U10213 (N_10213,N_9375,N_9434);
nor U10214 (N_10214,N_9230,N_9193);
or U10215 (N_10215,N_9374,N_9520);
nor U10216 (N_10216,N_9732,N_9356);
and U10217 (N_10217,N_9151,N_9268);
and U10218 (N_10218,N_9181,N_9512);
and U10219 (N_10219,N_9388,N_9113);
nor U10220 (N_10220,N_9549,N_9683);
nand U10221 (N_10221,N_9290,N_9174);
and U10222 (N_10222,N_9211,N_9599);
or U10223 (N_10223,N_9224,N_9607);
nand U10224 (N_10224,N_9202,N_9533);
and U10225 (N_10225,N_9527,N_9728);
or U10226 (N_10226,N_9014,N_9621);
nor U10227 (N_10227,N_9713,N_9503);
nand U10228 (N_10228,N_9627,N_9446);
and U10229 (N_10229,N_9709,N_9579);
or U10230 (N_10230,N_9188,N_9559);
nor U10231 (N_10231,N_9733,N_9362);
and U10232 (N_10232,N_9127,N_9437);
nor U10233 (N_10233,N_9092,N_9157);
or U10234 (N_10234,N_9330,N_9042);
nand U10235 (N_10235,N_9014,N_9046);
or U10236 (N_10236,N_9367,N_9205);
or U10237 (N_10237,N_9041,N_9691);
nor U10238 (N_10238,N_9364,N_9663);
or U10239 (N_10239,N_9492,N_9539);
nor U10240 (N_10240,N_9299,N_9485);
nor U10241 (N_10241,N_9416,N_9559);
or U10242 (N_10242,N_9673,N_9274);
or U10243 (N_10243,N_9578,N_9482);
or U10244 (N_10244,N_9463,N_9513);
and U10245 (N_10245,N_9085,N_9407);
nor U10246 (N_10246,N_9027,N_9224);
and U10247 (N_10247,N_9748,N_9581);
and U10248 (N_10248,N_9453,N_9596);
nand U10249 (N_10249,N_9437,N_9277);
nor U10250 (N_10250,N_9493,N_9030);
or U10251 (N_10251,N_9572,N_9609);
and U10252 (N_10252,N_9219,N_9457);
or U10253 (N_10253,N_9200,N_9148);
xnor U10254 (N_10254,N_9466,N_9563);
or U10255 (N_10255,N_9693,N_9623);
nand U10256 (N_10256,N_9281,N_9460);
xor U10257 (N_10257,N_9637,N_9588);
or U10258 (N_10258,N_9321,N_9249);
or U10259 (N_10259,N_9504,N_9376);
xor U10260 (N_10260,N_9588,N_9418);
nand U10261 (N_10261,N_9687,N_9436);
nor U10262 (N_10262,N_9369,N_9245);
nand U10263 (N_10263,N_9609,N_9553);
nand U10264 (N_10264,N_9044,N_9579);
nor U10265 (N_10265,N_9705,N_9541);
nor U10266 (N_10266,N_9543,N_9635);
or U10267 (N_10267,N_9396,N_9491);
xor U10268 (N_10268,N_9285,N_9641);
nand U10269 (N_10269,N_9493,N_9264);
and U10270 (N_10270,N_9051,N_9191);
or U10271 (N_10271,N_9119,N_9490);
and U10272 (N_10272,N_9473,N_9018);
xnor U10273 (N_10273,N_9453,N_9480);
or U10274 (N_10274,N_9457,N_9122);
nor U10275 (N_10275,N_9372,N_9273);
or U10276 (N_10276,N_9382,N_9103);
nor U10277 (N_10277,N_9196,N_9330);
nand U10278 (N_10278,N_9202,N_9666);
xnor U10279 (N_10279,N_9285,N_9615);
nor U10280 (N_10280,N_9702,N_9479);
nor U10281 (N_10281,N_9561,N_9180);
nand U10282 (N_10282,N_9258,N_9541);
nand U10283 (N_10283,N_9258,N_9186);
and U10284 (N_10284,N_9063,N_9290);
nor U10285 (N_10285,N_9168,N_9210);
or U10286 (N_10286,N_9510,N_9706);
and U10287 (N_10287,N_9288,N_9510);
nand U10288 (N_10288,N_9032,N_9694);
or U10289 (N_10289,N_9296,N_9267);
nand U10290 (N_10290,N_9260,N_9390);
or U10291 (N_10291,N_9062,N_9318);
and U10292 (N_10292,N_9004,N_9120);
or U10293 (N_10293,N_9224,N_9231);
nand U10294 (N_10294,N_9269,N_9217);
nand U10295 (N_10295,N_9719,N_9009);
nand U10296 (N_10296,N_9182,N_9469);
and U10297 (N_10297,N_9216,N_9303);
and U10298 (N_10298,N_9176,N_9666);
nor U10299 (N_10299,N_9692,N_9615);
nand U10300 (N_10300,N_9637,N_9714);
nor U10301 (N_10301,N_9552,N_9147);
or U10302 (N_10302,N_9329,N_9679);
or U10303 (N_10303,N_9293,N_9690);
or U10304 (N_10304,N_9635,N_9146);
and U10305 (N_10305,N_9406,N_9125);
nand U10306 (N_10306,N_9199,N_9020);
nor U10307 (N_10307,N_9038,N_9746);
nand U10308 (N_10308,N_9448,N_9188);
and U10309 (N_10309,N_9634,N_9664);
nand U10310 (N_10310,N_9088,N_9636);
nand U10311 (N_10311,N_9259,N_9717);
and U10312 (N_10312,N_9657,N_9636);
xnor U10313 (N_10313,N_9366,N_9349);
nor U10314 (N_10314,N_9177,N_9645);
nor U10315 (N_10315,N_9239,N_9300);
nor U10316 (N_10316,N_9365,N_9078);
nor U10317 (N_10317,N_9747,N_9246);
nor U10318 (N_10318,N_9598,N_9165);
and U10319 (N_10319,N_9281,N_9739);
nor U10320 (N_10320,N_9512,N_9705);
nor U10321 (N_10321,N_9538,N_9670);
and U10322 (N_10322,N_9426,N_9465);
nor U10323 (N_10323,N_9592,N_9331);
and U10324 (N_10324,N_9474,N_9455);
or U10325 (N_10325,N_9262,N_9376);
and U10326 (N_10326,N_9095,N_9727);
nand U10327 (N_10327,N_9400,N_9503);
or U10328 (N_10328,N_9718,N_9400);
xor U10329 (N_10329,N_9025,N_9489);
nand U10330 (N_10330,N_9293,N_9037);
and U10331 (N_10331,N_9345,N_9142);
and U10332 (N_10332,N_9407,N_9563);
and U10333 (N_10333,N_9191,N_9699);
nand U10334 (N_10334,N_9016,N_9235);
nand U10335 (N_10335,N_9176,N_9094);
and U10336 (N_10336,N_9181,N_9133);
and U10337 (N_10337,N_9177,N_9260);
nand U10338 (N_10338,N_9148,N_9330);
xor U10339 (N_10339,N_9068,N_9244);
xor U10340 (N_10340,N_9456,N_9162);
xor U10341 (N_10341,N_9723,N_9222);
or U10342 (N_10342,N_9074,N_9456);
or U10343 (N_10343,N_9315,N_9691);
or U10344 (N_10344,N_9208,N_9246);
and U10345 (N_10345,N_9112,N_9318);
nor U10346 (N_10346,N_9232,N_9120);
nor U10347 (N_10347,N_9171,N_9452);
or U10348 (N_10348,N_9488,N_9490);
or U10349 (N_10349,N_9200,N_9481);
nand U10350 (N_10350,N_9262,N_9719);
nand U10351 (N_10351,N_9067,N_9497);
nand U10352 (N_10352,N_9144,N_9400);
and U10353 (N_10353,N_9016,N_9194);
nand U10354 (N_10354,N_9248,N_9615);
or U10355 (N_10355,N_9076,N_9738);
nand U10356 (N_10356,N_9619,N_9066);
or U10357 (N_10357,N_9694,N_9072);
or U10358 (N_10358,N_9305,N_9391);
nand U10359 (N_10359,N_9454,N_9073);
nor U10360 (N_10360,N_9573,N_9309);
nor U10361 (N_10361,N_9683,N_9059);
or U10362 (N_10362,N_9028,N_9559);
xor U10363 (N_10363,N_9749,N_9399);
and U10364 (N_10364,N_9490,N_9682);
and U10365 (N_10365,N_9098,N_9533);
or U10366 (N_10366,N_9089,N_9307);
nand U10367 (N_10367,N_9283,N_9481);
nor U10368 (N_10368,N_9366,N_9033);
nor U10369 (N_10369,N_9615,N_9086);
nor U10370 (N_10370,N_9562,N_9299);
and U10371 (N_10371,N_9237,N_9715);
or U10372 (N_10372,N_9436,N_9738);
nand U10373 (N_10373,N_9649,N_9401);
or U10374 (N_10374,N_9123,N_9125);
or U10375 (N_10375,N_9452,N_9238);
nand U10376 (N_10376,N_9066,N_9141);
nor U10377 (N_10377,N_9749,N_9675);
nor U10378 (N_10378,N_9630,N_9400);
nand U10379 (N_10379,N_9525,N_9468);
nand U10380 (N_10380,N_9046,N_9467);
nand U10381 (N_10381,N_9242,N_9183);
or U10382 (N_10382,N_9448,N_9072);
and U10383 (N_10383,N_9302,N_9527);
xnor U10384 (N_10384,N_9536,N_9704);
xor U10385 (N_10385,N_9470,N_9218);
nor U10386 (N_10386,N_9679,N_9237);
nor U10387 (N_10387,N_9461,N_9409);
or U10388 (N_10388,N_9479,N_9213);
and U10389 (N_10389,N_9485,N_9060);
xnor U10390 (N_10390,N_9217,N_9117);
nor U10391 (N_10391,N_9164,N_9380);
nor U10392 (N_10392,N_9716,N_9283);
nand U10393 (N_10393,N_9587,N_9341);
or U10394 (N_10394,N_9135,N_9245);
nand U10395 (N_10395,N_9011,N_9410);
xnor U10396 (N_10396,N_9537,N_9744);
nor U10397 (N_10397,N_9019,N_9520);
xnor U10398 (N_10398,N_9540,N_9572);
nor U10399 (N_10399,N_9714,N_9040);
nand U10400 (N_10400,N_9574,N_9031);
or U10401 (N_10401,N_9378,N_9396);
or U10402 (N_10402,N_9442,N_9496);
nor U10403 (N_10403,N_9352,N_9294);
or U10404 (N_10404,N_9665,N_9152);
and U10405 (N_10405,N_9227,N_9293);
xnor U10406 (N_10406,N_9703,N_9258);
nand U10407 (N_10407,N_9575,N_9512);
or U10408 (N_10408,N_9111,N_9425);
and U10409 (N_10409,N_9074,N_9415);
and U10410 (N_10410,N_9202,N_9640);
and U10411 (N_10411,N_9284,N_9399);
or U10412 (N_10412,N_9208,N_9404);
or U10413 (N_10413,N_9435,N_9417);
and U10414 (N_10414,N_9125,N_9059);
xnor U10415 (N_10415,N_9405,N_9310);
nand U10416 (N_10416,N_9298,N_9692);
and U10417 (N_10417,N_9203,N_9171);
or U10418 (N_10418,N_9352,N_9034);
or U10419 (N_10419,N_9216,N_9096);
and U10420 (N_10420,N_9291,N_9003);
nor U10421 (N_10421,N_9241,N_9104);
and U10422 (N_10422,N_9348,N_9354);
nand U10423 (N_10423,N_9623,N_9316);
and U10424 (N_10424,N_9523,N_9491);
nor U10425 (N_10425,N_9174,N_9671);
nand U10426 (N_10426,N_9523,N_9247);
nand U10427 (N_10427,N_9550,N_9626);
nor U10428 (N_10428,N_9424,N_9594);
or U10429 (N_10429,N_9167,N_9525);
nand U10430 (N_10430,N_9559,N_9545);
xnor U10431 (N_10431,N_9207,N_9690);
nor U10432 (N_10432,N_9645,N_9256);
or U10433 (N_10433,N_9161,N_9651);
nor U10434 (N_10434,N_9321,N_9502);
and U10435 (N_10435,N_9360,N_9744);
nor U10436 (N_10436,N_9528,N_9406);
or U10437 (N_10437,N_9507,N_9151);
and U10438 (N_10438,N_9310,N_9276);
and U10439 (N_10439,N_9332,N_9671);
and U10440 (N_10440,N_9253,N_9472);
or U10441 (N_10441,N_9587,N_9677);
xnor U10442 (N_10442,N_9044,N_9532);
nor U10443 (N_10443,N_9063,N_9671);
or U10444 (N_10444,N_9724,N_9509);
or U10445 (N_10445,N_9302,N_9656);
nor U10446 (N_10446,N_9625,N_9217);
and U10447 (N_10447,N_9419,N_9465);
nand U10448 (N_10448,N_9723,N_9123);
nand U10449 (N_10449,N_9163,N_9437);
nand U10450 (N_10450,N_9433,N_9538);
nand U10451 (N_10451,N_9339,N_9174);
and U10452 (N_10452,N_9546,N_9491);
and U10453 (N_10453,N_9690,N_9356);
nor U10454 (N_10454,N_9358,N_9375);
nor U10455 (N_10455,N_9222,N_9102);
or U10456 (N_10456,N_9571,N_9530);
nor U10457 (N_10457,N_9422,N_9658);
nor U10458 (N_10458,N_9261,N_9536);
and U10459 (N_10459,N_9127,N_9497);
or U10460 (N_10460,N_9182,N_9517);
xor U10461 (N_10461,N_9092,N_9469);
nand U10462 (N_10462,N_9365,N_9718);
or U10463 (N_10463,N_9662,N_9655);
nor U10464 (N_10464,N_9031,N_9616);
or U10465 (N_10465,N_9013,N_9451);
nor U10466 (N_10466,N_9720,N_9364);
xor U10467 (N_10467,N_9173,N_9179);
or U10468 (N_10468,N_9196,N_9296);
and U10469 (N_10469,N_9368,N_9682);
and U10470 (N_10470,N_9010,N_9657);
nor U10471 (N_10471,N_9632,N_9337);
nor U10472 (N_10472,N_9481,N_9601);
nor U10473 (N_10473,N_9548,N_9292);
nor U10474 (N_10474,N_9601,N_9327);
nand U10475 (N_10475,N_9439,N_9634);
nor U10476 (N_10476,N_9339,N_9417);
xnor U10477 (N_10477,N_9134,N_9411);
and U10478 (N_10478,N_9597,N_9539);
nand U10479 (N_10479,N_9573,N_9634);
or U10480 (N_10480,N_9496,N_9545);
nand U10481 (N_10481,N_9064,N_9388);
or U10482 (N_10482,N_9437,N_9550);
and U10483 (N_10483,N_9183,N_9147);
and U10484 (N_10484,N_9519,N_9440);
and U10485 (N_10485,N_9143,N_9710);
or U10486 (N_10486,N_9046,N_9580);
nand U10487 (N_10487,N_9477,N_9035);
or U10488 (N_10488,N_9245,N_9705);
and U10489 (N_10489,N_9412,N_9129);
and U10490 (N_10490,N_9506,N_9591);
and U10491 (N_10491,N_9481,N_9237);
nand U10492 (N_10492,N_9037,N_9185);
and U10493 (N_10493,N_9005,N_9447);
and U10494 (N_10494,N_9344,N_9342);
or U10495 (N_10495,N_9116,N_9428);
nor U10496 (N_10496,N_9696,N_9136);
nand U10497 (N_10497,N_9450,N_9673);
nor U10498 (N_10498,N_9010,N_9569);
or U10499 (N_10499,N_9098,N_9609);
or U10500 (N_10500,N_10270,N_10202);
xnor U10501 (N_10501,N_10470,N_10387);
and U10502 (N_10502,N_10115,N_10171);
nand U10503 (N_10503,N_9801,N_10004);
nor U10504 (N_10504,N_10277,N_10183);
and U10505 (N_10505,N_10136,N_10335);
or U10506 (N_10506,N_10355,N_10449);
nor U10507 (N_10507,N_10426,N_9880);
nand U10508 (N_10508,N_10305,N_10489);
or U10509 (N_10509,N_10460,N_9833);
or U10510 (N_10510,N_9988,N_9889);
and U10511 (N_10511,N_9952,N_10195);
and U10512 (N_10512,N_9793,N_10349);
or U10513 (N_10513,N_9873,N_10315);
nor U10514 (N_10514,N_10022,N_10000);
or U10515 (N_10515,N_10238,N_10239);
nand U10516 (N_10516,N_10056,N_9967);
nand U10517 (N_10517,N_10257,N_10256);
or U10518 (N_10518,N_10247,N_10416);
nor U10519 (N_10519,N_9807,N_10274);
nand U10520 (N_10520,N_10401,N_9887);
nor U10521 (N_10521,N_9893,N_10388);
or U10522 (N_10522,N_10142,N_9787);
or U10523 (N_10523,N_10437,N_10495);
nor U10524 (N_10524,N_10095,N_10389);
nor U10525 (N_10525,N_9957,N_9827);
and U10526 (N_10526,N_9817,N_9913);
nor U10527 (N_10527,N_10366,N_9914);
or U10528 (N_10528,N_10310,N_10243);
and U10529 (N_10529,N_9795,N_10353);
and U10530 (N_10530,N_9768,N_10396);
or U10531 (N_10531,N_10427,N_9978);
nand U10532 (N_10532,N_10032,N_10314);
nor U10533 (N_10533,N_10438,N_10329);
and U10534 (N_10534,N_9916,N_10258);
and U10535 (N_10535,N_10473,N_10161);
xor U10536 (N_10536,N_10205,N_10128);
nand U10537 (N_10537,N_10444,N_10230);
and U10538 (N_10538,N_9792,N_9941);
nand U10539 (N_10539,N_10367,N_10319);
nand U10540 (N_10540,N_9810,N_10178);
xnor U10541 (N_10541,N_10499,N_10420);
nor U10542 (N_10542,N_10005,N_10244);
nor U10543 (N_10543,N_10200,N_9970);
nand U10544 (N_10544,N_9861,N_9750);
nor U10545 (N_10545,N_10141,N_9960);
xor U10546 (N_10546,N_10359,N_10053);
nor U10547 (N_10547,N_9896,N_10098);
or U10548 (N_10548,N_9879,N_9797);
xnor U10549 (N_10549,N_10482,N_10446);
nand U10550 (N_10550,N_9919,N_10198);
or U10551 (N_10551,N_10370,N_9975);
xnor U10552 (N_10552,N_9777,N_9942);
nand U10553 (N_10553,N_10307,N_9950);
or U10554 (N_10554,N_10155,N_10260);
nand U10555 (N_10555,N_9872,N_10087);
and U10556 (N_10556,N_10113,N_10081);
and U10557 (N_10557,N_9876,N_9943);
xor U10558 (N_10558,N_10386,N_9951);
and U10559 (N_10559,N_9858,N_10273);
xor U10560 (N_10560,N_10292,N_9806);
or U10561 (N_10561,N_9830,N_10408);
nor U10562 (N_10562,N_10413,N_9969);
nor U10563 (N_10563,N_9984,N_9865);
nor U10564 (N_10564,N_10104,N_10042);
nor U10565 (N_10565,N_9869,N_9963);
nor U10566 (N_10566,N_10333,N_10368);
and U10567 (N_10567,N_10194,N_9771);
nor U10568 (N_10568,N_10397,N_10031);
xor U10569 (N_10569,N_10044,N_10174);
nand U10570 (N_10570,N_9853,N_9953);
nand U10571 (N_10571,N_10160,N_10447);
nor U10572 (N_10572,N_10210,N_10463);
nor U10573 (N_10573,N_10085,N_10207);
or U10574 (N_10574,N_10219,N_9832);
and U10575 (N_10575,N_9915,N_10334);
nor U10576 (N_10576,N_10414,N_10491);
nand U10577 (N_10577,N_10126,N_10191);
nand U10578 (N_10578,N_10124,N_10343);
nand U10579 (N_10579,N_9757,N_10279);
nand U10580 (N_10580,N_9995,N_9874);
or U10581 (N_10581,N_10094,N_9881);
nor U10582 (N_10582,N_9979,N_10357);
nor U10583 (N_10583,N_10203,N_9791);
or U10584 (N_10584,N_9997,N_9905);
nand U10585 (N_10585,N_9985,N_10339);
nor U10586 (N_10586,N_9994,N_9839);
nor U10587 (N_10587,N_9760,N_10372);
nor U10588 (N_10588,N_10129,N_9980);
nor U10589 (N_10589,N_10430,N_9933);
nand U10590 (N_10590,N_10362,N_10132);
nand U10591 (N_10591,N_10208,N_10336);
and U10592 (N_10592,N_10411,N_10045);
nand U10593 (N_10593,N_9931,N_10278);
nand U10594 (N_10594,N_9772,N_10046);
nand U10595 (N_10595,N_9877,N_10285);
nor U10596 (N_10596,N_10309,N_9849);
nand U10597 (N_10597,N_9909,N_10109);
or U10598 (N_10598,N_9822,N_10096);
or U10599 (N_10599,N_9770,N_10374);
or U10600 (N_10600,N_10140,N_9815);
nor U10601 (N_10601,N_10267,N_10209);
or U10602 (N_10602,N_10035,N_9785);
and U10603 (N_10603,N_10373,N_9870);
nor U10604 (N_10604,N_10297,N_9821);
or U10605 (N_10605,N_10454,N_10488);
and U10606 (N_10606,N_10262,N_10007);
or U10607 (N_10607,N_10240,N_10189);
or U10608 (N_10608,N_10119,N_10120);
nor U10609 (N_10609,N_10296,N_10330);
or U10610 (N_10610,N_10038,N_9754);
and U10611 (N_10611,N_10407,N_10047);
nand U10612 (N_10612,N_9856,N_9888);
nand U10613 (N_10613,N_10057,N_10102);
and U10614 (N_10614,N_10347,N_10168);
nand U10615 (N_10615,N_9912,N_10254);
and U10616 (N_10616,N_10400,N_9867);
xnor U10617 (N_10617,N_9945,N_10215);
xnor U10618 (N_10618,N_10114,N_9751);
nand U10619 (N_10619,N_9819,N_10105);
or U10620 (N_10620,N_9923,N_10139);
or U10621 (N_10621,N_10301,N_10332);
and U10622 (N_10622,N_10293,N_10058);
and U10623 (N_10623,N_9904,N_9886);
nor U10624 (N_10624,N_9755,N_10423);
or U10625 (N_10625,N_9940,N_9983);
or U10626 (N_10626,N_9971,N_9902);
and U10627 (N_10627,N_9925,N_10322);
or U10628 (N_10628,N_10013,N_10036);
nor U10629 (N_10629,N_9884,N_10276);
nand U10630 (N_10630,N_9911,N_9929);
and U10631 (N_10631,N_10037,N_10049);
nor U10632 (N_10632,N_10172,N_10006);
nand U10633 (N_10633,N_10492,N_10398);
nor U10634 (N_10634,N_9901,N_9938);
xnor U10635 (N_10635,N_9993,N_10497);
nor U10636 (N_10636,N_10375,N_10421);
xnor U10637 (N_10637,N_10030,N_10227);
nand U10638 (N_10638,N_10248,N_10312);
nor U10639 (N_10639,N_9762,N_10441);
nand U10640 (N_10640,N_9966,N_10148);
nand U10641 (N_10641,N_10442,N_10236);
nor U10642 (N_10642,N_10402,N_10064);
nand U10643 (N_10643,N_9763,N_10253);
nor U10644 (N_10644,N_10241,N_10364);
xor U10645 (N_10645,N_10014,N_9972);
nor U10646 (N_10646,N_10299,N_10156);
and U10647 (N_10647,N_10121,N_10275);
nand U10648 (N_10648,N_10212,N_10061);
xnor U10649 (N_10649,N_10453,N_9859);
nand U10650 (N_10650,N_10452,N_10471);
and U10651 (N_10651,N_9855,N_9835);
nand U10652 (N_10652,N_10425,N_10249);
and U10653 (N_10653,N_10079,N_9885);
or U10654 (N_10654,N_10196,N_10050);
and U10655 (N_10655,N_9934,N_10108);
or U10656 (N_10656,N_10147,N_10481);
nor U10657 (N_10657,N_10154,N_10478);
and U10658 (N_10658,N_10010,N_10218);
xor U10659 (N_10659,N_10112,N_10034);
nand U10660 (N_10660,N_9803,N_10487);
and U10661 (N_10661,N_10175,N_9774);
or U10662 (N_10662,N_10327,N_10484);
and U10663 (N_10663,N_10211,N_10251);
or U10664 (N_10664,N_10180,N_10237);
and U10665 (N_10665,N_10226,N_10342);
and U10666 (N_10666,N_9955,N_9823);
nor U10667 (N_10667,N_10476,N_10229);
xnor U10668 (N_10668,N_9898,N_10451);
nand U10669 (N_10669,N_10039,N_9782);
nor U10670 (N_10670,N_10371,N_10068);
nand U10671 (N_10671,N_10158,N_10077);
nor U10672 (N_10672,N_9899,N_9977);
or U10673 (N_10673,N_10135,N_10479);
or U10674 (N_10674,N_10418,N_9892);
nand U10675 (N_10675,N_9799,N_10067);
xnor U10676 (N_10676,N_9965,N_9878);
nand U10677 (N_10677,N_10337,N_10358);
and U10678 (N_10678,N_10019,N_10001);
and U10679 (N_10679,N_10341,N_9820);
nor U10680 (N_10680,N_10338,N_10252);
xnor U10681 (N_10681,N_9761,N_9783);
nor U10682 (N_10682,N_9753,N_9825);
or U10683 (N_10683,N_10016,N_10026);
or U10684 (N_10684,N_9800,N_9860);
and U10685 (N_10685,N_10093,N_10302);
nor U10686 (N_10686,N_10151,N_10048);
and U10687 (N_10687,N_9921,N_9779);
nand U10688 (N_10688,N_10385,N_10092);
or U10689 (N_10689,N_9780,N_10179);
nand U10690 (N_10690,N_10163,N_10352);
and U10691 (N_10691,N_10281,N_10410);
and U10692 (N_10692,N_10106,N_9922);
nand U10693 (N_10693,N_9805,N_9852);
nand U10694 (N_10694,N_10246,N_10440);
nor U10695 (N_10695,N_10474,N_9796);
nand U10696 (N_10696,N_10103,N_9842);
xor U10697 (N_10697,N_10023,N_9949);
nand U10698 (N_10698,N_10055,N_9834);
or U10699 (N_10699,N_10231,N_10138);
or U10700 (N_10700,N_10017,N_10433);
and U10701 (N_10701,N_10214,N_10008);
or U10702 (N_10702,N_10417,N_10321);
or U10703 (N_10703,N_9871,N_10284);
and U10704 (N_10704,N_9890,N_10043);
nor U10705 (N_10705,N_9811,N_10477);
and U10706 (N_10706,N_9866,N_9851);
and U10707 (N_10707,N_10428,N_10080);
xnor U10708 (N_10708,N_9891,N_9818);
nor U10709 (N_10709,N_10261,N_10294);
and U10710 (N_10710,N_10395,N_10025);
nand U10711 (N_10711,N_10369,N_9790);
and U10712 (N_10712,N_10378,N_10271);
nor U10713 (N_10713,N_10409,N_9764);
nand U10714 (N_10714,N_10099,N_9864);
nand U10715 (N_10715,N_10146,N_9927);
nor U10716 (N_10716,N_10286,N_10118);
nor U10717 (N_10717,N_10197,N_10117);
nor U10718 (N_10718,N_10051,N_10456);
xnor U10719 (N_10719,N_10110,N_9895);
and U10720 (N_10720,N_10265,N_10468);
nor U10721 (N_10721,N_10176,N_10165);
or U10722 (N_10722,N_10455,N_9986);
or U10723 (N_10723,N_10052,N_10394);
nor U10724 (N_10724,N_10065,N_10062);
or U10725 (N_10725,N_10266,N_10496);
nand U10726 (N_10726,N_10101,N_9981);
nand U10727 (N_10727,N_10054,N_10184);
and U10728 (N_10728,N_9778,N_10439);
or U10729 (N_10729,N_9808,N_9752);
or U10730 (N_10730,N_10199,N_9917);
xnor U10731 (N_10731,N_10066,N_10340);
xnor U10732 (N_10732,N_9918,N_10018);
nand U10733 (N_10733,N_10003,N_9784);
or U10734 (N_10734,N_9857,N_9926);
and U10735 (N_10735,N_10193,N_10072);
or U10736 (N_10736,N_10268,N_10134);
xor U10737 (N_10737,N_9845,N_10185);
nand U10738 (N_10738,N_10393,N_10328);
nand U10739 (N_10739,N_9840,N_10224);
xor U10740 (N_10740,N_9765,N_9798);
nand U10741 (N_10741,N_9850,N_10177);
nor U10742 (N_10742,N_9767,N_10429);
and U10743 (N_10743,N_10269,N_10461);
nand U10744 (N_10744,N_10075,N_9946);
nor U10745 (N_10745,N_9920,N_9990);
nor U10746 (N_10746,N_10405,N_10311);
and U10747 (N_10747,N_9862,N_10404);
or U10748 (N_10748,N_10498,N_10221);
xor U10749 (N_10749,N_9837,N_10071);
nor U10750 (N_10750,N_10318,N_10377);
nor U10751 (N_10751,N_10325,N_9958);
xnor U10752 (N_10752,N_10348,N_9847);
or U10753 (N_10753,N_10084,N_10308);
nor U10754 (N_10754,N_9907,N_9826);
or U10755 (N_10755,N_10291,N_10091);
or U10756 (N_10756,N_10365,N_9908);
nor U10757 (N_10757,N_10028,N_10317);
nand U10758 (N_10758,N_10033,N_10467);
nand U10759 (N_10759,N_10169,N_10263);
nand U10760 (N_10760,N_9814,N_9848);
nand U10761 (N_10761,N_10070,N_10458);
and U10762 (N_10762,N_10020,N_10152);
nand U10763 (N_10763,N_10272,N_9991);
or U10764 (N_10764,N_9900,N_9935);
nor U10765 (N_10765,N_10086,N_10345);
nand U10766 (N_10766,N_10406,N_10344);
and U10767 (N_10767,N_9846,N_9996);
and U10768 (N_10768,N_10173,N_9776);
or U10769 (N_10769,N_9956,N_9910);
and U10770 (N_10770,N_10331,N_9936);
or U10771 (N_10771,N_10107,N_9831);
nor U10772 (N_10772,N_9989,N_10379);
or U10773 (N_10773,N_9947,N_10116);
nand U10774 (N_10774,N_9992,N_9903);
nand U10775 (N_10775,N_9794,N_9843);
and U10776 (N_10776,N_9781,N_9944);
xor U10777 (N_10777,N_10204,N_10029);
nand U10778 (N_10778,N_10242,N_9786);
and U10779 (N_10779,N_10100,N_9804);
or U10780 (N_10780,N_9788,N_10384);
or U10781 (N_10781,N_10153,N_10361);
nor U10782 (N_10782,N_10445,N_10475);
and U10783 (N_10783,N_10354,N_9829);
and U10784 (N_10784,N_9968,N_10181);
or U10785 (N_10785,N_9836,N_9883);
or U10786 (N_10786,N_9863,N_10078);
and U10787 (N_10787,N_9759,N_10376);
and U10788 (N_10788,N_10448,N_9906);
nand U10789 (N_10789,N_10351,N_9882);
nand U10790 (N_10790,N_9932,N_10422);
and U10791 (N_10791,N_10002,N_10295);
nor U10792 (N_10792,N_10415,N_10381);
nor U10793 (N_10793,N_10245,N_10490);
nand U10794 (N_10794,N_10316,N_9789);
nand U10795 (N_10795,N_10186,N_10290);
nand U10796 (N_10796,N_10125,N_10466);
nand U10797 (N_10797,N_9838,N_10346);
xor U10798 (N_10798,N_9775,N_10465);
nand U10799 (N_10799,N_9964,N_10063);
xor U10800 (N_10800,N_10170,N_10123);
xor U10801 (N_10801,N_10187,N_10073);
nand U10802 (N_10802,N_10360,N_10289);
nand U10803 (N_10803,N_10419,N_10060);
nor U10804 (N_10804,N_10083,N_9813);
and U10805 (N_10805,N_9868,N_10304);
nor U10806 (N_10806,N_10356,N_10233);
or U10807 (N_10807,N_10391,N_10399);
xnor U10808 (N_10808,N_9824,N_10443);
nand U10809 (N_10809,N_10166,N_9875);
nand U10810 (N_10810,N_10090,N_10216);
nor U10811 (N_10811,N_10076,N_10283);
nor U10812 (N_10812,N_9841,N_10074);
nor U10813 (N_10813,N_10167,N_10288);
or U10814 (N_10814,N_10350,N_10024);
nor U10815 (N_10815,N_9959,N_10225);
or U10816 (N_10816,N_10082,N_10015);
nand U10817 (N_10817,N_9854,N_10383);
xnor U10818 (N_10818,N_9894,N_9769);
or U10819 (N_10819,N_10464,N_9758);
xor U10820 (N_10820,N_10059,N_10469);
and U10821 (N_10821,N_9961,N_10259);
nand U10822 (N_10822,N_10303,N_10127);
nand U10823 (N_10823,N_10457,N_9974);
and U10824 (N_10824,N_10217,N_10235);
or U10825 (N_10825,N_10150,N_10392);
nor U10826 (N_10826,N_10232,N_10213);
nand U10827 (N_10827,N_10201,N_10264);
and U10828 (N_10828,N_10012,N_10472);
xor U10829 (N_10829,N_10390,N_10041);
nand U10830 (N_10830,N_10403,N_10190);
nor U10831 (N_10831,N_10250,N_9939);
or U10832 (N_10832,N_10220,N_9962);
and U10833 (N_10833,N_9828,N_9773);
nor U10834 (N_10834,N_9998,N_9954);
nand U10835 (N_10835,N_10122,N_10111);
or U10836 (N_10836,N_10228,N_10144);
nand U10837 (N_10837,N_10040,N_9976);
and U10838 (N_10838,N_10450,N_9937);
or U10839 (N_10839,N_10088,N_10382);
nor U10840 (N_10840,N_9973,N_10192);
nor U10841 (N_10841,N_10222,N_10486);
nor U10842 (N_10842,N_9924,N_10432);
nor U10843 (N_10843,N_10280,N_10069);
nand U10844 (N_10844,N_10133,N_10326);
xnor U10845 (N_10845,N_10424,N_10089);
and U10846 (N_10846,N_10097,N_10320);
nand U10847 (N_10847,N_10157,N_10412);
xnor U10848 (N_10848,N_9766,N_10435);
or U10849 (N_10849,N_9948,N_9928);
nor U10850 (N_10850,N_10011,N_10483);
or U10851 (N_10851,N_10431,N_10143);
xor U10852 (N_10852,N_10306,N_10182);
nor U10853 (N_10853,N_10459,N_10313);
nand U10854 (N_10854,N_10282,N_9756);
nand U10855 (N_10855,N_9809,N_10494);
nor U10856 (N_10856,N_10434,N_10324);
nor U10857 (N_10857,N_10223,N_9999);
nor U10858 (N_10858,N_10188,N_10323);
and U10859 (N_10859,N_9982,N_10363);
and U10860 (N_10860,N_10462,N_10480);
or U10861 (N_10861,N_10021,N_9930);
nor U10862 (N_10862,N_10485,N_9816);
xnor U10863 (N_10863,N_10137,N_10164);
nor U10864 (N_10864,N_9844,N_10206);
nor U10865 (N_10865,N_10131,N_9897);
xnor U10866 (N_10866,N_10436,N_10149);
and U10867 (N_10867,N_9802,N_10380);
xnor U10868 (N_10868,N_10300,N_10255);
nand U10869 (N_10869,N_10287,N_10145);
or U10870 (N_10870,N_10027,N_10298);
nor U10871 (N_10871,N_10162,N_10009);
or U10872 (N_10872,N_10234,N_9987);
xor U10873 (N_10873,N_10130,N_10493);
nand U10874 (N_10874,N_10159,N_9812);
and U10875 (N_10875,N_9930,N_10156);
xor U10876 (N_10876,N_9868,N_10027);
nand U10877 (N_10877,N_10198,N_9884);
nor U10878 (N_10878,N_9873,N_10023);
and U10879 (N_10879,N_10225,N_10153);
or U10880 (N_10880,N_10097,N_10252);
nor U10881 (N_10881,N_9837,N_9752);
nor U10882 (N_10882,N_10233,N_10000);
nor U10883 (N_10883,N_10288,N_10346);
and U10884 (N_10884,N_10197,N_9829);
nand U10885 (N_10885,N_9989,N_9803);
or U10886 (N_10886,N_10144,N_10480);
or U10887 (N_10887,N_9817,N_10119);
and U10888 (N_10888,N_9850,N_9835);
nor U10889 (N_10889,N_9787,N_10223);
or U10890 (N_10890,N_10137,N_9930);
or U10891 (N_10891,N_10293,N_9972);
nor U10892 (N_10892,N_9910,N_10213);
or U10893 (N_10893,N_9913,N_10493);
nand U10894 (N_10894,N_10181,N_9826);
or U10895 (N_10895,N_9812,N_10135);
or U10896 (N_10896,N_9908,N_9942);
and U10897 (N_10897,N_10414,N_10422);
and U10898 (N_10898,N_9788,N_10399);
or U10899 (N_10899,N_9909,N_10233);
or U10900 (N_10900,N_9933,N_10234);
nand U10901 (N_10901,N_9999,N_10018);
nor U10902 (N_10902,N_9786,N_10442);
nor U10903 (N_10903,N_10287,N_9912);
nand U10904 (N_10904,N_10424,N_10452);
nor U10905 (N_10905,N_10240,N_10010);
or U10906 (N_10906,N_9984,N_9900);
and U10907 (N_10907,N_10085,N_10113);
nand U10908 (N_10908,N_9835,N_10321);
nor U10909 (N_10909,N_10085,N_10328);
and U10910 (N_10910,N_9841,N_10473);
or U10911 (N_10911,N_9859,N_10333);
and U10912 (N_10912,N_10054,N_10003);
or U10913 (N_10913,N_10219,N_10276);
or U10914 (N_10914,N_9984,N_9850);
nor U10915 (N_10915,N_10026,N_10268);
or U10916 (N_10916,N_10363,N_10139);
nor U10917 (N_10917,N_9852,N_10186);
or U10918 (N_10918,N_10285,N_9990);
or U10919 (N_10919,N_9965,N_9876);
nor U10920 (N_10920,N_9998,N_10375);
nor U10921 (N_10921,N_10284,N_9773);
or U10922 (N_10922,N_10129,N_10290);
nor U10923 (N_10923,N_10174,N_10327);
or U10924 (N_10924,N_9884,N_10208);
nor U10925 (N_10925,N_10157,N_10133);
or U10926 (N_10926,N_9813,N_10470);
nand U10927 (N_10927,N_10080,N_10325);
xnor U10928 (N_10928,N_10047,N_10326);
or U10929 (N_10929,N_9950,N_10110);
and U10930 (N_10930,N_10460,N_9901);
and U10931 (N_10931,N_10379,N_10479);
xor U10932 (N_10932,N_10245,N_10443);
xnor U10933 (N_10933,N_10134,N_10272);
nor U10934 (N_10934,N_10423,N_10068);
or U10935 (N_10935,N_9950,N_9956);
nor U10936 (N_10936,N_10192,N_10053);
and U10937 (N_10937,N_9991,N_9862);
or U10938 (N_10938,N_10180,N_10069);
nand U10939 (N_10939,N_10463,N_9986);
or U10940 (N_10940,N_9913,N_10205);
and U10941 (N_10941,N_9975,N_9810);
and U10942 (N_10942,N_9878,N_10059);
and U10943 (N_10943,N_9874,N_10074);
or U10944 (N_10944,N_10143,N_10390);
nor U10945 (N_10945,N_10188,N_10394);
xor U10946 (N_10946,N_9873,N_10125);
or U10947 (N_10947,N_9893,N_10185);
and U10948 (N_10948,N_9935,N_10003);
or U10949 (N_10949,N_10145,N_10261);
and U10950 (N_10950,N_9956,N_9851);
nor U10951 (N_10951,N_9808,N_9922);
nand U10952 (N_10952,N_10245,N_10243);
nand U10953 (N_10953,N_10442,N_10448);
or U10954 (N_10954,N_10053,N_9990);
nor U10955 (N_10955,N_9879,N_10264);
nor U10956 (N_10956,N_10380,N_10032);
or U10957 (N_10957,N_9768,N_9774);
and U10958 (N_10958,N_10110,N_9893);
xor U10959 (N_10959,N_10327,N_9938);
nand U10960 (N_10960,N_9890,N_10451);
or U10961 (N_10961,N_10322,N_10216);
or U10962 (N_10962,N_9867,N_9839);
and U10963 (N_10963,N_9933,N_10116);
nor U10964 (N_10964,N_10138,N_9770);
xnor U10965 (N_10965,N_10282,N_10459);
nand U10966 (N_10966,N_10042,N_10145);
nand U10967 (N_10967,N_9831,N_9859);
and U10968 (N_10968,N_9979,N_10125);
nor U10969 (N_10969,N_9964,N_9956);
nand U10970 (N_10970,N_10397,N_10111);
and U10971 (N_10971,N_9825,N_9788);
xor U10972 (N_10972,N_10303,N_10089);
xor U10973 (N_10973,N_10220,N_10074);
or U10974 (N_10974,N_10271,N_9853);
nand U10975 (N_10975,N_10421,N_9775);
nand U10976 (N_10976,N_10433,N_10058);
or U10977 (N_10977,N_10015,N_10141);
nor U10978 (N_10978,N_9919,N_9797);
nor U10979 (N_10979,N_10277,N_10444);
and U10980 (N_10980,N_10439,N_10194);
or U10981 (N_10981,N_10279,N_9837);
or U10982 (N_10982,N_10262,N_10037);
xnor U10983 (N_10983,N_10089,N_10160);
or U10984 (N_10984,N_10376,N_10343);
or U10985 (N_10985,N_10475,N_10054);
and U10986 (N_10986,N_10472,N_10370);
nor U10987 (N_10987,N_10268,N_10355);
nand U10988 (N_10988,N_9787,N_9906);
nand U10989 (N_10989,N_9974,N_10375);
and U10990 (N_10990,N_9960,N_9949);
nor U10991 (N_10991,N_9980,N_10090);
or U10992 (N_10992,N_10481,N_10346);
and U10993 (N_10993,N_10379,N_10294);
or U10994 (N_10994,N_10400,N_9800);
and U10995 (N_10995,N_10127,N_10189);
nor U10996 (N_10996,N_10275,N_10016);
nand U10997 (N_10997,N_9813,N_10221);
or U10998 (N_10998,N_9896,N_10456);
nor U10999 (N_10999,N_10020,N_10433);
nand U11000 (N_11000,N_9955,N_9910);
nand U11001 (N_11001,N_10318,N_10218);
or U11002 (N_11002,N_10355,N_10455);
or U11003 (N_11003,N_10258,N_10286);
or U11004 (N_11004,N_9920,N_9817);
nand U11005 (N_11005,N_10295,N_10007);
or U11006 (N_11006,N_9799,N_10235);
nand U11007 (N_11007,N_9975,N_9988);
nand U11008 (N_11008,N_10315,N_10442);
nand U11009 (N_11009,N_10214,N_10065);
or U11010 (N_11010,N_10061,N_10369);
and U11011 (N_11011,N_9784,N_10092);
nor U11012 (N_11012,N_10321,N_10054);
xnor U11013 (N_11013,N_9923,N_9790);
and U11014 (N_11014,N_10001,N_10486);
or U11015 (N_11015,N_9869,N_10248);
nor U11016 (N_11016,N_9945,N_10409);
nand U11017 (N_11017,N_9837,N_10350);
and U11018 (N_11018,N_10225,N_10087);
or U11019 (N_11019,N_9835,N_9758);
nand U11020 (N_11020,N_10420,N_9810);
nor U11021 (N_11021,N_10047,N_10107);
or U11022 (N_11022,N_10291,N_10462);
or U11023 (N_11023,N_10140,N_9891);
nor U11024 (N_11024,N_10244,N_10359);
and U11025 (N_11025,N_10184,N_10327);
nand U11026 (N_11026,N_10105,N_10238);
nor U11027 (N_11027,N_10425,N_10014);
nor U11028 (N_11028,N_10250,N_10024);
and U11029 (N_11029,N_9995,N_9927);
and U11030 (N_11030,N_9920,N_10134);
and U11031 (N_11031,N_10058,N_9817);
nand U11032 (N_11032,N_10480,N_10196);
or U11033 (N_11033,N_10072,N_10225);
or U11034 (N_11034,N_10027,N_10230);
or U11035 (N_11035,N_9965,N_9886);
or U11036 (N_11036,N_10040,N_10098);
or U11037 (N_11037,N_10040,N_10283);
nand U11038 (N_11038,N_10446,N_10421);
nor U11039 (N_11039,N_10371,N_10182);
or U11040 (N_11040,N_10400,N_10286);
nor U11041 (N_11041,N_10380,N_9779);
or U11042 (N_11042,N_10097,N_9948);
or U11043 (N_11043,N_10028,N_10067);
or U11044 (N_11044,N_9980,N_10230);
and U11045 (N_11045,N_10004,N_10248);
xnor U11046 (N_11046,N_9795,N_9810);
or U11047 (N_11047,N_9889,N_10269);
or U11048 (N_11048,N_9971,N_10365);
or U11049 (N_11049,N_9971,N_10386);
nand U11050 (N_11050,N_10115,N_10144);
and U11051 (N_11051,N_9878,N_10388);
xnor U11052 (N_11052,N_10412,N_10097);
nand U11053 (N_11053,N_9991,N_10271);
xnor U11054 (N_11054,N_10279,N_10030);
nand U11055 (N_11055,N_10058,N_10077);
nor U11056 (N_11056,N_10476,N_10233);
nand U11057 (N_11057,N_10212,N_10098);
xor U11058 (N_11058,N_9892,N_10137);
or U11059 (N_11059,N_10421,N_10155);
and U11060 (N_11060,N_10136,N_10404);
or U11061 (N_11061,N_10196,N_9929);
and U11062 (N_11062,N_9939,N_10193);
nor U11063 (N_11063,N_10402,N_10285);
nor U11064 (N_11064,N_9963,N_10221);
or U11065 (N_11065,N_10183,N_10481);
nand U11066 (N_11066,N_10292,N_9750);
xnor U11067 (N_11067,N_10164,N_10323);
nand U11068 (N_11068,N_10387,N_10059);
nor U11069 (N_11069,N_9994,N_10290);
nor U11070 (N_11070,N_10470,N_10168);
or U11071 (N_11071,N_9840,N_10035);
nand U11072 (N_11072,N_9949,N_10245);
or U11073 (N_11073,N_9956,N_10294);
nor U11074 (N_11074,N_10092,N_9982);
and U11075 (N_11075,N_10491,N_10019);
nand U11076 (N_11076,N_10343,N_10109);
nor U11077 (N_11077,N_10039,N_10000);
or U11078 (N_11078,N_10495,N_10178);
nand U11079 (N_11079,N_9860,N_9880);
and U11080 (N_11080,N_9898,N_10395);
nand U11081 (N_11081,N_10426,N_9953);
or U11082 (N_11082,N_10207,N_9955);
nor U11083 (N_11083,N_10161,N_10373);
and U11084 (N_11084,N_9894,N_10297);
and U11085 (N_11085,N_9761,N_9975);
or U11086 (N_11086,N_9970,N_10380);
or U11087 (N_11087,N_10315,N_10069);
and U11088 (N_11088,N_9966,N_9793);
or U11089 (N_11089,N_9859,N_9974);
nand U11090 (N_11090,N_10323,N_10076);
nor U11091 (N_11091,N_9991,N_10139);
and U11092 (N_11092,N_9813,N_10317);
nor U11093 (N_11093,N_9857,N_9936);
nand U11094 (N_11094,N_10036,N_10136);
or U11095 (N_11095,N_10369,N_10084);
xnor U11096 (N_11096,N_9982,N_9903);
and U11097 (N_11097,N_10348,N_9806);
nor U11098 (N_11098,N_10076,N_9875);
nor U11099 (N_11099,N_10290,N_10130);
nor U11100 (N_11100,N_10094,N_9877);
or U11101 (N_11101,N_10060,N_10204);
and U11102 (N_11102,N_10233,N_10228);
nor U11103 (N_11103,N_10477,N_10249);
and U11104 (N_11104,N_9834,N_9865);
xor U11105 (N_11105,N_10151,N_9827);
or U11106 (N_11106,N_10345,N_9880);
nor U11107 (N_11107,N_10048,N_9930);
nor U11108 (N_11108,N_10420,N_10096);
nor U11109 (N_11109,N_10030,N_10003);
or U11110 (N_11110,N_9855,N_9939);
nor U11111 (N_11111,N_9919,N_9920);
and U11112 (N_11112,N_9809,N_9979);
nand U11113 (N_11113,N_9790,N_10286);
nand U11114 (N_11114,N_10381,N_10001);
and U11115 (N_11115,N_10051,N_10198);
nor U11116 (N_11116,N_10067,N_10431);
nand U11117 (N_11117,N_10102,N_9959);
nand U11118 (N_11118,N_10184,N_9827);
xnor U11119 (N_11119,N_10399,N_10453);
or U11120 (N_11120,N_10197,N_10438);
and U11121 (N_11121,N_10069,N_10325);
nand U11122 (N_11122,N_10192,N_10201);
or U11123 (N_11123,N_9787,N_10192);
nor U11124 (N_11124,N_10475,N_9886);
or U11125 (N_11125,N_9859,N_10395);
xor U11126 (N_11126,N_10458,N_9839);
or U11127 (N_11127,N_10253,N_10029);
or U11128 (N_11128,N_10372,N_10333);
nand U11129 (N_11129,N_10447,N_9886);
nor U11130 (N_11130,N_10402,N_9907);
and U11131 (N_11131,N_9776,N_10286);
and U11132 (N_11132,N_10106,N_10292);
nand U11133 (N_11133,N_9783,N_10108);
nor U11134 (N_11134,N_10021,N_10422);
nor U11135 (N_11135,N_9854,N_10363);
nor U11136 (N_11136,N_10103,N_10249);
and U11137 (N_11137,N_10490,N_10191);
nand U11138 (N_11138,N_10343,N_10106);
nand U11139 (N_11139,N_10442,N_10106);
and U11140 (N_11140,N_9896,N_10499);
and U11141 (N_11141,N_10219,N_10418);
nor U11142 (N_11142,N_10021,N_10454);
or U11143 (N_11143,N_10209,N_10396);
nor U11144 (N_11144,N_10210,N_10221);
or U11145 (N_11145,N_9830,N_9951);
nor U11146 (N_11146,N_9779,N_10051);
nor U11147 (N_11147,N_9777,N_10219);
nand U11148 (N_11148,N_10187,N_10120);
and U11149 (N_11149,N_10110,N_9909);
and U11150 (N_11150,N_10086,N_9984);
nand U11151 (N_11151,N_9921,N_9974);
nor U11152 (N_11152,N_10360,N_10116);
xor U11153 (N_11153,N_10213,N_10150);
nor U11154 (N_11154,N_9803,N_10413);
or U11155 (N_11155,N_10484,N_9781);
and U11156 (N_11156,N_10350,N_9768);
and U11157 (N_11157,N_10304,N_10368);
and U11158 (N_11158,N_10200,N_10333);
or U11159 (N_11159,N_10414,N_10120);
xnor U11160 (N_11160,N_10191,N_9907);
and U11161 (N_11161,N_9801,N_10093);
nand U11162 (N_11162,N_10356,N_9831);
and U11163 (N_11163,N_10117,N_9866);
nor U11164 (N_11164,N_10078,N_10135);
nor U11165 (N_11165,N_10146,N_9825);
and U11166 (N_11166,N_10186,N_10193);
and U11167 (N_11167,N_9992,N_10037);
and U11168 (N_11168,N_10401,N_9847);
and U11169 (N_11169,N_10492,N_10093);
and U11170 (N_11170,N_10354,N_10285);
and U11171 (N_11171,N_10071,N_10106);
and U11172 (N_11172,N_10350,N_10101);
and U11173 (N_11173,N_10286,N_10049);
nand U11174 (N_11174,N_10060,N_9806);
and U11175 (N_11175,N_9893,N_10072);
xor U11176 (N_11176,N_9996,N_9861);
nand U11177 (N_11177,N_9789,N_10337);
nor U11178 (N_11178,N_10482,N_9986);
nor U11179 (N_11179,N_10259,N_9944);
xor U11180 (N_11180,N_9756,N_10314);
xnor U11181 (N_11181,N_10090,N_9846);
xnor U11182 (N_11182,N_10296,N_10344);
and U11183 (N_11183,N_9940,N_10021);
and U11184 (N_11184,N_9819,N_10284);
nand U11185 (N_11185,N_10170,N_9995);
nand U11186 (N_11186,N_9779,N_9871);
or U11187 (N_11187,N_9917,N_10097);
xor U11188 (N_11188,N_10013,N_10413);
nand U11189 (N_11189,N_10022,N_10036);
and U11190 (N_11190,N_9943,N_10123);
or U11191 (N_11191,N_9831,N_9931);
and U11192 (N_11192,N_9944,N_9915);
nor U11193 (N_11193,N_10334,N_9852);
nand U11194 (N_11194,N_9994,N_10387);
nor U11195 (N_11195,N_9831,N_10005);
and U11196 (N_11196,N_10098,N_9893);
nor U11197 (N_11197,N_10344,N_10163);
and U11198 (N_11198,N_10259,N_10278);
and U11199 (N_11199,N_10418,N_9802);
nor U11200 (N_11200,N_10411,N_9893);
and U11201 (N_11201,N_10459,N_10203);
and U11202 (N_11202,N_10216,N_10142);
nand U11203 (N_11203,N_10387,N_9792);
or U11204 (N_11204,N_10198,N_10234);
nand U11205 (N_11205,N_10289,N_10343);
or U11206 (N_11206,N_10184,N_9902);
and U11207 (N_11207,N_10370,N_10050);
or U11208 (N_11208,N_9957,N_10409);
nor U11209 (N_11209,N_10378,N_10082);
xnor U11210 (N_11210,N_9837,N_10317);
nand U11211 (N_11211,N_10256,N_10244);
nand U11212 (N_11212,N_9810,N_10394);
or U11213 (N_11213,N_9902,N_9944);
nor U11214 (N_11214,N_10485,N_10175);
and U11215 (N_11215,N_10440,N_10133);
and U11216 (N_11216,N_9934,N_9990);
and U11217 (N_11217,N_10393,N_9842);
nor U11218 (N_11218,N_10369,N_9771);
nand U11219 (N_11219,N_10176,N_10291);
nand U11220 (N_11220,N_10426,N_10472);
nor U11221 (N_11221,N_10302,N_10088);
nor U11222 (N_11222,N_9987,N_10065);
nand U11223 (N_11223,N_10470,N_9992);
and U11224 (N_11224,N_10068,N_9993);
and U11225 (N_11225,N_9905,N_9907);
nor U11226 (N_11226,N_10468,N_10410);
nor U11227 (N_11227,N_10341,N_10206);
nor U11228 (N_11228,N_10124,N_9991);
or U11229 (N_11229,N_10429,N_10202);
nand U11230 (N_11230,N_10245,N_9779);
xor U11231 (N_11231,N_10210,N_10418);
xnor U11232 (N_11232,N_10379,N_10003);
and U11233 (N_11233,N_9935,N_10103);
or U11234 (N_11234,N_10455,N_10481);
or U11235 (N_11235,N_10083,N_10269);
and U11236 (N_11236,N_9867,N_9972);
nor U11237 (N_11237,N_10402,N_10379);
or U11238 (N_11238,N_10317,N_9989);
or U11239 (N_11239,N_9815,N_10356);
xnor U11240 (N_11240,N_10184,N_10268);
or U11241 (N_11241,N_10406,N_10103);
xnor U11242 (N_11242,N_10446,N_9879);
or U11243 (N_11243,N_10240,N_10388);
or U11244 (N_11244,N_10408,N_10344);
and U11245 (N_11245,N_10385,N_9850);
nor U11246 (N_11246,N_10480,N_9938);
and U11247 (N_11247,N_9871,N_10058);
nor U11248 (N_11248,N_10055,N_10479);
nand U11249 (N_11249,N_10355,N_10388);
or U11250 (N_11250,N_10813,N_10727);
or U11251 (N_11251,N_11039,N_10565);
or U11252 (N_11252,N_11116,N_10633);
or U11253 (N_11253,N_10780,N_10882);
nor U11254 (N_11254,N_11122,N_10522);
nor U11255 (N_11255,N_11031,N_10975);
nand U11256 (N_11256,N_10541,N_10993);
nand U11257 (N_11257,N_10763,N_10619);
nor U11258 (N_11258,N_11146,N_10746);
and U11259 (N_11259,N_10737,N_10970);
xnor U11260 (N_11260,N_10659,N_10538);
nor U11261 (N_11261,N_10706,N_11075);
or U11262 (N_11262,N_10604,N_10969);
or U11263 (N_11263,N_10729,N_10535);
or U11264 (N_11264,N_10556,N_10733);
or U11265 (N_11265,N_10503,N_11103);
nand U11266 (N_11266,N_10918,N_11248);
and U11267 (N_11267,N_11038,N_10721);
or U11268 (N_11268,N_10516,N_10870);
or U11269 (N_11269,N_10548,N_11026);
nand U11270 (N_11270,N_10759,N_10853);
nor U11271 (N_11271,N_10812,N_10952);
nand U11272 (N_11272,N_10588,N_11180);
or U11273 (N_11273,N_10521,N_11048);
xnor U11274 (N_11274,N_10893,N_11136);
nand U11275 (N_11275,N_11092,N_10776);
or U11276 (N_11276,N_11037,N_10640);
and U11277 (N_11277,N_10719,N_11137);
or U11278 (N_11278,N_10520,N_10947);
or U11279 (N_11279,N_10898,N_11174);
nand U11280 (N_11280,N_10753,N_10740);
or U11281 (N_11281,N_11047,N_11155);
and U11282 (N_11282,N_10707,N_10809);
nand U11283 (N_11283,N_10515,N_11093);
nand U11284 (N_11284,N_10666,N_10713);
nand U11285 (N_11285,N_10816,N_11023);
nor U11286 (N_11286,N_10747,N_10803);
and U11287 (N_11287,N_10658,N_11040);
and U11288 (N_11288,N_11134,N_11114);
and U11289 (N_11289,N_10940,N_11125);
or U11290 (N_11290,N_11034,N_10547);
and U11291 (N_11291,N_11020,N_10755);
nor U11292 (N_11292,N_10966,N_10814);
or U11293 (N_11293,N_11132,N_11220);
nand U11294 (N_11294,N_10656,N_10980);
and U11295 (N_11295,N_11097,N_11249);
nand U11296 (N_11296,N_11215,N_11107);
and U11297 (N_11297,N_10766,N_10684);
nor U11298 (N_11298,N_10871,N_10907);
nor U11299 (N_11299,N_10900,N_10828);
and U11300 (N_11300,N_10876,N_10630);
nor U11301 (N_11301,N_10854,N_11230);
or U11302 (N_11302,N_10661,N_10800);
nor U11303 (N_11303,N_11153,N_11113);
and U11304 (N_11304,N_11140,N_10601);
nor U11305 (N_11305,N_11007,N_10745);
or U11306 (N_11306,N_11193,N_10612);
or U11307 (N_11307,N_11124,N_11123);
nand U11308 (N_11308,N_11160,N_11130);
or U11309 (N_11309,N_11211,N_10892);
nand U11310 (N_11310,N_10570,N_10978);
and U11311 (N_11311,N_10829,N_11086);
nand U11312 (N_11312,N_10883,N_10714);
or U11313 (N_11313,N_11110,N_10916);
nor U11314 (N_11314,N_10586,N_10956);
and U11315 (N_11315,N_10960,N_11027);
nor U11316 (N_11316,N_10525,N_11012);
and U11317 (N_11317,N_11005,N_10648);
nor U11318 (N_11318,N_10912,N_10678);
or U11319 (N_11319,N_11222,N_11147);
nand U11320 (N_11320,N_10996,N_11170);
nand U11321 (N_11321,N_10873,N_10575);
nand U11322 (N_11322,N_11043,N_10577);
nor U11323 (N_11323,N_11120,N_11068);
nand U11324 (N_11324,N_10815,N_10731);
or U11325 (N_11325,N_10657,N_10668);
or U11326 (N_11326,N_11176,N_11212);
xnor U11327 (N_11327,N_11008,N_10518);
or U11328 (N_11328,N_10616,N_10781);
nor U11329 (N_11329,N_11101,N_10748);
nor U11330 (N_11330,N_10810,N_10880);
nor U11331 (N_11331,N_10506,N_10514);
nand U11332 (N_11332,N_10718,N_10942);
or U11333 (N_11333,N_10935,N_10730);
and U11334 (N_11334,N_10574,N_11017);
or U11335 (N_11335,N_10885,N_10700);
nand U11336 (N_11336,N_10712,N_10624);
and U11337 (N_11337,N_11002,N_10922);
and U11338 (N_11338,N_11148,N_11121);
and U11339 (N_11339,N_11221,N_10799);
or U11340 (N_11340,N_10894,N_11161);
or U11341 (N_11341,N_11219,N_10910);
and U11342 (N_11342,N_10599,N_10953);
or U11343 (N_11343,N_11083,N_10724);
nor U11344 (N_11344,N_11003,N_10569);
or U11345 (N_11345,N_11033,N_10795);
nor U11346 (N_11346,N_11018,N_10777);
xor U11347 (N_11347,N_10558,N_11173);
nor U11348 (N_11348,N_10682,N_10929);
or U11349 (N_11349,N_10536,N_10673);
nand U11350 (N_11350,N_10618,N_11213);
nor U11351 (N_11351,N_11025,N_11228);
nor U11352 (N_11352,N_10895,N_10505);
nor U11353 (N_11353,N_10623,N_10842);
nor U11354 (N_11354,N_11057,N_10634);
and U11355 (N_11355,N_11157,N_10797);
nand U11356 (N_11356,N_11062,N_11142);
nor U11357 (N_11357,N_10621,N_10778);
or U11358 (N_11358,N_10819,N_10647);
nor U11359 (N_11359,N_10787,N_10957);
and U11360 (N_11360,N_10717,N_11090);
and U11361 (N_11361,N_11095,N_10651);
nor U11362 (N_11362,N_10664,N_10944);
and U11363 (N_11363,N_10836,N_10632);
or U11364 (N_11364,N_11245,N_10674);
or U11365 (N_11365,N_10627,N_10681);
or U11366 (N_11366,N_10686,N_11001);
nor U11367 (N_11367,N_10846,N_11060);
xnor U11368 (N_11368,N_10702,N_10841);
nor U11369 (N_11369,N_10961,N_11016);
and U11370 (N_11370,N_10923,N_10798);
xor U11371 (N_11371,N_10555,N_11227);
nor U11372 (N_11372,N_10560,N_11195);
and U11373 (N_11373,N_10948,N_10637);
nand U11374 (N_11374,N_11183,N_11021);
xor U11375 (N_11375,N_10524,N_10999);
nand U11376 (N_11376,N_10594,N_10915);
xor U11377 (N_11377,N_11158,N_10603);
xnor U11378 (N_11378,N_11079,N_10869);
nand U11379 (N_11379,N_10597,N_10789);
or U11380 (N_11380,N_10862,N_11013);
and U11381 (N_11381,N_10790,N_10844);
nand U11382 (N_11382,N_11128,N_10550);
and U11383 (N_11383,N_10954,N_10701);
and U11384 (N_11384,N_10742,N_11105);
or U11385 (N_11385,N_11156,N_10582);
or U11386 (N_11386,N_10711,N_10551);
nor U11387 (N_11387,N_10765,N_11085);
or U11388 (N_11388,N_11196,N_11131);
and U11389 (N_11389,N_11035,N_11081);
and U11390 (N_11390,N_10855,N_10704);
or U11391 (N_11391,N_10868,N_11053);
or U11392 (N_11392,N_11224,N_10509);
or U11393 (N_11393,N_10553,N_10972);
nand U11394 (N_11394,N_10584,N_10937);
nand U11395 (N_11395,N_10794,N_10734);
or U11396 (N_11396,N_10965,N_11056);
nor U11397 (N_11397,N_10533,N_10866);
and U11398 (N_11398,N_10650,N_10938);
or U11399 (N_11399,N_11202,N_10837);
xnor U11400 (N_11400,N_10840,N_10884);
and U11401 (N_11401,N_11169,N_11238);
or U11402 (N_11402,N_11192,N_11234);
nand U11403 (N_11403,N_10585,N_11045);
xnor U11404 (N_11404,N_10826,N_10743);
nor U11405 (N_11405,N_10901,N_10615);
and U11406 (N_11406,N_10693,N_11209);
and U11407 (N_11407,N_10971,N_10998);
nor U11408 (N_11408,N_11189,N_10926);
and U11409 (N_11409,N_10783,N_10824);
nor U11410 (N_11410,N_10654,N_11135);
or U11411 (N_11411,N_10888,N_11139);
and U11412 (N_11412,N_10631,N_11054);
or U11413 (N_11413,N_10958,N_10517);
or U11414 (N_11414,N_10874,N_11190);
or U11415 (N_11415,N_10950,N_10967);
nand U11416 (N_11416,N_10646,N_11076);
nand U11417 (N_11417,N_11077,N_11216);
or U11418 (N_11418,N_10908,N_11091);
nand U11419 (N_11419,N_10739,N_10825);
or U11420 (N_11420,N_11150,N_10990);
nor U11421 (N_11421,N_10580,N_11127);
or U11422 (N_11422,N_11009,N_10896);
nor U11423 (N_11423,N_10987,N_10641);
or U11424 (N_11424,N_10775,N_10904);
and U11425 (N_11425,N_10933,N_10663);
or U11426 (N_11426,N_10749,N_11080);
and U11427 (N_11427,N_10504,N_11100);
or U11428 (N_11428,N_10939,N_11214);
or U11429 (N_11429,N_10802,N_10848);
and U11430 (N_11430,N_10757,N_10767);
or U11431 (N_11431,N_10690,N_10576);
or U11432 (N_11432,N_11171,N_10805);
nand U11433 (N_11433,N_11066,N_10983);
nand U11434 (N_11434,N_11164,N_10692);
nor U11435 (N_11435,N_10531,N_11032);
nand U11436 (N_11436,N_10530,N_10823);
or U11437 (N_11437,N_10644,N_10608);
nand U11438 (N_11438,N_10583,N_10566);
and U11439 (N_11439,N_10986,N_10741);
and U11440 (N_11440,N_10736,N_10785);
xor U11441 (N_11441,N_11232,N_11145);
nor U11442 (N_11442,N_10500,N_11204);
or U11443 (N_11443,N_10512,N_10716);
nand U11444 (N_11444,N_10914,N_11236);
and U11445 (N_11445,N_11197,N_11072);
and U11446 (N_11446,N_10924,N_10930);
or U11447 (N_11447,N_10945,N_10527);
nor U11448 (N_11448,N_10979,N_10807);
and U11449 (N_11449,N_10697,N_10959);
xor U11450 (N_11450,N_10784,N_11200);
and U11451 (N_11451,N_11133,N_11041);
xor U11452 (N_11452,N_10911,N_10991);
and U11453 (N_11453,N_10542,N_10688);
and U11454 (N_11454,N_10699,N_10786);
nor U11455 (N_11455,N_11205,N_10773);
or U11456 (N_11456,N_11098,N_11179);
nor U11457 (N_11457,N_10887,N_10984);
nand U11458 (N_11458,N_10595,N_11186);
xor U11459 (N_11459,N_10501,N_11225);
xnor U11460 (N_11460,N_10642,N_10528);
nand U11461 (N_11461,N_11050,N_11203);
and U11462 (N_11462,N_10897,N_10662);
nand U11463 (N_11463,N_10720,N_10859);
or U11464 (N_11464,N_10562,N_10981);
nand U11465 (N_11465,N_10899,N_11069);
nor U11466 (N_11466,N_10994,N_10683);
nand U11467 (N_11467,N_11104,N_10903);
or U11468 (N_11468,N_10564,N_10863);
nand U11469 (N_11469,N_10964,N_10593);
nand U11470 (N_11470,N_10913,N_10665);
nand U11471 (N_11471,N_11089,N_10676);
nand U11472 (N_11472,N_10610,N_10818);
or U11473 (N_11473,N_10974,N_10635);
nand U11474 (N_11474,N_11096,N_10968);
or U11475 (N_11475,N_11094,N_10526);
or U11476 (N_11476,N_10928,N_11108);
nor U11477 (N_11477,N_11051,N_11210);
nand U11478 (N_11478,N_11118,N_11244);
and U11479 (N_11479,N_10620,N_10936);
xor U11480 (N_11480,N_10507,N_11078);
nor U11481 (N_11481,N_10833,N_11182);
and U11482 (N_11482,N_10796,N_10756);
nor U11483 (N_11483,N_11058,N_10817);
nor U11484 (N_11484,N_10614,N_10687);
nand U11485 (N_11485,N_10752,N_10949);
and U11486 (N_11486,N_11191,N_11082);
and U11487 (N_11487,N_11199,N_10804);
xor U11488 (N_11488,N_11006,N_11198);
and U11489 (N_11489,N_10587,N_10617);
or U11490 (N_11490,N_10625,N_10792);
and U11491 (N_11491,N_10502,N_10544);
or U11492 (N_11492,N_10579,N_10605);
nand U11493 (N_11493,N_10590,N_11099);
and U11494 (N_11494,N_10639,N_11052);
xor U11495 (N_11495,N_10955,N_11181);
nor U11496 (N_11496,N_10529,N_11119);
nor U11497 (N_11497,N_10649,N_10875);
nand U11498 (N_11498,N_10655,N_10689);
nor U11499 (N_11499,N_10925,N_11177);
nor U11500 (N_11500,N_10782,N_10976);
nand U11501 (N_11501,N_11102,N_10744);
nor U11502 (N_11502,N_11242,N_10951);
and U11503 (N_11503,N_11109,N_10638);
xnor U11504 (N_11504,N_11106,N_10801);
xnor U11505 (N_11505,N_11046,N_11172);
nor U11506 (N_11506,N_10667,N_11055);
nand U11507 (N_11507,N_10758,N_10738);
nor U11508 (N_11508,N_11159,N_10771);
nand U11509 (N_11509,N_10698,N_11014);
xnor U11510 (N_11510,N_10572,N_10872);
nand U11511 (N_11511,N_10806,N_10852);
or U11512 (N_11512,N_10920,N_11246);
nand U11513 (N_11513,N_11241,N_10890);
nand U11514 (N_11514,N_10629,N_10760);
nor U11515 (N_11515,N_10578,N_10754);
nand U11516 (N_11516,N_10679,N_10830);
or U11517 (N_11517,N_10857,N_10653);
and U11518 (N_11518,N_10680,N_11201);
and U11519 (N_11519,N_10573,N_10858);
or U11520 (N_11520,N_10877,N_10927);
or U11521 (N_11521,N_11024,N_10723);
nor U11522 (N_11522,N_11154,N_10879);
nor U11523 (N_11523,N_10710,N_10675);
nor U11524 (N_11524,N_10865,N_10772);
and U11525 (N_11525,N_10670,N_10768);
xnor U11526 (N_11526,N_11117,N_10695);
nor U11527 (N_11527,N_10808,N_10660);
and U11528 (N_11528,N_10946,N_10669);
nor U11529 (N_11529,N_10891,N_11071);
xor U11530 (N_11530,N_10581,N_11028);
or U11531 (N_11531,N_10793,N_10596);
xnor U11532 (N_11532,N_10609,N_10820);
nand U11533 (N_11533,N_10561,N_11070);
or U11534 (N_11534,N_10557,N_11141);
or U11535 (N_11535,N_10791,N_11152);
nand U11536 (N_11536,N_11064,N_10537);
nand U11537 (N_11537,N_11187,N_11088);
nand U11538 (N_11538,N_10510,N_10691);
nor U11539 (N_11539,N_10864,N_11087);
xor U11540 (N_11540,N_10932,N_11044);
or U11541 (N_11541,N_10788,N_10636);
or U11542 (N_11542,N_10770,N_10889);
nand U11543 (N_11543,N_10628,N_10532);
nor U11544 (N_11544,N_10671,N_10977);
xnor U11545 (N_11545,N_11239,N_10821);
or U11546 (N_11546,N_10705,N_11184);
nand U11547 (N_11547,N_10769,N_11111);
nor U11548 (N_11548,N_11067,N_10921);
xor U11549 (N_11549,N_11175,N_10592);
nand U11550 (N_11550,N_10850,N_10992);
or U11551 (N_11551,N_11178,N_10861);
and U11552 (N_11552,N_10726,N_10982);
nor U11553 (N_11553,N_11237,N_10905);
nor U11554 (N_11554,N_11208,N_10831);
and U11555 (N_11555,N_10934,N_11218);
and U11556 (N_11556,N_10941,N_10811);
and U11557 (N_11557,N_10779,N_10708);
and U11558 (N_11558,N_10989,N_10735);
nor U11559 (N_11559,N_10902,N_10917);
nand U11560 (N_11560,N_11084,N_10761);
and U11561 (N_11561,N_11029,N_11166);
nor U11562 (N_11562,N_10613,N_10513);
and U11563 (N_11563,N_11226,N_10709);
or U11564 (N_11564,N_10963,N_10643);
nand U11565 (N_11565,N_11065,N_10834);
or U11566 (N_11566,N_11231,N_11149);
nor U11567 (N_11567,N_11010,N_10827);
and U11568 (N_11568,N_11063,N_10886);
and U11569 (N_11569,N_10860,N_10645);
nand U11570 (N_11570,N_10832,N_10559);
or U11571 (N_11571,N_10508,N_10995);
nor U11572 (N_11572,N_10600,N_11019);
or U11573 (N_11573,N_10973,N_10626);
and U11574 (N_11574,N_10652,N_10540);
and U11575 (N_11575,N_10985,N_11167);
nand U11576 (N_11576,N_10997,N_11229);
xor U11577 (N_11577,N_10591,N_11194);
nand U11578 (N_11578,N_10523,N_10988);
nand U11579 (N_11579,N_10567,N_10728);
nand U11580 (N_11580,N_10703,N_11049);
xnor U11581 (N_11581,N_10847,N_10838);
and U11582 (N_11582,N_11030,N_11138);
nor U11583 (N_11583,N_10856,N_11073);
nand U11584 (N_11584,N_10598,N_10762);
nand U11585 (N_11585,N_10774,N_10606);
and U11586 (N_11586,N_10909,N_11129);
nand U11587 (N_11587,N_10677,N_10881);
or U11588 (N_11588,N_11126,N_11243);
nand U11589 (N_11589,N_11206,N_10519);
and U11590 (N_11590,N_11059,N_10919);
nor U11591 (N_11591,N_10546,N_11235);
or U11592 (N_11592,N_10845,N_11143);
nor U11593 (N_11593,N_10722,N_10694);
xnor U11594 (N_11594,N_10835,N_10549);
and U11595 (N_11595,N_11233,N_10851);
nor U11596 (N_11596,N_10545,N_10602);
nand U11597 (N_11597,N_11247,N_10839);
or U11598 (N_11598,N_10611,N_10906);
nor U11599 (N_11599,N_10715,N_10511);
or U11600 (N_11600,N_11223,N_11022);
nand U11601 (N_11601,N_10552,N_10589);
nand U11602 (N_11602,N_11168,N_10962);
and U11603 (N_11603,N_11004,N_10571);
nand U11604 (N_11604,N_10843,N_10685);
nand U11605 (N_11605,N_10622,N_10534);
xor U11606 (N_11606,N_11188,N_10822);
nor U11607 (N_11607,N_10943,N_11115);
and U11608 (N_11608,N_10732,N_11074);
nand U11609 (N_11609,N_10554,N_11151);
nor U11610 (N_11610,N_11162,N_10878);
and U11611 (N_11611,N_10607,N_11163);
nor U11612 (N_11612,N_10750,N_10867);
nand U11613 (N_11613,N_10764,N_11165);
nand U11614 (N_11614,N_11240,N_11217);
and U11615 (N_11615,N_10725,N_10672);
xnor U11616 (N_11616,N_11015,N_10849);
nand U11617 (N_11617,N_10539,N_10751);
nand U11618 (N_11618,N_10696,N_11000);
nand U11619 (N_11619,N_11011,N_11036);
nor U11620 (N_11620,N_11144,N_10563);
nand U11621 (N_11621,N_10931,N_11061);
or U11622 (N_11622,N_11207,N_10543);
and U11623 (N_11623,N_11042,N_11112);
and U11624 (N_11624,N_11185,N_10568);
and U11625 (N_11625,N_11159,N_10784);
nor U11626 (N_11626,N_10735,N_11131);
xnor U11627 (N_11627,N_10945,N_10939);
and U11628 (N_11628,N_10685,N_10943);
nor U11629 (N_11629,N_10907,N_10944);
and U11630 (N_11630,N_10848,N_10928);
and U11631 (N_11631,N_11009,N_10650);
nor U11632 (N_11632,N_10536,N_11171);
nor U11633 (N_11633,N_11045,N_10819);
nand U11634 (N_11634,N_10646,N_10662);
nor U11635 (N_11635,N_10707,N_10732);
and U11636 (N_11636,N_10749,N_11237);
nand U11637 (N_11637,N_10736,N_10511);
nor U11638 (N_11638,N_11016,N_10967);
nor U11639 (N_11639,N_10985,N_10988);
and U11640 (N_11640,N_10556,N_10529);
nor U11641 (N_11641,N_10657,N_11225);
or U11642 (N_11642,N_10949,N_10853);
or U11643 (N_11643,N_11022,N_10979);
and U11644 (N_11644,N_10548,N_10771);
nand U11645 (N_11645,N_10886,N_10504);
nand U11646 (N_11646,N_10592,N_10942);
xnor U11647 (N_11647,N_10577,N_10630);
and U11648 (N_11648,N_10614,N_10720);
nor U11649 (N_11649,N_10538,N_11121);
or U11650 (N_11650,N_10814,N_10950);
nor U11651 (N_11651,N_10924,N_10786);
nand U11652 (N_11652,N_11083,N_10555);
nor U11653 (N_11653,N_10549,N_10954);
nand U11654 (N_11654,N_10698,N_11160);
nor U11655 (N_11655,N_11183,N_10975);
nand U11656 (N_11656,N_10864,N_10853);
or U11657 (N_11657,N_10972,N_11196);
or U11658 (N_11658,N_10922,N_10813);
nor U11659 (N_11659,N_10928,N_10932);
nand U11660 (N_11660,N_10771,N_11092);
and U11661 (N_11661,N_10732,N_11223);
nand U11662 (N_11662,N_10660,N_10522);
nand U11663 (N_11663,N_10518,N_10589);
nor U11664 (N_11664,N_10882,N_10858);
nor U11665 (N_11665,N_11178,N_10737);
nand U11666 (N_11666,N_10671,N_11036);
nor U11667 (N_11667,N_10808,N_10815);
or U11668 (N_11668,N_10712,N_10984);
nor U11669 (N_11669,N_11170,N_10592);
xor U11670 (N_11670,N_11028,N_10746);
and U11671 (N_11671,N_11226,N_11061);
and U11672 (N_11672,N_10682,N_10566);
or U11673 (N_11673,N_11019,N_11129);
or U11674 (N_11674,N_10996,N_10823);
or U11675 (N_11675,N_10671,N_10688);
nand U11676 (N_11676,N_10799,N_11220);
nor U11677 (N_11677,N_10818,N_10681);
nand U11678 (N_11678,N_10573,N_10955);
or U11679 (N_11679,N_10996,N_10871);
nand U11680 (N_11680,N_10646,N_10538);
nor U11681 (N_11681,N_10947,N_11218);
nand U11682 (N_11682,N_10745,N_11213);
or U11683 (N_11683,N_10766,N_10624);
nand U11684 (N_11684,N_10863,N_10583);
nand U11685 (N_11685,N_10746,N_10722);
and U11686 (N_11686,N_10932,N_10739);
xor U11687 (N_11687,N_11060,N_10643);
nor U11688 (N_11688,N_11178,N_10643);
nand U11689 (N_11689,N_11243,N_11077);
xor U11690 (N_11690,N_10801,N_10514);
and U11691 (N_11691,N_10583,N_11053);
xnor U11692 (N_11692,N_10576,N_10547);
and U11693 (N_11693,N_11117,N_10895);
nand U11694 (N_11694,N_10830,N_10629);
nand U11695 (N_11695,N_10885,N_11025);
or U11696 (N_11696,N_10900,N_10646);
or U11697 (N_11697,N_10730,N_10989);
and U11698 (N_11698,N_11243,N_10623);
nor U11699 (N_11699,N_10602,N_10701);
nand U11700 (N_11700,N_10729,N_11182);
nand U11701 (N_11701,N_10829,N_10998);
xor U11702 (N_11702,N_10740,N_10903);
nor U11703 (N_11703,N_10609,N_11048);
nand U11704 (N_11704,N_10859,N_10907);
or U11705 (N_11705,N_11211,N_11065);
or U11706 (N_11706,N_10570,N_10798);
nor U11707 (N_11707,N_11094,N_11055);
or U11708 (N_11708,N_10802,N_11163);
or U11709 (N_11709,N_10582,N_10630);
and U11710 (N_11710,N_10786,N_11159);
and U11711 (N_11711,N_11014,N_10500);
nor U11712 (N_11712,N_10518,N_11183);
and U11713 (N_11713,N_10585,N_11031);
and U11714 (N_11714,N_11102,N_11104);
nor U11715 (N_11715,N_11145,N_10645);
and U11716 (N_11716,N_11069,N_11104);
or U11717 (N_11717,N_11110,N_11207);
nand U11718 (N_11718,N_11151,N_11103);
and U11719 (N_11719,N_10565,N_10872);
nand U11720 (N_11720,N_11035,N_11063);
and U11721 (N_11721,N_11156,N_10946);
nor U11722 (N_11722,N_11155,N_11242);
nand U11723 (N_11723,N_11030,N_10543);
nand U11724 (N_11724,N_10810,N_11136);
nand U11725 (N_11725,N_10558,N_10573);
xor U11726 (N_11726,N_10852,N_10836);
nand U11727 (N_11727,N_10723,N_11136);
and U11728 (N_11728,N_10639,N_10758);
and U11729 (N_11729,N_10997,N_10659);
nor U11730 (N_11730,N_10654,N_10772);
or U11731 (N_11731,N_11142,N_11225);
and U11732 (N_11732,N_11070,N_10854);
xnor U11733 (N_11733,N_11029,N_11168);
or U11734 (N_11734,N_10688,N_11025);
and U11735 (N_11735,N_10839,N_11037);
or U11736 (N_11736,N_10866,N_11055);
or U11737 (N_11737,N_10736,N_10545);
and U11738 (N_11738,N_11151,N_11079);
nand U11739 (N_11739,N_10662,N_10710);
and U11740 (N_11740,N_10621,N_10901);
xnor U11741 (N_11741,N_10839,N_10712);
or U11742 (N_11742,N_10590,N_10799);
xnor U11743 (N_11743,N_10598,N_11035);
and U11744 (N_11744,N_11183,N_11172);
and U11745 (N_11745,N_10955,N_10700);
xnor U11746 (N_11746,N_10558,N_11184);
nor U11747 (N_11747,N_11014,N_10520);
nand U11748 (N_11748,N_11222,N_10982);
nand U11749 (N_11749,N_11062,N_10787);
or U11750 (N_11750,N_11121,N_11135);
and U11751 (N_11751,N_10521,N_11001);
nand U11752 (N_11752,N_11172,N_10560);
or U11753 (N_11753,N_11236,N_11156);
and U11754 (N_11754,N_10817,N_11006);
nand U11755 (N_11755,N_11248,N_11079);
and U11756 (N_11756,N_10638,N_10972);
and U11757 (N_11757,N_10541,N_11083);
nand U11758 (N_11758,N_10993,N_11084);
nor U11759 (N_11759,N_11031,N_10708);
or U11760 (N_11760,N_10602,N_10790);
or U11761 (N_11761,N_10571,N_10820);
or U11762 (N_11762,N_11013,N_10776);
or U11763 (N_11763,N_11225,N_10549);
and U11764 (N_11764,N_11170,N_11075);
and U11765 (N_11765,N_11082,N_11118);
nor U11766 (N_11766,N_10880,N_10858);
and U11767 (N_11767,N_10698,N_10769);
and U11768 (N_11768,N_11102,N_11192);
and U11769 (N_11769,N_10511,N_10836);
nor U11770 (N_11770,N_10662,N_11125);
nor U11771 (N_11771,N_11205,N_10804);
or U11772 (N_11772,N_10596,N_10787);
nand U11773 (N_11773,N_11195,N_10627);
nand U11774 (N_11774,N_10655,N_10944);
nand U11775 (N_11775,N_11213,N_10797);
nand U11776 (N_11776,N_11011,N_11227);
or U11777 (N_11777,N_11139,N_10589);
xor U11778 (N_11778,N_10786,N_10705);
and U11779 (N_11779,N_10924,N_10925);
nand U11780 (N_11780,N_10885,N_11053);
and U11781 (N_11781,N_10839,N_10940);
xor U11782 (N_11782,N_10878,N_11189);
nor U11783 (N_11783,N_10755,N_11196);
nor U11784 (N_11784,N_10746,N_10602);
or U11785 (N_11785,N_10614,N_10719);
or U11786 (N_11786,N_10822,N_10800);
and U11787 (N_11787,N_11215,N_10865);
and U11788 (N_11788,N_10774,N_11125);
and U11789 (N_11789,N_10792,N_10691);
xor U11790 (N_11790,N_11247,N_10657);
nor U11791 (N_11791,N_10732,N_10812);
and U11792 (N_11792,N_10661,N_10968);
and U11793 (N_11793,N_11077,N_10911);
or U11794 (N_11794,N_11016,N_10914);
xor U11795 (N_11795,N_10746,N_10837);
and U11796 (N_11796,N_10555,N_10745);
or U11797 (N_11797,N_10748,N_11214);
nor U11798 (N_11798,N_11247,N_10943);
nand U11799 (N_11799,N_10875,N_11018);
and U11800 (N_11800,N_11177,N_10793);
and U11801 (N_11801,N_11110,N_10734);
nor U11802 (N_11802,N_10817,N_10504);
or U11803 (N_11803,N_10824,N_11115);
nor U11804 (N_11804,N_10736,N_11189);
xnor U11805 (N_11805,N_10512,N_10998);
nor U11806 (N_11806,N_10886,N_10953);
nand U11807 (N_11807,N_10717,N_10941);
xor U11808 (N_11808,N_11130,N_10618);
xnor U11809 (N_11809,N_10866,N_10635);
or U11810 (N_11810,N_11050,N_10821);
nand U11811 (N_11811,N_11229,N_10820);
or U11812 (N_11812,N_10760,N_10522);
nand U11813 (N_11813,N_10732,N_11110);
or U11814 (N_11814,N_10756,N_10938);
or U11815 (N_11815,N_10999,N_11058);
nand U11816 (N_11816,N_10718,N_10708);
and U11817 (N_11817,N_10893,N_10955);
nand U11818 (N_11818,N_10872,N_10931);
or U11819 (N_11819,N_10645,N_10794);
nor U11820 (N_11820,N_10798,N_11198);
nor U11821 (N_11821,N_10832,N_11001);
and U11822 (N_11822,N_10534,N_10712);
nand U11823 (N_11823,N_10521,N_10612);
or U11824 (N_11824,N_11179,N_10524);
and U11825 (N_11825,N_10812,N_10609);
and U11826 (N_11826,N_11075,N_10887);
nand U11827 (N_11827,N_10611,N_10840);
nor U11828 (N_11828,N_11002,N_11134);
and U11829 (N_11829,N_10912,N_10888);
nand U11830 (N_11830,N_10815,N_10519);
and U11831 (N_11831,N_10940,N_11095);
nor U11832 (N_11832,N_10598,N_10512);
nand U11833 (N_11833,N_11094,N_11186);
nand U11834 (N_11834,N_11200,N_11054);
and U11835 (N_11835,N_10844,N_10785);
xnor U11836 (N_11836,N_10522,N_10513);
or U11837 (N_11837,N_10804,N_10571);
and U11838 (N_11838,N_10628,N_10724);
nand U11839 (N_11839,N_10781,N_10610);
or U11840 (N_11840,N_10843,N_11167);
nor U11841 (N_11841,N_10764,N_10818);
xnor U11842 (N_11842,N_10646,N_10511);
nand U11843 (N_11843,N_10899,N_10662);
nor U11844 (N_11844,N_11187,N_11071);
and U11845 (N_11845,N_10958,N_10518);
nor U11846 (N_11846,N_10636,N_11037);
nor U11847 (N_11847,N_10826,N_11003);
nor U11848 (N_11848,N_11158,N_10597);
nor U11849 (N_11849,N_11075,N_11167);
or U11850 (N_11850,N_10612,N_10959);
and U11851 (N_11851,N_11123,N_10627);
nand U11852 (N_11852,N_10919,N_10678);
nor U11853 (N_11853,N_10800,N_11148);
nor U11854 (N_11854,N_10983,N_10922);
nor U11855 (N_11855,N_10867,N_10516);
xor U11856 (N_11856,N_10787,N_10501);
nor U11857 (N_11857,N_11228,N_10963);
nand U11858 (N_11858,N_10893,N_10675);
or U11859 (N_11859,N_10785,N_10829);
xor U11860 (N_11860,N_10667,N_10715);
nor U11861 (N_11861,N_10885,N_10616);
nor U11862 (N_11862,N_11058,N_10625);
xor U11863 (N_11863,N_11096,N_10802);
nor U11864 (N_11864,N_10830,N_10622);
nor U11865 (N_11865,N_10843,N_11040);
nor U11866 (N_11866,N_11124,N_10603);
nor U11867 (N_11867,N_10929,N_10554);
nor U11868 (N_11868,N_10978,N_10952);
or U11869 (N_11869,N_10873,N_10823);
or U11870 (N_11870,N_10999,N_11168);
and U11871 (N_11871,N_11081,N_10687);
and U11872 (N_11872,N_11052,N_10878);
or U11873 (N_11873,N_10640,N_11196);
nand U11874 (N_11874,N_10978,N_11200);
and U11875 (N_11875,N_10793,N_10759);
and U11876 (N_11876,N_10712,N_10701);
or U11877 (N_11877,N_10924,N_10519);
nand U11878 (N_11878,N_10668,N_10790);
or U11879 (N_11879,N_10632,N_11050);
or U11880 (N_11880,N_11032,N_10850);
nor U11881 (N_11881,N_11112,N_11234);
nand U11882 (N_11882,N_10987,N_11181);
and U11883 (N_11883,N_10625,N_10715);
nor U11884 (N_11884,N_10882,N_10848);
xnor U11885 (N_11885,N_10862,N_10713);
and U11886 (N_11886,N_10635,N_10964);
or U11887 (N_11887,N_10808,N_10575);
nand U11888 (N_11888,N_11171,N_10569);
nand U11889 (N_11889,N_10999,N_10738);
or U11890 (N_11890,N_10622,N_11174);
or U11891 (N_11891,N_10686,N_11046);
nor U11892 (N_11892,N_10767,N_10955);
xor U11893 (N_11893,N_11105,N_10661);
nand U11894 (N_11894,N_10573,N_10700);
and U11895 (N_11895,N_10901,N_11083);
nand U11896 (N_11896,N_11181,N_10631);
or U11897 (N_11897,N_11178,N_10841);
and U11898 (N_11898,N_10810,N_11221);
xnor U11899 (N_11899,N_11244,N_10599);
nand U11900 (N_11900,N_11042,N_11204);
nand U11901 (N_11901,N_11177,N_11163);
or U11902 (N_11902,N_11196,N_10696);
and U11903 (N_11903,N_11086,N_10882);
or U11904 (N_11904,N_11212,N_10966);
or U11905 (N_11905,N_11202,N_10695);
nand U11906 (N_11906,N_10842,N_10755);
nor U11907 (N_11907,N_10518,N_10900);
and U11908 (N_11908,N_11204,N_10771);
or U11909 (N_11909,N_10672,N_10616);
nand U11910 (N_11910,N_11023,N_10599);
xnor U11911 (N_11911,N_10800,N_10734);
xor U11912 (N_11912,N_10992,N_10931);
or U11913 (N_11913,N_10516,N_10535);
nand U11914 (N_11914,N_11230,N_10702);
nand U11915 (N_11915,N_10624,N_10600);
or U11916 (N_11916,N_10790,N_10811);
and U11917 (N_11917,N_10676,N_10672);
nand U11918 (N_11918,N_10618,N_10898);
or U11919 (N_11919,N_10707,N_11191);
xor U11920 (N_11920,N_10560,N_10758);
xnor U11921 (N_11921,N_11139,N_10936);
or U11922 (N_11922,N_10607,N_11179);
nor U11923 (N_11923,N_10517,N_11189);
nor U11924 (N_11924,N_10623,N_10995);
and U11925 (N_11925,N_11117,N_10981);
and U11926 (N_11926,N_10796,N_11248);
nor U11927 (N_11927,N_10853,N_11067);
nor U11928 (N_11928,N_10889,N_10775);
nor U11929 (N_11929,N_10692,N_10815);
and U11930 (N_11930,N_11114,N_11172);
or U11931 (N_11931,N_10981,N_11114);
or U11932 (N_11932,N_11040,N_10650);
nor U11933 (N_11933,N_11229,N_11080);
and U11934 (N_11934,N_10987,N_11212);
or U11935 (N_11935,N_10776,N_10854);
or U11936 (N_11936,N_10997,N_10812);
or U11937 (N_11937,N_10836,N_10983);
or U11938 (N_11938,N_11186,N_10983);
xnor U11939 (N_11939,N_11142,N_10972);
nand U11940 (N_11940,N_11079,N_11116);
and U11941 (N_11941,N_10639,N_11054);
xor U11942 (N_11942,N_10943,N_10636);
or U11943 (N_11943,N_11202,N_10955);
nand U11944 (N_11944,N_11136,N_11119);
and U11945 (N_11945,N_10600,N_10900);
nand U11946 (N_11946,N_10699,N_10716);
nand U11947 (N_11947,N_11245,N_10570);
nor U11948 (N_11948,N_10795,N_10863);
or U11949 (N_11949,N_10537,N_10705);
nand U11950 (N_11950,N_11212,N_11128);
nor U11951 (N_11951,N_11055,N_11130);
nand U11952 (N_11952,N_11009,N_10800);
nand U11953 (N_11953,N_11110,N_10874);
and U11954 (N_11954,N_11195,N_10948);
nor U11955 (N_11955,N_10818,N_10518);
xnor U11956 (N_11956,N_10639,N_11051);
xor U11957 (N_11957,N_10766,N_10912);
or U11958 (N_11958,N_10733,N_11125);
nor U11959 (N_11959,N_10837,N_10547);
or U11960 (N_11960,N_11114,N_10674);
and U11961 (N_11961,N_11181,N_10584);
and U11962 (N_11962,N_10552,N_11186);
nor U11963 (N_11963,N_10644,N_10605);
nand U11964 (N_11964,N_11024,N_10638);
and U11965 (N_11965,N_10951,N_11098);
nor U11966 (N_11966,N_11052,N_11209);
and U11967 (N_11967,N_11198,N_10504);
xnor U11968 (N_11968,N_10517,N_11169);
nand U11969 (N_11969,N_10951,N_10555);
nand U11970 (N_11970,N_10513,N_10710);
nand U11971 (N_11971,N_11137,N_10577);
nand U11972 (N_11972,N_10818,N_10896);
nand U11973 (N_11973,N_10981,N_11037);
and U11974 (N_11974,N_11074,N_10979);
and U11975 (N_11975,N_10626,N_10833);
and U11976 (N_11976,N_10976,N_10548);
nand U11977 (N_11977,N_10836,N_10755);
and U11978 (N_11978,N_10771,N_10675);
nand U11979 (N_11979,N_11028,N_11036);
nand U11980 (N_11980,N_10896,N_10723);
and U11981 (N_11981,N_10895,N_10890);
or U11982 (N_11982,N_11124,N_10993);
and U11983 (N_11983,N_10893,N_10521);
and U11984 (N_11984,N_11103,N_10783);
xnor U11985 (N_11985,N_11079,N_11118);
and U11986 (N_11986,N_10865,N_11086);
nand U11987 (N_11987,N_10529,N_11193);
and U11988 (N_11988,N_10546,N_10991);
nor U11989 (N_11989,N_11078,N_10724);
xor U11990 (N_11990,N_11099,N_10658);
and U11991 (N_11991,N_11248,N_10988);
and U11992 (N_11992,N_11184,N_10727);
or U11993 (N_11993,N_10954,N_10703);
nor U11994 (N_11994,N_11022,N_10995);
or U11995 (N_11995,N_10507,N_10927);
nand U11996 (N_11996,N_11054,N_10866);
or U11997 (N_11997,N_10852,N_10510);
nor U11998 (N_11998,N_10672,N_10881);
xnor U11999 (N_11999,N_11150,N_10603);
nand U12000 (N_12000,N_11256,N_11262);
nand U12001 (N_12001,N_11670,N_11924);
nor U12002 (N_12002,N_11523,N_11749);
xor U12003 (N_12003,N_11475,N_11326);
or U12004 (N_12004,N_11503,N_11562);
and U12005 (N_12005,N_11261,N_11297);
nand U12006 (N_12006,N_11993,N_11458);
and U12007 (N_12007,N_11837,N_11449);
or U12008 (N_12008,N_11917,N_11799);
and U12009 (N_12009,N_11428,N_11581);
nand U12010 (N_12010,N_11396,N_11653);
and U12011 (N_12011,N_11448,N_11401);
nor U12012 (N_12012,N_11651,N_11622);
or U12013 (N_12013,N_11641,N_11520);
xnor U12014 (N_12014,N_11443,N_11934);
nand U12015 (N_12015,N_11388,N_11666);
or U12016 (N_12016,N_11358,N_11915);
or U12017 (N_12017,N_11509,N_11865);
and U12018 (N_12018,N_11943,N_11422);
nand U12019 (N_12019,N_11854,N_11790);
nand U12020 (N_12020,N_11892,N_11834);
and U12021 (N_12021,N_11384,N_11619);
nand U12022 (N_12022,N_11379,N_11411);
or U12023 (N_12023,N_11480,N_11997);
or U12024 (N_12024,N_11374,N_11766);
and U12025 (N_12025,N_11404,N_11894);
or U12026 (N_12026,N_11492,N_11642);
and U12027 (N_12027,N_11360,N_11484);
and U12028 (N_12028,N_11822,N_11727);
nor U12029 (N_12029,N_11890,N_11946);
nand U12030 (N_12030,N_11494,N_11335);
nor U12031 (N_12031,N_11489,N_11561);
or U12032 (N_12032,N_11763,N_11381);
and U12033 (N_12033,N_11913,N_11788);
or U12034 (N_12034,N_11330,N_11873);
nand U12035 (N_12035,N_11795,N_11327);
nand U12036 (N_12036,N_11811,N_11539);
nor U12037 (N_12037,N_11307,N_11944);
and U12038 (N_12038,N_11424,N_11988);
nand U12039 (N_12039,N_11293,N_11706);
or U12040 (N_12040,N_11688,N_11356);
nor U12041 (N_12041,N_11765,N_11252);
nand U12042 (N_12042,N_11856,N_11710);
nor U12043 (N_12043,N_11703,N_11536);
nor U12044 (N_12044,N_11729,N_11732);
nor U12045 (N_12045,N_11349,N_11544);
nor U12046 (N_12046,N_11957,N_11800);
nor U12047 (N_12047,N_11324,N_11276);
nand U12048 (N_12048,N_11928,N_11620);
nor U12049 (N_12049,N_11310,N_11580);
and U12050 (N_12050,N_11578,N_11771);
or U12051 (N_12051,N_11624,N_11987);
or U12052 (N_12052,N_11785,N_11901);
and U12053 (N_12053,N_11724,N_11332);
or U12054 (N_12054,N_11515,N_11251);
or U12055 (N_12055,N_11806,N_11504);
nor U12056 (N_12056,N_11370,N_11627);
nand U12057 (N_12057,N_11826,N_11468);
nor U12058 (N_12058,N_11419,N_11522);
or U12059 (N_12059,N_11886,N_11889);
nand U12060 (N_12060,N_11745,N_11643);
nand U12061 (N_12061,N_11345,N_11664);
and U12062 (N_12062,N_11748,N_11958);
nor U12063 (N_12063,N_11417,N_11258);
nor U12064 (N_12064,N_11777,N_11275);
nand U12065 (N_12065,N_11658,N_11339);
nand U12066 (N_12066,N_11851,N_11630);
nor U12067 (N_12067,N_11833,N_11662);
or U12068 (N_12068,N_11780,N_11585);
and U12069 (N_12069,N_11798,N_11714);
or U12070 (N_12070,N_11552,N_11968);
nand U12071 (N_12071,N_11316,N_11413);
nand U12072 (N_12072,N_11974,N_11859);
nor U12073 (N_12073,N_11451,N_11789);
or U12074 (N_12074,N_11648,N_11699);
nand U12075 (N_12075,N_11996,N_11399);
xnor U12076 (N_12076,N_11902,N_11885);
or U12077 (N_12077,N_11555,N_11493);
xor U12078 (N_12078,N_11830,N_11803);
and U12079 (N_12079,N_11908,N_11846);
xnor U12080 (N_12080,N_11808,N_11738);
nor U12081 (N_12081,N_11589,N_11464);
and U12082 (N_12082,N_11511,N_11352);
nand U12083 (N_12083,N_11867,N_11774);
nor U12084 (N_12084,N_11739,N_11270);
or U12085 (N_12085,N_11740,N_11977);
nor U12086 (N_12086,N_11866,N_11966);
nand U12087 (N_12087,N_11880,N_11827);
nor U12088 (N_12088,N_11805,N_11418);
nand U12089 (N_12089,N_11440,N_11392);
nor U12090 (N_12090,N_11538,N_11435);
or U12091 (N_12091,N_11845,N_11758);
nor U12092 (N_12092,N_11632,N_11962);
or U12093 (N_12093,N_11274,N_11896);
nand U12094 (N_12094,N_11753,N_11817);
or U12095 (N_12095,N_11454,N_11259);
nand U12096 (N_12096,N_11593,N_11558);
or U12097 (N_12097,N_11663,N_11487);
nor U12098 (N_12098,N_11576,N_11537);
and U12099 (N_12099,N_11628,N_11441);
or U12100 (N_12100,N_11855,N_11989);
nand U12101 (N_12101,N_11991,N_11704);
xor U12102 (N_12102,N_11255,N_11891);
and U12103 (N_12103,N_11807,N_11495);
nand U12104 (N_12104,N_11960,N_11718);
nand U12105 (N_12105,N_11410,N_11400);
and U12106 (N_12106,N_11540,N_11810);
nand U12107 (N_12107,N_11969,N_11707);
and U12108 (N_12108,N_11348,N_11265);
nor U12109 (N_12109,N_11906,N_11457);
nand U12110 (N_12110,N_11271,N_11661);
and U12111 (N_12111,N_11814,N_11868);
or U12112 (N_12112,N_11331,N_11336);
xor U12113 (N_12113,N_11932,N_11722);
nand U12114 (N_12114,N_11687,N_11847);
nor U12115 (N_12115,N_11741,N_11883);
nand U12116 (N_12116,N_11824,N_11306);
nand U12117 (N_12117,N_11382,N_11542);
nand U12118 (N_12118,N_11927,N_11362);
nor U12119 (N_12119,N_11416,N_11998);
xnor U12120 (N_12120,N_11541,N_11647);
or U12121 (N_12121,N_11559,N_11754);
or U12122 (N_12122,N_11782,N_11858);
or U12123 (N_12123,N_11947,N_11922);
nor U12124 (N_12124,N_11796,N_11264);
and U12125 (N_12125,N_11923,N_11668);
or U12126 (N_12126,N_11629,N_11994);
and U12127 (N_12127,N_11534,N_11823);
and U12128 (N_12128,N_11900,N_11446);
nor U12129 (N_12129,N_11528,N_11587);
nand U12130 (N_12130,N_11412,N_11967);
and U12131 (N_12131,N_11592,N_11321);
and U12132 (N_12132,N_11529,N_11548);
and U12133 (N_12133,N_11965,N_11978);
or U12134 (N_12134,N_11683,N_11471);
nor U12135 (N_12135,N_11533,N_11547);
and U12136 (N_12136,N_11402,N_11756);
nand U12137 (N_12137,N_11616,N_11819);
and U12138 (N_12138,N_11999,N_11870);
nand U12139 (N_12139,N_11301,N_11941);
nor U12140 (N_12140,N_11831,N_11575);
nor U12141 (N_12141,N_11359,N_11848);
nand U12142 (N_12142,N_11801,N_11617);
and U12143 (N_12143,N_11346,N_11496);
nand U12144 (N_12144,N_11815,N_11295);
nand U12145 (N_12145,N_11672,N_11570);
or U12146 (N_12146,N_11595,N_11689);
nand U12147 (N_12147,N_11383,N_11611);
nor U12148 (N_12148,N_11925,N_11787);
nor U12149 (N_12149,N_11296,N_11692);
or U12150 (N_12150,N_11828,N_11566);
nand U12151 (N_12151,N_11311,N_11737);
and U12152 (N_12152,N_11884,N_11604);
nand U12153 (N_12153,N_11899,N_11260);
nor U12154 (N_12154,N_11843,N_11577);
and U12155 (N_12155,N_11931,N_11371);
or U12156 (N_12156,N_11476,N_11638);
and U12157 (N_12157,N_11726,N_11283);
or U12158 (N_12158,N_11304,N_11567);
or U12159 (N_12159,N_11733,N_11744);
nand U12160 (N_12160,N_11527,N_11409);
nand U12161 (N_12161,N_11463,N_11612);
and U12162 (N_12162,N_11660,N_11677);
and U12163 (N_12163,N_11635,N_11711);
or U12164 (N_12164,N_11693,N_11488);
nor U12165 (N_12165,N_11450,N_11333);
or U12166 (N_12166,N_11709,N_11277);
and U12167 (N_12167,N_11818,N_11361);
and U12168 (N_12168,N_11905,N_11783);
nand U12169 (N_12169,N_11775,N_11387);
or U12170 (N_12170,N_11602,N_11621);
and U12171 (N_12171,N_11586,N_11747);
or U12172 (N_12172,N_11970,N_11505);
xnor U12173 (N_12173,N_11861,N_11469);
and U12174 (N_12174,N_11712,N_11961);
nor U12175 (N_12175,N_11702,N_11369);
or U12176 (N_12176,N_11483,N_11742);
or U12177 (N_12177,N_11445,N_11626);
nand U12178 (N_12178,N_11420,N_11809);
or U12179 (N_12179,N_11600,N_11973);
or U12180 (N_12180,N_11608,N_11317);
or U12181 (N_12181,N_11948,N_11355);
or U12182 (N_12182,N_11376,N_11279);
and U12183 (N_12183,N_11940,N_11564);
xor U12184 (N_12184,N_11303,N_11736);
or U12185 (N_12185,N_11408,N_11531);
and U12186 (N_12186,N_11907,N_11514);
or U12187 (N_12187,N_11954,N_11474);
and U12188 (N_12188,N_11287,N_11601);
nand U12189 (N_12189,N_11414,N_11588);
nand U12190 (N_12190,N_11983,N_11305);
nand U12191 (N_12191,N_11556,N_11308);
nand U12192 (N_12192,N_11390,N_11452);
nor U12193 (N_12193,N_11486,N_11583);
nor U12194 (N_12194,N_11779,N_11300);
or U12195 (N_12195,N_11521,N_11984);
and U12196 (N_12196,N_11263,N_11502);
and U12197 (N_12197,N_11309,N_11568);
nor U12198 (N_12198,N_11746,N_11398);
nor U12199 (N_12199,N_11266,N_11813);
or U12200 (N_12200,N_11357,N_11980);
nor U12201 (N_12201,N_11553,N_11656);
or U12202 (N_12202,N_11426,N_11910);
and U12203 (N_12203,N_11453,N_11281);
or U12204 (N_12204,N_11519,N_11462);
and U12205 (N_12205,N_11708,N_11278);
or U12206 (N_12206,N_11770,N_11875);
or U12207 (N_12207,N_11344,N_11691);
nand U12208 (N_12208,N_11513,N_11280);
or U12209 (N_12209,N_11425,N_11772);
nor U12210 (N_12210,N_11778,N_11955);
and U12211 (N_12211,N_11431,N_11935);
nor U12212 (N_12212,N_11895,N_11294);
nand U12213 (N_12213,N_11298,N_11904);
and U12214 (N_12214,N_11872,N_11951);
nor U12215 (N_12215,N_11760,N_11761);
or U12216 (N_12216,N_11609,N_11535);
nor U12217 (N_12217,N_11341,N_11717);
and U12218 (N_12218,N_11517,N_11860);
or U12219 (N_12219,N_11715,N_11821);
nor U12220 (N_12220,N_11322,N_11914);
nand U12221 (N_12221,N_11794,N_11490);
nor U12222 (N_12222,N_11597,N_11734);
nand U12223 (N_12223,N_11942,N_11518);
nor U12224 (N_12224,N_11838,N_11606);
nor U12225 (N_12225,N_11500,N_11871);
nand U12226 (N_12226,N_11288,N_11945);
or U12227 (N_12227,N_11700,N_11912);
or U12228 (N_12228,N_11675,N_11716);
and U12229 (N_12229,N_11603,N_11459);
or U12230 (N_12230,N_11897,N_11764);
or U12231 (N_12231,N_11719,N_11992);
or U12232 (N_12232,N_11768,N_11743);
nand U12233 (N_12233,N_11524,N_11353);
nand U12234 (N_12234,N_11644,N_11573);
nor U12235 (N_12235,N_11507,N_11841);
xor U12236 (N_12236,N_11427,N_11781);
and U12237 (N_12237,N_11437,N_11645);
nand U12238 (N_12238,N_11366,N_11497);
nand U12239 (N_12239,N_11921,N_11659);
and U12240 (N_12240,N_11466,N_11313);
nor U12241 (N_12241,N_11268,N_11721);
nor U12242 (N_12242,N_11590,N_11351);
nand U12243 (N_12243,N_11930,N_11730);
or U12244 (N_12244,N_11257,N_11607);
nand U12245 (N_12245,N_11926,N_11793);
nor U12246 (N_12246,N_11972,N_11543);
xor U12247 (N_12247,N_11920,N_11421);
nor U12248 (N_12248,N_11574,N_11325);
or U12249 (N_12249,N_11887,N_11472);
and U12250 (N_12250,N_11516,N_11591);
nor U12251 (N_12251,N_11916,N_11731);
or U12252 (N_12252,N_11852,N_11698);
nor U12253 (N_12253,N_11423,N_11334);
and U12254 (N_12254,N_11874,N_11684);
nor U12255 (N_12255,N_11671,N_11757);
or U12256 (N_12256,N_11415,N_11338);
nand U12257 (N_12257,N_11579,N_11499);
nor U12258 (N_12258,N_11784,N_11665);
nor U12259 (N_12259,N_11532,N_11498);
or U12260 (N_12260,N_11669,N_11836);
nand U12261 (N_12261,N_11640,N_11971);
or U12262 (N_12262,N_11269,N_11705);
nand U12263 (N_12263,N_11939,N_11876);
nand U12264 (N_12264,N_11995,N_11862);
and U12265 (N_12265,N_11981,N_11986);
xnor U12266 (N_12266,N_11582,N_11444);
or U12267 (N_12267,N_11956,N_11633);
xor U12268 (N_12268,N_11302,N_11596);
nor U12269 (N_12269,N_11485,N_11755);
nand U12270 (N_12270,N_11686,N_11888);
nand U12271 (N_12271,N_11253,N_11864);
nand U12272 (N_12272,N_11657,N_11695);
nor U12273 (N_12273,N_11364,N_11639);
xnor U12274 (N_12274,N_11403,N_11701);
xnor U12275 (N_12275,N_11812,N_11312);
or U12276 (N_12276,N_11685,N_11508);
nand U12277 (N_12277,N_11501,N_11563);
nand U12278 (N_12278,N_11386,N_11975);
or U12279 (N_12279,N_11918,N_11636);
nor U12280 (N_12280,N_11328,N_11337);
nand U12281 (N_12281,N_11898,N_11530);
and U12282 (N_12282,N_11769,N_11365);
xor U12283 (N_12283,N_11882,N_11526);
or U12284 (N_12284,N_11938,N_11985);
and U12285 (N_12285,N_11982,N_11825);
or U12286 (N_12286,N_11525,N_11751);
and U12287 (N_12287,N_11797,N_11546);
nand U12288 (N_12288,N_11272,N_11844);
and U12289 (N_12289,N_11456,N_11903);
nor U12290 (N_12290,N_11491,N_11373);
and U12291 (N_12291,N_11694,N_11990);
nand U12292 (N_12292,N_11850,N_11682);
nor U12293 (N_12293,N_11649,N_11853);
nor U12294 (N_12294,N_11510,N_11438);
and U12295 (N_12295,N_11678,N_11479);
or U12296 (N_12296,N_11584,N_11477);
and U12297 (N_12297,N_11342,N_11953);
nand U12298 (N_12298,N_11637,N_11460);
and U12299 (N_12299,N_11285,N_11447);
nand U12300 (N_12300,N_11439,N_11832);
nor U12301 (N_12301,N_11565,N_11389);
or U12302 (N_12302,N_11470,N_11461);
and U12303 (N_12303,N_11613,N_11594);
nor U12304 (N_12304,N_11433,N_11676);
nor U12305 (N_12305,N_11720,N_11929);
or U12306 (N_12306,N_11634,N_11654);
and U12307 (N_12307,N_11254,N_11250);
or U12308 (N_12308,N_11842,N_11963);
nand U12309 (N_12309,N_11723,N_11347);
xor U12310 (N_12310,N_11372,N_11323);
nand U12311 (N_12311,N_11354,N_11292);
nand U12312 (N_12312,N_11393,N_11482);
xor U12313 (N_12313,N_11652,N_11395);
nor U12314 (N_12314,N_11933,N_11318);
nor U12315 (N_12315,N_11314,N_11877);
nor U12316 (N_12316,N_11377,N_11599);
or U12317 (N_12317,N_11697,N_11735);
nor U12318 (N_12318,N_11713,N_11911);
nor U12319 (N_12319,N_11467,N_11950);
nand U12320 (N_12320,N_11976,N_11610);
nor U12321 (N_12321,N_11407,N_11598);
and U12322 (N_12322,N_11350,N_11397);
or U12323 (N_12323,N_11367,N_11340);
nor U12324 (N_12324,N_11979,N_11655);
nor U12325 (N_12325,N_11762,N_11290);
or U12326 (N_12326,N_11455,N_11319);
nand U12327 (N_12327,N_11646,N_11478);
or U12328 (N_12328,N_11863,N_11696);
nor U12329 (N_12329,N_11273,N_11792);
and U12330 (N_12330,N_11674,N_11571);
nand U12331 (N_12331,N_11752,N_11681);
and U12332 (N_12332,N_11430,N_11909);
nand U12333 (N_12333,N_11442,N_11791);
nor U12334 (N_12334,N_11820,N_11949);
and U12335 (N_12335,N_11569,N_11767);
and U12336 (N_12336,N_11572,N_11405);
nor U12337 (N_12337,N_11385,N_11465);
or U12338 (N_12338,N_11614,N_11728);
or U12339 (N_12339,N_11759,N_11690);
and U12340 (N_12340,N_11786,N_11299);
and U12341 (N_12341,N_11406,N_11673);
or U12342 (N_12342,N_11879,N_11554);
or U12343 (N_12343,N_11429,N_11919);
nor U12344 (N_12344,N_11380,N_11804);
nor U12345 (N_12345,N_11631,N_11802);
nor U12346 (N_12346,N_11329,N_11835);
nor U12347 (N_12347,N_11605,N_11680);
nor U12348 (N_12348,N_11506,N_11291);
nor U12349 (N_12349,N_11849,N_11282);
nor U12350 (N_12350,N_11964,N_11625);
nor U12351 (N_12351,N_11667,N_11952);
nand U12352 (N_12352,N_11375,N_11679);
nand U12353 (N_12353,N_11551,N_11394);
and U12354 (N_12354,N_11857,N_11869);
and U12355 (N_12355,N_11839,N_11615);
nor U12356 (N_12356,N_11473,N_11436);
nand U12357 (N_12357,N_11286,N_11560);
or U12358 (N_12358,N_11550,N_11937);
or U12359 (N_12359,N_11267,N_11289);
or U12360 (N_12360,N_11512,N_11893);
nor U12361 (N_12361,N_11363,N_11650);
or U12362 (N_12362,N_11725,N_11959);
and U12363 (N_12363,N_11284,N_11881);
or U12364 (N_12364,N_11391,N_11816);
or U12365 (N_12365,N_11545,N_11378);
and U12366 (N_12366,N_11776,N_11829);
or U12367 (N_12367,N_11773,N_11343);
and U12368 (N_12368,N_11315,N_11623);
or U12369 (N_12369,N_11549,N_11840);
or U12370 (N_12370,N_11368,N_11320);
or U12371 (N_12371,N_11481,N_11557);
or U12372 (N_12372,N_11618,N_11750);
nor U12373 (N_12373,N_11936,N_11878);
nor U12374 (N_12374,N_11432,N_11434);
or U12375 (N_12375,N_11487,N_11711);
or U12376 (N_12376,N_11706,N_11492);
nand U12377 (N_12377,N_11829,N_11760);
nand U12378 (N_12378,N_11842,N_11380);
and U12379 (N_12379,N_11465,N_11555);
and U12380 (N_12380,N_11864,N_11260);
xnor U12381 (N_12381,N_11286,N_11550);
nor U12382 (N_12382,N_11534,N_11377);
or U12383 (N_12383,N_11488,N_11309);
nor U12384 (N_12384,N_11695,N_11988);
and U12385 (N_12385,N_11473,N_11458);
and U12386 (N_12386,N_11522,N_11278);
or U12387 (N_12387,N_11598,N_11375);
nand U12388 (N_12388,N_11542,N_11358);
nor U12389 (N_12389,N_11367,N_11787);
or U12390 (N_12390,N_11547,N_11796);
and U12391 (N_12391,N_11914,N_11704);
nor U12392 (N_12392,N_11296,N_11998);
nor U12393 (N_12393,N_11288,N_11737);
nand U12394 (N_12394,N_11533,N_11646);
nor U12395 (N_12395,N_11384,N_11365);
and U12396 (N_12396,N_11970,N_11723);
xor U12397 (N_12397,N_11286,N_11754);
nor U12398 (N_12398,N_11893,N_11399);
xor U12399 (N_12399,N_11389,N_11269);
nor U12400 (N_12400,N_11280,N_11746);
nor U12401 (N_12401,N_11526,N_11670);
and U12402 (N_12402,N_11441,N_11501);
nor U12403 (N_12403,N_11322,N_11552);
or U12404 (N_12404,N_11921,N_11924);
or U12405 (N_12405,N_11893,N_11462);
and U12406 (N_12406,N_11260,N_11832);
and U12407 (N_12407,N_11596,N_11945);
nand U12408 (N_12408,N_11642,N_11980);
and U12409 (N_12409,N_11795,N_11620);
nor U12410 (N_12410,N_11537,N_11413);
nand U12411 (N_12411,N_11755,N_11370);
xor U12412 (N_12412,N_11353,N_11962);
and U12413 (N_12413,N_11458,N_11843);
or U12414 (N_12414,N_11419,N_11815);
nor U12415 (N_12415,N_11445,N_11942);
and U12416 (N_12416,N_11278,N_11613);
nand U12417 (N_12417,N_11621,N_11834);
nor U12418 (N_12418,N_11631,N_11572);
and U12419 (N_12419,N_11467,N_11378);
nand U12420 (N_12420,N_11600,N_11873);
nor U12421 (N_12421,N_11335,N_11513);
xor U12422 (N_12422,N_11920,N_11562);
nor U12423 (N_12423,N_11266,N_11697);
and U12424 (N_12424,N_11669,N_11823);
nor U12425 (N_12425,N_11561,N_11894);
nor U12426 (N_12426,N_11590,N_11960);
nor U12427 (N_12427,N_11854,N_11986);
nand U12428 (N_12428,N_11784,N_11592);
nand U12429 (N_12429,N_11677,N_11926);
nand U12430 (N_12430,N_11728,N_11973);
and U12431 (N_12431,N_11340,N_11437);
nand U12432 (N_12432,N_11469,N_11634);
xor U12433 (N_12433,N_11639,N_11308);
and U12434 (N_12434,N_11261,N_11412);
and U12435 (N_12435,N_11410,N_11986);
or U12436 (N_12436,N_11647,N_11674);
nand U12437 (N_12437,N_11792,N_11937);
nor U12438 (N_12438,N_11644,N_11328);
and U12439 (N_12439,N_11918,N_11789);
and U12440 (N_12440,N_11353,N_11489);
or U12441 (N_12441,N_11893,N_11911);
nor U12442 (N_12442,N_11941,N_11450);
and U12443 (N_12443,N_11482,N_11676);
or U12444 (N_12444,N_11567,N_11826);
and U12445 (N_12445,N_11835,N_11998);
or U12446 (N_12446,N_11983,N_11380);
nand U12447 (N_12447,N_11625,N_11408);
nand U12448 (N_12448,N_11612,N_11768);
nand U12449 (N_12449,N_11493,N_11399);
and U12450 (N_12450,N_11426,N_11796);
xnor U12451 (N_12451,N_11552,N_11960);
and U12452 (N_12452,N_11434,N_11374);
nand U12453 (N_12453,N_11435,N_11937);
and U12454 (N_12454,N_11375,N_11861);
nor U12455 (N_12455,N_11661,N_11495);
and U12456 (N_12456,N_11935,N_11765);
nand U12457 (N_12457,N_11392,N_11669);
nand U12458 (N_12458,N_11396,N_11545);
or U12459 (N_12459,N_11415,N_11552);
and U12460 (N_12460,N_11539,N_11932);
nand U12461 (N_12461,N_11342,N_11769);
or U12462 (N_12462,N_11741,N_11570);
or U12463 (N_12463,N_11555,N_11972);
nand U12464 (N_12464,N_11395,N_11573);
or U12465 (N_12465,N_11377,N_11949);
nor U12466 (N_12466,N_11449,N_11783);
and U12467 (N_12467,N_11926,N_11610);
or U12468 (N_12468,N_11703,N_11689);
and U12469 (N_12469,N_11337,N_11282);
nand U12470 (N_12470,N_11484,N_11411);
nor U12471 (N_12471,N_11552,N_11634);
or U12472 (N_12472,N_11447,N_11291);
or U12473 (N_12473,N_11276,N_11666);
nor U12474 (N_12474,N_11535,N_11468);
nor U12475 (N_12475,N_11590,N_11933);
nor U12476 (N_12476,N_11304,N_11637);
nand U12477 (N_12477,N_11634,N_11477);
and U12478 (N_12478,N_11588,N_11792);
or U12479 (N_12479,N_11856,N_11694);
nor U12480 (N_12480,N_11318,N_11361);
xor U12481 (N_12481,N_11412,N_11820);
or U12482 (N_12482,N_11467,N_11644);
nor U12483 (N_12483,N_11459,N_11306);
and U12484 (N_12484,N_11782,N_11627);
and U12485 (N_12485,N_11397,N_11336);
or U12486 (N_12486,N_11995,N_11551);
and U12487 (N_12487,N_11511,N_11775);
nor U12488 (N_12488,N_11470,N_11284);
nor U12489 (N_12489,N_11552,N_11444);
nor U12490 (N_12490,N_11727,N_11816);
and U12491 (N_12491,N_11818,N_11794);
nor U12492 (N_12492,N_11526,N_11483);
and U12493 (N_12493,N_11803,N_11387);
nor U12494 (N_12494,N_11581,N_11845);
nand U12495 (N_12495,N_11425,N_11919);
xnor U12496 (N_12496,N_11583,N_11386);
nand U12497 (N_12497,N_11385,N_11660);
xnor U12498 (N_12498,N_11599,N_11806);
nand U12499 (N_12499,N_11464,N_11697);
nor U12500 (N_12500,N_11622,N_11809);
and U12501 (N_12501,N_11676,N_11880);
nand U12502 (N_12502,N_11924,N_11909);
nand U12503 (N_12503,N_11530,N_11801);
or U12504 (N_12504,N_11939,N_11652);
or U12505 (N_12505,N_11883,N_11822);
nor U12506 (N_12506,N_11736,N_11811);
nand U12507 (N_12507,N_11638,N_11831);
nand U12508 (N_12508,N_11599,N_11572);
nor U12509 (N_12509,N_11742,N_11513);
and U12510 (N_12510,N_11564,N_11848);
xnor U12511 (N_12511,N_11345,N_11765);
xnor U12512 (N_12512,N_11422,N_11343);
nand U12513 (N_12513,N_11397,N_11671);
nand U12514 (N_12514,N_11353,N_11525);
nor U12515 (N_12515,N_11793,N_11665);
and U12516 (N_12516,N_11810,N_11677);
or U12517 (N_12517,N_11777,N_11738);
nor U12518 (N_12518,N_11549,N_11893);
nor U12519 (N_12519,N_11656,N_11304);
or U12520 (N_12520,N_11990,N_11473);
nand U12521 (N_12521,N_11722,N_11774);
or U12522 (N_12522,N_11333,N_11504);
or U12523 (N_12523,N_11566,N_11475);
nor U12524 (N_12524,N_11986,N_11662);
nor U12525 (N_12525,N_11424,N_11446);
or U12526 (N_12526,N_11928,N_11346);
nor U12527 (N_12527,N_11375,N_11876);
nor U12528 (N_12528,N_11653,N_11329);
and U12529 (N_12529,N_11979,N_11735);
and U12530 (N_12530,N_11623,N_11544);
nor U12531 (N_12531,N_11570,N_11730);
xnor U12532 (N_12532,N_11469,N_11670);
or U12533 (N_12533,N_11424,N_11594);
or U12534 (N_12534,N_11778,N_11416);
or U12535 (N_12535,N_11698,N_11986);
nand U12536 (N_12536,N_11883,N_11746);
or U12537 (N_12537,N_11311,N_11695);
nor U12538 (N_12538,N_11339,N_11556);
and U12539 (N_12539,N_11680,N_11640);
or U12540 (N_12540,N_11285,N_11402);
nor U12541 (N_12541,N_11656,N_11516);
nand U12542 (N_12542,N_11702,N_11631);
nor U12543 (N_12543,N_11476,N_11682);
nor U12544 (N_12544,N_11334,N_11930);
or U12545 (N_12545,N_11841,N_11749);
nor U12546 (N_12546,N_11753,N_11326);
or U12547 (N_12547,N_11404,N_11688);
or U12548 (N_12548,N_11691,N_11539);
or U12549 (N_12549,N_11254,N_11922);
nor U12550 (N_12550,N_11826,N_11618);
and U12551 (N_12551,N_11547,N_11259);
and U12552 (N_12552,N_11593,N_11681);
nor U12553 (N_12553,N_11625,N_11843);
nor U12554 (N_12554,N_11773,N_11600);
nand U12555 (N_12555,N_11496,N_11830);
nand U12556 (N_12556,N_11500,N_11289);
nand U12557 (N_12557,N_11395,N_11576);
nor U12558 (N_12558,N_11296,N_11899);
and U12559 (N_12559,N_11718,N_11939);
nor U12560 (N_12560,N_11663,N_11388);
nor U12561 (N_12561,N_11905,N_11509);
and U12562 (N_12562,N_11408,N_11942);
or U12563 (N_12563,N_11787,N_11751);
nand U12564 (N_12564,N_11421,N_11404);
or U12565 (N_12565,N_11704,N_11753);
xnor U12566 (N_12566,N_11543,N_11415);
and U12567 (N_12567,N_11675,N_11504);
or U12568 (N_12568,N_11719,N_11599);
xor U12569 (N_12569,N_11620,N_11327);
and U12570 (N_12570,N_11506,N_11468);
or U12571 (N_12571,N_11776,N_11635);
nand U12572 (N_12572,N_11730,N_11978);
nor U12573 (N_12573,N_11384,N_11885);
or U12574 (N_12574,N_11315,N_11344);
nand U12575 (N_12575,N_11448,N_11287);
or U12576 (N_12576,N_11348,N_11324);
nand U12577 (N_12577,N_11879,N_11852);
nand U12578 (N_12578,N_11982,N_11481);
nand U12579 (N_12579,N_11615,N_11755);
and U12580 (N_12580,N_11869,N_11706);
and U12581 (N_12581,N_11431,N_11551);
nor U12582 (N_12582,N_11383,N_11592);
or U12583 (N_12583,N_11846,N_11431);
and U12584 (N_12584,N_11778,N_11263);
or U12585 (N_12585,N_11343,N_11742);
and U12586 (N_12586,N_11728,N_11277);
nor U12587 (N_12587,N_11967,N_11472);
nand U12588 (N_12588,N_11578,N_11756);
nand U12589 (N_12589,N_11855,N_11916);
or U12590 (N_12590,N_11909,N_11758);
and U12591 (N_12591,N_11857,N_11286);
and U12592 (N_12592,N_11649,N_11891);
or U12593 (N_12593,N_11870,N_11558);
or U12594 (N_12594,N_11436,N_11542);
nand U12595 (N_12595,N_11853,N_11990);
and U12596 (N_12596,N_11953,N_11960);
or U12597 (N_12597,N_11422,N_11650);
or U12598 (N_12598,N_11641,N_11910);
and U12599 (N_12599,N_11871,N_11453);
or U12600 (N_12600,N_11869,N_11448);
nor U12601 (N_12601,N_11644,N_11607);
xor U12602 (N_12602,N_11905,N_11829);
nand U12603 (N_12603,N_11728,N_11942);
xor U12604 (N_12604,N_11864,N_11839);
or U12605 (N_12605,N_11674,N_11605);
xor U12606 (N_12606,N_11266,N_11747);
or U12607 (N_12607,N_11966,N_11819);
nand U12608 (N_12608,N_11451,N_11511);
and U12609 (N_12609,N_11340,N_11875);
nor U12610 (N_12610,N_11299,N_11268);
or U12611 (N_12611,N_11844,N_11280);
nand U12612 (N_12612,N_11497,N_11438);
nor U12613 (N_12613,N_11542,N_11352);
nand U12614 (N_12614,N_11820,N_11609);
or U12615 (N_12615,N_11976,N_11775);
nand U12616 (N_12616,N_11959,N_11288);
and U12617 (N_12617,N_11314,N_11372);
or U12618 (N_12618,N_11625,N_11333);
nor U12619 (N_12619,N_11841,N_11502);
nor U12620 (N_12620,N_11533,N_11294);
xnor U12621 (N_12621,N_11323,N_11596);
nor U12622 (N_12622,N_11278,N_11914);
nor U12623 (N_12623,N_11942,N_11622);
or U12624 (N_12624,N_11646,N_11318);
and U12625 (N_12625,N_11254,N_11417);
and U12626 (N_12626,N_11390,N_11740);
or U12627 (N_12627,N_11267,N_11780);
xor U12628 (N_12628,N_11780,N_11899);
nand U12629 (N_12629,N_11556,N_11323);
or U12630 (N_12630,N_11287,N_11356);
nor U12631 (N_12631,N_11250,N_11397);
and U12632 (N_12632,N_11695,N_11975);
or U12633 (N_12633,N_11945,N_11688);
nor U12634 (N_12634,N_11741,N_11668);
xnor U12635 (N_12635,N_11521,N_11523);
or U12636 (N_12636,N_11318,N_11799);
nand U12637 (N_12637,N_11671,N_11596);
or U12638 (N_12638,N_11742,N_11539);
nand U12639 (N_12639,N_11824,N_11561);
and U12640 (N_12640,N_11992,N_11926);
and U12641 (N_12641,N_11790,N_11875);
or U12642 (N_12642,N_11289,N_11527);
nor U12643 (N_12643,N_11863,N_11520);
nand U12644 (N_12644,N_11549,N_11947);
and U12645 (N_12645,N_11792,N_11647);
nand U12646 (N_12646,N_11529,N_11719);
and U12647 (N_12647,N_11734,N_11934);
and U12648 (N_12648,N_11938,N_11501);
and U12649 (N_12649,N_11693,N_11922);
nand U12650 (N_12650,N_11307,N_11411);
nor U12651 (N_12651,N_11840,N_11640);
nor U12652 (N_12652,N_11648,N_11837);
nand U12653 (N_12653,N_11572,N_11983);
or U12654 (N_12654,N_11924,N_11257);
and U12655 (N_12655,N_11389,N_11638);
xnor U12656 (N_12656,N_11375,N_11360);
or U12657 (N_12657,N_11539,N_11297);
or U12658 (N_12658,N_11617,N_11669);
xnor U12659 (N_12659,N_11961,N_11292);
or U12660 (N_12660,N_11945,N_11593);
or U12661 (N_12661,N_11305,N_11947);
nand U12662 (N_12662,N_11319,N_11369);
and U12663 (N_12663,N_11351,N_11446);
nor U12664 (N_12664,N_11825,N_11693);
or U12665 (N_12665,N_11512,N_11359);
nand U12666 (N_12666,N_11924,N_11585);
nand U12667 (N_12667,N_11466,N_11820);
nand U12668 (N_12668,N_11644,N_11533);
nor U12669 (N_12669,N_11437,N_11690);
xnor U12670 (N_12670,N_11909,N_11714);
and U12671 (N_12671,N_11984,N_11787);
nor U12672 (N_12672,N_11539,N_11418);
nand U12673 (N_12673,N_11298,N_11838);
nor U12674 (N_12674,N_11577,N_11526);
nand U12675 (N_12675,N_11412,N_11330);
nand U12676 (N_12676,N_11474,N_11904);
and U12677 (N_12677,N_11387,N_11497);
or U12678 (N_12678,N_11381,N_11910);
nand U12679 (N_12679,N_11716,N_11961);
and U12680 (N_12680,N_11332,N_11552);
or U12681 (N_12681,N_11630,N_11956);
xnor U12682 (N_12682,N_11551,N_11996);
and U12683 (N_12683,N_11860,N_11317);
or U12684 (N_12684,N_11923,N_11876);
nand U12685 (N_12685,N_11396,N_11833);
nor U12686 (N_12686,N_11761,N_11848);
nand U12687 (N_12687,N_11387,N_11991);
and U12688 (N_12688,N_11527,N_11920);
nand U12689 (N_12689,N_11560,N_11729);
nor U12690 (N_12690,N_11674,N_11740);
xnor U12691 (N_12691,N_11581,N_11993);
or U12692 (N_12692,N_11389,N_11472);
xor U12693 (N_12693,N_11628,N_11445);
nand U12694 (N_12694,N_11286,N_11263);
and U12695 (N_12695,N_11901,N_11823);
and U12696 (N_12696,N_11430,N_11326);
and U12697 (N_12697,N_11642,N_11549);
xnor U12698 (N_12698,N_11620,N_11551);
or U12699 (N_12699,N_11498,N_11991);
nor U12700 (N_12700,N_11840,N_11544);
or U12701 (N_12701,N_11269,N_11982);
and U12702 (N_12702,N_11435,N_11516);
nand U12703 (N_12703,N_11478,N_11666);
nor U12704 (N_12704,N_11463,N_11685);
nand U12705 (N_12705,N_11299,N_11987);
nand U12706 (N_12706,N_11682,N_11686);
nand U12707 (N_12707,N_11598,N_11275);
or U12708 (N_12708,N_11408,N_11261);
and U12709 (N_12709,N_11874,N_11944);
nand U12710 (N_12710,N_11731,N_11857);
and U12711 (N_12711,N_11744,N_11638);
or U12712 (N_12712,N_11656,N_11768);
and U12713 (N_12713,N_11840,N_11540);
nor U12714 (N_12714,N_11403,N_11267);
and U12715 (N_12715,N_11889,N_11619);
nand U12716 (N_12716,N_11526,N_11621);
nand U12717 (N_12717,N_11671,N_11393);
nand U12718 (N_12718,N_11317,N_11978);
and U12719 (N_12719,N_11904,N_11843);
and U12720 (N_12720,N_11688,N_11386);
or U12721 (N_12721,N_11654,N_11467);
nor U12722 (N_12722,N_11468,N_11974);
or U12723 (N_12723,N_11503,N_11561);
or U12724 (N_12724,N_11407,N_11866);
or U12725 (N_12725,N_11686,N_11439);
nand U12726 (N_12726,N_11265,N_11688);
or U12727 (N_12727,N_11409,N_11402);
xor U12728 (N_12728,N_11777,N_11458);
and U12729 (N_12729,N_11820,N_11487);
nor U12730 (N_12730,N_11906,N_11888);
and U12731 (N_12731,N_11401,N_11763);
or U12732 (N_12732,N_11836,N_11924);
nor U12733 (N_12733,N_11452,N_11760);
or U12734 (N_12734,N_11306,N_11991);
xor U12735 (N_12735,N_11957,N_11380);
or U12736 (N_12736,N_11301,N_11486);
nor U12737 (N_12737,N_11623,N_11991);
nor U12738 (N_12738,N_11870,N_11905);
or U12739 (N_12739,N_11813,N_11323);
nor U12740 (N_12740,N_11387,N_11288);
nand U12741 (N_12741,N_11650,N_11365);
and U12742 (N_12742,N_11614,N_11438);
or U12743 (N_12743,N_11370,N_11272);
nand U12744 (N_12744,N_11708,N_11308);
nand U12745 (N_12745,N_11874,N_11640);
and U12746 (N_12746,N_11599,N_11919);
and U12747 (N_12747,N_11857,N_11837);
or U12748 (N_12748,N_11716,N_11737);
or U12749 (N_12749,N_11500,N_11376);
or U12750 (N_12750,N_12259,N_12715);
nand U12751 (N_12751,N_12134,N_12096);
nor U12752 (N_12752,N_12670,N_12025);
xnor U12753 (N_12753,N_12466,N_12445);
and U12754 (N_12754,N_12462,N_12268);
or U12755 (N_12755,N_12142,N_12453);
or U12756 (N_12756,N_12610,N_12523);
nand U12757 (N_12757,N_12588,N_12289);
nand U12758 (N_12758,N_12544,N_12382);
nand U12759 (N_12759,N_12069,N_12214);
nor U12760 (N_12760,N_12372,N_12590);
and U12761 (N_12761,N_12529,N_12723);
xnor U12762 (N_12762,N_12235,N_12149);
nor U12763 (N_12763,N_12126,N_12180);
or U12764 (N_12764,N_12007,N_12402);
or U12765 (N_12765,N_12426,N_12266);
or U12766 (N_12766,N_12575,N_12632);
xor U12767 (N_12767,N_12179,N_12373);
nand U12768 (N_12768,N_12004,N_12495);
nand U12769 (N_12769,N_12295,N_12562);
nand U12770 (N_12770,N_12192,N_12601);
nor U12771 (N_12771,N_12571,N_12036);
xor U12772 (N_12772,N_12077,N_12135);
or U12773 (N_12773,N_12094,N_12371);
or U12774 (N_12774,N_12404,N_12207);
or U12775 (N_12775,N_12538,N_12366);
nor U12776 (N_12776,N_12370,N_12284);
and U12777 (N_12777,N_12731,N_12668);
nand U12778 (N_12778,N_12725,N_12425);
nor U12779 (N_12779,N_12526,N_12704);
nor U12780 (N_12780,N_12212,N_12068);
xnor U12781 (N_12781,N_12262,N_12394);
or U12782 (N_12782,N_12248,N_12100);
or U12783 (N_12783,N_12654,N_12010);
nor U12784 (N_12784,N_12117,N_12434);
and U12785 (N_12785,N_12230,N_12319);
or U12786 (N_12786,N_12300,N_12688);
and U12787 (N_12787,N_12076,N_12258);
nand U12788 (N_12788,N_12664,N_12124);
or U12789 (N_12789,N_12237,N_12563);
and U12790 (N_12790,N_12532,N_12517);
nor U12791 (N_12791,N_12278,N_12458);
nand U12792 (N_12792,N_12287,N_12270);
xnor U12793 (N_12793,N_12357,N_12000);
nor U12794 (N_12794,N_12543,N_12414);
nor U12795 (N_12795,N_12607,N_12323);
or U12796 (N_12796,N_12053,N_12442);
nor U12797 (N_12797,N_12566,N_12113);
nor U12798 (N_12798,N_12129,N_12141);
and U12799 (N_12799,N_12683,N_12701);
nor U12800 (N_12800,N_12556,N_12012);
nand U12801 (N_12801,N_12661,N_12732);
and U12802 (N_12802,N_12673,N_12712);
nand U12803 (N_12803,N_12509,N_12595);
and U12804 (N_12804,N_12167,N_12491);
or U12805 (N_12805,N_12619,N_12573);
and U12806 (N_12806,N_12084,N_12653);
or U12807 (N_12807,N_12220,N_12545);
nor U12808 (N_12808,N_12487,N_12616);
nand U12809 (N_12809,N_12226,N_12471);
and U12810 (N_12810,N_12508,N_12255);
or U12811 (N_12811,N_12185,N_12318);
or U12812 (N_12812,N_12660,N_12009);
xor U12813 (N_12813,N_12044,N_12510);
and U12814 (N_12814,N_12024,N_12379);
nand U12815 (N_12815,N_12005,N_12490);
nor U12816 (N_12816,N_12480,N_12349);
or U12817 (N_12817,N_12519,N_12639);
xnor U12818 (N_12818,N_12746,N_12038);
and U12819 (N_12819,N_12177,N_12350);
nor U12820 (N_12820,N_12125,N_12552);
nor U12821 (N_12821,N_12525,N_12209);
or U12822 (N_12822,N_12470,N_12283);
or U12823 (N_12823,N_12354,N_12612);
and U12824 (N_12824,N_12298,N_12099);
or U12825 (N_12825,N_12506,N_12536);
xnor U12826 (N_12826,N_12273,N_12111);
nand U12827 (N_12827,N_12496,N_12676);
or U12828 (N_12828,N_12606,N_12296);
or U12829 (N_12829,N_12033,N_12098);
xnor U12830 (N_12830,N_12474,N_12674);
nor U12831 (N_12831,N_12446,N_12368);
nand U12832 (N_12832,N_12320,N_12420);
nand U12833 (N_12833,N_12342,N_12229);
nand U12834 (N_12834,N_12339,N_12157);
nor U12835 (N_12835,N_12161,N_12691);
nor U12836 (N_12836,N_12333,N_12589);
xnor U12837 (N_12837,N_12375,N_12472);
nor U12838 (N_12838,N_12559,N_12473);
and U12839 (N_12839,N_12070,N_12669);
or U12840 (N_12840,N_12680,N_12586);
or U12841 (N_12841,N_12202,N_12694);
and U12842 (N_12842,N_12039,N_12436);
nand U12843 (N_12843,N_12223,N_12022);
nor U12844 (N_12844,N_12104,N_12599);
or U12845 (N_12845,N_12102,N_12416);
nor U12846 (N_12846,N_12254,N_12271);
or U12847 (N_12847,N_12103,N_12380);
nand U12848 (N_12848,N_12611,N_12358);
or U12849 (N_12849,N_12400,N_12017);
or U12850 (N_12850,N_12479,N_12282);
or U12851 (N_12851,N_12264,N_12250);
and U12852 (N_12852,N_12484,N_12689);
nand U12853 (N_12853,N_12722,N_12120);
and U12854 (N_12854,N_12640,N_12521);
or U12855 (N_12855,N_12208,N_12587);
nand U12856 (N_12856,N_12615,N_12585);
nand U12857 (N_12857,N_12363,N_12336);
and U12858 (N_12858,N_12636,N_12463);
and U12859 (N_12859,N_12686,N_12092);
nor U12860 (N_12860,N_12217,N_12073);
and U12861 (N_12861,N_12720,N_12170);
or U12862 (N_12862,N_12513,N_12156);
or U12863 (N_12863,N_12401,N_12623);
xor U12864 (N_12864,N_12216,N_12469);
and U12865 (N_12865,N_12430,N_12499);
nand U12866 (N_12866,N_12211,N_12376);
nand U12867 (N_12867,N_12071,N_12256);
nand U12868 (N_12868,N_12449,N_12485);
and U12869 (N_12869,N_12147,N_12742);
or U12870 (N_12870,N_12065,N_12291);
nand U12871 (N_12871,N_12310,N_12205);
nor U12872 (N_12872,N_12238,N_12154);
nand U12873 (N_12873,N_12191,N_12049);
or U12874 (N_12874,N_12501,N_12594);
or U12875 (N_12875,N_12066,N_12608);
nor U12876 (N_12876,N_12743,N_12429);
nor U12877 (N_12877,N_12634,N_12663);
nor U12878 (N_12878,N_12707,N_12037);
or U12879 (N_12879,N_12047,N_12643);
nand U12880 (N_12880,N_12432,N_12072);
and U12881 (N_12881,N_12215,N_12570);
nor U12882 (N_12882,N_12105,N_12711);
nand U12883 (N_12883,N_12080,N_12322);
and U12884 (N_12884,N_12582,N_12201);
nor U12885 (N_12885,N_12306,N_12034);
or U12886 (N_12886,N_12493,N_12130);
or U12887 (N_12887,N_12252,N_12609);
or U12888 (N_12888,N_12410,N_12074);
nand U12889 (N_12889,N_12651,N_12277);
and U12890 (N_12890,N_12138,N_12687);
nor U12891 (N_12891,N_12118,N_12326);
nand U12892 (N_12892,N_12194,N_12602);
nor U12893 (N_12893,N_12574,N_12627);
or U12894 (N_12894,N_12231,N_12481);
or U12895 (N_12895,N_12316,N_12015);
and U12896 (N_12896,N_12576,N_12247);
nand U12897 (N_12897,N_12564,N_12709);
or U12898 (N_12898,N_12655,N_12335);
or U12899 (N_12899,N_12507,N_12003);
and U12900 (N_12900,N_12435,N_12406);
or U12901 (N_12901,N_12657,N_12500);
nand U12902 (N_12902,N_12315,N_12112);
and U12903 (N_12903,N_12397,N_12269);
nand U12904 (N_12904,N_12378,N_12717);
nor U12905 (N_12905,N_12512,N_12514);
or U12906 (N_12906,N_12528,N_12160);
nand U12907 (N_12907,N_12232,N_12504);
nor U12908 (N_12908,N_12249,N_12520);
nand U12909 (N_12909,N_12679,N_12438);
nand U12910 (N_12910,N_12002,N_12530);
nand U12911 (N_12911,N_12304,N_12360);
and U12912 (N_12912,N_12086,N_12128);
nor U12913 (N_12913,N_12391,N_12275);
nand U12914 (N_12914,N_12693,N_12078);
nor U12915 (N_12915,N_12567,N_12046);
and U12916 (N_12916,N_12101,N_12381);
or U12917 (N_12917,N_12396,N_12293);
and U12918 (N_12918,N_12503,N_12557);
and U12919 (N_12919,N_12132,N_12210);
nor U12920 (N_12920,N_12516,N_12681);
xor U12921 (N_12921,N_12642,N_12219);
and U12922 (N_12922,N_12169,N_12303);
nor U12923 (N_12923,N_12706,N_12168);
xnor U12924 (N_12924,N_12454,N_12023);
and U12925 (N_12925,N_12427,N_12387);
and U12926 (N_12926,N_12240,N_12478);
nor U12927 (N_12927,N_12555,N_12183);
or U12928 (N_12928,N_12656,N_12345);
or U12929 (N_12929,N_12367,N_12311);
nand U12930 (N_12930,N_12716,N_12228);
nand U12931 (N_12931,N_12422,N_12285);
nor U12932 (N_12932,N_12062,N_12136);
xnor U12933 (N_12933,N_12647,N_12119);
nor U12934 (N_12934,N_12174,N_12253);
nor U12935 (N_12935,N_12001,N_12452);
nor U12936 (N_12936,N_12390,N_12659);
and U12937 (N_12937,N_12204,N_12551);
nor U12938 (N_12938,N_12153,N_12239);
and U12939 (N_12939,N_12419,N_12451);
or U12940 (N_12940,N_12173,N_12620);
nand U12941 (N_12941,N_12067,N_12733);
xor U12942 (N_12942,N_12748,N_12355);
and U12943 (N_12943,N_12286,N_12121);
xnor U12944 (N_12944,N_12677,N_12393);
and U12945 (N_12945,N_12637,N_12139);
nand U12946 (N_12946,N_12030,N_12534);
nor U12947 (N_12947,N_12464,N_12597);
or U12948 (N_12948,N_12714,N_12447);
and U12949 (N_12949,N_12302,N_12411);
nor U12950 (N_12950,N_12016,N_12644);
nand U12951 (N_12951,N_12383,N_12392);
xnor U12952 (N_12952,N_12362,N_12352);
nor U12953 (N_12953,N_12635,N_12106);
or U12954 (N_12954,N_12618,N_12245);
and U12955 (N_12955,N_12337,N_12133);
or U12956 (N_12956,N_12041,N_12054);
nor U12957 (N_12957,N_12417,N_12568);
or U12958 (N_12958,N_12386,N_12241);
nor U12959 (N_12959,N_12407,N_12384);
or U12960 (N_12960,N_12629,N_12537);
nand U12961 (N_12961,N_12163,N_12624);
and U12962 (N_12962,N_12553,N_12307);
or U12963 (N_12963,N_12389,N_12724);
nor U12964 (N_12964,N_12622,N_12482);
or U12965 (N_12965,N_12081,N_12581);
nand U12966 (N_12966,N_12043,N_12539);
or U12967 (N_12967,N_12364,N_12088);
nor U12968 (N_12968,N_12527,N_12515);
nor U12969 (N_12969,N_12408,N_12008);
xnor U12970 (N_12970,N_12189,N_12329);
nand U12971 (N_12971,N_12361,N_12308);
nor U12972 (N_12972,N_12540,N_12467);
or U12973 (N_12973,N_12684,N_12492);
or U12974 (N_12974,N_12421,N_12511);
nand U12975 (N_12975,N_12460,N_12164);
and U12976 (N_12976,N_12747,N_12730);
and U12977 (N_12977,N_12468,N_12261);
xor U12978 (N_12978,N_12475,N_12292);
and U12979 (N_12979,N_12060,N_12018);
nor U12980 (N_12980,N_12107,N_12267);
nor U12981 (N_12981,N_12621,N_12083);
nand U12982 (N_12982,N_12744,N_12699);
or U12983 (N_12983,N_12144,N_12328);
and U12984 (N_12984,N_12448,N_12726);
and U12985 (N_12985,N_12423,N_12524);
nor U12986 (N_12986,N_12522,N_12341);
nand U12987 (N_12987,N_12064,N_12171);
nor U12988 (N_12988,N_12351,N_12583);
and U12989 (N_12989,N_12176,N_12734);
nand U12990 (N_12990,N_12705,N_12288);
or U12991 (N_12991,N_12572,N_12184);
and U12992 (N_12992,N_12330,N_12741);
or U12993 (N_12993,N_12110,N_12166);
and U12994 (N_12994,N_12641,N_12646);
nor U12995 (N_12995,N_12388,N_12692);
and U12996 (N_12996,N_12721,N_12200);
and U12997 (N_12997,N_12549,N_12405);
or U12998 (N_12998,N_12672,N_12159);
or U12999 (N_12999,N_12444,N_12035);
xor U13000 (N_13000,N_12122,N_12152);
nand U13001 (N_13001,N_12398,N_12281);
xor U13002 (N_13002,N_12151,N_12045);
nand U13003 (N_13003,N_12127,N_12598);
nor U13004 (N_13004,N_12150,N_12658);
and U13005 (N_13005,N_12505,N_12497);
or U13006 (N_13006,N_12145,N_12312);
or U13007 (N_13007,N_12093,N_12225);
or U13008 (N_13008,N_12666,N_12195);
and U13009 (N_13009,N_12346,N_12090);
nor U13010 (N_13010,N_12014,N_12662);
nand U13011 (N_13011,N_12050,N_12645);
nand U13012 (N_13012,N_12456,N_12187);
or U13013 (N_13013,N_12580,N_12206);
nand U13014 (N_13014,N_12413,N_12535);
nor U13015 (N_13015,N_12246,N_12338);
nor U13016 (N_13016,N_12309,N_12546);
and U13017 (N_13017,N_12652,N_12548);
nand U13018 (N_13018,N_12085,N_12675);
and U13019 (N_13019,N_12181,N_12224);
or U13020 (N_13020,N_12440,N_12502);
nand U13021 (N_13021,N_12332,N_12542);
nand U13022 (N_13022,N_12087,N_12600);
nand U13023 (N_13023,N_12531,N_12011);
nand U13024 (N_13024,N_12604,N_12115);
xnor U13025 (N_13025,N_12348,N_12097);
or U13026 (N_13026,N_12584,N_12075);
nor U13027 (N_13027,N_12745,N_12353);
nor U13028 (N_13028,N_12441,N_12554);
nand U13029 (N_13029,N_12199,N_12671);
or U13030 (N_13030,N_12457,N_12146);
xnor U13031 (N_13031,N_12137,N_12317);
nand U13032 (N_13032,N_12737,N_12148);
nand U13033 (N_13033,N_12477,N_12028);
nand U13034 (N_13034,N_12603,N_12061);
or U13035 (N_13035,N_12158,N_12213);
and U13036 (N_13036,N_12299,N_12729);
nor U13037 (N_13037,N_12412,N_12057);
and U13038 (N_13038,N_12243,N_12667);
nand U13039 (N_13039,N_12428,N_12578);
nand U13040 (N_13040,N_12029,N_12665);
xnor U13041 (N_13041,N_12569,N_12633);
nor U13042 (N_13042,N_12626,N_12131);
and U13043 (N_13043,N_12631,N_12344);
nand U13044 (N_13044,N_12082,N_12718);
nand U13045 (N_13045,N_12091,N_12280);
or U13046 (N_13046,N_12221,N_12533);
nand U13047 (N_13047,N_12385,N_12109);
and U13048 (N_13048,N_12596,N_12260);
and U13049 (N_13049,N_12347,N_12026);
nor U13050 (N_13050,N_12359,N_12042);
and U13051 (N_13051,N_12749,N_12314);
xor U13052 (N_13052,N_12162,N_12728);
nand U13053 (N_13053,N_12695,N_12565);
or U13054 (N_13054,N_12019,N_12331);
or U13055 (N_13055,N_12678,N_12196);
and U13056 (N_13056,N_12648,N_12058);
nor U13057 (N_13057,N_12172,N_12403);
nand U13058 (N_13058,N_12251,N_12186);
and U13059 (N_13059,N_12579,N_12418);
and U13060 (N_13060,N_12356,N_12739);
and U13061 (N_13061,N_12188,N_12297);
nand U13062 (N_13062,N_12052,N_12257);
nor U13063 (N_13063,N_12031,N_12374);
xor U13064 (N_13064,N_12272,N_12461);
nand U13065 (N_13065,N_12108,N_12305);
nor U13066 (N_13066,N_12114,N_12279);
and U13067 (N_13067,N_12301,N_12321);
or U13068 (N_13068,N_12040,N_12313);
nor U13069 (N_13069,N_12055,N_12193);
nand U13070 (N_13070,N_12409,N_12494);
nor U13071 (N_13071,N_12630,N_12614);
and U13072 (N_13072,N_12095,N_12577);
and U13073 (N_13073,N_12327,N_12738);
or U13074 (N_13074,N_12592,N_12274);
nand U13075 (N_13075,N_12561,N_12735);
or U13076 (N_13076,N_12431,N_12365);
nand U13077 (N_13077,N_12051,N_12116);
nor U13078 (N_13078,N_12708,N_12476);
nand U13079 (N_13079,N_12605,N_12343);
nand U13080 (N_13080,N_12027,N_12340);
or U13081 (N_13081,N_12056,N_12294);
nand U13082 (N_13082,N_12190,N_12020);
nand U13083 (N_13083,N_12740,N_12593);
and U13084 (N_13084,N_12334,N_12560);
nand U13085 (N_13085,N_12182,N_12483);
nand U13086 (N_13086,N_12702,N_12063);
and U13087 (N_13087,N_12059,N_12465);
nand U13088 (N_13088,N_12227,N_12222);
or U13089 (N_13089,N_12625,N_12617);
and U13090 (N_13090,N_12234,N_12650);
nand U13091 (N_13091,N_12591,N_12518);
and U13092 (N_13092,N_12123,N_12710);
nand U13093 (N_13093,N_12486,N_12489);
or U13094 (N_13094,N_12558,N_12263);
nand U13095 (N_13095,N_12175,N_12424);
and U13096 (N_13096,N_12218,N_12415);
or U13097 (N_13097,N_12233,N_12439);
nor U13098 (N_13098,N_12165,N_12433);
nand U13099 (N_13099,N_12155,N_12703);
nor U13100 (N_13100,N_12638,N_12399);
nor U13101 (N_13101,N_12443,N_12547);
nor U13102 (N_13102,N_12140,N_12048);
nand U13103 (N_13103,N_12455,N_12541);
nand U13104 (N_13104,N_12325,N_12628);
and U13105 (N_13105,N_12324,N_12719);
xor U13106 (N_13106,N_12143,N_12682);
xor U13107 (N_13107,N_12488,N_12613);
xnor U13108 (N_13108,N_12203,N_12032);
and U13109 (N_13109,N_12685,N_12696);
and U13110 (N_13110,N_12021,N_12197);
nand U13111 (N_13111,N_12698,N_12713);
and U13112 (N_13112,N_12697,N_12178);
nor U13113 (N_13113,N_12089,N_12727);
nor U13114 (N_13114,N_12198,N_12450);
nor U13115 (N_13115,N_12369,N_12690);
nand U13116 (N_13116,N_12276,N_12006);
nor U13117 (N_13117,N_12550,N_12244);
xor U13118 (N_13118,N_12437,N_12242);
nor U13119 (N_13119,N_12459,N_12265);
xnor U13120 (N_13120,N_12736,N_12649);
or U13121 (N_13121,N_12236,N_12290);
xnor U13122 (N_13122,N_12377,N_12498);
nand U13123 (N_13123,N_12079,N_12395);
xnor U13124 (N_13124,N_12013,N_12700);
and U13125 (N_13125,N_12341,N_12688);
or U13126 (N_13126,N_12746,N_12650);
nor U13127 (N_13127,N_12320,N_12158);
or U13128 (N_13128,N_12501,N_12210);
or U13129 (N_13129,N_12746,N_12318);
nand U13130 (N_13130,N_12471,N_12684);
nor U13131 (N_13131,N_12326,N_12373);
xnor U13132 (N_13132,N_12062,N_12708);
and U13133 (N_13133,N_12711,N_12517);
xor U13134 (N_13134,N_12316,N_12620);
nor U13135 (N_13135,N_12494,N_12495);
or U13136 (N_13136,N_12181,N_12354);
or U13137 (N_13137,N_12319,N_12564);
nor U13138 (N_13138,N_12297,N_12540);
or U13139 (N_13139,N_12222,N_12009);
nand U13140 (N_13140,N_12505,N_12715);
nand U13141 (N_13141,N_12309,N_12621);
xnor U13142 (N_13142,N_12092,N_12429);
nor U13143 (N_13143,N_12635,N_12334);
nand U13144 (N_13144,N_12699,N_12622);
or U13145 (N_13145,N_12192,N_12184);
and U13146 (N_13146,N_12669,N_12259);
and U13147 (N_13147,N_12733,N_12249);
and U13148 (N_13148,N_12512,N_12288);
nor U13149 (N_13149,N_12426,N_12614);
and U13150 (N_13150,N_12300,N_12682);
nand U13151 (N_13151,N_12709,N_12204);
nand U13152 (N_13152,N_12275,N_12410);
and U13153 (N_13153,N_12254,N_12430);
and U13154 (N_13154,N_12065,N_12668);
nand U13155 (N_13155,N_12415,N_12003);
nand U13156 (N_13156,N_12111,N_12394);
or U13157 (N_13157,N_12028,N_12202);
or U13158 (N_13158,N_12336,N_12285);
xnor U13159 (N_13159,N_12657,N_12139);
nand U13160 (N_13160,N_12542,N_12476);
xnor U13161 (N_13161,N_12183,N_12308);
xor U13162 (N_13162,N_12532,N_12672);
or U13163 (N_13163,N_12650,N_12345);
nand U13164 (N_13164,N_12514,N_12714);
or U13165 (N_13165,N_12455,N_12317);
nor U13166 (N_13166,N_12045,N_12399);
nor U13167 (N_13167,N_12747,N_12621);
or U13168 (N_13168,N_12156,N_12567);
xnor U13169 (N_13169,N_12496,N_12722);
or U13170 (N_13170,N_12445,N_12131);
nor U13171 (N_13171,N_12294,N_12321);
xnor U13172 (N_13172,N_12682,N_12156);
nor U13173 (N_13173,N_12547,N_12410);
nand U13174 (N_13174,N_12001,N_12305);
and U13175 (N_13175,N_12593,N_12293);
nand U13176 (N_13176,N_12024,N_12146);
and U13177 (N_13177,N_12115,N_12360);
xnor U13178 (N_13178,N_12062,N_12020);
and U13179 (N_13179,N_12735,N_12515);
and U13180 (N_13180,N_12502,N_12718);
nand U13181 (N_13181,N_12251,N_12344);
or U13182 (N_13182,N_12259,N_12713);
and U13183 (N_13183,N_12535,N_12106);
nand U13184 (N_13184,N_12636,N_12233);
or U13185 (N_13185,N_12434,N_12672);
xnor U13186 (N_13186,N_12085,N_12266);
nand U13187 (N_13187,N_12291,N_12098);
nand U13188 (N_13188,N_12306,N_12450);
xnor U13189 (N_13189,N_12376,N_12069);
nand U13190 (N_13190,N_12481,N_12645);
xor U13191 (N_13191,N_12420,N_12428);
nand U13192 (N_13192,N_12177,N_12670);
nor U13193 (N_13193,N_12346,N_12032);
or U13194 (N_13194,N_12548,N_12427);
nand U13195 (N_13195,N_12694,N_12291);
nor U13196 (N_13196,N_12176,N_12177);
nor U13197 (N_13197,N_12632,N_12572);
nand U13198 (N_13198,N_12502,N_12451);
nor U13199 (N_13199,N_12156,N_12204);
nor U13200 (N_13200,N_12516,N_12032);
and U13201 (N_13201,N_12315,N_12221);
nor U13202 (N_13202,N_12540,N_12572);
and U13203 (N_13203,N_12366,N_12498);
and U13204 (N_13204,N_12298,N_12590);
nand U13205 (N_13205,N_12390,N_12675);
or U13206 (N_13206,N_12396,N_12459);
nor U13207 (N_13207,N_12329,N_12732);
nand U13208 (N_13208,N_12388,N_12744);
nor U13209 (N_13209,N_12676,N_12026);
nor U13210 (N_13210,N_12285,N_12114);
or U13211 (N_13211,N_12709,N_12397);
nor U13212 (N_13212,N_12012,N_12040);
nor U13213 (N_13213,N_12615,N_12213);
or U13214 (N_13214,N_12249,N_12614);
nand U13215 (N_13215,N_12137,N_12486);
nand U13216 (N_13216,N_12251,N_12309);
nor U13217 (N_13217,N_12613,N_12645);
and U13218 (N_13218,N_12537,N_12683);
nand U13219 (N_13219,N_12008,N_12738);
nand U13220 (N_13220,N_12309,N_12090);
or U13221 (N_13221,N_12535,N_12107);
and U13222 (N_13222,N_12526,N_12198);
nor U13223 (N_13223,N_12601,N_12478);
and U13224 (N_13224,N_12444,N_12111);
and U13225 (N_13225,N_12000,N_12375);
and U13226 (N_13226,N_12528,N_12413);
or U13227 (N_13227,N_12069,N_12319);
nor U13228 (N_13228,N_12580,N_12438);
or U13229 (N_13229,N_12641,N_12407);
xor U13230 (N_13230,N_12744,N_12359);
and U13231 (N_13231,N_12421,N_12207);
and U13232 (N_13232,N_12394,N_12376);
nand U13233 (N_13233,N_12041,N_12731);
or U13234 (N_13234,N_12470,N_12538);
or U13235 (N_13235,N_12368,N_12667);
nor U13236 (N_13236,N_12584,N_12701);
nor U13237 (N_13237,N_12041,N_12245);
and U13238 (N_13238,N_12143,N_12116);
nand U13239 (N_13239,N_12493,N_12405);
nand U13240 (N_13240,N_12009,N_12507);
nand U13241 (N_13241,N_12667,N_12719);
xor U13242 (N_13242,N_12693,N_12040);
nand U13243 (N_13243,N_12075,N_12478);
or U13244 (N_13244,N_12124,N_12097);
nor U13245 (N_13245,N_12094,N_12682);
and U13246 (N_13246,N_12195,N_12062);
and U13247 (N_13247,N_12167,N_12448);
xnor U13248 (N_13248,N_12590,N_12156);
xor U13249 (N_13249,N_12303,N_12322);
nand U13250 (N_13250,N_12546,N_12533);
or U13251 (N_13251,N_12347,N_12293);
or U13252 (N_13252,N_12650,N_12748);
or U13253 (N_13253,N_12605,N_12237);
nor U13254 (N_13254,N_12544,N_12047);
nor U13255 (N_13255,N_12602,N_12184);
nor U13256 (N_13256,N_12278,N_12066);
or U13257 (N_13257,N_12066,N_12320);
nand U13258 (N_13258,N_12586,N_12204);
or U13259 (N_13259,N_12687,N_12028);
xnor U13260 (N_13260,N_12118,N_12035);
or U13261 (N_13261,N_12371,N_12262);
or U13262 (N_13262,N_12058,N_12277);
or U13263 (N_13263,N_12732,N_12411);
or U13264 (N_13264,N_12746,N_12268);
or U13265 (N_13265,N_12172,N_12284);
xor U13266 (N_13266,N_12217,N_12513);
nor U13267 (N_13267,N_12427,N_12267);
and U13268 (N_13268,N_12580,N_12602);
or U13269 (N_13269,N_12349,N_12269);
or U13270 (N_13270,N_12659,N_12213);
nor U13271 (N_13271,N_12728,N_12060);
xor U13272 (N_13272,N_12144,N_12578);
and U13273 (N_13273,N_12477,N_12601);
nand U13274 (N_13274,N_12546,N_12481);
and U13275 (N_13275,N_12024,N_12054);
xor U13276 (N_13276,N_12392,N_12655);
nand U13277 (N_13277,N_12331,N_12296);
nor U13278 (N_13278,N_12432,N_12711);
or U13279 (N_13279,N_12100,N_12632);
and U13280 (N_13280,N_12438,N_12589);
nor U13281 (N_13281,N_12455,N_12428);
and U13282 (N_13282,N_12206,N_12160);
nand U13283 (N_13283,N_12311,N_12312);
and U13284 (N_13284,N_12733,N_12047);
nor U13285 (N_13285,N_12604,N_12526);
nor U13286 (N_13286,N_12039,N_12560);
or U13287 (N_13287,N_12712,N_12605);
or U13288 (N_13288,N_12358,N_12641);
or U13289 (N_13289,N_12515,N_12037);
nor U13290 (N_13290,N_12296,N_12325);
nor U13291 (N_13291,N_12613,N_12299);
nor U13292 (N_13292,N_12644,N_12467);
nor U13293 (N_13293,N_12653,N_12326);
or U13294 (N_13294,N_12422,N_12277);
nand U13295 (N_13295,N_12273,N_12159);
nor U13296 (N_13296,N_12302,N_12156);
and U13297 (N_13297,N_12693,N_12158);
nor U13298 (N_13298,N_12356,N_12162);
or U13299 (N_13299,N_12024,N_12537);
nor U13300 (N_13300,N_12450,N_12647);
nand U13301 (N_13301,N_12242,N_12253);
nor U13302 (N_13302,N_12076,N_12560);
nor U13303 (N_13303,N_12071,N_12487);
xor U13304 (N_13304,N_12423,N_12092);
nor U13305 (N_13305,N_12005,N_12672);
and U13306 (N_13306,N_12563,N_12293);
nand U13307 (N_13307,N_12530,N_12682);
or U13308 (N_13308,N_12337,N_12548);
nand U13309 (N_13309,N_12578,N_12080);
and U13310 (N_13310,N_12406,N_12480);
or U13311 (N_13311,N_12129,N_12545);
nor U13312 (N_13312,N_12028,N_12198);
or U13313 (N_13313,N_12000,N_12344);
nor U13314 (N_13314,N_12506,N_12636);
nor U13315 (N_13315,N_12523,N_12469);
and U13316 (N_13316,N_12277,N_12151);
or U13317 (N_13317,N_12548,N_12565);
nor U13318 (N_13318,N_12724,N_12485);
nand U13319 (N_13319,N_12494,N_12147);
and U13320 (N_13320,N_12506,N_12571);
xor U13321 (N_13321,N_12315,N_12050);
nor U13322 (N_13322,N_12047,N_12632);
xnor U13323 (N_13323,N_12007,N_12018);
xor U13324 (N_13324,N_12042,N_12080);
or U13325 (N_13325,N_12124,N_12121);
or U13326 (N_13326,N_12247,N_12079);
and U13327 (N_13327,N_12312,N_12023);
and U13328 (N_13328,N_12648,N_12380);
or U13329 (N_13329,N_12596,N_12509);
nand U13330 (N_13330,N_12737,N_12107);
or U13331 (N_13331,N_12337,N_12583);
or U13332 (N_13332,N_12115,N_12695);
nor U13333 (N_13333,N_12017,N_12505);
nor U13334 (N_13334,N_12609,N_12026);
or U13335 (N_13335,N_12047,N_12662);
xor U13336 (N_13336,N_12401,N_12422);
and U13337 (N_13337,N_12634,N_12520);
nor U13338 (N_13338,N_12075,N_12109);
and U13339 (N_13339,N_12077,N_12440);
or U13340 (N_13340,N_12261,N_12274);
and U13341 (N_13341,N_12536,N_12154);
nand U13342 (N_13342,N_12515,N_12039);
and U13343 (N_13343,N_12605,N_12699);
or U13344 (N_13344,N_12083,N_12691);
or U13345 (N_13345,N_12434,N_12438);
and U13346 (N_13346,N_12377,N_12626);
xnor U13347 (N_13347,N_12493,N_12315);
and U13348 (N_13348,N_12614,N_12143);
and U13349 (N_13349,N_12596,N_12295);
or U13350 (N_13350,N_12506,N_12542);
nor U13351 (N_13351,N_12502,N_12120);
or U13352 (N_13352,N_12570,N_12387);
nand U13353 (N_13353,N_12033,N_12572);
xnor U13354 (N_13354,N_12312,N_12564);
xor U13355 (N_13355,N_12608,N_12263);
and U13356 (N_13356,N_12029,N_12232);
nand U13357 (N_13357,N_12519,N_12383);
and U13358 (N_13358,N_12413,N_12265);
or U13359 (N_13359,N_12593,N_12185);
and U13360 (N_13360,N_12739,N_12189);
nand U13361 (N_13361,N_12444,N_12278);
and U13362 (N_13362,N_12296,N_12498);
or U13363 (N_13363,N_12294,N_12359);
and U13364 (N_13364,N_12529,N_12514);
nor U13365 (N_13365,N_12336,N_12581);
and U13366 (N_13366,N_12633,N_12643);
nor U13367 (N_13367,N_12098,N_12644);
nand U13368 (N_13368,N_12293,N_12052);
nor U13369 (N_13369,N_12353,N_12192);
nor U13370 (N_13370,N_12728,N_12030);
nor U13371 (N_13371,N_12715,N_12217);
xnor U13372 (N_13372,N_12413,N_12433);
and U13373 (N_13373,N_12042,N_12268);
and U13374 (N_13374,N_12118,N_12551);
or U13375 (N_13375,N_12227,N_12628);
xor U13376 (N_13376,N_12051,N_12416);
xor U13377 (N_13377,N_12193,N_12062);
and U13378 (N_13378,N_12130,N_12302);
nand U13379 (N_13379,N_12208,N_12411);
nor U13380 (N_13380,N_12153,N_12629);
nand U13381 (N_13381,N_12551,N_12518);
nor U13382 (N_13382,N_12412,N_12611);
xnor U13383 (N_13383,N_12379,N_12000);
nand U13384 (N_13384,N_12123,N_12110);
or U13385 (N_13385,N_12025,N_12150);
and U13386 (N_13386,N_12415,N_12724);
or U13387 (N_13387,N_12147,N_12311);
or U13388 (N_13388,N_12136,N_12605);
and U13389 (N_13389,N_12428,N_12352);
nand U13390 (N_13390,N_12460,N_12136);
nor U13391 (N_13391,N_12057,N_12054);
nand U13392 (N_13392,N_12146,N_12663);
nor U13393 (N_13393,N_12420,N_12021);
nor U13394 (N_13394,N_12681,N_12465);
nand U13395 (N_13395,N_12545,N_12287);
or U13396 (N_13396,N_12723,N_12694);
or U13397 (N_13397,N_12525,N_12000);
nor U13398 (N_13398,N_12464,N_12728);
and U13399 (N_13399,N_12330,N_12666);
and U13400 (N_13400,N_12696,N_12488);
or U13401 (N_13401,N_12187,N_12279);
nand U13402 (N_13402,N_12044,N_12715);
or U13403 (N_13403,N_12749,N_12719);
nand U13404 (N_13404,N_12261,N_12354);
nand U13405 (N_13405,N_12110,N_12480);
or U13406 (N_13406,N_12422,N_12429);
nand U13407 (N_13407,N_12092,N_12056);
nand U13408 (N_13408,N_12048,N_12649);
nor U13409 (N_13409,N_12116,N_12583);
nand U13410 (N_13410,N_12044,N_12368);
and U13411 (N_13411,N_12080,N_12736);
nand U13412 (N_13412,N_12175,N_12235);
xnor U13413 (N_13413,N_12076,N_12586);
nand U13414 (N_13414,N_12329,N_12505);
nand U13415 (N_13415,N_12327,N_12255);
nor U13416 (N_13416,N_12633,N_12543);
nor U13417 (N_13417,N_12530,N_12545);
nand U13418 (N_13418,N_12021,N_12154);
nor U13419 (N_13419,N_12021,N_12063);
and U13420 (N_13420,N_12498,N_12742);
and U13421 (N_13421,N_12037,N_12577);
or U13422 (N_13422,N_12628,N_12163);
or U13423 (N_13423,N_12010,N_12260);
and U13424 (N_13424,N_12661,N_12136);
nor U13425 (N_13425,N_12085,N_12227);
or U13426 (N_13426,N_12156,N_12741);
nand U13427 (N_13427,N_12673,N_12547);
nor U13428 (N_13428,N_12108,N_12663);
or U13429 (N_13429,N_12086,N_12303);
nand U13430 (N_13430,N_12494,N_12306);
nand U13431 (N_13431,N_12206,N_12127);
and U13432 (N_13432,N_12053,N_12620);
nand U13433 (N_13433,N_12116,N_12662);
or U13434 (N_13434,N_12079,N_12003);
xnor U13435 (N_13435,N_12723,N_12584);
nand U13436 (N_13436,N_12714,N_12707);
or U13437 (N_13437,N_12738,N_12238);
and U13438 (N_13438,N_12148,N_12178);
or U13439 (N_13439,N_12550,N_12285);
nor U13440 (N_13440,N_12254,N_12574);
or U13441 (N_13441,N_12384,N_12150);
nand U13442 (N_13442,N_12170,N_12390);
or U13443 (N_13443,N_12613,N_12699);
xor U13444 (N_13444,N_12098,N_12510);
and U13445 (N_13445,N_12435,N_12428);
nor U13446 (N_13446,N_12016,N_12238);
and U13447 (N_13447,N_12742,N_12680);
and U13448 (N_13448,N_12062,N_12524);
and U13449 (N_13449,N_12366,N_12488);
nand U13450 (N_13450,N_12191,N_12319);
xor U13451 (N_13451,N_12459,N_12665);
and U13452 (N_13452,N_12719,N_12742);
nand U13453 (N_13453,N_12376,N_12441);
or U13454 (N_13454,N_12259,N_12010);
nand U13455 (N_13455,N_12151,N_12495);
nor U13456 (N_13456,N_12511,N_12312);
xor U13457 (N_13457,N_12371,N_12035);
nand U13458 (N_13458,N_12240,N_12632);
nor U13459 (N_13459,N_12418,N_12629);
or U13460 (N_13460,N_12197,N_12191);
and U13461 (N_13461,N_12180,N_12314);
nor U13462 (N_13462,N_12504,N_12371);
and U13463 (N_13463,N_12031,N_12255);
nor U13464 (N_13464,N_12481,N_12662);
or U13465 (N_13465,N_12496,N_12113);
or U13466 (N_13466,N_12108,N_12454);
and U13467 (N_13467,N_12307,N_12317);
nor U13468 (N_13468,N_12604,N_12045);
and U13469 (N_13469,N_12496,N_12639);
nor U13470 (N_13470,N_12648,N_12402);
nor U13471 (N_13471,N_12724,N_12232);
xnor U13472 (N_13472,N_12746,N_12705);
or U13473 (N_13473,N_12165,N_12266);
or U13474 (N_13474,N_12558,N_12405);
nor U13475 (N_13475,N_12007,N_12458);
nor U13476 (N_13476,N_12065,N_12636);
nor U13477 (N_13477,N_12736,N_12269);
and U13478 (N_13478,N_12748,N_12312);
nand U13479 (N_13479,N_12293,N_12336);
or U13480 (N_13480,N_12439,N_12711);
nor U13481 (N_13481,N_12579,N_12299);
nand U13482 (N_13482,N_12302,N_12341);
nand U13483 (N_13483,N_12403,N_12602);
nand U13484 (N_13484,N_12520,N_12255);
and U13485 (N_13485,N_12275,N_12451);
or U13486 (N_13486,N_12546,N_12462);
xor U13487 (N_13487,N_12705,N_12340);
and U13488 (N_13488,N_12733,N_12185);
nor U13489 (N_13489,N_12285,N_12163);
xor U13490 (N_13490,N_12538,N_12402);
nand U13491 (N_13491,N_12160,N_12219);
nand U13492 (N_13492,N_12635,N_12162);
nor U13493 (N_13493,N_12359,N_12698);
and U13494 (N_13494,N_12584,N_12201);
nor U13495 (N_13495,N_12116,N_12059);
and U13496 (N_13496,N_12266,N_12370);
nor U13497 (N_13497,N_12241,N_12465);
and U13498 (N_13498,N_12512,N_12076);
nor U13499 (N_13499,N_12382,N_12146);
nand U13500 (N_13500,N_12758,N_13395);
nor U13501 (N_13501,N_13011,N_12808);
nor U13502 (N_13502,N_12843,N_13465);
nand U13503 (N_13503,N_13073,N_13091);
nand U13504 (N_13504,N_12786,N_13057);
or U13505 (N_13505,N_13228,N_12753);
or U13506 (N_13506,N_12809,N_12761);
nand U13507 (N_13507,N_12989,N_13229);
nor U13508 (N_13508,N_13356,N_13428);
nand U13509 (N_13509,N_13315,N_12764);
nor U13510 (N_13510,N_12958,N_13263);
xor U13511 (N_13511,N_12838,N_13481);
or U13512 (N_13512,N_13497,N_13137);
nand U13513 (N_13513,N_12842,N_12861);
or U13514 (N_13514,N_13443,N_12840);
nand U13515 (N_13515,N_13201,N_13109);
and U13516 (N_13516,N_13043,N_13096);
and U13517 (N_13517,N_13289,N_13028);
nor U13518 (N_13518,N_13132,N_12961);
or U13519 (N_13519,N_13247,N_13006);
and U13520 (N_13520,N_13189,N_13184);
and U13521 (N_13521,N_13400,N_13479);
or U13522 (N_13522,N_13188,N_12994);
xnor U13523 (N_13523,N_13143,N_13203);
nand U13524 (N_13524,N_13482,N_13080);
nor U13525 (N_13525,N_12879,N_12960);
nor U13526 (N_13526,N_12763,N_12990);
or U13527 (N_13527,N_13179,N_12798);
or U13528 (N_13528,N_13357,N_12965);
and U13529 (N_13529,N_13217,N_12897);
or U13530 (N_13530,N_13471,N_12797);
nand U13531 (N_13531,N_12848,N_13025);
or U13532 (N_13532,N_13204,N_13024);
or U13533 (N_13533,N_13301,N_13077);
nor U13534 (N_13534,N_13379,N_13216);
nor U13535 (N_13535,N_12818,N_12765);
or U13536 (N_13536,N_13448,N_12777);
nand U13537 (N_13537,N_13139,N_12854);
nand U13538 (N_13538,N_13238,N_13361);
or U13539 (N_13539,N_13036,N_13276);
nor U13540 (N_13540,N_13150,N_13198);
xor U13541 (N_13541,N_13283,N_13153);
and U13542 (N_13542,N_13351,N_12756);
xor U13543 (N_13543,N_13230,N_12956);
and U13544 (N_13544,N_13103,N_13222);
nor U13545 (N_13545,N_12948,N_12817);
and U13546 (N_13546,N_13224,N_12874);
nor U13547 (N_13547,N_12906,N_12849);
nor U13548 (N_13548,N_13031,N_13061);
and U13549 (N_13549,N_12853,N_13253);
and U13550 (N_13550,N_13429,N_13082);
nor U13551 (N_13551,N_13450,N_12917);
or U13552 (N_13552,N_13377,N_13368);
nor U13553 (N_13553,N_13492,N_13172);
nand U13554 (N_13554,N_12949,N_12912);
or U13555 (N_13555,N_13250,N_13162);
nor U13556 (N_13556,N_13393,N_12881);
or U13557 (N_13557,N_13176,N_13020);
xor U13558 (N_13558,N_13272,N_12770);
nand U13559 (N_13559,N_13474,N_13107);
nor U13560 (N_13560,N_12884,N_12785);
nor U13561 (N_13561,N_12776,N_12779);
and U13562 (N_13562,N_12830,N_13273);
or U13563 (N_13563,N_13427,N_12875);
or U13564 (N_13564,N_12913,N_13062);
nand U13565 (N_13565,N_13420,N_13262);
and U13566 (N_13566,N_13047,N_12922);
nor U13567 (N_13567,N_13072,N_12782);
nor U13568 (N_13568,N_13241,N_13209);
and U13569 (N_13569,N_13392,N_13175);
nand U13570 (N_13570,N_13329,N_13015);
nor U13571 (N_13571,N_13453,N_12919);
nor U13572 (N_13572,N_13245,N_12951);
nand U13573 (N_13573,N_13292,N_12970);
nor U13574 (N_13574,N_13088,N_13434);
or U13575 (N_13575,N_12821,N_13307);
or U13576 (N_13576,N_12997,N_12751);
nor U13577 (N_13577,N_13449,N_12939);
nand U13578 (N_13578,N_13168,N_12787);
nand U13579 (N_13579,N_13439,N_13341);
and U13580 (N_13580,N_12932,N_12992);
nand U13581 (N_13581,N_13063,N_12986);
nand U13582 (N_13582,N_12841,N_13322);
and U13583 (N_13583,N_13375,N_13042);
nand U13584 (N_13584,N_13323,N_12819);
xnor U13585 (N_13585,N_13312,N_12898);
nand U13586 (N_13586,N_13067,N_13265);
or U13587 (N_13587,N_12893,N_13141);
and U13588 (N_13588,N_13051,N_13009);
nor U13589 (N_13589,N_13462,N_12952);
and U13590 (N_13590,N_13214,N_13249);
and U13591 (N_13591,N_13074,N_12928);
nor U13592 (N_13592,N_13252,N_12868);
nand U13593 (N_13593,N_13333,N_13338);
nand U13594 (N_13594,N_12988,N_13394);
or U13595 (N_13595,N_13331,N_13019);
nor U13596 (N_13596,N_13306,N_13156);
xor U13597 (N_13597,N_13363,N_12971);
nor U13598 (N_13598,N_13076,N_13342);
and U13599 (N_13599,N_12832,N_13003);
nand U13600 (N_13600,N_13018,N_13084);
and U13601 (N_13601,N_12903,N_12945);
and U13602 (N_13602,N_13410,N_13382);
nor U13603 (N_13603,N_13012,N_13258);
or U13604 (N_13604,N_13405,N_13447);
xnor U13605 (N_13605,N_12882,N_12752);
or U13606 (N_13606,N_13220,N_13336);
nand U13607 (N_13607,N_13367,N_12966);
nor U13608 (N_13608,N_13475,N_12845);
and U13609 (N_13609,N_13346,N_12839);
or U13610 (N_13610,N_12804,N_12826);
and U13611 (N_13611,N_13381,N_13083);
or U13612 (N_13612,N_12806,N_12831);
nand U13613 (N_13613,N_13494,N_12857);
xor U13614 (N_13614,N_12967,N_13303);
nor U13615 (N_13615,N_13264,N_13243);
and U13616 (N_13616,N_13463,N_12944);
and U13617 (N_13617,N_12869,N_13488);
xor U13618 (N_13618,N_12978,N_13399);
and U13619 (N_13619,N_13149,N_13235);
nand U13620 (N_13620,N_12864,N_13455);
or U13621 (N_13621,N_13196,N_13040);
nor U13622 (N_13622,N_13498,N_13456);
nor U13623 (N_13623,N_13483,N_12921);
nor U13624 (N_13624,N_13060,N_13349);
nor U13625 (N_13625,N_13069,N_13218);
nand U13626 (N_13626,N_13070,N_13099);
and U13627 (N_13627,N_13111,N_13305);
or U13628 (N_13628,N_13105,N_13412);
nand U13629 (N_13629,N_13360,N_13202);
and U13630 (N_13630,N_12969,N_12955);
or U13631 (N_13631,N_13293,N_13138);
nor U13632 (N_13632,N_13350,N_13219);
xnor U13633 (N_13633,N_13387,N_12825);
nand U13634 (N_13634,N_13248,N_13325);
nor U13635 (N_13635,N_13454,N_12995);
xor U13636 (N_13636,N_13476,N_13207);
and U13637 (N_13637,N_13499,N_12911);
nand U13638 (N_13638,N_13423,N_12982);
nor U13639 (N_13639,N_13424,N_13376);
and U13640 (N_13640,N_13173,N_13255);
and U13641 (N_13641,N_13421,N_13416);
nand U13642 (N_13642,N_13390,N_13308);
and U13643 (N_13643,N_13092,N_13407);
nand U13644 (N_13644,N_13195,N_13186);
nand U13645 (N_13645,N_13436,N_13371);
xor U13646 (N_13646,N_13147,N_13413);
and U13647 (N_13647,N_12866,N_13284);
and U13648 (N_13648,N_13116,N_13237);
and U13649 (N_13649,N_13050,N_12933);
nand U13650 (N_13650,N_13117,N_13151);
and U13651 (N_13651,N_13389,N_13268);
nand U13652 (N_13652,N_13190,N_13496);
nor U13653 (N_13653,N_13213,N_13348);
and U13654 (N_13654,N_13089,N_13300);
nand U13655 (N_13655,N_13364,N_13441);
nand U13656 (N_13656,N_13016,N_13226);
nor U13657 (N_13657,N_13282,N_13317);
nand U13658 (N_13658,N_12867,N_12800);
or U13659 (N_13659,N_13052,N_13490);
nor U13660 (N_13660,N_13267,N_13032);
nor U13661 (N_13661,N_13459,N_13221);
nand U13662 (N_13662,N_13145,N_12943);
nor U13663 (N_13663,N_13347,N_13055);
or U13664 (N_13664,N_13468,N_13417);
nor U13665 (N_13665,N_13337,N_12996);
or U13666 (N_13666,N_13155,N_12810);
or U13667 (N_13667,N_13166,N_13039);
nand U13668 (N_13668,N_13098,N_13435);
nand U13669 (N_13669,N_13286,N_13440);
or U13670 (N_13670,N_13005,N_13075);
nand U13671 (N_13671,N_13194,N_13071);
and U13672 (N_13672,N_12811,N_12894);
nor U13673 (N_13673,N_13287,N_13438);
and U13674 (N_13674,N_13451,N_12936);
nor U13675 (N_13675,N_13174,N_13004);
xnor U13676 (N_13676,N_13081,N_13053);
nand U13677 (N_13677,N_13185,N_13345);
nand U13678 (N_13678,N_12915,N_12851);
nor U13679 (N_13679,N_13119,N_12780);
or U13680 (N_13680,N_12883,N_13373);
nor U13681 (N_13681,N_12937,N_13232);
and U13682 (N_13682,N_12895,N_12759);
nand U13683 (N_13683,N_13113,N_13008);
nor U13684 (N_13684,N_13260,N_13285);
nor U13685 (N_13685,N_13157,N_13118);
and U13686 (N_13686,N_13415,N_12794);
nand U13687 (N_13687,N_13326,N_13383);
or U13688 (N_13688,N_13487,N_12999);
or U13689 (N_13689,N_13414,N_12834);
nor U13690 (N_13690,N_13123,N_13135);
and U13691 (N_13691,N_13034,N_13396);
xor U13692 (N_13692,N_13161,N_13340);
nor U13693 (N_13693,N_13128,N_12892);
xor U13694 (N_13694,N_13183,N_13058);
or U13695 (N_13695,N_13000,N_13457);
nand U13696 (N_13696,N_13140,N_13205);
nand U13697 (N_13697,N_13130,N_13495);
xnor U13698 (N_13698,N_12899,N_13320);
or U13699 (N_13699,N_13104,N_13355);
xor U13700 (N_13700,N_12750,N_13261);
nand U13701 (N_13701,N_13425,N_13484);
and U13702 (N_13702,N_13313,N_12773);
and U13703 (N_13703,N_12812,N_12799);
nor U13704 (N_13704,N_13225,N_13171);
and U13705 (N_13705,N_12896,N_12822);
or U13706 (N_13706,N_13002,N_13419);
xor U13707 (N_13707,N_13134,N_13056);
nand U13708 (N_13708,N_13120,N_12791);
nor U13709 (N_13709,N_12938,N_12946);
nand U13710 (N_13710,N_12863,N_13299);
nor U13711 (N_13711,N_13402,N_13266);
nor U13712 (N_13712,N_13352,N_13404);
nand U13713 (N_13713,N_12934,N_13170);
and U13714 (N_13714,N_12846,N_13027);
or U13715 (N_13715,N_12918,N_12950);
or U13716 (N_13716,N_13411,N_12998);
or U13717 (N_13717,N_12796,N_12959);
nor U13718 (N_13718,N_13023,N_12901);
nand U13719 (N_13719,N_13038,N_12844);
nor U13720 (N_13720,N_13281,N_12766);
nor U13721 (N_13721,N_13452,N_13131);
nor U13722 (N_13722,N_13021,N_12859);
or U13723 (N_13723,N_13277,N_12823);
nor U13724 (N_13724,N_13246,N_12813);
or U13725 (N_13725,N_12914,N_12803);
nor U13726 (N_13726,N_12940,N_12957);
nor U13727 (N_13727,N_13279,N_13146);
or U13728 (N_13728,N_13328,N_12762);
or U13729 (N_13729,N_12908,N_12792);
nand U13730 (N_13730,N_12916,N_12835);
nor U13731 (N_13731,N_13254,N_12755);
nand U13732 (N_13732,N_12870,N_13234);
nor U13733 (N_13733,N_12850,N_13065);
nor U13734 (N_13734,N_12980,N_13469);
xor U13735 (N_13735,N_13112,N_12828);
and U13736 (N_13736,N_12953,N_12991);
nor U13737 (N_13737,N_13491,N_12860);
nor U13738 (N_13738,N_12816,N_13339);
nor U13739 (N_13739,N_13477,N_12983);
and U13740 (N_13740,N_13401,N_13485);
nor U13741 (N_13741,N_13212,N_12981);
and U13742 (N_13742,N_12923,N_13354);
nor U13743 (N_13743,N_12880,N_13197);
or U13744 (N_13744,N_13374,N_12772);
xor U13745 (N_13745,N_12941,N_13295);
and U13746 (N_13746,N_13180,N_12836);
nor U13747 (N_13747,N_12963,N_13480);
nand U13748 (N_13748,N_13100,N_12907);
or U13749 (N_13749,N_13126,N_13291);
nand U13750 (N_13750,N_13288,N_13433);
nor U13751 (N_13751,N_12873,N_13101);
and U13752 (N_13752,N_13125,N_12972);
nand U13753 (N_13753,N_13369,N_12784);
and U13754 (N_13754,N_12962,N_12886);
or U13755 (N_13755,N_13208,N_12814);
nor U13756 (N_13756,N_12977,N_13398);
and U13757 (N_13757,N_13037,N_12775);
nor U13758 (N_13758,N_13473,N_13041);
nand U13759 (N_13759,N_13122,N_12942);
or U13760 (N_13760,N_13359,N_13259);
and U13761 (N_13761,N_13311,N_13330);
or U13762 (N_13762,N_13085,N_13432);
nand U13763 (N_13763,N_13159,N_13193);
or U13764 (N_13764,N_13403,N_13233);
xor U13765 (N_13765,N_13178,N_13321);
nand U13766 (N_13766,N_13182,N_13437);
xor U13767 (N_13767,N_13310,N_12891);
or U13768 (N_13768,N_12789,N_13046);
and U13769 (N_13769,N_13385,N_13114);
nand U13770 (N_13770,N_12769,N_12909);
nor U13771 (N_13771,N_12820,N_13271);
nand U13772 (N_13772,N_12872,N_13332);
and U13773 (N_13773,N_13489,N_13422);
nor U13774 (N_13774,N_13380,N_13418);
and U13775 (N_13775,N_13470,N_13211);
nand U13776 (N_13776,N_13270,N_13094);
and U13777 (N_13777,N_12760,N_13378);
and U13778 (N_13778,N_13033,N_13242);
xor U13779 (N_13779,N_12968,N_12887);
and U13780 (N_13780,N_12829,N_13054);
xnor U13781 (N_13781,N_13294,N_13239);
nor U13782 (N_13782,N_13090,N_13318);
nand U13783 (N_13783,N_12795,N_13466);
nor U13784 (N_13784,N_13030,N_13335);
nand U13785 (N_13785,N_13129,N_13160);
xnor U13786 (N_13786,N_13158,N_12774);
nand U13787 (N_13787,N_13210,N_12757);
nand U13788 (N_13788,N_13014,N_12805);
or U13789 (N_13789,N_13296,N_12973);
or U13790 (N_13790,N_12993,N_13464);
nor U13791 (N_13791,N_12947,N_13044);
nor U13792 (N_13792,N_13215,N_13256);
nand U13793 (N_13793,N_13165,N_13409);
nand U13794 (N_13794,N_12871,N_12771);
or U13795 (N_13795,N_13244,N_12904);
nand U13796 (N_13796,N_13251,N_13314);
or U13797 (N_13797,N_13372,N_13115);
or U13798 (N_13798,N_12890,N_13257);
nand U13799 (N_13799,N_13064,N_12802);
and U13800 (N_13800,N_12768,N_12862);
or U13801 (N_13801,N_12865,N_13431);
nor U13802 (N_13802,N_12927,N_13017);
and U13803 (N_13803,N_13493,N_13446);
nor U13804 (N_13804,N_13384,N_12815);
nand U13805 (N_13805,N_12926,N_13144);
nor U13806 (N_13806,N_12793,N_13154);
nand U13807 (N_13807,N_13366,N_13280);
or U13808 (N_13808,N_13007,N_13124);
and U13809 (N_13809,N_13269,N_13049);
or U13810 (N_13810,N_12976,N_13467);
and U13811 (N_13811,N_12778,N_12888);
nor U13812 (N_13812,N_13444,N_13133);
nor U13813 (N_13813,N_13231,N_13048);
nor U13814 (N_13814,N_13045,N_13461);
nand U13815 (N_13815,N_12889,N_13309);
and U13816 (N_13816,N_12827,N_13426);
or U13817 (N_13817,N_12783,N_13079);
xor U13818 (N_13818,N_12858,N_12985);
nor U13819 (N_13819,N_13121,N_13035);
nor U13820 (N_13820,N_13106,N_13386);
nand U13821 (N_13821,N_12856,N_13164);
and U13822 (N_13822,N_12935,N_12984);
or U13823 (N_13823,N_13302,N_12931);
and U13824 (N_13824,N_13066,N_12974);
nand U13825 (N_13825,N_13191,N_12807);
nor U13826 (N_13826,N_13142,N_13319);
and U13827 (N_13827,N_12788,N_13458);
nand U13828 (N_13828,N_13199,N_13324);
or U13829 (N_13829,N_13127,N_13148);
nand U13830 (N_13830,N_13278,N_12900);
and U13831 (N_13831,N_13478,N_13353);
or U13832 (N_13832,N_13223,N_12878);
nand U13833 (N_13833,N_12979,N_13022);
and U13834 (N_13834,N_13445,N_12824);
nor U13835 (N_13835,N_13472,N_13068);
or U13836 (N_13836,N_13290,N_12975);
or U13837 (N_13837,N_12964,N_13391);
nand U13838 (N_13838,N_12930,N_13181);
xor U13839 (N_13839,N_12885,N_12837);
or U13840 (N_13840,N_12855,N_13152);
xnor U13841 (N_13841,N_13240,N_13343);
and U13842 (N_13842,N_13406,N_13236);
nand U13843 (N_13843,N_13327,N_13274);
and U13844 (N_13844,N_12754,N_13200);
or U13845 (N_13845,N_12910,N_13334);
or U13846 (N_13846,N_13086,N_13460);
and U13847 (N_13847,N_13227,N_12924);
and U13848 (N_13848,N_12902,N_12833);
nand U13849 (N_13849,N_13408,N_13187);
nand U13850 (N_13850,N_13097,N_13026);
nor U13851 (N_13851,N_12790,N_12905);
and U13852 (N_13852,N_13304,N_13430);
xnor U13853 (N_13853,N_12954,N_12801);
nand U13854 (N_13854,N_13177,N_13275);
or U13855 (N_13855,N_12987,N_12781);
nand U13856 (N_13856,N_13059,N_13362);
nor U13857 (N_13857,N_13365,N_12876);
and U13858 (N_13858,N_13316,N_13108);
or U13859 (N_13859,N_13167,N_13136);
nand U13860 (N_13860,N_13442,N_13093);
nand U13861 (N_13861,N_13001,N_12852);
nand U13862 (N_13862,N_13169,N_13486);
and U13863 (N_13863,N_13029,N_13192);
and U13864 (N_13864,N_13397,N_13370);
nor U13865 (N_13865,N_13102,N_13110);
nand U13866 (N_13866,N_13344,N_12925);
and U13867 (N_13867,N_12929,N_13078);
xnor U13868 (N_13868,N_13388,N_13095);
nor U13869 (N_13869,N_13298,N_13297);
or U13870 (N_13870,N_13163,N_12877);
or U13871 (N_13871,N_13087,N_13013);
nor U13872 (N_13872,N_13358,N_13010);
xor U13873 (N_13873,N_13206,N_12847);
nor U13874 (N_13874,N_12767,N_12920);
or U13875 (N_13875,N_12757,N_13215);
nand U13876 (N_13876,N_12917,N_13175);
xor U13877 (N_13877,N_13214,N_13442);
nand U13878 (N_13878,N_13212,N_12904);
nand U13879 (N_13879,N_12767,N_13459);
nor U13880 (N_13880,N_13436,N_13123);
and U13881 (N_13881,N_13003,N_12836);
xor U13882 (N_13882,N_12938,N_13334);
xnor U13883 (N_13883,N_13169,N_13027);
or U13884 (N_13884,N_13163,N_13330);
nor U13885 (N_13885,N_13148,N_13315);
and U13886 (N_13886,N_13078,N_13449);
nor U13887 (N_13887,N_13374,N_13255);
and U13888 (N_13888,N_13248,N_13260);
xnor U13889 (N_13889,N_12948,N_13090);
and U13890 (N_13890,N_13301,N_13237);
nor U13891 (N_13891,N_13386,N_13442);
nand U13892 (N_13892,N_13102,N_13270);
nor U13893 (N_13893,N_13038,N_12786);
and U13894 (N_13894,N_12986,N_13331);
nor U13895 (N_13895,N_13294,N_13189);
and U13896 (N_13896,N_13196,N_13200);
and U13897 (N_13897,N_13397,N_13410);
nor U13898 (N_13898,N_12755,N_12838);
nand U13899 (N_13899,N_12793,N_13122);
or U13900 (N_13900,N_13178,N_13291);
xnor U13901 (N_13901,N_13203,N_13223);
nor U13902 (N_13902,N_12971,N_12909);
or U13903 (N_13903,N_12797,N_13267);
nor U13904 (N_13904,N_13406,N_12839);
or U13905 (N_13905,N_13278,N_12853);
nor U13906 (N_13906,N_13479,N_13078);
and U13907 (N_13907,N_12940,N_13410);
nor U13908 (N_13908,N_12786,N_12825);
and U13909 (N_13909,N_13467,N_13246);
nor U13910 (N_13910,N_13475,N_13493);
nand U13911 (N_13911,N_13398,N_13434);
or U13912 (N_13912,N_13033,N_13020);
xnor U13913 (N_13913,N_13048,N_13054);
xor U13914 (N_13914,N_13444,N_13104);
or U13915 (N_13915,N_13363,N_13195);
nand U13916 (N_13916,N_13300,N_13211);
nand U13917 (N_13917,N_12844,N_12785);
nor U13918 (N_13918,N_13496,N_13474);
xnor U13919 (N_13919,N_12900,N_13353);
and U13920 (N_13920,N_13203,N_13051);
nor U13921 (N_13921,N_13302,N_13258);
and U13922 (N_13922,N_13134,N_13307);
nand U13923 (N_13923,N_12921,N_12996);
nor U13924 (N_13924,N_12944,N_13167);
or U13925 (N_13925,N_12793,N_13091);
or U13926 (N_13926,N_13157,N_13243);
or U13927 (N_13927,N_13156,N_12941);
and U13928 (N_13928,N_12848,N_13362);
nor U13929 (N_13929,N_13162,N_13313);
and U13930 (N_13930,N_13302,N_12850);
nand U13931 (N_13931,N_12979,N_12974);
or U13932 (N_13932,N_13150,N_12822);
xor U13933 (N_13933,N_12992,N_12908);
nor U13934 (N_13934,N_12815,N_12988);
and U13935 (N_13935,N_13020,N_13128);
and U13936 (N_13936,N_12947,N_13045);
and U13937 (N_13937,N_13182,N_13166);
nand U13938 (N_13938,N_13284,N_12841);
nand U13939 (N_13939,N_13461,N_12988);
nand U13940 (N_13940,N_12986,N_13150);
nor U13941 (N_13941,N_12767,N_13007);
nand U13942 (N_13942,N_13223,N_13346);
nor U13943 (N_13943,N_13030,N_13152);
and U13944 (N_13944,N_12815,N_13216);
and U13945 (N_13945,N_13482,N_13189);
nor U13946 (N_13946,N_13238,N_13170);
and U13947 (N_13947,N_13483,N_13056);
xnor U13948 (N_13948,N_13265,N_13079);
or U13949 (N_13949,N_13241,N_13198);
or U13950 (N_13950,N_13078,N_12851);
nor U13951 (N_13951,N_13441,N_13387);
nor U13952 (N_13952,N_13341,N_13053);
nand U13953 (N_13953,N_13050,N_13385);
or U13954 (N_13954,N_13099,N_12928);
and U13955 (N_13955,N_13302,N_12820);
or U13956 (N_13956,N_13412,N_12784);
xor U13957 (N_13957,N_13244,N_13066);
or U13958 (N_13958,N_13490,N_13141);
nand U13959 (N_13959,N_12782,N_13053);
xnor U13960 (N_13960,N_13006,N_12873);
and U13961 (N_13961,N_13156,N_13099);
and U13962 (N_13962,N_13389,N_13273);
and U13963 (N_13963,N_12990,N_12764);
and U13964 (N_13964,N_13047,N_13113);
and U13965 (N_13965,N_12967,N_12763);
nor U13966 (N_13966,N_13141,N_13360);
xnor U13967 (N_13967,N_13003,N_12922);
xor U13968 (N_13968,N_13194,N_12992);
nor U13969 (N_13969,N_13089,N_13113);
nor U13970 (N_13970,N_13318,N_13423);
nor U13971 (N_13971,N_12993,N_13183);
xor U13972 (N_13972,N_12836,N_13421);
nor U13973 (N_13973,N_13324,N_12994);
and U13974 (N_13974,N_12778,N_13498);
nor U13975 (N_13975,N_13252,N_13393);
or U13976 (N_13976,N_13017,N_13124);
xnor U13977 (N_13977,N_13018,N_13182);
xor U13978 (N_13978,N_12890,N_12926);
and U13979 (N_13979,N_12803,N_12906);
nor U13980 (N_13980,N_13122,N_13355);
and U13981 (N_13981,N_13015,N_13397);
nor U13982 (N_13982,N_13280,N_13236);
or U13983 (N_13983,N_12933,N_13460);
or U13984 (N_13984,N_13415,N_12878);
or U13985 (N_13985,N_12951,N_12997);
nor U13986 (N_13986,N_13125,N_13432);
nor U13987 (N_13987,N_13136,N_12842);
and U13988 (N_13988,N_13457,N_13393);
and U13989 (N_13989,N_13285,N_13402);
xnor U13990 (N_13990,N_12993,N_13031);
or U13991 (N_13991,N_12798,N_13003);
nand U13992 (N_13992,N_12917,N_13019);
and U13993 (N_13993,N_13410,N_13238);
nand U13994 (N_13994,N_13470,N_13365);
and U13995 (N_13995,N_13495,N_12904);
nand U13996 (N_13996,N_13471,N_12841);
nor U13997 (N_13997,N_12991,N_13303);
and U13998 (N_13998,N_13350,N_12765);
nand U13999 (N_13999,N_12949,N_13233);
nand U14000 (N_14000,N_13129,N_13367);
or U14001 (N_14001,N_13040,N_13306);
or U14002 (N_14002,N_13109,N_12832);
xor U14003 (N_14003,N_13021,N_12840);
nand U14004 (N_14004,N_13161,N_13191);
and U14005 (N_14005,N_13243,N_13309);
and U14006 (N_14006,N_13167,N_13424);
and U14007 (N_14007,N_12776,N_13105);
and U14008 (N_14008,N_13038,N_13333);
or U14009 (N_14009,N_13004,N_13039);
or U14010 (N_14010,N_13449,N_13408);
nor U14011 (N_14011,N_13274,N_13034);
or U14012 (N_14012,N_13472,N_13171);
and U14013 (N_14013,N_13062,N_13069);
nand U14014 (N_14014,N_13019,N_13418);
or U14015 (N_14015,N_13119,N_13212);
nand U14016 (N_14016,N_13376,N_13269);
or U14017 (N_14017,N_13487,N_13295);
nand U14018 (N_14018,N_12837,N_13309);
nor U14019 (N_14019,N_13402,N_13100);
and U14020 (N_14020,N_12844,N_13108);
and U14021 (N_14021,N_13029,N_13007);
nor U14022 (N_14022,N_13495,N_13180);
nor U14023 (N_14023,N_13105,N_13167);
and U14024 (N_14024,N_13106,N_13187);
or U14025 (N_14025,N_13188,N_12879);
and U14026 (N_14026,N_13141,N_12763);
and U14027 (N_14027,N_13375,N_13356);
and U14028 (N_14028,N_12875,N_12787);
nor U14029 (N_14029,N_12985,N_13451);
nand U14030 (N_14030,N_13198,N_13349);
nand U14031 (N_14031,N_12820,N_13390);
nor U14032 (N_14032,N_13124,N_13481);
nand U14033 (N_14033,N_13088,N_12879);
xor U14034 (N_14034,N_12790,N_12772);
or U14035 (N_14035,N_13218,N_12984);
and U14036 (N_14036,N_12880,N_12888);
and U14037 (N_14037,N_12788,N_12782);
or U14038 (N_14038,N_12863,N_12841);
or U14039 (N_14039,N_12858,N_13059);
or U14040 (N_14040,N_13378,N_13328);
nor U14041 (N_14041,N_12779,N_13341);
or U14042 (N_14042,N_12947,N_12889);
and U14043 (N_14043,N_13335,N_13272);
nand U14044 (N_14044,N_13154,N_13285);
xor U14045 (N_14045,N_12814,N_13188);
and U14046 (N_14046,N_13489,N_13161);
nand U14047 (N_14047,N_13256,N_13388);
or U14048 (N_14048,N_13305,N_13276);
nor U14049 (N_14049,N_13204,N_12909);
nand U14050 (N_14050,N_13460,N_13041);
and U14051 (N_14051,N_13071,N_13145);
nor U14052 (N_14052,N_13153,N_12904);
nand U14053 (N_14053,N_13194,N_13032);
nor U14054 (N_14054,N_12781,N_13031);
nor U14055 (N_14055,N_13057,N_13104);
nor U14056 (N_14056,N_13441,N_12990);
nand U14057 (N_14057,N_12900,N_12997);
nand U14058 (N_14058,N_12974,N_12793);
or U14059 (N_14059,N_12808,N_13215);
or U14060 (N_14060,N_13313,N_12966);
or U14061 (N_14061,N_13436,N_12952);
or U14062 (N_14062,N_12846,N_13465);
nor U14063 (N_14063,N_12893,N_12814);
nor U14064 (N_14064,N_13438,N_12850);
or U14065 (N_14065,N_13261,N_12772);
or U14066 (N_14066,N_13474,N_12845);
or U14067 (N_14067,N_13418,N_13003);
nand U14068 (N_14068,N_13488,N_12953);
nor U14069 (N_14069,N_13042,N_12898);
or U14070 (N_14070,N_13457,N_13134);
nor U14071 (N_14071,N_13062,N_12879);
xor U14072 (N_14072,N_12967,N_12877);
and U14073 (N_14073,N_13469,N_12775);
nand U14074 (N_14074,N_12999,N_13452);
and U14075 (N_14075,N_12761,N_13491);
or U14076 (N_14076,N_13035,N_13113);
nor U14077 (N_14077,N_13255,N_13084);
nand U14078 (N_14078,N_12997,N_13317);
and U14079 (N_14079,N_13408,N_13137);
nor U14080 (N_14080,N_13416,N_13254);
nand U14081 (N_14081,N_13153,N_12835);
or U14082 (N_14082,N_13406,N_13105);
and U14083 (N_14083,N_13423,N_12896);
xnor U14084 (N_14084,N_13324,N_12888);
nor U14085 (N_14085,N_13461,N_13117);
or U14086 (N_14086,N_13118,N_12867);
nand U14087 (N_14087,N_13379,N_13231);
and U14088 (N_14088,N_13097,N_13496);
nor U14089 (N_14089,N_13163,N_13257);
nand U14090 (N_14090,N_12864,N_13407);
and U14091 (N_14091,N_13496,N_13038);
or U14092 (N_14092,N_12892,N_13410);
and U14093 (N_14093,N_12969,N_12755);
nor U14094 (N_14094,N_13011,N_13417);
or U14095 (N_14095,N_12881,N_13088);
nand U14096 (N_14096,N_13451,N_13327);
and U14097 (N_14097,N_13213,N_13303);
or U14098 (N_14098,N_13087,N_12811);
or U14099 (N_14099,N_13082,N_12939);
and U14100 (N_14100,N_13165,N_13428);
nand U14101 (N_14101,N_13024,N_13375);
and U14102 (N_14102,N_13099,N_13296);
and U14103 (N_14103,N_12807,N_13015);
nand U14104 (N_14104,N_13068,N_13181);
or U14105 (N_14105,N_13119,N_13307);
xor U14106 (N_14106,N_12980,N_13078);
nand U14107 (N_14107,N_13220,N_12967);
nand U14108 (N_14108,N_13142,N_12836);
nor U14109 (N_14109,N_13252,N_13349);
or U14110 (N_14110,N_13365,N_13293);
and U14111 (N_14111,N_13076,N_13014);
xor U14112 (N_14112,N_13283,N_13222);
nand U14113 (N_14113,N_12922,N_12997);
or U14114 (N_14114,N_13030,N_13445);
and U14115 (N_14115,N_13495,N_13270);
or U14116 (N_14116,N_13034,N_12785);
and U14117 (N_14117,N_13232,N_13031);
or U14118 (N_14118,N_12846,N_13209);
or U14119 (N_14119,N_13327,N_12855);
nand U14120 (N_14120,N_13359,N_12935);
nand U14121 (N_14121,N_13175,N_12881);
nor U14122 (N_14122,N_12814,N_12829);
and U14123 (N_14123,N_13234,N_13074);
or U14124 (N_14124,N_13401,N_12802);
and U14125 (N_14125,N_13020,N_13385);
or U14126 (N_14126,N_13433,N_13099);
and U14127 (N_14127,N_13423,N_12917);
nand U14128 (N_14128,N_13478,N_12795);
xor U14129 (N_14129,N_13142,N_13271);
or U14130 (N_14130,N_13497,N_12851);
and U14131 (N_14131,N_12794,N_13012);
or U14132 (N_14132,N_13084,N_12832);
or U14133 (N_14133,N_13012,N_13259);
nor U14134 (N_14134,N_12756,N_13495);
xor U14135 (N_14135,N_13198,N_13000);
xnor U14136 (N_14136,N_13455,N_12966);
nand U14137 (N_14137,N_12985,N_13492);
and U14138 (N_14138,N_13071,N_12888);
nor U14139 (N_14139,N_13308,N_12832);
nand U14140 (N_14140,N_13389,N_12804);
nor U14141 (N_14141,N_13362,N_12807);
or U14142 (N_14142,N_13366,N_12838);
and U14143 (N_14143,N_12995,N_13440);
and U14144 (N_14144,N_13132,N_12932);
or U14145 (N_14145,N_13152,N_13198);
nand U14146 (N_14146,N_13487,N_13240);
or U14147 (N_14147,N_12996,N_12817);
xor U14148 (N_14148,N_12924,N_13167);
or U14149 (N_14149,N_12786,N_13263);
nand U14150 (N_14150,N_13330,N_13099);
nand U14151 (N_14151,N_12882,N_12879);
nor U14152 (N_14152,N_13473,N_13323);
nor U14153 (N_14153,N_13076,N_12761);
nor U14154 (N_14154,N_13328,N_13010);
nor U14155 (N_14155,N_13079,N_12758);
nor U14156 (N_14156,N_13176,N_13115);
nor U14157 (N_14157,N_12822,N_13408);
or U14158 (N_14158,N_12859,N_13465);
and U14159 (N_14159,N_13175,N_13011);
and U14160 (N_14160,N_12755,N_12934);
and U14161 (N_14161,N_13019,N_13249);
nor U14162 (N_14162,N_13143,N_13208);
and U14163 (N_14163,N_13495,N_13388);
nand U14164 (N_14164,N_13283,N_13329);
nor U14165 (N_14165,N_12941,N_13032);
nand U14166 (N_14166,N_13314,N_12818);
or U14167 (N_14167,N_12967,N_13479);
and U14168 (N_14168,N_13374,N_13062);
and U14169 (N_14169,N_13234,N_12956);
nor U14170 (N_14170,N_13375,N_13108);
or U14171 (N_14171,N_13354,N_13098);
and U14172 (N_14172,N_13128,N_13405);
or U14173 (N_14173,N_13237,N_13451);
nor U14174 (N_14174,N_13391,N_13480);
xor U14175 (N_14175,N_13328,N_12750);
and U14176 (N_14176,N_13230,N_12808);
or U14177 (N_14177,N_12898,N_13440);
or U14178 (N_14178,N_13356,N_13383);
xnor U14179 (N_14179,N_13441,N_13428);
xor U14180 (N_14180,N_12794,N_12943);
and U14181 (N_14181,N_13313,N_13474);
and U14182 (N_14182,N_13198,N_13061);
or U14183 (N_14183,N_13034,N_12931);
xor U14184 (N_14184,N_12802,N_13405);
nand U14185 (N_14185,N_13016,N_12751);
or U14186 (N_14186,N_13431,N_12802);
nand U14187 (N_14187,N_13059,N_12857);
and U14188 (N_14188,N_13257,N_12786);
or U14189 (N_14189,N_12832,N_13126);
or U14190 (N_14190,N_13316,N_13110);
or U14191 (N_14191,N_12875,N_13329);
and U14192 (N_14192,N_13186,N_12834);
nor U14193 (N_14193,N_13374,N_13051);
and U14194 (N_14194,N_13276,N_12948);
nand U14195 (N_14195,N_13256,N_12819);
or U14196 (N_14196,N_13463,N_13420);
nor U14197 (N_14197,N_12845,N_13246);
nand U14198 (N_14198,N_13449,N_13445);
nor U14199 (N_14199,N_13186,N_13293);
xnor U14200 (N_14200,N_12916,N_12909);
and U14201 (N_14201,N_13418,N_13487);
nand U14202 (N_14202,N_13461,N_13331);
nor U14203 (N_14203,N_13276,N_13079);
and U14204 (N_14204,N_13381,N_13472);
and U14205 (N_14205,N_12914,N_13253);
nand U14206 (N_14206,N_13021,N_12878);
nand U14207 (N_14207,N_13319,N_13400);
and U14208 (N_14208,N_12932,N_12985);
nor U14209 (N_14209,N_13038,N_13058);
xor U14210 (N_14210,N_12811,N_12895);
or U14211 (N_14211,N_12795,N_12813);
and U14212 (N_14212,N_13341,N_13495);
nand U14213 (N_14213,N_13345,N_12866);
xnor U14214 (N_14214,N_13312,N_13277);
and U14215 (N_14215,N_12840,N_13285);
or U14216 (N_14216,N_13485,N_13146);
nor U14217 (N_14217,N_13243,N_13225);
or U14218 (N_14218,N_13113,N_13495);
nor U14219 (N_14219,N_12969,N_13066);
and U14220 (N_14220,N_12816,N_12963);
or U14221 (N_14221,N_12825,N_13336);
nand U14222 (N_14222,N_13120,N_13164);
xnor U14223 (N_14223,N_12754,N_13003);
nor U14224 (N_14224,N_13158,N_12835);
nor U14225 (N_14225,N_13265,N_13251);
nor U14226 (N_14226,N_13308,N_13113);
nand U14227 (N_14227,N_12996,N_13396);
and U14228 (N_14228,N_12756,N_13018);
and U14229 (N_14229,N_12927,N_12838);
and U14230 (N_14230,N_12798,N_13157);
or U14231 (N_14231,N_13327,N_13061);
or U14232 (N_14232,N_13206,N_13045);
and U14233 (N_14233,N_13319,N_13345);
nor U14234 (N_14234,N_13320,N_13230);
nand U14235 (N_14235,N_13477,N_12970);
nor U14236 (N_14236,N_12949,N_13368);
or U14237 (N_14237,N_13223,N_13020);
nor U14238 (N_14238,N_13488,N_13210);
nor U14239 (N_14239,N_13218,N_13015);
nand U14240 (N_14240,N_13482,N_13287);
and U14241 (N_14241,N_13310,N_13012);
nor U14242 (N_14242,N_12853,N_12880);
xor U14243 (N_14243,N_13115,N_13243);
or U14244 (N_14244,N_12982,N_12917);
nor U14245 (N_14245,N_13189,N_12901);
or U14246 (N_14246,N_13009,N_12911);
and U14247 (N_14247,N_13119,N_13053);
xnor U14248 (N_14248,N_12945,N_12929);
and U14249 (N_14249,N_13345,N_13499);
and U14250 (N_14250,N_14119,N_13870);
or U14251 (N_14251,N_13943,N_13923);
nor U14252 (N_14252,N_14227,N_13929);
or U14253 (N_14253,N_13796,N_13700);
and U14254 (N_14254,N_13793,N_13734);
or U14255 (N_14255,N_13656,N_14208);
and U14256 (N_14256,N_13890,N_13524);
nand U14257 (N_14257,N_13722,N_13758);
nor U14258 (N_14258,N_13939,N_13748);
nand U14259 (N_14259,N_14017,N_14078);
xor U14260 (N_14260,N_13540,N_13692);
or U14261 (N_14261,N_13837,N_14077);
or U14262 (N_14262,N_13761,N_14135);
or U14263 (N_14263,N_13736,N_13717);
nor U14264 (N_14264,N_13694,N_14029);
nor U14265 (N_14265,N_13500,N_13725);
and U14266 (N_14266,N_13671,N_13518);
or U14267 (N_14267,N_13538,N_14195);
and U14268 (N_14268,N_13760,N_13888);
or U14269 (N_14269,N_13655,N_13836);
and U14270 (N_14270,N_14101,N_13969);
nand U14271 (N_14271,N_14187,N_13823);
nor U14272 (N_14272,N_14116,N_13997);
nor U14273 (N_14273,N_13642,N_13513);
nand U14274 (N_14274,N_13814,N_14231);
or U14275 (N_14275,N_13665,N_13653);
or U14276 (N_14276,N_14000,N_13530);
nand U14277 (N_14277,N_13921,N_13644);
nor U14278 (N_14278,N_13527,N_14100);
and U14279 (N_14279,N_14160,N_14164);
nand U14280 (N_14280,N_14028,N_13844);
or U14281 (N_14281,N_13894,N_14030);
or U14282 (N_14282,N_13983,N_14144);
xor U14283 (N_14283,N_14201,N_14234);
nor U14284 (N_14284,N_13855,N_14243);
or U14285 (N_14285,N_14180,N_13766);
xor U14286 (N_14286,N_14052,N_14131);
nor U14287 (N_14287,N_13534,N_13895);
nand U14288 (N_14288,N_13554,N_13613);
or U14289 (N_14289,N_14018,N_13541);
or U14290 (N_14290,N_14040,N_13509);
and U14291 (N_14291,N_13910,N_14200);
and U14292 (N_14292,N_13614,N_14129);
nor U14293 (N_14293,N_13931,N_13581);
nand U14294 (N_14294,N_13909,N_13868);
nor U14295 (N_14295,N_13946,N_13740);
nor U14296 (N_14296,N_13815,N_14042);
or U14297 (N_14297,N_13628,N_14056);
and U14298 (N_14298,N_13750,N_13537);
and U14299 (N_14299,N_13713,N_14229);
or U14300 (N_14300,N_13543,N_13617);
and U14301 (N_14301,N_13912,N_13627);
nor U14302 (N_14302,N_14176,N_14013);
nor U14303 (N_14303,N_13712,N_14206);
nand U14304 (N_14304,N_14038,N_14133);
or U14305 (N_14305,N_13634,N_13589);
and U14306 (N_14306,N_14218,N_13755);
or U14307 (N_14307,N_13775,N_13745);
xnor U14308 (N_14308,N_13687,N_14202);
and U14309 (N_14309,N_13859,N_13579);
and U14310 (N_14310,N_14062,N_14241);
nor U14311 (N_14311,N_14105,N_13732);
xnor U14312 (N_14312,N_13697,N_13788);
and U14313 (N_14313,N_13676,N_13737);
xnor U14314 (N_14314,N_13677,N_13879);
nand U14315 (N_14315,N_13630,N_13695);
nand U14316 (N_14316,N_13952,N_14041);
nand U14317 (N_14317,N_13528,N_13647);
nor U14318 (N_14318,N_13922,N_13776);
or U14319 (N_14319,N_13520,N_14089);
nor U14320 (N_14320,N_14205,N_13757);
or U14321 (N_14321,N_13860,N_13516);
nor U14322 (N_14322,N_14107,N_13612);
or U14323 (N_14323,N_13526,N_13723);
or U14324 (N_14324,N_14068,N_13916);
and U14325 (N_14325,N_13730,N_13986);
nand U14326 (N_14326,N_13993,N_13684);
xnor U14327 (N_14327,N_13531,N_13831);
xnor U14328 (N_14328,N_14118,N_14172);
nor U14329 (N_14329,N_13587,N_13762);
and U14330 (N_14330,N_14183,N_14124);
nor U14331 (N_14331,N_14113,N_14177);
xor U14332 (N_14332,N_13575,N_14002);
or U14333 (N_14333,N_13768,N_14248);
or U14334 (N_14334,N_14071,N_13544);
and U14335 (N_14335,N_13556,N_13953);
xor U14336 (N_14336,N_13877,N_13600);
nor U14337 (N_14337,N_14184,N_14021);
nand U14338 (N_14338,N_13738,N_13871);
and U14339 (N_14339,N_14209,N_13756);
nand U14340 (N_14340,N_13535,N_14193);
nand U14341 (N_14341,N_13662,N_13830);
nor U14342 (N_14342,N_13705,N_13974);
or U14343 (N_14343,N_13838,N_14009);
nor U14344 (N_14344,N_13563,N_13812);
nand U14345 (N_14345,N_14165,N_14233);
or U14346 (N_14346,N_14019,N_13959);
nor U14347 (N_14347,N_13521,N_14125);
nand U14348 (N_14348,N_14099,N_13893);
nor U14349 (N_14349,N_13794,N_13739);
or U14350 (N_14350,N_13972,N_13801);
nor U14351 (N_14351,N_13661,N_14049);
or U14352 (N_14352,N_14091,N_14120);
nor U14353 (N_14353,N_13821,N_13558);
nor U14354 (N_14354,N_13674,N_13511);
and U14355 (N_14355,N_13948,N_13876);
or U14356 (N_14356,N_13551,N_13637);
or U14357 (N_14357,N_13817,N_14236);
nand U14358 (N_14358,N_13787,N_13584);
nand U14359 (N_14359,N_13593,N_13779);
and U14360 (N_14360,N_13803,N_14197);
and U14361 (N_14361,N_13994,N_13660);
or U14362 (N_14362,N_14235,N_13790);
nor U14363 (N_14363,N_14054,N_13696);
and U14364 (N_14364,N_13670,N_14242);
and U14365 (N_14365,N_13685,N_14083);
nand U14366 (N_14366,N_13666,N_13865);
or U14367 (N_14367,N_14142,N_13678);
and U14368 (N_14368,N_14210,N_13915);
nor U14369 (N_14369,N_13576,N_14065);
or U14370 (N_14370,N_14214,N_13845);
nand U14371 (N_14371,N_13564,N_13566);
nand U14372 (N_14372,N_13623,N_14121);
and U14373 (N_14373,N_14001,N_13763);
and U14374 (N_14374,N_13769,N_13512);
nand U14375 (N_14375,N_13650,N_14152);
nand U14376 (N_14376,N_14198,N_14156);
xor U14377 (N_14377,N_13805,N_13610);
and U14378 (N_14378,N_14104,N_14066);
nand U14379 (N_14379,N_14162,N_13914);
nor U14380 (N_14380,N_14194,N_13691);
nor U14381 (N_14381,N_13924,N_13847);
nor U14382 (N_14382,N_13846,N_14145);
or U14383 (N_14383,N_13832,N_13829);
and U14384 (N_14384,N_13795,N_14084);
nor U14385 (N_14385,N_13574,N_13588);
nor U14386 (N_14386,N_13663,N_13827);
or U14387 (N_14387,N_13622,N_14005);
nor U14388 (N_14388,N_14207,N_14217);
or U14389 (N_14389,N_14102,N_14050);
nor U14390 (N_14390,N_13645,N_13773);
nand U14391 (N_14391,N_13913,N_14146);
or U14392 (N_14392,N_14239,N_13873);
nor U14393 (N_14393,N_13560,N_13780);
and U14394 (N_14394,N_13652,N_13605);
nor U14395 (N_14395,N_13679,N_14039);
or U14396 (N_14396,N_13602,N_14189);
nor U14397 (N_14397,N_13604,N_14059);
or U14398 (N_14398,N_13596,N_13771);
nor U14399 (N_14399,N_14226,N_14134);
nor U14400 (N_14400,N_14097,N_13896);
nor U14401 (N_14401,N_14025,N_13822);
and U14402 (N_14402,N_13802,N_14190);
and U14403 (N_14403,N_13930,N_13954);
or U14404 (N_14404,N_13571,N_13508);
or U14405 (N_14405,N_13862,N_14117);
or U14406 (N_14406,N_14088,N_14137);
or U14407 (N_14407,N_13716,N_13562);
nor U14408 (N_14408,N_13784,N_13742);
nor U14409 (N_14409,N_13651,N_14112);
or U14410 (N_14410,N_14157,N_14219);
or U14411 (N_14411,N_14114,N_14095);
nor U14412 (N_14412,N_14159,N_14203);
nand U14413 (N_14413,N_13599,N_13568);
and U14414 (N_14414,N_14060,N_14058);
nand U14415 (N_14415,N_13777,N_14244);
xor U14416 (N_14416,N_13759,N_13702);
or U14417 (N_14417,N_14181,N_13547);
and U14418 (N_14418,N_13843,N_13505);
and U14419 (N_14419,N_13704,N_13973);
and U14420 (N_14420,N_14169,N_13861);
nor U14421 (N_14421,N_13863,N_14222);
nand U14422 (N_14422,N_13741,N_13928);
and U14423 (N_14423,N_14188,N_14004);
nor U14424 (N_14424,N_14151,N_14034);
or U14425 (N_14425,N_13586,N_13884);
or U14426 (N_14426,N_13631,N_14149);
nand U14427 (N_14427,N_14237,N_13878);
nor U14428 (N_14428,N_14007,N_13782);
xnor U14429 (N_14429,N_13615,N_13731);
nor U14430 (N_14430,N_13626,N_14111);
or U14431 (N_14431,N_13849,N_13958);
or U14432 (N_14432,N_14153,N_13609);
and U14433 (N_14433,N_13724,N_13885);
and U14434 (N_14434,N_13992,N_14106);
nand U14435 (N_14435,N_14185,N_14215);
or U14436 (N_14436,N_13714,N_13866);
or U14437 (N_14437,N_14143,N_13937);
and U14438 (N_14438,N_13657,N_13743);
nor U14439 (N_14439,N_14094,N_13919);
nor U14440 (N_14440,N_13851,N_13950);
or U14441 (N_14441,N_13770,N_13525);
and U14442 (N_14442,N_13698,N_13681);
xnor U14443 (N_14443,N_13559,N_14128);
nand U14444 (N_14444,N_13979,N_13533);
nor U14445 (N_14445,N_14057,N_14110);
nand U14446 (N_14446,N_13529,N_13852);
nand U14447 (N_14447,N_14064,N_13826);
and U14448 (N_14448,N_13553,N_13625);
or U14449 (N_14449,N_14196,N_13778);
nand U14450 (N_14450,N_13754,N_13848);
xnor U14451 (N_14451,N_14182,N_13565);
xnor U14452 (N_14452,N_13920,N_14044);
nand U14453 (N_14453,N_13639,N_13791);
and U14454 (N_14454,N_14011,N_13585);
or U14455 (N_14455,N_13956,N_13985);
nand U14456 (N_14456,N_13809,N_13548);
or U14457 (N_14457,N_14171,N_13872);
and U14458 (N_14458,N_13841,N_13818);
xor U14459 (N_14459,N_13785,N_13897);
nor U14460 (N_14460,N_13601,N_13620);
nor U14461 (N_14461,N_13942,N_14070);
nor U14462 (N_14462,N_13898,N_13810);
xnor U14463 (N_14463,N_13889,N_14224);
xor U14464 (N_14464,N_13892,N_13598);
xnor U14465 (N_14465,N_13635,N_13975);
and U14466 (N_14466,N_13899,N_14126);
or U14467 (N_14467,N_13686,N_13706);
xor U14468 (N_14468,N_14090,N_13690);
nand U14469 (N_14469,N_13998,N_14220);
nor U14470 (N_14470,N_14053,N_13545);
nand U14471 (N_14471,N_13867,N_14199);
or U14472 (N_14472,N_13813,N_13798);
and U14473 (N_14473,N_13995,N_13514);
or U14474 (N_14474,N_14067,N_13887);
nor U14475 (N_14475,N_14173,N_13984);
or U14476 (N_14476,N_13804,N_13834);
or U14477 (N_14477,N_14026,N_14008);
nand U14478 (N_14478,N_13669,N_13675);
and U14479 (N_14479,N_13934,N_14170);
nand U14480 (N_14480,N_13774,N_13550);
nand U14481 (N_14481,N_13819,N_13567);
nand U14482 (N_14482,N_13792,N_13944);
nand U14483 (N_14483,N_13597,N_13940);
or U14484 (N_14484,N_13502,N_13659);
or U14485 (N_14485,N_13557,N_13753);
nand U14486 (N_14486,N_13951,N_14015);
and U14487 (N_14487,N_13546,N_14246);
and U14488 (N_14488,N_14216,N_14166);
nor U14489 (N_14489,N_13835,N_13881);
nand U14490 (N_14490,N_14247,N_13965);
and U14491 (N_14491,N_13970,N_13968);
or U14492 (N_14492,N_13747,N_13811);
and U14493 (N_14493,N_14204,N_13964);
nand U14494 (N_14494,N_13976,N_14098);
nor U14495 (N_14495,N_13619,N_14221);
nor U14496 (N_14496,N_14161,N_13720);
xor U14497 (N_14497,N_13522,N_14087);
and U14498 (N_14498,N_14081,N_13632);
xor U14499 (N_14499,N_14213,N_13901);
and U14500 (N_14500,N_13927,N_13891);
nand U14501 (N_14501,N_14072,N_14082);
or U14502 (N_14502,N_13523,N_13797);
nor U14503 (N_14503,N_14148,N_14154);
or U14504 (N_14504,N_13582,N_13590);
or U14505 (N_14505,N_14014,N_14155);
or U14506 (N_14506,N_13683,N_13905);
and U14507 (N_14507,N_13746,N_13971);
or U14508 (N_14508,N_13710,N_13786);
nor U14509 (N_14509,N_13515,N_14023);
nand U14510 (N_14510,N_13850,N_13733);
and U14511 (N_14511,N_13806,N_13987);
or U14512 (N_14512,N_14069,N_13886);
and U14513 (N_14513,N_13555,N_13978);
and U14514 (N_14514,N_13869,N_13990);
xor U14515 (N_14515,N_13783,N_13961);
or U14516 (N_14516,N_13820,N_13606);
xnor U14517 (N_14517,N_13772,N_14033);
or U14518 (N_14518,N_13751,N_13902);
or U14519 (N_14519,N_14024,N_13577);
nand U14520 (N_14520,N_14136,N_13808);
or U14521 (N_14521,N_14178,N_13699);
or U14522 (N_14522,N_13800,N_14035);
or U14523 (N_14523,N_13573,N_13680);
and U14524 (N_14524,N_14175,N_14115);
nand U14525 (N_14525,N_13689,N_14086);
nand U14526 (N_14526,N_13947,N_13646);
and U14527 (N_14527,N_14179,N_13962);
nor U14528 (N_14528,N_13727,N_13693);
nand U14529 (N_14529,N_14045,N_14016);
xnor U14530 (N_14530,N_13532,N_14240);
and U14531 (N_14531,N_13611,N_13967);
nor U14532 (N_14532,N_14211,N_13536);
or U14533 (N_14533,N_13977,N_13949);
nor U14534 (N_14534,N_13833,N_14132);
nor U14535 (N_14535,N_13840,N_13856);
and U14536 (N_14536,N_13932,N_13616);
and U14537 (N_14537,N_13595,N_13688);
and U14538 (N_14538,N_14036,N_13510);
and U14539 (N_14539,N_13519,N_14075);
nand U14540 (N_14540,N_14076,N_13542);
and U14541 (N_14541,N_13874,N_13664);
nor U14542 (N_14542,N_13807,N_14073);
and U14543 (N_14543,N_14192,N_13752);
and U14544 (N_14544,N_14061,N_13933);
nand U14545 (N_14545,N_13980,N_14108);
and U14546 (N_14546,N_13816,N_14228);
nand U14547 (N_14547,N_13999,N_14051);
nand U14548 (N_14548,N_13667,N_14043);
and U14549 (N_14549,N_13578,N_13982);
or U14550 (N_14550,N_13507,N_13701);
nand U14551 (N_14551,N_14047,N_13991);
or U14552 (N_14552,N_14020,N_13672);
nor U14553 (N_14553,N_13648,N_13721);
and U14554 (N_14554,N_13709,N_13882);
or U14555 (N_14555,N_13858,N_13824);
nor U14556 (N_14556,N_14150,N_13883);
or U14557 (N_14557,N_14123,N_13842);
and U14558 (N_14558,N_14048,N_14245);
nand U14559 (N_14559,N_14225,N_13765);
or U14560 (N_14560,N_13517,N_14186);
nand U14561 (N_14561,N_13594,N_13825);
and U14562 (N_14562,N_14130,N_14006);
or U14563 (N_14563,N_14138,N_13649);
nor U14564 (N_14564,N_13789,N_13749);
nand U14565 (N_14565,N_13828,N_14230);
nor U14566 (N_14566,N_13767,N_13941);
and U14567 (N_14567,N_14022,N_13580);
nor U14568 (N_14568,N_14093,N_14096);
or U14569 (N_14569,N_14147,N_13569);
nor U14570 (N_14570,N_14141,N_13864);
nand U14571 (N_14571,N_13591,N_13506);
and U14572 (N_14572,N_13629,N_13908);
nand U14573 (N_14573,N_14092,N_14158);
and U14574 (N_14574,N_13641,N_13853);
nor U14575 (N_14575,N_14223,N_13764);
and U14576 (N_14576,N_13799,N_13854);
or U14577 (N_14577,N_13726,N_13539);
nand U14578 (N_14578,N_13839,N_14055);
or U14579 (N_14579,N_13708,N_14031);
or U14580 (N_14580,N_13640,N_13857);
and U14581 (N_14581,N_13633,N_13875);
xnor U14582 (N_14582,N_13607,N_14003);
nor U14583 (N_14583,N_14080,N_13658);
nand U14584 (N_14584,N_13711,N_14027);
or U14585 (N_14585,N_13707,N_13719);
nand U14586 (N_14586,N_13624,N_13638);
xnor U14587 (N_14587,N_14085,N_13503);
xnor U14588 (N_14588,N_13936,N_13880);
and U14589 (N_14589,N_14103,N_13728);
nand U14590 (N_14590,N_13981,N_13904);
nand U14591 (N_14591,N_14032,N_13945);
nor U14592 (N_14592,N_13552,N_13572);
or U14593 (N_14593,N_14238,N_14074);
nand U14594 (N_14594,N_13989,N_14168);
nor U14595 (N_14595,N_13900,N_13966);
or U14596 (N_14596,N_13781,N_13996);
or U14597 (N_14597,N_13925,N_14037);
or U14598 (N_14598,N_13668,N_14046);
nor U14599 (N_14599,N_14139,N_13654);
nand U14600 (N_14600,N_14212,N_13570);
or U14601 (N_14601,N_14010,N_13938);
nor U14602 (N_14602,N_13718,N_13673);
or U14603 (N_14603,N_13903,N_13935);
nand U14604 (N_14604,N_13735,N_13955);
nor U14605 (N_14605,N_13960,N_13963);
or U14606 (N_14606,N_13621,N_13549);
and U14607 (N_14607,N_13729,N_14063);
and U14608 (N_14608,N_14232,N_13988);
nor U14609 (N_14609,N_13682,N_14167);
and U14610 (N_14610,N_13918,N_13744);
and U14611 (N_14611,N_13715,N_13603);
and U14612 (N_14612,N_14140,N_13703);
nor U14613 (N_14613,N_13561,N_14122);
nand U14614 (N_14614,N_13618,N_14127);
or U14615 (N_14615,N_14012,N_13504);
xor U14616 (N_14616,N_14079,N_13907);
nor U14617 (N_14617,N_13917,N_13911);
or U14618 (N_14618,N_14249,N_13643);
and U14619 (N_14619,N_14109,N_13583);
nor U14620 (N_14620,N_13636,N_13608);
and U14621 (N_14621,N_13501,N_14163);
or U14622 (N_14622,N_14174,N_13592);
nand U14623 (N_14623,N_14191,N_13906);
nor U14624 (N_14624,N_13957,N_13926);
nand U14625 (N_14625,N_14223,N_13742);
nand U14626 (N_14626,N_13834,N_14208);
or U14627 (N_14627,N_14197,N_13808);
or U14628 (N_14628,N_13701,N_13578);
xnor U14629 (N_14629,N_14081,N_14071);
nand U14630 (N_14630,N_13804,N_13961);
and U14631 (N_14631,N_13839,N_13802);
or U14632 (N_14632,N_13953,N_14220);
nor U14633 (N_14633,N_13837,N_14170);
xor U14634 (N_14634,N_13589,N_13892);
nor U14635 (N_14635,N_13537,N_13969);
or U14636 (N_14636,N_14198,N_13950);
nor U14637 (N_14637,N_13792,N_13553);
or U14638 (N_14638,N_14077,N_13930);
and U14639 (N_14639,N_13952,N_13968);
or U14640 (N_14640,N_13917,N_13748);
nor U14641 (N_14641,N_13959,N_13719);
nor U14642 (N_14642,N_13879,N_13553);
and U14643 (N_14643,N_13758,N_13740);
nand U14644 (N_14644,N_13831,N_13839);
nand U14645 (N_14645,N_13955,N_13714);
or U14646 (N_14646,N_13597,N_14218);
and U14647 (N_14647,N_14097,N_14064);
or U14648 (N_14648,N_13673,N_13591);
nand U14649 (N_14649,N_13886,N_13904);
or U14650 (N_14650,N_14033,N_13807);
nor U14651 (N_14651,N_13850,N_13582);
or U14652 (N_14652,N_13640,N_14150);
xnor U14653 (N_14653,N_13948,N_14067);
nor U14654 (N_14654,N_13546,N_14115);
and U14655 (N_14655,N_14236,N_13695);
nand U14656 (N_14656,N_14217,N_13850);
nand U14657 (N_14657,N_13706,N_14153);
nand U14658 (N_14658,N_13955,N_13559);
xor U14659 (N_14659,N_13876,N_13875);
xor U14660 (N_14660,N_13902,N_14162);
nor U14661 (N_14661,N_13614,N_14077);
and U14662 (N_14662,N_14116,N_13721);
and U14663 (N_14663,N_13798,N_13705);
and U14664 (N_14664,N_13598,N_13566);
nand U14665 (N_14665,N_13831,N_13621);
nor U14666 (N_14666,N_13671,N_13899);
xnor U14667 (N_14667,N_13536,N_13957);
or U14668 (N_14668,N_13639,N_14072);
and U14669 (N_14669,N_14076,N_13801);
nor U14670 (N_14670,N_13917,N_13582);
and U14671 (N_14671,N_13855,N_14056);
nor U14672 (N_14672,N_13720,N_13815);
nand U14673 (N_14673,N_14249,N_13963);
or U14674 (N_14674,N_14032,N_13760);
and U14675 (N_14675,N_14045,N_13615);
or U14676 (N_14676,N_14197,N_14184);
nor U14677 (N_14677,N_14113,N_13819);
nand U14678 (N_14678,N_14180,N_13948);
nand U14679 (N_14679,N_14118,N_14234);
nor U14680 (N_14680,N_13597,N_13933);
xnor U14681 (N_14681,N_13797,N_13783);
or U14682 (N_14682,N_13654,N_13892);
and U14683 (N_14683,N_13521,N_13700);
nor U14684 (N_14684,N_14076,N_13860);
nand U14685 (N_14685,N_13514,N_14207);
nand U14686 (N_14686,N_13815,N_14128);
or U14687 (N_14687,N_13698,N_13644);
nor U14688 (N_14688,N_13865,N_13609);
nor U14689 (N_14689,N_13929,N_13601);
or U14690 (N_14690,N_13936,N_13894);
and U14691 (N_14691,N_13548,N_14249);
nor U14692 (N_14692,N_14018,N_13558);
and U14693 (N_14693,N_13959,N_14077);
nor U14694 (N_14694,N_14089,N_13709);
nand U14695 (N_14695,N_14156,N_13601);
and U14696 (N_14696,N_13712,N_13511);
or U14697 (N_14697,N_13672,N_13858);
and U14698 (N_14698,N_13912,N_13670);
or U14699 (N_14699,N_13696,N_13931);
nor U14700 (N_14700,N_13621,N_14240);
and U14701 (N_14701,N_13884,N_13772);
and U14702 (N_14702,N_13982,N_14018);
nor U14703 (N_14703,N_14209,N_13518);
nand U14704 (N_14704,N_13616,N_14168);
and U14705 (N_14705,N_13566,N_13698);
nor U14706 (N_14706,N_13567,N_13505);
and U14707 (N_14707,N_13795,N_14176);
and U14708 (N_14708,N_14182,N_13870);
nand U14709 (N_14709,N_14147,N_13750);
and U14710 (N_14710,N_14207,N_14214);
nor U14711 (N_14711,N_13770,N_13626);
and U14712 (N_14712,N_13620,N_13822);
and U14713 (N_14713,N_13826,N_13516);
xor U14714 (N_14714,N_13906,N_13610);
nor U14715 (N_14715,N_13685,N_13908);
and U14716 (N_14716,N_13601,N_14035);
or U14717 (N_14717,N_13740,N_14073);
and U14718 (N_14718,N_13905,N_14097);
nor U14719 (N_14719,N_13699,N_13655);
and U14720 (N_14720,N_13953,N_13628);
or U14721 (N_14721,N_13789,N_13842);
xnor U14722 (N_14722,N_13890,N_13563);
and U14723 (N_14723,N_14226,N_13628);
nor U14724 (N_14724,N_13617,N_13667);
and U14725 (N_14725,N_13705,N_13657);
or U14726 (N_14726,N_14146,N_14016);
nand U14727 (N_14727,N_13568,N_13727);
nor U14728 (N_14728,N_13687,N_14230);
or U14729 (N_14729,N_14086,N_13954);
nand U14730 (N_14730,N_14240,N_13948);
and U14731 (N_14731,N_14151,N_14088);
or U14732 (N_14732,N_14068,N_14165);
nand U14733 (N_14733,N_13707,N_13655);
or U14734 (N_14734,N_14134,N_13897);
nand U14735 (N_14735,N_13675,N_13994);
nor U14736 (N_14736,N_13991,N_13597);
or U14737 (N_14737,N_13761,N_13678);
xor U14738 (N_14738,N_13680,N_13525);
nor U14739 (N_14739,N_13716,N_13798);
nand U14740 (N_14740,N_14063,N_14135);
nand U14741 (N_14741,N_13982,N_13597);
nor U14742 (N_14742,N_14106,N_14002);
or U14743 (N_14743,N_13656,N_14002);
or U14744 (N_14744,N_13683,N_13654);
and U14745 (N_14745,N_14074,N_13792);
and U14746 (N_14746,N_14249,N_13603);
nand U14747 (N_14747,N_14156,N_13675);
xnor U14748 (N_14748,N_14059,N_13649);
and U14749 (N_14749,N_14174,N_14204);
nand U14750 (N_14750,N_13667,N_14084);
and U14751 (N_14751,N_14095,N_13640);
or U14752 (N_14752,N_13801,N_13900);
nor U14753 (N_14753,N_14201,N_13709);
nand U14754 (N_14754,N_13655,N_14071);
xnor U14755 (N_14755,N_14107,N_13735);
nand U14756 (N_14756,N_14101,N_13725);
nor U14757 (N_14757,N_13578,N_14117);
nor U14758 (N_14758,N_13808,N_13673);
nand U14759 (N_14759,N_14079,N_13625);
nand U14760 (N_14760,N_13564,N_13803);
nor U14761 (N_14761,N_13608,N_13570);
nor U14762 (N_14762,N_14110,N_13820);
xor U14763 (N_14763,N_13937,N_14033);
or U14764 (N_14764,N_14105,N_14132);
nor U14765 (N_14765,N_13515,N_13544);
nor U14766 (N_14766,N_14014,N_14060);
xor U14767 (N_14767,N_14142,N_13648);
and U14768 (N_14768,N_13770,N_14146);
nand U14769 (N_14769,N_14123,N_13988);
nand U14770 (N_14770,N_13652,N_13969);
xnor U14771 (N_14771,N_14162,N_13898);
and U14772 (N_14772,N_14243,N_14061);
or U14773 (N_14773,N_13868,N_13665);
and U14774 (N_14774,N_13930,N_13677);
nor U14775 (N_14775,N_13957,N_14227);
or U14776 (N_14776,N_13653,N_14047);
nor U14777 (N_14777,N_13988,N_14058);
or U14778 (N_14778,N_14011,N_13579);
nand U14779 (N_14779,N_13798,N_14080);
nand U14780 (N_14780,N_13638,N_13505);
or U14781 (N_14781,N_13913,N_14164);
and U14782 (N_14782,N_13519,N_14004);
and U14783 (N_14783,N_13708,N_13724);
nand U14784 (N_14784,N_13555,N_13564);
or U14785 (N_14785,N_13674,N_13690);
or U14786 (N_14786,N_13739,N_13534);
and U14787 (N_14787,N_13527,N_14122);
and U14788 (N_14788,N_13831,N_13906);
nor U14789 (N_14789,N_13945,N_13703);
nand U14790 (N_14790,N_14071,N_13773);
or U14791 (N_14791,N_14060,N_13763);
or U14792 (N_14792,N_14185,N_13713);
or U14793 (N_14793,N_14062,N_13757);
and U14794 (N_14794,N_13922,N_13989);
nand U14795 (N_14795,N_14042,N_14047);
nand U14796 (N_14796,N_14213,N_14176);
and U14797 (N_14797,N_14231,N_14161);
nor U14798 (N_14798,N_13761,N_13939);
and U14799 (N_14799,N_13878,N_13900);
nand U14800 (N_14800,N_13661,N_14213);
and U14801 (N_14801,N_13671,N_13517);
xnor U14802 (N_14802,N_13812,N_13707);
nand U14803 (N_14803,N_13672,N_13675);
nand U14804 (N_14804,N_13727,N_13922);
and U14805 (N_14805,N_13731,N_13694);
xnor U14806 (N_14806,N_13556,N_14016);
nand U14807 (N_14807,N_13564,N_14101);
or U14808 (N_14808,N_13849,N_14090);
nor U14809 (N_14809,N_14176,N_13766);
and U14810 (N_14810,N_14098,N_13955);
xor U14811 (N_14811,N_14097,N_14200);
and U14812 (N_14812,N_14249,N_14172);
nor U14813 (N_14813,N_14187,N_13958);
and U14814 (N_14814,N_13939,N_13724);
nand U14815 (N_14815,N_13691,N_14005);
nor U14816 (N_14816,N_13683,N_14173);
nand U14817 (N_14817,N_13554,N_14177);
xor U14818 (N_14818,N_13504,N_13724);
nor U14819 (N_14819,N_13587,N_13690);
nor U14820 (N_14820,N_13837,N_13616);
xor U14821 (N_14821,N_13551,N_13662);
or U14822 (N_14822,N_13513,N_13865);
nand U14823 (N_14823,N_13983,N_13837);
nand U14824 (N_14824,N_14165,N_14196);
nand U14825 (N_14825,N_14220,N_13542);
nor U14826 (N_14826,N_14171,N_13919);
or U14827 (N_14827,N_13665,N_14119);
nand U14828 (N_14828,N_13727,N_13882);
nor U14829 (N_14829,N_14121,N_13605);
and U14830 (N_14830,N_14139,N_13868);
nor U14831 (N_14831,N_14211,N_13998);
xnor U14832 (N_14832,N_13937,N_13908);
nor U14833 (N_14833,N_13724,N_13508);
nor U14834 (N_14834,N_13639,N_13815);
or U14835 (N_14835,N_14047,N_14241);
or U14836 (N_14836,N_13707,N_13511);
nand U14837 (N_14837,N_13517,N_13944);
nand U14838 (N_14838,N_13704,N_13934);
and U14839 (N_14839,N_13768,N_13886);
nand U14840 (N_14840,N_13996,N_14093);
xor U14841 (N_14841,N_13664,N_13502);
xnor U14842 (N_14842,N_13921,N_13815);
or U14843 (N_14843,N_14154,N_14089);
or U14844 (N_14844,N_13593,N_13575);
xnor U14845 (N_14845,N_14103,N_13670);
or U14846 (N_14846,N_14218,N_13765);
nor U14847 (N_14847,N_14131,N_13732);
nor U14848 (N_14848,N_14052,N_14072);
or U14849 (N_14849,N_14216,N_13526);
nand U14850 (N_14850,N_14091,N_14147);
or U14851 (N_14851,N_13767,N_13769);
and U14852 (N_14852,N_14229,N_13704);
or U14853 (N_14853,N_14193,N_14109);
nand U14854 (N_14854,N_14199,N_14038);
xnor U14855 (N_14855,N_14170,N_13908);
and U14856 (N_14856,N_14030,N_13535);
and U14857 (N_14857,N_14091,N_14248);
nor U14858 (N_14858,N_13532,N_13919);
or U14859 (N_14859,N_13545,N_13510);
or U14860 (N_14860,N_14225,N_13720);
or U14861 (N_14861,N_14052,N_13538);
nor U14862 (N_14862,N_14015,N_14032);
or U14863 (N_14863,N_14140,N_13993);
and U14864 (N_14864,N_13525,N_14011);
and U14865 (N_14865,N_13896,N_13925);
and U14866 (N_14866,N_13697,N_14003);
or U14867 (N_14867,N_13960,N_14243);
and U14868 (N_14868,N_13804,N_14143);
or U14869 (N_14869,N_14088,N_13976);
or U14870 (N_14870,N_14176,N_13636);
and U14871 (N_14871,N_13614,N_14063);
nor U14872 (N_14872,N_13795,N_13700);
and U14873 (N_14873,N_13586,N_13956);
or U14874 (N_14874,N_14142,N_13915);
and U14875 (N_14875,N_13691,N_13961);
and U14876 (N_14876,N_13630,N_13919);
nor U14877 (N_14877,N_13819,N_13964);
and U14878 (N_14878,N_13983,N_13635);
xnor U14879 (N_14879,N_13795,N_13647);
nor U14880 (N_14880,N_13943,N_13630);
and U14881 (N_14881,N_13653,N_14082);
nand U14882 (N_14882,N_14096,N_13985);
or U14883 (N_14883,N_13786,N_14000);
or U14884 (N_14884,N_14244,N_13845);
nand U14885 (N_14885,N_14180,N_14091);
and U14886 (N_14886,N_13825,N_13808);
nand U14887 (N_14887,N_13682,N_13964);
nor U14888 (N_14888,N_13565,N_13655);
and U14889 (N_14889,N_14146,N_13537);
nor U14890 (N_14890,N_13964,N_13667);
nand U14891 (N_14891,N_14217,N_13649);
or U14892 (N_14892,N_13873,N_13896);
xnor U14893 (N_14893,N_14200,N_13538);
and U14894 (N_14894,N_14216,N_13826);
and U14895 (N_14895,N_13986,N_13770);
nor U14896 (N_14896,N_13861,N_13722);
or U14897 (N_14897,N_13681,N_14246);
or U14898 (N_14898,N_13540,N_14152);
and U14899 (N_14899,N_13589,N_13897);
nand U14900 (N_14900,N_14152,N_13564);
nand U14901 (N_14901,N_13997,N_14050);
nor U14902 (N_14902,N_14118,N_13918);
nor U14903 (N_14903,N_13837,N_14246);
and U14904 (N_14904,N_13979,N_14205);
nor U14905 (N_14905,N_14091,N_14078);
xnor U14906 (N_14906,N_14160,N_13519);
xnor U14907 (N_14907,N_13726,N_14195);
or U14908 (N_14908,N_14051,N_13837);
and U14909 (N_14909,N_13651,N_13658);
xnor U14910 (N_14910,N_13569,N_14235);
and U14911 (N_14911,N_13926,N_13989);
or U14912 (N_14912,N_13824,N_13594);
nand U14913 (N_14913,N_13764,N_13716);
or U14914 (N_14914,N_13568,N_14146);
xnor U14915 (N_14915,N_13701,N_13685);
xnor U14916 (N_14916,N_14144,N_14112);
nor U14917 (N_14917,N_13895,N_13706);
nand U14918 (N_14918,N_14169,N_13573);
or U14919 (N_14919,N_14055,N_13628);
nand U14920 (N_14920,N_13996,N_13901);
nand U14921 (N_14921,N_13628,N_13832);
nor U14922 (N_14922,N_14043,N_14222);
nor U14923 (N_14923,N_13866,N_13667);
and U14924 (N_14924,N_13899,N_14105);
or U14925 (N_14925,N_13567,N_13890);
or U14926 (N_14926,N_13926,N_13811);
or U14927 (N_14927,N_14106,N_13528);
nor U14928 (N_14928,N_13969,N_14025);
or U14929 (N_14929,N_13784,N_14013);
or U14930 (N_14930,N_13818,N_13669);
or U14931 (N_14931,N_13564,N_13510);
nand U14932 (N_14932,N_13581,N_13598);
nand U14933 (N_14933,N_13512,N_14227);
nor U14934 (N_14934,N_13748,N_13878);
or U14935 (N_14935,N_13713,N_13725);
nand U14936 (N_14936,N_13872,N_14230);
and U14937 (N_14937,N_13971,N_13613);
or U14938 (N_14938,N_13539,N_14189);
xnor U14939 (N_14939,N_13947,N_13585);
and U14940 (N_14940,N_13760,N_13748);
and U14941 (N_14941,N_13653,N_14158);
and U14942 (N_14942,N_13657,N_13545);
and U14943 (N_14943,N_13717,N_13554);
nand U14944 (N_14944,N_14084,N_13549);
nand U14945 (N_14945,N_13670,N_13856);
xor U14946 (N_14946,N_14118,N_13810);
xor U14947 (N_14947,N_14107,N_13707);
nand U14948 (N_14948,N_13546,N_13924);
nand U14949 (N_14949,N_14124,N_13932);
nor U14950 (N_14950,N_13910,N_14041);
or U14951 (N_14951,N_13850,N_13588);
and U14952 (N_14952,N_14077,N_13531);
nand U14953 (N_14953,N_13831,N_13979);
and U14954 (N_14954,N_13650,N_13663);
and U14955 (N_14955,N_13882,N_13513);
or U14956 (N_14956,N_14241,N_13875);
and U14957 (N_14957,N_14241,N_13640);
or U14958 (N_14958,N_13964,N_13506);
nand U14959 (N_14959,N_13817,N_13956);
xnor U14960 (N_14960,N_13902,N_14176);
nand U14961 (N_14961,N_13515,N_13530);
nor U14962 (N_14962,N_14051,N_14195);
or U14963 (N_14963,N_14180,N_13585);
or U14964 (N_14964,N_13660,N_13903);
nand U14965 (N_14965,N_13527,N_14224);
and U14966 (N_14966,N_14097,N_14101);
or U14967 (N_14967,N_13980,N_14226);
nor U14968 (N_14968,N_13582,N_13545);
or U14969 (N_14969,N_14105,N_13854);
nand U14970 (N_14970,N_14201,N_13919);
or U14971 (N_14971,N_14167,N_13822);
and U14972 (N_14972,N_13832,N_14017);
nor U14973 (N_14973,N_13643,N_13639);
nor U14974 (N_14974,N_13671,N_13761);
and U14975 (N_14975,N_14156,N_14022);
nand U14976 (N_14976,N_13694,N_13505);
or U14977 (N_14977,N_13614,N_13723);
nor U14978 (N_14978,N_14197,N_13707);
nor U14979 (N_14979,N_13894,N_14171);
nor U14980 (N_14980,N_14154,N_13634);
nand U14981 (N_14981,N_13714,N_13689);
xnor U14982 (N_14982,N_13623,N_14059);
nand U14983 (N_14983,N_14029,N_13934);
and U14984 (N_14984,N_13979,N_13885);
and U14985 (N_14985,N_13808,N_13562);
and U14986 (N_14986,N_13970,N_13886);
or U14987 (N_14987,N_13688,N_13887);
nor U14988 (N_14988,N_13923,N_13772);
nor U14989 (N_14989,N_13680,N_13605);
xnor U14990 (N_14990,N_13668,N_13684);
or U14991 (N_14991,N_13533,N_14104);
or U14992 (N_14992,N_14076,N_13773);
or U14993 (N_14993,N_13706,N_14207);
or U14994 (N_14994,N_14161,N_13708);
or U14995 (N_14995,N_13768,N_13942);
xor U14996 (N_14996,N_13713,N_13926);
and U14997 (N_14997,N_14099,N_13698);
or U14998 (N_14998,N_13723,N_13696);
nand U14999 (N_14999,N_13897,N_13817);
nand UO_0 (O_0,N_14560,N_14407);
and UO_1 (O_1,N_14441,N_14589);
or UO_2 (O_2,N_14490,N_14878);
or UO_3 (O_3,N_14499,N_14507);
and UO_4 (O_4,N_14926,N_14682);
nor UO_5 (O_5,N_14669,N_14437);
xor UO_6 (O_6,N_14973,N_14330);
or UO_7 (O_7,N_14621,N_14559);
and UO_8 (O_8,N_14769,N_14617);
nand UO_9 (O_9,N_14797,N_14486);
nand UO_10 (O_10,N_14664,N_14981);
nor UO_11 (O_11,N_14483,N_14562);
nor UO_12 (O_12,N_14366,N_14281);
nor UO_13 (O_13,N_14752,N_14896);
nor UO_14 (O_14,N_14556,N_14945);
nor UO_15 (O_15,N_14683,N_14755);
nor UO_16 (O_16,N_14550,N_14667);
nand UO_17 (O_17,N_14909,N_14553);
nand UO_18 (O_18,N_14999,N_14466);
nand UO_19 (O_19,N_14271,N_14604);
nor UO_20 (O_20,N_14998,N_14933);
nand UO_21 (O_21,N_14855,N_14842);
nor UO_22 (O_22,N_14343,N_14458);
or UO_23 (O_23,N_14648,N_14658);
and UO_24 (O_24,N_14767,N_14943);
and UO_25 (O_25,N_14401,N_14868);
nand UO_26 (O_26,N_14696,N_14530);
nand UO_27 (O_27,N_14914,N_14512);
nor UO_28 (O_28,N_14776,N_14285);
nand UO_29 (O_29,N_14390,N_14480);
nor UO_30 (O_30,N_14850,N_14256);
and UO_31 (O_31,N_14418,N_14760);
nand UO_32 (O_32,N_14375,N_14740);
xor UO_33 (O_33,N_14870,N_14582);
nand UO_34 (O_34,N_14475,N_14558);
and UO_35 (O_35,N_14781,N_14662);
or UO_36 (O_36,N_14303,N_14893);
xor UO_37 (O_37,N_14978,N_14277);
and UO_38 (O_38,N_14810,N_14779);
nor UO_39 (O_39,N_14503,N_14546);
or UO_40 (O_40,N_14424,N_14554);
nor UO_41 (O_41,N_14257,N_14615);
and UO_42 (O_42,N_14987,N_14997);
nand UO_43 (O_43,N_14660,N_14629);
and UO_44 (O_44,N_14304,N_14314);
and UO_45 (O_45,N_14880,N_14731);
nor UO_46 (O_46,N_14516,N_14548);
nand UO_47 (O_47,N_14789,N_14610);
and UO_48 (O_48,N_14645,N_14625);
nand UO_49 (O_49,N_14495,N_14885);
nor UO_50 (O_50,N_14489,N_14672);
xor UO_51 (O_51,N_14439,N_14848);
or UO_52 (O_52,N_14677,N_14812);
and UO_53 (O_53,N_14688,N_14864);
and UO_54 (O_54,N_14768,N_14491);
and UO_55 (O_55,N_14649,N_14345);
nand UO_56 (O_56,N_14590,N_14942);
and UO_57 (O_57,N_14921,N_14989);
nand UO_58 (O_58,N_14592,N_14340);
nor UO_59 (O_59,N_14720,N_14828);
nand UO_60 (O_60,N_14958,N_14521);
nand UO_61 (O_61,N_14829,N_14421);
xnor UO_62 (O_62,N_14598,N_14840);
or UO_63 (O_63,N_14965,N_14944);
nand UO_64 (O_64,N_14392,N_14427);
nand UO_65 (O_65,N_14352,N_14759);
nand UO_66 (O_66,N_14936,N_14849);
xor UO_67 (O_67,N_14920,N_14860);
and UO_68 (O_68,N_14659,N_14370);
and UO_69 (O_69,N_14750,N_14467);
nor UO_70 (O_70,N_14518,N_14739);
and UO_71 (O_71,N_14916,N_14524);
or UO_72 (O_72,N_14297,N_14723);
nand UO_73 (O_73,N_14357,N_14784);
or UO_74 (O_74,N_14379,N_14798);
or UO_75 (O_75,N_14317,N_14552);
and UO_76 (O_76,N_14320,N_14957);
nor UO_77 (O_77,N_14968,N_14890);
nand UO_78 (O_78,N_14875,N_14959);
and UO_79 (O_79,N_14974,N_14572);
nand UO_80 (O_80,N_14701,N_14538);
nand UO_81 (O_81,N_14396,N_14844);
or UO_82 (O_82,N_14627,N_14416);
xnor UO_83 (O_83,N_14874,N_14377);
and UO_84 (O_84,N_14535,N_14811);
nor UO_85 (O_85,N_14851,N_14924);
nand UO_86 (O_86,N_14476,N_14895);
nor UO_87 (O_87,N_14286,N_14459);
or UO_88 (O_88,N_14255,N_14887);
nor UO_89 (O_89,N_14673,N_14346);
or UO_90 (O_90,N_14472,N_14670);
nor UO_91 (O_91,N_14671,N_14732);
and UO_92 (O_92,N_14948,N_14821);
nor UO_93 (O_93,N_14643,N_14708);
nor UO_94 (O_94,N_14818,N_14384);
nand UO_95 (O_95,N_14774,N_14497);
nand UO_96 (O_96,N_14743,N_14704);
and UO_97 (O_97,N_14910,N_14272);
nor UO_98 (O_98,N_14742,N_14832);
nor UO_99 (O_99,N_14907,N_14908);
or UO_100 (O_100,N_14536,N_14730);
and UO_101 (O_101,N_14254,N_14638);
or UO_102 (O_102,N_14680,N_14498);
or UO_103 (O_103,N_14494,N_14517);
nand UO_104 (O_104,N_14325,N_14266);
and UO_105 (O_105,N_14533,N_14406);
nor UO_106 (O_106,N_14904,N_14350);
nand UO_107 (O_107,N_14527,N_14251);
nor UO_108 (O_108,N_14534,N_14465);
nor UO_109 (O_109,N_14292,N_14700);
nand UO_110 (O_110,N_14446,N_14865);
nand UO_111 (O_111,N_14367,N_14316);
nand UO_112 (O_112,N_14337,N_14970);
or UO_113 (O_113,N_14381,N_14616);
or UO_114 (O_114,N_14531,N_14508);
and UO_115 (O_115,N_14461,N_14854);
nor UO_116 (O_116,N_14596,N_14445);
and UO_117 (O_117,N_14310,N_14770);
or UO_118 (O_118,N_14478,N_14713);
and UO_119 (O_119,N_14744,N_14448);
nand UO_120 (O_120,N_14425,N_14541);
or UO_121 (O_121,N_14915,N_14695);
nand UO_122 (O_122,N_14994,N_14819);
or UO_123 (O_123,N_14585,N_14358);
nor UO_124 (O_124,N_14996,N_14253);
xnor UO_125 (O_125,N_14455,N_14258);
or UO_126 (O_126,N_14555,N_14603);
nor UO_127 (O_127,N_14709,N_14333);
nor UO_128 (O_128,N_14252,N_14565);
or UO_129 (O_129,N_14631,N_14298);
or UO_130 (O_130,N_14332,N_14485);
and UO_131 (O_131,N_14815,N_14846);
or UO_132 (O_132,N_14576,N_14463);
xor UO_133 (O_133,N_14793,N_14632);
nand UO_134 (O_134,N_14540,N_14727);
nor UO_135 (O_135,N_14808,N_14542);
or UO_136 (O_136,N_14305,N_14288);
nor UO_137 (O_137,N_14468,N_14872);
xor UO_138 (O_138,N_14983,N_14666);
and UO_139 (O_139,N_14619,N_14452);
and UO_140 (O_140,N_14827,N_14278);
and UO_141 (O_141,N_14510,N_14597);
and UO_142 (O_142,N_14280,N_14609);
xor UO_143 (O_143,N_14279,N_14741);
nor UO_144 (O_144,N_14993,N_14359);
nand UO_145 (O_145,N_14805,N_14397);
nor UO_146 (O_146,N_14873,N_14923);
and UO_147 (O_147,N_14500,N_14734);
nand UO_148 (O_148,N_14869,N_14967);
xor UO_149 (O_149,N_14665,N_14436);
nor UO_150 (O_150,N_14313,N_14833);
nand UO_151 (O_151,N_14733,N_14593);
xor UO_152 (O_152,N_14365,N_14567);
nand UO_153 (O_153,N_14566,N_14826);
nor UO_154 (O_154,N_14698,N_14917);
nor UO_155 (O_155,N_14702,N_14426);
nand UO_156 (O_156,N_14898,N_14900);
nor UO_157 (O_157,N_14939,N_14949);
or UO_158 (O_158,N_14646,N_14434);
or UO_159 (O_159,N_14640,N_14913);
nand UO_160 (O_160,N_14675,N_14299);
and UO_161 (O_161,N_14432,N_14492);
or UO_162 (O_162,N_14644,N_14382);
or UO_163 (O_163,N_14804,N_14290);
nand UO_164 (O_164,N_14349,N_14372);
nand UO_165 (O_165,N_14988,N_14449);
nor UO_166 (O_166,N_14543,N_14716);
nor UO_167 (O_167,N_14816,N_14883);
and UO_168 (O_168,N_14663,N_14888);
nor UO_169 (O_169,N_14712,N_14335);
nor UO_170 (O_170,N_14626,N_14311);
nor UO_171 (O_171,N_14674,N_14766);
and UO_172 (O_172,N_14570,N_14886);
nor UO_173 (O_173,N_14462,N_14928);
nand UO_174 (O_174,N_14790,N_14302);
and UO_175 (O_175,N_14661,N_14636);
or UO_176 (O_176,N_14338,N_14308);
nand UO_177 (O_177,N_14746,N_14353);
or UO_178 (O_178,N_14685,N_14364);
and UO_179 (O_179,N_14705,N_14971);
and UO_180 (O_180,N_14783,N_14327);
nor UO_181 (O_181,N_14919,N_14802);
xor UO_182 (O_182,N_14391,N_14841);
or UO_183 (O_183,N_14795,N_14504);
nor UO_184 (O_184,N_14788,N_14265);
or UO_185 (O_185,N_14532,N_14642);
nand UO_186 (O_186,N_14903,N_14754);
nand UO_187 (O_187,N_14947,N_14514);
nand UO_188 (O_188,N_14830,N_14451);
and UO_189 (O_189,N_14726,N_14259);
or UO_190 (O_190,N_14992,N_14929);
nor UO_191 (O_191,N_14980,N_14502);
nor UO_192 (O_192,N_14778,N_14454);
nand UO_193 (O_193,N_14889,N_14506);
nor UO_194 (O_194,N_14599,N_14402);
nand UO_195 (O_195,N_14487,N_14505);
or UO_196 (O_196,N_14395,N_14263);
or UO_197 (O_197,N_14691,N_14655);
xnor UO_198 (O_198,N_14956,N_14736);
nor UO_199 (O_199,N_14293,N_14689);
nand UO_200 (O_200,N_14569,N_14405);
xnor UO_201 (O_201,N_14267,N_14547);
nor UO_202 (O_202,N_14474,N_14803);
xor UO_203 (O_203,N_14300,N_14728);
nand UO_204 (O_204,N_14457,N_14719);
xor UO_205 (O_205,N_14836,N_14417);
and UO_206 (O_206,N_14551,N_14525);
nor UO_207 (O_207,N_14264,N_14481);
xor UO_208 (O_208,N_14792,N_14964);
nor UO_209 (O_209,N_14261,N_14544);
nor UO_210 (O_210,N_14668,N_14694);
or UO_211 (O_211,N_14412,N_14686);
or UO_212 (O_212,N_14336,N_14955);
nor UO_213 (O_213,N_14322,N_14523);
nor UO_214 (O_214,N_14715,N_14801);
or UO_215 (O_215,N_14982,N_14820);
or UO_216 (O_216,N_14953,N_14881);
or UO_217 (O_217,N_14678,N_14753);
nor UO_218 (O_218,N_14932,N_14876);
and UO_219 (O_219,N_14930,N_14399);
or UO_220 (O_220,N_14488,N_14845);
nand UO_221 (O_221,N_14780,N_14371);
and UO_222 (O_222,N_14834,N_14513);
nor UO_223 (O_223,N_14564,N_14545);
nor UO_224 (O_224,N_14413,N_14977);
and UO_225 (O_225,N_14952,N_14435);
and UO_226 (O_226,N_14785,N_14289);
nand UO_227 (O_227,N_14250,N_14937);
and UO_228 (O_228,N_14813,N_14351);
nor UO_229 (O_229,N_14976,N_14654);
nor UO_230 (O_230,N_14356,N_14653);
and UO_231 (O_231,N_14931,N_14641);
and UO_232 (O_232,N_14707,N_14511);
nor UO_233 (O_233,N_14270,N_14990);
or UO_234 (O_234,N_14422,N_14637);
xnor UO_235 (O_235,N_14268,N_14986);
xnor UO_236 (O_236,N_14493,N_14925);
nand UO_237 (O_237,N_14318,N_14941);
xnor UO_238 (O_238,N_14339,N_14706);
or UO_239 (O_239,N_14954,N_14823);
nand UO_240 (O_240,N_14773,N_14331);
or UO_241 (O_241,N_14963,N_14612);
or UO_242 (O_242,N_14595,N_14312);
xnor UO_243 (O_243,N_14369,N_14853);
nor UO_244 (O_244,N_14765,N_14433);
or UO_245 (O_245,N_14938,N_14806);
or UO_246 (O_246,N_14835,N_14862);
nand UO_247 (O_247,N_14758,N_14423);
or UO_248 (O_248,N_14275,N_14717);
xor UO_249 (O_249,N_14960,N_14394);
xnor UO_250 (O_250,N_14577,N_14415);
and UO_251 (O_251,N_14972,N_14722);
nand UO_252 (O_252,N_14342,N_14579);
nand UO_253 (O_253,N_14838,N_14613);
nor UO_254 (O_254,N_14323,N_14867);
xnor UO_255 (O_255,N_14647,N_14630);
and UO_256 (O_256,N_14469,N_14796);
or UO_257 (O_257,N_14309,N_14962);
nand UO_258 (O_258,N_14568,N_14639);
nor UO_259 (O_259,N_14324,N_14484);
or UO_260 (O_260,N_14807,N_14341);
nand UO_261 (O_261,N_14347,N_14618);
nand UO_262 (O_262,N_14857,N_14456);
and UO_263 (O_263,N_14697,N_14496);
nand UO_264 (O_264,N_14620,N_14749);
nand UO_265 (O_265,N_14319,N_14825);
and UO_266 (O_266,N_14262,N_14573);
or UO_267 (O_267,N_14334,N_14703);
or UO_268 (O_268,N_14877,N_14561);
and UO_269 (O_269,N_14583,N_14306);
nor UO_270 (O_270,N_14471,N_14607);
xnor UO_271 (O_271,N_14772,N_14699);
or UO_272 (O_272,N_14526,N_14519);
nand UO_273 (O_273,N_14725,N_14969);
nand UO_274 (O_274,N_14651,N_14387);
and UO_275 (O_275,N_14847,N_14363);
or UO_276 (O_276,N_14283,N_14737);
nor UO_277 (O_277,N_14757,N_14622);
and UO_278 (O_278,N_14676,N_14563);
and UO_279 (O_279,N_14771,N_14906);
and UO_280 (O_280,N_14681,N_14419);
nand UO_281 (O_281,N_14315,N_14307);
and UO_282 (O_282,N_14373,N_14692);
or UO_283 (O_283,N_14403,N_14408);
or UO_284 (O_284,N_14539,N_14591);
or UO_285 (O_285,N_14411,N_14360);
nor UO_286 (O_286,N_14824,N_14839);
and UO_287 (O_287,N_14383,N_14440);
xnor UO_288 (O_288,N_14438,N_14354);
nor UO_289 (O_289,N_14374,N_14501);
and UO_290 (O_290,N_14652,N_14587);
nor UO_291 (O_291,N_14984,N_14473);
nor UO_292 (O_292,N_14444,N_14863);
and UO_293 (O_293,N_14748,N_14528);
xnor UO_294 (O_294,N_14326,N_14301);
nand UO_295 (O_295,N_14388,N_14782);
nor UO_296 (O_296,N_14884,N_14380);
xor UO_297 (O_297,N_14633,N_14775);
or UO_298 (O_298,N_14430,N_14282);
nand UO_299 (O_299,N_14410,N_14389);
nor UO_300 (O_300,N_14273,N_14656);
and UO_301 (O_301,N_14866,N_14764);
nor UO_302 (O_302,N_14328,N_14581);
xor UO_303 (O_303,N_14761,N_14464);
nand UO_304 (O_304,N_14991,N_14745);
or UO_305 (O_305,N_14608,N_14393);
or UO_306 (O_306,N_14791,N_14871);
and UO_307 (O_307,N_14861,N_14276);
xnor UO_308 (O_308,N_14786,N_14602);
and UO_309 (O_309,N_14911,N_14584);
nand UO_310 (O_310,N_14940,N_14950);
or UO_311 (O_311,N_14344,N_14287);
nor UO_312 (O_312,N_14902,N_14571);
xnor UO_313 (O_313,N_14482,N_14409);
and UO_314 (O_314,N_14628,N_14296);
nor UO_315 (O_315,N_14578,N_14814);
or UO_316 (O_316,N_14624,N_14460);
nand UO_317 (O_317,N_14751,N_14594);
nand UO_318 (O_318,N_14574,N_14348);
or UO_319 (O_319,N_14549,N_14894);
nand UO_320 (O_320,N_14634,N_14817);
or UO_321 (O_321,N_14586,N_14800);
and UO_322 (O_322,N_14843,N_14918);
or UO_323 (O_323,N_14735,N_14657);
nand UO_324 (O_324,N_14291,N_14856);
nand UO_325 (O_325,N_14443,N_14450);
or UO_326 (O_326,N_14605,N_14718);
and UO_327 (O_327,N_14442,N_14927);
nand UO_328 (O_328,N_14635,N_14901);
nor UO_329 (O_329,N_14600,N_14479);
nand UO_330 (O_330,N_14477,N_14985);
xor UO_331 (O_331,N_14321,N_14922);
and UO_332 (O_332,N_14979,N_14274);
nor UO_333 (O_333,N_14724,N_14809);
nand UO_334 (O_334,N_14762,N_14269);
nor UO_335 (O_335,N_14738,N_14899);
and UO_336 (O_336,N_14368,N_14580);
or UO_337 (O_337,N_14515,N_14891);
nor UO_338 (O_338,N_14946,N_14687);
nand UO_339 (O_339,N_14859,N_14522);
nand UO_340 (O_340,N_14614,N_14611);
and UO_341 (O_341,N_14756,N_14376);
and UO_342 (O_342,N_14447,N_14588);
nor UO_343 (O_343,N_14747,N_14537);
or UO_344 (O_344,N_14879,N_14837);
nand UO_345 (O_345,N_14362,N_14710);
and UO_346 (O_346,N_14361,N_14431);
nand UO_347 (O_347,N_14852,N_14414);
nand UO_348 (O_348,N_14529,N_14693);
or UO_349 (O_349,N_14470,N_14453);
nand UO_350 (O_350,N_14404,N_14787);
nand UO_351 (O_351,N_14714,N_14799);
or UO_352 (O_352,N_14995,N_14295);
nor UO_353 (O_353,N_14386,N_14355);
or UO_354 (O_354,N_14329,N_14935);
and UO_355 (O_355,N_14260,N_14420);
and UO_356 (O_356,N_14882,N_14711);
or UO_357 (O_357,N_14294,N_14429);
nand UO_358 (O_358,N_14905,N_14575);
and UO_359 (O_359,N_14606,N_14794);
nor UO_360 (O_360,N_14601,N_14897);
nor UO_361 (O_361,N_14892,N_14858);
nand UO_362 (O_362,N_14690,N_14378);
or UO_363 (O_363,N_14509,N_14912);
nor UO_364 (O_364,N_14966,N_14961);
nor UO_365 (O_365,N_14428,N_14721);
xor UO_366 (O_366,N_14520,N_14729);
nand UO_367 (O_367,N_14650,N_14975);
nand UO_368 (O_368,N_14398,N_14934);
or UO_369 (O_369,N_14385,N_14951);
nand UO_370 (O_370,N_14684,N_14400);
or UO_371 (O_371,N_14763,N_14831);
and UO_372 (O_372,N_14822,N_14284);
and UO_373 (O_373,N_14679,N_14557);
nand UO_374 (O_374,N_14623,N_14777);
or UO_375 (O_375,N_14896,N_14707);
and UO_376 (O_376,N_14803,N_14603);
or UO_377 (O_377,N_14536,N_14784);
nand UO_378 (O_378,N_14603,N_14906);
xor UO_379 (O_379,N_14386,N_14535);
nand UO_380 (O_380,N_14571,N_14657);
nor UO_381 (O_381,N_14612,N_14793);
xor UO_382 (O_382,N_14383,N_14327);
or UO_383 (O_383,N_14935,N_14655);
xnor UO_384 (O_384,N_14935,N_14626);
and UO_385 (O_385,N_14403,N_14332);
nand UO_386 (O_386,N_14373,N_14847);
nand UO_387 (O_387,N_14277,N_14463);
or UO_388 (O_388,N_14277,N_14391);
nand UO_389 (O_389,N_14769,N_14588);
nand UO_390 (O_390,N_14253,N_14955);
nor UO_391 (O_391,N_14302,N_14284);
nand UO_392 (O_392,N_14478,N_14924);
nor UO_393 (O_393,N_14319,N_14878);
or UO_394 (O_394,N_14949,N_14579);
or UO_395 (O_395,N_14920,N_14397);
nand UO_396 (O_396,N_14302,N_14846);
nor UO_397 (O_397,N_14561,N_14317);
and UO_398 (O_398,N_14749,N_14929);
and UO_399 (O_399,N_14879,N_14398);
and UO_400 (O_400,N_14490,N_14975);
xnor UO_401 (O_401,N_14349,N_14600);
and UO_402 (O_402,N_14252,N_14503);
xor UO_403 (O_403,N_14581,N_14623);
nand UO_404 (O_404,N_14643,N_14479);
or UO_405 (O_405,N_14799,N_14881);
and UO_406 (O_406,N_14288,N_14419);
or UO_407 (O_407,N_14989,N_14696);
or UO_408 (O_408,N_14333,N_14523);
nand UO_409 (O_409,N_14503,N_14751);
and UO_410 (O_410,N_14898,N_14709);
and UO_411 (O_411,N_14557,N_14304);
nand UO_412 (O_412,N_14666,N_14378);
nand UO_413 (O_413,N_14730,N_14515);
or UO_414 (O_414,N_14933,N_14962);
or UO_415 (O_415,N_14664,N_14864);
nor UO_416 (O_416,N_14624,N_14951);
or UO_417 (O_417,N_14475,N_14796);
nor UO_418 (O_418,N_14777,N_14951);
nand UO_419 (O_419,N_14763,N_14876);
xor UO_420 (O_420,N_14824,N_14369);
nand UO_421 (O_421,N_14605,N_14608);
nor UO_422 (O_422,N_14362,N_14416);
and UO_423 (O_423,N_14379,N_14935);
or UO_424 (O_424,N_14776,N_14700);
and UO_425 (O_425,N_14257,N_14933);
or UO_426 (O_426,N_14865,N_14579);
nand UO_427 (O_427,N_14862,N_14387);
and UO_428 (O_428,N_14520,N_14720);
or UO_429 (O_429,N_14279,N_14314);
nor UO_430 (O_430,N_14919,N_14651);
or UO_431 (O_431,N_14662,N_14344);
xor UO_432 (O_432,N_14982,N_14552);
or UO_433 (O_433,N_14534,N_14520);
nor UO_434 (O_434,N_14389,N_14607);
nand UO_435 (O_435,N_14722,N_14536);
xor UO_436 (O_436,N_14995,N_14297);
and UO_437 (O_437,N_14609,N_14392);
and UO_438 (O_438,N_14497,N_14929);
nand UO_439 (O_439,N_14480,N_14628);
or UO_440 (O_440,N_14670,N_14353);
nand UO_441 (O_441,N_14365,N_14877);
nand UO_442 (O_442,N_14658,N_14764);
nor UO_443 (O_443,N_14752,N_14436);
nor UO_444 (O_444,N_14385,N_14312);
xnor UO_445 (O_445,N_14659,N_14340);
nor UO_446 (O_446,N_14837,N_14423);
and UO_447 (O_447,N_14898,N_14259);
or UO_448 (O_448,N_14673,N_14571);
xor UO_449 (O_449,N_14498,N_14684);
nor UO_450 (O_450,N_14760,N_14954);
or UO_451 (O_451,N_14578,N_14563);
or UO_452 (O_452,N_14459,N_14432);
nor UO_453 (O_453,N_14786,N_14361);
xor UO_454 (O_454,N_14361,N_14553);
and UO_455 (O_455,N_14878,N_14948);
or UO_456 (O_456,N_14428,N_14529);
nor UO_457 (O_457,N_14802,N_14822);
nand UO_458 (O_458,N_14454,N_14660);
nand UO_459 (O_459,N_14619,N_14649);
nand UO_460 (O_460,N_14393,N_14983);
and UO_461 (O_461,N_14651,N_14555);
nand UO_462 (O_462,N_14506,N_14499);
nor UO_463 (O_463,N_14869,N_14594);
or UO_464 (O_464,N_14419,N_14300);
and UO_465 (O_465,N_14877,N_14534);
or UO_466 (O_466,N_14982,N_14812);
and UO_467 (O_467,N_14406,N_14823);
and UO_468 (O_468,N_14480,N_14858);
or UO_469 (O_469,N_14791,N_14554);
nor UO_470 (O_470,N_14514,N_14594);
and UO_471 (O_471,N_14748,N_14851);
nor UO_472 (O_472,N_14484,N_14315);
and UO_473 (O_473,N_14906,N_14605);
or UO_474 (O_474,N_14675,N_14302);
and UO_475 (O_475,N_14291,N_14496);
nor UO_476 (O_476,N_14484,N_14794);
xor UO_477 (O_477,N_14846,N_14655);
nor UO_478 (O_478,N_14613,N_14513);
nand UO_479 (O_479,N_14853,N_14287);
xnor UO_480 (O_480,N_14344,N_14447);
and UO_481 (O_481,N_14344,N_14320);
or UO_482 (O_482,N_14735,N_14722);
and UO_483 (O_483,N_14972,N_14539);
and UO_484 (O_484,N_14366,N_14765);
nor UO_485 (O_485,N_14373,N_14382);
nor UO_486 (O_486,N_14422,N_14313);
and UO_487 (O_487,N_14436,N_14270);
nand UO_488 (O_488,N_14820,N_14357);
and UO_489 (O_489,N_14413,N_14354);
nor UO_490 (O_490,N_14954,N_14366);
or UO_491 (O_491,N_14453,N_14773);
or UO_492 (O_492,N_14637,N_14680);
and UO_493 (O_493,N_14372,N_14806);
nand UO_494 (O_494,N_14346,N_14922);
or UO_495 (O_495,N_14532,N_14757);
xnor UO_496 (O_496,N_14700,N_14556);
nor UO_497 (O_497,N_14787,N_14603);
nand UO_498 (O_498,N_14870,N_14721);
and UO_499 (O_499,N_14662,N_14554);
nand UO_500 (O_500,N_14417,N_14796);
nand UO_501 (O_501,N_14654,N_14874);
xor UO_502 (O_502,N_14633,N_14498);
nand UO_503 (O_503,N_14633,N_14955);
or UO_504 (O_504,N_14547,N_14431);
and UO_505 (O_505,N_14603,N_14381);
nor UO_506 (O_506,N_14731,N_14926);
and UO_507 (O_507,N_14348,N_14588);
nand UO_508 (O_508,N_14304,N_14624);
nor UO_509 (O_509,N_14710,N_14844);
xnor UO_510 (O_510,N_14863,N_14753);
and UO_511 (O_511,N_14316,N_14831);
xor UO_512 (O_512,N_14659,N_14413);
nor UO_513 (O_513,N_14319,N_14562);
nor UO_514 (O_514,N_14270,N_14552);
and UO_515 (O_515,N_14987,N_14253);
nor UO_516 (O_516,N_14559,N_14334);
or UO_517 (O_517,N_14614,N_14780);
or UO_518 (O_518,N_14738,N_14460);
nand UO_519 (O_519,N_14714,N_14892);
or UO_520 (O_520,N_14292,N_14389);
nor UO_521 (O_521,N_14809,N_14891);
xnor UO_522 (O_522,N_14774,N_14653);
xor UO_523 (O_523,N_14841,N_14567);
nor UO_524 (O_524,N_14658,N_14973);
or UO_525 (O_525,N_14859,N_14627);
nor UO_526 (O_526,N_14361,N_14909);
nand UO_527 (O_527,N_14591,N_14422);
xor UO_528 (O_528,N_14438,N_14655);
or UO_529 (O_529,N_14813,N_14799);
and UO_530 (O_530,N_14890,N_14974);
nor UO_531 (O_531,N_14436,N_14326);
xnor UO_532 (O_532,N_14702,N_14560);
or UO_533 (O_533,N_14288,N_14804);
xor UO_534 (O_534,N_14908,N_14363);
nand UO_535 (O_535,N_14306,N_14852);
or UO_536 (O_536,N_14342,N_14500);
nand UO_537 (O_537,N_14406,N_14977);
nor UO_538 (O_538,N_14887,N_14719);
or UO_539 (O_539,N_14350,N_14270);
and UO_540 (O_540,N_14436,N_14512);
nor UO_541 (O_541,N_14781,N_14660);
nor UO_542 (O_542,N_14894,N_14743);
and UO_543 (O_543,N_14705,N_14547);
xnor UO_544 (O_544,N_14783,N_14784);
nand UO_545 (O_545,N_14623,N_14703);
and UO_546 (O_546,N_14510,N_14842);
and UO_547 (O_547,N_14815,N_14582);
and UO_548 (O_548,N_14957,N_14938);
and UO_549 (O_549,N_14854,N_14473);
nand UO_550 (O_550,N_14665,N_14520);
or UO_551 (O_551,N_14522,N_14455);
nand UO_552 (O_552,N_14778,N_14769);
or UO_553 (O_553,N_14503,N_14323);
nor UO_554 (O_554,N_14752,N_14881);
or UO_555 (O_555,N_14479,N_14785);
and UO_556 (O_556,N_14524,N_14722);
and UO_557 (O_557,N_14626,N_14319);
nor UO_558 (O_558,N_14978,N_14668);
and UO_559 (O_559,N_14707,N_14331);
or UO_560 (O_560,N_14542,N_14712);
nand UO_561 (O_561,N_14810,N_14409);
nand UO_562 (O_562,N_14735,N_14636);
nand UO_563 (O_563,N_14472,N_14492);
nand UO_564 (O_564,N_14557,N_14414);
nand UO_565 (O_565,N_14406,N_14770);
or UO_566 (O_566,N_14792,N_14748);
and UO_567 (O_567,N_14485,N_14890);
nand UO_568 (O_568,N_14915,N_14988);
xor UO_569 (O_569,N_14927,N_14632);
nor UO_570 (O_570,N_14432,N_14607);
and UO_571 (O_571,N_14326,N_14600);
or UO_572 (O_572,N_14728,N_14851);
and UO_573 (O_573,N_14895,N_14563);
and UO_574 (O_574,N_14263,N_14385);
and UO_575 (O_575,N_14807,N_14928);
or UO_576 (O_576,N_14284,N_14614);
and UO_577 (O_577,N_14379,N_14711);
and UO_578 (O_578,N_14440,N_14962);
or UO_579 (O_579,N_14475,N_14943);
and UO_580 (O_580,N_14664,N_14872);
or UO_581 (O_581,N_14583,N_14425);
or UO_582 (O_582,N_14600,N_14566);
and UO_583 (O_583,N_14766,N_14304);
nor UO_584 (O_584,N_14517,N_14587);
or UO_585 (O_585,N_14657,N_14966);
nand UO_586 (O_586,N_14633,N_14482);
nor UO_587 (O_587,N_14277,N_14558);
and UO_588 (O_588,N_14467,N_14343);
nor UO_589 (O_589,N_14289,N_14483);
nand UO_590 (O_590,N_14275,N_14917);
nand UO_591 (O_591,N_14674,N_14656);
and UO_592 (O_592,N_14256,N_14343);
xor UO_593 (O_593,N_14294,N_14946);
or UO_594 (O_594,N_14347,N_14912);
or UO_595 (O_595,N_14931,N_14355);
nor UO_596 (O_596,N_14764,N_14530);
nor UO_597 (O_597,N_14749,N_14920);
nand UO_598 (O_598,N_14278,N_14934);
nand UO_599 (O_599,N_14426,N_14964);
nand UO_600 (O_600,N_14958,N_14910);
nor UO_601 (O_601,N_14304,N_14992);
or UO_602 (O_602,N_14318,N_14736);
and UO_603 (O_603,N_14619,N_14657);
or UO_604 (O_604,N_14295,N_14669);
and UO_605 (O_605,N_14383,N_14890);
nand UO_606 (O_606,N_14941,N_14710);
and UO_607 (O_607,N_14615,N_14817);
nand UO_608 (O_608,N_14256,N_14273);
nand UO_609 (O_609,N_14958,N_14634);
or UO_610 (O_610,N_14289,N_14998);
nor UO_611 (O_611,N_14327,N_14803);
nor UO_612 (O_612,N_14757,N_14991);
nand UO_613 (O_613,N_14280,N_14611);
nor UO_614 (O_614,N_14598,N_14439);
xor UO_615 (O_615,N_14420,N_14903);
nand UO_616 (O_616,N_14803,N_14326);
and UO_617 (O_617,N_14952,N_14753);
and UO_618 (O_618,N_14883,N_14781);
and UO_619 (O_619,N_14487,N_14628);
and UO_620 (O_620,N_14426,N_14322);
nor UO_621 (O_621,N_14350,N_14710);
nand UO_622 (O_622,N_14368,N_14871);
nor UO_623 (O_623,N_14602,N_14357);
nand UO_624 (O_624,N_14625,N_14290);
or UO_625 (O_625,N_14804,N_14312);
or UO_626 (O_626,N_14982,N_14275);
or UO_627 (O_627,N_14620,N_14508);
nor UO_628 (O_628,N_14519,N_14731);
nand UO_629 (O_629,N_14422,N_14628);
and UO_630 (O_630,N_14768,N_14776);
nor UO_631 (O_631,N_14686,N_14614);
xnor UO_632 (O_632,N_14386,N_14818);
xor UO_633 (O_633,N_14859,N_14600);
xor UO_634 (O_634,N_14693,N_14912);
or UO_635 (O_635,N_14822,N_14463);
nand UO_636 (O_636,N_14611,N_14286);
or UO_637 (O_637,N_14899,N_14755);
and UO_638 (O_638,N_14341,N_14999);
nand UO_639 (O_639,N_14737,N_14663);
nor UO_640 (O_640,N_14777,N_14753);
xnor UO_641 (O_641,N_14556,N_14276);
nor UO_642 (O_642,N_14279,N_14902);
nor UO_643 (O_643,N_14975,N_14500);
xnor UO_644 (O_644,N_14443,N_14358);
or UO_645 (O_645,N_14842,N_14834);
nor UO_646 (O_646,N_14811,N_14337);
nor UO_647 (O_647,N_14792,N_14985);
and UO_648 (O_648,N_14974,N_14878);
nor UO_649 (O_649,N_14343,N_14817);
and UO_650 (O_650,N_14584,N_14441);
nor UO_651 (O_651,N_14652,N_14692);
and UO_652 (O_652,N_14438,N_14797);
or UO_653 (O_653,N_14802,N_14791);
nand UO_654 (O_654,N_14941,N_14384);
nor UO_655 (O_655,N_14301,N_14539);
nor UO_656 (O_656,N_14659,N_14470);
nand UO_657 (O_657,N_14315,N_14270);
nor UO_658 (O_658,N_14520,N_14993);
nor UO_659 (O_659,N_14804,N_14258);
or UO_660 (O_660,N_14315,N_14278);
nor UO_661 (O_661,N_14642,N_14724);
and UO_662 (O_662,N_14572,N_14801);
nor UO_663 (O_663,N_14518,N_14746);
and UO_664 (O_664,N_14747,N_14495);
or UO_665 (O_665,N_14775,N_14403);
nor UO_666 (O_666,N_14387,N_14629);
nand UO_667 (O_667,N_14300,N_14681);
nand UO_668 (O_668,N_14717,N_14660);
xor UO_669 (O_669,N_14426,N_14439);
or UO_670 (O_670,N_14297,N_14816);
xor UO_671 (O_671,N_14539,N_14433);
and UO_672 (O_672,N_14537,N_14851);
xor UO_673 (O_673,N_14771,N_14510);
nor UO_674 (O_674,N_14689,N_14299);
xnor UO_675 (O_675,N_14346,N_14364);
or UO_676 (O_676,N_14704,N_14480);
nand UO_677 (O_677,N_14599,N_14637);
nor UO_678 (O_678,N_14682,N_14487);
or UO_679 (O_679,N_14917,N_14541);
or UO_680 (O_680,N_14725,N_14302);
nor UO_681 (O_681,N_14336,N_14750);
xor UO_682 (O_682,N_14256,N_14875);
and UO_683 (O_683,N_14870,N_14827);
nor UO_684 (O_684,N_14319,N_14691);
and UO_685 (O_685,N_14901,N_14845);
or UO_686 (O_686,N_14740,N_14451);
nand UO_687 (O_687,N_14288,N_14834);
or UO_688 (O_688,N_14448,N_14967);
and UO_689 (O_689,N_14971,N_14349);
nand UO_690 (O_690,N_14586,N_14994);
nand UO_691 (O_691,N_14718,N_14848);
xnor UO_692 (O_692,N_14378,N_14266);
nor UO_693 (O_693,N_14829,N_14814);
nor UO_694 (O_694,N_14621,N_14722);
nand UO_695 (O_695,N_14765,N_14662);
and UO_696 (O_696,N_14661,N_14333);
or UO_697 (O_697,N_14774,N_14338);
or UO_698 (O_698,N_14931,N_14862);
nand UO_699 (O_699,N_14338,N_14959);
nand UO_700 (O_700,N_14301,N_14963);
nor UO_701 (O_701,N_14873,N_14607);
nor UO_702 (O_702,N_14510,N_14791);
nor UO_703 (O_703,N_14724,N_14828);
and UO_704 (O_704,N_14884,N_14934);
or UO_705 (O_705,N_14751,N_14611);
and UO_706 (O_706,N_14595,N_14523);
or UO_707 (O_707,N_14909,N_14522);
nor UO_708 (O_708,N_14716,N_14653);
nand UO_709 (O_709,N_14425,N_14485);
nand UO_710 (O_710,N_14492,N_14839);
nand UO_711 (O_711,N_14896,N_14918);
nor UO_712 (O_712,N_14960,N_14571);
or UO_713 (O_713,N_14493,N_14903);
nand UO_714 (O_714,N_14659,N_14282);
or UO_715 (O_715,N_14563,N_14632);
nor UO_716 (O_716,N_14814,N_14381);
or UO_717 (O_717,N_14495,N_14932);
nor UO_718 (O_718,N_14796,N_14797);
nor UO_719 (O_719,N_14430,N_14427);
or UO_720 (O_720,N_14762,N_14496);
nor UO_721 (O_721,N_14651,N_14854);
nor UO_722 (O_722,N_14324,N_14990);
or UO_723 (O_723,N_14668,N_14667);
or UO_724 (O_724,N_14277,N_14816);
and UO_725 (O_725,N_14473,N_14683);
nand UO_726 (O_726,N_14662,N_14522);
or UO_727 (O_727,N_14253,N_14507);
or UO_728 (O_728,N_14927,N_14314);
and UO_729 (O_729,N_14778,N_14424);
nand UO_730 (O_730,N_14794,N_14369);
and UO_731 (O_731,N_14423,N_14335);
or UO_732 (O_732,N_14479,N_14376);
or UO_733 (O_733,N_14778,N_14751);
nor UO_734 (O_734,N_14991,N_14539);
and UO_735 (O_735,N_14715,N_14349);
and UO_736 (O_736,N_14421,N_14687);
xnor UO_737 (O_737,N_14489,N_14254);
xnor UO_738 (O_738,N_14681,N_14667);
and UO_739 (O_739,N_14958,N_14956);
xnor UO_740 (O_740,N_14615,N_14912);
nand UO_741 (O_741,N_14787,N_14944);
and UO_742 (O_742,N_14757,N_14497);
and UO_743 (O_743,N_14914,N_14367);
nand UO_744 (O_744,N_14535,N_14741);
nor UO_745 (O_745,N_14767,N_14806);
or UO_746 (O_746,N_14866,N_14437);
or UO_747 (O_747,N_14875,N_14771);
nand UO_748 (O_748,N_14837,N_14369);
or UO_749 (O_749,N_14947,N_14289);
nand UO_750 (O_750,N_14712,N_14740);
nand UO_751 (O_751,N_14365,N_14989);
xor UO_752 (O_752,N_14695,N_14970);
or UO_753 (O_753,N_14563,N_14912);
nand UO_754 (O_754,N_14853,N_14530);
nand UO_755 (O_755,N_14778,N_14432);
and UO_756 (O_756,N_14729,N_14791);
or UO_757 (O_757,N_14582,N_14980);
nor UO_758 (O_758,N_14792,N_14263);
nor UO_759 (O_759,N_14595,N_14306);
xor UO_760 (O_760,N_14517,N_14763);
nand UO_761 (O_761,N_14333,N_14660);
nor UO_762 (O_762,N_14950,N_14300);
nor UO_763 (O_763,N_14861,N_14524);
nand UO_764 (O_764,N_14348,N_14370);
nor UO_765 (O_765,N_14955,N_14722);
or UO_766 (O_766,N_14583,N_14447);
nor UO_767 (O_767,N_14859,N_14994);
nand UO_768 (O_768,N_14889,N_14625);
nand UO_769 (O_769,N_14373,N_14875);
and UO_770 (O_770,N_14598,N_14554);
or UO_771 (O_771,N_14632,N_14400);
and UO_772 (O_772,N_14691,N_14719);
or UO_773 (O_773,N_14786,N_14416);
and UO_774 (O_774,N_14576,N_14733);
or UO_775 (O_775,N_14295,N_14573);
or UO_776 (O_776,N_14565,N_14272);
xor UO_777 (O_777,N_14470,N_14759);
or UO_778 (O_778,N_14902,N_14469);
and UO_779 (O_779,N_14826,N_14568);
nor UO_780 (O_780,N_14837,N_14302);
nand UO_781 (O_781,N_14890,N_14421);
nand UO_782 (O_782,N_14502,N_14393);
nand UO_783 (O_783,N_14956,N_14657);
and UO_784 (O_784,N_14389,N_14775);
and UO_785 (O_785,N_14757,N_14859);
or UO_786 (O_786,N_14992,N_14576);
xor UO_787 (O_787,N_14433,N_14375);
or UO_788 (O_788,N_14644,N_14774);
nand UO_789 (O_789,N_14349,N_14850);
or UO_790 (O_790,N_14715,N_14611);
nand UO_791 (O_791,N_14720,N_14644);
xor UO_792 (O_792,N_14976,N_14921);
nand UO_793 (O_793,N_14694,N_14804);
nand UO_794 (O_794,N_14836,N_14761);
nor UO_795 (O_795,N_14868,N_14341);
nand UO_796 (O_796,N_14534,N_14589);
xnor UO_797 (O_797,N_14357,N_14503);
nand UO_798 (O_798,N_14925,N_14962);
and UO_799 (O_799,N_14491,N_14472);
or UO_800 (O_800,N_14612,N_14683);
nand UO_801 (O_801,N_14515,N_14671);
or UO_802 (O_802,N_14316,N_14796);
nand UO_803 (O_803,N_14677,N_14990);
nand UO_804 (O_804,N_14456,N_14317);
nor UO_805 (O_805,N_14689,N_14960);
nor UO_806 (O_806,N_14420,N_14528);
or UO_807 (O_807,N_14994,N_14390);
nor UO_808 (O_808,N_14337,N_14861);
nand UO_809 (O_809,N_14908,N_14334);
or UO_810 (O_810,N_14598,N_14266);
xor UO_811 (O_811,N_14669,N_14601);
and UO_812 (O_812,N_14633,N_14819);
and UO_813 (O_813,N_14867,N_14672);
and UO_814 (O_814,N_14807,N_14609);
nor UO_815 (O_815,N_14546,N_14489);
or UO_816 (O_816,N_14929,N_14630);
and UO_817 (O_817,N_14550,N_14885);
nand UO_818 (O_818,N_14481,N_14422);
or UO_819 (O_819,N_14668,N_14597);
xnor UO_820 (O_820,N_14668,N_14315);
and UO_821 (O_821,N_14482,N_14790);
and UO_822 (O_822,N_14378,N_14750);
nand UO_823 (O_823,N_14258,N_14786);
or UO_824 (O_824,N_14656,N_14312);
nor UO_825 (O_825,N_14767,N_14505);
or UO_826 (O_826,N_14494,N_14510);
or UO_827 (O_827,N_14718,N_14970);
nand UO_828 (O_828,N_14655,N_14882);
nor UO_829 (O_829,N_14632,N_14559);
or UO_830 (O_830,N_14276,N_14641);
and UO_831 (O_831,N_14305,N_14522);
nand UO_832 (O_832,N_14464,N_14360);
nor UO_833 (O_833,N_14848,N_14820);
nor UO_834 (O_834,N_14583,N_14382);
or UO_835 (O_835,N_14960,N_14440);
and UO_836 (O_836,N_14662,N_14338);
and UO_837 (O_837,N_14842,N_14711);
nor UO_838 (O_838,N_14267,N_14756);
or UO_839 (O_839,N_14873,N_14452);
or UO_840 (O_840,N_14752,N_14575);
nand UO_841 (O_841,N_14946,N_14362);
nand UO_842 (O_842,N_14455,N_14695);
and UO_843 (O_843,N_14756,N_14613);
nor UO_844 (O_844,N_14776,N_14281);
and UO_845 (O_845,N_14918,N_14793);
xor UO_846 (O_846,N_14888,N_14607);
nor UO_847 (O_847,N_14481,N_14978);
or UO_848 (O_848,N_14736,N_14772);
or UO_849 (O_849,N_14596,N_14688);
or UO_850 (O_850,N_14700,N_14738);
nor UO_851 (O_851,N_14839,N_14349);
and UO_852 (O_852,N_14423,N_14328);
nand UO_853 (O_853,N_14899,N_14953);
or UO_854 (O_854,N_14907,N_14472);
and UO_855 (O_855,N_14830,N_14980);
or UO_856 (O_856,N_14694,N_14891);
nand UO_857 (O_857,N_14261,N_14759);
nor UO_858 (O_858,N_14337,N_14339);
nand UO_859 (O_859,N_14582,N_14539);
or UO_860 (O_860,N_14947,N_14624);
xor UO_861 (O_861,N_14408,N_14330);
nor UO_862 (O_862,N_14343,N_14606);
nand UO_863 (O_863,N_14415,N_14370);
xnor UO_864 (O_864,N_14660,N_14560);
nand UO_865 (O_865,N_14993,N_14384);
or UO_866 (O_866,N_14785,N_14669);
nand UO_867 (O_867,N_14672,N_14393);
or UO_868 (O_868,N_14541,N_14828);
or UO_869 (O_869,N_14523,N_14798);
xnor UO_870 (O_870,N_14702,N_14599);
and UO_871 (O_871,N_14334,N_14522);
and UO_872 (O_872,N_14758,N_14269);
and UO_873 (O_873,N_14517,N_14498);
nand UO_874 (O_874,N_14672,N_14827);
or UO_875 (O_875,N_14858,N_14994);
xnor UO_876 (O_876,N_14919,N_14896);
nor UO_877 (O_877,N_14503,N_14439);
and UO_878 (O_878,N_14605,N_14728);
nor UO_879 (O_879,N_14357,N_14345);
or UO_880 (O_880,N_14589,N_14737);
xnor UO_881 (O_881,N_14682,N_14850);
nor UO_882 (O_882,N_14277,N_14494);
nand UO_883 (O_883,N_14827,N_14598);
xnor UO_884 (O_884,N_14526,N_14860);
nand UO_885 (O_885,N_14756,N_14769);
and UO_886 (O_886,N_14557,N_14694);
and UO_887 (O_887,N_14320,N_14493);
nand UO_888 (O_888,N_14656,N_14615);
nand UO_889 (O_889,N_14752,N_14352);
or UO_890 (O_890,N_14581,N_14468);
or UO_891 (O_891,N_14662,N_14268);
nand UO_892 (O_892,N_14577,N_14992);
nor UO_893 (O_893,N_14802,N_14704);
nand UO_894 (O_894,N_14722,N_14858);
nand UO_895 (O_895,N_14533,N_14362);
or UO_896 (O_896,N_14359,N_14408);
nand UO_897 (O_897,N_14284,N_14813);
or UO_898 (O_898,N_14921,N_14639);
nand UO_899 (O_899,N_14523,N_14418);
nand UO_900 (O_900,N_14490,N_14724);
and UO_901 (O_901,N_14796,N_14554);
nand UO_902 (O_902,N_14316,N_14982);
or UO_903 (O_903,N_14553,N_14365);
and UO_904 (O_904,N_14787,N_14283);
xor UO_905 (O_905,N_14613,N_14781);
xnor UO_906 (O_906,N_14372,N_14871);
nor UO_907 (O_907,N_14513,N_14829);
nor UO_908 (O_908,N_14611,N_14443);
xnor UO_909 (O_909,N_14806,N_14404);
nand UO_910 (O_910,N_14296,N_14284);
and UO_911 (O_911,N_14902,N_14521);
nor UO_912 (O_912,N_14997,N_14259);
and UO_913 (O_913,N_14640,N_14783);
and UO_914 (O_914,N_14939,N_14657);
and UO_915 (O_915,N_14608,N_14567);
nor UO_916 (O_916,N_14488,N_14414);
or UO_917 (O_917,N_14889,N_14710);
nor UO_918 (O_918,N_14599,N_14384);
and UO_919 (O_919,N_14313,N_14385);
nor UO_920 (O_920,N_14313,N_14462);
nor UO_921 (O_921,N_14862,N_14579);
and UO_922 (O_922,N_14920,N_14740);
and UO_923 (O_923,N_14929,N_14914);
and UO_924 (O_924,N_14691,N_14961);
or UO_925 (O_925,N_14390,N_14385);
nor UO_926 (O_926,N_14841,N_14403);
and UO_927 (O_927,N_14917,N_14440);
and UO_928 (O_928,N_14947,N_14826);
nand UO_929 (O_929,N_14706,N_14469);
or UO_930 (O_930,N_14707,N_14356);
nand UO_931 (O_931,N_14304,N_14991);
nand UO_932 (O_932,N_14442,N_14440);
nand UO_933 (O_933,N_14744,N_14346);
nor UO_934 (O_934,N_14282,N_14402);
nand UO_935 (O_935,N_14365,N_14255);
or UO_936 (O_936,N_14685,N_14669);
xor UO_937 (O_937,N_14631,N_14865);
or UO_938 (O_938,N_14824,N_14442);
xnor UO_939 (O_939,N_14379,N_14550);
xor UO_940 (O_940,N_14917,N_14726);
or UO_941 (O_941,N_14904,N_14872);
nor UO_942 (O_942,N_14362,N_14687);
nand UO_943 (O_943,N_14782,N_14752);
nor UO_944 (O_944,N_14313,N_14805);
nand UO_945 (O_945,N_14399,N_14316);
xnor UO_946 (O_946,N_14772,N_14877);
nand UO_947 (O_947,N_14255,N_14945);
and UO_948 (O_948,N_14658,N_14310);
and UO_949 (O_949,N_14863,N_14976);
or UO_950 (O_950,N_14860,N_14685);
and UO_951 (O_951,N_14709,N_14371);
or UO_952 (O_952,N_14505,N_14765);
nand UO_953 (O_953,N_14363,N_14412);
and UO_954 (O_954,N_14282,N_14914);
nor UO_955 (O_955,N_14371,N_14891);
nand UO_956 (O_956,N_14734,N_14451);
and UO_957 (O_957,N_14483,N_14793);
nor UO_958 (O_958,N_14790,N_14564);
and UO_959 (O_959,N_14351,N_14734);
and UO_960 (O_960,N_14721,N_14803);
or UO_961 (O_961,N_14828,N_14435);
and UO_962 (O_962,N_14265,N_14701);
or UO_963 (O_963,N_14954,N_14886);
and UO_964 (O_964,N_14548,N_14483);
nand UO_965 (O_965,N_14577,N_14458);
and UO_966 (O_966,N_14774,N_14670);
nand UO_967 (O_967,N_14762,N_14353);
and UO_968 (O_968,N_14795,N_14285);
nand UO_969 (O_969,N_14585,N_14697);
nor UO_970 (O_970,N_14386,N_14974);
nor UO_971 (O_971,N_14362,N_14830);
nand UO_972 (O_972,N_14289,N_14861);
nor UO_973 (O_973,N_14653,N_14490);
nor UO_974 (O_974,N_14280,N_14797);
or UO_975 (O_975,N_14422,N_14503);
nand UO_976 (O_976,N_14817,N_14664);
or UO_977 (O_977,N_14896,N_14717);
nor UO_978 (O_978,N_14447,N_14960);
xor UO_979 (O_979,N_14362,N_14769);
and UO_980 (O_980,N_14468,N_14495);
or UO_981 (O_981,N_14424,N_14361);
nor UO_982 (O_982,N_14303,N_14858);
and UO_983 (O_983,N_14762,N_14704);
nor UO_984 (O_984,N_14612,N_14894);
nand UO_985 (O_985,N_14736,N_14564);
nor UO_986 (O_986,N_14538,N_14540);
nand UO_987 (O_987,N_14866,N_14468);
nand UO_988 (O_988,N_14817,N_14659);
or UO_989 (O_989,N_14573,N_14983);
or UO_990 (O_990,N_14865,N_14789);
and UO_991 (O_991,N_14440,N_14272);
xnor UO_992 (O_992,N_14740,N_14782);
nor UO_993 (O_993,N_14425,N_14718);
nor UO_994 (O_994,N_14379,N_14664);
nor UO_995 (O_995,N_14809,N_14396);
nand UO_996 (O_996,N_14726,N_14885);
or UO_997 (O_997,N_14791,N_14837);
nand UO_998 (O_998,N_14718,N_14683);
nand UO_999 (O_999,N_14969,N_14628);
or UO_1000 (O_1000,N_14828,N_14956);
and UO_1001 (O_1001,N_14531,N_14853);
and UO_1002 (O_1002,N_14356,N_14560);
or UO_1003 (O_1003,N_14657,N_14875);
or UO_1004 (O_1004,N_14285,N_14717);
xnor UO_1005 (O_1005,N_14582,N_14666);
nor UO_1006 (O_1006,N_14446,N_14593);
or UO_1007 (O_1007,N_14704,N_14597);
nand UO_1008 (O_1008,N_14503,N_14874);
and UO_1009 (O_1009,N_14322,N_14858);
and UO_1010 (O_1010,N_14374,N_14838);
nor UO_1011 (O_1011,N_14786,N_14610);
nand UO_1012 (O_1012,N_14934,N_14494);
and UO_1013 (O_1013,N_14271,N_14529);
nand UO_1014 (O_1014,N_14295,N_14546);
nor UO_1015 (O_1015,N_14826,N_14573);
and UO_1016 (O_1016,N_14957,N_14548);
and UO_1017 (O_1017,N_14467,N_14517);
nand UO_1018 (O_1018,N_14572,N_14362);
nand UO_1019 (O_1019,N_14485,N_14612);
xor UO_1020 (O_1020,N_14761,N_14699);
nor UO_1021 (O_1021,N_14329,N_14994);
nor UO_1022 (O_1022,N_14298,N_14375);
nand UO_1023 (O_1023,N_14392,N_14826);
xor UO_1024 (O_1024,N_14310,N_14408);
nor UO_1025 (O_1025,N_14982,N_14287);
or UO_1026 (O_1026,N_14382,N_14672);
or UO_1027 (O_1027,N_14946,N_14848);
nand UO_1028 (O_1028,N_14429,N_14948);
and UO_1029 (O_1029,N_14906,N_14746);
nor UO_1030 (O_1030,N_14959,N_14417);
or UO_1031 (O_1031,N_14710,N_14960);
and UO_1032 (O_1032,N_14381,N_14361);
or UO_1033 (O_1033,N_14756,N_14329);
nor UO_1034 (O_1034,N_14614,N_14745);
nand UO_1035 (O_1035,N_14689,N_14436);
xnor UO_1036 (O_1036,N_14852,N_14939);
nand UO_1037 (O_1037,N_14597,N_14474);
and UO_1038 (O_1038,N_14928,N_14346);
and UO_1039 (O_1039,N_14575,N_14573);
nand UO_1040 (O_1040,N_14270,N_14357);
or UO_1041 (O_1041,N_14797,N_14563);
or UO_1042 (O_1042,N_14271,N_14482);
nand UO_1043 (O_1043,N_14980,N_14913);
and UO_1044 (O_1044,N_14441,N_14951);
or UO_1045 (O_1045,N_14456,N_14990);
nand UO_1046 (O_1046,N_14670,N_14344);
nor UO_1047 (O_1047,N_14284,N_14467);
or UO_1048 (O_1048,N_14807,N_14254);
nand UO_1049 (O_1049,N_14818,N_14457);
nor UO_1050 (O_1050,N_14387,N_14420);
or UO_1051 (O_1051,N_14400,N_14678);
or UO_1052 (O_1052,N_14505,N_14714);
nand UO_1053 (O_1053,N_14988,N_14785);
and UO_1054 (O_1054,N_14415,N_14806);
nand UO_1055 (O_1055,N_14823,N_14537);
nand UO_1056 (O_1056,N_14470,N_14679);
nand UO_1057 (O_1057,N_14993,N_14452);
nand UO_1058 (O_1058,N_14295,N_14375);
and UO_1059 (O_1059,N_14456,N_14292);
nor UO_1060 (O_1060,N_14982,N_14903);
and UO_1061 (O_1061,N_14882,N_14349);
or UO_1062 (O_1062,N_14638,N_14840);
or UO_1063 (O_1063,N_14536,N_14309);
nand UO_1064 (O_1064,N_14795,N_14287);
and UO_1065 (O_1065,N_14761,N_14924);
and UO_1066 (O_1066,N_14497,N_14286);
nand UO_1067 (O_1067,N_14385,N_14702);
and UO_1068 (O_1068,N_14394,N_14660);
and UO_1069 (O_1069,N_14678,N_14767);
xnor UO_1070 (O_1070,N_14388,N_14724);
and UO_1071 (O_1071,N_14559,N_14808);
or UO_1072 (O_1072,N_14348,N_14662);
nand UO_1073 (O_1073,N_14956,N_14693);
xor UO_1074 (O_1074,N_14831,N_14609);
and UO_1075 (O_1075,N_14343,N_14935);
or UO_1076 (O_1076,N_14660,N_14866);
nand UO_1077 (O_1077,N_14325,N_14550);
and UO_1078 (O_1078,N_14826,N_14831);
and UO_1079 (O_1079,N_14523,N_14299);
or UO_1080 (O_1080,N_14350,N_14820);
nand UO_1081 (O_1081,N_14649,N_14982);
nand UO_1082 (O_1082,N_14357,N_14504);
or UO_1083 (O_1083,N_14536,N_14455);
and UO_1084 (O_1084,N_14893,N_14308);
and UO_1085 (O_1085,N_14791,N_14456);
nor UO_1086 (O_1086,N_14920,N_14642);
nand UO_1087 (O_1087,N_14787,N_14592);
nor UO_1088 (O_1088,N_14759,N_14354);
and UO_1089 (O_1089,N_14594,N_14263);
and UO_1090 (O_1090,N_14936,N_14863);
or UO_1091 (O_1091,N_14379,N_14299);
or UO_1092 (O_1092,N_14590,N_14992);
or UO_1093 (O_1093,N_14951,N_14850);
or UO_1094 (O_1094,N_14865,N_14316);
nand UO_1095 (O_1095,N_14609,N_14538);
and UO_1096 (O_1096,N_14744,N_14601);
and UO_1097 (O_1097,N_14308,N_14587);
or UO_1098 (O_1098,N_14708,N_14820);
or UO_1099 (O_1099,N_14981,N_14811);
or UO_1100 (O_1100,N_14397,N_14863);
or UO_1101 (O_1101,N_14873,N_14838);
nor UO_1102 (O_1102,N_14781,N_14488);
and UO_1103 (O_1103,N_14740,N_14268);
nand UO_1104 (O_1104,N_14829,N_14318);
or UO_1105 (O_1105,N_14780,N_14606);
nor UO_1106 (O_1106,N_14679,N_14543);
nand UO_1107 (O_1107,N_14557,N_14906);
nand UO_1108 (O_1108,N_14425,N_14311);
or UO_1109 (O_1109,N_14270,N_14908);
nor UO_1110 (O_1110,N_14972,N_14426);
nor UO_1111 (O_1111,N_14722,N_14602);
nand UO_1112 (O_1112,N_14336,N_14537);
nor UO_1113 (O_1113,N_14871,N_14806);
nand UO_1114 (O_1114,N_14533,N_14521);
and UO_1115 (O_1115,N_14379,N_14922);
and UO_1116 (O_1116,N_14914,N_14527);
xor UO_1117 (O_1117,N_14975,N_14988);
nand UO_1118 (O_1118,N_14998,N_14319);
or UO_1119 (O_1119,N_14569,N_14912);
or UO_1120 (O_1120,N_14457,N_14764);
nor UO_1121 (O_1121,N_14691,N_14401);
xnor UO_1122 (O_1122,N_14373,N_14463);
or UO_1123 (O_1123,N_14271,N_14386);
or UO_1124 (O_1124,N_14784,N_14632);
nand UO_1125 (O_1125,N_14878,N_14344);
nand UO_1126 (O_1126,N_14326,N_14800);
and UO_1127 (O_1127,N_14713,N_14668);
or UO_1128 (O_1128,N_14940,N_14555);
and UO_1129 (O_1129,N_14374,N_14300);
and UO_1130 (O_1130,N_14901,N_14537);
and UO_1131 (O_1131,N_14808,N_14667);
nand UO_1132 (O_1132,N_14850,N_14375);
nor UO_1133 (O_1133,N_14328,N_14697);
nand UO_1134 (O_1134,N_14509,N_14723);
nand UO_1135 (O_1135,N_14444,N_14922);
nand UO_1136 (O_1136,N_14588,N_14886);
and UO_1137 (O_1137,N_14929,N_14709);
and UO_1138 (O_1138,N_14929,N_14369);
nor UO_1139 (O_1139,N_14309,N_14367);
and UO_1140 (O_1140,N_14702,N_14391);
or UO_1141 (O_1141,N_14811,N_14498);
nor UO_1142 (O_1142,N_14568,N_14413);
and UO_1143 (O_1143,N_14552,N_14632);
nor UO_1144 (O_1144,N_14703,N_14957);
nor UO_1145 (O_1145,N_14407,N_14940);
and UO_1146 (O_1146,N_14613,N_14990);
nand UO_1147 (O_1147,N_14994,N_14812);
nor UO_1148 (O_1148,N_14519,N_14310);
nor UO_1149 (O_1149,N_14960,N_14564);
nor UO_1150 (O_1150,N_14285,N_14740);
nand UO_1151 (O_1151,N_14534,N_14987);
nand UO_1152 (O_1152,N_14642,N_14644);
nor UO_1153 (O_1153,N_14408,N_14978);
nor UO_1154 (O_1154,N_14631,N_14425);
nor UO_1155 (O_1155,N_14329,N_14325);
or UO_1156 (O_1156,N_14370,N_14376);
and UO_1157 (O_1157,N_14373,N_14357);
xor UO_1158 (O_1158,N_14332,N_14341);
and UO_1159 (O_1159,N_14955,N_14901);
nor UO_1160 (O_1160,N_14819,N_14389);
or UO_1161 (O_1161,N_14564,N_14643);
or UO_1162 (O_1162,N_14430,N_14589);
and UO_1163 (O_1163,N_14450,N_14389);
nand UO_1164 (O_1164,N_14383,N_14377);
or UO_1165 (O_1165,N_14493,N_14666);
and UO_1166 (O_1166,N_14571,N_14662);
or UO_1167 (O_1167,N_14637,N_14579);
and UO_1168 (O_1168,N_14952,N_14330);
or UO_1169 (O_1169,N_14437,N_14738);
nand UO_1170 (O_1170,N_14607,N_14758);
and UO_1171 (O_1171,N_14999,N_14861);
nor UO_1172 (O_1172,N_14805,N_14488);
and UO_1173 (O_1173,N_14435,N_14535);
xnor UO_1174 (O_1174,N_14304,N_14739);
and UO_1175 (O_1175,N_14297,N_14851);
or UO_1176 (O_1176,N_14545,N_14505);
or UO_1177 (O_1177,N_14809,N_14824);
and UO_1178 (O_1178,N_14970,N_14547);
nand UO_1179 (O_1179,N_14713,N_14302);
nand UO_1180 (O_1180,N_14474,N_14480);
xnor UO_1181 (O_1181,N_14837,N_14792);
and UO_1182 (O_1182,N_14323,N_14849);
or UO_1183 (O_1183,N_14844,N_14486);
nand UO_1184 (O_1184,N_14619,N_14819);
nor UO_1185 (O_1185,N_14631,N_14907);
and UO_1186 (O_1186,N_14352,N_14263);
nor UO_1187 (O_1187,N_14832,N_14911);
or UO_1188 (O_1188,N_14483,N_14450);
nand UO_1189 (O_1189,N_14918,N_14449);
and UO_1190 (O_1190,N_14984,N_14603);
nand UO_1191 (O_1191,N_14596,N_14720);
and UO_1192 (O_1192,N_14883,N_14876);
nor UO_1193 (O_1193,N_14521,N_14905);
xor UO_1194 (O_1194,N_14879,N_14829);
nand UO_1195 (O_1195,N_14555,N_14686);
or UO_1196 (O_1196,N_14372,N_14797);
and UO_1197 (O_1197,N_14953,N_14284);
and UO_1198 (O_1198,N_14718,N_14463);
nor UO_1199 (O_1199,N_14781,N_14448);
xor UO_1200 (O_1200,N_14376,N_14983);
nand UO_1201 (O_1201,N_14290,N_14796);
nor UO_1202 (O_1202,N_14664,N_14987);
and UO_1203 (O_1203,N_14714,N_14974);
nand UO_1204 (O_1204,N_14484,N_14741);
or UO_1205 (O_1205,N_14620,N_14698);
nor UO_1206 (O_1206,N_14429,N_14695);
xnor UO_1207 (O_1207,N_14268,N_14295);
xor UO_1208 (O_1208,N_14476,N_14377);
or UO_1209 (O_1209,N_14253,N_14936);
nand UO_1210 (O_1210,N_14654,N_14716);
and UO_1211 (O_1211,N_14426,N_14553);
or UO_1212 (O_1212,N_14693,N_14965);
nor UO_1213 (O_1213,N_14962,N_14282);
xor UO_1214 (O_1214,N_14967,N_14764);
and UO_1215 (O_1215,N_14963,N_14305);
nor UO_1216 (O_1216,N_14489,N_14898);
and UO_1217 (O_1217,N_14873,N_14987);
nor UO_1218 (O_1218,N_14772,N_14273);
or UO_1219 (O_1219,N_14927,N_14446);
nand UO_1220 (O_1220,N_14997,N_14581);
nand UO_1221 (O_1221,N_14390,N_14526);
or UO_1222 (O_1222,N_14595,N_14307);
or UO_1223 (O_1223,N_14815,N_14516);
and UO_1224 (O_1224,N_14623,N_14687);
and UO_1225 (O_1225,N_14537,N_14547);
xnor UO_1226 (O_1226,N_14299,N_14763);
or UO_1227 (O_1227,N_14382,N_14437);
or UO_1228 (O_1228,N_14730,N_14942);
nor UO_1229 (O_1229,N_14942,N_14394);
nor UO_1230 (O_1230,N_14510,N_14775);
or UO_1231 (O_1231,N_14397,N_14617);
nor UO_1232 (O_1232,N_14568,N_14945);
and UO_1233 (O_1233,N_14615,N_14737);
nor UO_1234 (O_1234,N_14389,N_14397);
and UO_1235 (O_1235,N_14379,N_14676);
xnor UO_1236 (O_1236,N_14419,N_14936);
nand UO_1237 (O_1237,N_14790,N_14935);
nand UO_1238 (O_1238,N_14725,N_14716);
xor UO_1239 (O_1239,N_14270,N_14264);
xnor UO_1240 (O_1240,N_14914,N_14595);
or UO_1241 (O_1241,N_14564,N_14909);
nor UO_1242 (O_1242,N_14549,N_14668);
nor UO_1243 (O_1243,N_14525,N_14611);
xnor UO_1244 (O_1244,N_14419,N_14503);
nor UO_1245 (O_1245,N_14958,N_14435);
and UO_1246 (O_1246,N_14808,N_14709);
or UO_1247 (O_1247,N_14331,N_14966);
nor UO_1248 (O_1248,N_14467,N_14877);
nand UO_1249 (O_1249,N_14820,N_14516);
or UO_1250 (O_1250,N_14989,N_14632);
nor UO_1251 (O_1251,N_14586,N_14402);
nor UO_1252 (O_1252,N_14505,N_14630);
nor UO_1253 (O_1253,N_14738,N_14836);
or UO_1254 (O_1254,N_14535,N_14628);
or UO_1255 (O_1255,N_14630,N_14590);
and UO_1256 (O_1256,N_14449,N_14610);
xor UO_1257 (O_1257,N_14932,N_14251);
nor UO_1258 (O_1258,N_14959,N_14536);
and UO_1259 (O_1259,N_14998,N_14280);
or UO_1260 (O_1260,N_14494,N_14659);
nand UO_1261 (O_1261,N_14299,N_14493);
and UO_1262 (O_1262,N_14751,N_14951);
or UO_1263 (O_1263,N_14403,N_14360);
nand UO_1264 (O_1264,N_14568,N_14772);
and UO_1265 (O_1265,N_14633,N_14536);
and UO_1266 (O_1266,N_14494,N_14582);
nand UO_1267 (O_1267,N_14741,N_14271);
nor UO_1268 (O_1268,N_14421,N_14281);
nor UO_1269 (O_1269,N_14474,N_14905);
and UO_1270 (O_1270,N_14752,N_14302);
nand UO_1271 (O_1271,N_14839,N_14970);
nand UO_1272 (O_1272,N_14787,N_14448);
nand UO_1273 (O_1273,N_14525,N_14746);
nand UO_1274 (O_1274,N_14885,N_14863);
nand UO_1275 (O_1275,N_14955,N_14475);
nand UO_1276 (O_1276,N_14981,N_14790);
and UO_1277 (O_1277,N_14441,N_14600);
and UO_1278 (O_1278,N_14806,N_14282);
xnor UO_1279 (O_1279,N_14864,N_14521);
xnor UO_1280 (O_1280,N_14596,N_14614);
nand UO_1281 (O_1281,N_14851,N_14313);
nand UO_1282 (O_1282,N_14552,N_14665);
xnor UO_1283 (O_1283,N_14336,N_14994);
and UO_1284 (O_1284,N_14577,N_14580);
and UO_1285 (O_1285,N_14859,N_14796);
nand UO_1286 (O_1286,N_14804,N_14825);
and UO_1287 (O_1287,N_14399,N_14797);
nand UO_1288 (O_1288,N_14978,N_14888);
nand UO_1289 (O_1289,N_14627,N_14965);
or UO_1290 (O_1290,N_14710,N_14781);
nand UO_1291 (O_1291,N_14732,N_14412);
or UO_1292 (O_1292,N_14978,N_14405);
nand UO_1293 (O_1293,N_14965,N_14651);
nor UO_1294 (O_1294,N_14326,N_14918);
and UO_1295 (O_1295,N_14931,N_14498);
or UO_1296 (O_1296,N_14996,N_14468);
nor UO_1297 (O_1297,N_14614,N_14484);
xor UO_1298 (O_1298,N_14661,N_14259);
xnor UO_1299 (O_1299,N_14260,N_14278);
nand UO_1300 (O_1300,N_14735,N_14466);
or UO_1301 (O_1301,N_14293,N_14575);
and UO_1302 (O_1302,N_14625,N_14453);
and UO_1303 (O_1303,N_14884,N_14959);
or UO_1304 (O_1304,N_14720,N_14554);
nor UO_1305 (O_1305,N_14775,N_14465);
nand UO_1306 (O_1306,N_14994,N_14722);
nor UO_1307 (O_1307,N_14995,N_14508);
nand UO_1308 (O_1308,N_14782,N_14280);
xor UO_1309 (O_1309,N_14500,N_14843);
or UO_1310 (O_1310,N_14915,N_14379);
xor UO_1311 (O_1311,N_14713,N_14441);
and UO_1312 (O_1312,N_14761,N_14412);
or UO_1313 (O_1313,N_14809,N_14270);
nand UO_1314 (O_1314,N_14482,N_14859);
and UO_1315 (O_1315,N_14582,N_14271);
nor UO_1316 (O_1316,N_14691,N_14391);
or UO_1317 (O_1317,N_14320,N_14591);
nor UO_1318 (O_1318,N_14968,N_14710);
nor UO_1319 (O_1319,N_14873,N_14332);
or UO_1320 (O_1320,N_14356,N_14844);
nand UO_1321 (O_1321,N_14911,N_14731);
or UO_1322 (O_1322,N_14808,N_14513);
or UO_1323 (O_1323,N_14584,N_14862);
or UO_1324 (O_1324,N_14933,N_14863);
and UO_1325 (O_1325,N_14434,N_14375);
and UO_1326 (O_1326,N_14897,N_14899);
nor UO_1327 (O_1327,N_14466,N_14544);
nand UO_1328 (O_1328,N_14841,N_14684);
nor UO_1329 (O_1329,N_14829,N_14604);
nor UO_1330 (O_1330,N_14426,N_14332);
or UO_1331 (O_1331,N_14453,N_14556);
nor UO_1332 (O_1332,N_14585,N_14338);
nand UO_1333 (O_1333,N_14824,N_14755);
xnor UO_1334 (O_1334,N_14305,N_14287);
nand UO_1335 (O_1335,N_14973,N_14937);
or UO_1336 (O_1336,N_14900,N_14794);
nor UO_1337 (O_1337,N_14780,N_14384);
nand UO_1338 (O_1338,N_14664,N_14787);
and UO_1339 (O_1339,N_14882,N_14386);
and UO_1340 (O_1340,N_14629,N_14797);
and UO_1341 (O_1341,N_14727,N_14451);
nand UO_1342 (O_1342,N_14857,N_14411);
and UO_1343 (O_1343,N_14588,N_14544);
and UO_1344 (O_1344,N_14743,N_14514);
nand UO_1345 (O_1345,N_14689,N_14400);
nand UO_1346 (O_1346,N_14550,N_14648);
nor UO_1347 (O_1347,N_14967,N_14555);
nor UO_1348 (O_1348,N_14914,N_14298);
and UO_1349 (O_1349,N_14306,N_14940);
or UO_1350 (O_1350,N_14507,N_14615);
nor UO_1351 (O_1351,N_14710,N_14790);
nor UO_1352 (O_1352,N_14985,N_14481);
or UO_1353 (O_1353,N_14755,N_14628);
or UO_1354 (O_1354,N_14654,N_14328);
nor UO_1355 (O_1355,N_14708,N_14676);
nand UO_1356 (O_1356,N_14562,N_14499);
or UO_1357 (O_1357,N_14871,N_14270);
nor UO_1358 (O_1358,N_14478,N_14307);
nor UO_1359 (O_1359,N_14891,N_14459);
and UO_1360 (O_1360,N_14613,N_14696);
xnor UO_1361 (O_1361,N_14345,N_14388);
and UO_1362 (O_1362,N_14485,N_14738);
nor UO_1363 (O_1363,N_14834,N_14677);
nand UO_1364 (O_1364,N_14513,N_14877);
nand UO_1365 (O_1365,N_14407,N_14790);
or UO_1366 (O_1366,N_14282,N_14322);
nand UO_1367 (O_1367,N_14794,N_14568);
or UO_1368 (O_1368,N_14852,N_14797);
xor UO_1369 (O_1369,N_14761,N_14870);
nor UO_1370 (O_1370,N_14413,N_14799);
and UO_1371 (O_1371,N_14721,N_14740);
nor UO_1372 (O_1372,N_14776,N_14869);
nor UO_1373 (O_1373,N_14598,N_14577);
xnor UO_1374 (O_1374,N_14735,N_14358);
nor UO_1375 (O_1375,N_14955,N_14314);
or UO_1376 (O_1376,N_14374,N_14653);
nand UO_1377 (O_1377,N_14733,N_14454);
and UO_1378 (O_1378,N_14756,N_14711);
nand UO_1379 (O_1379,N_14279,N_14580);
nand UO_1380 (O_1380,N_14488,N_14740);
nand UO_1381 (O_1381,N_14680,N_14930);
nor UO_1382 (O_1382,N_14897,N_14392);
and UO_1383 (O_1383,N_14872,N_14318);
xor UO_1384 (O_1384,N_14343,N_14911);
nand UO_1385 (O_1385,N_14821,N_14593);
nand UO_1386 (O_1386,N_14831,N_14495);
nor UO_1387 (O_1387,N_14401,N_14595);
nand UO_1388 (O_1388,N_14850,N_14404);
nand UO_1389 (O_1389,N_14920,N_14861);
or UO_1390 (O_1390,N_14916,N_14277);
nand UO_1391 (O_1391,N_14473,N_14341);
or UO_1392 (O_1392,N_14551,N_14608);
nand UO_1393 (O_1393,N_14561,N_14468);
nor UO_1394 (O_1394,N_14331,N_14553);
and UO_1395 (O_1395,N_14526,N_14540);
nand UO_1396 (O_1396,N_14590,N_14360);
or UO_1397 (O_1397,N_14339,N_14549);
nand UO_1398 (O_1398,N_14641,N_14386);
nand UO_1399 (O_1399,N_14499,N_14864);
nor UO_1400 (O_1400,N_14440,N_14433);
xor UO_1401 (O_1401,N_14687,N_14327);
nand UO_1402 (O_1402,N_14910,N_14437);
nor UO_1403 (O_1403,N_14344,N_14767);
nor UO_1404 (O_1404,N_14612,N_14365);
xnor UO_1405 (O_1405,N_14401,N_14764);
and UO_1406 (O_1406,N_14672,N_14936);
xnor UO_1407 (O_1407,N_14257,N_14793);
nor UO_1408 (O_1408,N_14347,N_14420);
and UO_1409 (O_1409,N_14279,N_14283);
nor UO_1410 (O_1410,N_14352,N_14816);
nor UO_1411 (O_1411,N_14503,N_14270);
and UO_1412 (O_1412,N_14845,N_14463);
nand UO_1413 (O_1413,N_14278,N_14908);
nand UO_1414 (O_1414,N_14407,N_14399);
and UO_1415 (O_1415,N_14532,N_14802);
nand UO_1416 (O_1416,N_14421,N_14883);
and UO_1417 (O_1417,N_14425,N_14958);
and UO_1418 (O_1418,N_14627,N_14861);
nand UO_1419 (O_1419,N_14578,N_14300);
or UO_1420 (O_1420,N_14681,N_14701);
or UO_1421 (O_1421,N_14999,N_14550);
nand UO_1422 (O_1422,N_14487,N_14755);
nand UO_1423 (O_1423,N_14250,N_14502);
and UO_1424 (O_1424,N_14688,N_14726);
or UO_1425 (O_1425,N_14382,N_14434);
or UO_1426 (O_1426,N_14683,N_14730);
xnor UO_1427 (O_1427,N_14909,N_14996);
nand UO_1428 (O_1428,N_14904,N_14842);
xor UO_1429 (O_1429,N_14340,N_14990);
xnor UO_1430 (O_1430,N_14831,N_14701);
and UO_1431 (O_1431,N_14755,N_14344);
xnor UO_1432 (O_1432,N_14275,N_14271);
nor UO_1433 (O_1433,N_14591,N_14730);
xor UO_1434 (O_1434,N_14792,N_14565);
and UO_1435 (O_1435,N_14584,N_14421);
and UO_1436 (O_1436,N_14646,N_14760);
and UO_1437 (O_1437,N_14938,N_14647);
or UO_1438 (O_1438,N_14860,N_14943);
nor UO_1439 (O_1439,N_14909,N_14925);
nor UO_1440 (O_1440,N_14437,N_14568);
or UO_1441 (O_1441,N_14673,N_14375);
and UO_1442 (O_1442,N_14993,N_14758);
and UO_1443 (O_1443,N_14823,N_14372);
nor UO_1444 (O_1444,N_14608,N_14569);
and UO_1445 (O_1445,N_14934,N_14692);
xor UO_1446 (O_1446,N_14718,N_14281);
and UO_1447 (O_1447,N_14699,N_14611);
or UO_1448 (O_1448,N_14944,N_14613);
xor UO_1449 (O_1449,N_14283,N_14329);
or UO_1450 (O_1450,N_14356,N_14970);
and UO_1451 (O_1451,N_14611,N_14564);
nor UO_1452 (O_1452,N_14650,N_14359);
nand UO_1453 (O_1453,N_14549,N_14682);
or UO_1454 (O_1454,N_14447,N_14397);
nand UO_1455 (O_1455,N_14725,N_14801);
nor UO_1456 (O_1456,N_14689,N_14637);
or UO_1457 (O_1457,N_14406,N_14567);
and UO_1458 (O_1458,N_14590,N_14411);
nor UO_1459 (O_1459,N_14978,N_14410);
and UO_1460 (O_1460,N_14256,N_14483);
nand UO_1461 (O_1461,N_14598,N_14779);
or UO_1462 (O_1462,N_14614,N_14984);
or UO_1463 (O_1463,N_14842,N_14455);
or UO_1464 (O_1464,N_14857,N_14727);
and UO_1465 (O_1465,N_14295,N_14434);
nor UO_1466 (O_1466,N_14263,N_14876);
or UO_1467 (O_1467,N_14373,N_14404);
nor UO_1468 (O_1468,N_14701,N_14691);
and UO_1469 (O_1469,N_14650,N_14632);
xnor UO_1470 (O_1470,N_14708,N_14409);
nand UO_1471 (O_1471,N_14779,N_14564);
nor UO_1472 (O_1472,N_14477,N_14703);
nor UO_1473 (O_1473,N_14788,N_14421);
and UO_1474 (O_1474,N_14253,N_14473);
and UO_1475 (O_1475,N_14950,N_14402);
and UO_1476 (O_1476,N_14323,N_14504);
nand UO_1477 (O_1477,N_14998,N_14579);
or UO_1478 (O_1478,N_14661,N_14824);
and UO_1479 (O_1479,N_14860,N_14366);
and UO_1480 (O_1480,N_14981,N_14514);
xnor UO_1481 (O_1481,N_14334,N_14954);
nand UO_1482 (O_1482,N_14562,N_14340);
nand UO_1483 (O_1483,N_14623,N_14848);
nor UO_1484 (O_1484,N_14850,N_14296);
and UO_1485 (O_1485,N_14494,N_14419);
nand UO_1486 (O_1486,N_14618,N_14541);
nand UO_1487 (O_1487,N_14919,N_14307);
nor UO_1488 (O_1488,N_14630,N_14840);
or UO_1489 (O_1489,N_14256,N_14928);
and UO_1490 (O_1490,N_14902,N_14515);
xor UO_1491 (O_1491,N_14696,N_14783);
nor UO_1492 (O_1492,N_14792,N_14712);
nor UO_1493 (O_1493,N_14455,N_14943);
and UO_1494 (O_1494,N_14687,N_14307);
xor UO_1495 (O_1495,N_14748,N_14978);
nor UO_1496 (O_1496,N_14329,N_14921);
nor UO_1497 (O_1497,N_14814,N_14389);
and UO_1498 (O_1498,N_14730,N_14385);
or UO_1499 (O_1499,N_14702,N_14327);
or UO_1500 (O_1500,N_14374,N_14743);
or UO_1501 (O_1501,N_14339,N_14772);
nor UO_1502 (O_1502,N_14588,N_14631);
nand UO_1503 (O_1503,N_14559,N_14653);
or UO_1504 (O_1504,N_14717,N_14575);
nand UO_1505 (O_1505,N_14581,N_14616);
and UO_1506 (O_1506,N_14439,N_14328);
and UO_1507 (O_1507,N_14423,N_14507);
nand UO_1508 (O_1508,N_14938,N_14683);
and UO_1509 (O_1509,N_14876,N_14831);
nand UO_1510 (O_1510,N_14473,N_14339);
or UO_1511 (O_1511,N_14254,N_14729);
nand UO_1512 (O_1512,N_14510,N_14923);
and UO_1513 (O_1513,N_14690,N_14850);
nor UO_1514 (O_1514,N_14737,N_14336);
or UO_1515 (O_1515,N_14385,N_14899);
and UO_1516 (O_1516,N_14262,N_14299);
and UO_1517 (O_1517,N_14268,N_14449);
nand UO_1518 (O_1518,N_14716,N_14890);
or UO_1519 (O_1519,N_14790,N_14621);
nor UO_1520 (O_1520,N_14790,N_14300);
nor UO_1521 (O_1521,N_14787,N_14413);
and UO_1522 (O_1522,N_14584,N_14949);
and UO_1523 (O_1523,N_14534,N_14619);
or UO_1524 (O_1524,N_14488,N_14750);
nand UO_1525 (O_1525,N_14748,N_14258);
or UO_1526 (O_1526,N_14473,N_14586);
and UO_1527 (O_1527,N_14950,N_14641);
xnor UO_1528 (O_1528,N_14311,N_14669);
and UO_1529 (O_1529,N_14404,N_14807);
nand UO_1530 (O_1530,N_14837,N_14466);
and UO_1531 (O_1531,N_14273,N_14998);
and UO_1532 (O_1532,N_14578,N_14935);
or UO_1533 (O_1533,N_14970,N_14371);
nand UO_1534 (O_1534,N_14771,N_14743);
nand UO_1535 (O_1535,N_14797,N_14374);
nand UO_1536 (O_1536,N_14788,N_14955);
xor UO_1537 (O_1537,N_14255,N_14286);
and UO_1538 (O_1538,N_14710,N_14463);
xnor UO_1539 (O_1539,N_14578,N_14901);
or UO_1540 (O_1540,N_14879,N_14887);
and UO_1541 (O_1541,N_14414,N_14667);
nand UO_1542 (O_1542,N_14556,N_14459);
and UO_1543 (O_1543,N_14841,N_14402);
nor UO_1544 (O_1544,N_14770,N_14892);
and UO_1545 (O_1545,N_14511,N_14762);
or UO_1546 (O_1546,N_14704,N_14778);
nor UO_1547 (O_1547,N_14579,N_14259);
nand UO_1548 (O_1548,N_14905,N_14499);
or UO_1549 (O_1549,N_14597,N_14348);
or UO_1550 (O_1550,N_14474,N_14802);
nor UO_1551 (O_1551,N_14728,N_14494);
xnor UO_1552 (O_1552,N_14756,N_14798);
or UO_1553 (O_1553,N_14863,N_14433);
or UO_1554 (O_1554,N_14743,N_14726);
and UO_1555 (O_1555,N_14396,N_14832);
nand UO_1556 (O_1556,N_14462,N_14910);
nor UO_1557 (O_1557,N_14709,N_14787);
nand UO_1558 (O_1558,N_14972,N_14607);
nor UO_1559 (O_1559,N_14948,N_14260);
and UO_1560 (O_1560,N_14488,N_14972);
or UO_1561 (O_1561,N_14278,N_14358);
nor UO_1562 (O_1562,N_14761,N_14686);
or UO_1563 (O_1563,N_14869,N_14334);
or UO_1564 (O_1564,N_14592,N_14491);
nand UO_1565 (O_1565,N_14913,N_14911);
and UO_1566 (O_1566,N_14825,N_14369);
nor UO_1567 (O_1567,N_14843,N_14705);
nor UO_1568 (O_1568,N_14607,N_14563);
and UO_1569 (O_1569,N_14441,N_14620);
nor UO_1570 (O_1570,N_14487,N_14276);
nand UO_1571 (O_1571,N_14643,N_14375);
or UO_1572 (O_1572,N_14775,N_14883);
nand UO_1573 (O_1573,N_14490,N_14745);
and UO_1574 (O_1574,N_14505,N_14755);
or UO_1575 (O_1575,N_14443,N_14874);
nand UO_1576 (O_1576,N_14967,N_14626);
and UO_1577 (O_1577,N_14785,N_14989);
or UO_1578 (O_1578,N_14317,N_14625);
nand UO_1579 (O_1579,N_14511,N_14267);
xnor UO_1580 (O_1580,N_14301,N_14719);
and UO_1581 (O_1581,N_14285,N_14852);
nor UO_1582 (O_1582,N_14964,N_14829);
nand UO_1583 (O_1583,N_14341,N_14905);
nand UO_1584 (O_1584,N_14958,N_14540);
and UO_1585 (O_1585,N_14657,N_14385);
nand UO_1586 (O_1586,N_14975,N_14919);
nor UO_1587 (O_1587,N_14650,N_14304);
or UO_1588 (O_1588,N_14661,N_14281);
nor UO_1589 (O_1589,N_14996,N_14870);
nand UO_1590 (O_1590,N_14966,N_14830);
nor UO_1591 (O_1591,N_14724,N_14860);
or UO_1592 (O_1592,N_14466,N_14750);
and UO_1593 (O_1593,N_14510,N_14353);
and UO_1594 (O_1594,N_14266,N_14918);
nand UO_1595 (O_1595,N_14257,N_14976);
or UO_1596 (O_1596,N_14814,N_14804);
nand UO_1597 (O_1597,N_14315,N_14370);
or UO_1598 (O_1598,N_14855,N_14958);
or UO_1599 (O_1599,N_14715,N_14811);
nor UO_1600 (O_1600,N_14892,N_14444);
nor UO_1601 (O_1601,N_14875,N_14348);
xnor UO_1602 (O_1602,N_14356,N_14355);
nor UO_1603 (O_1603,N_14325,N_14832);
or UO_1604 (O_1604,N_14407,N_14672);
and UO_1605 (O_1605,N_14405,N_14878);
xnor UO_1606 (O_1606,N_14495,N_14895);
nand UO_1607 (O_1607,N_14331,N_14339);
and UO_1608 (O_1608,N_14414,N_14495);
and UO_1609 (O_1609,N_14330,N_14275);
nand UO_1610 (O_1610,N_14275,N_14784);
nor UO_1611 (O_1611,N_14436,N_14386);
nor UO_1612 (O_1612,N_14740,N_14902);
or UO_1613 (O_1613,N_14458,N_14821);
nor UO_1614 (O_1614,N_14769,N_14328);
nand UO_1615 (O_1615,N_14929,N_14281);
nand UO_1616 (O_1616,N_14315,N_14776);
nor UO_1617 (O_1617,N_14467,N_14352);
or UO_1618 (O_1618,N_14379,N_14772);
and UO_1619 (O_1619,N_14773,N_14879);
nand UO_1620 (O_1620,N_14347,N_14398);
nor UO_1621 (O_1621,N_14668,N_14712);
nor UO_1622 (O_1622,N_14447,N_14688);
nor UO_1623 (O_1623,N_14619,N_14775);
or UO_1624 (O_1624,N_14480,N_14370);
xnor UO_1625 (O_1625,N_14917,N_14276);
nand UO_1626 (O_1626,N_14591,N_14560);
xor UO_1627 (O_1627,N_14528,N_14832);
nor UO_1628 (O_1628,N_14761,N_14714);
nand UO_1629 (O_1629,N_14512,N_14257);
nand UO_1630 (O_1630,N_14893,N_14617);
or UO_1631 (O_1631,N_14855,N_14574);
and UO_1632 (O_1632,N_14711,N_14336);
or UO_1633 (O_1633,N_14319,N_14866);
and UO_1634 (O_1634,N_14317,N_14519);
or UO_1635 (O_1635,N_14364,N_14759);
or UO_1636 (O_1636,N_14836,N_14463);
nand UO_1637 (O_1637,N_14419,N_14735);
or UO_1638 (O_1638,N_14578,N_14823);
nand UO_1639 (O_1639,N_14577,N_14948);
and UO_1640 (O_1640,N_14912,N_14301);
or UO_1641 (O_1641,N_14674,N_14440);
nand UO_1642 (O_1642,N_14666,N_14391);
nor UO_1643 (O_1643,N_14333,N_14671);
or UO_1644 (O_1644,N_14587,N_14349);
or UO_1645 (O_1645,N_14943,N_14497);
nand UO_1646 (O_1646,N_14305,N_14787);
nor UO_1647 (O_1647,N_14637,N_14511);
nor UO_1648 (O_1648,N_14904,N_14410);
or UO_1649 (O_1649,N_14293,N_14888);
nor UO_1650 (O_1650,N_14411,N_14268);
or UO_1651 (O_1651,N_14440,N_14331);
nand UO_1652 (O_1652,N_14684,N_14772);
nand UO_1653 (O_1653,N_14579,N_14307);
or UO_1654 (O_1654,N_14936,N_14571);
nor UO_1655 (O_1655,N_14261,N_14934);
and UO_1656 (O_1656,N_14917,N_14777);
and UO_1657 (O_1657,N_14810,N_14511);
or UO_1658 (O_1658,N_14451,N_14687);
xnor UO_1659 (O_1659,N_14724,N_14655);
nand UO_1660 (O_1660,N_14494,N_14930);
or UO_1661 (O_1661,N_14757,N_14920);
or UO_1662 (O_1662,N_14790,N_14681);
or UO_1663 (O_1663,N_14506,N_14706);
and UO_1664 (O_1664,N_14348,N_14549);
nand UO_1665 (O_1665,N_14972,N_14675);
nor UO_1666 (O_1666,N_14963,N_14752);
nand UO_1667 (O_1667,N_14761,N_14403);
and UO_1668 (O_1668,N_14843,N_14932);
nor UO_1669 (O_1669,N_14393,N_14650);
nand UO_1670 (O_1670,N_14354,N_14706);
nor UO_1671 (O_1671,N_14274,N_14808);
and UO_1672 (O_1672,N_14840,N_14495);
and UO_1673 (O_1673,N_14416,N_14993);
or UO_1674 (O_1674,N_14469,N_14258);
or UO_1675 (O_1675,N_14830,N_14342);
nand UO_1676 (O_1676,N_14715,N_14549);
nand UO_1677 (O_1677,N_14599,N_14465);
nor UO_1678 (O_1678,N_14532,N_14694);
nor UO_1679 (O_1679,N_14705,N_14619);
nand UO_1680 (O_1680,N_14548,N_14795);
nand UO_1681 (O_1681,N_14333,N_14800);
and UO_1682 (O_1682,N_14654,N_14251);
nor UO_1683 (O_1683,N_14323,N_14861);
nand UO_1684 (O_1684,N_14950,N_14579);
or UO_1685 (O_1685,N_14606,N_14268);
and UO_1686 (O_1686,N_14938,N_14398);
and UO_1687 (O_1687,N_14964,N_14652);
or UO_1688 (O_1688,N_14931,N_14662);
or UO_1689 (O_1689,N_14915,N_14547);
nand UO_1690 (O_1690,N_14325,N_14369);
nor UO_1691 (O_1691,N_14879,N_14492);
nand UO_1692 (O_1692,N_14992,N_14713);
and UO_1693 (O_1693,N_14709,N_14988);
and UO_1694 (O_1694,N_14491,N_14562);
nand UO_1695 (O_1695,N_14406,N_14949);
nor UO_1696 (O_1696,N_14471,N_14746);
and UO_1697 (O_1697,N_14389,N_14269);
nor UO_1698 (O_1698,N_14511,N_14332);
xor UO_1699 (O_1699,N_14970,N_14716);
and UO_1700 (O_1700,N_14945,N_14969);
or UO_1701 (O_1701,N_14616,N_14878);
nor UO_1702 (O_1702,N_14744,N_14849);
nor UO_1703 (O_1703,N_14527,N_14586);
nand UO_1704 (O_1704,N_14906,N_14401);
or UO_1705 (O_1705,N_14923,N_14863);
and UO_1706 (O_1706,N_14738,N_14314);
nor UO_1707 (O_1707,N_14807,N_14909);
nor UO_1708 (O_1708,N_14411,N_14335);
or UO_1709 (O_1709,N_14452,N_14588);
nor UO_1710 (O_1710,N_14828,N_14570);
or UO_1711 (O_1711,N_14534,N_14815);
and UO_1712 (O_1712,N_14772,N_14495);
nand UO_1713 (O_1713,N_14899,N_14987);
and UO_1714 (O_1714,N_14908,N_14411);
nor UO_1715 (O_1715,N_14286,N_14972);
or UO_1716 (O_1716,N_14981,N_14832);
or UO_1717 (O_1717,N_14815,N_14271);
nor UO_1718 (O_1718,N_14982,N_14398);
nand UO_1719 (O_1719,N_14976,N_14604);
nor UO_1720 (O_1720,N_14384,N_14805);
xor UO_1721 (O_1721,N_14773,N_14256);
and UO_1722 (O_1722,N_14553,N_14816);
nor UO_1723 (O_1723,N_14463,N_14496);
or UO_1724 (O_1724,N_14423,N_14757);
and UO_1725 (O_1725,N_14752,N_14700);
nor UO_1726 (O_1726,N_14735,N_14406);
nor UO_1727 (O_1727,N_14480,N_14845);
and UO_1728 (O_1728,N_14991,N_14684);
nand UO_1729 (O_1729,N_14590,N_14733);
or UO_1730 (O_1730,N_14580,N_14933);
and UO_1731 (O_1731,N_14891,N_14779);
and UO_1732 (O_1732,N_14315,N_14403);
nor UO_1733 (O_1733,N_14669,N_14683);
nor UO_1734 (O_1734,N_14766,N_14749);
and UO_1735 (O_1735,N_14722,N_14694);
nand UO_1736 (O_1736,N_14268,N_14518);
nand UO_1737 (O_1737,N_14712,N_14294);
nor UO_1738 (O_1738,N_14778,N_14718);
or UO_1739 (O_1739,N_14802,N_14625);
and UO_1740 (O_1740,N_14687,N_14570);
nor UO_1741 (O_1741,N_14875,N_14933);
nand UO_1742 (O_1742,N_14379,N_14387);
nor UO_1743 (O_1743,N_14792,N_14459);
nor UO_1744 (O_1744,N_14957,N_14448);
xor UO_1745 (O_1745,N_14779,N_14282);
nor UO_1746 (O_1746,N_14431,N_14581);
xor UO_1747 (O_1747,N_14467,N_14321);
xnor UO_1748 (O_1748,N_14786,N_14417);
nand UO_1749 (O_1749,N_14274,N_14709);
nand UO_1750 (O_1750,N_14395,N_14436);
nor UO_1751 (O_1751,N_14917,N_14632);
or UO_1752 (O_1752,N_14524,N_14426);
nand UO_1753 (O_1753,N_14341,N_14887);
and UO_1754 (O_1754,N_14795,N_14802);
nand UO_1755 (O_1755,N_14846,N_14910);
or UO_1756 (O_1756,N_14475,N_14301);
nand UO_1757 (O_1757,N_14361,N_14812);
nand UO_1758 (O_1758,N_14410,N_14498);
and UO_1759 (O_1759,N_14906,N_14995);
nor UO_1760 (O_1760,N_14716,N_14447);
or UO_1761 (O_1761,N_14633,N_14320);
nor UO_1762 (O_1762,N_14873,N_14571);
or UO_1763 (O_1763,N_14503,N_14434);
nand UO_1764 (O_1764,N_14935,N_14508);
xor UO_1765 (O_1765,N_14800,N_14806);
nor UO_1766 (O_1766,N_14416,N_14895);
nor UO_1767 (O_1767,N_14449,N_14882);
or UO_1768 (O_1768,N_14672,N_14394);
nor UO_1769 (O_1769,N_14746,N_14663);
nand UO_1770 (O_1770,N_14618,N_14958);
nor UO_1771 (O_1771,N_14281,N_14713);
or UO_1772 (O_1772,N_14553,N_14620);
or UO_1773 (O_1773,N_14726,N_14303);
or UO_1774 (O_1774,N_14607,N_14740);
or UO_1775 (O_1775,N_14842,N_14828);
nor UO_1776 (O_1776,N_14344,N_14676);
and UO_1777 (O_1777,N_14654,N_14434);
xnor UO_1778 (O_1778,N_14848,N_14466);
or UO_1779 (O_1779,N_14731,N_14979);
or UO_1780 (O_1780,N_14970,N_14899);
xnor UO_1781 (O_1781,N_14549,N_14486);
and UO_1782 (O_1782,N_14743,N_14458);
and UO_1783 (O_1783,N_14564,N_14699);
nand UO_1784 (O_1784,N_14991,N_14488);
nand UO_1785 (O_1785,N_14875,N_14734);
nand UO_1786 (O_1786,N_14632,N_14682);
nor UO_1787 (O_1787,N_14852,N_14795);
and UO_1788 (O_1788,N_14870,N_14451);
or UO_1789 (O_1789,N_14926,N_14889);
and UO_1790 (O_1790,N_14922,N_14919);
and UO_1791 (O_1791,N_14944,N_14607);
nand UO_1792 (O_1792,N_14767,N_14980);
or UO_1793 (O_1793,N_14641,N_14582);
or UO_1794 (O_1794,N_14443,N_14704);
nand UO_1795 (O_1795,N_14887,N_14575);
or UO_1796 (O_1796,N_14878,N_14460);
xnor UO_1797 (O_1797,N_14962,N_14757);
or UO_1798 (O_1798,N_14694,N_14329);
xnor UO_1799 (O_1799,N_14384,N_14907);
or UO_1800 (O_1800,N_14856,N_14622);
and UO_1801 (O_1801,N_14337,N_14614);
and UO_1802 (O_1802,N_14720,N_14418);
or UO_1803 (O_1803,N_14590,N_14834);
and UO_1804 (O_1804,N_14878,N_14790);
and UO_1805 (O_1805,N_14706,N_14926);
and UO_1806 (O_1806,N_14278,N_14805);
nand UO_1807 (O_1807,N_14474,N_14771);
and UO_1808 (O_1808,N_14833,N_14379);
or UO_1809 (O_1809,N_14378,N_14988);
nand UO_1810 (O_1810,N_14381,N_14364);
nor UO_1811 (O_1811,N_14910,N_14840);
or UO_1812 (O_1812,N_14922,N_14731);
and UO_1813 (O_1813,N_14851,N_14686);
and UO_1814 (O_1814,N_14331,N_14401);
nand UO_1815 (O_1815,N_14415,N_14700);
nand UO_1816 (O_1816,N_14575,N_14557);
or UO_1817 (O_1817,N_14716,N_14372);
or UO_1818 (O_1818,N_14633,N_14931);
and UO_1819 (O_1819,N_14661,N_14624);
and UO_1820 (O_1820,N_14607,N_14745);
nor UO_1821 (O_1821,N_14491,N_14752);
and UO_1822 (O_1822,N_14838,N_14949);
or UO_1823 (O_1823,N_14623,N_14522);
or UO_1824 (O_1824,N_14505,N_14932);
nand UO_1825 (O_1825,N_14709,N_14822);
and UO_1826 (O_1826,N_14812,N_14549);
nor UO_1827 (O_1827,N_14748,N_14510);
xor UO_1828 (O_1828,N_14821,N_14599);
nor UO_1829 (O_1829,N_14763,N_14748);
and UO_1830 (O_1830,N_14406,N_14757);
or UO_1831 (O_1831,N_14412,N_14488);
nand UO_1832 (O_1832,N_14444,N_14565);
xnor UO_1833 (O_1833,N_14446,N_14877);
and UO_1834 (O_1834,N_14766,N_14679);
nand UO_1835 (O_1835,N_14390,N_14290);
nand UO_1836 (O_1836,N_14840,N_14576);
nand UO_1837 (O_1837,N_14994,N_14765);
nand UO_1838 (O_1838,N_14910,N_14914);
nor UO_1839 (O_1839,N_14297,N_14863);
nand UO_1840 (O_1840,N_14892,N_14865);
nand UO_1841 (O_1841,N_14567,N_14620);
and UO_1842 (O_1842,N_14329,N_14825);
and UO_1843 (O_1843,N_14730,N_14978);
and UO_1844 (O_1844,N_14993,N_14914);
xnor UO_1845 (O_1845,N_14292,N_14343);
or UO_1846 (O_1846,N_14418,N_14293);
or UO_1847 (O_1847,N_14915,N_14983);
nand UO_1848 (O_1848,N_14747,N_14681);
nand UO_1849 (O_1849,N_14948,N_14255);
nand UO_1850 (O_1850,N_14349,N_14311);
nor UO_1851 (O_1851,N_14365,N_14440);
nor UO_1852 (O_1852,N_14273,N_14649);
and UO_1853 (O_1853,N_14335,N_14823);
nor UO_1854 (O_1854,N_14720,N_14692);
nor UO_1855 (O_1855,N_14650,N_14850);
or UO_1856 (O_1856,N_14535,N_14897);
or UO_1857 (O_1857,N_14495,N_14957);
nand UO_1858 (O_1858,N_14384,N_14440);
nor UO_1859 (O_1859,N_14760,N_14834);
or UO_1860 (O_1860,N_14292,N_14455);
nand UO_1861 (O_1861,N_14931,N_14295);
and UO_1862 (O_1862,N_14942,N_14770);
or UO_1863 (O_1863,N_14887,N_14568);
nor UO_1864 (O_1864,N_14706,N_14701);
nor UO_1865 (O_1865,N_14276,N_14553);
or UO_1866 (O_1866,N_14636,N_14738);
and UO_1867 (O_1867,N_14538,N_14628);
nor UO_1868 (O_1868,N_14812,N_14627);
and UO_1869 (O_1869,N_14703,N_14341);
nor UO_1870 (O_1870,N_14576,N_14963);
and UO_1871 (O_1871,N_14517,N_14352);
xor UO_1872 (O_1872,N_14781,N_14901);
nand UO_1873 (O_1873,N_14961,N_14593);
and UO_1874 (O_1874,N_14278,N_14529);
nor UO_1875 (O_1875,N_14833,N_14820);
nand UO_1876 (O_1876,N_14541,N_14410);
nand UO_1877 (O_1877,N_14938,N_14947);
nor UO_1878 (O_1878,N_14371,N_14470);
nor UO_1879 (O_1879,N_14785,N_14702);
nor UO_1880 (O_1880,N_14340,N_14250);
nand UO_1881 (O_1881,N_14710,N_14785);
or UO_1882 (O_1882,N_14297,N_14761);
or UO_1883 (O_1883,N_14481,N_14756);
nor UO_1884 (O_1884,N_14479,N_14261);
and UO_1885 (O_1885,N_14667,N_14410);
nor UO_1886 (O_1886,N_14357,N_14667);
nor UO_1887 (O_1887,N_14879,N_14493);
nor UO_1888 (O_1888,N_14475,N_14627);
nor UO_1889 (O_1889,N_14612,N_14481);
xor UO_1890 (O_1890,N_14336,N_14404);
nand UO_1891 (O_1891,N_14738,N_14768);
or UO_1892 (O_1892,N_14756,N_14304);
and UO_1893 (O_1893,N_14818,N_14445);
and UO_1894 (O_1894,N_14258,N_14431);
nor UO_1895 (O_1895,N_14874,N_14533);
nand UO_1896 (O_1896,N_14639,N_14765);
or UO_1897 (O_1897,N_14411,N_14313);
or UO_1898 (O_1898,N_14697,N_14787);
xor UO_1899 (O_1899,N_14946,N_14281);
and UO_1900 (O_1900,N_14972,N_14682);
nand UO_1901 (O_1901,N_14865,N_14543);
xnor UO_1902 (O_1902,N_14499,N_14590);
or UO_1903 (O_1903,N_14692,N_14837);
nand UO_1904 (O_1904,N_14872,N_14647);
or UO_1905 (O_1905,N_14922,N_14437);
or UO_1906 (O_1906,N_14981,N_14474);
or UO_1907 (O_1907,N_14259,N_14666);
nand UO_1908 (O_1908,N_14984,N_14266);
and UO_1909 (O_1909,N_14260,N_14805);
nor UO_1910 (O_1910,N_14651,N_14761);
nor UO_1911 (O_1911,N_14378,N_14831);
and UO_1912 (O_1912,N_14541,N_14621);
or UO_1913 (O_1913,N_14916,N_14403);
and UO_1914 (O_1914,N_14542,N_14639);
nand UO_1915 (O_1915,N_14650,N_14829);
and UO_1916 (O_1916,N_14344,N_14330);
nor UO_1917 (O_1917,N_14338,N_14936);
or UO_1918 (O_1918,N_14296,N_14779);
nand UO_1919 (O_1919,N_14458,N_14475);
and UO_1920 (O_1920,N_14480,N_14630);
nor UO_1921 (O_1921,N_14507,N_14597);
xor UO_1922 (O_1922,N_14470,N_14944);
nor UO_1923 (O_1923,N_14622,N_14411);
or UO_1924 (O_1924,N_14715,N_14737);
nor UO_1925 (O_1925,N_14324,N_14321);
nand UO_1926 (O_1926,N_14511,N_14501);
or UO_1927 (O_1927,N_14420,N_14995);
nor UO_1928 (O_1928,N_14625,N_14393);
or UO_1929 (O_1929,N_14878,N_14993);
or UO_1930 (O_1930,N_14877,N_14478);
nand UO_1931 (O_1931,N_14327,N_14800);
nand UO_1932 (O_1932,N_14276,N_14692);
or UO_1933 (O_1933,N_14688,N_14527);
nor UO_1934 (O_1934,N_14660,N_14293);
or UO_1935 (O_1935,N_14644,N_14374);
nand UO_1936 (O_1936,N_14459,N_14616);
and UO_1937 (O_1937,N_14838,N_14577);
xnor UO_1938 (O_1938,N_14915,N_14797);
nor UO_1939 (O_1939,N_14923,N_14549);
xor UO_1940 (O_1940,N_14515,N_14781);
and UO_1941 (O_1941,N_14518,N_14813);
nor UO_1942 (O_1942,N_14756,N_14677);
nor UO_1943 (O_1943,N_14534,N_14583);
or UO_1944 (O_1944,N_14461,N_14940);
or UO_1945 (O_1945,N_14500,N_14714);
or UO_1946 (O_1946,N_14935,N_14931);
nor UO_1947 (O_1947,N_14344,N_14915);
and UO_1948 (O_1948,N_14943,N_14978);
nor UO_1949 (O_1949,N_14320,N_14778);
nor UO_1950 (O_1950,N_14587,N_14254);
and UO_1951 (O_1951,N_14316,N_14937);
nor UO_1952 (O_1952,N_14901,N_14709);
nor UO_1953 (O_1953,N_14449,N_14977);
and UO_1954 (O_1954,N_14290,N_14448);
nand UO_1955 (O_1955,N_14909,N_14973);
and UO_1956 (O_1956,N_14385,N_14399);
or UO_1957 (O_1957,N_14456,N_14932);
nor UO_1958 (O_1958,N_14677,N_14852);
or UO_1959 (O_1959,N_14387,N_14432);
and UO_1960 (O_1960,N_14784,N_14514);
and UO_1961 (O_1961,N_14673,N_14613);
nor UO_1962 (O_1962,N_14746,N_14974);
nor UO_1963 (O_1963,N_14284,N_14497);
and UO_1964 (O_1964,N_14485,N_14344);
nor UO_1965 (O_1965,N_14803,N_14533);
or UO_1966 (O_1966,N_14469,N_14754);
nand UO_1967 (O_1967,N_14594,N_14983);
xor UO_1968 (O_1968,N_14871,N_14492);
nor UO_1969 (O_1969,N_14563,N_14785);
nand UO_1970 (O_1970,N_14336,N_14786);
and UO_1971 (O_1971,N_14717,N_14436);
nor UO_1972 (O_1972,N_14728,N_14502);
nand UO_1973 (O_1973,N_14385,N_14842);
and UO_1974 (O_1974,N_14802,N_14614);
nor UO_1975 (O_1975,N_14527,N_14795);
or UO_1976 (O_1976,N_14813,N_14672);
nor UO_1977 (O_1977,N_14919,N_14448);
nor UO_1978 (O_1978,N_14284,N_14478);
nor UO_1979 (O_1979,N_14477,N_14377);
nand UO_1980 (O_1980,N_14263,N_14312);
and UO_1981 (O_1981,N_14943,N_14884);
xor UO_1982 (O_1982,N_14276,N_14568);
or UO_1983 (O_1983,N_14356,N_14256);
and UO_1984 (O_1984,N_14396,N_14646);
nand UO_1985 (O_1985,N_14648,N_14282);
and UO_1986 (O_1986,N_14996,N_14345);
or UO_1987 (O_1987,N_14512,N_14850);
and UO_1988 (O_1988,N_14256,N_14283);
or UO_1989 (O_1989,N_14493,N_14372);
or UO_1990 (O_1990,N_14454,N_14366);
nand UO_1991 (O_1991,N_14587,N_14601);
and UO_1992 (O_1992,N_14803,N_14308);
xor UO_1993 (O_1993,N_14734,N_14369);
nand UO_1994 (O_1994,N_14864,N_14734);
nor UO_1995 (O_1995,N_14361,N_14845);
and UO_1996 (O_1996,N_14527,N_14434);
nor UO_1997 (O_1997,N_14398,N_14933);
and UO_1998 (O_1998,N_14919,N_14721);
nor UO_1999 (O_1999,N_14357,N_14724);
endmodule