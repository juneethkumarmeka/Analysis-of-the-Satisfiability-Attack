module basic_500_3000_500_15_levels_1xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_184,In_459);
and U1 (N_1,In_150,In_138);
nand U2 (N_2,In_386,In_30);
nand U3 (N_3,In_497,In_324);
or U4 (N_4,In_6,In_415);
and U5 (N_5,In_132,In_108);
nand U6 (N_6,In_383,In_455);
nor U7 (N_7,In_406,In_261);
or U8 (N_8,In_378,In_14);
nand U9 (N_9,In_338,In_149);
nor U10 (N_10,In_167,In_25);
xor U11 (N_11,In_39,In_279);
nand U12 (N_12,In_281,In_164);
and U13 (N_13,In_487,In_353);
or U14 (N_14,In_152,In_142);
or U15 (N_15,In_8,In_440);
and U16 (N_16,In_436,In_175);
and U17 (N_17,In_450,In_496);
or U18 (N_18,In_79,In_411);
nor U19 (N_19,In_80,In_205);
and U20 (N_20,In_92,In_171);
or U21 (N_21,In_376,In_29);
and U22 (N_22,In_260,In_488);
nand U23 (N_23,In_468,In_412);
nand U24 (N_24,In_162,In_188);
or U25 (N_25,In_443,In_354);
nand U26 (N_26,In_417,In_348);
or U27 (N_27,In_469,In_221);
or U28 (N_28,In_283,In_114);
nand U29 (N_29,In_20,In_262);
nor U30 (N_30,In_356,In_52);
and U31 (N_31,In_256,In_477);
nor U32 (N_32,In_312,In_360);
nor U33 (N_33,In_105,In_75);
or U34 (N_34,In_15,In_264);
nor U35 (N_35,In_151,In_453);
xor U36 (N_36,In_207,In_185);
and U37 (N_37,In_50,In_17);
or U38 (N_38,In_196,In_209);
nand U39 (N_39,In_267,In_115);
and U40 (N_40,In_431,In_27);
nor U41 (N_41,In_282,In_219);
nand U42 (N_42,In_110,In_45);
nor U43 (N_43,In_389,In_339);
and U44 (N_44,In_401,In_350);
nor U45 (N_45,In_367,In_74);
and U46 (N_46,In_212,In_63);
and U47 (N_47,In_374,In_64);
nor U48 (N_48,In_143,In_457);
and U49 (N_49,In_420,In_181);
or U50 (N_50,In_494,In_355);
or U51 (N_51,In_272,In_31);
nand U52 (N_52,In_358,In_93);
nor U53 (N_53,In_315,In_409);
nand U54 (N_54,In_476,In_69);
nor U55 (N_55,In_331,In_271);
and U56 (N_56,In_294,In_357);
and U57 (N_57,In_144,In_439);
nand U58 (N_58,In_435,In_446);
nor U59 (N_59,In_291,In_368);
nor U60 (N_60,In_347,In_90);
nor U61 (N_61,In_273,In_430);
or U62 (N_62,In_301,In_429);
and U63 (N_63,In_22,In_43);
nor U64 (N_64,In_396,In_202);
or U65 (N_65,In_67,In_106);
and U66 (N_66,In_274,In_421);
and U67 (N_67,In_322,In_452);
nand U68 (N_68,In_85,In_183);
or U69 (N_69,In_465,In_55);
nand U70 (N_70,In_266,In_191);
and U71 (N_71,In_329,In_489);
nand U72 (N_72,In_319,In_161);
and U73 (N_73,In_180,In_302);
and U74 (N_74,In_210,In_280);
nor U75 (N_75,In_333,In_133);
and U76 (N_76,In_381,In_449);
or U77 (N_77,In_81,In_37);
nand U78 (N_78,In_466,In_148);
nand U79 (N_79,In_42,In_444);
and U80 (N_80,In_235,In_275);
or U81 (N_81,In_399,In_165);
nor U82 (N_82,In_159,In_117);
and U83 (N_83,In_177,In_438);
or U84 (N_84,In_400,In_134);
nand U85 (N_85,In_458,In_38);
and U86 (N_86,In_427,In_157);
nor U87 (N_87,In_286,In_237);
nand U88 (N_88,In_344,In_491);
and U89 (N_89,In_222,In_326);
nand U90 (N_90,In_451,In_385);
nor U91 (N_91,In_73,In_464);
and U92 (N_92,In_23,In_53);
or U93 (N_93,In_293,In_335);
or U94 (N_94,In_363,In_36);
or U95 (N_95,In_332,In_57);
or U96 (N_96,In_240,In_41);
nand U97 (N_97,In_475,In_220);
and U98 (N_98,In_277,In_352);
or U99 (N_99,In_408,In_0);
or U100 (N_100,In_380,In_16);
nor U101 (N_101,In_113,In_7);
and U102 (N_102,In_316,In_131);
nor U103 (N_103,In_231,In_284);
and U104 (N_104,In_249,In_122);
and U105 (N_105,In_426,In_123);
or U106 (N_106,In_236,In_238);
nor U107 (N_107,In_395,In_269);
nand U108 (N_108,In_300,In_102);
and U109 (N_109,In_78,In_84);
nor U110 (N_110,In_428,In_182);
nand U111 (N_111,In_480,In_160);
and U112 (N_112,In_351,In_285);
nor U113 (N_113,In_425,In_382);
or U114 (N_114,In_225,In_490);
and U115 (N_115,In_118,In_214);
and U116 (N_116,In_158,In_4);
nor U117 (N_117,In_215,In_481);
and U118 (N_118,In_369,In_343);
and U119 (N_119,In_28,In_198);
nor U120 (N_120,In_65,In_244);
nor U121 (N_121,In_201,In_47);
nor U122 (N_122,In_402,In_461);
or U123 (N_123,In_68,In_330);
nand U124 (N_124,In_145,In_166);
nand U125 (N_125,In_479,In_247);
nor U126 (N_126,In_11,In_86);
and U127 (N_127,In_309,In_141);
or U128 (N_128,In_96,In_288);
nor U129 (N_129,In_189,In_361);
nor U130 (N_130,In_72,In_250);
or U131 (N_131,In_192,In_49);
nand U132 (N_132,In_454,In_233);
and U133 (N_133,In_448,In_125);
or U134 (N_134,In_456,In_48);
nand U135 (N_135,In_276,In_317);
and U136 (N_136,In_441,In_246);
or U137 (N_137,In_362,In_471);
and U138 (N_138,In_397,In_100);
nor U139 (N_139,In_259,In_394);
nor U140 (N_140,In_146,In_199);
or U141 (N_141,In_71,In_486);
or U142 (N_142,In_54,In_217);
and U143 (N_143,In_239,In_254);
or U144 (N_144,In_392,In_371);
or U145 (N_145,In_320,In_414);
and U146 (N_146,In_365,In_391);
nand U147 (N_147,In_24,In_218);
and U148 (N_148,In_186,In_478);
or U149 (N_149,In_470,In_327);
or U150 (N_150,In_107,In_359);
nand U151 (N_151,In_372,In_432);
and U152 (N_152,In_304,In_194);
and U153 (N_153,In_334,In_445);
nor U154 (N_154,In_342,In_190);
or U155 (N_155,In_140,In_227);
nor U156 (N_156,In_307,In_228);
nand U157 (N_157,In_1,In_139);
and U158 (N_158,In_137,In_21);
and U159 (N_159,In_156,In_398);
or U160 (N_160,In_59,In_245);
nor U161 (N_161,In_314,In_88);
nor U162 (N_162,In_230,In_268);
or U163 (N_163,In_482,In_169);
and U164 (N_164,In_126,In_40);
and U165 (N_165,In_111,In_163);
nand U166 (N_166,In_419,In_384);
nor U167 (N_167,In_19,In_91);
and U168 (N_168,In_98,In_147);
nor U169 (N_169,In_127,In_252);
or U170 (N_170,In_336,In_193);
nor U171 (N_171,In_3,In_213);
and U172 (N_172,In_136,In_35);
nand U173 (N_173,In_340,In_234);
or U174 (N_174,In_216,In_311);
and U175 (N_175,In_116,In_462);
and U176 (N_176,In_423,In_255);
nor U177 (N_177,In_223,In_424);
or U178 (N_178,In_66,In_257);
or U179 (N_179,In_377,In_173);
or U180 (N_180,In_128,In_104);
and U181 (N_181,In_306,In_130);
nand U182 (N_182,In_94,In_413);
or U183 (N_183,In_99,In_226);
and U184 (N_184,In_18,In_2);
xor U185 (N_185,In_287,In_321);
nand U186 (N_186,In_387,In_119);
nand U187 (N_187,In_407,In_153);
and U188 (N_188,In_168,In_83);
nor U189 (N_189,In_121,In_345);
nand U190 (N_190,In_296,In_295);
nor U191 (N_191,In_437,In_103);
and U192 (N_192,In_10,In_46);
and U193 (N_193,In_498,In_232);
or U194 (N_194,In_242,In_292);
or U195 (N_195,In_101,In_473);
nand U196 (N_196,In_416,In_404);
and U197 (N_197,In_77,In_325);
nor U198 (N_198,In_61,In_278);
or U199 (N_199,In_393,In_433);
nand U200 (N_200,N_40,In_410);
nand U201 (N_201,In_170,N_39);
nor U202 (N_202,N_92,N_193);
nand U203 (N_203,N_131,In_112);
or U204 (N_204,In_474,N_198);
nor U205 (N_205,N_140,N_46);
nand U206 (N_206,N_158,N_114);
or U207 (N_207,N_45,N_199);
or U208 (N_208,N_138,N_159);
nor U209 (N_209,N_119,N_91);
nor U210 (N_210,N_5,In_172);
or U211 (N_211,In_434,N_23);
and U212 (N_212,In_258,In_493);
nand U213 (N_213,N_145,N_73);
nand U214 (N_214,N_0,N_178);
nor U215 (N_215,In_34,N_67);
nor U216 (N_216,In_303,In_248);
and U217 (N_217,N_25,N_148);
nand U218 (N_218,N_143,In_82);
nor U219 (N_219,In_460,In_265);
or U220 (N_220,N_123,N_120);
nand U221 (N_221,N_1,N_181);
nand U222 (N_222,N_54,N_11);
or U223 (N_223,N_163,N_51);
or U224 (N_224,N_174,N_49);
or U225 (N_225,N_17,N_4);
or U226 (N_226,N_35,In_499);
or U227 (N_227,In_229,In_154);
and U228 (N_228,N_42,In_197);
or U229 (N_229,N_157,N_153);
or U230 (N_230,N_14,In_442);
or U231 (N_231,N_3,N_124);
and U232 (N_232,In_109,N_41);
or U233 (N_233,N_105,N_172);
and U234 (N_234,N_112,In_51);
and U235 (N_235,In_349,N_66);
or U236 (N_236,N_60,N_8);
or U237 (N_237,In_323,In_485);
nand U238 (N_238,N_20,In_203);
nand U239 (N_239,N_58,N_129);
nand U240 (N_240,N_70,N_104);
or U241 (N_241,In_204,N_72);
or U242 (N_242,N_166,N_116);
nand U243 (N_243,N_156,N_33);
nor U244 (N_244,N_167,N_50);
or U245 (N_245,In_56,N_52);
and U246 (N_246,In_418,N_7);
or U247 (N_247,N_81,In_62);
nor U248 (N_248,N_192,N_90);
or U249 (N_249,In_224,N_83);
and U250 (N_250,In_241,N_84);
and U251 (N_251,N_82,N_188);
and U252 (N_252,N_27,In_405);
or U253 (N_253,In_97,N_136);
nor U254 (N_254,N_118,N_182);
and U255 (N_255,N_189,In_179);
nor U256 (N_256,N_176,N_150);
or U257 (N_257,N_177,In_495);
nand U258 (N_258,N_133,N_44);
or U259 (N_259,In_328,In_370);
nand U260 (N_260,N_71,N_151);
nand U261 (N_261,In_60,In_313);
nand U262 (N_262,In_290,N_85);
nor U263 (N_263,In_289,N_180);
or U264 (N_264,In_187,In_379);
nand U265 (N_265,N_43,In_447);
and U266 (N_266,N_141,In_178);
xor U267 (N_267,In_206,N_30);
and U268 (N_268,In_9,In_76);
nor U269 (N_269,N_19,N_154);
nor U270 (N_270,In_346,N_137);
nor U271 (N_271,N_125,In_297);
or U272 (N_272,N_47,N_24);
and U273 (N_273,N_121,In_70);
nand U274 (N_274,N_126,N_117);
nand U275 (N_275,In_253,N_144);
and U276 (N_276,N_155,N_169);
nor U277 (N_277,In_341,In_375);
nor U278 (N_278,In_299,N_32);
or U279 (N_279,N_75,N_142);
or U280 (N_280,In_422,In_129);
or U281 (N_281,N_194,In_388);
and U282 (N_282,In_492,N_196);
nor U283 (N_283,N_190,N_161);
and U284 (N_284,N_76,In_310);
and U285 (N_285,N_21,N_165);
nor U286 (N_286,N_63,N_18);
nor U287 (N_287,N_170,N_130);
nand U288 (N_288,N_22,N_139);
nand U289 (N_289,N_61,N_168);
or U290 (N_290,N_183,N_103);
nor U291 (N_291,In_208,N_134);
nor U292 (N_292,In_298,In_12);
nor U293 (N_293,N_110,N_87);
and U294 (N_294,N_37,In_366);
and U295 (N_295,In_308,N_171);
nor U296 (N_296,In_251,In_195);
nand U297 (N_297,N_197,N_162);
or U298 (N_298,N_146,In_270);
nand U299 (N_299,In_5,N_64);
or U300 (N_300,N_38,N_184);
nor U301 (N_301,N_59,N_160);
and U302 (N_302,In_120,N_186);
and U303 (N_303,N_88,N_65);
or U304 (N_304,N_93,N_79);
nor U305 (N_305,In_472,In_95);
and U306 (N_306,N_173,N_100);
nand U307 (N_307,N_97,N_12);
nor U308 (N_308,N_179,In_463);
nand U309 (N_309,N_99,N_107);
or U310 (N_310,In_263,N_113);
nor U311 (N_311,N_109,N_31);
or U312 (N_312,N_147,N_6);
nor U313 (N_313,N_48,In_243);
nand U314 (N_314,N_89,N_195);
and U315 (N_315,N_57,N_94);
and U316 (N_316,In_467,N_2);
or U317 (N_317,N_122,N_191);
nor U318 (N_318,In_483,In_337);
or U319 (N_319,N_77,N_26);
or U320 (N_320,In_174,N_96);
or U321 (N_321,In_44,In_58);
nor U322 (N_322,In_135,In_124);
and U323 (N_323,N_74,In_403);
nor U324 (N_324,In_364,In_318);
nand U325 (N_325,N_36,In_176);
or U326 (N_326,N_28,N_106);
nand U327 (N_327,N_53,N_95);
nor U328 (N_328,N_127,N_164);
nor U329 (N_329,N_101,N_149);
nor U330 (N_330,N_175,N_15);
and U331 (N_331,In_211,N_187);
nand U332 (N_332,N_86,N_152);
or U333 (N_333,N_29,In_155);
and U334 (N_334,In_33,In_13);
and U335 (N_335,In_26,In_484);
nor U336 (N_336,N_68,In_89);
nor U337 (N_337,N_55,N_10);
nand U338 (N_338,N_128,N_132);
and U339 (N_339,N_62,N_13);
nand U340 (N_340,In_32,N_111);
nand U341 (N_341,N_69,N_34);
and U342 (N_342,N_80,N_98);
or U343 (N_343,N_56,N_108);
xnor U344 (N_344,N_185,In_390);
or U345 (N_345,In_87,In_305);
and U346 (N_346,N_135,N_115);
nand U347 (N_347,N_16,In_200);
or U348 (N_348,In_373,N_102);
and U349 (N_349,N_78,N_9);
nor U350 (N_350,N_142,N_5);
or U351 (N_351,In_305,N_79);
or U352 (N_352,N_104,N_87);
nor U353 (N_353,N_26,N_144);
and U354 (N_354,N_2,N_67);
and U355 (N_355,N_165,N_59);
or U356 (N_356,In_373,N_141);
or U357 (N_357,N_20,N_172);
nor U358 (N_358,N_69,N_49);
nor U359 (N_359,In_297,N_136);
or U360 (N_360,N_69,N_146);
nor U361 (N_361,In_328,N_117);
nor U362 (N_362,N_139,In_13);
or U363 (N_363,N_118,N_169);
and U364 (N_364,In_12,N_35);
or U365 (N_365,N_4,N_95);
nor U366 (N_366,N_100,In_248);
or U367 (N_367,In_472,N_130);
nand U368 (N_368,In_70,In_124);
nand U369 (N_369,In_493,N_111);
nor U370 (N_370,N_116,N_25);
or U371 (N_371,N_185,N_15);
nor U372 (N_372,In_474,In_390);
and U373 (N_373,N_196,N_67);
nor U374 (N_374,In_58,N_88);
and U375 (N_375,N_12,N_174);
nand U376 (N_376,N_119,N_107);
nor U377 (N_377,N_111,In_229);
nand U378 (N_378,N_43,In_174);
nand U379 (N_379,In_467,N_113);
or U380 (N_380,In_251,In_290);
nand U381 (N_381,N_108,In_299);
or U382 (N_382,N_105,N_42);
or U383 (N_383,N_194,N_64);
nand U384 (N_384,In_467,N_110);
nand U385 (N_385,N_64,N_70);
nor U386 (N_386,In_187,N_87);
or U387 (N_387,N_101,In_463);
or U388 (N_388,N_175,N_52);
nand U389 (N_389,N_190,N_11);
nor U390 (N_390,N_32,N_153);
or U391 (N_391,N_169,N_167);
nor U392 (N_392,N_56,N_82);
nand U393 (N_393,N_44,N_196);
or U394 (N_394,In_289,N_172);
nand U395 (N_395,N_118,N_188);
nor U396 (N_396,N_174,In_484);
or U397 (N_397,N_149,N_196);
or U398 (N_398,N_49,In_308);
or U399 (N_399,N_154,N_27);
or U400 (N_400,N_254,N_384);
or U401 (N_401,N_389,N_390);
nor U402 (N_402,N_314,N_328);
nand U403 (N_403,N_270,N_355);
nand U404 (N_404,N_294,N_242);
nand U405 (N_405,N_209,N_305);
nand U406 (N_406,N_340,N_298);
or U407 (N_407,N_245,N_378);
nor U408 (N_408,N_286,N_344);
nor U409 (N_409,N_338,N_381);
nor U410 (N_410,N_259,N_238);
or U411 (N_411,N_313,N_386);
or U412 (N_412,N_276,N_218);
and U413 (N_413,N_249,N_337);
or U414 (N_414,N_203,N_205);
nand U415 (N_415,N_388,N_222);
or U416 (N_416,N_393,N_370);
nor U417 (N_417,N_334,N_374);
or U418 (N_418,N_364,N_397);
nor U419 (N_419,N_351,N_301);
nand U420 (N_420,N_219,N_280);
nor U421 (N_421,N_296,N_202);
nor U422 (N_422,N_387,N_320);
nand U423 (N_423,N_317,N_315);
or U424 (N_424,N_367,N_247);
nor U425 (N_425,N_365,N_256);
or U426 (N_426,N_327,N_215);
nor U427 (N_427,N_221,N_233);
or U428 (N_428,N_382,N_360);
nor U429 (N_429,N_288,N_200);
nand U430 (N_430,N_368,N_321);
nand U431 (N_431,N_293,N_361);
or U432 (N_432,N_309,N_323);
nand U433 (N_433,N_394,N_252);
or U434 (N_434,N_376,N_335);
or U435 (N_435,N_204,N_295);
or U436 (N_436,N_380,N_358);
or U437 (N_437,N_263,N_239);
nand U438 (N_438,N_354,N_230);
nor U439 (N_439,N_267,N_348);
nor U440 (N_440,N_325,N_359);
or U441 (N_441,N_342,N_223);
nand U442 (N_442,N_326,N_278);
nor U443 (N_443,N_211,N_345);
nor U444 (N_444,N_307,N_274);
nor U445 (N_445,N_308,N_285);
nand U446 (N_446,N_227,N_290);
nand U447 (N_447,N_329,N_312);
or U448 (N_448,N_206,N_322);
nand U449 (N_449,N_346,N_371);
and U450 (N_450,N_234,N_398);
and U451 (N_451,N_302,N_210);
nand U452 (N_452,N_369,N_392);
or U453 (N_453,N_268,N_356);
nor U454 (N_454,N_332,N_217);
and U455 (N_455,N_347,N_257);
and U456 (N_456,N_214,N_319);
nand U457 (N_457,N_303,N_224);
nor U458 (N_458,N_250,N_324);
nand U459 (N_459,N_248,N_300);
or U460 (N_460,N_212,N_275);
nor U461 (N_461,N_213,N_281);
or U462 (N_462,N_373,N_260);
and U463 (N_463,N_366,N_277);
or U464 (N_464,N_282,N_253);
or U465 (N_465,N_310,N_266);
nand U466 (N_466,N_291,N_241);
nand U467 (N_467,N_383,N_385);
and U468 (N_468,N_297,N_353);
nand U469 (N_469,N_235,N_283);
nand U470 (N_470,N_336,N_220);
nor U471 (N_471,N_255,N_316);
nor U472 (N_472,N_269,N_229);
or U473 (N_473,N_262,N_349);
nor U474 (N_474,N_246,N_372);
and U475 (N_475,N_237,N_375);
or U476 (N_476,N_395,N_306);
or U477 (N_477,N_207,N_399);
nand U478 (N_478,N_339,N_362);
and U479 (N_479,N_216,N_352);
or U480 (N_480,N_264,N_272);
nand U481 (N_481,N_341,N_377);
or U482 (N_482,N_350,N_273);
and U483 (N_483,N_228,N_226);
nand U484 (N_484,N_232,N_258);
nor U485 (N_485,N_331,N_201);
nor U486 (N_486,N_208,N_357);
nand U487 (N_487,N_304,N_271);
and U488 (N_488,N_311,N_279);
nand U489 (N_489,N_333,N_231);
and U490 (N_490,N_236,N_251);
or U491 (N_491,N_379,N_225);
or U492 (N_492,N_396,N_391);
nor U493 (N_493,N_292,N_287);
nand U494 (N_494,N_261,N_330);
nand U495 (N_495,N_343,N_243);
or U496 (N_496,N_318,N_363);
nor U497 (N_497,N_289,N_284);
nor U498 (N_498,N_240,N_299);
nor U499 (N_499,N_244,N_265);
or U500 (N_500,N_299,N_217);
nand U501 (N_501,N_327,N_208);
nor U502 (N_502,N_357,N_390);
nor U503 (N_503,N_389,N_311);
nand U504 (N_504,N_208,N_345);
nor U505 (N_505,N_206,N_348);
nor U506 (N_506,N_380,N_294);
nand U507 (N_507,N_277,N_210);
nand U508 (N_508,N_212,N_247);
nand U509 (N_509,N_386,N_307);
or U510 (N_510,N_329,N_284);
nand U511 (N_511,N_272,N_310);
nand U512 (N_512,N_298,N_235);
and U513 (N_513,N_366,N_244);
nor U514 (N_514,N_258,N_215);
and U515 (N_515,N_259,N_389);
or U516 (N_516,N_324,N_312);
and U517 (N_517,N_342,N_344);
or U518 (N_518,N_399,N_289);
or U519 (N_519,N_266,N_274);
nor U520 (N_520,N_200,N_334);
and U521 (N_521,N_245,N_293);
or U522 (N_522,N_218,N_229);
or U523 (N_523,N_266,N_390);
nand U524 (N_524,N_341,N_272);
nand U525 (N_525,N_281,N_348);
or U526 (N_526,N_356,N_240);
or U527 (N_527,N_362,N_370);
and U528 (N_528,N_314,N_207);
nand U529 (N_529,N_375,N_317);
nand U530 (N_530,N_267,N_205);
and U531 (N_531,N_381,N_269);
nor U532 (N_532,N_266,N_247);
or U533 (N_533,N_236,N_252);
nor U534 (N_534,N_392,N_224);
nand U535 (N_535,N_205,N_309);
nand U536 (N_536,N_306,N_361);
nand U537 (N_537,N_287,N_324);
nand U538 (N_538,N_301,N_242);
or U539 (N_539,N_278,N_292);
nor U540 (N_540,N_339,N_242);
or U541 (N_541,N_208,N_289);
nand U542 (N_542,N_227,N_381);
or U543 (N_543,N_288,N_323);
nor U544 (N_544,N_381,N_261);
or U545 (N_545,N_354,N_341);
or U546 (N_546,N_370,N_258);
nor U547 (N_547,N_311,N_288);
nand U548 (N_548,N_392,N_258);
or U549 (N_549,N_355,N_201);
or U550 (N_550,N_339,N_272);
nor U551 (N_551,N_272,N_380);
nand U552 (N_552,N_200,N_311);
nand U553 (N_553,N_293,N_392);
nor U554 (N_554,N_303,N_307);
nor U555 (N_555,N_329,N_396);
nor U556 (N_556,N_233,N_208);
nand U557 (N_557,N_320,N_311);
nor U558 (N_558,N_202,N_211);
or U559 (N_559,N_338,N_239);
nor U560 (N_560,N_248,N_235);
nand U561 (N_561,N_259,N_282);
or U562 (N_562,N_297,N_340);
or U563 (N_563,N_240,N_351);
or U564 (N_564,N_324,N_220);
and U565 (N_565,N_275,N_224);
and U566 (N_566,N_211,N_299);
and U567 (N_567,N_377,N_244);
nand U568 (N_568,N_231,N_263);
nand U569 (N_569,N_208,N_201);
and U570 (N_570,N_221,N_356);
nand U571 (N_571,N_345,N_223);
or U572 (N_572,N_207,N_321);
nor U573 (N_573,N_380,N_365);
or U574 (N_574,N_311,N_318);
or U575 (N_575,N_239,N_206);
nor U576 (N_576,N_219,N_378);
nand U577 (N_577,N_252,N_339);
and U578 (N_578,N_203,N_378);
or U579 (N_579,N_366,N_389);
nand U580 (N_580,N_267,N_386);
and U581 (N_581,N_247,N_279);
nand U582 (N_582,N_360,N_385);
nor U583 (N_583,N_269,N_324);
and U584 (N_584,N_307,N_378);
nand U585 (N_585,N_302,N_219);
and U586 (N_586,N_395,N_384);
or U587 (N_587,N_201,N_269);
nor U588 (N_588,N_350,N_231);
and U589 (N_589,N_221,N_237);
nor U590 (N_590,N_262,N_313);
and U591 (N_591,N_305,N_394);
nand U592 (N_592,N_313,N_370);
nand U593 (N_593,N_285,N_298);
and U594 (N_594,N_220,N_263);
or U595 (N_595,N_286,N_301);
nor U596 (N_596,N_240,N_256);
and U597 (N_597,N_372,N_204);
nand U598 (N_598,N_286,N_285);
or U599 (N_599,N_333,N_337);
nor U600 (N_600,N_514,N_418);
nor U601 (N_601,N_573,N_521);
or U602 (N_602,N_594,N_516);
nand U603 (N_603,N_477,N_448);
nand U604 (N_604,N_482,N_506);
and U605 (N_605,N_478,N_596);
nand U606 (N_606,N_413,N_454);
and U607 (N_607,N_430,N_440);
or U608 (N_608,N_533,N_589);
nand U609 (N_609,N_502,N_542);
and U610 (N_610,N_563,N_495);
nor U611 (N_611,N_547,N_500);
and U612 (N_612,N_496,N_535);
and U613 (N_613,N_554,N_544);
or U614 (N_614,N_576,N_420);
nand U615 (N_615,N_458,N_403);
or U616 (N_616,N_451,N_488);
or U617 (N_617,N_592,N_443);
and U618 (N_618,N_597,N_577);
nand U619 (N_619,N_434,N_505);
nor U620 (N_620,N_417,N_582);
nor U621 (N_621,N_459,N_517);
or U622 (N_622,N_524,N_433);
nand U623 (N_623,N_476,N_531);
and U624 (N_624,N_485,N_472);
or U625 (N_625,N_461,N_400);
nor U626 (N_626,N_537,N_431);
nor U627 (N_627,N_479,N_526);
or U628 (N_628,N_515,N_401);
nand U629 (N_629,N_405,N_583);
and U630 (N_630,N_491,N_539);
or U631 (N_631,N_538,N_522);
and U632 (N_632,N_412,N_540);
and U633 (N_633,N_572,N_559);
nor U634 (N_634,N_429,N_591);
and U635 (N_635,N_578,N_530);
and U636 (N_636,N_548,N_501);
nand U637 (N_637,N_450,N_410);
or U638 (N_638,N_409,N_407);
nor U639 (N_639,N_446,N_511);
nand U640 (N_640,N_422,N_503);
and U641 (N_641,N_408,N_556);
nand U642 (N_642,N_427,N_453);
or U643 (N_643,N_490,N_421);
nor U644 (N_644,N_571,N_460);
or U645 (N_645,N_444,N_509);
nand U646 (N_646,N_411,N_579);
nor U647 (N_647,N_492,N_402);
or U648 (N_648,N_425,N_465);
nor U649 (N_649,N_534,N_580);
or U650 (N_650,N_428,N_549);
nand U651 (N_651,N_587,N_493);
and U652 (N_652,N_406,N_471);
nand U653 (N_653,N_439,N_512);
or U654 (N_654,N_564,N_463);
and U655 (N_655,N_543,N_470);
or U656 (N_656,N_510,N_436);
nand U657 (N_657,N_593,N_487);
nand U658 (N_658,N_584,N_585);
xor U659 (N_659,N_513,N_550);
or U660 (N_660,N_404,N_536);
nor U661 (N_661,N_546,N_468);
nand U662 (N_662,N_499,N_532);
nor U663 (N_663,N_424,N_586);
nor U664 (N_664,N_525,N_560);
and U665 (N_665,N_447,N_552);
or U666 (N_666,N_442,N_473);
and U667 (N_667,N_445,N_494);
or U668 (N_668,N_416,N_545);
and U669 (N_669,N_504,N_574);
or U670 (N_670,N_441,N_529);
nand U671 (N_671,N_581,N_497);
and U672 (N_672,N_527,N_562);
and U673 (N_673,N_568,N_565);
nand U674 (N_674,N_518,N_575);
and U675 (N_675,N_519,N_423);
nand U676 (N_676,N_561,N_466);
nand U677 (N_677,N_590,N_541);
and U678 (N_678,N_462,N_599);
nor U679 (N_679,N_457,N_426);
or U680 (N_680,N_553,N_456);
and U681 (N_681,N_435,N_438);
nor U682 (N_682,N_588,N_523);
and U683 (N_683,N_566,N_483);
nor U684 (N_684,N_569,N_555);
nand U685 (N_685,N_484,N_415);
nand U686 (N_686,N_480,N_455);
nor U687 (N_687,N_464,N_437);
and U688 (N_688,N_419,N_474);
or U689 (N_689,N_475,N_570);
nor U690 (N_690,N_498,N_452);
nor U691 (N_691,N_489,N_557);
nor U692 (N_692,N_449,N_469);
and U693 (N_693,N_432,N_595);
or U694 (N_694,N_551,N_414);
nand U695 (N_695,N_481,N_486);
or U696 (N_696,N_520,N_598);
nand U697 (N_697,N_507,N_467);
nor U698 (N_698,N_567,N_528);
or U699 (N_699,N_558,N_508);
and U700 (N_700,N_445,N_429);
nor U701 (N_701,N_414,N_400);
or U702 (N_702,N_501,N_418);
and U703 (N_703,N_555,N_523);
or U704 (N_704,N_548,N_580);
nand U705 (N_705,N_556,N_429);
or U706 (N_706,N_470,N_508);
and U707 (N_707,N_482,N_595);
or U708 (N_708,N_427,N_531);
nand U709 (N_709,N_582,N_595);
and U710 (N_710,N_532,N_591);
or U711 (N_711,N_496,N_534);
nor U712 (N_712,N_580,N_490);
or U713 (N_713,N_556,N_576);
or U714 (N_714,N_567,N_410);
nand U715 (N_715,N_448,N_492);
or U716 (N_716,N_499,N_449);
and U717 (N_717,N_478,N_501);
and U718 (N_718,N_454,N_452);
and U719 (N_719,N_520,N_480);
and U720 (N_720,N_487,N_584);
or U721 (N_721,N_594,N_532);
nor U722 (N_722,N_524,N_555);
nand U723 (N_723,N_513,N_574);
or U724 (N_724,N_559,N_583);
nand U725 (N_725,N_515,N_419);
nor U726 (N_726,N_577,N_459);
and U727 (N_727,N_435,N_573);
or U728 (N_728,N_454,N_594);
and U729 (N_729,N_428,N_490);
nor U730 (N_730,N_463,N_464);
or U731 (N_731,N_578,N_473);
and U732 (N_732,N_408,N_552);
and U733 (N_733,N_492,N_521);
nand U734 (N_734,N_404,N_544);
nand U735 (N_735,N_521,N_577);
nor U736 (N_736,N_406,N_419);
nor U737 (N_737,N_410,N_537);
nand U738 (N_738,N_451,N_401);
or U739 (N_739,N_551,N_544);
nand U740 (N_740,N_490,N_427);
xnor U741 (N_741,N_528,N_544);
and U742 (N_742,N_415,N_567);
and U743 (N_743,N_482,N_496);
nor U744 (N_744,N_549,N_539);
nor U745 (N_745,N_524,N_558);
nand U746 (N_746,N_468,N_588);
nand U747 (N_747,N_484,N_561);
and U748 (N_748,N_417,N_569);
and U749 (N_749,N_538,N_463);
and U750 (N_750,N_555,N_577);
nor U751 (N_751,N_424,N_445);
or U752 (N_752,N_574,N_534);
nor U753 (N_753,N_570,N_548);
and U754 (N_754,N_511,N_453);
or U755 (N_755,N_400,N_407);
nor U756 (N_756,N_476,N_518);
or U757 (N_757,N_512,N_586);
nand U758 (N_758,N_417,N_479);
nor U759 (N_759,N_407,N_567);
nor U760 (N_760,N_517,N_508);
nor U761 (N_761,N_529,N_593);
nand U762 (N_762,N_445,N_548);
and U763 (N_763,N_586,N_578);
nor U764 (N_764,N_597,N_573);
nor U765 (N_765,N_549,N_446);
or U766 (N_766,N_540,N_523);
nand U767 (N_767,N_461,N_440);
nor U768 (N_768,N_484,N_459);
and U769 (N_769,N_425,N_477);
nand U770 (N_770,N_437,N_587);
and U771 (N_771,N_409,N_468);
and U772 (N_772,N_462,N_452);
and U773 (N_773,N_403,N_505);
nor U774 (N_774,N_513,N_524);
or U775 (N_775,N_567,N_599);
nand U776 (N_776,N_434,N_410);
xor U777 (N_777,N_483,N_598);
nor U778 (N_778,N_507,N_570);
nand U779 (N_779,N_548,N_578);
or U780 (N_780,N_529,N_517);
nor U781 (N_781,N_572,N_580);
and U782 (N_782,N_498,N_525);
or U783 (N_783,N_510,N_428);
or U784 (N_784,N_528,N_503);
nor U785 (N_785,N_503,N_425);
nand U786 (N_786,N_419,N_535);
nand U787 (N_787,N_499,N_488);
nand U788 (N_788,N_527,N_472);
nand U789 (N_789,N_537,N_571);
and U790 (N_790,N_507,N_495);
and U791 (N_791,N_472,N_495);
nand U792 (N_792,N_531,N_431);
or U793 (N_793,N_497,N_447);
and U794 (N_794,N_560,N_483);
nand U795 (N_795,N_503,N_579);
nor U796 (N_796,N_470,N_567);
nor U797 (N_797,N_523,N_453);
and U798 (N_798,N_476,N_550);
and U799 (N_799,N_539,N_560);
nor U800 (N_800,N_708,N_692);
or U801 (N_801,N_758,N_681);
or U802 (N_802,N_770,N_765);
or U803 (N_803,N_714,N_752);
nor U804 (N_804,N_639,N_719);
and U805 (N_805,N_631,N_780);
nand U806 (N_806,N_742,N_670);
and U807 (N_807,N_712,N_612);
or U808 (N_808,N_761,N_690);
nand U809 (N_809,N_617,N_777);
nand U810 (N_810,N_771,N_687);
and U811 (N_811,N_721,N_730);
or U812 (N_812,N_695,N_682);
nand U813 (N_813,N_688,N_666);
nor U814 (N_814,N_672,N_627);
nor U815 (N_815,N_665,N_636);
or U816 (N_816,N_610,N_654);
or U817 (N_817,N_602,N_652);
nor U818 (N_818,N_679,N_727);
and U819 (N_819,N_608,N_671);
or U820 (N_820,N_711,N_607);
nand U821 (N_821,N_728,N_662);
nor U822 (N_822,N_774,N_701);
nand U823 (N_823,N_675,N_732);
and U824 (N_824,N_704,N_798);
and U825 (N_825,N_667,N_792);
and U826 (N_826,N_615,N_789);
and U827 (N_827,N_788,N_753);
or U828 (N_828,N_733,N_673);
nand U829 (N_829,N_710,N_632);
nor U830 (N_830,N_678,N_751);
and U831 (N_831,N_637,N_737);
and U832 (N_832,N_717,N_677);
nor U833 (N_833,N_643,N_787);
nand U834 (N_834,N_713,N_745);
or U835 (N_835,N_658,N_656);
or U836 (N_836,N_760,N_781);
and U837 (N_837,N_778,N_629);
nand U838 (N_838,N_791,N_657);
and U839 (N_839,N_739,N_649);
nor U840 (N_840,N_763,N_647);
nand U841 (N_841,N_619,N_779);
or U842 (N_842,N_715,N_621);
nand U843 (N_843,N_640,N_769);
nand U844 (N_844,N_766,N_685);
xor U845 (N_845,N_716,N_724);
nand U846 (N_846,N_624,N_738);
nor U847 (N_847,N_703,N_691);
nor U848 (N_848,N_686,N_706);
or U849 (N_849,N_726,N_622);
or U850 (N_850,N_795,N_749);
nand U851 (N_851,N_669,N_694);
or U852 (N_852,N_729,N_600);
nand U853 (N_853,N_720,N_611);
nand U854 (N_854,N_783,N_744);
and U855 (N_855,N_635,N_759);
nand U856 (N_856,N_773,N_683);
or U857 (N_857,N_768,N_660);
or U858 (N_858,N_723,N_653);
nor U859 (N_859,N_775,N_734);
nand U860 (N_860,N_799,N_609);
nor U861 (N_861,N_796,N_772);
or U862 (N_862,N_693,N_603);
nand U863 (N_863,N_782,N_741);
nor U864 (N_864,N_757,N_630);
nand U865 (N_865,N_623,N_606);
and U866 (N_866,N_756,N_628);
nand U867 (N_867,N_731,N_605);
nand U868 (N_868,N_700,N_645);
or U869 (N_869,N_743,N_702);
nor U870 (N_870,N_750,N_784);
nor U871 (N_871,N_776,N_655);
or U872 (N_872,N_663,N_755);
or U873 (N_873,N_718,N_705);
or U874 (N_874,N_668,N_725);
nor U875 (N_875,N_659,N_793);
nor U876 (N_876,N_620,N_797);
nor U877 (N_877,N_764,N_664);
or U878 (N_878,N_633,N_709);
nand U879 (N_879,N_785,N_650);
nand U880 (N_880,N_680,N_746);
and U881 (N_881,N_648,N_641);
and U882 (N_882,N_634,N_754);
nor U883 (N_883,N_748,N_786);
nor U884 (N_884,N_626,N_676);
and U885 (N_885,N_722,N_689);
nand U886 (N_886,N_747,N_740);
nor U887 (N_887,N_651,N_697);
nor U888 (N_888,N_646,N_638);
nand U889 (N_889,N_767,N_614);
and U890 (N_890,N_696,N_642);
nor U891 (N_891,N_735,N_699);
nor U892 (N_892,N_794,N_674);
or U893 (N_893,N_684,N_613);
nor U894 (N_894,N_736,N_762);
and U895 (N_895,N_616,N_707);
and U896 (N_896,N_644,N_661);
nand U897 (N_897,N_625,N_790);
or U898 (N_898,N_698,N_604);
or U899 (N_899,N_601,N_618);
or U900 (N_900,N_755,N_779);
nor U901 (N_901,N_679,N_745);
nand U902 (N_902,N_705,N_640);
nor U903 (N_903,N_794,N_703);
nand U904 (N_904,N_754,N_612);
nand U905 (N_905,N_624,N_779);
or U906 (N_906,N_747,N_656);
or U907 (N_907,N_747,N_634);
or U908 (N_908,N_729,N_791);
nor U909 (N_909,N_741,N_730);
nor U910 (N_910,N_779,N_794);
and U911 (N_911,N_782,N_663);
and U912 (N_912,N_653,N_676);
nor U913 (N_913,N_683,N_650);
nor U914 (N_914,N_682,N_617);
or U915 (N_915,N_798,N_613);
or U916 (N_916,N_689,N_790);
or U917 (N_917,N_792,N_765);
and U918 (N_918,N_761,N_609);
or U919 (N_919,N_703,N_686);
or U920 (N_920,N_607,N_762);
and U921 (N_921,N_626,N_603);
or U922 (N_922,N_605,N_617);
nor U923 (N_923,N_786,N_792);
and U924 (N_924,N_789,N_614);
nor U925 (N_925,N_697,N_645);
or U926 (N_926,N_799,N_727);
nand U927 (N_927,N_729,N_639);
or U928 (N_928,N_794,N_610);
nor U929 (N_929,N_698,N_794);
or U930 (N_930,N_694,N_642);
and U931 (N_931,N_646,N_751);
and U932 (N_932,N_682,N_619);
and U933 (N_933,N_612,N_725);
and U934 (N_934,N_719,N_724);
or U935 (N_935,N_648,N_693);
nor U936 (N_936,N_776,N_618);
or U937 (N_937,N_778,N_645);
or U938 (N_938,N_739,N_717);
and U939 (N_939,N_718,N_609);
or U940 (N_940,N_692,N_747);
or U941 (N_941,N_735,N_635);
nor U942 (N_942,N_755,N_720);
nand U943 (N_943,N_715,N_672);
or U944 (N_944,N_724,N_791);
nand U945 (N_945,N_643,N_663);
nor U946 (N_946,N_660,N_691);
or U947 (N_947,N_766,N_679);
or U948 (N_948,N_710,N_732);
nand U949 (N_949,N_796,N_757);
or U950 (N_950,N_653,N_603);
and U951 (N_951,N_622,N_603);
nand U952 (N_952,N_660,N_739);
nand U953 (N_953,N_660,N_765);
and U954 (N_954,N_687,N_720);
nand U955 (N_955,N_716,N_742);
nand U956 (N_956,N_606,N_788);
and U957 (N_957,N_750,N_730);
nor U958 (N_958,N_741,N_636);
nand U959 (N_959,N_687,N_767);
and U960 (N_960,N_657,N_716);
and U961 (N_961,N_728,N_613);
nand U962 (N_962,N_707,N_622);
or U963 (N_963,N_665,N_752);
or U964 (N_964,N_660,N_748);
nor U965 (N_965,N_706,N_761);
nor U966 (N_966,N_744,N_750);
or U967 (N_967,N_610,N_668);
nor U968 (N_968,N_769,N_751);
and U969 (N_969,N_793,N_759);
nand U970 (N_970,N_626,N_675);
or U971 (N_971,N_621,N_657);
nand U972 (N_972,N_687,N_662);
nor U973 (N_973,N_748,N_691);
nand U974 (N_974,N_799,N_682);
xnor U975 (N_975,N_625,N_668);
nor U976 (N_976,N_738,N_751);
nand U977 (N_977,N_659,N_704);
or U978 (N_978,N_649,N_726);
nand U979 (N_979,N_607,N_648);
or U980 (N_980,N_678,N_622);
and U981 (N_981,N_794,N_626);
nand U982 (N_982,N_606,N_782);
and U983 (N_983,N_662,N_604);
or U984 (N_984,N_614,N_711);
or U985 (N_985,N_614,N_686);
and U986 (N_986,N_608,N_765);
or U987 (N_987,N_798,N_706);
nor U988 (N_988,N_735,N_610);
or U989 (N_989,N_737,N_670);
or U990 (N_990,N_749,N_663);
nor U991 (N_991,N_709,N_782);
or U992 (N_992,N_720,N_773);
nand U993 (N_993,N_733,N_601);
or U994 (N_994,N_602,N_732);
and U995 (N_995,N_783,N_718);
or U996 (N_996,N_783,N_731);
nor U997 (N_997,N_631,N_794);
or U998 (N_998,N_706,N_677);
or U999 (N_999,N_673,N_772);
nand U1000 (N_1000,N_998,N_889);
nand U1001 (N_1001,N_977,N_870);
nor U1002 (N_1002,N_837,N_836);
or U1003 (N_1003,N_873,N_875);
or U1004 (N_1004,N_860,N_980);
and U1005 (N_1005,N_902,N_880);
or U1006 (N_1006,N_964,N_927);
or U1007 (N_1007,N_845,N_821);
and U1008 (N_1008,N_916,N_812);
or U1009 (N_1009,N_993,N_918);
nand U1010 (N_1010,N_835,N_908);
nand U1011 (N_1011,N_804,N_800);
nor U1012 (N_1012,N_921,N_997);
nand U1013 (N_1013,N_868,N_862);
xor U1014 (N_1014,N_859,N_952);
nor U1015 (N_1015,N_935,N_941);
nand U1016 (N_1016,N_817,N_929);
or U1017 (N_1017,N_815,N_891);
nor U1018 (N_1018,N_966,N_915);
nor U1019 (N_1019,N_940,N_852);
or U1020 (N_1020,N_976,N_841);
and U1021 (N_1021,N_933,N_828);
or U1022 (N_1022,N_819,N_970);
and U1023 (N_1023,N_951,N_959);
and U1024 (N_1024,N_999,N_842);
or U1025 (N_1025,N_864,N_810);
nor U1026 (N_1026,N_856,N_809);
nand U1027 (N_1027,N_851,N_896);
nand U1028 (N_1028,N_876,N_914);
nor U1029 (N_1029,N_863,N_991);
nor U1030 (N_1030,N_811,N_960);
and U1031 (N_1031,N_801,N_982);
nor U1032 (N_1032,N_942,N_995);
nor U1033 (N_1033,N_932,N_832);
nor U1034 (N_1034,N_963,N_978);
or U1035 (N_1035,N_979,N_866);
or U1036 (N_1036,N_986,N_827);
nand U1037 (N_1037,N_949,N_988);
nor U1038 (N_1038,N_840,N_838);
nand U1039 (N_1039,N_816,N_881);
nor U1040 (N_1040,N_983,N_895);
nor U1041 (N_1041,N_846,N_922);
and U1042 (N_1042,N_967,N_853);
and U1043 (N_1043,N_944,N_822);
or U1044 (N_1044,N_912,N_877);
and U1045 (N_1045,N_945,N_826);
nand U1046 (N_1046,N_901,N_861);
xnor U1047 (N_1047,N_934,N_913);
or U1048 (N_1048,N_962,N_939);
or U1049 (N_1049,N_961,N_965);
or U1050 (N_1050,N_931,N_928);
or U1051 (N_1051,N_865,N_987);
nor U1052 (N_1052,N_981,N_971);
and U1053 (N_1053,N_930,N_955);
and U1054 (N_1054,N_806,N_894);
nand U1055 (N_1055,N_917,N_974);
nor U1056 (N_1056,N_886,N_885);
and U1057 (N_1057,N_813,N_968);
and U1058 (N_1058,N_957,N_936);
nand U1059 (N_1059,N_887,N_858);
or U1060 (N_1060,N_989,N_892);
and U1061 (N_1061,N_871,N_973);
and U1062 (N_1062,N_818,N_893);
or U1063 (N_1063,N_805,N_969);
nor U1064 (N_1064,N_847,N_996);
and U1065 (N_1065,N_899,N_882);
nor U1066 (N_1066,N_920,N_807);
or U1067 (N_1067,N_950,N_898);
or U1068 (N_1068,N_975,N_872);
nand U1069 (N_1069,N_829,N_867);
and U1070 (N_1070,N_903,N_948);
and U1071 (N_1071,N_909,N_958);
or U1072 (N_1072,N_937,N_904);
and U1073 (N_1073,N_833,N_831);
or U1074 (N_1074,N_947,N_924);
or U1075 (N_1075,N_839,N_869);
and U1076 (N_1076,N_900,N_992);
and U1077 (N_1077,N_884,N_857);
or U1078 (N_1078,N_954,N_985);
and U1079 (N_1079,N_814,N_919);
nor U1080 (N_1080,N_926,N_820);
or U1081 (N_1081,N_938,N_907);
or U1082 (N_1082,N_994,N_956);
nand U1083 (N_1083,N_925,N_803);
and U1084 (N_1084,N_825,N_874);
nor U1085 (N_1085,N_802,N_972);
nand U1086 (N_1086,N_946,N_879);
and U1087 (N_1087,N_854,N_883);
or U1088 (N_1088,N_850,N_844);
and U1089 (N_1089,N_984,N_849);
and U1090 (N_1090,N_824,N_855);
nor U1091 (N_1091,N_911,N_943);
and U1092 (N_1092,N_905,N_808);
nor U1093 (N_1093,N_848,N_990);
or U1094 (N_1094,N_897,N_878);
or U1095 (N_1095,N_888,N_823);
nand U1096 (N_1096,N_890,N_843);
or U1097 (N_1097,N_910,N_953);
nand U1098 (N_1098,N_923,N_834);
and U1099 (N_1099,N_830,N_906);
or U1100 (N_1100,N_870,N_906);
and U1101 (N_1101,N_853,N_840);
nand U1102 (N_1102,N_996,N_925);
and U1103 (N_1103,N_893,N_937);
nor U1104 (N_1104,N_821,N_870);
and U1105 (N_1105,N_924,N_830);
nor U1106 (N_1106,N_924,N_867);
and U1107 (N_1107,N_821,N_948);
nor U1108 (N_1108,N_985,N_818);
or U1109 (N_1109,N_884,N_908);
nand U1110 (N_1110,N_993,N_942);
nor U1111 (N_1111,N_830,N_948);
and U1112 (N_1112,N_989,N_826);
or U1113 (N_1113,N_823,N_918);
nand U1114 (N_1114,N_919,N_984);
and U1115 (N_1115,N_871,N_936);
and U1116 (N_1116,N_813,N_863);
nand U1117 (N_1117,N_847,N_831);
and U1118 (N_1118,N_879,N_872);
and U1119 (N_1119,N_992,N_924);
nand U1120 (N_1120,N_927,N_876);
nor U1121 (N_1121,N_888,N_999);
nor U1122 (N_1122,N_994,N_890);
nor U1123 (N_1123,N_812,N_966);
and U1124 (N_1124,N_834,N_805);
nand U1125 (N_1125,N_883,N_861);
nand U1126 (N_1126,N_821,N_988);
and U1127 (N_1127,N_911,N_872);
nor U1128 (N_1128,N_933,N_953);
or U1129 (N_1129,N_909,N_820);
nand U1130 (N_1130,N_955,N_849);
and U1131 (N_1131,N_925,N_958);
nor U1132 (N_1132,N_819,N_985);
and U1133 (N_1133,N_905,N_826);
or U1134 (N_1134,N_835,N_837);
nor U1135 (N_1135,N_858,N_853);
nor U1136 (N_1136,N_933,N_954);
or U1137 (N_1137,N_942,N_892);
nor U1138 (N_1138,N_993,N_904);
nor U1139 (N_1139,N_940,N_914);
or U1140 (N_1140,N_891,N_961);
nand U1141 (N_1141,N_846,N_952);
or U1142 (N_1142,N_988,N_982);
nand U1143 (N_1143,N_876,N_835);
nand U1144 (N_1144,N_943,N_953);
or U1145 (N_1145,N_805,N_998);
xor U1146 (N_1146,N_825,N_952);
or U1147 (N_1147,N_954,N_992);
nor U1148 (N_1148,N_998,N_829);
nand U1149 (N_1149,N_843,N_934);
or U1150 (N_1150,N_942,N_831);
and U1151 (N_1151,N_805,N_926);
nand U1152 (N_1152,N_874,N_885);
and U1153 (N_1153,N_830,N_956);
nor U1154 (N_1154,N_975,N_868);
and U1155 (N_1155,N_927,N_836);
and U1156 (N_1156,N_970,N_987);
or U1157 (N_1157,N_859,N_821);
and U1158 (N_1158,N_828,N_983);
nor U1159 (N_1159,N_898,N_863);
and U1160 (N_1160,N_862,N_843);
and U1161 (N_1161,N_854,N_843);
and U1162 (N_1162,N_900,N_957);
nor U1163 (N_1163,N_868,N_911);
nand U1164 (N_1164,N_993,N_810);
nor U1165 (N_1165,N_816,N_872);
nand U1166 (N_1166,N_801,N_827);
or U1167 (N_1167,N_896,N_979);
nand U1168 (N_1168,N_943,N_891);
nor U1169 (N_1169,N_959,N_936);
nor U1170 (N_1170,N_922,N_971);
nand U1171 (N_1171,N_972,N_872);
and U1172 (N_1172,N_992,N_804);
and U1173 (N_1173,N_959,N_848);
and U1174 (N_1174,N_890,N_897);
nor U1175 (N_1175,N_826,N_814);
and U1176 (N_1176,N_956,N_885);
nand U1177 (N_1177,N_951,N_839);
and U1178 (N_1178,N_867,N_958);
and U1179 (N_1179,N_853,N_857);
or U1180 (N_1180,N_915,N_939);
nor U1181 (N_1181,N_868,N_950);
and U1182 (N_1182,N_889,N_849);
or U1183 (N_1183,N_982,N_870);
and U1184 (N_1184,N_862,N_985);
nor U1185 (N_1185,N_936,N_856);
or U1186 (N_1186,N_935,N_888);
or U1187 (N_1187,N_984,N_827);
and U1188 (N_1188,N_997,N_910);
nand U1189 (N_1189,N_843,N_976);
and U1190 (N_1190,N_952,N_831);
nor U1191 (N_1191,N_942,N_820);
or U1192 (N_1192,N_896,N_925);
or U1193 (N_1193,N_881,N_983);
nand U1194 (N_1194,N_958,N_852);
or U1195 (N_1195,N_970,N_851);
or U1196 (N_1196,N_876,N_923);
or U1197 (N_1197,N_911,N_818);
and U1198 (N_1198,N_903,N_961);
and U1199 (N_1199,N_866,N_822);
or U1200 (N_1200,N_1047,N_1014);
nor U1201 (N_1201,N_1112,N_1097);
nor U1202 (N_1202,N_1022,N_1025);
nand U1203 (N_1203,N_1144,N_1042);
nor U1204 (N_1204,N_1069,N_1123);
or U1205 (N_1205,N_1080,N_1137);
nor U1206 (N_1206,N_1039,N_1045);
or U1207 (N_1207,N_1121,N_1119);
nand U1208 (N_1208,N_1020,N_1138);
nor U1209 (N_1209,N_1191,N_1125);
or U1210 (N_1210,N_1050,N_1098);
nor U1211 (N_1211,N_1064,N_1141);
nor U1212 (N_1212,N_1183,N_1120);
nor U1213 (N_1213,N_1133,N_1167);
and U1214 (N_1214,N_1149,N_1044);
nand U1215 (N_1215,N_1082,N_1172);
nand U1216 (N_1216,N_1102,N_1100);
nand U1217 (N_1217,N_1109,N_1142);
nor U1218 (N_1218,N_1040,N_1037);
nand U1219 (N_1219,N_1083,N_1115);
or U1220 (N_1220,N_1128,N_1159);
nor U1221 (N_1221,N_1156,N_1004);
nand U1222 (N_1222,N_1184,N_1085);
or U1223 (N_1223,N_1150,N_1088);
and U1224 (N_1224,N_1027,N_1181);
nor U1225 (N_1225,N_1010,N_1171);
nor U1226 (N_1226,N_1067,N_1170);
or U1227 (N_1227,N_1023,N_1074);
or U1228 (N_1228,N_1180,N_1066);
or U1229 (N_1229,N_1145,N_1158);
nand U1230 (N_1230,N_1173,N_1190);
nand U1231 (N_1231,N_1081,N_1110);
and U1232 (N_1232,N_1084,N_1054);
or U1233 (N_1233,N_1032,N_1174);
and U1234 (N_1234,N_1058,N_1197);
nand U1235 (N_1235,N_1101,N_1105);
nor U1236 (N_1236,N_1162,N_1015);
nand U1237 (N_1237,N_1016,N_1087);
nor U1238 (N_1238,N_1068,N_1099);
nor U1239 (N_1239,N_1148,N_1187);
nor U1240 (N_1240,N_1001,N_1053);
nand U1241 (N_1241,N_1072,N_1029);
or U1242 (N_1242,N_1033,N_1008);
nand U1243 (N_1243,N_1143,N_1002);
or U1244 (N_1244,N_1062,N_1117);
and U1245 (N_1245,N_1094,N_1086);
and U1246 (N_1246,N_1196,N_1089);
nand U1247 (N_1247,N_1005,N_1107);
nor U1248 (N_1248,N_1051,N_1134);
or U1249 (N_1249,N_1006,N_1135);
and U1250 (N_1250,N_1147,N_1030);
nor U1251 (N_1251,N_1118,N_1021);
nand U1252 (N_1252,N_1160,N_1146);
nor U1253 (N_1253,N_1056,N_1127);
nand U1254 (N_1254,N_1113,N_1161);
or U1255 (N_1255,N_1052,N_1041);
or U1256 (N_1256,N_1034,N_1177);
nor U1257 (N_1257,N_1152,N_1075);
nand U1258 (N_1258,N_1108,N_1186);
and U1259 (N_1259,N_1059,N_1019);
or U1260 (N_1260,N_1078,N_1169);
and U1261 (N_1261,N_1060,N_1017);
nor U1262 (N_1262,N_1035,N_1028);
or U1263 (N_1263,N_1061,N_1093);
and U1264 (N_1264,N_1114,N_1049);
nor U1265 (N_1265,N_1139,N_1168);
or U1266 (N_1266,N_1018,N_1165);
nor U1267 (N_1267,N_1195,N_1124);
nand U1268 (N_1268,N_1154,N_1091);
nand U1269 (N_1269,N_1063,N_1038);
nand U1270 (N_1270,N_1153,N_1007);
and U1271 (N_1271,N_1009,N_1155);
nand U1272 (N_1272,N_1036,N_1000);
and U1273 (N_1273,N_1048,N_1013);
and U1274 (N_1274,N_1031,N_1026);
or U1275 (N_1275,N_1199,N_1126);
or U1276 (N_1276,N_1136,N_1095);
and U1277 (N_1277,N_1179,N_1178);
nor U1278 (N_1278,N_1192,N_1193);
and U1279 (N_1279,N_1157,N_1073);
nand U1280 (N_1280,N_1185,N_1003);
nand U1281 (N_1281,N_1055,N_1092);
nor U1282 (N_1282,N_1012,N_1129);
and U1283 (N_1283,N_1198,N_1106);
nand U1284 (N_1284,N_1194,N_1046);
and U1285 (N_1285,N_1076,N_1103);
nand U1286 (N_1286,N_1057,N_1096);
nand U1287 (N_1287,N_1043,N_1071);
nor U1288 (N_1288,N_1065,N_1140);
nor U1289 (N_1289,N_1077,N_1070);
xnor U1290 (N_1290,N_1090,N_1163);
nor U1291 (N_1291,N_1111,N_1188);
nand U1292 (N_1292,N_1182,N_1104);
nor U1293 (N_1293,N_1189,N_1011);
nand U1294 (N_1294,N_1164,N_1175);
nand U1295 (N_1295,N_1131,N_1116);
nand U1296 (N_1296,N_1151,N_1024);
nand U1297 (N_1297,N_1130,N_1132);
nand U1298 (N_1298,N_1079,N_1176);
or U1299 (N_1299,N_1122,N_1166);
or U1300 (N_1300,N_1016,N_1119);
or U1301 (N_1301,N_1071,N_1008);
and U1302 (N_1302,N_1129,N_1104);
or U1303 (N_1303,N_1167,N_1061);
nand U1304 (N_1304,N_1145,N_1186);
nand U1305 (N_1305,N_1170,N_1099);
nand U1306 (N_1306,N_1039,N_1100);
nand U1307 (N_1307,N_1010,N_1054);
and U1308 (N_1308,N_1199,N_1179);
nor U1309 (N_1309,N_1162,N_1187);
nor U1310 (N_1310,N_1131,N_1117);
nor U1311 (N_1311,N_1021,N_1070);
or U1312 (N_1312,N_1097,N_1002);
nand U1313 (N_1313,N_1093,N_1122);
and U1314 (N_1314,N_1082,N_1176);
and U1315 (N_1315,N_1167,N_1126);
and U1316 (N_1316,N_1016,N_1145);
and U1317 (N_1317,N_1164,N_1099);
or U1318 (N_1318,N_1120,N_1195);
nand U1319 (N_1319,N_1013,N_1028);
nor U1320 (N_1320,N_1118,N_1065);
or U1321 (N_1321,N_1135,N_1167);
nand U1322 (N_1322,N_1119,N_1057);
or U1323 (N_1323,N_1006,N_1008);
nor U1324 (N_1324,N_1146,N_1159);
or U1325 (N_1325,N_1078,N_1175);
nor U1326 (N_1326,N_1180,N_1027);
nor U1327 (N_1327,N_1103,N_1087);
nand U1328 (N_1328,N_1029,N_1117);
nand U1329 (N_1329,N_1014,N_1171);
or U1330 (N_1330,N_1100,N_1029);
and U1331 (N_1331,N_1108,N_1103);
or U1332 (N_1332,N_1043,N_1127);
nor U1333 (N_1333,N_1145,N_1121);
or U1334 (N_1334,N_1104,N_1069);
or U1335 (N_1335,N_1026,N_1184);
and U1336 (N_1336,N_1128,N_1157);
or U1337 (N_1337,N_1194,N_1158);
nand U1338 (N_1338,N_1086,N_1027);
nor U1339 (N_1339,N_1178,N_1058);
and U1340 (N_1340,N_1110,N_1010);
and U1341 (N_1341,N_1105,N_1178);
nand U1342 (N_1342,N_1054,N_1123);
nand U1343 (N_1343,N_1038,N_1179);
nor U1344 (N_1344,N_1015,N_1164);
nand U1345 (N_1345,N_1085,N_1191);
nor U1346 (N_1346,N_1059,N_1101);
and U1347 (N_1347,N_1092,N_1171);
or U1348 (N_1348,N_1077,N_1112);
nor U1349 (N_1349,N_1123,N_1003);
nor U1350 (N_1350,N_1155,N_1039);
nand U1351 (N_1351,N_1154,N_1180);
nor U1352 (N_1352,N_1071,N_1096);
or U1353 (N_1353,N_1151,N_1022);
nand U1354 (N_1354,N_1064,N_1070);
and U1355 (N_1355,N_1065,N_1188);
nor U1356 (N_1356,N_1061,N_1134);
or U1357 (N_1357,N_1046,N_1148);
or U1358 (N_1358,N_1020,N_1011);
and U1359 (N_1359,N_1177,N_1067);
nand U1360 (N_1360,N_1136,N_1155);
nor U1361 (N_1361,N_1044,N_1156);
and U1362 (N_1362,N_1121,N_1193);
or U1363 (N_1363,N_1095,N_1138);
or U1364 (N_1364,N_1098,N_1165);
and U1365 (N_1365,N_1078,N_1185);
nand U1366 (N_1366,N_1081,N_1091);
or U1367 (N_1367,N_1161,N_1020);
or U1368 (N_1368,N_1095,N_1052);
or U1369 (N_1369,N_1068,N_1111);
nor U1370 (N_1370,N_1061,N_1136);
nand U1371 (N_1371,N_1070,N_1162);
nand U1372 (N_1372,N_1130,N_1103);
and U1373 (N_1373,N_1119,N_1135);
or U1374 (N_1374,N_1061,N_1039);
or U1375 (N_1375,N_1130,N_1020);
and U1376 (N_1376,N_1074,N_1016);
nor U1377 (N_1377,N_1002,N_1131);
and U1378 (N_1378,N_1154,N_1105);
and U1379 (N_1379,N_1137,N_1143);
nor U1380 (N_1380,N_1033,N_1165);
nand U1381 (N_1381,N_1150,N_1112);
nand U1382 (N_1382,N_1191,N_1119);
nor U1383 (N_1383,N_1061,N_1169);
nand U1384 (N_1384,N_1069,N_1087);
nand U1385 (N_1385,N_1199,N_1032);
and U1386 (N_1386,N_1184,N_1155);
nor U1387 (N_1387,N_1045,N_1099);
and U1388 (N_1388,N_1065,N_1167);
or U1389 (N_1389,N_1107,N_1136);
and U1390 (N_1390,N_1145,N_1196);
or U1391 (N_1391,N_1105,N_1024);
nand U1392 (N_1392,N_1133,N_1126);
and U1393 (N_1393,N_1046,N_1159);
nand U1394 (N_1394,N_1181,N_1138);
and U1395 (N_1395,N_1037,N_1053);
nor U1396 (N_1396,N_1176,N_1097);
nand U1397 (N_1397,N_1153,N_1061);
nand U1398 (N_1398,N_1033,N_1032);
nand U1399 (N_1399,N_1050,N_1190);
and U1400 (N_1400,N_1326,N_1274);
or U1401 (N_1401,N_1213,N_1269);
or U1402 (N_1402,N_1238,N_1207);
nor U1403 (N_1403,N_1302,N_1303);
or U1404 (N_1404,N_1385,N_1257);
and U1405 (N_1405,N_1321,N_1256);
nand U1406 (N_1406,N_1245,N_1393);
nor U1407 (N_1407,N_1305,N_1211);
and U1408 (N_1408,N_1248,N_1365);
and U1409 (N_1409,N_1296,N_1231);
and U1410 (N_1410,N_1251,N_1223);
nand U1411 (N_1411,N_1299,N_1233);
nor U1412 (N_1412,N_1328,N_1335);
and U1413 (N_1413,N_1225,N_1373);
and U1414 (N_1414,N_1208,N_1398);
and U1415 (N_1415,N_1347,N_1341);
and U1416 (N_1416,N_1244,N_1228);
or U1417 (N_1417,N_1376,N_1348);
nand U1418 (N_1418,N_1202,N_1312);
nand U1419 (N_1419,N_1285,N_1290);
or U1420 (N_1420,N_1295,N_1236);
and U1421 (N_1421,N_1345,N_1291);
or U1422 (N_1422,N_1230,N_1252);
nand U1423 (N_1423,N_1304,N_1241);
or U1424 (N_1424,N_1359,N_1374);
nand U1425 (N_1425,N_1286,N_1298);
nor U1426 (N_1426,N_1382,N_1300);
nor U1427 (N_1427,N_1352,N_1350);
nor U1428 (N_1428,N_1320,N_1356);
nor U1429 (N_1429,N_1219,N_1392);
nor U1430 (N_1430,N_1314,N_1323);
and U1431 (N_1431,N_1340,N_1380);
or U1432 (N_1432,N_1292,N_1266);
and U1433 (N_1433,N_1394,N_1229);
and U1434 (N_1434,N_1310,N_1271);
nor U1435 (N_1435,N_1265,N_1361);
and U1436 (N_1436,N_1212,N_1346);
nor U1437 (N_1437,N_1210,N_1282);
or U1438 (N_1438,N_1330,N_1397);
nor U1439 (N_1439,N_1332,N_1258);
nand U1440 (N_1440,N_1388,N_1288);
and U1441 (N_1441,N_1201,N_1343);
nor U1442 (N_1442,N_1364,N_1370);
nand U1443 (N_1443,N_1276,N_1216);
and U1444 (N_1444,N_1293,N_1367);
nand U1445 (N_1445,N_1351,N_1342);
or U1446 (N_1446,N_1249,N_1203);
or U1447 (N_1447,N_1217,N_1336);
or U1448 (N_1448,N_1319,N_1260);
and U1449 (N_1449,N_1227,N_1237);
nand U1450 (N_1450,N_1289,N_1360);
and U1451 (N_1451,N_1246,N_1270);
nand U1452 (N_1452,N_1337,N_1389);
nor U1453 (N_1453,N_1371,N_1220);
nor U1454 (N_1454,N_1262,N_1390);
nor U1455 (N_1455,N_1369,N_1387);
or U1456 (N_1456,N_1355,N_1200);
or U1457 (N_1457,N_1278,N_1333);
nand U1458 (N_1458,N_1309,N_1268);
nand U1459 (N_1459,N_1287,N_1322);
or U1460 (N_1460,N_1399,N_1315);
nand U1461 (N_1461,N_1267,N_1239);
nor U1462 (N_1462,N_1221,N_1279);
or U1463 (N_1463,N_1259,N_1206);
nor U1464 (N_1464,N_1277,N_1384);
and U1465 (N_1465,N_1224,N_1357);
or U1466 (N_1466,N_1391,N_1334);
nor U1467 (N_1467,N_1329,N_1313);
and U1468 (N_1468,N_1209,N_1331);
nand U1469 (N_1469,N_1205,N_1344);
or U1470 (N_1470,N_1235,N_1324);
nor U1471 (N_1471,N_1215,N_1254);
nor U1472 (N_1472,N_1386,N_1306);
and U1473 (N_1473,N_1327,N_1396);
and U1474 (N_1474,N_1243,N_1325);
and U1475 (N_1475,N_1318,N_1297);
or U1476 (N_1476,N_1354,N_1349);
nand U1477 (N_1477,N_1275,N_1273);
nand U1478 (N_1478,N_1338,N_1253);
and U1479 (N_1479,N_1261,N_1339);
or U1480 (N_1480,N_1316,N_1381);
or U1481 (N_1481,N_1232,N_1204);
xnor U1482 (N_1482,N_1226,N_1363);
or U1483 (N_1483,N_1247,N_1263);
and U1484 (N_1484,N_1368,N_1377);
and U1485 (N_1485,N_1317,N_1311);
and U1486 (N_1486,N_1280,N_1379);
or U1487 (N_1487,N_1358,N_1375);
nor U1488 (N_1488,N_1281,N_1395);
and U1489 (N_1489,N_1301,N_1242);
nand U1490 (N_1490,N_1366,N_1255);
or U1491 (N_1491,N_1264,N_1240);
nor U1492 (N_1492,N_1353,N_1234);
nor U1493 (N_1493,N_1272,N_1218);
or U1494 (N_1494,N_1378,N_1222);
nor U1495 (N_1495,N_1308,N_1307);
or U1496 (N_1496,N_1372,N_1284);
and U1497 (N_1497,N_1362,N_1383);
nand U1498 (N_1498,N_1294,N_1214);
or U1499 (N_1499,N_1250,N_1283);
nor U1500 (N_1500,N_1273,N_1321);
and U1501 (N_1501,N_1249,N_1396);
and U1502 (N_1502,N_1329,N_1247);
nand U1503 (N_1503,N_1333,N_1343);
or U1504 (N_1504,N_1256,N_1282);
or U1505 (N_1505,N_1355,N_1234);
nand U1506 (N_1506,N_1395,N_1383);
nand U1507 (N_1507,N_1285,N_1376);
and U1508 (N_1508,N_1297,N_1350);
xor U1509 (N_1509,N_1227,N_1347);
nor U1510 (N_1510,N_1229,N_1241);
and U1511 (N_1511,N_1268,N_1212);
nand U1512 (N_1512,N_1323,N_1229);
or U1513 (N_1513,N_1254,N_1319);
nand U1514 (N_1514,N_1275,N_1254);
nor U1515 (N_1515,N_1238,N_1315);
and U1516 (N_1516,N_1315,N_1348);
nor U1517 (N_1517,N_1305,N_1240);
or U1518 (N_1518,N_1207,N_1270);
nand U1519 (N_1519,N_1209,N_1385);
and U1520 (N_1520,N_1309,N_1371);
and U1521 (N_1521,N_1218,N_1355);
or U1522 (N_1522,N_1371,N_1311);
nor U1523 (N_1523,N_1366,N_1299);
and U1524 (N_1524,N_1392,N_1362);
nor U1525 (N_1525,N_1314,N_1282);
nor U1526 (N_1526,N_1258,N_1213);
and U1527 (N_1527,N_1221,N_1204);
and U1528 (N_1528,N_1369,N_1323);
nor U1529 (N_1529,N_1310,N_1205);
and U1530 (N_1530,N_1314,N_1385);
nand U1531 (N_1531,N_1263,N_1396);
nor U1532 (N_1532,N_1201,N_1347);
and U1533 (N_1533,N_1371,N_1224);
and U1534 (N_1534,N_1229,N_1220);
or U1535 (N_1535,N_1300,N_1303);
or U1536 (N_1536,N_1266,N_1386);
nand U1537 (N_1537,N_1292,N_1204);
nor U1538 (N_1538,N_1223,N_1237);
nand U1539 (N_1539,N_1275,N_1226);
or U1540 (N_1540,N_1305,N_1354);
and U1541 (N_1541,N_1397,N_1350);
and U1542 (N_1542,N_1321,N_1292);
and U1543 (N_1543,N_1335,N_1203);
xnor U1544 (N_1544,N_1313,N_1391);
and U1545 (N_1545,N_1352,N_1372);
nand U1546 (N_1546,N_1258,N_1222);
nor U1547 (N_1547,N_1234,N_1202);
nand U1548 (N_1548,N_1333,N_1209);
or U1549 (N_1549,N_1261,N_1201);
or U1550 (N_1550,N_1342,N_1387);
and U1551 (N_1551,N_1282,N_1238);
nor U1552 (N_1552,N_1312,N_1286);
or U1553 (N_1553,N_1324,N_1341);
or U1554 (N_1554,N_1316,N_1267);
nor U1555 (N_1555,N_1285,N_1297);
and U1556 (N_1556,N_1341,N_1258);
nand U1557 (N_1557,N_1386,N_1284);
nor U1558 (N_1558,N_1313,N_1286);
nand U1559 (N_1559,N_1381,N_1249);
or U1560 (N_1560,N_1347,N_1292);
nand U1561 (N_1561,N_1324,N_1380);
nor U1562 (N_1562,N_1268,N_1241);
or U1563 (N_1563,N_1318,N_1343);
nand U1564 (N_1564,N_1388,N_1331);
or U1565 (N_1565,N_1334,N_1389);
nand U1566 (N_1566,N_1313,N_1236);
and U1567 (N_1567,N_1360,N_1200);
nand U1568 (N_1568,N_1325,N_1301);
and U1569 (N_1569,N_1234,N_1298);
and U1570 (N_1570,N_1221,N_1367);
and U1571 (N_1571,N_1331,N_1249);
and U1572 (N_1572,N_1376,N_1292);
nor U1573 (N_1573,N_1327,N_1386);
nand U1574 (N_1574,N_1252,N_1232);
nor U1575 (N_1575,N_1248,N_1322);
nor U1576 (N_1576,N_1288,N_1263);
and U1577 (N_1577,N_1268,N_1393);
or U1578 (N_1578,N_1324,N_1326);
or U1579 (N_1579,N_1207,N_1323);
nor U1580 (N_1580,N_1302,N_1280);
nor U1581 (N_1581,N_1230,N_1210);
nor U1582 (N_1582,N_1335,N_1323);
or U1583 (N_1583,N_1346,N_1273);
nand U1584 (N_1584,N_1338,N_1341);
nand U1585 (N_1585,N_1389,N_1280);
or U1586 (N_1586,N_1397,N_1378);
nor U1587 (N_1587,N_1381,N_1386);
or U1588 (N_1588,N_1253,N_1302);
nand U1589 (N_1589,N_1344,N_1270);
nor U1590 (N_1590,N_1212,N_1313);
and U1591 (N_1591,N_1293,N_1218);
nor U1592 (N_1592,N_1365,N_1242);
nor U1593 (N_1593,N_1359,N_1210);
and U1594 (N_1594,N_1306,N_1293);
and U1595 (N_1595,N_1368,N_1248);
nand U1596 (N_1596,N_1305,N_1202);
or U1597 (N_1597,N_1270,N_1355);
or U1598 (N_1598,N_1206,N_1285);
or U1599 (N_1599,N_1339,N_1247);
nand U1600 (N_1600,N_1518,N_1487);
and U1601 (N_1601,N_1527,N_1423);
and U1602 (N_1602,N_1508,N_1550);
nand U1603 (N_1603,N_1591,N_1474);
nand U1604 (N_1604,N_1528,N_1446);
nand U1605 (N_1605,N_1429,N_1431);
or U1606 (N_1606,N_1466,N_1480);
and U1607 (N_1607,N_1561,N_1417);
nor U1608 (N_1608,N_1519,N_1441);
nor U1609 (N_1609,N_1439,N_1544);
nand U1610 (N_1610,N_1483,N_1465);
and U1611 (N_1611,N_1420,N_1411);
nor U1612 (N_1612,N_1587,N_1452);
or U1613 (N_1613,N_1581,N_1408);
nand U1614 (N_1614,N_1500,N_1486);
and U1615 (N_1615,N_1514,N_1510);
or U1616 (N_1616,N_1547,N_1576);
or U1617 (N_1617,N_1526,N_1590);
nand U1618 (N_1618,N_1492,N_1568);
nor U1619 (N_1619,N_1462,N_1574);
nand U1620 (N_1620,N_1421,N_1534);
nand U1621 (N_1621,N_1471,N_1582);
or U1622 (N_1622,N_1584,N_1554);
nor U1623 (N_1623,N_1538,N_1577);
or U1624 (N_1624,N_1541,N_1535);
or U1625 (N_1625,N_1539,N_1578);
nand U1626 (N_1626,N_1445,N_1506);
or U1627 (N_1627,N_1489,N_1498);
nand U1628 (N_1628,N_1455,N_1593);
nor U1629 (N_1629,N_1488,N_1502);
nor U1630 (N_1630,N_1545,N_1477);
nor U1631 (N_1631,N_1512,N_1548);
nor U1632 (N_1632,N_1438,N_1497);
nand U1633 (N_1633,N_1557,N_1425);
nand U1634 (N_1634,N_1469,N_1546);
or U1635 (N_1635,N_1515,N_1583);
nor U1636 (N_1636,N_1482,N_1413);
and U1637 (N_1637,N_1529,N_1428);
and U1638 (N_1638,N_1418,N_1433);
nand U1639 (N_1639,N_1569,N_1566);
nand U1640 (N_1640,N_1414,N_1406);
and U1641 (N_1641,N_1533,N_1473);
nand U1642 (N_1642,N_1559,N_1580);
and U1643 (N_1643,N_1404,N_1531);
nor U1644 (N_1644,N_1504,N_1571);
nand U1645 (N_1645,N_1437,N_1463);
or U1646 (N_1646,N_1427,N_1494);
nor U1647 (N_1647,N_1499,N_1460);
or U1648 (N_1648,N_1434,N_1560);
nor U1649 (N_1649,N_1572,N_1495);
or U1650 (N_1650,N_1505,N_1588);
and U1651 (N_1651,N_1485,N_1552);
or U1652 (N_1652,N_1467,N_1407);
and U1653 (N_1653,N_1517,N_1507);
and U1654 (N_1654,N_1573,N_1564);
nor U1655 (N_1655,N_1558,N_1450);
and U1656 (N_1656,N_1448,N_1525);
and U1657 (N_1657,N_1403,N_1530);
or U1658 (N_1658,N_1449,N_1436);
nand U1659 (N_1659,N_1589,N_1509);
and U1660 (N_1660,N_1410,N_1520);
nor U1661 (N_1661,N_1402,N_1513);
nand U1662 (N_1662,N_1444,N_1567);
or U1663 (N_1663,N_1409,N_1594);
nand U1664 (N_1664,N_1598,N_1555);
or U1665 (N_1665,N_1516,N_1522);
and U1666 (N_1666,N_1562,N_1457);
nor U1667 (N_1667,N_1579,N_1405);
nand U1668 (N_1668,N_1412,N_1586);
nor U1669 (N_1669,N_1511,N_1456);
or U1670 (N_1670,N_1481,N_1468);
nand U1671 (N_1671,N_1472,N_1521);
nor U1672 (N_1672,N_1543,N_1563);
nand U1673 (N_1673,N_1435,N_1426);
and U1674 (N_1674,N_1493,N_1575);
or U1675 (N_1675,N_1490,N_1501);
and U1676 (N_1676,N_1419,N_1553);
or U1677 (N_1677,N_1570,N_1537);
and U1678 (N_1678,N_1565,N_1416);
and U1679 (N_1679,N_1461,N_1478);
nor U1680 (N_1680,N_1447,N_1476);
or U1681 (N_1681,N_1532,N_1540);
nand U1682 (N_1682,N_1597,N_1454);
and U1683 (N_1683,N_1415,N_1585);
nor U1684 (N_1684,N_1542,N_1442);
nand U1685 (N_1685,N_1551,N_1549);
or U1686 (N_1686,N_1432,N_1523);
and U1687 (N_1687,N_1459,N_1400);
nand U1688 (N_1688,N_1440,N_1599);
or U1689 (N_1689,N_1458,N_1596);
nor U1690 (N_1690,N_1592,N_1503);
or U1691 (N_1691,N_1464,N_1595);
nor U1692 (N_1692,N_1424,N_1422);
and U1693 (N_1693,N_1475,N_1430);
and U1694 (N_1694,N_1401,N_1524);
nand U1695 (N_1695,N_1451,N_1496);
and U1696 (N_1696,N_1443,N_1479);
and U1697 (N_1697,N_1491,N_1453);
nor U1698 (N_1698,N_1484,N_1536);
and U1699 (N_1699,N_1470,N_1556);
and U1700 (N_1700,N_1469,N_1441);
or U1701 (N_1701,N_1575,N_1489);
nand U1702 (N_1702,N_1465,N_1455);
nor U1703 (N_1703,N_1406,N_1537);
nor U1704 (N_1704,N_1465,N_1595);
nor U1705 (N_1705,N_1516,N_1507);
or U1706 (N_1706,N_1524,N_1432);
or U1707 (N_1707,N_1506,N_1490);
and U1708 (N_1708,N_1593,N_1416);
or U1709 (N_1709,N_1514,N_1485);
or U1710 (N_1710,N_1592,N_1563);
or U1711 (N_1711,N_1473,N_1424);
xor U1712 (N_1712,N_1412,N_1535);
or U1713 (N_1713,N_1545,N_1458);
or U1714 (N_1714,N_1557,N_1526);
and U1715 (N_1715,N_1507,N_1465);
or U1716 (N_1716,N_1594,N_1513);
and U1717 (N_1717,N_1530,N_1432);
nand U1718 (N_1718,N_1495,N_1598);
and U1719 (N_1719,N_1491,N_1577);
nor U1720 (N_1720,N_1544,N_1572);
or U1721 (N_1721,N_1574,N_1545);
nand U1722 (N_1722,N_1506,N_1580);
or U1723 (N_1723,N_1564,N_1529);
or U1724 (N_1724,N_1543,N_1456);
nand U1725 (N_1725,N_1447,N_1441);
nor U1726 (N_1726,N_1535,N_1529);
or U1727 (N_1727,N_1535,N_1569);
or U1728 (N_1728,N_1451,N_1556);
or U1729 (N_1729,N_1485,N_1429);
or U1730 (N_1730,N_1439,N_1501);
nor U1731 (N_1731,N_1487,N_1412);
and U1732 (N_1732,N_1560,N_1425);
or U1733 (N_1733,N_1560,N_1543);
or U1734 (N_1734,N_1536,N_1565);
and U1735 (N_1735,N_1402,N_1474);
nand U1736 (N_1736,N_1483,N_1548);
nand U1737 (N_1737,N_1474,N_1425);
and U1738 (N_1738,N_1527,N_1441);
nor U1739 (N_1739,N_1522,N_1582);
or U1740 (N_1740,N_1513,N_1430);
and U1741 (N_1741,N_1591,N_1543);
nand U1742 (N_1742,N_1486,N_1432);
and U1743 (N_1743,N_1551,N_1511);
nand U1744 (N_1744,N_1510,N_1447);
or U1745 (N_1745,N_1441,N_1500);
and U1746 (N_1746,N_1572,N_1524);
or U1747 (N_1747,N_1505,N_1562);
or U1748 (N_1748,N_1413,N_1475);
nor U1749 (N_1749,N_1430,N_1400);
nor U1750 (N_1750,N_1556,N_1568);
nand U1751 (N_1751,N_1514,N_1547);
nand U1752 (N_1752,N_1425,N_1447);
nor U1753 (N_1753,N_1442,N_1489);
nand U1754 (N_1754,N_1467,N_1587);
and U1755 (N_1755,N_1587,N_1407);
nor U1756 (N_1756,N_1528,N_1525);
nor U1757 (N_1757,N_1593,N_1438);
nor U1758 (N_1758,N_1572,N_1461);
or U1759 (N_1759,N_1550,N_1456);
or U1760 (N_1760,N_1564,N_1418);
xnor U1761 (N_1761,N_1499,N_1493);
and U1762 (N_1762,N_1599,N_1505);
and U1763 (N_1763,N_1476,N_1545);
or U1764 (N_1764,N_1575,N_1437);
or U1765 (N_1765,N_1538,N_1491);
nand U1766 (N_1766,N_1517,N_1473);
or U1767 (N_1767,N_1454,N_1482);
or U1768 (N_1768,N_1539,N_1459);
or U1769 (N_1769,N_1468,N_1442);
nand U1770 (N_1770,N_1592,N_1482);
nor U1771 (N_1771,N_1409,N_1577);
nor U1772 (N_1772,N_1443,N_1560);
and U1773 (N_1773,N_1406,N_1419);
and U1774 (N_1774,N_1562,N_1512);
nor U1775 (N_1775,N_1532,N_1519);
or U1776 (N_1776,N_1543,N_1478);
nor U1777 (N_1777,N_1408,N_1557);
or U1778 (N_1778,N_1541,N_1523);
and U1779 (N_1779,N_1593,N_1459);
and U1780 (N_1780,N_1527,N_1558);
nor U1781 (N_1781,N_1429,N_1537);
and U1782 (N_1782,N_1465,N_1546);
nand U1783 (N_1783,N_1558,N_1590);
or U1784 (N_1784,N_1528,N_1504);
nor U1785 (N_1785,N_1432,N_1528);
and U1786 (N_1786,N_1598,N_1433);
nand U1787 (N_1787,N_1585,N_1401);
or U1788 (N_1788,N_1458,N_1409);
nor U1789 (N_1789,N_1587,N_1422);
nand U1790 (N_1790,N_1507,N_1403);
or U1791 (N_1791,N_1473,N_1528);
nor U1792 (N_1792,N_1419,N_1424);
nand U1793 (N_1793,N_1430,N_1583);
xnor U1794 (N_1794,N_1525,N_1465);
nor U1795 (N_1795,N_1486,N_1400);
nor U1796 (N_1796,N_1515,N_1543);
nor U1797 (N_1797,N_1515,N_1560);
nand U1798 (N_1798,N_1466,N_1507);
nor U1799 (N_1799,N_1451,N_1567);
nor U1800 (N_1800,N_1642,N_1675);
nor U1801 (N_1801,N_1612,N_1763);
nor U1802 (N_1802,N_1738,N_1646);
and U1803 (N_1803,N_1796,N_1783);
nand U1804 (N_1804,N_1741,N_1739);
nor U1805 (N_1805,N_1755,N_1600);
or U1806 (N_1806,N_1672,N_1784);
or U1807 (N_1807,N_1635,N_1699);
or U1808 (N_1808,N_1713,N_1614);
nor U1809 (N_1809,N_1789,N_1715);
or U1810 (N_1810,N_1643,N_1712);
or U1811 (N_1811,N_1762,N_1648);
nand U1812 (N_1812,N_1621,N_1616);
and U1813 (N_1813,N_1742,N_1617);
or U1814 (N_1814,N_1744,N_1702);
nor U1815 (N_1815,N_1627,N_1787);
nand U1816 (N_1816,N_1639,N_1706);
nor U1817 (N_1817,N_1710,N_1774);
nor U1818 (N_1818,N_1729,N_1606);
xor U1819 (N_1819,N_1775,N_1727);
and U1820 (N_1820,N_1740,N_1694);
or U1821 (N_1821,N_1633,N_1632);
nand U1822 (N_1822,N_1743,N_1749);
nor U1823 (N_1823,N_1766,N_1652);
or U1824 (N_1824,N_1665,N_1769);
and U1825 (N_1825,N_1625,N_1777);
nand U1826 (N_1826,N_1771,N_1683);
nor U1827 (N_1827,N_1759,N_1797);
and U1828 (N_1828,N_1676,N_1737);
and U1829 (N_1829,N_1658,N_1731);
and U1830 (N_1830,N_1619,N_1747);
nor U1831 (N_1831,N_1767,N_1788);
or U1832 (N_1832,N_1640,N_1605);
or U1833 (N_1833,N_1768,N_1705);
and U1834 (N_1834,N_1781,N_1692);
or U1835 (N_1835,N_1723,N_1650);
and U1836 (N_1836,N_1611,N_1687);
or U1837 (N_1837,N_1779,N_1603);
nand U1838 (N_1838,N_1657,N_1645);
nor U1839 (N_1839,N_1656,N_1798);
or U1840 (N_1840,N_1682,N_1716);
or U1841 (N_1841,N_1709,N_1610);
nand U1842 (N_1842,N_1688,N_1756);
nand U1843 (N_1843,N_1677,N_1717);
nor U1844 (N_1844,N_1689,N_1753);
nand U1845 (N_1845,N_1636,N_1602);
nand U1846 (N_1846,N_1674,N_1719);
nand U1847 (N_1847,N_1733,N_1697);
or U1848 (N_1848,N_1649,N_1748);
and U1849 (N_1849,N_1714,N_1700);
or U1850 (N_1850,N_1698,N_1790);
nor U1851 (N_1851,N_1654,N_1628);
or U1852 (N_1852,N_1780,N_1662);
or U1853 (N_1853,N_1693,N_1792);
nand U1854 (N_1854,N_1609,N_1680);
or U1855 (N_1855,N_1695,N_1604);
or U1856 (N_1856,N_1765,N_1673);
nor U1857 (N_1857,N_1696,N_1623);
nor U1858 (N_1858,N_1791,N_1690);
and U1859 (N_1859,N_1685,N_1746);
and U1860 (N_1860,N_1655,N_1663);
nand U1861 (N_1861,N_1708,N_1618);
nor U1862 (N_1862,N_1730,N_1678);
nand U1863 (N_1863,N_1671,N_1728);
nand U1864 (N_1864,N_1726,N_1638);
and U1865 (N_1865,N_1626,N_1659);
nor U1866 (N_1866,N_1770,N_1637);
nor U1867 (N_1867,N_1707,N_1653);
nand U1868 (N_1868,N_1778,N_1745);
nand U1869 (N_1869,N_1799,N_1666);
or U1870 (N_1870,N_1629,N_1615);
or U1871 (N_1871,N_1622,N_1721);
nand U1872 (N_1872,N_1647,N_1681);
nor U1873 (N_1873,N_1776,N_1704);
nand U1874 (N_1874,N_1794,N_1686);
or U1875 (N_1875,N_1711,N_1684);
and U1876 (N_1876,N_1601,N_1608);
and U1877 (N_1877,N_1725,N_1751);
or U1878 (N_1878,N_1651,N_1691);
nor U1879 (N_1879,N_1773,N_1644);
nor U1880 (N_1880,N_1764,N_1722);
nand U1881 (N_1881,N_1786,N_1634);
nand U1882 (N_1882,N_1701,N_1624);
nor U1883 (N_1883,N_1732,N_1718);
and U1884 (N_1884,N_1757,N_1607);
nand U1885 (N_1885,N_1720,N_1641);
or U1886 (N_1886,N_1793,N_1761);
nand U1887 (N_1887,N_1703,N_1661);
or U1888 (N_1888,N_1734,N_1735);
nor U1889 (N_1889,N_1724,N_1630);
nand U1890 (N_1890,N_1785,N_1772);
nor U1891 (N_1891,N_1613,N_1736);
nand U1892 (N_1892,N_1620,N_1758);
and U1893 (N_1893,N_1750,N_1752);
or U1894 (N_1894,N_1754,N_1795);
or U1895 (N_1895,N_1679,N_1669);
nor U1896 (N_1896,N_1668,N_1670);
and U1897 (N_1897,N_1660,N_1760);
nand U1898 (N_1898,N_1631,N_1667);
and U1899 (N_1899,N_1664,N_1782);
and U1900 (N_1900,N_1722,N_1626);
nor U1901 (N_1901,N_1765,N_1634);
and U1902 (N_1902,N_1692,N_1616);
nand U1903 (N_1903,N_1642,N_1645);
or U1904 (N_1904,N_1773,N_1793);
or U1905 (N_1905,N_1746,N_1795);
nor U1906 (N_1906,N_1613,N_1653);
nor U1907 (N_1907,N_1638,N_1606);
and U1908 (N_1908,N_1713,N_1650);
and U1909 (N_1909,N_1750,N_1605);
nor U1910 (N_1910,N_1628,N_1694);
or U1911 (N_1911,N_1641,N_1656);
and U1912 (N_1912,N_1682,N_1644);
nor U1913 (N_1913,N_1790,N_1797);
nand U1914 (N_1914,N_1732,N_1695);
or U1915 (N_1915,N_1605,N_1745);
and U1916 (N_1916,N_1616,N_1618);
nand U1917 (N_1917,N_1736,N_1660);
or U1918 (N_1918,N_1760,N_1723);
and U1919 (N_1919,N_1737,N_1610);
or U1920 (N_1920,N_1653,N_1755);
nand U1921 (N_1921,N_1616,N_1797);
or U1922 (N_1922,N_1714,N_1675);
or U1923 (N_1923,N_1719,N_1687);
nand U1924 (N_1924,N_1756,N_1750);
nand U1925 (N_1925,N_1609,N_1782);
nand U1926 (N_1926,N_1635,N_1625);
or U1927 (N_1927,N_1792,N_1727);
and U1928 (N_1928,N_1640,N_1723);
or U1929 (N_1929,N_1726,N_1657);
nand U1930 (N_1930,N_1718,N_1766);
nor U1931 (N_1931,N_1614,N_1759);
nor U1932 (N_1932,N_1779,N_1709);
nor U1933 (N_1933,N_1642,N_1612);
nand U1934 (N_1934,N_1770,N_1785);
nor U1935 (N_1935,N_1719,N_1662);
nor U1936 (N_1936,N_1770,N_1780);
or U1937 (N_1937,N_1734,N_1666);
nand U1938 (N_1938,N_1709,N_1673);
or U1939 (N_1939,N_1614,N_1640);
nor U1940 (N_1940,N_1796,N_1657);
xor U1941 (N_1941,N_1652,N_1716);
or U1942 (N_1942,N_1727,N_1746);
nor U1943 (N_1943,N_1638,N_1719);
or U1944 (N_1944,N_1795,N_1652);
or U1945 (N_1945,N_1619,N_1790);
and U1946 (N_1946,N_1780,N_1684);
nand U1947 (N_1947,N_1625,N_1617);
nor U1948 (N_1948,N_1670,N_1752);
and U1949 (N_1949,N_1608,N_1605);
nand U1950 (N_1950,N_1713,N_1646);
nor U1951 (N_1951,N_1750,N_1723);
nand U1952 (N_1952,N_1794,N_1758);
nand U1953 (N_1953,N_1754,N_1629);
or U1954 (N_1954,N_1611,N_1712);
nand U1955 (N_1955,N_1693,N_1763);
or U1956 (N_1956,N_1638,N_1728);
nor U1957 (N_1957,N_1769,N_1631);
nand U1958 (N_1958,N_1671,N_1757);
and U1959 (N_1959,N_1731,N_1757);
and U1960 (N_1960,N_1614,N_1631);
and U1961 (N_1961,N_1769,N_1780);
or U1962 (N_1962,N_1770,N_1713);
or U1963 (N_1963,N_1757,N_1792);
xnor U1964 (N_1964,N_1622,N_1617);
nor U1965 (N_1965,N_1796,N_1731);
or U1966 (N_1966,N_1667,N_1611);
nor U1967 (N_1967,N_1629,N_1610);
and U1968 (N_1968,N_1647,N_1630);
nor U1969 (N_1969,N_1751,N_1651);
nor U1970 (N_1970,N_1603,N_1719);
nor U1971 (N_1971,N_1752,N_1606);
and U1972 (N_1972,N_1693,N_1746);
nor U1973 (N_1973,N_1731,N_1752);
nor U1974 (N_1974,N_1794,N_1690);
or U1975 (N_1975,N_1659,N_1650);
and U1976 (N_1976,N_1605,N_1761);
and U1977 (N_1977,N_1755,N_1643);
nand U1978 (N_1978,N_1649,N_1618);
and U1979 (N_1979,N_1652,N_1718);
and U1980 (N_1980,N_1752,N_1733);
and U1981 (N_1981,N_1670,N_1749);
or U1982 (N_1982,N_1653,N_1790);
nand U1983 (N_1983,N_1654,N_1611);
or U1984 (N_1984,N_1656,N_1631);
and U1985 (N_1985,N_1621,N_1778);
and U1986 (N_1986,N_1629,N_1605);
and U1987 (N_1987,N_1699,N_1695);
or U1988 (N_1988,N_1733,N_1616);
nor U1989 (N_1989,N_1634,N_1787);
and U1990 (N_1990,N_1711,N_1772);
nand U1991 (N_1991,N_1653,N_1765);
or U1992 (N_1992,N_1769,N_1716);
nor U1993 (N_1993,N_1636,N_1708);
nor U1994 (N_1994,N_1715,N_1636);
nor U1995 (N_1995,N_1729,N_1645);
nand U1996 (N_1996,N_1727,N_1694);
and U1997 (N_1997,N_1696,N_1772);
and U1998 (N_1998,N_1608,N_1771);
nor U1999 (N_1999,N_1621,N_1726);
or U2000 (N_2000,N_1848,N_1879);
and U2001 (N_2001,N_1885,N_1981);
or U2002 (N_2002,N_1933,N_1810);
or U2003 (N_2003,N_1955,N_1833);
xor U2004 (N_2004,N_1807,N_1866);
nand U2005 (N_2005,N_1819,N_1898);
nand U2006 (N_2006,N_1859,N_1985);
nand U2007 (N_2007,N_1944,N_1992);
or U2008 (N_2008,N_1871,N_1946);
nor U2009 (N_2009,N_1897,N_1987);
nor U2010 (N_2010,N_1829,N_1989);
nor U2011 (N_2011,N_1801,N_1821);
nand U2012 (N_2012,N_1974,N_1941);
or U2013 (N_2013,N_1943,N_1969);
nand U2014 (N_2014,N_1891,N_1870);
nor U2015 (N_2015,N_1945,N_1972);
and U2016 (N_2016,N_1834,N_1906);
nand U2017 (N_2017,N_1966,N_1903);
or U2018 (N_2018,N_1922,N_1934);
or U2019 (N_2019,N_1947,N_1917);
or U2020 (N_2020,N_1949,N_1867);
nor U2021 (N_2021,N_1800,N_1875);
nand U2022 (N_2022,N_1900,N_1827);
and U2023 (N_2023,N_1923,N_1993);
nand U2024 (N_2024,N_1872,N_1857);
nand U2025 (N_2025,N_1911,N_1953);
and U2026 (N_2026,N_1977,N_1811);
and U2027 (N_2027,N_1995,N_1901);
and U2028 (N_2028,N_1828,N_1958);
nand U2029 (N_2029,N_1825,N_1861);
nor U2030 (N_2030,N_1932,N_1889);
or U2031 (N_2031,N_1840,N_1920);
or U2032 (N_2032,N_1845,N_1978);
and U2033 (N_2033,N_1971,N_1930);
nand U2034 (N_2034,N_1914,N_1976);
or U2035 (N_2035,N_1880,N_1893);
or U2036 (N_2036,N_1817,N_1869);
and U2037 (N_2037,N_1999,N_1863);
nor U2038 (N_2038,N_1878,N_1950);
nand U2039 (N_2039,N_1894,N_1855);
and U2040 (N_2040,N_1803,N_1935);
nand U2041 (N_2041,N_1938,N_1998);
nand U2042 (N_2042,N_1984,N_1983);
and U2043 (N_2043,N_1862,N_1826);
or U2044 (N_2044,N_1838,N_1886);
or U2045 (N_2045,N_1994,N_1846);
or U2046 (N_2046,N_1888,N_1970);
and U2047 (N_2047,N_1876,N_1830);
and U2048 (N_2048,N_1837,N_1921);
or U2049 (N_2049,N_1956,N_1865);
nor U2050 (N_2050,N_1925,N_1823);
nand U2051 (N_2051,N_1882,N_1832);
or U2052 (N_2052,N_1982,N_1942);
nand U2053 (N_2053,N_1818,N_1909);
nand U2054 (N_2054,N_1836,N_1802);
or U2055 (N_2055,N_1961,N_1812);
nand U2056 (N_2056,N_1814,N_1899);
or U2057 (N_2057,N_1931,N_1990);
and U2058 (N_2058,N_1937,N_1831);
and U2059 (N_2059,N_1820,N_1868);
nand U2060 (N_2060,N_1928,N_1874);
and U2061 (N_2061,N_1915,N_1926);
and U2062 (N_2062,N_1884,N_1940);
nor U2063 (N_2063,N_1809,N_1912);
xor U2064 (N_2064,N_1858,N_1905);
nor U2065 (N_2065,N_1959,N_1996);
nor U2066 (N_2066,N_1948,N_1856);
or U2067 (N_2067,N_1997,N_1951);
or U2068 (N_2068,N_1939,N_1853);
or U2069 (N_2069,N_1919,N_1895);
or U2070 (N_2070,N_1881,N_1849);
nor U2071 (N_2071,N_1822,N_1815);
nand U2072 (N_2072,N_1887,N_1973);
or U2073 (N_2073,N_1883,N_1988);
nand U2074 (N_2074,N_1924,N_1907);
or U2075 (N_2075,N_1844,N_1890);
nand U2076 (N_2076,N_1960,N_1804);
and U2077 (N_2077,N_1929,N_1963);
and U2078 (N_2078,N_1908,N_1980);
nor U2079 (N_2079,N_1916,N_1927);
nor U2080 (N_2080,N_1986,N_1806);
or U2081 (N_2081,N_1892,N_1965);
nand U2082 (N_2082,N_1841,N_1913);
or U2083 (N_2083,N_1936,N_1864);
nor U2084 (N_2084,N_1860,N_1877);
nand U2085 (N_2085,N_1918,N_1843);
and U2086 (N_2086,N_1805,N_1850);
and U2087 (N_2087,N_1851,N_1842);
nand U2088 (N_2088,N_1957,N_1835);
or U2089 (N_2089,N_1968,N_1964);
and U2090 (N_2090,N_1902,N_1816);
nor U2091 (N_2091,N_1847,N_1813);
nand U2092 (N_2092,N_1854,N_1954);
nand U2093 (N_2093,N_1991,N_1839);
nand U2094 (N_2094,N_1852,N_1824);
and U2095 (N_2095,N_1952,N_1896);
nand U2096 (N_2096,N_1904,N_1962);
nand U2097 (N_2097,N_1873,N_1979);
nand U2098 (N_2098,N_1975,N_1967);
or U2099 (N_2099,N_1910,N_1808);
nand U2100 (N_2100,N_1996,N_1953);
nor U2101 (N_2101,N_1932,N_1946);
or U2102 (N_2102,N_1897,N_1993);
nand U2103 (N_2103,N_1942,N_1922);
nand U2104 (N_2104,N_1988,N_1872);
nand U2105 (N_2105,N_1903,N_1876);
nand U2106 (N_2106,N_1939,N_1816);
nand U2107 (N_2107,N_1942,N_1888);
nand U2108 (N_2108,N_1902,N_1866);
nor U2109 (N_2109,N_1913,N_1852);
and U2110 (N_2110,N_1818,N_1811);
nor U2111 (N_2111,N_1888,N_1836);
and U2112 (N_2112,N_1855,N_1945);
nand U2113 (N_2113,N_1844,N_1869);
nand U2114 (N_2114,N_1878,N_1846);
nor U2115 (N_2115,N_1903,N_1867);
xnor U2116 (N_2116,N_1934,N_1890);
nand U2117 (N_2117,N_1859,N_1818);
and U2118 (N_2118,N_1962,N_1907);
nand U2119 (N_2119,N_1842,N_1878);
nand U2120 (N_2120,N_1816,N_1854);
nor U2121 (N_2121,N_1867,N_1940);
or U2122 (N_2122,N_1873,N_1846);
and U2123 (N_2123,N_1854,N_1946);
nor U2124 (N_2124,N_1840,N_1878);
or U2125 (N_2125,N_1818,N_1866);
and U2126 (N_2126,N_1806,N_1994);
or U2127 (N_2127,N_1952,N_1919);
or U2128 (N_2128,N_1879,N_1972);
and U2129 (N_2129,N_1938,N_1820);
or U2130 (N_2130,N_1921,N_1911);
nor U2131 (N_2131,N_1858,N_1935);
nor U2132 (N_2132,N_1931,N_1991);
nor U2133 (N_2133,N_1977,N_1837);
nand U2134 (N_2134,N_1936,N_1945);
xnor U2135 (N_2135,N_1879,N_1981);
and U2136 (N_2136,N_1838,N_1892);
nor U2137 (N_2137,N_1883,N_1860);
xor U2138 (N_2138,N_1846,N_1972);
nand U2139 (N_2139,N_1877,N_1955);
and U2140 (N_2140,N_1837,N_1989);
nand U2141 (N_2141,N_1949,N_1906);
nand U2142 (N_2142,N_1801,N_1830);
or U2143 (N_2143,N_1930,N_1904);
nor U2144 (N_2144,N_1996,N_1964);
and U2145 (N_2145,N_1900,N_1929);
and U2146 (N_2146,N_1965,N_1819);
and U2147 (N_2147,N_1895,N_1889);
nand U2148 (N_2148,N_1922,N_1958);
nor U2149 (N_2149,N_1858,N_1876);
or U2150 (N_2150,N_1982,N_1969);
and U2151 (N_2151,N_1929,N_1920);
nand U2152 (N_2152,N_1973,N_1880);
nor U2153 (N_2153,N_1893,N_1805);
and U2154 (N_2154,N_1804,N_1834);
nand U2155 (N_2155,N_1854,N_1940);
nor U2156 (N_2156,N_1935,N_1998);
or U2157 (N_2157,N_1894,N_1896);
nor U2158 (N_2158,N_1878,N_1907);
nor U2159 (N_2159,N_1867,N_1945);
and U2160 (N_2160,N_1899,N_1878);
and U2161 (N_2161,N_1823,N_1818);
and U2162 (N_2162,N_1895,N_1955);
or U2163 (N_2163,N_1984,N_1852);
or U2164 (N_2164,N_1906,N_1808);
and U2165 (N_2165,N_1982,N_1801);
and U2166 (N_2166,N_1842,N_1974);
or U2167 (N_2167,N_1988,N_1894);
nor U2168 (N_2168,N_1919,N_1908);
and U2169 (N_2169,N_1817,N_1807);
nand U2170 (N_2170,N_1933,N_1946);
or U2171 (N_2171,N_1999,N_1936);
nand U2172 (N_2172,N_1827,N_1965);
nor U2173 (N_2173,N_1845,N_1873);
and U2174 (N_2174,N_1806,N_1902);
nand U2175 (N_2175,N_1988,N_1993);
or U2176 (N_2176,N_1817,N_1858);
nor U2177 (N_2177,N_1897,N_1853);
or U2178 (N_2178,N_1889,N_1945);
or U2179 (N_2179,N_1920,N_1987);
nor U2180 (N_2180,N_1869,N_1994);
nand U2181 (N_2181,N_1889,N_1869);
nor U2182 (N_2182,N_1889,N_1971);
and U2183 (N_2183,N_1886,N_1820);
and U2184 (N_2184,N_1843,N_1996);
and U2185 (N_2185,N_1875,N_1828);
nor U2186 (N_2186,N_1879,N_1855);
nand U2187 (N_2187,N_1981,N_1978);
and U2188 (N_2188,N_1903,N_1999);
and U2189 (N_2189,N_1873,N_1818);
nand U2190 (N_2190,N_1891,N_1924);
or U2191 (N_2191,N_1886,N_1827);
or U2192 (N_2192,N_1958,N_1921);
nand U2193 (N_2193,N_1980,N_1828);
or U2194 (N_2194,N_1814,N_1977);
nand U2195 (N_2195,N_1922,N_1878);
and U2196 (N_2196,N_1972,N_1873);
nor U2197 (N_2197,N_1939,N_1886);
nand U2198 (N_2198,N_1914,N_1850);
or U2199 (N_2199,N_1966,N_1958);
and U2200 (N_2200,N_2132,N_2049);
nor U2201 (N_2201,N_2166,N_2156);
and U2202 (N_2202,N_2163,N_2088);
nor U2203 (N_2203,N_2004,N_2152);
nand U2204 (N_2204,N_2170,N_2102);
or U2205 (N_2205,N_2181,N_2172);
nand U2206 (N_2206,N_2182,N_2120);
or U2207 (N_2207,N_2020,N_2112);
nor U2208 (N_2208,N_2174,N_2150);
nand U2209 (N_2209,N_2012,N_2117);
nor U2210 (N_2210,N_2057,N_2127);
or U2211 (N_2211,N_2066,N_2041);
and U2212 (N_2212,N_2128,N_2025);
and U2213 (N_2213,N_2177,N_2090);
nand U2214 (N_2214,N_2139,N_2089);
or U2215 (N_2215,N_2035,N_2131);
and U2216 (N_2216,N_2153,N_2019);
nor U2217 (N_2217,N_2155,N_2122);
and U2218 (N_2218,N_2038,N_2101);
nor U2219 (N_2219,N_2017,N_2058);
nand U2220 (N_2220,N_2029,N_2118);
nand U2221 (N_2221,N_2055,N_2093);
nand U2222 (N_2222,N_2162,N_2081);
nand U2223 (N_2223,N_2107,N_2008);
or U2224 (N_2224,N_2042,N_2046);
and U2225 (N_2225,N_2037,N_2005);
nor U2226 (N_2226,N_2065,N_2098);
nand U2227 (N_2227,N_2073,N_2068);
nand U2228 (N_2228,N_2087,N_2146);
nand U2229 (N_2229,N_2144,N_2056);
or U2230 (N_2230,N_2115,N_2064);
and U2231 (N_2231,N_2001,N_2157);
nand U2232 (N_2232,N_2014,N_2100);
and U2233 (N_2233,N_2135,N_2137);
and U2234 (N_2234,N_2136,N_2036);
or U2235 (N_2235,N_2133,N_2124);
or U2236 (N_2236,N_2032,N_2193);
nand U2237 (N_2237,N_2197,N_2050);
nor U2238 (N_2238,N_2013,N_2175);
and U2239 (N_2239,N_2160,N_2018);
and U2240 (N_2240,N_2159,N_2097);
or U2241 (N_2241,N_2126,N_2104);
and U2242 (N_2242,N_2059,N_2026);
nor U2243 (N_2243,N_2173,N_2063);
nand U2244 (N_2244,N_2007,N_2189);
nand U2245 (N_2245,N_2084,N_2141);
nand U2246 (N_2246,N_2192,N_2062);
or U2247 (N_2247,N_2054,N_2031);
nand U2248 (N_2248,N_2143,N_2096);
and U2249 (N_2249,N_2142,N_2138);
or U2250 (N_2250,N_2196,N_2176);
nand U2251 (N_2251,N_2076,N_2185);
or U2252 (N_2252,N_2109,N_2024);
or U2253 (N_2253,N_2186,N_2078);
or U2254 (N_2254,N_2129,N_2198);
and U2255 (N_2255,N_2022,N_2034);
or U2256 (N_2256,N_2040,N_2003);
and U2257 (N_2257,N_2069,N_2091);
or U2258 (N_2258,N_2010,N_2119);
and U2259 (N_2259,N_2080,N_2171);
nand U2260 (N_2260,N_2154,N_2116);
and U2261 (N_2261,N_2039,N_2106);
or U2262 (N_2262,N_2067,N_2082);
or U2263 (N_2263,N_2021,N_2016);
and U2264 (N_2264,N_2147,N_2103);
and U2265 (N_2265,N_2167,N_2077);
nor U2266 (N_2266,N_2114,N_2072);
or U2267 (N_2267,N_2009,N_2151);
and U2268 (N_2268,N_2187,N_2190);
nand U2269 (N_2269,N_2092,N_2149);
and U2270 (N_2270,N_2180,N_2111);
nor U2271 (N_2271,N_2178,N_2121);
and U2272 (N_2272,N_2195,N_2113);
or U2273 (N_2273,N_2134,N_2071);
and U2274 (N_2274,N_2052,N_2086);
and U2275 (N_2275,N_2075,N_2051);
xnor U2276 (N_2276,N_2169,N_2099);
or U2277 (N_2277,N_2125,N_2123);
and U2278 (N_2278,N_2002,N_2085);
and U2279 (N_2279,N_2148,N_2033);
nor U2280 (N_2280,N_2061,N_2095);
and U2281 (N_2281,N_2105,N_2079);
nand U2282 (N_2282,N_2047,N_2184);
nand U2283 (N_2283,N_2199,N_2060);
xnor U2284 (N_2284,N_2158,N_2094);
or U2285 (N_2285,N_2130,N_2191);
nor U2286 (N_2286,N_2006,N_2044);
nor U2287 (N_2287,N_2194,N_2000);
nand U2288 (N_2288,N_2145,N_2161);
and U2289 (N_2289,N_2011,N_2030);
or U2290 (N_2290,N_2048,N_2188);
or U2291 (N_2291,N_2165,N_2028);
and U2292 (N_2292,N_2108,N_2164);
or U2293 (N_2293,N_2043,N_2045);
nor U2294 (N_2294,N_2070,N_2053);
and U2295 (N_2295,N_2074,N_2179);
nor U2296 (N_2296,N_2027,N_2015);
or U2297 (N_2297,N_2140,N_2183);
nand U2298 (N_2298,N_2023,N_2110);
or U2299 (N_2299,N_2083,N_2168);
or U2300 (N_2300,N_2052,N_2060);
or U2301 (N_2301,N_2030,N_2066);
nand U2302 (N_2302,N_2099,N_2166);
and U2303 (N_2303,N_2155,N_2061);
nor U2304 (N_2304,N_2099,N_2197);
nor U2305 (N_2305,N_2115,N_2075);
and U2306 (N_2306,N_2034,N_2014);
nor U2307 (N_2307,N_2030,N_2055);
nor U2308 (N_2308,N_2043,N_2196);
xor U2309 (N_2309,N_2073,N_2122);
and U2310 (N_2310,N_2001,N_2134);
and U2311 (N_2311,N_2035,N_2082);
nand U2312 (N_2312,N_2086,N_2091);
nor U2313 (N_2313,N_2000,N_2161);
and U2314 (N_2314,N_2058,N_2160);
nor U2315 (N_2315,N_2112,N_2095);
or U2316 (N_2316,N_2183,N_2130);
or U2317 (N_2317,N_2055,N_2191);
or U2318 (N_2318,N_2166,N_2153);
or U2319 (N_2319,N_2106,N_2183);
nand U2320 (N_2320,N_2098,N_2177);
nor U2321 (N_2321,N_2155,N_2055);
and U2322 (N_2322,N_2129,N_2167);
nand U2323 (N_2323,N_2196,N_2038);
and U2324 (N_2324,N_2030,N_2058);
nand U2325 (N_2325,N_2109,N_2081);
and U2326 (N_2326,N_2131,N_2068);
nand U2327 (N_2327,N_2050,N_2053);
nor U2328 (N_2328,N_2050,N_2021);
or U2329 (N_2329,N_2119,N_2012);
or U2330 (N_2330,N_2015,N_2123);
and U2331 (N_2331,N_2059,N_2122);
or U2332 (N_2332,N_2106,N_2041);
nor U2333 (N_2333,N_2134,N_2123);
nor U2334 (N_2334,N_2094,N_2062);
or U2335 (N_2335,N_2025,N_2058);
nand U2336 (N_2336,N_2190,N_2078);
and U2337 (N_2337,N_2154,N_2113);
nand U2338 (N_2338,N_2193,N_2182);
or U2339 (N_2339,N_2081,N_2138);
nor U2340 (N_2340,N_2079,N_2038);
and U2341 (N_2341,N_2001,N_2077);
xor U2342 (N_2342,N_2094,N_2095);
and U2343 (N_2343,N_2135,N_2129);
and U2344 (N_2344,N_2146,N_2179);
and U2345 (N_2345,N_2010,N_2199);
nor U2346 (N_2346,N_2041,N_2137);
nor U2347 (N_2347,N_2107,N_2033);
or U2348 (N_2348,N_2062,N_2069);
and U2349 (N_2349,N_2162,N_2137);
nor U2350 (N_2350,N_2065,N_2090);
or U2351 (N_2351,N_2026,N_2168);
nor U2352 (N_2352,N_2130,N_2128);
and U2353 (N_2353,N_2024,N_2103);
or U2354 (N_2354,N_2038,N_2064);
and U2355 (N_2355,N_2084,N_2042);
nand U2356 (N_2356,N_2100,N_2007);
xnor U2357 (N_2357,N_2082,N_2063);
or U2358 (N_2358,N_2180,N_2130);
or U2359 (N_2359,N_2140,N_2101);
nand U2360 (N_2360,N_2064,N_2020);
or U2361 (N_2361,N_2105,N_2052);
or U2362 (N_2362,N_2008,N_2122);
and U2363 (N_2363,N_2141,N_2002);
and U2364 (N_2364,N_2196,N_2124);
nor U2365 (N_2365,N_2117,N_2054);
or U2366 (N_2366,N_2091,N_2075);
nand U2367 (N_2367,N_2038,N_2035);
or U2368 (N_2368,N_2122,N_2039);
nand U2369 (N_2369,N_2191,N_2156);
or U2370 (N_2370,N_2049,N_2001);
or U2371 (N_2371,N_2109,N_2193);
nor U2372 (N_2372,N_2149,N_2047);
nor U2373 (N_2373,N_2048,N_2081);
and U2374 (N_2374,N_2019,N_2115);
or U2375 (N_2375,N_2086,N_2174);
or U2376 (N_2376,N_2095,N_2160);
and U2377 (N_2377,N_2187,N_2068);
nand U2378 (N_2378,N_2144,N_2195);
nand U2379 (N_2379,N_2088,N_2019);
nor U2380 (N_2380,N_2093,N_2010);
nor U2381 (N_2381,N_2064,N_2109);
and U2382 (N_2382,N_2085,N_2190);
nand U2383 (N_2383,N_2115,N_2044);
nor U2384 (N_2384,N_2016,N_2115);
and U2385 (N_2385,N_2017,N_2124);
nor U2386 (N_2386,N_2064,N_2119);
nand U2387 (N_2387,N_2042,N_2016);
or U2388 (N_2388,N_2005,N_2169);
nand U2389 (N_2389,N_2016,N_2084);
or U2390 (N_2390,N_2135,N_2097);
nor U2391 (N_2391,N_2153,N_2116);
nand U2392 (N_2392,N_2060,N_2140);
nand U2393 (N_2393,N_2080,N_2011);
nand U2394 (N_2394,N_2117,N_2016);
and U2395 (N_2395,N_2041,N_2158);
or U2396 (N_2396,N_2159,N_2197);
nor U2397 (N_2397,N_2151,N_2195);
nand U2398 (N_2398,N_2119,N_2175);
nor U2399 (N_2399,N_2189,N_2018);
and U2400 (N_2400,N_2329,N_2201);
or U2401 (N_2401,N_2225,N_2279);
or U2402 (N_2402,N_2378,N_2390);
xor U2403 (N_2403,N_2376,N_2289);
and U2404 (N_2404,N_2313,N_2317);
nor U2405 (N_2405,N_2364,N_2354);
nand U2406 (N_2406,N_2224,N_2291);
and U2407 (N_2407,N_2310,N_2237);
and U2408 (N_2408,N_2287,N_2311);
or U2409 (N_2409,N_2211,N_2315);
and U2410 (N_2410,N_2242,N_2300);
and U2411 (N_2411,N_2223,N_2268);
and U2412 (N_2412,N_2233,N_2236);
nand U2413 (N_2413,N_2336,N_2254);
and U2414 (N_2414,N_2320,N_2245);
or U2415 (N_2415,N_2202,N_2206);
nand U2416 (N_2416,N_2334,N_2399);
nand U2417 (N_2417,N_2257,N_2398);
or U2418 (N_2418,N_2288,N_2340);
and U2419 (N_2419,N_2278,N_2203);
nor U2420 (N_2420,N_2333,N_2284);
and U2421 (N_2421,N_2234,N_2301);
or U2422 (N_2422,N_2360,N_2273);
nor U2423 (N_2423,N_2235,N_2316);
nor U2424 (N_2424,N_2297,N_2389);
and U2425 (N_2425,N_2290,N_2332);
or U2426 (N_2426,N_2325,N_2298);
and U2427 (N_2427,N_2270,N_2255);
nand U2428 (N_2428,N_2261,N_2339);
and U2429 (N_2429,N_2260,N_2210);
nor U2430 (N_2430,N_2209,N_2356);
nand U2431 (N_2431,N_2205,N_2265);
or U2432 (N_2432,N_2244,N_2347);
or U2433 (N_2433,N_2359,N_2246);
nor U2434 (N_2434,N_2324,N_2294);
nand U2435 (N_2435,N_2241,N_2282);
and U2436 (N_2436,N_2343,N_2330);
nand U2437 (N_2437,N_2228,N_2213);
nand U2438 (N_2438,N_2350,N_2387);
nor U2439 (N_2439,N_2338,N_2370);
and U2440 (N_2440,N_2331,N_2314);
nand U2441 (N_2441,N_2362,N_2258);
nand U2442 (N_2442,N_2299,N_2295);
nand U2443 (N_2443,N_2271,N_2304);
nor U2444 (N_2444,N_2238,N_2272);
nor U2445 (N_2445,N_2379,N_2217);
nor U2446 (N_2446,N_2321,N_2207);
nor U2447 (N_2447,N_2256,N_2342);
and U2448 (N_2448,N_2226,N_2312);
or U2449 (N_2449,N_2227,N_2369);
and U2450 (N_2450,N_2280,N_2253);
nor U2451 (N_2451,N_2323,N_2309);
nand U2452 (N_2452,N_2373,N_2353);
nor U2453 (N_2453,N_2395,N_2326);
nand U2454 (N_2454,N_2303,N_2388);
or U2455 (N_2455,N_2381,N_2204);
or U2456 (N_2456,N_2219,N_2231);
and U2457 (N_2457,N_2335,N_2322);
nand U2458 (N_2458,N_2220,N_2357);
and U2459 (N_2459,N_2248,N_2383);
or U2460 (N_2460,N_2264,N_2267);
nand U2461 (N_2461,N_2348,N_2346);
nand U2462 (N_2462,N_2345,N_2293);
nor U2463 (N_2463,N_2372,N_2239);
nand U2464 (N_2464,N_2263,N_2266);
or U2465 (N_2465,N_2212,N_2361);
nor U2466 (N_2466,N_2276,N_2384);
nand U2467 (N_2467,N_2277,N_2218);
or U2468 (N_2468,N_2281,N_2394);
or U2469 (N_2469,N_2355,N_2274);
nor U2470 (N_2470,N_2328,N_2349);
and U2471 (N_2471,N_2230,N_2243);
nor U2472 (N_2472,N_2229,N_2363);
nor U2473 (N_2473,N_2327,N_2380);
and U2474 (N_2474,N_2318,N_2344);
or U2475 (N_2475,N_2371,N_2337);
or U2476 (N_2476,N_2382,N_2296);
and U2477 (N_2477,N_2200,N_2375);
nor U2478 (N_2478,N_2251,N_2215);
nor U2479 (N_2479,N_2358,N_2305);
or U2480 (N_2480,N_2307,N_2275);
nor U2481 (N_2481,N_2262,N_2214);
nand U2482 (N_2482,N_2259,N_2368);
and U2483 (N_2483,N_2250,N_2221);
nand U2484 (N_2484,N_2319,N_2341);
and U2485 (N_2485,N_2366,N_2374);
nor U2486 (N_2486,N_2249,N_2351);
or U2487 (N_2487,N_2367,N_2377);
and U2488 (N_2488,N_2292,N_2308);
and U2489 (N_2489,N_2386,N_2302);
nand U2490 (N_2490,N_2240,N_2306);
nor U2491 (N_2491,N_2232,N_2222);
or U2492 (N_2492,N_2285,N_2252);
or U2493 (N_2493,N_2396,N_2283);
nor U2494 (N_2494,N_2397,N_2247);
nor U2495 (N_2495,N_2269,N_2352);
or U2496 (N_2496,N_2286,N_2216);
or U2497 (N_2497,N_2385,N_2208);
and U2498 (N_2498,N_2392,N_2365);
and U2499 (N_2499,N_2393,N_2391);
or U2500 (N_2500,N_2314,N_2380);
or U2501 (N_2501,N_2379,N_2251);
or U2502 (N_2502,N_2357,N_2386);
and U2503 (N_2503,N_2262,N_2282);
nor U2504 (N_2504,N_2310,N_2241);
nand U2505 (N_2505,N_2305,N_2288);
nor U2506 (N_2506,N_2232,N_2310);
nand U2507 (N_2507,N_2388,N_2255);
and U2508 (N_2508,N_2352,N_2297);
nand U2509 (N_2509,N_2226,N_2377);
and U2510 (N_2510,N_2240,N_2348);
nand U2511 (N_2511,N_2219,N_2248);
nand U2512 (N_2512,N_2234,N_2337);
or U2513 (N_2513,N_2261,N_2371);
or U2514 (N_2514,N_2303,N_2301);
nand U2515 (N_2515,N_2269,N_2396);
or U2516 (N_2516,N_2361,N_2275);
nor U2517 (N_2517,N_2303,N_2386);
nor U2518 (N_2518,N_2326,N_2365);
nor U2519 (N_2519,N_2235,N_2343);
nand U2520 (N_2520,N_2321,N_2291);
nor U2521 (N_2521,N_2209,N_2313);
nor U2522 (N_2522,N_2328,N_2264);
or U2523 (N_2523,N_2345,N_2367);
and U2524 (N_2524,N_2235,N_2240);
or U2525 (N_2525,N_2332,N_2203);
nor U2526 (N_2526,N_2399,N_2215);
nor U2527 (N_2527,N_2367,N_2216);
and U2528 (N_2528,N_2294,N_2386);
and U2529 (N_2529,N_2203,N_2231);
nand U2530 (N_2530,N_2270,N_2399);
and U2531 (N_2531,N_2260,N_2330);
or U2532 (N_2532,N_2375,N_2250);
and U2533 (N_2533,N_2361,N_2297);
nand U2534 (N_2534,N_2280,N_2250);
or U2535 (N_2535,N_2294,N_2224);
and U2536 (N_2536,N_2266,N_2206);
or U2537 (N_2537,N_2390,N_2248);
nand U2538 (N_2538,N_2222,N_2297);
nand U2539 (N_2539,N_2273,N_2290);
and U2540 (N_2540,N_2304,N_2317);
nor U2541 (N_2541,N_2242,N_2372);
nand U2542 (N_2542,N_2290,N_2216);
or U2543 (N_2543,N_2243,N_2200);
and U2544 (N_2544,N_2262,N_2244);
nor U2545 (N_2545,N_2295,N_2240);
nor U2546 (N_2546,N_2228,N_2274);
and U2547 (N_2547,N_2379,N_2235);
or U2548 (N_2548,N_2289,N_2250);
and U2549 (N_2549,N_2239,N_2352);
or U2550 (N_2550,N_2385,N_2324);
and U2551 (N_2551,N_2233,N_2353);
nor U2552 (N_2552,N_2355,N_2324);
xnor U2553 (N_2553,N_2282,N_2320);
or U2554 (N_2554,N_2247,N_2250);
and U2555 (N_2555,N_2300,N_2380);
nand U2556 (N_2556,N_2293,N_2359);
nand U2557 (N_2557,N_2387,N_2268);
nand U2558 (N_2558,N_2280,N_2240);
xor U2559 (N_2559,N_2325,N_2263);
nand U2560 (N_2560,N_2349,N_2304);
and U2561 (N_2561,N_2394,N_2239);
nor U2562 (N_2562,N_2227,N_2375);
and U2563 (N_2563,N_2367,N_2217);
or U2564 (N_2564,N_2233,N_2305);
nor U2565 (N_2565,N_2293,N_2367);
nand U2566 (N_2566,N_2202,N_2329);
and U2567 (N_2567,N_2348,N_2217);
nor U2568 (N_2568,N_2348,N_2393);
nand U2569 (N_2569,N_2258,N_2326);
and U2570 (N_2570,N_2317,N_2230);
nor U2571 (N_2571,N_2287,N_2331);
and U2572 (N_2572,N_2396,N_2321);
nor U2573 (N_2573,N_2335,N_2273);
and U2574 (N_2574,N_2367,N_2374);
nand U2575 (N_2575,N_2276,N_2235);
and U2576 (N_2576,N_2306,N_2264);
nand U2577 (N_2577,N_2255,N_2326);
and U2578 (N_2578,N_2233,N_2289);
or U2579 (N_2579,N_2229,N_2318);
nand U2580 (N_2580,N_2384,N_2325);
nand U2581 (N_2581,N_2349,N_2379);
or U2582 (N_2582,N_2364,N_2345);
nand U2583 (N_2583,N_2326,N_2376);
xor U2584 (N_2584,N_2386,N_2201);
nor U2585 (N_2585,N_2369,N_2268);
or U2586 (N_2586,N_2365,N_2371);
or U2587 (N_2587,N_2251,N_2378);
and U2588 (N_2588,N_2378,N_2229);
and U2589 (N_2589,N_2345,N_2224);
and U2590 (N_2590,N_2272,N_2294);
and U2591 (N_2591,N_2372,N_2315);
or U2592 (N_2592,N_2361,N_2203);
nor U2593 (N_2593,N_2292,N_2338);
or U2594 (N_2594,N_2241,N_2398);
nand U2595 (N_2595,N_2214,N_2306);
nand U2596 (N_2596,N_2237,N_2334);
or U2597 (N_2597,N_2209,N_2274);
nand U2598 (N_2598,N_2318,N_2350);
xor U2599 (N_2599,N_2322,N_2332);
nand U2600 (N_2600,N_2432,N_2420);
and U2601 (N_2601,N_2440,N_2522);
nand U2602 (N_2602,N_2494,N_2410);
and U2603 (N_2603,N_2530,N_2442);
or U2604 (N_2604,N_2457,N_2458);
or U2605 (N_2605,N_2470,N_2571);
or U2606 (N_2606,N_2417,N_2456);
nand U2607 (N_2607,N_2445,N_2452);
nand U2608 (N_2608,N_2472,N_2558);
and U2609 (N_2609,N_2537,N_2562);
nor U2610 (N_2610,N_2513,N_2489);
nand U2611 (N_2611,N_2597,N_2565);
and U2612 (N_2612,N_2401,N_2435);
nor U2613 (N_2613,N_2583,N_2408);
and U2614 (N_2614,N_2478,N_2575);
and U2615 (N_2615,N_2477,N_2591);
nand U2616 (N_2616,N_2403,N_2517);
or U2617 (N_2617,N_2579,N_2539);
or U2618 (N_2618,N_2501,N_2423);
nand U2619 (N_2619,N_2535,N_2505);
or U2620 (N_2620,N_2511,N_2464);
or U2621 (N_2621,N_2459,N_2553);
and U2622 (N_2622,N_2506,N_2484);
or U2623 (N_2623,N_2434,N_2424);
nand U2624 (N_2624,N_2599,N_2534);
nor U2625 (N_2625,N_2454,N_2520);
and U2626 (N_2626,N_2497,N_2431);
nor U2627 (N_2627,N_2402,N_2418);
and U2628 (N_2628,N_2487,N_2468);
nand U2629 (N_2629,N_2427,N_2588);
nand U2630 (N_2630,N_2594,N_2563);
or U2631 (N_2631,N_2578,N_2473);
or U2632 (N_2632,N_2481,N_2550);
or U2633 (N_2633,N_2476,N_2480);
or U2634 (N_2634,N_2462,N_2572);
or U2635 (N_2635,N_2504,N_2507);
or U2636 (N_2636,N_2465,N_2586);
or U2637 (N_2637,N_2540,N_2439);
nand U2638 (N_2638,N_2584,N_2433);
nand U2639 (N_2639,N_2425,N_2449);
nor U2640 (N_2640,N_2598,N_2536);
or U2641 (N_2641,N_2544,N_2546);
nor U2642 (N_2642,N_2528,N_2595);
nor U2643 (N_2643,N_2547,N_2491);
nand U2644 (N_2644,N_2526,N_2587);
nor U2645 (N_2645,N_2589,N_2561);
and U2646 (N_2646,N_2446,N_2461);
nand U2647 (N_2647,N_2585,N_2512);
or U2648 (N_2648,N_2523,N_2525);
nor U2649 (N_2649,N_2437,N_2519);
nand U2650 (N_2650,N_2500,N_2593);
nand U2651 (N_2651,N_2436,N_2463);
or U2652 (N_2652,N_2411,N_2490);
and U2653 (N_2653,N_2404,N_2430);
nor U2654 (N_2654,N_2551,N_2426);
nor U2655 (N_2655,N_2407,N_2475);
nor U2656 (N_2656,N_2444,N_2568);
or U2657 (N_2657,N_2429,N_2533);
nor U2658 (N_2658,N_2543,N_2479);
nand U2659 (N_2659,N_2566,N_2560);
and U2660 (N_2660,N_2567,N_2559);
xor U2661 (N_2661,N_2556,N_2474);
and U2662 (N_2662,N_2557,N_2453);
nor U2663 (N_2663,N_2531,N_2412);
nand U2664 (N_2664,N_2460,N_2516);
and U2665 (N_2665,N_2485,N_2569);
nor U2666 (N_2666,N_2448,N_2555);
or U2667 (N_2667,N_2492,N_2469);
and U2668 (N_2668,N_2451,N_2545);
and U2669 (N_2669,N_2428,N_2502);
nand U2670 (N_2670,N_2483,N_2421);
and U2671 (N_2671,N_2413,N_2405);
and U2672 (N_2672,N_2518,N_2510);
nand U2673 (N_2673,N_2438,N_2542);
or U2674 (N_2674,N_2582,N_2592);
or U2675 (N_2675,N_2416,N_2419);
or U2676 (N_2676,N_2554,N_2496);
nor U2677 (N_2677,N_2415,N_2581);
nor U2678 (N_2678,N_2580,N_2552);
and U2679 (N_2679,N_2482,N_2422);
nor U2680 (N_2680,N_2574,N_2495);
nand U2681 (N_2681,N_2409,N_2400);
nand U2682 (N_2682,N_2548,N_2503);
and U2683 (N_2683,N_2406,N_2576);
nand U2684 (N_2684,N_2467,N_2466);
nand U2685 (N_2685,N_2590,N_2527);
nand U2686 (N_2686,N_2443,N_2486);
and U2687 (N_2687,N_2499,N_2532);
nand U2688 (N_2688,N_2521,N_2509);
nand U2689 (N_2689,N_2515,N_2529);
nand U2690 (N_2690,N_2447,N_2471);
or U2691 (N_2691,N_2524,N_2596);
nor U2692 (N_2692,N_2549,N_2441);
nand U2693 (N_2693,N_2508,N_2573);
and U2694 (N_2694,N_2493,N_2455);
nor U2695 (N_2695,N_2488,N_2450);
and U2696 (N_2696,N_2538,N_2570);
nand U2697 (N_2697,N_2564,N_2414);
nor U2698 (N_2698,N_2498,N_2577);
and U2699 (N_2699,N_2514,N_2541);
or U2700 (N_2700,N_2568,N_2413);
nor U2701 (N_2701,N_2423,N_2529);
nand U2702 (N_2702,N_2590,N_2499);
nor U2703 (N_2703,N_2577,N_2568);
and U2704 (N_2704,N_2577,N_2472);
nor U2705 (N_2705,N_2506,N_2595);
or U2706 (N_2706,N_2598,N_2511);
nand U2707 (N_2707,N_2543,N_2431);
or U2708 (N_2708,N_2525,N_2401);
and U2709 (N_2709,N_2449,N_2427);
and U2710 (N_2710,N_2445,N_2597);
or U2711 (N_2711,N_2462,N_2511);
nor U2712 (N_2712,N_2500,N_2451);
or U2713 (N_2713,N_2492,N_2599);
nand U2714 (N_2714,N_2583,N_2503);
and U2715 (N_2715,N_2590,N_2569);
or U2716 (N_2716,N_2426,N_2465);
and U2717 (N_2717,N_2421,N_2547);
or U2718 (N_2718,N_2572,N_2471);
nor U2719 (N_2719,N_2427,N_2430);
or U2720 (N_2720,N_2584,N_2557);
xor U2721 (N_2721,N_2576,N_2506);
and U2722 (N_2722,N_2590,N_2498);
nand U2723 (N_2723,N_2591,N_2500);
nand U2724 (N_2724,N_2540,N_2512);
nand U2725 (N_2725,N_2476,N_2419);
or U2726 (N_2726,N_2516,N_2432);
and U2727 (N_2727,N_2543,N_2423);
nand U2728 (N_2728,N_2566,N_2417);
nor U2729 (N_2729,N_2509,N_2425);
nand U2730 (N_2730,N_2445,N_2575);
nand U2731 (N_2731,N_2400,N_2550);
or U2732 (N_2732,N_2457,N_2440);
nand U2733 (N_2733,N_2586,N_2562);
or U2734 (N_2734,N_2499,N_2564);
nand U2735 (N_2735,N_2596,N_2402);
and U2736 (N_2736,N_2564,N_2548);
nor U2737 (N_2737,N_2488,N_2550);
and U2738 (N_2738,N_2490,N_2473);
nand U2739 (N_2739,N_2481,N_2588);
or U2740 (N_2740,N_2540,N_2497);
or U2741 (N_2741,N_2456,N_2427);
nand U2742 (N_2742,N_2522,N_2408);
xnor U2743 (N_2743,N_2474,N_2440);
xnor U2744 (N_2744,N_2504,N_2581);
and U2745 (N_2745,N_2488,N_2435);
nand U2746 (N_2746,N_2458,N_2472);
and U2747 (N_2747,N_2534,N_2523);
nor U2748 (N_2748,N_2587,N_2593);
nand U2749 (N_2749,N_2454,N_2551);
nor U2750 (N_2750,N_2554,N_2413);
nand U2751 (N_2751,N_2405,N_2526);
xnor U2752 (N_2752,N_2481,N_2506);
nand U2753 (N_2753,N_2486,N_2552);
and U2754 (N_2754,N_2474,N_2579);
nand U2755 (N_2755,N_2553,N_2455);
and U2756 (N_2756,N_2439,N_2464);
nor U2757 (N_2757,N_2554,N_2432);
and U2758 (N_2758,N_2435,N_2501);
nand U2759 (N_2759,N_2544,N_2592);
or U2760 (N_2760,N_2519,N_2411);
nand U2761 (N_2761,N_2599,N_2474);
nand U2762 (N_2762,N_2582,N_2415);
nand U2763 (N_2763,N_2444,N_2563);
or U2764 (N_2764,N_2405,N_2448);
nor U2765 (N_2765,N_2572,N_2476);
and U2766 (N_2766,N_2460,N_2429);
or U2767 (N_2767,N_2483,N_2580);
or U2768 (N_2768,N_2413,N_2548);
or U2769 (N_2769,N_2597,N_2411);
or U2770 (N_2770,N_2588,N_2465);
nand U2771 (N_2771,N_2544,N_2448);
nand U2772 (N_2772,N_2486,N_2475);
nor U2773 (N_2773,N_2506,N_2415);
and U2774 (N_2774,N_2514,N_2451);
and U2775 (N_2775,N_2456,N_2558);
nand U2776 (N_2776,N_2462,N_2546);
nand U2777 (N_2777,N_2505,N_2478);
nand U2778 (N_2778,N_2458,N_2431);
nand U2779 (N_2779,N_2432,N_2581);
and U2780 (N_2780,N_2451,N_2524);
or U2781 (N_2781,N_2451,N_2582);
nand U2782 (N_2782,N_2556,N_2558);
nand U2783 (N_2783,N_2568,N_2557);
and U2784 (N_2784,N_2467,N_2415);
and U2785 (N_2785,N_2541,N_2533);
nor U2786 (N_2786,N_2479,N_2464);
or U2787 (N_2787,N_2574,N_2510);
and U2788 (N_2788,N_2526,N_2403);
nor U2789 (N_2789,N_2479,N_2547);
nor U2790 (N_2790,N_2543,N_2485);
nor U2791 (N_2791,N_2448,N_2499);
or U2792 (N_2792,N_2409,N_2554);
and U2793 (N_2793,N_2454,N_2585);
and U2794 (N_2794,N_2585,N_2559);
nor U2795 (N_2795,N_2570,N_2597);
nand U2796 (N_2796,N_2419,N_2406);
or U2797 (N_2797,N_2437,N_2595);
nor U2798 (N_2798,N_2414,N_2589);
nand U2799 (N_2799,N_2535,N_2508);
nand U2800 (N_2800,N_2651,N_2614);
nor U2801 (N_2801,N_2666,N_2671);
nand U2802 (N_2802,N_2660,N_2628);
or U2803 (N_2803,N_2616,N_2692);
and U2804 (N_2804,N_2745,N_2639);
and U2805 (N_2805,N_2749,N_2683);
nand U2806 (N_2806,N_2687,N_2633);
nand U2807 (N_2807,N_2640,N_2731);
nor U2808 (N_2808,N_2714,N_2681);
or U2809 (N_2809,N_2631,N_2600);
or U2810 (N_2810,N_2622,N_2663);
nor U2811 (N_2811,N_2762,N_2799);
or U2812 (N_2812,N_2779,N_2647);
nand U2813 (N_2813,N_2739,N_2643);
nor U2814 (N_2814,N_2775,N_2763);
and U2815 (N_2815,N_2790,N_2690);
or U2816 (N_2816,N_2684,N_2727);
and U2817 (N_2817,N_2755,N_2612);
or U2818 (N_2818,N_2703,N_2746);
and U2819 (N_2819,N_2637,N_2758);
or U2820 (N_2820,N_2736,N_2735);
and U2821 (N_2821,N_2734,N_2604);
or U2822 (N_2822,N_2765,N_2636);
and U2823 (N_2823,N_2642,N_2773);
or U2824 (N_2824,N_2757,N_2621);
nand U2825 (N_2825,N_2783,N_2764);
nand U2826 (N_2826,N_2786,N_2602);
and U2827 (N_2827,N_2717,N_2635);
nand U2828 (N_2828,N_2619,N_2759);
and U2829 (N_2829,N_2748,N_2705);
nor U2830 (N_2830,N_2613,N_2654);
nor U2831 (N_2831,N_2719,N_2625);
or U2832 (N_2832,N_2794,N_2627);
nor U2833 (N_2833,N_2784,N_2725);
xnor U2834 (N_2834,N_2675,N_2653);
nand U2835 (N_2835,N_2618,N_2667);
nand U2836 (N_2836,N_2655,N_2712);
or U2837 (N_2837,N_2788,N_2668);
and U2838 (N_2838,N_2610,N_2742);
or U2839 (N_2839,N_2697,N_2669);
or U2840 (N_2840,N_2724,N_2650);
nor U2841 (N_2841,N_2718,N_2673);
and U2842 (N_2842,N_2608,N_2658);
and U2843 (N_2843,N_2728,N_2760);
and U2844 (N_2844,N_2617,N_2713);
nand U2845 (N_2845,N_2709,N_2743);
or U2846 (N_2846,N_2656,N_2756);
nand U2847 (N_2847,N_2787,N_2630);
or U2848 (N_2848,N_2751,N_2664);
and U2849 (N_2849,N_2708,N_2737);
and U2850 (N_2850,N_2605,N_2792);
xor U2851 (N_2851,N_2721,N_2691);
or U2852 (N_2852,N_2624,N_2798);
nor U2853 (N_2853,N_2670,N_2665);
and U2854 (N_2854,N_2766,N_2676);
nand U2855 (N_2855,N_2609,N_2699);
nor U2856 (N_2856,N_2701,N_2620);
and U2857 (N_2857,N_2603,N_2682);
nand U2858 (N_2858,N_2770,N_2780);
nor U2859 (N_2859,N_2679,N_2644);
nor U2860 (N_2860,N_2776,N_2767);
nor U2861 (N_2861,N_2626,N_2791);
nor U2862 (N_2862,N_2674,N_2629);
nor U2863 (N_2863,N_2657,N_2795);
or U2864 (N_2864,N_2648,N_2781);
nor U2865 (N_2865,N_2772,N_2611);
nor U2866 (N_2866,N_2672,N_2778);
nand U2867 (N_2867,N_2649,N_2710);
or U2868 (N_2868,N_2771,N_2738);
or U2869 (N_2869,N_2706,N_2615);
or U2870 (N_2870,N_2607,N_2659);
or U2871 (N_2871,N_2774,N_2686);
nor U2872 (N_2872,N_2696,N_2740);
and U2873 (N_2873,N_2761,N_2646);
and U2874 (N_2874,N_2711,N_2730);
or U2875 (N_2875,N_2685,N_2747);
and U2876 (N_2876,N_2688,N_2716);
or U2877 (N_2877,N_2634,N_2732);
or U2878 (N_2878,N_2606,N_2645);
nor U2879 (N_2879,N_2652,N_2693);
and U2880 (N_2880,N_2785,N_2641);
nor U2881 (N_2881,N_2750,N_2733);
nor U2882 (N_2882,N_2704,N_2797);
nor U2883 (N_2883,N_2777,N_2698);
and U2884 (N_2884,N_2715,N_2769);
or U2885 (N_2885,N_2789,N_2723);
nand U2886 (N_2886,N_2678,N_2768);
nor U2887 (N_2887,N_2741,N_2695);
nand U2888 (N_2888,N_2689,N_2753);
and U2889 (N_2889,N_2754,N_2782);
nand U2890 (N_2890,N_2601,N_2694);
or U2891 (N_2891,N_2662,N_2623);
or U2892 (N_2892,N_2752,N_2632);
or U2893 (N_2893,N_2700,N_2726);
nor U2894 (N_2894,N_2677,N_2638);
and U2895 (N_2895,N_2722,N_2729);
nand U2896 (N_2896,N_2720,N_2707);
or U2897 (N_2897,N_2793,N_2796);
nor U2898 (N_2898,N_2680,N_2744);
or U2899 (N_2899,N_2702,N_2661);
nor U2900 (N_2900,N_2684,N_2674);
nor U2901 (N_2901,N_2773,N_2617);
nand U2902 (N_2902,N_2797,N_2701);
or U2903 (N_2903,N_2670,N_2702);
and U2904 (N_2904,N_2796,N_2744);
and U2905 (N_2905,N_2662,N_2766);
nor U2906 (N_2906,N_2786,N_2788);
and U2907 (N_2907,N_2698,N_2651);
and U2908 (N_2908,N_2636,N_2752);
nand U2909 (N_2909,N_2661,N_2743);
and U2910 (N_2910,N_2719,N_2668);
or U2911 (N_2911,N_2742,N_2646);
nor U2912 (N_2912,N_2729,N_2747);
nor U2913 (N_2913,N_2797,N_2739);
nand U2914 (N_2914,N_2619,N_2781);
nor U2915 (N_2915,N_2783,N_2762);
nor U2916 (N_2916,N_2617,N_2677);
or U2917 (N_2917,N_2633,N_2634);
and U2918 (N_2918,N_2763,N_2691);
or U2919 (N_2919,N_2644,N_2776);
or U2920 (N_2920,N_2675,N_2609);
and U2921 (N_2921,N_2741,N_2677);
nand U2922 (N_2922,N_2789,N_2708);
or U2923 (N_2923,N_2719,N_2616);
nand U2924 (N_2924,N_2659,N_2620);
nand U2925 (N_2925,N_2783,N_2627);
nor U2926 (N_2926,N_2722,N_2742);
nor U2927 (N_2927,N_2657,N_2635);
nand U2928 (N_2928,N_2638,N_2695);
nor U2929 (N_2929,N_2744,N_2740);
or U2930 (N_2930,N_2796,N_2708);
and U2931 (N_2931,N_2624,N_2710);
nand U2932 (N_2932,N_2653,N_2686);
nor U2933 (N_2933,N_2658,N_2717);
or U2934 (N_2934,N_2794,N_2608);
or U2935 (N_2935,N_2653,N_2641);
nand U2936 (N_2936,N_2678,N_2774);
and U2937 (N_2937,N_2768,N_2754);
nand U2938 (N_2938,N_2621,N_2642);
or U2939 (N_2939,N_2680,N_2767);
and U2940 (N_2940,N_2716,N_2659);
nor U2941 (N_2941,N_2642,N_2672);
or U2942 (N_2942,N_2673,N_2638);
or U2943 (N_2943,N_2742,N_2618);
nand U2944 (N_2944,N_2629,N_2707);
nand U2945 (N_2945,N_2620,N_2682);
or U2946 (N_2946,N_2679,N_2799);
and U2947 (N_2947,N_2652,N_2788);
nand U2948 (N_2948,N_2764,N_2695);
nand U2949 (N_2949,N_2693,N_2658);
or U2950 (N_2950,N_2713,N_2740);
and U2951 (N_2951,N_2636,N_2697);
and U2952 (N_2952,N_2706,N_2601);
and U2953 (N_2953,N_2600,N_2602);
nand U2954 (N_2954,N_2665,N_2664);
nor U2955 (N_2955,N_2721,N_2777);
or U2956 (N_2956,N_2623,N_2726);
or U2957 (N_2957,N_2760,N_2791);
or U2958 (N_2958,N_2622,N_2614);
and U2959 (N_2959,N_2688,N_2643);
nand U2960 (N_2960,N_2760,N_2701);
or U2961 (N_2961,N_2630,N_2673);
nand U2962 (N_2962,N_2666,N_2673);
or U2963 (N_2963,N_2698,N_2778);
and U2964 (N_2964,N_2741,N_2681);
nor U2965 (N_2965,N_2666,N_2770);
or U2966 (N_2966,N_2704,N_2764);
nor U2967 (N_2967,N_2789,N_2755);
nand U2968 (N_2968,N_2630,N_2749);
nand U2969 (N_2969,N_2723,N_2629);
and U2970 (N_2970,N_2721,N_2768);
nand U2971 (N_2971,N_2780,N_2754);
nand U2972 (N_2972,N_2717,N_2604);
or U2973 (N_2973,N_2687,N_2786);
nand U2974 (N_2974,N_2729,N_2659);
or U2975 (N_2975,N_2797,N_2628);
nand U2976 (N_2976,N_2748,N_2678);
nand U2977 (N_2977,N_2656,N_2655);
and U2978 (N_2978,N_2777,N_2626);
nand U2979 (N_2979,N_2726,N_2769);
nor U2980 (N_2980,N_2687,N_2793);
nand U2981 (N_2981,N_2779,N_2716);
nor U2982 (N_2982,N_2738,N_2661);
nor U2983 (N_2983,N_2691,N_2689);
and U2984 (N_2984,N_2761,N_2754);
and U2985 (N_2985,N_2784,N_2625);
and U2986 (N_2986,N_2644,N_2625);
or U2987 (N_2987,N_2757,N_2744);
and U2988 (N_2988,N_2634,N_2741);
nor U2989 (N_2989,N_2652,N_2714);
nand U2990 (N_2990,N_2690,N_2651);
and U2991 (N_2991,N_2608,N_2719);
nand U2992 (N_2992,N_2614,N_2749);
nor U2993 (N_2993,N_2672,N_2752);
nand U2994 (N_2994,N_2617,N_2765);
nor U2995 (N_2995,N_2694,N_2665);
nor U2996 (N_2996,N_2638,N_2620);
or U2997 (N_2997,N_2799,N_2797);
and U2998 (N_2998,N_2795,N_2677);
nand U2999 (N_2999,N_2795,N_2649);
or UO_0 (O_0,N_2997,N_2942);
nor UO_1 (O_1,N_2821,N_2914);
nand UO_2 (O_2,N_2874,N_2905);
or UO_3 (O_3,N_2812,N_2846);
or UO_4 (O_4,N_2946,N_2885);
and UO_5 (O_5,N_2969,N_2860);
or UO_6 (O_6,N_2919,N_2987);
and UO_7 (O_7,N_2840,N_2981);
or UO_8 (O_8,N_2916,N_2810);
nor UO_9 (O_9,N_2959,N_2937);
nor UO_10 (O_10,N_2983,N_2901);
nor UO_11 (O_11,N_2972,N_2865);
nand UO_12 (O_12,N_2825,N_2859);
and UO_13 (O_13,N_2961,N_2973);
or UO_14 (O_14,N_2968,N_2828);
nand UO_15 (O_15,N_2802,N_2814);
or UO_16 (O_16,N_2945,N_2858);
nor UO_17 (O_17,N_2925,N_2890);
or UO_18 (O_18,N_2984,N_2941);
or UO_19 (O_19,N_2808,N_2831);
or UO_20 (O_20,N_2949,N_2966);
or UO_21 (O_21,N_2801,N_2803);
nand UO_22 (O_22,N_2882,N_2926);
or UO_23 (O_23,N_2857,N_2913);
or UO_24 (O_24,N_2958,N_2823);
and UO_25 (O_25,N_2832,N_2988);
or UO_26 (O_26,N_2982,N_2998);
and UO_27 (O_27,N_2985,N_2893);
nand UO_28 (O_28,N_2939,N_2889);
or UO_29 (O_29,N_2922,N_2903);
and UO_30 (O_30,N_2943,N_2904);
nor UO_31 (O_31,N_2956,N_2954);
and UO_32 (O_32,N_2870,N_2979);
nand UO_33 (O_33,N_2848,N_2886);
nand UO_34 (O_34,N_2978,N_2871);
nand UO_35 (O_35,N_2842,N_2824);
nor UO_36 (O_36,N_2932,N_2990);
nand UO_37 (O_37,N_2887,N_2809);
or UO_38 (O_38,N_2816,N_2999);
and UO_39 (O_39,N_2837,N_2918);
nand UO_40 (O_40,N_2834,N_2955);
nand UO_41 (O_41,N_2891,N_2856);
nor UO_42 (O_42,N_2888,N_2829);
or UO_43 (O_43,N_2854,N_2881);
and UO_44 (O_44,N_2951,N_2872);
or UO_45 (O_45,N_2957,N_2867);
and UO_46 (O_46,N_2950,N_2953);
nor UO_47 (O_47,N_2895,N_2996);
or UO_48 (O_48,N_2965,N_2868);
nand UO_49 (O_49,N_2838,N_2944);
nor UO_50 (O_50,N_2976,N_2819);
nor UO_51 (O_51,N_2804,N_2928);
nor UO_52 (O_52,N_2836,N_2866);
nand UO_53 (O_53,N_2835,N_2947);
and UO_54 (O_54,N_2806,N_2898);
nand UO_55 (O_55,N_2911,N_2934);
or UO_56 (O_56,N_2995,N_2864);
nor UO_57 (O_57,N_2967,N_2818);
nand UO_58 (O_58,N_2894,N_2879);
nand UO_59 (O_59,N_2853,N_2845);
and UO_60 (O_60,N_2813,N_2991);
or UO_61 (O_61,N_2923,N_2974);
or UO_62 (O_62,N_2964,N_2920);
nand UO_63 (O_63,N_2921,N_2929);
nor UO_64 (O_64,N_2855,N_2847);
nor UO_65 (O_65,N_2940,N_2852);
and UO_66 (O_66,N_2899,N_2910);
or UO_67 (O_67,N_2862,N_2849);
and UO_68 (O_68,N_2875,N_2839);
nor UO_69 (O_69,N_2936,N_2843);
and UO_70 (O_70,N_2924,N_2822);
nor UO_71 (O_71,N_2850,N_2909);
nor UO_72 (O_72,N_2927,N_2908);
nor UO_73 (O_73,N_2963,N_2915);
and UO_74 (O_74,N_2977,N_2931);
or UO_75 (O_75,N_2933,N_2897);
nand UO_76 (O_76,N_2960,N_2878);
nor UO_77 (O_77,N_2962,N_2877);
or UO_78 (O_78,N_2851,N_2906);
nand UO_79 (O_79,N_2883,N_2986);
and UO_80 (O_80,N_2869,N_2952);
nor UO_81 (O_81,N_2830,N_2930);
and UO_82 (O_82,N_2815,N_2861);
and UO_83 (O_83,N_2807,N_2892);
nand UO_84 (O_84,N_2989,N_2917);
or UO_85 (O_85,N_2884,N_2863);
or UO_86 (O_86,N_2900,N_2975);
and UO_87 (O_87,N_2844,N_2820);
nor UO_88 (O_88,N_2907,N_2902);
or UO_89 (O_89,N_2896,N_2876);
and UO_90 (O_90,N_2971,N_2827);
nand UO_91 (O_91,N_2994,N_2970);
or UO_92 (O_92,N_2811,N_2880);
and UO_93 (O_93,N_2841,N_2993);
nand UO_94 (O_94,N_2826,N_2948);
and UO_95 (O_95,N_2935,N_2912);
or UO_96 (O_96,N_2938,N_2980);
or UO_97 (O_97,N_2833,N_2873);
and UO_98 (O_98,N_2800,N_2817);
or UO_99 (O_99,N_2992,N_2805);
nor UO_100 (O_100,N_2847,N_2808);
nor UO_101 (O_101,N_2869,N_2989);
or UO_102 (O_102,N_2897,N_2834);
and UO_103 (O_103,N_2935,N_2886);
nand UO_104 (O_104,N_2963,N_2877);
and UO_105 (O_105,N_2848,N_2913);
nand UO_106 (O_106,N_2852,N_2892);
or UO_107 (O_107,N_2861,N_2961);
nand UO_108 (O_108,N_2910,N_2813);
nand UO_109 (O_109,N_2834,N_2863);
and UO_110 (O_110,N_2840,N_2985);
or UO_111 (O_111,N_2961,N_2980);
and UO_112 (O_112,N_2883,N_2810);
nor UO_113 (O_113,N_2870,N_2844);
nor UO_114 (O_114,N_2883,N_2837);
nand UO_115 (O_115,N_2805,N_2918);
and UO_116 (O_116,N_2830,N_2919);
nor UO_117 (O_117,N_2929,N_2925);
and UO_118 (O_118,N_2868,N_2840);
nand UO_119 (O_119,N_2819,N_2975);
nand UO_120 (O_120,N_2854,N_2837);
or UO_121 (O_121,N_2892,N_2808);
or UO_122 (O_122,N_2914,N_2933);
nor UO_123 (O_123,N_2851,N_2970);
nand UO_124 (O_124,N_2830,N_2860);
nand UO_125 (O_125,N_2848,N_2888);
nor UO_126 (O_126,N_2897,N_2883);
nand UO_127 (O_127,N_2936,N_2829);
nor UO_128 (O_128,N_2903,N_2964);
nand UO_129 (O_129,N_2856,N_2990);
or UO_130 (O_130,N_2903,N_2870);
nand UO_131 (O_131,N_2971,N_2891);
and UO_132 (O_132,N_2930,N_2858);
and UO_133 (O_133,N_2926,N_2902);
nor UO_134 (O_134,N_2866,N_2829);
nand UO_135 (O_135,N_2922,N_2803);
nand UO_136 (O_136,N_2853,N_2810);
nand UO_137 (O_137,N_2973,N_2915);
and UO_138 (O_138,N_2965,N_2860);
nand UO_139 (O_139,N_2963,N_2826);
nand UO_140 (O_140,N_2895,N_2949);
and UO_141 (O_141,N_2835,N_2940);
or UO_142 (O_142,N_2828,N_2889);
or UO_143 (O_143,N_2939,N_2811);
nand UO_144 (O_144,N_2812,N_2972);
or UO_145 (O_145,N_2939,N_2873);
and UO_146 (O_146,N_2866,N_2805);
and UO_147 (O_147,N_2903,N_2800);
nand UO_148 (O_148,N_2967,N_2868);
nor UO_149 (O_149,N_2823,N_2832);
or UO_150 (O_150,N_2901,N_2924);
or UO_151 (O_151,N_2814,N_2951);
or UO_152 (O_152,N_2908,N_2961);
or UO_153 (O_153,N_2993,N_2831);
and UO_154 (O_154,N_2906,N_2855);
nand UO_155 (O_155,N_2978,N_2926);
nand UO_156 (O_156,N_2815,N_2873);
nand UO_157 (O_157,N_2887,N_2906);
nand UO_158 (O_158,N_2903,N_2876);
nand UO_159 (O_159,N_2958,N_2946);
and UO_160 (O_160,N_2880,N_2994);
or UO_161 (O_161,N_2967,N_2937);
nand UO_162 (O_162,N_2894,N_2809);
nand UO_163 (O_163,N_2869,N_2931);
nor UO_164 (O_164,N_2926,N_2854);
and UO_165 (O_165,N_2949,N_2857);
nor UO_166 (O_166,N_2965,N_2824);
nand UO_167 (O_167,N_2986,N_2801);
or UO_168 (O_168,N_2993,N_2963);
or UO_169 (O_169,N_2925,N_2816);
or UO_170 (O_170,N_2989,N_2901);
nor UO_171 (O_171,N_2876,N_2836);
or UO_172 (O_172,N_2839,N_2808);
and UO_173 (O_173,N_2916,N_2905);
nand UO_174 (O_174,N_2969,N_2852);
nor UO_175 (O_175,N_2961,N_2844);
nor UO_176 (O_176,N_2838,N_2813);
or UO_177 (O_177,N_2901,N_2965);
nand UO_178 (O_178,N_2959,N_2802);
or UO_179 (O_179,N_2826,N_2966);
nand UO_180 (O_180,N_2907,N_2886);
or UO_181 (O_181,N_2934,N_2896);
or UO_182 (O_182,N_2995,N_2932);
or UO_183 (O_183,N_2856,N_2860);
nand UO_184 (O_184,N_2855,N_2852);
nor UO_185 (O_185,N_2800,N_2938);
or UO_186 (O_186,N_2959,N_2891);
or UO_187 (O_187,N_2882,N_2879);
or UO_188 (O_188,N_2922,N_2853);
and UO_189 (O_189,N_2917,N_2935);
nand UO_190 (O_190,N_2813,N_2831);
nor UO_191 (O_191,N_2932,N_2919);
or UO_192 (O_192,N_2987,N_2976);
nor UO_193 (O_193,N_2971,N_2820);
nand UO_194 (O_194,N_2985,N_2822);
nand UO_195 (O_195,N_2844,N_2828);
or UO_196 (O_196,N_2899,N_2941);
or UO_197 (O_197,N_2850,N_2994);
and UO_198 (O_198,N_2806,N_2889);
or UO_199 (O_199,N_2843,N_2927);
and UO_200 (O_200,N_2871,N_2986);
and UO_201 (O_201,N_2931,N_2875);
nand UO_202 (O_202,N_2910,N_2954);
and UO_203 (O_203,N_2839,N_2817);
nand UO_204 (O_204,N_2850,N_2807);
nand UO_205 (O_205,N_2852,N_2860);
or UO_206 (O_206,N_2980,N_2933);
nand UO_207 (O_207,N_2833,N_2934);
and UO_208 (O_208,N_2813,N_2805);
nor UO_209 (O_209,N_2833,N_2944);
and UO_210 (O_210,N_2978,N_2802);
nand UO_211 (O_211,N_2954,N_2978);
nand UO_212 (O_212,N_2864,N_2815);
nor UO_213 (O_213,N_2861,N_2812);
or UO_214 (O_214,N_2940,N_2998);
nand UO_215 (O_215,N_2871,N_2947);
nand UO_216 (O_216,N_2895,N_2871);
nand UO_217 (O_217,N_2909,N_2864);
and UO_218 (O_218,N_2810,N_2855);
and UO_219 (O_219,N_2993,N_2852);
and UO_220 (O_220,N_2913,N_2961);
or UO_221 (O_221,N_2930,N_2984);
nand UO_222 (O_222,N_2854,N_2821);
or UO_223 (O_223,N_2886,N_2960);
nand UO_224 (O_224,N_2841,N_2808);
and UO_225 (O_225,N_2938,N_2885);
and UO_226 (O_226,N_2921,N_2992);
and UO_227 (O_227,N_2886,N_2941);
nand UO_228 (O_228,N_2866,N_2953);
nand UO_229 (O_229,N_2869,N_2959);
and UO_230 (O_230,N_2852,N_2815);
and UO_231 (O_231,N_2992,N_2944);
nor UO_232 (O_232,N_2864,N_2932);
nand UO_233 (O_233,N_2805,N_2882);
or UO_234 (O_234,N_2876,N_2878);
nor UO_235 (O_235,N_2820,N_2954);
nor UO_236 (O_236,N_2955,N_2833);
and UO_237 (O_237,N_2820,N_2982);
or UO_238 (O_238,N_2842,N_2882);
nor UO_239 (O_239,N_2909,N_2875);
and UO_240 (O_240,N_2949,N_2914);
or UO_241 (O_241,N_2830,N_2965);
nor UO_242 (O_242,N_2897,N_2926);
and UO_243 (O_243,N_2936,N_2867);
or UO_244 (O_244,N_2866,N_2989);
or UO_245 (O_245,N_2870,N_2907);
nor UO_246 (O_246,N_2890,N_2846);
and UO_247 (O_247,N_2933,N_2833);
nand UO_248 (O_248,N_2902,N_2852);
or UO_249 (O_249,N_2814,N_2820);
nand UO_250 (O_250,N_2802,N_2817);
nand UO_251 (O_251,N_2898,N_2867);
nand UO_252 (O_252,N_2929,N_2875);
or UO_253 (O_253,N_2914,N_2827);
and UO_254 (O_254,N_2825,N_2847);
or UO_255 (O_255,N_2815,N_2814);
nand UO_256 (O_256,N_2864,N_2812);
or UO_257 (O_257,N_2936,N_2840);
nand UO_258 (O_258,N_2915,N_2944);
and UO_259 (O_259,N_2920,N_2996);
nor UO_260 (O_260,N_2941,N_2913);
nand UO_261 (O_261,N_2823,N_2928);
and UO_262 (O_262,N_2977,N_2888);
and UO_263 (O_263,N_2922,N_2926);
nor UO_264 (O_264,N_2994,N_2893);
and UO_265 (O_265,N_2861,N_2830);
nand UO_266 (O_266,N_2915,N_2913);
nor UO_267 (O_267,N_2849,N_2963);
nand UO_268 (O_268,N_2920,N_2891);
and UO_269 (O_269,N_2962,N_2978);
or UO_270 (O_270,N_2899,N_2896);
nor UO_271 (O_271,N_2831,N_2957);
nand UO_272 (O_272,N_2847,N_2820);
or UO_273 (O_273,N_2959,N_2941);
nor UO_274 (O_274,N_2954,N_2865);
nor UO_275 (O_275,N_2805,N_2865);
or UO_276 (O_276,N_2946,N_2840);
nor UO_277 (O_277,N_2905,N_2991);
or UO_278 (O_278,N_2982,N_2837);
nand UO_279 (O_279,N_2979,N_2863);
or UO_280 (O_280,N_2812,N_2954);
nor UO_281 (O_281,N_2909,N_2870);
or UO_282 (O_282,N_2958,N_2948);
and UO_283 (O_283,N_2927,N_2969);
or UO_284 (O_284,N_2890,N_2849);
and UO_285 (O_285,N_2803,N_2989);
and UO_286 (O_286,N_2929,N_2817);
nor UO_287 (O_287,N_2958,N_2982);
nor UO_288 (O_288,N_2879,N_2841);
or UO_289 (O_289,N_2824,N_2941);
and UO_290 (O_290,N_2925,N_2951);
and UO_291 (O_291,N_2884,N_2862);
and UO_292 (O_292,N_2955,N_2871);
nor UO_293 (O_293,N_2971,N_2879);
and UO_294 (O_294,N_2990,N_2823);
nor UO_295 (O_295,N_2832,N_2961);
nand UO_296 (O_296,N_2969,N_2877);
or UO_297 (O_297,N_2923,N_2848);
and UO_298 (O_298,N_2879,N_2898);
or UO_299 (O_299,N_2903,N_2875);
nand UO_300 (O_300,N_2997,N_2988);
nor UO_301 (O_301,N_2814,N_2955);
nand UO_302 (O_302,N_2838,N_2830);
nand UO_303 (O_303,N_2836,N_2924);
and UO_304 (O_304,N_2845,N_2897);
nor UO_305 (O_305,N_2853,N_2873);
or UO_306 (O_306,N_2879,N_2895);
nand UO_307 (O_307,N_2859,N_2930);
nor UO_308 (O_308,N_2926,N_2901);
nand UO_309 (O_309,N_2833,N_2846);
or UO_310 (O_310,N_2811,N_2883);
nor UO_311 (O_311,N_2819,N_2930);
nor UO_312 (O_312,N_2834,N_2908);
nand UO_313 (O_313,N_2906,N_2967);
or UO_314 (O_314,N_2893,N_2832);
nor UO_315 (O_315,N_2824,N_2855);
nor UO_316 (O_316,N_2959,N_2899);
nor UO_317 (O_317,N_2835,N_2901);
or UO_318 (O_318,N_2950,N_2994);
or UO_319 (O_319,N_2831,N_2935);
or UO_320 (O_320,N_2928,N_2884);
nand UO_321 (O_321,N_2813,N_2992);
or UO_322 (O_322,N_2963,N_2975);
or UO_323 (O_323,N_2842,N_2933);
or UO_324 (O_324,N_2995,N_2979);
or UO_325 (O_325,N_2804,N_2988);
or UO_326 (O_326,N_2844,N_2838);
and UO_327 (O_327,N_2993,N_2926);
or UO_328 (O_328,N_2994,N_2993);
and UO_329 (O_329,N_2921,N_2955);
nor UO_330 (O_330,N_2921,N_2959);
and UO_331 (O_331,N_2930,N_2970);
or UO_332 (O_332,N_2997,N_2828);
and UO_333 (O_333,N_2893,N_2901);
or UO_334 (O_334,N_2886,N_2873);
nand UO_335 (O_335,N_2961,N_2946);
and UO_336 (O_336,N_2828,N_2864);
and UO_337 (O_337,N_2838,N_2864);
nand UO_338 (O_338,N_2957,N_2975);
nand UO_339 (O_339,N_2814,N_2985);
nand UO_340 (O_340,N_2846,N_2983);
or UO_341 (O_341,N_2885,N_2852);
or UO_342 (O_342,N_2940,N_2947);
nor UO_343 (O_343,N_2883,N_2914);
and UO_344 (O_344,N_2959,N_2945);
nand UO_345 (O_345,N_2841,N_2891);
or UO_346 (O_346,N_2956,N_2965);
nand UO_347 (O_347,N_2952,N_2905);
and UO_348 (O_348,N_2905,N_2805);
or UO_349 (O_349,N_2995,N_2868);
or UO_350 (O_350,N_2902,N_2971);
nor UO_351 (O_351,N_2922,N_2813);
and UO_352 (O_352,N_2831,N_2942);
and UO_353 (O_353,N_2804,N_2912);
nor UO_354 (O_354,N_2930,N_2936);
nand UO_355 (O_355,N_2855,N_2983);
nand UO_356 (O_356,N_2899,N_2876);
and UO_357 (O_357,N_2984,N_2910);
and UO_358 (O_358,N_2884,N_2967);
nor UO_359 (O_359,N_2870,N_2915);
nand UO_360 (O_360,N_2807,N_2982);
nor UO_361 (O_361,N_2887,N_2913);
nand UO_362 (O_362,N_2884,N_2910);
nand UO_363 (O_363,N_2910,N_2944);
and UO_364 (O_364,N_2877,N_2940);
nand UO_365 (O_365,N_2892,N_2840);
nand UO_366 (O_366,N_2931,N_2909);
or UO_367 (O_367,N_2974,N_2876);
nand UO_368 (O_368,N_2956,N_2857);
or UO_369 (O_369,N_2969,N_2995);
or UO_370 (O_370,N_2961,N_2885);
or UO_371 (O_371,N_2910,N_2938);
nand UO_372 (O_372,N_2900,N_2938);
nor UO_373 (O_373,N_2983,N_2987);
nand UO_374 (O_374,N_2997,N_2820);
and UO_375 (O_375,N_2949,N_2952);
nor UO_376 (O_376,N_2878,N_2937);
nand UO_377 (O_377,N_2981,N_2980);
or UO_378 (O_378,N_2901,N_2889);
or UO_379 (O_379,N_2923,N_2882);
or UO_380 (O_380,N_2959,N_2882);
and UO_381 (O_381,N_2886,N_2804);
nor UO_382 (O_382,N_2837,N_2936);
nor UO_383 (O_383,N_2808,N_2919);
nor UO_384 (O_384,N_2846,N_2940);
nor UO_385 (O_385,N_2947,N_2904);
or UO_386 (O_386,N_2956,N_2871);
or UO_387 (O_387,N_2812,N_2890);
nor UO_388 (O_388,N_2881,N_2889);
nand UO_389 (O_389,N_2944,N_2873);
nand UO_390 (O_390,N_2821,N_2838);
nor UO_391 (O_391,N_2955,N_2943);
or UO_392 (O_392,N_2922,N_2837);
and UO_393 (O_393,N_2844,N_2909);
or UO_394 (O_394,N_2874,N_2958);
nor UO_395 (O_395,N_2800,N_2978);
nand UO_396 (O_396,N_2882,N_2920);
nor UO_397 (O_397,N_2945,N_2979);
nor UO_398 (O_398,N_2941,N_2891);
nand UO_399 (O_399,N_2894,N_2991);
nor UO_400 (O_400,N_2968,N_2923);
and UO_401 (O_401,N_2921,N_2980);
or UO_402 (O_402,N_2863,N_2909);
or UO_403 (O_403,N_2833,N_2870);
or UO_404 (O_404,N_2827,N_2892);
nor UO_405 (O_405,N_2893,N_2992);
nor UO_406 (O_406,N_2963,N_2927);
nand UO_407 (O_407,N_2808,N_2976);
nor UO_408 (O_408,N_2904,N_2901);
nor UO_409 (O_409,N_2822,N_2947);
nor UO_410 (O_410,N_2816,N_2990);
or UO_411 (O_411,N_2927,N_2987);
and UO_412 (O_412,N_2840,N_2989);
and UO_413 (O_413,N_2975,N_2815);
or UO_414 (O_414,N_2832,N_2836);
and UO_415 (O_415,N_2900,N_2995);
nand UO_416 (O_416,N_2905,N_2989);
nor UO_417 (O_417,N_2810,N_2911);
nand UO_418 (O_418,N_2885,N_2823);
nor UO_419 (O_419,N_2865,N_2903);
or UO_420 (O_420,N_2923,N_2880);
nand UO_421 (O_421,N_2968,N_2838);
or UO_422 (O_422,N_2958,N_2867);
or UO_423 (O_423,N_2822,N_2900);
nor UO_424 (O_424,N_2994,N_2841);
and UO_425 (O_425,N_2949,N_2919);
and UO_426 (O_426,N_2918,N_2957);
or UO_427 (O_427,N_2843,N_2925);
and UO_428 (O_428,N_2984,N_2828);
or UO_429 (O_429,N_2968,N_2927);
nand UO_430 (O_430,N_2881,N_2866);
nand UO_431 (O_431,N_2875,N_2958);
nand UO_432 (O_432,N_2995,N_2989);
and UO_433 (O_433,N_2867,N_2860);
or UO_434 (O_434,N_2974,N_2875);
and UO_435 (O_435,N_2812,N_2883);
nand UO_436 (O_436,N_2983,N_2972);
nand UO_437 (O_437,N_2907,N_2943);
nand UO_438 (O_438,N_2855,N_2961);
nor UO_439 (O_439,N_2973,N_2992);
nand UO_440 (O_440,N_2805,N_2815);
or UO_441 (O_441,N_2987,N_2991);
or UO_442 (O_442,N_2934,N_2936);
and UO_443 (O_443,N_2853,N_2887);
or UO_444 (O_444,N_2973,N_2809);
or UO_445 (O_445,N_2934,N_2996);
and UO_446 (O_446,N_2833,N_2903);
and UO_447 (O_447,N_2998,N_2805);
nor UO_448 (O_448,N_2949,N_2827);
nand UO_449 (O_449,N_2954,N_2881);
nor UO_450 (O_450,N_2993,N_2819);
and UO_451 (O_451,N_2857,N_2997);
xnor UO_452 (O_452,N_2836,N_2993);
nor UO_453 (O_453,N_2802,N_2982);
nor UO_454 (O_454,N_2961,N_2847);
and UO_455 (O_455,N_2830,N_2883);
or UO_456 (O_456,N_2949,N_2965);
or UO_457 (O_457,N_2932,N_2872);
nand UO_458 (O_458,N_2916,N_2953);
nor UO_459 (O_459,N_2988,N_2959);
and UO_460 (O_460,N_2876,N_2993);
nor UO_461 (O_461,N_2855,N_2888);
or UO_462 (O_462,N_2951,N_2987);
and UO_463 (O_463,N_2961,N_2821);
nand UO_464 (O_464,N_2929,N_2937);
nand UO_465 (O_465,N_2945,N_2824);
nor UO_466 (O_466,N_2947,N_2920);
nor UO_467 (O_467,N_2948,N_2978);
nor UO_468 (O_468,N_2869,N_2957);
or UO_469 (O_469,N_2924,N_2928);
nand UO_470 (O_470,N_2814,N_2965);
nand UO_471 (O_471,N_2990,N_2929);
or UO_472 (O_472,N_2969,N_2998);
and UO_473 (O_473,N_2901,N_2894);
nand UO_474 (O_474,N_2859,N_2994);
or UO_475 (O_475,N_2809,N_2869);
nor UO_476 (O_476,N_2889,N_2815);
or UO_477 (O_477,N_2941,N_2820);
nor UO_478 (O_478,N_2818,N_2915);
nand UO_479 (O_479,N_2904,N_2823);
and UO_480 (O_480,N_2932,N_2863);
and UO_481 (O_481,N_2901,N_2982);
nor UO_482 (O_482,N_2940,N_2882);
nand UO_483 (O_483,N_2804,N_2932);
nand UO_484 (O_484,N_2991,N_2950);
nand UO_485 (O_485,N_2880,N_2955);
nand UO_486 (O_486,N_2874,N_2846);
and UO_487 (O_487,N_2867,N_2864);
nand UO_488 (O_488,N_2915,N_2843);
nor UO_489 (O_489,N_2808,N_2828);
nor UO_490 (O_490,N_2906,N_2953);
nor UO_491 (O_491,N_2803,N_2967);
or UO_492 (O_492,N_2930,N_2963);
nor UO_493 (O_493,N_2840,N_2885);
and UO_494 (O_494,N_2897,N_2964);
nor UO_495 (O_495,N_2881,N_2822);
nor UO_496 (O_496,N_2882,N_2891);
or UO_497 (O_497,N_2807,N_2811);
or UO_498 (O_498,N_2942,N_2952);
and UO_499 (O_499,N_2945,N_2923);
endmodule