module basic_1000_10000_1500_5_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
xor U0 (N_0,In_350,In_921);
and U1 (N_1,In_108,In_263);
nor U2 (N_2,In_101,In_120);
nand U3 (N_3,In_897,In_713);
xor U4 (N_4,In_388,In_430);
and U5 (N_5,In_714,In_462);
and U6 (N_6,In_300,In_222);
xor U7 (N_7,In_335,In_759);
xnor U8 (N_8,In_236,In_203);
nor U9 (N_9,In_737,In_984);
nand U10 (N_10,In_319,In_329);
and U11 (N_11,In_52,In_751);
or U12 (N_12,In_231,In_40);
xor U13 (N_13,In_461,In_410);
nor U14 (N_14,In_696,In_559);
nor U15 (N_15,In_7,In_772);
and U16 (N_16,In_411,In_637);
nand U17 (N_17,In_389,In_578);
nand U18 (N_18,In_249,In_378);
and U19 (N_19,In_692,In_164);
xor U20 (N_20,In_936,In_910);
and U21 (N_21,In_434,In_975);
nor U22 (N_22,In_178,In_163);
or U23 (N_23,In_351,In_254);
nand U24 (N_24,In_546,In_720);
nor U25 (N_25,In_962,In_602);
xor U26 (N_26,In_556,In_938);
or U27 (N_27,In_153,In_133);
xnor U28 (N_28,In_683,In_827);
nor U29 (N_29,In_986,In_483);
xor U30 (N_30,In_68,In_707);
and U31 (N_31,In_767,In_186);
or U32 (N_32,In_193,In_402);
and U33 (N_33,In_87,In_875);
and U34 (N_34,In_640,In_492);
nand U35 (N_35,In_477,In_849);
and U36 (N_36,In_860,In_668);
or U37 (N_37,In_927,In_204);
and U38 (N_38,In_960,In_816);
xnor U39 (N_39,In_491,In_784);
nand U40 (N_40,In_903,In_673);
nor U41 (N_41,In_13,In_45);
nor U42 (N_42,In_62,In_294);
xnor U43 (N_43,In_829,In_918);
nor U44 (N_44,In_939,In_850);
xor U45 (N_45,In_213,In_722);
and U46 (N_46,In_252,In_919);
or U47 (N_47,In_914,In_297);
or U48 (N_48,In_83,In_620);
and U49 (N_49,In_451,In_316);
or U50 (N_50,In_349,In_266);
or U51 (N_51,In_224,In_457);
and U52 (N_52,In_409,In_991);
nor U53 (N_53,In_216,In_736);
xnor U54 (N_54,In_745,In_848);
nor U55 (N_55,In_876,In_900);
nand U56 (N_56,In_616,In_332);
or U57 (N_57,In_306,In_398);
and U58 (N_58,In_889,In_902);
nor U59 (N_59,In_522,In_576);
nand U60 (N_60,In_301,In_77);
and U61 (N_61,In_499,In_156);
or U62 (N_62,In_128,In_192);
nand U63 (N_63,In_700,In_519);
xor U64 (N_64,In_652,In_479);
nor U65 (N_65,In_75,In_412);
or U66 (N_66,In_752,In_78);
nand U67 (N_67,In_29,In_787);
or U68 (N_68,In_670,In_183);
nand U69 (N_69,In_452,In_314);
xnor U70 (N_70,In_196,In_702);
or U71 (N_71,In_25,In_654);
and U72 (N_72,In_417,In_563);
and U73 (N_73,In_917,In_210);
or U74 (N_74,In_436,In_84);
or U75 (N_75,In_539,In_221);
nand U76 (N_76,In_633,In_564);
nor U77 (N_77,In_425,In_964);
and U78 (N_78,In_107,In_968);
nor U79 (N_79,In_413,In_624);
nor U80 (N_80,In_494,In_414);
and U81 (N_81,In_540,In_998);
xnor U82 (N_82,In_172,In_923);
nand U83 (N_83,In_21,In_106);
nand U84 (N_84,In_17,In_547);
nand U85 (N_85,In_854,In_873);
and U86 (N_86,In_131,In_869);
nor U87 (N_87,In_138,In_116);
xor U88 (N_88,In_646,In_308);
or U89 (N_89,In_315,In_608);
or U90 (N_90,In_650,In_542);
nand U91 (N_91,In_994,In_996);
or U92 (N_92,In_672,In_733);
xor U93 (N_93,In_43,In_112);
xor U94 (N_94,In_46,In_580);
and U95 (N_95,In_780,In_235);
nor U96 (N_96,In_292,In_606);
nand U97 (N_97,In_230,In_219);
xnor U98 (N_98,In_495,In_201);
or U99 (N_99,In_225,In_88);
and U100 (N_100,In_730,In_568);
nand U101 (N_101,In_475,In_282);
nand U102 (N_102,In_326,In_42);
xnor U103 (N_103,In_992,In_480);
nor U104 (N_104,In_358,In_956);
nor U105 (N_105,In_125,In_803);
or U106 (N_106,In_701,In_603);
xnor U107 (N_107,In_129,In_93);
and U108 (N_108,In_949,In_528);
and U109 (N_109,In_792,In_171);
xor U110 (N_110,In_864,In_508);
and U111 (N_111,In_521,In_699);
nor U112 (N_112,In_832,In_643);
and U113 (N_113,In_360,In_940);
xnor U114 (N_114,In_657,In_317);
nand U115 (N_115,In_506,In_122);
nand U116 (N_116,In_989,In_238);
nand U117 (N_117,In_498,In_882);
xor U118 (N_118,In_888,In_9);
xor U119 (N_119,In_53,In_309);
xnor U120 (N_120,In_271,In_515);
xnor U121 (N_121,In_373,In_143);
nand U122 (N_122,In_887,In_245);
or U123 (N_123,In_912,In_340);
or U124 (N_124,In_159,In_783);
xor U125 (N_125,In_232,In_132);
or U126 (N_126,In_770,In_950);
xnor U127 (N_127,In_323,In_92);
and U128 (N_128,In_154,In_200);
nand U129 (N_129,In_435,In_740);
xor U130 (N_130,In_146,In_313);
nand U131 (N_131,In_771,In_706);
nor U132 (N_132,In_255,In_845);
nor U133 (N_133,In_680,In_202);
and U134 (N_134,In_513,In_27);
nor U135 (N_135,In_212,In_644);
and U136 (N_136,In_913,In_575);
nor U137 (N_137,In_874,In_325);
nor U138 (N_138,In_113,In_932);
nand U139 (N_139,In_48,In_839);
or U140 (N_140,In_518,In_344);
nor U141 (N_141,In_166,In_541);
nor U142 (N_142,In_181,In_781);
nand U143 (N_143,In_215,In_432);
nor U144 (N_144,In_127,In_507);
and U145 (N_145,In_291,In_898);
and U146 (N_146,In_367,In_584);
and U147 (N_147,In_961,In_558);
nand U148 (N_148,In_35,In_866);
and U149 (N_149,In_26,In_243);
nor U150 (N_150,In_195,In_459);
and U151 (N_151,In_175,In_555);
xnor U152 (N_152,In_844,In_334);
and U153 (N_153,In_90,In_32);
xor U154 (N_154,In_247,In_237);
nor U155 (N_155,In_81,In_636);
xor U156 (N_156,In_762,In_658);
xnor U157 (N_157,In_299,In_551);
nor U158 (N_158,In_867,In_728);
or U159 (N_159,In_375,In_86);
and U160 (N_160,In_988,In_211);
or U161 (N_161,In_597,In_524);
xor U162 (N_162,In_532,In_741);
xor U163 (N_163,In_843,In_727);
xor U164 (N_164,In_865,In_951);
nand U165 (N_165,In_152,In_520);
and U166 (N_166,In_614,In_69);
nand U167 (N_167,In_331,In_416);
xnor U168 (N_168,In_993,In_579);
or U169 (N_169,In_905,In_831);
or U170 (N_170,In_3,In_997);
and U171 (N_171,In_486,In_530);
or U172 (N_172,In_681,In_338);
and U173 (N_173,In_362,In_943);
or U174 (N_174,In_320,In_944);
nor U175 (N_175,In_565,In_408);
xor U176 (N_176,In_871,In_621);
nand U177 (N_177,In_695,In_777);
nand U178 (N_178,In_383,In_611);
or U179 (N_179,In_123,In_447);
or U180 (N_180,In_667,In_110);
or U181 (N_181,In_440,In_798);
and U182 (N_182,In_158,In_478);
nor U183 (N_183,In_769,In_509);
nand U184 (N_184,In_420,In_969);
nor U185 (N_185,In_885,In_191);
xor U186 (N_186,In_339,In_180);
and U187 (N_187,In_895,In_501);
nand U188 (N_188,In_41,In_293);
or U189 (N_189,In_909,In_703);
nor U190 (N_190,In_439,In_76);
nand U191 (N_191,In_795,In_653);
xnor U192 (N_192,In_16,In_856);
and U193 (N_193,In_742,In_296);
xor U194 (N_194,In_725,In_708);
nand U195 (N_195,In_226,In_645);
nor U196 (N_196,In_954,In_719);
nor U197 (N_197,In_259,In_37);
nor U198 (N_198,In_791,In_374);
nor U199 (N_199,In_91,In_970);
nor U200 (N_200,In_270,In_709);
nand U201 (N_201,In_666,In_162);
or U202 (N_202,In_405,In_881);
or U203 (N_203,In_361,In_626);
nor U204 (N_204,In_96,In_89);
nor U205 (N_205,In_295,In_161);
and U206 (N_206,In_935,In_277);
nand U207 (N_207,In_734,In_472);
or U208 (N_208,In_167,In_582);
nor U209 (N_209,In_899,In_952);
nand U210 (N_210,In_863,In_444);
and U211 (N_211,In_2,In_80);
xnor U212 (N_212,In_466,In_47);
nor U213 (N_213,In_258,In_922);
and U214 (N_214,In_214,In_104);
and U215 (N_215,In_925,In_594);
nor U216 (N_216,In_124,In_766);
nand U217 (N_217,In_613,In_851);
nand U218 (N_218,In_688,In_468);
xor U219 (N_219,In_286,In_911);
or U220 (N_220,In_945,In_396);
xnor U221 (N_221,In_879,In_647);
nand U222 (N_222,In_930,In_12);
nand U223 (N_223,In_562,In_363);
xnor U224 (N_224,In_841,In_233);
and U225 (N_225,In_639,In_959);
nor U226 (N_226,In_70,In_431);
xor U227 (N_227,In_890,In_729);
and U228 (N_228,In_712,In_241);
nor U229 (N_229,In_693,In_946);
nor U230 (N_230,In_407,In_982);
and U231 (N_231,In_976,In_567);
and U232 (N_232,In_983,In_469);
xnor U233 (N_233,In_625,In_460);
or U234 (N_234,In_144,In_303);
or U235 (N_235,In_797,In_114);
nor U236 (N_236,In_785,In_561);
xnor U237 (N_237,In_817,In_768);
nand U238 (N_238,In_607,In_30);
xnor U239 (N_239,In_5,In_929);
or U240 (N_240,In_760,In_638);
or U241 (N_241,In_788,In_280);
xnor U242 (N_242,In_310,In_800);
and U243 (N_243,In_596,In_371);
and U244 (N_244,In_738,In_281);
and U245 (N_245,In_6,In_105);
xor U246 (N_246,In_268,In_49);
nor U247 (N_247,In_557,In_324);
xor U248 (N_248,In_206,In_907);
xor U249 (N_249,In_786,In_58);
or U250 (N_250,In_586,In_406);
nand U251 (N_251,In_789,In_823);
or U252 (N_252,In_333,In_208);
xnor U253 (N_253,In_691,In_599);
nor U254 (N_254,In_168,In_641);
or U255 (N_255,In_117,In_73);
nand U256 (N_256,In_525,In_775);
nand U257 (N_257,In_972,In_239);
nor U258 (N_258,In_187,In_763);
and U259 (N_259,In_481,In_651);
or U260 (N_260,In_753,In_779);
nand U261 (N_261,In_31,In_353);
xor U262 (N_262,In_391,In_676);
and U263 (N_263,In_610,In_23);
xnor U264 (N_264,In_537,In_504);
nor U265 (N_265,In_977,In_790);
or U266 (N_266,In_318,In_279);
nand U267 (N_267,In_227,In_514);
and U268 (N_268,In_446,In_445);
nor U269 (N_269,In_357,In_174);
nor U270 (N_270,In_442,In_978);
xor U271 (N_271,In_746,In_853);
nor U272 (N_272,In_56,In_176);
nor U273 (N_273,In_529,In_99);
and U274 (N_274,In_473,In_773);
xor U275 (N_275,In_822,In_137);
and U276 (N_276,In_838,In_593);
nand U277 (N_277,In_679,In_601);
and U278 (N_278,In_312,In_937);
and U279 (N_279,In_517,In_39);
and U280 (N_280,In_355,In_552);
and U281 (N_281,In_828,In_534);
xnor U282 (N_282,In_207,In_502);
or U283 (N_283,In_415,In_732);
xor U284 (N_284,In_140,In_242);
nand U285 (N_285,In_18,In_20);
and U286 (N_286,In_503,In_560);
and U287 (N_287,In_595,In_482);
and U288 (N_288,In_674,In_980);
xnor U289 (N_289,In_179,In_750);
and U290 (N_290,In_628,In_22);
and U291 (N_291,In_554,In_543);
nor U292 (N_292,In_450,In_678);
nor U293 (N_293,In_967,In_382);
xor U294 (N_294,In_920,In_218);
or U295 (N_295,In_648,In_404);
or U296 (N_296,In_527,In_883);
or U297 (N_297,In_392,In_669);
and U298 (N_298,In_878,In_928);
and U299 (N_299,In_393,In_684);
nand U300 (N_300,In_533,In_585);
xnor U301 (N_301,In_663,In_72);
nand U302 (N_302,In_948,In_427);
nand U303 (N_303,In_642,In_223);
nand U304 (N_304,In_687,In_453);
nor U305 (N_305,In_199,In_184);
nand U306 (N_306,In_896,In_609);
nor U307 (N_307,In_169,In_372);
or U308 (N_308,In_799,In_685);
nor U309 (N_309,In_71,In_627);
nand U310 (N_310,In_130,In_465);
xnor U311 (N_311,In_493,In_535);
or U312 (N_312,In_100,In_135);
and U313 (N_313,In_150,In_868);
and U314 (N_314,In_573,In_671);
nor U315 (N_315,In_1,In_188);
and U316 (N_316,In_328,In_51);
or U317 (N_317,In_198,In_748);
xnor U318 (N_318,In_209,In_605);
nor U319 (N_319,In_892,In_464);
or U320 (N_320,In_302,In_136);
xnor U321 (N_321,In_428,In_587);
nor U322 (N_322,In_583,In_805);
nor U323 (N_323,In_19,In_471);
or U324 (N_324,In_833,In_723);
and U325 (N_325,In_111,In_754);
and U326 (N_326,In_103,In_272);
xnor U327 (N_327,In_757,In_484);
xnor U328 (N_328,In_656,In_617);
nand U329 (N_329,In_505,In_689);
xor U330 (N_330,In_148,In_500);
or U331 (N_331,In_747,In_488);
or U332 (N_332,In_884,In_433);
and U333 (N_333,In_386,In_267);
xor U334 (N_334,In_682,In_731);
and U335 (N_335,In_716,In_155);
xor U336 (N_336,In_995,In_458);
xnor U337 (N_337,In_631,In_476);
xor U338 (N_338,In_283,In_229);
or U339 (N_339,In_470,In_830);
xnor U340 (N_340,In_749,In_61);
and U341 (N_341,In_837,In_804);
xor U342 (N_342,In_244,In_194);
xnor U343 (N_343,In_630,In_836);
nor U344 (N_344,In_955,In_387);
nor U345 (N_345,In_441,In_973);
nand U346 (N_346,In_304,In_926);
xor U347 (N_347,In_74,In_661);
and U348 (N_348,In_801,In_15);
nand U349 (N_349,In_36,In_429);
or U350 (N_350,In_764,In_10);
nor U351 (N_351,In_510,In_877);
xor U352 (N_352,In_342,In_177);
xnor U353 (N_353,In_275,In_311);
nand U354 (N_354,In_958,In_102);
and U355 (N_355,In_336,In_818);
or U356 (N_356,In_343,In_377);
and U357 (N_357,In_705,In_234);
nand U358 (N_358,In_619,In_717);
xor U359 (N_359,In_821,In_807);
and U360 (N_360,In_965,In_577);
or U361 (N_361,In_197,In_173);
nor U362 (N_362,In_690,In_953);
nand U363 (N_363,In_812,In_697);
and U364 (N_364,In_901,In_893);
nand U365 (N_365,In_571,In_497);
or U366 (N_366,In_966,In_276);
nand U367 (N_367,In_835,In_778);
nand U368 (N_368,In_395,In_842);
nand U369 (N_369,In_126,In_886);
nor U370 (N_370,In_285,In_813);
and U371 (N_371,In_793,In_635);
and U372 (N_372,In_947,In_257);
xor U373 (N_373,In_54,In_721);
nor U374 (N_374,In_544,In_44);
or U375 (N_375,In_134,In_660);
or U376 (N_376,In_981,In_744);
and U377 (N_377,In_489,In_456);
nand U378 (N_378,In_858,In_756);
nand U379 (N_379,In_999,In_906);
xor U380 (N_380,In_846,In_354);
nand U381 (N_381,In_327,In_776);
and U382 (N_382,In_589,In_347);
nor U383 (N_383,In_265,In_57);
or U384 (N_384,In_824,In_806);
xor U385 (N_385,In_485,In_401);
xnor U386 (N_386,In_248,In_287);
nor U387 (N_387,In_284,In_550);
nand U388 (N_388,In_380,In_337);
or U389 (N_389,In_810,In_298);
and U390 (N_390,In_145,In_189);
nand U391 (N_391,In_139,In_151);
xor U392 (N_392,In_278,In_394);
and U393 (N_393,In_261,In_384);
nor U394 (N_394,In_437,In_85);
or U395 (N_395,In_761,In_686);
nor U396 (N_396,In_63,In_979);
xnor U397 (N_397,In_59,In_400);
or U398 (N_398,In_809,In_369);
and U399 (N_399,In_160,In_185);
or U400 (N_400,In_79,In_264);
nand U401 (N_401,In_659,In_904);
xor U402 (N_402,In_418,In_675);
and U403 (N_403,In_811,In_538);
or U404 (N_404,In_352,In_205);
and U405 (N_405,In_894,In_574);
or U406 (N_406,In_289,In_694);
xor U407 (N_407,In_64,In_253);
and U408 (N_408,In_794,In_825);
nand U409 (N_409,In_840,In_269);
nand U410 (N_410,In_545,In_115);
xnor U411 (N_411,In_739,In_512);
and U412 (N_412,In_14,In_33);
xor U413 (N_413,In_250,In_322);
nand U414 (N_414,In_632,In_649);
and U415 (N_415,In_397,In_516);
nand U416 (N_416,In_119,In_872);
and U417 (N_417,In_487,In_572);
xnor U418 (N_418,In_370,In_755);
nor U419 (N_419,In_50,In_399);
or U420 (N_420,In_288,In_251);
xnor U421 (N_421,In_655,In_665);
nor U422 (N_422,In_847,In_861);
xor U423 (N_423,In_743,In_455);
nand U424 (N_424,In_422,In_403);
nand U425 (N_425,In_622,In_536);
nor U426 (N_426,In_726,In_782);
or U427 (N_427,In_467,In_165);
xnor U428 (N_428,In_11,In_870);
xor U429 (N_429,In_933,In_570);
xnor U430 (N_430,In_364,In_274);
nand U431 (N_431,In_4,In_141);
nor U432 (N_432,In_862,In_941);
xnor U433 (N_433,In_94,In_109);
nand U434 (N_434,In_256,In_618);
and U435 (N_435,In_97,In_985);
and U436 (N_436,In_931,In_463);
and U437 (N_437,In_423,In_758);
nor U438 (N_438,In_548,In_710);
or U439 (N_439,In_365,In_600);
and U440 (N_440,In_149,In_915);
or U441 (N_441,In_808,In_379);
xnor U442 (N_442,In_341,In_170);
nand U443 (N_443,In_490,In_531);
and U444 (N_444,In_449,In_591);
nor U445 (N_445,In_924,In_346);
or U446 (N_446,In_217,In_942);
xnor U447 (N_447,In_348,In_549);
and U448 (N_448,In_859,In_60);
xnor U449 (N_449,In_424,In_95);
and U450 (N_450,In_55,In_240);
or U451 (N_451,In_834,In_511);
nor U452 (N_452,In_366,In_704);
nand U453 (N_453,In_629,In_443);
or U454 (N_454,In_8,In_880);
nand U455 (N_455,In_677,In_774);
xnor U456 (N_456,In_82,In_474);
nand U457 (N_457,In_796,In_290);
nor U458 (N_458,In_523,In_228);
xnor U459 (N_459,In_971,In_496);
xor U460 (N_460,In_592,In_765);
or U461 (N_461,In_569,In_246);
or U462 (N_462,In_65,In_987);
xnor U463 (N_463,In_623,In_157);
or U464 (N_464,In_916,In_934);
and U465 (N_465,In_454,In_990);
nand U466 (N_466,In_34,In_0);
nor U467 (N_467,In_664,In_28);
and U468 (N_468,In_67,In_121);
nand U469 (N_469,In_735,In_38);
nand U470 (N_470,In_826,In_526);
nand U471 (N_471,In_260,In_852);
nor U472 (N_472,In_385,In_820);
xnor U473 (N_473,In_356,In_553);
and U474 (N_474,In_590,In_66);
xnor U475 (N_475,In_390,In_345);
nand U476 (N_476,In_815,In_963);
xor U477 (N_477,In_24,In_724);
nand U478 (N_478,In_448,In_718);
and U479 (N_479,In_305,In_802);
and U480 (N_480,In_598,In_190);
xnor U481 (N_481,In_98,In_604);
nor U482 (N_482,In_588,In_974);
nand U483 (N_483,In_891,In_612);
and U484 (N_484,In_142,In_814);
xnor U485 (N_485,In_438,In_698);
xnor U486 (N_486,In_419,In_634);
or U487 (N_487,In_857,In_321);
xor U488 (N_488,In_957,In_855);
and U489 (N_489,In_662,In_381);
and U490 (N_490,In_182,In_262);
nand U491 (N_491,In_581,In_220);
nand U492 (N_492,In_715,In_118);
nand U493 (N_493,In_330,In_368);
nor U494 (N_494,In_359,In_711);
nor U495 (N_495,In_908,In_421);
xor U496 (N_496,In_147,In_376);
nor U497 (N_497,In_819,In_426);
xnor U498 (N_498,In_273,In_615);
nor U499 (N_499,In_307,In_566);
nand U500 (N_500,In_682,In_30);
or U501 (N_501,In_446,In_959);
and U502 (N_502,In_231,In_464);
and U503 (N_503,In_761,In_99);
nand U504 (N_504,In_550,In_699);
and U505 (N_505,In_235,In_624);
nand U506 (N_506,In_182,In_479);
nor U507 (N_507,In_629,In_803);
nor U508 (N_508,In_174,In_607);
nor U509 (N_509,In_363,In_640);
xnor U510 (N_510,In_433,In_911);
nor U511 (N_511,In_862,In_566);
or U512 (N_512,In_780,In_75);
nor U513 (N_513,In_249,In_159);
nand U514 (N_514,In_212,In_916);
and U515 (N_515,In_124,In_73);
nand U516 (N_516,In_714,In_628);
nand U517 (N_517,In_879,In_111);
and U518 (N_518,In_224,In_135);
xor U519 (N_519,In_904,In_935);
and U520 (N_520,In_162,In_427);
nand U521 (N_521,In_226,In_559);
nor U522 (N_522,In_279,In_112);
and U523 (N_523,In_397,In_626);
and U524 (N_524,In_990,In_481);
nand U525 (N_525,In_257,In_138);
nor U526 (N_526,In_574,In_34);
or U527 (N_527,In_754,In_976);
nor U528 (N_528,In_746,In_975);
or U529 (N_529,In_691,In_59);
nand U530 (N_530,In_970,In_622);
xnor U531 (N_531,In_393,In_108);
and U532 (N_532,In_609,In_30);
xor U533 (N_533,In_840,In_674);
nor U534 (N_534,In_491,In_663);
nand U535 (N_535,In_501,In_284);
xnor U536 (N_536,In_776,In_840);
nand U537 (N_537,In_741,In_539);
and U538 (N_538,In_63,In_495);
nand U539 (N_539,In_390,In_836);
nor U540 (N_540,In_482,In_277);
nand U541 (N_541,In_221,In_882);
or U542 (N_542,In_528,In_696);
nor U543 (N_543,In_386,In_973);
nor U544 (N_544,In_274,In_311);
nor U545 (N_545,In_15,In_342);
xor U546 (N_546,In_332,In_473);
and U547 (N_547,In_779,In_750);
and U548 (N_548,In_943,In_870);
and U549 (N_549,In_336,In_51);
xnor U550 (N_550,In_903,In_113);
xor U551 (N_551,In_376,In_445);
xnor U552 (N_552,In_61,In_81);
and U553 (N_553,In_568,In_29);
or U554 (N_554,In_52,In_282);
and U555 (N_555,In_190,In_894);
and U556 (N_556,In_178,In_654);
nor U557 (N_557,In_770,In_96);
and U558 (N_558,In_104,In_17);
or U559 (N_559,In_67,In_865);
and U560 (N_560,In_515,In_394);
nor U561 (N_561,In_506,In_29);
or U562 (N_562,In_259,In_469);
and U563 (N_563,In_588,In_552);
nor U564 (N_564,In_877,In_225);
nand U565 (N_565,In_363,In_98);
and U566 (N_566,In_10,In_944);
nor U567 (N_567,In_189,In_161);
or U568 (N_568,In_407,In_672);
or U569 (N_569,In_827,In_913);
and U570 (N_570,In_242,In_770);
or U571 (N_571,In_501,In_567);
and U572 (N_572,In_262,In_506);
or U573 (N_573,In_463,In_154);
xor U574 (N_574,In_711,In_251);
xnor U575 (N_575,In_701,In_229);
and U576 (N_576,In_791,In_487);
nand U577 (N_577,In_965,In_172);
nand U578 (N_578,In_296,In_117);
xnor U579 (N_579,In_518,In_692);
nor U580 (N_580,In_642,In_189);
or U581 (N_581,In_306,In_685);
or U582 (N_582,In_764,In_343);
and U583 (N_583,In_978,In_936);
nor U584 (N_584,In_164,In_507);
or U585 (N_585,In_460,In_61);
xor U586 (N_586,In_853,In_647);
nor U587 (N_587,In_166,In_869);
and U588 (N_588,In_238,In_769);
nand U589 (N_589,In_645,In_361);
nand U590 (N_590,In_725,In_961);
and U591 (N_591,In_34,In_192);
nand U592 (N_592,In_365,In_47);
nor U593 (N_593,In_272,In_294);
xnor U594 (N_594,In_971,In_611);
nand U595 (N_595,In_860,In_176);
or U596 (N_596,In_110,In_517);
nor U597 (N_597,In_651,In_589);
xnor U598 (N_598,In_134,In_74);
nor U599 (N_599,In_320,In_891);
or U600 (N_600,In_875,In_608);
nor U601 (N_601,In_610,In_419);
nand U602 (N_602,In_520,In_471);
nand U603 (N_603,In_215,In_861);
nor U604 (N_604,In_504,In_499);
nor U605 (N_605,In_185,In_801);
or U606 (N_606,In_988,In_3);
xnor U607 (N_607,In_250,In_575);
or U608 (N_608,In_987,In_676);
and U609 (N_609,In_870,In_570);
nor U610 (N_610,In_282,In_380);
xor U611 (N_611,In_818,In_507);
nor U612 (N_612,In_63,In_123);
and U613 (N_613,In_470,In_675);
xnor U614 (N_614,In_795,In_407);
nand U615 (N_615,In_899,In_687);
and U616 (N_616,In_40,In_270);
and U617 (N_617,In_200,In_253);
xnor U618 (N_618,In_959,In_770);
or U619 (N_619,In_199,In_403);
nor U620 (N_620,In_721,In_987);
or U621 (N_621,In_227,In_654);
and U622 (N_622,In_305,In_93);
nor U623 (N_623,In_503,In_473);
or U624 (N_624,In_252,In_391);
nor U625 (N_625,In_832,In_512);
and U626 (N_626,In_368,In_197);
nand U627 (N_627,In_884,In_349);
nand U628 (N_628,In_534,In_528);
and U629 (N_629,In_468,In_862);
or U630 (N_630,In_511,In_903);
or U631 (N_631,In_142,In_350);
nor U632 (N_632,In_501,In_411);
nor U633 (N_633,In_900,In_943);
and U634 (N_634,In_951,In_916);
and U635 (N_635,In_194,In_393);
and U636 (N_636,In_84,In_262);
xnor U637 (N_637,In_323,In_714);
or U638 (N_638,In_802,In_611);
nand U639 (N_639,In_735,In_89);
nor U640 (N_640,In_649,In_325);
xnor U641 (N_641,In_700,In_240);
and U642 (N_642,In_981,In_906);
xnor U643 (N_643,In_275,In_749);
nand U644 (N_644,In_896,In_213);
and U645 (N_645,In_155,In_783);
nand U646 (N_646,In_871,In_319);
nand U647 (N_647,In_498,In_378);
or U648 (N_648,In_210,In_192);
or U649 (N_649,In_695,In_980);
or U650 (N_650,In_310,In_170);
nand U651 (N_651,In_795,In_354);
xor U652 (N_652,In_626,In_51);
and U653 (N_653,In_262,In_570);
nand U654 (N_654,In_117,In_102);
or U655 (N_655,In_78,In_909);
or U656 (N_656,In_434,In_69);
xor U657 (N_657,In_728,In_37);
or U658 (N_658,In_827,In_816);
xor U659 (N_659,In_607,In_878);
xor U660 (N_660,In_748,In_111);
nor U661 (N_661,In_87,In_859);
nand U662 (N_662,In_373,In_601);
or U663 (N_663,In_455,In_300);
and U664 (N_664,In_525,In_328);
or U665 (N_665,In_916,In_876);
nor U666 (N_666,In_550,In_113);
or U667 (N_667,In_819,In_519);
or U668 (N_668,In_697,In_134);
nand U669 (N_669,In_857,In_776);
nor U670 (N_670,In_169,In_76);
nand U671 (N_671,In_582,In_174);
nand U672 (N_672,In_868,In_713);
nor U673 (N_673,In_567,In_356);
and U674 (N_674,In_814,In_129);
nor U675 (N_675,In_808,In_473);
and U676 (N_676,In_456,In_746);
nor U677 (N_677,In_684,In_154);
nand U678 (N_678,In_596,In_101);
nand U679 (N_679,In_317,In_14);
or U680 (N_680,In_691,In_303);
or U681 (N_681,In_181,In_555);
nand U682 (N_682,In_678,In_760);
nand U683 (N_683,In_847,In_327);
or U684 (N_684,In_996,In_871);
nand U685 (N_685,In_402,In_302);
and U686 (N_686,In_968,In_511);
or U687 (N_687,In_124,In_826);
or U688 (N_688,In_430,In_164);
or U689 (N_689,In_789,In_69);
nand U690 (N_690,In_95,In_236);
and U691 (N_691,In_976,In_918);
or U692 (N_692,In_238,In_992);
xnor U693 (N_693,In_478,In_660);
or U694 (N_694,In_587,In_368);
nand U695 (N_695,In_13,In_919);
nand U696 (N_696,In_540,In_895);
xor U697 (N_697,In_977,In_561);
nor U698 (N_698,In_317,In_612);
and U699 (N_699,In_945,In_991);
and U700 (N_700,In_906,In_300);
and U701 (N_701,In_552,In_172);
nor U702 (N_702,In_295,In_418);
and U703 (N_703,In_866,In_659);
and U704 (N_704,In_359,In_265);
or U705 (N_705,In_999,In_618);
or U706 (N_706,In_203,In_869);
nor U707 (N_707,In_119,In_347);
or U708 (N_708,In_91,In_133);
nor U709 (N_709,In_855,In_44);
or U710 (N_710,In_994,In_71);
nand U711 (N_711,In_916,In_80);
nor U712 (N_712,In_397,In_259);
xor U713 (N_713,In_873,In_667);
nand U714 (N_714,In_830,In_212);
nand U715 (N_715,In_457,In_451);
nor U716 (N_716,In_135,In_158);
xnor U717 (N_717,In_728,In_268);
nand U718 (N_718,In_368,In_656);
or U719 (N_719,In_177,In_655);
nand U720 (N_720,In_107,In_825);
and U721 (N_721,In_792,In_912);
or U722 (N_722,In_345,In_910);
nor U723 (N_723,In_282,In_529);
and U724 (N_724,In_467,In_142);
or U725 (N_725,In_24,In_279);
nand U726 (N_726,In_153,In_124);
or U727 (N_727,In_466,In_323);
nor U728 (N_728,In_944,In_191);
or U729 (N_729,In_769,In_727);
and U730 (N_730,In_653,In_813);
xnor U731 (N_731,In_129,In_355);
nor U732 (N_732,In_317,In_912);
or U733 (N_733,In_439,In_854);
nor U734 (N_734,In_490,In_445);
nor U735 (N_735,In_33,In_676);
nor U736 (N_736,In_84,In_932);
xnor U737 (N_737,In_511,In_709);
nor U738 (N_738,In_389,In_129);
nand U739 (N_739,In_319,In_165);
nor U740 (N_740,In_938,In_247);
xor U741 (N_741,In_691,In_37);
xnor U742 (N_742,In_779,In_787);
xnor U743 (N_743,In_993,In_559);
nand U744 (N_744,In_143,In_665);
and U745 (N_745,In_707,In_300);
and U746 (N_746,In_760,In_637);
or U747 (N_747,In_892,In_133);
nand U748 (N_748,In_426,In_881);
xor U749 (N_749,In_535,In_398);
nand U750 (N_750,In_618,In_904);
nand U751 (N_751,In_550,In_666);
or U752 (N_752,In_344,In_599);
nor U753 (N_753,In_140,In_525);
and U754 (N_754,In_195,In_168);
nor U755 (N_755,In_315,In_1);
nor U756 (N_756,In_812,In_538);
and U757 (N_757,In_787,In_403);
nor U758 (N_758,In_835,In_327);
and U759 (N_759,In_51,In_242);
nor U760 (N_760,In_461,In_505);
nor U761 (N_761,In_471,In_247);
and U762 (N_762,In_600,In_140);
nand U763 (N_763,In_902,In_368);
nand U764 (N_764,In_300,In_457);
or U765 (N_765,In_498,In_402);
nand U766 (N_766,In_326,In_351);
and U767 (N_767,In_304,In_705);
xnor U768 (N_768,In_780,In_96);
nor U769 (N_769,In_739,In_988);
and U770 (N_770,In_39,In_180);
and U771 (N_771,In_171,In_878);
and U772 (N_772,In_208,In_232);
or U773 (N_773,In_14,In_80);
or U774 (N_774,In_234,In_849);
or U775 (N_775,In_48,In_674);
xnor U776 (N_776,In_134,In_635);
and U777 (N_777,In_737,In_408);
xnor U778 (N_778,In_935,In_956);
and U779 (N_779,In_373,In_758);
nor U780 (N_780,In_92,In_593);
xor U781 (N_781,In_128,In_170);
or U782 (N_782,In_293,In_653);
and U783 (N_783,In_966,In_840);
nor U784 (N_784,In_100,In_368);
nor U785 (N_785,In_25,In_968);
xnor U786 (N_786,In_659,In_195);
or U787 (N_787,In_834,In_162);
nor U788 (N_788,In_538,In_621);
xor U789 (N_789,In_582,In_362);
or U790 (N_790,In_75,In_244);
or U791 (N_791,In_967,In_205);
xor U792 (N_792,In_958,In_196);
and U793 (N_793,In_522,In_833);
xnor U794 (N_794,In_632,In_862);
or U795 (N_795,In_987,In_291);
and U796 (N_796,In_635,In_493);
nand U797 (N_797,In_596,In_38);
nor U798 (N_798,In_157,In_40);
and U799 (N_799,In_611,In_246);
and U800 (N_800,In_187,In_727);
and U801 (N_801,In_16,In_114);
nand U802 (N_802,In_219,In_427);
nor U803 (N_803,In_676,In_468);
nand U804 (N_804,In_84,In_616);
nor U805 (N_805,In_68,In_52);
nor U806 (N_806,In_608,In_171);
nand U807 (N_807,In_167,In_254);
nor U808 (N_808,In_799,In_639);
xnor U809 (N_809,In_668,In_578);
or U810 (N_810,In_622,In_234);
or U811 (N_811,In_488,In_541);
xor U812 (N_812,In_253,In_168);
or U813 (N_813,In_847,In_602);
or U814 (N_814,In_905,In_728);
or U815 (N_815,In_283,In_226);
and U816 (N_816,In_278,In_977);
or U817 (N_817,In_22,In_938);
nor U818 (N_818,In_154,In_339);
xor U819 (N_819,In_721,In_889);
nor U820 (N_820,In_235,In_470);
nand U821 (N_821,In_90,In_819);
nor U822 (N_822,In_205,In_424);
nor U823 (N_823,In_783,In_914);
nor U824 (N_824,In_126,In_903);
nand U825 (N_825,In_636,In_647);
nand U826 (N_826,In_788,In_831);
nand U827 (N_827,In_570,In_76);
and U828 (N_828,In_570,In_37);
or U829 (N_829,In_895,In_977);
xor U830 (N_830,In_245,In_600);
and U831 (N_831,In_888,In_320);
nor U832 (N_832,In_570,In_887);
and U833 (N_833,In_674,In_569);
and U834 (N_834,In_894,In_386);
or U835 (N_835,In_117,In_141);
nand U836 (N_836,In_291,In_534);
nor U837 (N_837,In_309,In_952);
nand U838 (N_838,In_252,In_60);
or U839 (N_839,In_273,In_311);
or U840 (N_840,In_155,In_580);
and U841 (N_841,In_897,In_650);
and U842 (N_842,In_467,In_979);
nor U843 (N_843,In_38,In_661);
xnor U844 (N_844,In_637,In_486);
xor U845 (N_845,In_79,In_765);
xor U846 (N_846,In_200,In_801);
xor U847 (N_847,In_556,In_144);
and U848 (N_848,In_871,In_116);
nor U849 (N_849,In_340,In_564);
or U850 (N_850,In_856,In_359);
xor U851 (N_851,In_649,In_574);
and U852 (N_852,In_796,In_437);
xnor U853 (N_853,In_207,In_791);
xnor U854 (N_854,In_717,In_470);
nand U855 (N_855,In_457,In_39);
nor U856 (N_856,In_537,In_559);
and U857 (N_857,In_935,In_443);
nor U858 (N_858,In_358,In_853);
nor U859 (N_859,In_411,In_557);
nor U860 (N_860,In_330,In_743);
or U861 (N_861,In_282,In_547);
and U862 (N_862,In_100,In_5);
or U863 (N_863,In_655,In_656);
or U864 (N_864,In_627,In_110);
or U865 (N_865,In_2,In_783);
nand U866 (N_866,In_121,In_198);
nand U867 (N_867,In_789,In_2);
nor U868 (N_868,In_470,In_821);
xnor U869 (N_869,In_742,In_272);
or U870 (N_870,In_679,In_548);
or U871 (N_871,In_961,In_753);
nand U872 (N_872,In_946,In_939);
and U873 (N_873,In_358,In_186);
xnor U874 (N_874,In_722,In_698);
nand U875 (N_875,In_906,In_658);
or U876 (N_876,In_681,In_887);
nor U877 (N_877,In_412,In_471);
xor U878 (N_878,In_563,In_174);
xor U879 (N_879,In_155,In_320);
nor U880 (N_880,In_373,In_145);
nand U881 (N_881,In_558,In_768);
nand U882 (N_882,In_797,In_375);
xnor U883 (N_883,In_903,In_723);
and U884 (N_884,In_867,In_335);
and U885 (N_885,In_815,In_247);
nor U886 (N_886,In_533,In_970);
nand U887 (N_887,In_77,In_672);
nor U888 (N_888,In_686,In_314);
xnor U889 (N_889,In_719,In_705);
xor U890 (N_890,In_712,In_925);
nand U891 (N_891,In_389,In_623);
and U892 (N_892,In_474,In_719);
or U893 (N_893,In_558,In_744);
nor U894 (N_894,In_251,In_838);
and U895 (N_895,In_346,In_531);
and U896 (N_896,In_423,In_847);
or U897 (N_897,In_232,In_644);
nor U898 (N_898,In_480,In_368);
nand U899 (N_899,In_670,In_499);
or U900 (N_900,In_525,In_527);
and U901 (N_901,In_370,In_672);
nor U902 (N_902,In_911,In_943);
xor U903 (N_903,In_497,In_319);
and U904 (N_904,In_337,In_447);
or U905 (N_905,In_578,In_537);
and U906 (N_906,In_497,In_589);
and U907 (N_907,In_155,In_403);
and U908 (N_908,In_101,In_831);
or U909 (N_909,In_352,In_551);
or U910 (N_910,In_930,In_722);
nor U911 (N_911,In_697,In_140);
or U912 (N_912,In_241,In_709);
and U913 (N_913,In_549,In_522);
or U914 (N_914,In_95,In_834);
and U915 (N_915,In_340,In_397);
nor U916 (N_916,In_561,In_55);
or U917 (N_917,In_790,In_945);
nor U918 (N_918,In_32,In_651);
nand U919 (N_919,In_343,In_437);
xor U920 (N_920,In_18,In_456);
or U921 (N_921,In_822,In_306);
nand U922 (N_922,In_754,In_653);
nor U923 (N_923,In_330,In_25);
nand U924 (N_924,In_646,In_136);
and U925 (N_925,In_757,In_338);
nor U926 (N_926,In_478,In_159);
and U927 (N_927,In_620,In_20);
and U928 (N_928,In_80,In_62);
or U929 (N_929,In_40,In_371);
xor U930 (N_930,In_86,In_241);
nor U931 (N_931,In_380,In_364);
nor U932 (N_932,In_791,In_715);
nor U933 (N_933,In_183,In_56);
and U934 (N_934,In_722,In_412);
nand U935 (N_935,In_516,In_544);
or U936 (N_936,In_640,In_835);
nand U937 (N_937,In_630,In_176);
xor U938 (N_938,In_857,In_129);
or U939 (N_939,In_238,In_550);
or U940 (N_940,In_152,In_348);
or U941 (N_941,In_599,In_936);
nand U942 (N_942,In_348,In_138);
and U943 (N_943,In_112,In_870);
and U944 (N_944,In_102,In_655);
or U945 (N_945,In_50,In_445);
nor U946 (N_946,In_554,In_533);
nand U947 (N_947,In_10,In_747);
or U948 (N_948,In_241,In_187);
and U949 (N_949,In_818,In_329);
and U950 (N_950,In_105,In_257);
nor U951 (N_951,In_12,In_448);
nor U952 (N_952,In_233,In_261);
and U953 (N_953,In_646,In_823);
nor U954 (N_954,In_993,In_225);
nand U955 (N_955,In_489,In_845);
nand U956 (N_956,In_883,In_692);
nand U957 (N_957,In_914,In_986);
or U958 (N_958,In_106,In_707);
nand U959 (N_959,In_996,In_59);
and U960 (N_960,In_941,In_936);
and U961 (N_961,In_473,In_1);
and U962 (N_962,In_862,In_727);
and U963 (N_963,In_751,In_663);
and U964 (N_964,In_115,In_178);
nor U965 (N_965,In_761,In_303);
nand U966 (N_966,In_309,In_321);
nor U967 (N_967,In_459,In_181);
and U968 (N_968,In_91,In_431);
and U969 (N_969,In_758,In_99);
and U970 (N_970,In_475,In_571);
nor U971 (N_971,In_258,In_168);
or U972 (N_972,In_486,In_549);
or U973 (N_973,In_435,In_820);
and U974 (N_974,In_359,In_666);
nand U975 (N_975,In_770,In_153);
or U976 (N_976,In_884,In_627);
or U977 (N_977,In_979,In_348);
and U978 (N_978,In_66,In_913);
and U979 (N_979,In_532,In_357);
nand U980 (N_980,In_128,In_587);
nor U981 (N_981,In_355,In_483);
or U982 (N_982,In_18,In_431);
nand U983 (N_983,In_912,In_427);
and U984 (N_984,In_61,In_37);
nand U985 (N_985,In_328,In_240);
nand U986 (N_986,In_708,In_261);
nand U987 (N_987,In_590,In_857);
nor U988 (N_988,In_854,In_815);
xnor U989 (N_989,In_776,In_101);
or U990 (N_990,In_684,In_157);
and U991 (N_991,In_951,In_629);
xor U992 (N_992,In_20,In_939);
xor U993 (N_993,In_147,In_709);
xor U994 (N_994,In_582,In_741);
nand U995 (N_995,In_716,In_813);
or U996 (N_996,In_622,In_389);
nand U997 (N_997,In_106,In_475);
nand U998 (N_998,In_505,In_630);
and U999 (N_999,In_639,In_337);
or U1000 (N_1000,In_91,In_650);
xnor U1001 (N_1001,In_448,In_390);
and U1002 (N_1002,In_476,In_431);
and U1003 (N_1003,In_494,In_475);
and U1004 (N_1004,In_872,In_464);
and U1005 (N_1005,In_756,In_240);
or U1006 (N_1006,In_822,In_134);
and U1007 (N_1007,In_349,In_747);
nor U1008 (N_1008,In_814,In_686);
nand U1009 (N_1009,In_961,In_368);
nor U1010 (N_1010,In_909,In_398);
xnor U1011 (N_1011,In_448,In_315);
or U1012 (N_1012,In_862,In_989);
nor U1013 (N_1013,In_227,In_79);
xnor U1014 (N_1014,In_243,In_957);
and U1015 (N_1015,In_166,In_673);
and U1016 (N_1016,In_974,In_766);
nand U1017 (N_1017,In_279,In_580);
xnor U1018 (N_1018,In_833,In_339);
or U1019 (N_1019,In_704,In_316);
xor U1020 (N_1020,In_570,In_460);
xor U1021 (N_1021,In_282,In_953);
xor U1022 (N_1022,In_571,In_980);
nand U1023 (N_1023,In_100,In_968);
xnor U1024 (N_1024,In_306,In_333);
nor U1025 (N_1025,In_580,In_748);
and U1026 (N_1026,In_175,In_422);
xor U1027 (N_1027,In_694,In_682);
xor U1028 (N_1028,In_76,In_761);
nor U1029 (N_1029,In_573,In_827);
nand U1030 (N_1030,In_997,In_536);
or U1031 (N_1031,In_952,In_6);
nor U1032 (N_1032,In_990,In_160);
nor U1033 (N_1033,In_475,In_841);
and U1034 (N_1034,In_49,In_716);
or U1035 (N_1035,In_636,In_658);
or U1036 (N_1036,In_278,In_223);
nand U1037 (N_1037,In_82,In_896);
nand U1038 (N_1038,In_658,In_397);
xnor U1039 (N_1039,In_119,In_28);
nand U1040 (N_1040,In_78,In_664);
or U1041 (N_1041,In_278,In_532);
and U1042 (N_1042,In_74,In_494);
and U1043 (N_1043,In_97,In_544);
xnor U1044 (N_1044,In_973,In_784);
xnor U1045 (N_1045,In_337,In_997);
nor U1046 (N_1046,In_296,In_888);
xor U1047 (N_1047,In_745,In_46);
or U1048 (N_1048,In_539,In_153);
nor U1049 (N_1049,In_888,In_252);
or U1050 (N_1050,In_681,In_825);
xor U1051 (N_1051,In_219,In_124);
nor U1052 (N_1052,In_109,In_657);
or U1053 (N_1053,In_642,In_794);
nor U1054 (N_1054,In_987,In_972);
xor U1055 (N_1055,In_5,In_795);
or U1056 (N_1056,In_240,In_146);
and U1057 (N_1057,In_49,In_146);
and U1058 (N_1058,In_906,In_564);
nand U1059 (N_1059,In_947,In_853);
nand U1060 (N_1060,In_338,In_903);
nand U1061 (N_1061,In_485,In_727);
and U1062 (N_1062,In_49,In_927);
nor U1063 (N_1063,In_41,In_890);
xnor U1064 (N_1064,In_608,In_888);
or U1065 (N_1065,In_209,In_406);
or U1066 (N_1066,In_516,In_730);
nor U1067 (N_1067,In_519,In_64);
nand U1068 (N_1068,In_649,In_902);
nand U1069 (N_1069,In_774,In_694);
nor U1070 (N_1070,In_668,In_133);
nor U1071 (N_1071,In_91,In_270);
nor U1072 (N_1072,In_752,In_754);
and U1073 (N_1073,In_508,In_369);
nor U1074 (N_1074,In_50,In_340);
xnor U1075 (N_1075,In_95,In_564);
nand U1076 (N_1076,In_539,In_336);
xnor U1077 (N_1077,In_582,In_933);
nor U1078 (N_1078,In_368,In_588);
nand U1079 (N_1079,In_905,In_520);
or U1080 (N_1080,In_691,In_463);
and U1081 (N_1081,In_862,In_720);
and U1082 (N_1082,In_515,In_966);
nand U1083 (N_1083,In_189,In_83);
nor U1084 (N_1084,In_156,In_337);
and U1085 (N_1085,In_961,In_121);
or U1086 (N_1086,In_154,In_349);
xor U1087 (N_1087,In_137,In_60);
xor U1088 (N_1088,In_542,In_829);
and U1089 (N_1089,In_24,In_441);
or U1090 (N_1090,In_568,In_10);
nand U1091 (N_1091,In_886,In_342);
nand U1092 (N_1092,In_601,In_589);
xor U1093 (N_1093,In_457,In_733);
nand U1094 (N_1094,In_61,In_295);
and U1095 (N_1095,In_919,In_413);
xnor U1096 (N_1096,In_227,In_808);
or U1097 (N_1097,In_559,In_780);
or U1098 (N_1098,In_179,In_274);
and U1099 (N_1099,In_156,In_696);
and U1100 (N_1100,In_529,In_164);
nand U1101 (N_1101,In_669,In_381);
xnor U1102 (N_1102,In_283,In_382);
or U1103 (N_1103,In_308,In_470);
nor U1104 (N_1104,In_517,In_764);
nor U1105 (N_1105,In_694,In_212);
and U1106 (N_1106,In_326,In_937);
nor U1107 (N_1107,In_471,In_517);
nand U1108 (N_1108,In_467,In_534);
nand U1109 (N_1109,In_194,In_780);
and U1110 (N_1110,In_505,In_134);
nor U1111 (N_1111,In_585,In_401);
or U1112 (N_1112,In_434,In_100);
nand U1113 (N_1113,In_700,In_925);
and U1114 (N_1114,In_892,In_129);
nor U1115 (N_1115,In_742,In_25);
nand U1116 (N_1116,In_804,In_935);
nor U1117 (N_1117,In_478,In_101);
and U1118 (N_1118,In_243,In_368);
or U1119 (N_1119,In_175,In_272);
nand U1120 (N_1120,In_659,In_41);
xor U1121 (N_1121,In_460,In_986);
and U1122 (N_1122,In_848,In_723);
or U1123 (N_1123,In_628,In_129);
or U1124 (N_1124,In_561,In_646);
xnor U1125 (N_1125,In_195,In_692);
and U1126 (N_1126,In_412,In_794);
and U1127 (N_1127,In_63,In_642);
nand U1128 (N_1128,In_521,In_568);
nor U1129 (N_1129,In_466,In_455);
nand U1130 (N_1130,In_23,In_454);
or U1131 (N_1131,In_510,In_632);
xor U1132 (N_1132,In_168,In_230);
xor U1133 (N_1133,In_101,In_784);
nand U1134 (N_1134,In_876,In_177);
nor U1135 (N_1135,In_780,In_506);
and U1136 (N_1136,In_635,In_72);
nand U1137 (N_1137,In_675,In_976);
xnor U1138 (N_1138,In_380,In_833);
nor U1139 (N_1139,In_124,In_678);
xnor U1140 (N_1140,In_416,In_175);
nor U1141 (N_1141,In_420,In_844);
and U1142 (N_1142,In_925,In_446);
nor U1143 (N_1143,In_14,In_562);
xor U1144 (N_1144,In_650,In_572);
xnor U1145 (N_1145,In_391,In_915);
and U1146 (N_1146,In_127,In_976);
nand U1147 (N_1147,In_685,In_523);
nor U1148 (N_1148,In_985,In_232);
xnor U1149 (N_1149,In_718,In_618);
or U1150 (N_1150,In_740,In_630);
nand U1151 (N_1151,In_533,In_335);
xnor U1152 (N_1152,In_671,In_542);
nor U1153 (N_1153,In_324,In_495);
and U1154 (N_1154,In_726,In_631);
nor U1155 (N_1155,In_207,In_67);
xor U1156 (N_1156,In_349,In_831);
nand U1157 (N_1157,In_377,In_704);
or U1158 (N_1158,In_932,In_815);
and U1159 (N_1159,In_220,In_496);
xor U1160 (N_1160,In_820,In_13);
or U1161 (N_1161,In_459,In_624);
nand U1162 (N_1162,In_582,In_230);
and U1163 (N_1163,In_351,In_968);
or U1164 (N_1164,In_855,In_473);
nor U1165 (N_1165,In_299,In_29);
nand U1166 (N_1166,In_526,In_575);
nor U1167 (N_1167,In_841,In_126);
nand U1168 (N_1168,In_583,In_955);
xnor U1169 (N_1169,In_655,In_316);
nor U1170 (N_1170,In_982,In_782);
or U1171 (N_1171,In_819,In_648);
or U1172 (N_1172,In_104,In_686);
nor U1173 (N_1173,In_845,In_777);
and U1174 (N_1174,In_808,In_597);
nor U1175 (N_1175,In_49,In_108);
or U1176 (N_1176,In_445,In_956);
xnor U1177 (N_1177,In_629,In_51);
and U1178 (N_1178,In_897,In_810);
nand U1179 (N_1179,In_454,In_663);
xnor U1180 (N_1180,In_381,In_445);
nand U1181 (N_1181,In_988,In_770);
and U1182 (N_1182,In_787,In_559);
nor U1183 (N_1183,In_629,In_229);
nand U1184 (N_1184,In_187,In_980);
and U1185 (N_1185,In_773,In_431);
xnor U1186 (N_1186,In_424,In_41);
nand U1187 (N_1187,In_591,In_985);
xnor U1188 (N_1188,In_12,In_65);
xor U1189 (N_1189,In_648,In_592);
nand U1190 (N_1190,In_441,In_263);
nor U1191 (N_1191,In_296,In_690);
and U1192 (N_1192,In_557,In_447);
or U1193 (N_1193,In_494,In_309);
or U1194 (N_1194,In_46,In_974);
nand U1195 (N_1195,In_165,In_197);
nor U1196 (N_1196,In_994,In_346);
or U1197 (N_1197,In_158,In_968);
or U1198 (N_1198,In_510,In_298);
xor U1199 (N_1199,In_32,In_417);
or U1200 (N_1200,In_736,In_567);
xnor U1201 (N_1201,In_740,In_779);
xor U1202 (N_1202,In_540,In_307);
and U1203 (N_1203,In_492,In_846);
nor U1204 (N_1204,In_878,In_723);
xnor U1205 (N_1205,In_943,In_482);
xnor U1206 (N_1206,In_286,In_507);
xor U1207 (N_1207,In_288,In_194);
or U1208 (N_1208,In_406,In_175);
and U1209 (N_1209,In_843,In_258);
nand U1210 (N_1210,In_865,In_258);
or U1211 (N_1211,In_855,In_152);
xor U1212 (N_1212,In_811,In_581);
and U1213 (N_1213,In_974,In_708);
nor U1214 (N_1214,In_677,In_401);
nand U1215 (N_1215,In_58,In_671);
or U1216 (N_1216,In_203,In_158);
nor U1217 (N_1217,In_537,In_258);
nand U1218 (N_1218,In_412,In_250);
nand U1219 (N_1219,In_990,In_467);
nor U1220 (N_1220,In_811,In_847);
nor U1221 (N_1221,In_897,In_300);
xor U1222 (N_1222,In_905,In_206);
and U1223 (N_1223,In_765,In_391);
and U1224 (N_1224,In_985,In_728);
nor U1225 (N_1225,In_911,In_128);
xnor U1226 (N_1226,In_384,In_627);
nand U1227 (N_1227,In_808,In_983);
nand U1228 (N_1228,In_867,In_812);
nor U1229 (N_1229,In_97,In_15);
nor U1230 (N_1230,In_197,In_432);
nor U1231 (N_1231,In_853,In_752);
nand U1232 (N_1232,In_872,In_291);
nand U1233 (N_1233,In_248,In_580);
nor U1234 (N_1234,In_160,In_315);
xnor U1235 (N_1235,In_624,In_831);
nand U1236 (N_1236,In_438,In_297);
or U1237 (N_1237,In_421,In_783);
nor U1238 (N_1238,In_879,In_756);
nor U1239 (N_1239,In_708,In_276);
nor U1240 (N_1240,In_142,In_938);
and U1241 (N_1241,In_734,In_791);
xnor U1242 (N_1242,In_938,In_202);
or U1243 (N_1243,In_37,In_551);
and U1244 (N_1244,In_415,In_241);
nor U1245 (N_1245,In_268,In_197);
and U1246 (N_1246,In_93,In_290);
or U1247 (N_1247,In_302,In_365);
or U1248 (N_1248,In_144,In_743);
and U1249 (N_1249,In_443,In_416);
nor U1250 (N_1250,In_462,In_456);
nor U1251 (N_1251,In_655,In_325);
nand U1252 (N_1252,In_376,In_319);
xor U1253 (N_1253,In_551,In_901);
nand U1254 (N_1254,In_629,In_269);
and U1255 (N_1255,In_45,In_824);
nor U1256 (N_1256,In_316,In_345);
or U1257 (N_1257,In_844,In_361);
nor U1258 (N_1258,In_952,In_12);
nor U1259 (N_1259,In_118,In_434);
nor U1260 (N_1260,In_439,In_888);
xor U1261 (N_1261,In_524,In_475);
or U1262 (N_1262,In_36,In_843);
or U1263 (N_1263,In_276,In_824);
or U1264 (N_1264,In_191,In_158);
or U1265 (N_1265,In_566,In_183);
nand U1266 (N_1266,In_609,In_447);
and U1267 (N_1267,In_179,In_639);
xor U1268 (N_1268,In_831,In_752);
and U1269 (N_1269,In_330,In_376);
nor U1270 (N_1270,In_322,In_549);
and U1271 (N_1271,In_460,In_211);
or U1272 (N_1272,In_821,In_751);
nand U1273 (N_1273,In_124,In_549);
or U1274 (N_1274,In_132,In_88);
nand U1275 (N_1275,In_722,In_518);
xor U1276 (N_1276,In_107,In_991);
nor U1277 (N_1277,In_324,In_643);
and U1278 (N_1278,In_376,In_844);
nor U1279 (N_1279,In_428,In_3);
or U1280 (N_1280,In_718,In_178);
nor U1281 (N_1281,In_755,In_613);
xor U1282 (N_1282,In_462,In_748);
xnor U1283 (N_1283,In_7,In_951);
and U1284 (N_1284,In_260,In_338);
xnor U1285 (N_1285,In_323,In_464);
nand U1286 (N_1286,In_625,In_384);
nand U1287 (N_1287,In_977,In_346);
and U1288 (N_1288,In_0,In_908);
xor U1289 (N_1289,In_948,In_135);
nor U1290 (N_1290,In_16,In_225);
and U1291 (N_1291,In_777,In_570);
xnor U1292 (N_1292,In_240,In_377);
and U1293 (N_1293,In_213,In_205);
or U1294 (N_1294,In_869,In_92);
xor U1295 (N_1295,In_543,In_384);
xor U1296 (N_1296,In_533,In_854);
nor U1297 (N_1297,In_729,In_19);
and U1298 (N_1298,In_51,In_25);
nand U1299 (N_1299,In_554,In_580);
nand U1300 (N_1300,In_815,In_57);
and U1301 (N_1301,In_666,In_995);
xnor U1302 (N_1302,In_423,In_326);
or U1303 (N_1303,In_89,In_288);
nand U1304 (N_1304,In_774,In_751);
or U1305 (N_1305,In_198,In_439);
xnor U1306 (N_1306,In_373,In_384);
xnor U1307 (N_1307,In_313,In_3);
nand U1308 (N_1308,In_792,In_263);
nor U1309 (N_1309,In_476,In_481);
and U1310 (N_1310,In_519,In_648);
nor U1311 (N_1311,In_821,In_515);
nand U1312 (N_1312,In_73,In_546);
nor U1313 (N_1313,In_473,In_186);
or U1314 (N_1314,In_264,In_566);
xnor U1315 (N_1315,In_29,In_351);
nand U1316 (N_1316,In_67,In_545);
nor U1317 (N_1317,In_644,In_950);
xnor U1318 (N_1318,In_526,In_783);
nand U1319 (N_1319,In_111,In_990);
and U1320 (N_1320,In_360,In_336);
nand U1321 (N_1321,In_971,In_539);
xnor U1322 (N_1322,In_61,In_51);
nand U1323 (N_1323,In_835,In_123);
xor U1324 (N_1324,In_656,In_325);
xnor U1325 (N_1325,In_803,In_277);
nand U1326 (N_1326,In_326,In_49);
xor U1327 (N_1327,In_122,In_76);
nand U1328 (N_1328,In_736,In_207);
nand U1329 (N_1329,In_207,In_140);
nor U1330 (N_1330,In_688,In_702);
or U1331 (N_1331,In_974,In_727);
nand U1332 (N_1332,In_918,In_638);
nor U1333 (N_1333,In_545,In_924);
and U1334 (N_1334,In_77,In_607);
nand U1335 (N_1335,In_512,In_484);
and U1336 (N_1336,In_120,In_635);
nand U1337 (N_1337,In_779,In_271);
xor U1338 (N_1338,In_518,In_800);
xor U1339 (N_1339,In_22,In_413);
and U1340 (N_1340,In_897,In_233);
xnor U1341 (N_1341,In_839,In_948);
nor U1342 (N_1342,In_964,In_677);
nor U1343 (N_1343,In_614,In_727);
and U1344 (N_1344,In_564,In_255);
nand U1345 (N_1345,In_316,In_996);
xor U1346 (N_1346,In_986,In_707);
nor U1347 (N_1347,In_511,In_294);
or U1348 (N_1348,In_169,In_519);
and U1349 (N_1349,In_892,In_42);
nor U1350 (N_1350,In_457,In_540);
or U1351 (N_1351,In_386,In_259);
nor U1352 (N_1352,In_501,In_335);
and U1353 (N_1353,In_186,In_903);
nor U1354 (N_1354,In_295,In_73);
nand U1355 (N_1355,In_961,In_273);
nor U1356 (N_1356,In_865,In_941);
nor U1357 (N_1357,In_699,In_192);
nand U1358 (N_1358,In_361,In_601);
nor U1359 (N_1359,In_402,In_624);
and U1360 (N_1360,In_720,In_599);
nor U1361 (N_1361,In_780,In_801);
and U1362 (N_1362,In_338,In_367);
xor U1363 (N_1363,In_833,In_536);
nand U1364 (N_1364,In_949,In_400);
and U1365 (N_1365,In_346,In_216);
nor U1366 (N_1366,In_683,In_30);
or U1367 (N_1367,In_360,In_907);
nand U1368 (N_1368,In_342,In_526);
xor U1369 (N_1369,In_60,In_539);
xnor U1370 (N_1370,In_774,In_614);
nor U1371 (N_1371,In_846,In_197);
nand U1372 (N_1372,In_765,In_964);
xnor U1373 (N_1373,In_996,In_199);
nor U1374 (N_1374,In_375,In_734);
xor U1375 (N_1375,In_390,In_361);
xnor U1376 (N_1376,In_469,In_705);
xor U1377 (N_1377,In_708,In_134);
and U1378 (N_1378,In_334,In_110);
xnor U1379 (N_1379,In_81,In_530);
xnor U1380 (N_1380,In_864,In_711);
nor U1381 (N_1381,In_420,In_237);
nor U1382 (N_1382,In_945,In_63);
xnor U1383 (N_1383,In_181,In_460);
nand U1384 (N_1384,In_798,In_789);
nor U1385 (N_1385,In_8,In_542);
or U1386 (N_1386,In_893,In_277);
nor U1387 (N_1387,In_725,In_260);
xnor U1388 (N_1388,In_598,In_643);
nor U1389 (N_1389,In_386,In_297);
nand U1390 (N_1390,In_577,In_457);
or U1391 (N_1391,In_780,In_620);
and U1392 (N_1392,In_40,In_608);
nand U1393 (N_1393,In_713,In_574);
xnor U1394 (N_1394,In_826,In_868);
xnor U1395 (N_1395,In_938,In_144);
nor U1396 (N_1396,In_818,In_207);
or U1397 (N_1397,In_821,In_343);
nor U1398 (N_1398,In_850,In_466);
and U1399 (N_1399,In_692,In_355);
nand U1400 (N_1400,In_986,In_734);
nor U1401 (N_1401,In_529,In_552);
nand U1402 (N_1402,In_646,In_61);
or U1403 (N_1403,In_626,In_366);
or U1404 (N_1404,In_917,In_351);
or U1405 (N_1405,In_266,In_250);
nand U1406 (N_1406,In_274,In_86);
or U1407 (N_1407,In_115,In_567);
xor U1408 (N_1408,In_720,In_528);
or U1409 (N_1409,In_506,In_909);
nand U1410 (N_1410,In_422,In_359);
nand U1411 (N_1411,In_558,In_539);
nand U1412 (N_1412,In_772,In_533);
xor U1413 (N_1413,In_30,In_147);
xor U1414 (N_1414,In_704,In_25);
xnor U1415 (N_1415,In_367,In_912);
and U1416 (N_1416,In_62,In_778);
nand U1417 (N_1417,In_387,In_786);
xor U1418 (N_1418,In_367,In_376);
and U1419 (N_1419,In_727,In_747);
or U1420 (N_1420,In_443,In_841);
or U1421 (N_1421,In_322,In_368);
and U1422 (N_1422,In_436,In_359);
xnor U1423 (N_1423,In_88,In_166);
nor U1424 (N_1424,In_9,In_251);
nand U1425 (N_1425,In_994,In_203);
nor U1426 (N_1426,In_934,In_565);
xnor U1427 (N_1427,In_911,In_723);
nor U1428 (N_1428,In_793,In_576);
and U1429 (N_1429,In_837,In_62);
or U1430 (N_1430,In_476,In_50);
or U1431 (N_1431,In_236,In_208);
or U1432 (N_1432,In_960,In_399);
nand U1433 (N_1433,In_43,In_206);
and U1434 (N_1434,In_640,In_418);
nand U1435 (N_1435,In_813,In_71);
xor U1436 (N_1436,In_450,In_693);
or U1437 (N_1437,In_556,In_156);
xor U1438 (N_1438,In_161,In_121);
nor U1439 (N_1439,In_679,In_975);
and U1440 (N_1440,In_54,In_737);
and U1441 (N_1441,In_208,In_901);
xor U1442 (N_1442,In_378,In_825);
xor U1443 (N_1443,In_496,In_834);
and U1444 (N_1444,In_231,In_814);
nand U1445 (N_1445,In_392,In_179);
or U1446 (N_1446,In_993,In_946);
nand U1447 (N_1447,In_190,In_523);
or U1448 (N_1448,In_463,In_528);
or U1449 (N_1449,In_778,In_221);
and U1450 (N_1450,In_890,In_1);
or U1451 (N_1451,In_138,In_852);
nand U1452 (N_1452,In_572,In_991);
xor U1453 (N_1453,In_3,In_507);
nor U1454 (N_1454,In_748,In_186);
nand U1455 (N_1455,In_128,In_918);
or U1456 (N_1456,In_796,In_846);
and U1457 (N_1457,In_9,In_105);
nand U1458 (N_1458,In_749,In_244);
or U1459 (N_1459,In_737,In_896);
nand U1460 (N_1460,In_674,In_118);
nor U1461 (N_1461,In_242,In_842);
nand U1462 (N_1462,In_365,In_580);
nand U1463 (N_1463,In_185,In_575);
or U1464 (N_1464,In_683,In_487);
or U1465 (N_1465,In_312,In_495);
xor U1466 (N_1466,In_103,In_4);
or U1467 (N_1467,In_607,In_502);
or U1468 (N_1468,In_849,In_990);
xnor U1469 (N_1469,In_571,In_114);
nor U1470 (N_1470,In_682,In_446);
and U1471 (N_1471,In_573,In_987);
nand U1472 (N_1472,In_214,In_774);
and U1473 (N_1473,In_161,In_37);
xnor U1474 (N_1474,In_87,In_729);
xnor U1475 (N_1475,In_752,In_820);
nor U1476 (N_1476,In_381,In_66);
nor U1477 (N_1477,In_300,In_610);
and U1478 (N_1478,In_944,In_644);
nor U1479 (N_1479,In_665,In_913);
nor U1480 (N_1480,In_469,In_403);
and U1481 (N_1481,In_560,In_273);
xor U1482 (N_1482,In_136,In_927);
or U1483 (N_1483,In_810,In_72);
or U1484 (N_1484,In_795,In_152);
and U1485 (N_1485,In_718,In_986);
and U1486 (N_1486,In_925,In_74);
nor U1487 (N_1487,In_201,In_419);
nand U1488 (N_1488,In_154,In_694);
nand U1489 (N_1489,In_263,In_983);
and U1490 (N_1490,In_755,In_319);
or U1491 (N_1491,In_906,In_809);
nand U1492 (N_1492,In_240,In_496);
nand U1493 (N_1493,In_513,In_164);
xnor U1494 (N_1494,In_614,In_325);
xnor U1495 (N_1495,In_25,In_472);
nand U1496 (N_1496,In_525,In_287);
xnor U1497 (N_1497,In_175,In_21);
nor U1498 (N_1498,In_523,In_825);
nand U1499 (N_1499,In_814,In_317);
nand U1500 (N_1500,In_358,In_674);
and U1501 (N_1501,In_322,In_249);
and U1502 (N_1502,In_552,In_108);
nor U1503 (N_1503,In_626,In_127);
nand U1504 (N_1504,In_369,In_636);
or U1505 (N_1505,In_25,In_47);
nand U1506 (N_1506,In_472,In_635);
or U1507 (N_1507,In_797,In_859);
or U1508 (N_1508,In_969,In_326);
or U1509 (N_1509,In_149,In_839);
xnor U1510 (N_1510,In_545,In_744);
xnor U1511 (N_1511,In_957,In_699);
or U1512 (N_1512,In_807,In_792);
nand U1513 (N_1513,In_461,In_116);
xor U1514 (N_1514,In_271,In_841);
nor U1515 (N_1515,In_263,In_678);
xnor U1516 (N_1516,In_605,In_458);
or U1517 (N_1517,In_92,In_892);
xnor U1518 (N_1518,In_952,In_126);
xor U1519 (N_1519,In_181,In_501);
and U1520 (N_1520,In_976,In_968);
nand U1521 (N_1521,In_596,In_379);
and U1522 (N_1522,In_906,In_634);
or U1523 (N_1523,In_929,In_425);
or U1524 (N_1524,In_722,In_294);
nor U1525 (N_1525,In_653,In_77);
nand U1526 (N_1526,In_755,In_985);
xor U1527 (N_1527,In_626,In_578);
nand U1528 (N_1528,In_240,In_794);
nand U1529 (N_1529,In_852,In_674);
and U1530 (N_1530,In_309,In_41);
nor U1531 (N_1531,In_350,In_479);
nand U1532 (N_1532,In_322,In_723);
nand U1533 (N_1533,In_459,In_489);
nor U1534 (N_1534,In_918,In_919);
or U1535 (N_1535,In_777,In_870);
xnor U1536 (N_1536,In_627,In_885);
and U1537 (N_1537,In_628,In_190);
xor U1538 (N_1538,In_857,In_204);
and U1539 (N_1539,In_301,In_810);
and U1540 (N_1540,In_734,In_966);
nand U1541 (N_1541,In_628,In_917);
and U1542 (N_1542,In_894,In_920);
or U1543 (N_1543,In_321,In_787);
nor U1544 (N_1544,In_733,In_22);
nor U1545 (N_1545,In_19,In_407);
xor U1546 (N_1546,In_512,In_743);
nand U1547 (N_1547,In_337,In_687);
and U1548 (N_1548,In_865,In_492);
nand U1549 (N_1549,In_253,In_266);
and U1550 (N_1550,In_360,In_519);
or U1551 (N_1551,In_586,In_271);
and U1552 (N_1552,In_415,In_866);
or U1553 (N_1553,In_898,In_113);
xnor U1554 (N_1554,In_62,In_817);
nand U1555 (N_1555,In_937,In_348);
or U1556 (N_1556,In_118,In_416);
nand U1557 (N_1557,In_724,In_66);
or U1558 (N_1558,In_177,In_48);
xor U1559 (N_1559,In_266,In_300);
and U1560 (N_1560,In_885,In_688);
nand U1561 (N_1561,In_741,In_658);
xnor U1562 (N_1562,In_306,In_926);
and U1563 (N_1563,In_773,In_847);
and U1564 (N_1564,In_307,In_420);
or U1565 (N_1565,In_319,In_457);
nand U1566 (N_1566,In_300,In_574);
or U1567 (N_1567,In_953,In_667);
or U1568 (N_1568,In_37,In_469);
xor U1569 (N_1569,In_944,In_662);
and U1570 (N_1570,In_94,In_356);
xnor U1571 (N_1571,In_816,In_550);
xnor U1572 (N_1572,In_528,In_982);
and U1573 (N_1573,In_195,In_353);
nor U1574 (N_1574,In_996,In_793);
xor U1575 (N_1575,In_605,In_294);
or U1576 (N_1576,In_363,In_16);
nor U1577 (N_1577,In_964,In_57);
nand U1578 (N_1578,In_359,In_673);
nor U1579 (N_1579,In_642,In_604);
nor U1580 (N_1580,In_819,In_316);
nor U1581 (N_1581,In_664,In_689);
or U1582 (N_1582,In_846,In_189);
and U1583 (N_1583,In_251,In_421);
xor U1584 (N_1584,In_635,In_561);
xnor U1585 (N_1585,In_341,In_418);
or U1586 (N_1586,In_31,In_283);
or U1587 (N_1587,In_82,In_27);
nor U1588 (N_1588,In_713,In_688);
nor U1589 (N_1589,In_599,In_221);
nand U1590 (N_1590,In_233,In_872);
and U1591 (N_1591,In_564,In_581);
or U1592 (N_1592,In_379,In_714);
nor U1593 (N_1593,In_527,In_696);
xor U1594 (N_1594,In_84,In_716);
nor U1595 (N_1595,In_606,In_690);
nand U1596 (N_1596,In_143,In_808);
xor U1597 (N_1597,In_283,In_978);
or U1598 (N_1598,In_829,In_423);
nand U1599 (N_1599,In_355,In_397);
nor U1600 (N_1600,In_464,In_827);
nor U1601 (N_1601,In_993,In_90);
nand U1602 (N_1602,In_624,In_243);
xor U1603 (N_1603,In_956,In_437);
xor U1604 (N_1604,In_451,In_406);
nand U1605 (N_1605,In_762,In_560);
xnor U1606 (N_1606,In_437,In_849);
or U1607 (N_1607,In_586,In_422);
nand U1608 (N_1608,In_89,In_137);
nand U1609 (N_1609,In_857,In_520);
nand U1610 (N_1610,In_287,In_627);
nand U1611 (N_1611,In_643,In_692);
nand U1612 (N_1612,In_745,In_0);
xor U1613 (N_1613,In_72,In_54);
nor U1614 (N_1614,In_439,In_94);
nor U1615 (N_1615,In_82,In_445);
and U1616 (N_1616,In_609,In_785);
nor U1617 (N_1617,In_950,In_12);
and U1618 (N_1618,In_977,In_937);
and U1619 (N_1619,In_540,In_281);
nor U1620 (N_1620,In_220,In_477);
xor U1621 (N_1621,In_549,In_491);
xnor U1622 (N_1622,In_261,In_838);
and U1623 (N_1623,In_720,In_442);
and U1624 (N_1624,In_752,In_509);
or U1625 (N_1625,In_385,In_492);
or U1626 (N_1626,In_409,In_405);
or U1627 (N_1627,In_978,In_950);
xnor U1628 (N_1628,In_436,In_944);
or U1629 (N_1629,In_934,In_650);
or U1630 (N_1630,In_128,In_45);
or U1631 (N_1631,In_187,In_383);
nand U1632 (N_1632,In_253,In_718);
xor U1633 (N_1633,In_940,In_362);
and U1634 (N_1634,In_180,In_226);
nand U1635 (N_1635,In_788,In_265);
or U1636 (N_1636,In_298,In_70);
or U1637 (N_1637,In_911,In_21);
nor U1638 (N_1638,In_540,In_20);
xor U1639 (N_1639,In_845,In_540);
and U1640 (N_1640,In_952,In_279);
nor U1641 (N_1641,In_539,In_572);
nand U1642 (N_1642,In_926,In_240);
or U1643 (N_1643,In_425,In_605);
and U1644 (N_1644,In_163,In_454);
and U1645 (N_1645,In_595,In_861);
and U1646 (N_1646,In_910,In_169);
or U1647 (N_1647,In_396,In_16);
nor U1648 (N_1648,In_33,In_342);
xor U1649 (N_1649,In_248,In_979);
nor U1650 (N_1650,In_801,In_629);
and U1651 (N_1651,In_145,In_711);
xor U1652 (N_1652,In_890,In_970);
nand U1653 (N_1653,In_980,In_343);
nand U1654 (N_1654,In_225,In_949);
nor U1655 (N_1655,In_181,In_450);
xnor U1656 (N_1656,In_495,In_990);
nor U1657 (N_1657,In_8,In_623);
xor U1658 (N_1658,In_714,In_658);
nand U1659 (N_1659,In_707,In_349);
and U1660 (N_1660,In_11,In_653);
and U1661 (N_1661,In_642,In_947);
nor U1662 (N_1662,In_714,In_134);
nor U1663 (N_1663,In_139,In_94);
xor U1664 (N_1664,In_410,In_183);
or U1665 (N_1665,In_806,In_423);
or U1666 (N_1666,In_78,In_543);
and U1667 (N_1667,In_78,In_445);
xor U1668 (N_1668,In_186,In_290);
nor U1669 (N_1669,In_738,In_548);
nand U1670 (N_1670,In_131,In_856);
or U1671 (N_1671,In_431,In_879);
or U1672 (N_1672,In_795,In_330);
nand U1673 (N_1673,In_550,In_181);
nand U1674 (N_1674,In_925,In_550);
or U1675 (N_1675,In_372,In_875);
xnor U1676 (N_1676,In_558,In_509);
nand U1677 (N_1677,In_270,In_509);
nor U1678 (N_1678,In_34,In_123);
nand U1679 (N_1679,In_355,In_898);
xor U1680 (N_1680,In_796,In_898);
nor U1681 (N_1681,In_428,In_39);
nand U1682 (N_1682,In_148,In_766);
and U1683 (N_1683,In_664,In_866);
and U1684 (N_1684,In_436,In_980);
and U1685 (N_1685,In_343,In_843);
and U1686 (N_1686,In_350,In_37);
nand U1687 (N_1687,In_328,In_130);
and U1688 (N_1688,In_323,In_316);
xor U1689 (N_1689,In_764,In_992);
nand U1690 (N_1690,In_60,In_214);
nand U1691 (N_1691,In_473,In_485);
xor U1692 (N_1692,In_110,In_590);
xor U1693 (N_1693,In_318,In_870);
nor U1694 (N_1694,In_529,In_262);
nor U1695 (N_1695,In_318,In_143);
and U1696 (N_1696,In_595,In_702);
xnor U1697 (N_1697,In_597,In_151);
and U1698 (N_1698,In_442,In_139);
xor U1699 (N_1699,In_971,In_494);
nor U1700 (N_1700,In_259,In_550);
xnor U1701 (N_1701,In_943,In_66);
nor U1702 (N_1702,In_222,In_130);
nor U1703 (N_1703,In_307,In_936);
or U1704 (N_1704,In_169,In_422);
nor U1705 (N_1705,In_94,In_887);
or U1706 (N_1706,In_450,In_81);
nand U1707 (N_1707,In_663,In_732);
nor U1708 (N_1708,In_952,In_983);
or U1709 (N_1709,In_373,In_631);
or U1710 (N_1710,In_207,In_108);
or U1711 (N_1711,In_260,In_666);
nor U1712 (N_1712,In_284,In_366);
nor U1713 (N_1713,In_67,In_323);
xor U1714 (N_1714,In_101,In_153);
xnor U1715 (N_1715,In_342,In_319);
or U1716 (N_1716,In_707,In_212);
nor U1717 (N_1717,In_758,In_782);
nor U1718 (N_1718,In_799,In_658);
nand U1719 (N_1719,In_163,In_53);
and U1720 (N_1720,In_337,In_823);
nor U1721 (N_1721,In_1,In_102);
nand U1722 (N_1722,In_894,In_495);
and U1723 (N_1723,In_590,In_863);
nand U1724 (N_1724,In_970,In_884);
nor U1725 (N_1725,In_303,In_901);
nor U1726 (N_1726,In_330,In_352);
or U1727 (N_1727,In_754,In_173);
nand U1728 (N_1728,In_181,In_48);
xor U1729 (N_1729,In_547,In_324);
and U1730 (N_1730,In_707,In_610);
or U1731 (N_1731,In_212,In_340);
and U1732 (N_1732,In_749,In_703);
nor U1733 (N_1733,In_907,In_76);
nand U1734 (N_1734,In_491,In_419);
xnor U1735 (N_1735,In_295,In_252);
nor U1736 (N_1736,In_720,In_324);
nand U1737 (N_1737,In_566,In_887);
or U1738 (N_1738,In_161,In_860);
or U1739 (N_1739,In_722,In_706);
nor U1740 (N_1740,In_480,In_619);
and U1741 (N_1741,In_825,In_850);
nor U1742 (N_1742,In_149,In_521);
nand U1743 (N_1743,In_349,In_908);
nand U1744 (N_1744,In_465,In_927);
or U1745 (N_1745,In_142,In_177);
nand U1746 (N_1746,In_20,In_68);
and U1747 (N_1747,In_182,In_528);
and U1748 (N_1748,In_8,In_831);
nor U1749 (N_1749,In_810,In_764);
xnor U1750 (N_1750,In_30,In_499);
or U1751 (N_1751,In_811,In_290);
or U1752 (N_1752,In_72,In_876);
xor U1753 (N_1753,In_338,In_660);
and U1754 (N_1754,In_664,In_277);
nor U1755 (N_1755,In_620,In_108);
or U1756 (N_1756,In_887,In_446);
nor U1757 (N_1757,In_298,In_477);
xor U1758 (N_1758,In_726,In_641);
nand U1759 (N_1759,In_669,In_557);
xor U1760 (N_1760,In_78,In_383);
or U1761 (N_1761,In_932,In_635);
and U1762 (N_1762,In_18,In_526);
or U1763 (N_1763,In_630,In_546);
xnor U1764 (N_1764,In_470,In_147);
and U1765 (N_1765,In_60,In_413);
nor U1766 (N_1766,In_183,In_836);
or U1767 (N_1767,In_410,In_720);
xnor U1768 (N_1768,In_223,In_124);
or U1769 (N_1769,In_933,In_711);
nand U1770 (N_1770,In_422,In_51);
nand U1771 (N_1771,In_377,In_831);
nand U1772 (N_1772,In_703,In_626);
nand U1773 (N_1773,In_748,In_600);
nor U1774 (N_1774,In_488,In_225);
nand U1775 (N_1775,In_567,In_99);
and U1776 (N_1776,In_521,In_956);
and U1777 (N_1777,In_866,In_88);
and U1778 (N_1778,In_50,In_815);
or U1779 (N_1779,In_299,In_571);
nor U1780 (N_1780,In_276,In_711);
xnor U1781 (N_1781,In_148,In_970);
xor U1782 (N_1782,In_459,In_792);
or U1783 (N_1783,In_1,In_769);
nand U1784 (N_1784,In_872,In_46);
xnor U1785 (N_1785,In_855,In_349);
nand U1786 (N_1786,In_562,In_35);
or U1787 (N_1787,In_946,In_808);
or U1788 (N_1788,In_839,In_309);
or U1789 (N_1789,In_259,In_189);
nand U1790 (N_1790,In_701,In_282);
and U1791 (N_1791,In_675,In_184);
nand U1792 (N_1792,In_442,In_77);
or U1793 (N_1793,In_864,In_641);
nor U1794 (N_1794,In_805,In_967);
nor U1795 (N_1795,In_635,In_333);
and U1796 (N_1796,In_325,In_508);
nor U1797 (N_1797,In_493,In_480);
and U1798 (N_1798,In_150,In_400);
xnor U1799 (N_1799,In_588,In_142);
xor U1800 (N_1800,In_845,In_260);
and U1801 (N_1801,In_907,In_566);
or U1802 (N_1802,In_191,In_903);
and U1803 (N_1803,In_828,In_147);
nand U1804 (N_1804,In_119,In_246);
nor U1805 (N_1805,In_735,In_652);
or U1806 (N_1806,In_593,In_787);
and U1807 (N_1807,In_42,In_917);
nand U1808 (N_1808,In_149,In_360);
nand U1809 (N_1809,In_18,In_466);
xnor U1810 (N_1810,In_949,In_50);
nand U1811 (N_1811,In_75,In_46);
and U1812 (N_1812,In_860,In_891);
xnor U1813 (N_1813,In_370,In_458);
xor U1814 (N_1814,In_452,In_695);
nor U1815 (N_1815,In_84,In_560);
and U1816 (N_1816,In_841,In_286);
or U1817 (N_1817,In_445,In_30);
xor U1818 (N_1818,In_454,In_717);
nand U1819 (N_1819,In_908,In_742);
or U1820 (N_1820,In_485,In_113);
or U1821 (N_1821,In_286,In_870);
or U1822 (N_1822,In_528,In_8);
nand U1823 (N_1823,In_902,In_336);
nand U1824 (N_1824,In_836,In_110);
nor U1825 (N_1825,In_809,In_145);
nor U1826 (N_1826,In_88,In_404);
nand U1827 (N_1827,In_479,In_745);
and U1828 (N_1828,In_392,In_484);
and U1829 (N_1829,In_655,In_509);
nor U1830 (N_1830,In_540,In_431);
nor U1831 (N_1831,In_344,In_956);
or U1832 (N_1832,In_194,In_167);
and U1833 (N_1833,In_108,In_234);
nand U1834 (N_1834,In_842,In_272);
xor U1835 (N_1835,In_480,In_488);
and U1836 (N_1836,In_400,In_534);
nand U1837 (N_1837,In_853,In_356);
nor U1838 (N_1838,In_195,In_278);
or U1839 (N_1839,In_549,In_110);
xor U1840 (N_1840,In_964,In_272);
and U1841 (N_1841,In_271,In_312);
nor U1842 (N_1842,In_209,In_52);
nand U1843 (N_1843,In_379,In_722);
nand U1844 (N_1844,In_236,In_773);
nor U1845 (N_1845,In_624,In_183);
and U1846 (N_1846,In_515,In_381);
nor U1847 (N_1847,In_147,In_196);
nand U1848 (N_1848,In_165,In_882);
nand U1849 (N_1849,In_626,In_393);
and U1850 (N_1850,In_581,In_804);
xnor U1851 (N_1851,In_793,In_759);
nand U1852 (N_1852,In_478,In_877);
xnor U1853 (N_1853,In_719,In_903);
and U1854 (N_1854,In_575,In_339);
nor U1855 (N_1855,In_809,In_594);
and U1856 (N_1856,In_705,In_620);
and U1857 (N_1857,In_722,In_858);
or U1858 (N_1858,In_106,In_390);
and U1859 (N_1859,In_768,In_570);
nor U1860 (N_1860,In_236,In_395);
xnor U1861 (N_1861,In_249,In_991);
nand U1862 (N_1862,In_814,In_402);
nor U1863 (N_1863,In_426,In_31);
nor U1864 (N_1864,In_510,In_288);
or U1865 (N_1865,In_885,In_428);
nor U1866 (N_1866,In_671,In_825);
nor U1867 (N_1867,In_501,In_433);
and U1868 (N_1868,In_859,In_257);
xnor U1869 (N_1869,In_550,In_392);
nor U1870 (N_1870,In_652,In_86);
or U1871 (N_1871,In_791,In_474);
xnor U1872 (N_1872,In_788,In_234);
xnor U1873 (N_1873,In_754,In_920);
or U1874 (N_1874,In_137,In_14);
or U1875 (N_1875,In_61,In_724);
or U1876 (N_1876,In_207,In_606);
nand U1877 (N_1877,In_116,In_186);
xor U1878 (N_1878,In_79,In_423);
nor U1879 (N_1879,In_879,In_80);
nor U1880 (N_1880,In_279,In_893);
and U1881 (N_1881,In_332,In_14);
and U1882 (N_1882,In_139,In_384);
or U1883 (N_1883,In_629,In_513);
xor U1884 (N_1884,In_517,In_247);
and U1885 (N_1885,In_722,In_854);
nor U1886 (N_1886,In_941,In_986);
xnor U1887 (N_1887,In_878,In_780);
nor U1888 (N_1888,In_37,In_94);
and U1889 (N_1889,In_284,In_645);
and U1890 (N_1890,In_695,In_758);
xnor U1891 (N_1891,In_542,In_823);
or U1892 (N_1892,In_99,In_953);
or U1893 (N_1893,In_343,In_868);
xor U1894 (N_1894,In_939,In_84);
xor U1895 (N_1895,In_603,In_849);
nor U1896 (N_1896,In_844,In_848);
nor U1897 (N_1897,In_555,In_77);
or U1898 (N_1898,In_374,In_614);
or U1899 (N_1899,In_170,In_471);
and U1900 (N_1900,In_13,In_486);
nand U1901 (N_1901,In_876,In_710);
and U1902 (N_1902,In_141,In_26);
or U1903 (N_1903,In_762,In_872);
nand U1904 (N_1904,In_910,In_627);
xor U1905 (N_1905,In_711,In_929);
and U1906 (N_1906,In_578,In_559);
nor U1907 (N_1907,In_386,In_874);
or U1908 (N_1908,In_160,In_289);
xor U1909 (N_1909,In_332,In_857);
or U1910 (N_1910,In_729,In_546);
xnor U1911 (N_1911,In_672,In_543);
xnor U1912 (N_1912,In_76,In_782);
or U1913 (N_1913,In_187,In_374);
nor U1914 (N_1914,In_520,In_922);
xor U1915 (N_1915,In_200,In_632);
nand U1916 (N_1916,In_553,In_573);
nand U1917 (N_1917,In_888,In_828);
xor U1918 (N_1918,In_137,In_731);
nor U1919 (N_1919,In_985,In_670);
nand U1920 (N_1920,In_637,In_294);
and U1921 (N_1921,In_148,In_124);
or U1922 (N_1922,In_836,In_492);
xor U1923 (N_1923,In_971,In_637);
nand U1924 (N_1924,In_103,In_131);
or U1925 (N_1925,In_969,In_460);
nand U1926 (N_1926,In_810,In_788);
or U1927 (N_1927,In_100,In_48);
nand U1928 (N_1928,In_595,In_625);
nor U1929 (N_1929,In_607,In_478);
nand U1930 (N_1930,In_649,In_741);
nor U1931 (N_1931,In_819,In_76);
and U1932 (N_1932,In_891,In_336);
nor U1933 (N_1933,In_946,In_896);
nor U1934 (N_1934,In_553,In_387);
or U1935 (N_1935,In_359,In_379);
nand U1936 (N_1936,In_448,In_744);
or U1937 (N_1937,In_510,In_695);
nand U1938 (N_1938,In_873,In_623);
nor U1939 (N_1939,In_428,In_530);
nor U1940 (N_1940,In_623,In_418);
or U1941 (N_1941,In_439,In_146);
nand U1942 (N_1942,In_37,In_622);
nand U1943 (N_1943,In_670,In_257);
nand U1944 (N_1944,In_718,In_146);
nand U1945 (N_1945,In_112,In_661);
or U1946 (N_1946,In_232,In_935);
xnor U1947 (N_1947,In_758,In_824);
or U1948 (N_1948,In_657,In_995);
or U1949 (N_1949,In_384,In_909);
xnor U1950 (N_1950,In_188,In_738);
xnor U1951 (N_1951,In_18,In_310);
nor U1952 (N_1952,In_686,In_925);
nand U1953 (N_1953,In_653,In_62);
nand U1954 (N_1954,In_546,In_418);
nor U1955 (N_1955,In_16,In_243);
nor U1956 (N_1956,In_319,In_654);
nor U1957 (N_1957,In_495,In_956);
or U1958 (N_1958,In_416,In_382);
nor U1959 (N_1959,In_360,In_861);
or U1960 (N_1960,In_41,In_154);
nor U1961 (N_1961,In_482,In_107);
nand U1962 (N_1962,In_670,In_660);
nor U1963 (N_1963,In_305,In_515);
or U1964 (N_1964,In_447,In_819);
nor U1965 (N_1965,In_511,In_674);
and U1966 (N_1966,In_161,In_925);
nor U1967 (N_1967,In_294,In_454);
xor U1968 (N_1968,In_414,In_817);
xnor U1969 (N_1969,In_915,In_905);
nor U1970 (N_1970,In_937,In_753);
nor U1971 (N_1971,In_607,In_82);
nand U1972 (N_1972,In_200,In_198);
and U1973 (N_1973,In_482,In_779);
or U1974 (N_1974,In_237,In_658);
nor U1975 (N_1975,In_234,In_491);
nor U1976 (N_1976,In_716,In_292);
nand U1977 (N_1977,In_193,In_361);
nand U1978 (N_1978,In_722,In_396);
xor U1979 (N_1979,In_715,In_922);
and U1980 (N_1980,In_724,In_619);
nor U1981 (N_1981,In_617,In_387);
or U1982 (N_1982,In_116,In_971);
and U1983 (N_1983,In_935,In_975);
or U1984 (N_1984,In_733,In_216);
and U1985 (N_1985,In_864,In_888);
or U1986 (N_1986,In_106,In_555);
nand U1987 (N_1987,In_437,In_835);
or U1988 (N_1988,In_820,In_461);
xor U1989 (N_1989,In_864,In_791);
or U1990 (N_1990,In_851,In_673);
nor U1991 (N_1991,In_189,In_60);
xnor U1992 (N_1992,In_554,In_627);
and U1993 (N_1993,In_826,In_275);
nand U1994 (N_1994,In_215,In_964);
or U1995 (N_1995,In_438,In_238);
nand U1996 (N_1996,In_829,In_233);
nand U1997 (N_1997,In_85,In_9);
and U1998 (N_1998,In_977,In_564);
nor U1999 (N_1999,In_644,In_388);
nor U2000 (N_2000,N_1261,N_580);
or U2001 (N_2001,N_1571,N_1889);
and U2002 (N_2002,N_774,N_585);
xnor U2003 (N_2003,N_1290,N_1855);
nand U2004 (N_2004,N_571,N_511);
or U2005 (N_2005,N_625,N_226);
nand U2006 (N_2006,N_767,N_543);
nand U2007 (N_2007,N_1471,N_553);
nor U2008 (N_2008,N_312,N_1016);
nor U2009 (N_2009,N_151,N_1465);
xor U2010 (N_2010,N_1888,N_1627);
nor U2011 (N_2011,N_549,N_1552);
or U2012 (N_2012,N_1869,N_1864);
or U2013 (N_2013,N_1553,N_1061);
xnor U2014 (N_2014,N_956,N_1131);
nor U2015 (N_2015,N_1736,N_1017);
nor U2016 (N_2016,N_1718,N_375);
nor U2017 (N_2017,N_1455,N_1668);
or U2018 (N_2018,N_1582,N_902);
xor U2019 (N_2019,N_797,N_241);
and U2020 (N_2020,N_412,N_939);
nand U2021 (N_2021,N_411,N_1661);
and U2022 (N_2022,N_1273,N_1007);
nor U2023 (N_2023,N_1015,N_1699);
and U2024 (N_2024,N_1097,N_1228);
nor U2025 (N_2025,N_1789,N_1875);
or U2026 (N_2026,N_1049,N_666);
nand U2027 (N_2027,N_1883,N_1091);
nor U2028 (N_2028,N_1504,N_1766);
nand U2029 (N_2029,N_555,N_1986);
nor U2030 (N_2030,N_1164,N_1198);
or U2031 (N_2031,N_1113,N_1490);
nand U2032 (N_2032,N_1881,N_888);
nand U2033 (N_2033,N_20,N_1293);
or U2034 (N_2034,N_970,N_66);
or U2035 (N_2035,N_121,N_1344);
xor U2036 (N_2036,N_381,N_1363);
nand U2037 (N_2037,N_1054,N_367);
or U2038 (N_2038,N_1102,N_463);
nor U2039 (N_2039,N_660,N_1051);
and U2040 (N_2040,N_1080,N_1006);
nor U2041 (N_2041,N_1499,N_248);
nor U2042 (N_2042,N_1682,N_1480);
nand U2043 (N_2043,N_1897,N_1414);
nor U2044 (N_2044,N_649,N_1491);
nand U2045 (N_2045,N_793,N_1744);
or U2046 (N_2046,N_1133,N_250);
or U2047 (N_2047,N_910,N_1222);
nand U2048 (N_2048,N_328,N_1686);
or U2049 (N_2049,N_1128,N_1852);
nand U2050 (N_2050,N_990,N_1568);
and U2051 (N_2051,N_810,N_805);
or U2052 (N_2052,N_1443,N_1447);
xnor U2053 (N_2053,N_1655,N_1749);
and U2054 (N_2054,N_822,N_1650);
nand U2055 (N_2055,N_434,N_1757);
or U2056 (N_2056,N_1068,N_30);
xor U2057 (N_2057,N_304,N_1969);
nand U2058 (N_2058,N_841,N_1925);
nand U2059 (N_2059,N_1329,N_1468);
nor U2060 (N_2060,N_460,N_746);
or U2061 (N_2061,N_1478,N_994);
nor U2062 (N_2062,N_1115,N_1044);
or U2063 (N_2063,N_545,N_1274);
nor U2064 (N_2064,N_1625,N_1633);
and U2065 (N_2065,N_343,N_22);
or U2066 (N_2066,N_680,N_740);
nor U2067 (N_2067,N_1887,N_407);
xnor U2068 (N_2068,N_1385,N_1435);
nor U2069 (N_2069,N_64,N_1771);
and U2070 (N_2070,N_148,N_352);
and U2071 (N_2071,N_536,N_1278);
nor U2072 (N_2072,N_1166,N_642);
nor U2073 (N_2073,N_1246,N_708);
and U2074 (N_2074,N_441,N_11);
or U2075 (N_2075,N_1157,N_1907);
or U2076 (N_2076,N_1460,N_733);
nand U2077 (N_2077,N_4,N_648);
and U2078 (N_2078,N_1783,N_1482);
or U2079 (N_2079,N_1843,N_100);
nor U2080 (N_2080,N_1250,N_19);
and U2081 (N_2081,N_1900,N_1701);
xnor U2082 (N_2082,N_809,N_147);
or U2083 (N_2083,N_41,N_907);
and U2084 (N_2084,N_849,N_317);
nand U2085 (N_2085,N_1603,N_1972);
or U2086 (N_2086,N_567,N_1801);
and U2087 (N_2087,N_776,N_1241);
and U2088 (N_2088,N_815,N_1866);
xor U2089 (N_2089,N_1404,N_1782);
xor U2090 (N_2090,N_495,N_1464);
xnor U2091 (N_2091,N_1560,N_561);
nor U2092 (N_2092,N_1338,N_1658);
xor U2093 (N_2093,N_357,N_337);
or U2094 (N_2094,N_1013,N_679);
xnor U2095 (N_2095,N_1424,N_1963);
or U2096 (N_2096,N_1772,N_1470);
nand U2097 (N_2097,N_1187,N_506);
nor U2098 (N_2098,N_424,N_481);
and U2099 (N_2099,N_905,N_391);
or U2100 (N_2100,N_1743,N_627);
xnor U2101 (N_2101,N_880,N_1430);
xnor U2102 (N_2102,N_1590,N_759);
xnor U2103 (N_2103,N_425,N_1577);
nand U2104 (N_2104,N_1215,N_807);
and U2105 (N_2105,N_1253,N_1175);
nor U2106 (N_2106,N_1980,N_216);
nand U2107 (N_2107,N_1702,N_1269);
and U2108 (N_2108,N_593,N_1725);
and U2109 (N_2109,N_36,N_1971);
xnor U2110 (N_2110,N_341,N_1635);
nand U2111 (N_2111,N_632,N_431);
xor U2112 (N_2112,N_347,N_1506);
or U2113 (N_2113,N_871,N_96);
nor U2114 (N_2114,N_240,N_950);
nor U2115 (N_2115,N_227,N_535);
nand U2116 (N_2116,N_618,N_724);
nand U2117 (N_2117,N_450,N_484);
xnor U2118 (N_2118,N_894,N_1354);
nor U2119 (N_2119,N_854,N_1401);
xor U2120 (N_2120,N_1088,N_75);
and U2121 (N_2121,N_73,N_1310);
nand U2122 (N_2122,N_996,N_1275);
nand U2123 (N_2123,N_1585,N_1056);
xor U2124 (N_2124,N_438,N_262);
nor U2125 (N_2125,N_1217,N_6);
and U2126 (N_2126,N_541,N_1352);
nand U2127 (N_2127,N_1841,N_953);
and U2128 (N_2128,N_160,N_1377);
nor U2129 (N_2129,N_35,N_847);
or U2130 (N_2130,N_1285,N_1365);
or U2131 (N_2131,N_168,N_726);
nor U2132 (N_2132,N_1410,N_1838);
xor U2133 (N_2133,N_823,N_967);
nor U2134 (N_2134,N_1985,N_743);
xnor U2135 (N_2135,N_1437,N_417);
and U2136 (N_2136,N_436,N_1865);
nand U2137 (N_2137,N_1652,N_772);
xnor U2138 (N_2138,N_1878,N_808);
nand U2139 (N_2139,N_635,N_668);
or U2140 (N_2140,N_1555,N_1713);
and U2141 (N_2141,N_1676,N_579);
xor U2142 (N_2142,N_500,N_1512);
xnor U2143 (N_2143,N_863,N_951);
nand U2144 (N_2144,N_1067,N_1752);
nand U2145 (N_2145,N_1557,N_1545);
nor U2146 (N_2146,N_1669,N_255);
nand U2147 (N_2147,N_695,N_91);
or U2148 (N_2148,N_451,N_235);
or U2149 (N_2149,N_1353,N_1853);
xor U2150 (N_2150,N_249,N_470);
nor U2151 (N_2151,N_1589,N_99);
or U2152 (N_2152,N_758,N_1271);
xor U2153 (N_2153,N_1313,N_984);
nand U2154 (N_2154,N_1909,N_1305);
nor U2155 (N_2155,N_1847,N_496);
xnor U2156 (N_2156,N_442,N_886);
and U2157 (N_2157,N_1562,N_1340);
nor U2158 (N_2158,N_389,N_993);
or U2159 (N_2159,N_1683,N_229);
nand U2160 (N_2160,N_497,N_46);
and U2161 (N_2161,N_1674,N_275);
nor U2162 (N_2162,N_1476,N_912);
xnor U2163 (N_2163,N_669,N_1461);
xnor U2164 (N_2164,N_715,N_205);
nand U2165 (N_2165,N_1386,N_1192);
nand U2166 (N_2166,N_140,N_1330);
nor U2167 (N_2167,N_59,N_1180);
or U2168 (N_2168,N_1662,N_992);
nor U2169 (N_2169,N_1944,N_1910);
or U2170 (N_2170,N_298,N_1832);
nand U2171 (N_2171,N_1472,N_1096);
nor U2172 (N_2172,N_1953,N_489);
xnor U2173 (N_2173,N_1724,N_673);
nand U2174 (N_2174,N_801,N_1999);
nand U2175 (N_2175,N_1204,N_1009);
xnor U2176 (N_2176,N_1492,N_29);
and U2177 (N_2177,N_1197,N_1828);
and U2178 (N_2178,N_1341,N_1267);
or U2179 (N_2179,N_1272,N_1750);
nand U2180 (N_2180,N_507,N_1099);
xor U2181 (N_2181,N_640,N_595);
nor U2182 (N_2182,N_1554,N_1334);
xnor U2183 (N_2183,N_1418,N_641);
and U2184 (N_2184,N_385,N_980);
or U2185 (N_2185,N_725,N_1549);
nor U2186 (N_2186,N_603,N_409);
nor U2187 (N_2187,N_1628,N_1558);
nor U2188 (N_2188,N_1928,N_314);
nand U2189 (N_2189,N_1979,N_1758);
or U2190 (N_2190,N_303,N_1422);
or U2191 (N_2191,N_927,N_416);
nor U2192 (N_2192,N_614,N_1225);
nand U2193 (N_2193,N_524,N_1916);
and U2194 (N_2194,N_859,N_1439);
and U2195 (N_2195,N_1629,N_1020);
and U2196 (N_2196,N_1734,N_1729);
nand U2197 (N_2197,N_1135,N_582);
nand U2198 (N_2198,N_1587,N_97);
nor U2199 (N_2199,N_1178,N_1130);
xnor U2200 (N_2200,N_1011,N_1239);
or U2201 (N_2201,N_414,N_306);
nand U2202 (N_2202,N_1234,N_483);
xnor U2203 (N_2203,N_1389,N_1815);
nand U2204 (N_2204,N_435,N_187);
nor U2205 (N_2205,N_1369,N_1093);
or U2206 (N_2206,N_1935,N_1008);
and U2207 (N_2207,N_39,N_1646);
nor U2208 (N_2208,N_316,N_1173);
nor U2209 (N_2209,N_399,N_1203);
and U2210 (N_2210,N_891,N_1859);
nand U2211 (N_2211,N_1429,N_869);
xnor U2212 (N_2212,N_1988,N_1738);
nand U2213 (N_2213,N_1901,N_1580);
nor U2214 (N_2214,N_946,N_1446);
xor U2215 (N_2215,N_42,N_534);
or U2216 (N_2216,N_1235,N_1835);
nor U2217 (N_2217,N_51,N_761);
nor U2218 (N_2218,N_1947,N_210);
xor U2219 (N_2219,N_1136,N_792);
xor U2220 (N_2220,N_1825,N_853);
nand U2221 (N_2221,N_445,N_1371);
or U2222 (N_2222,N_1452,N_152);
nand U2223 (N_2223,N_1308,N_836);
or U2224 (N_2224,N_709,N_447);
nor U2225 (N_2225,N_736,N_1005);
or U2226 (N_2226,N_1882,N_1262);
nand U2227 (N_2227,N_1268,N_1026);
xnor U2228 (N_2228,N_831,N_1170);
or U2229 (N_2229,N_1551,N_1194);
xnor U2230 (N_2230,N_1638,N_134);
and U2231 (N_2231,N_1547,N_581);
and U2232 (N_2232,N_365,N_1681);
nand U2233 (N_2233,N_218,N_492);
nor U2234 (N_2234,N_1040,N_464);
xor U2235 (N_2235,N_1531,N_1861);
nand U2236 (N_2236,N_790,N_943);
or U2237 (N_2237,N_1599,N_1817);
or U2238 (N_2238,N_1448,N_1903);
or U2239 (N_2239,N_1886,N_26);
and U2240 (N_2240,N_881,N_1438);
xnor U2241 (N_2241,N_832,N_1937);
xor U2242 (N_2242,N_1231,N_1704);
or U2243 (N_2243,N_879,N_321);
nor U2244 (N_2244,N_1375,N_896);
and U2245 (N_2245,N_1821,N_128);
and U2246 (N_2246,N_1779,N_781);
xor U2247 (N_2247,N_565,N_141);
and U2248 (N_2248,N_1014,N_1189);
nand U2249 (N_2249,N_1107,N_1717);
xor U2250 (N_2250,N_634,N_56);
or U2251 (N_2251,N_1836,N_755);
nand U2252 (N_2252,N_514,N_393);
nand U2253 (N_2253,N_884,N_194);
or U2254 (N_2254,N_899,N_518);
nor U2255 (N_2255,N_1920,N_207);
and U2256 (N_2256,N_1383,N_629);
xnor U2257 (N_2257,N_1319,N_770);
nand U2258 (N_2258,N_966,N_1079);
and U2259 (N_2259,N_1679,N_728);
nor U2260 (N_2260,N_935,N_1915);
or U2261 (N_2261,N_475,N_558);
or U2262 (N_2262,N_164,N_1670);
or U2263 (N_2263,N_127,N_615);
nand U2264 (N_2264,N_1742,N_336);
and U2265 (N_2265,N_771,N_1110);
or U2266 (N_2266,N_833,N_1169);
and U2267 (N_2267,N_491,N_1588);
or U2268 (N_2268,N_1100,N_1024);
xnor U2269 (N_2269,N_319,N_1144);
nand U2270 (N_2270,N_1498,N_55);
nand U2271 (N_2271,N_1824,N_837);
nand U2272 (N_2272,N_1507,N_1756);
or U2273 (N_2273,N_1966,N_146);
or U2274 (N_2274,N_1707,N_397);
or U2275 (N_2275,N_114,N_1712);
nand U2276 (N_2276,N_1158,N_1733);
xnor U2277 (N_2277,N_201,N_546);
xnor U2278 (N_2278,N_313,N_1398);
nor U2279 (N_2279,N_707,N_247);
nand U2280 (N_2280,N_1373,N_1324);
xnor U2281 (N_2281,N_297,N_1450);
and U2282 (N_2282,N_50,N_130);
or U2283 (N_2283,N_1309,N_295);
nor U2284 (N_2284,N_92,N_1645);
xnor U2285 (N_2285,N_1703,N_1496);
nand U2286 (N_2286,N_145,N_1572);
nor U2287 (N_2287,N_530,N_60);
xor U2288 (N_2288,N_1412,N_1112);
nor U2289 (N_2289,N_1103,N_1109);
xor U2290 (N_2290,N_874,N_1207);
nand U2291 (N_2291,N_527,N_28);
and U2292 (N_2292,N_1322,N_637);
and U2293 (N_2293,N_499,N_2);
nor U2294 (N_2294,N_1312,N_1493);
and U2295 (N_2295,N_394,N_623);
or U2296 (N_2296,N_933,N_800);
xnor U2297 (N_2297,N_1095,N_320);
and U2298 (N_2298,N_296,N_1680);
nand U2299 (N_2299,N_83,N_911);
xor U2300 (N_2300,N_701,N_1163);
and U2301 (N_2301,N_311,N_37);
nand U2302 (N_2302,N_693,N_1974);
nor U2303 (N_2303,N_351,N_1238);
and U2304 (N_2304,N_165,N_1002);
or U2305 (N_2305,N_238,N_1863);
xor U2306 (N_2306,N_677,N_1047);
xor U2307 (N_2307,N_1069,N_12);
and U2308 (N_2308,N_813,N_508);
nor U2309 (N_2309,N_1797,N_504);
xnor U2310 (N_2310,N_428,N_193);
or U2311 (N_2311,N_291,N_1754);
nor U2312 (N_2312,N_1891,N_1101);
xor U2313 (N_2313,N_1519,N_1933);
and U2314 (N_2314,N_510,N_760);
nor U2315 (N_2315,N_178,N_1902);
xor U2316 (N_2316,N_163,N_835);
or U2317 (N_2317,N_877,N_584);
xnor U2318 (N_2318,N_117,N_1073);
xnor U2319 (N_2319,N_1800,N_1433);
or U2320 (N_2320,N_1081,N_554);
and U2321 (N_2321,N_1029,N_254);
nand U2322 (N_2322,N_1997,N_268);
xnor U2323 (N_2323,N_1129,N_1142);
xor U2324 (N_2324,N_1532,N_1610);
nand U2325 (N_2325,N_1297,N_1848);
xnor U2326 (N_2326,N_186,N_1030);
and U2327 (N_2327,N_1413,N_1708);
and U2328 (N_2328,N_1339,N_826);
nor U2329 (N_2329,N_1632,N_1172);
or U2330 (N_2330,N_969,N_1114);
nand U2331 (N_2331,N_155,N_78);
nor U2332 (N_2332,N_763,N_852);
nor U2333 (N_2333,N_222,N_1611);
nor U2334 (N_2334,N_1311,N_600);
or U2335 (N_2335,N_1584,N_1174);
nor U2336 (N_2336,N_62,N_202);
and U2337 (N_2337,N_1042,N_1380);
or U2338 (N_2338,N_479,N_748);
xor U2339 (N_2339,N_261,N_271);
and U2340 (N_2340,N_1417,N_941);
or U2341 (N_2341,N_702,N_1509);
xnor U2342 (N_2342,N_1539,N_1563);
nor U2343 (N_2343,N_875,N_1535);
or U2344 (N_2344,N_1479,N_775);
nor U2345 (N_2345,N_1576,N_1595);
xnor U2346 (N_2346,N_1762,N_591);
xnor U2347 (N_2347,N_1503,N_1591);
and U2348 (N_2348,N_1994,N_1242);
or U2349 (N_2349,N_1614,N_1899);
or U2350 (N_2350,N_1561,N_1475);
or U2351 (N_2351,N_821,N_686);
or U2352 (N_2352,N_1249,N_1892);
and U2353 (N_2353,N_1990,N_456);
and U2354 (N_2354,N_667,N_1487);
and U2355 (N_2355,N_1391,N_133);
xor U2356 (N_2356,N_267,N_348);
xnor U2357 (N_2357,N_1639,N_15);
or U2358 (N_2358,N_1653,N_1601);
nand U2359 (N_2359,N_681,N_895);
nor U2360 (N_2360,N_1155,N_1799);
nor U2361 (N_2361,N_1202,N_924);
nor U2362 (N_2362,N_1959,N_112);
or U2363 (N_2363,N_1667,N_806);
xnor U2364 (N_2364,N_960,N_936);
xnor U2365 (N_2365,N_277,N_851);
or U2366 (N_2366,N_1876,N_1457);
xnor U2367 (N_2367,N_929,N_270);
and U2368 (N_2368,N_1569,N_958);
or U2369 (N_2369,N_848,N_171);
or U2370 (N_2370,N_1001,N_1399);
xor U2371 (N_2371,N_1511,N_1540);
xor U2372 (N_2372,N_636,N_1279);
or U2373 (N_2373,N_997,N_1440);
xor U2374 (N_2374,N_377,N_1098);
nand U2375 (N_2375,N_477,N_104);
and U2376 (N_2376,N_1780,N_742);
xnor U2377 (N_2377,N_674,N_1908);
or U2378 (N_2378,N_116,N_1119);
nand U2379 (N_2379,N_283,N_949);
and U2380 (N_2380,N_1502,N_945);
nor U2381 (N_2381,N_1454,N_1181);
nand U2382 (N_2382,N_991,N_1488);
xor U2383 (N_2383,N_154,N_865);
nand U2384 (N_2384,N_1027,N_973);
or U2385 (N_2385,N_185,N_43);
xor U2386 (N_2386,N_289,N_1956);
xor U2387 (N_2387,N_1252,N_467);
nand U2388 (N_2388,N_687,N_690);
and U2389 (N_2389,N_1445,N_1153);
nor U2390 (N_2390,N_1931,N_1716);
nand U2391 (N_2391,N_1141,N_95);
or U2392 (N_2392,N_421,N_1776);
and U2393 (N_2393,N_111,N_883);
nor U2394 (N_2394,N_906,N_1400);
nor U2395 (N_2395,N_1695,N_1419);
xnor U2396 (N_2396,N_756,N_482);
xor U2397 (N_2397,N_979,N_211);
and U2398 (N_2398,N_1523,N_1760);
nand U2399 (N_2399,N_455,N_215);
or U2400 (N_2400,N_318,N_1431);
nor U2401 (N_2401,N_1199,N_70);
xor U2402 (N_2402,N_488,N_1379);
nand U2403 (N_2403,N_274,N_1602);
nand U2404 (N_2404,N_711,N_619);
or U2405 (N_2405,N_778,N_490);
nor U2406 (N_2406,N_714,N_1343);
xor U2407 (N_2407,N_1930,N_1402);
nand U2408 (N_2408,N_1781,N_374);
nand U2409 (N_2409,N_94,N_1684);
nand U2410 (N_2410,N_332,N_1062);
nand U2411 (N_2411,N_560,N_1996);
nand U2412 (N_2412,N_1162,N_444);
nor U2413 (N_2413,N_192,N_1317);
and U2414 (N_2414,N_878,N_61);
and U2415 (N_2415,N_1600,N_1849);
and U2416 (N_2416,N_818,N_1395);
xor U2417 (N_2417,N_175,N_1700);
or U2418 (N_2418,N_689,N_420);
or U2419 (N_2419,N_1301,N_1927);
xnor U2420 (N_2420,N_243,N_144);
xor U2421 (N_2421,N_184,N_74);
or U2422 (N_2422,N_1630,N_260);
xor U2423 (N_2423,N_360,N_696);
or U2424 (N_2424,N_676,N_1678);
and U2425 (N_2425,N_418,N_1046);
nand U2426 (N_2426,N_1578,N_376);
nor U2427 (N_2427,N_578,N_93);
and U2428 (N_2428,N_440,N_915);
and U2429 (N_2429,N_1583,N_744);
and U2430 (N_2430,N_1739,N_532);
nand U2431 (N_2431,N_1229,N_1436);
xor U2432 (N_2432,N_299,N_131);
and U2433 (N_2433,N_143,N_1723);
xor U2434 (N_2434,N_1518,N_498);
and U2435 (N_2435,N_137,N_404);
or U2436 (N_2436,N_392,N_181);
or U2437 (N_2437,N_388,N_1809);
xnor U2438 (N_2438,N_862,N_605);
xor U2439 (N_2439,N_1070,N_612);
nand U2440 (N_2440,N_1608,N_1906);
xnor U2441 (N_2441,N_176,N_938);
nor U2442 (N_2442,N_1884,N_1484);
nand U2443 (N_2443,N_802,N_1378);
or U2444 (N_2444,N_1209,N_24);
nand U2445 (N_2445,N_1307,N_1286);
or U2446 (N_2446,N_5,N_722);
and U2447 (N_2447,N_1367,N_1168);
nand U2448 (N_2448,N_236,N_16);
nor U2449 (N_2449,N_1387,N_1932);
and U2450 (N_2450,N_493,N_322);
and U2451 (N_2451,N_1634,N_426);
nor U2452 (N_2452,N_505,N_1082);
nand U2453 (N_2453,N_1818,N_570);
and U2454 (N_2454,N_452,N_564);
and U2455 (N_2455,N_780,N_1221);
xnor U2456 (N_2456,N_123,N_650);
and U2457 (N_2457,N_188,N_1872);
nor U2458 (N_2458,N_1698,N_1605);
or U2459 (N_2459,N_1137,N_1534);
nor U2460 (N_2460,N_63,N_1421);
xor U2461 (N_2461,N_480,N_982);
or U2462 (N_2462,N_525,N_1654);
and U2463 (N_2463,N_1566,N_1770);
and U2464 (N_2464,N_1374,N_860);
and U2465 (N_2465,N_45,N_342);
nor U2466 (N_2466,N_245,N_1620);
and U2467 (N_2467,N_150,N_7);
and U2468 (N_2468,N_937,N_975);
nor U2469 (N_2469,N_485,N_1300);
xnor U2470 (N_2470,N_1362,N_1598);
nand U2471 (N_2471,N_370,N_784);
or U2472 (N_2472,N_1793,N_827);
nor U2473 (N_2473,N_232,N_700);
nor U2474 (N_2474,N_1767,N_597);
nand U2475 (N_2475,N_177,N_1924);
nand U2476 (N_2476,N_972,N_526);
nand U2477 (N_2477,N_69,N_638);
or U2478 (N_2478,N_225,N_1525);
nor U2479 (N_2479,N_791,N_182);
and U2480 (N_2480,N_1923,N_1184);
xnor U2481 (N_2481,N_1328,N_577);
nor U2482 (N_2482,N_914,N_52);
xnor U2483 (N_2483,N_1983,N_1537);
and U2484 (N_2484,N_665,N_10);
xnor U2485 (N_2485,N_189,N_1366);
nand U2486 (N_2486,N_413,N_1453);
xor U2487 (N_2487,N_462,N_408);
and U2488 (N_2488,N_1057,N_473);
or U2489 (N_2489,N_1232,N_132);
or U2490 (N_2490,N_1810,N_346);
nand U2491 (N_2491,N_1121,N_279);
nand U2492 (N_2492,N_1403,N_1117);
xnor U2493 (N_2493,N_1579,N_1124);
xnor U2494 (N_2494,N_820,N_940);
or U2495 (N_2495,N_1945,N_1660);
or U2496 (N_2496,N_1053,N_622);
nand U2497 (N_2497,N_934,N_656);
or U2498 (N_2498,N_513,N_1467);
and U2499 (N_2499,N_655,N_1792);
xnor U2500 (N_2500,N_988,N_1710);
nor U2501 (N_2501,N_1500,N_1298);
nand U2502 (N_2502,N_1694,N_1182);
nor U2503 (N_2503,N_1473,N_1407);
xor U2504 (N_2504,N_1415,N_1621);
and U2505 (N_2505,N_1939,N_9);
nand U2506 (N_2506,N_1023,N_1977);
nand U2507 (N_2507,N_293,N_1874);
nand U2508 (N_2508,N_195,N_1466);
or U2509 (N_2509,N_1449,N_469);
nor U2510 (N_2510,N_1247,N_1485);
or U2511 (N_2511,N_98,N_1975);
nor U2512 (N_2512,N_691,N_1462);
or U2513 (N_2513,N_1641,N_1294);
xnor U2514 (N_2514,N_1753,N_1179);
nor U2515 (N_2515,N_1616,N_1992);
or U2516 (N_2516,N_387,N_520);
nor U2517 (N_2517,N_1200,N_1105);
nand U2518 (N_2518,N_1567,N_1880);
nand U2519 (N_2519,N_1954,N_356);
or U2520 (N_2520,N_276,N_1218);
xnor U2521 (N_2521,N_1636,N_183);
nor U2522 (N_2522,N_1149,N_657);
nor U2523 (N_2523,N_162,N_1786);
nand U2524 (N_2524,N_196,N_643);
nand U2525 (N_2525,N_1592,N_1885);
nor U2526 (N_2526,N_1230,N_926);
or U2527 (N_2527,N_105,N_864);
xor U2528 (N_2528,N_1648,N_824);
nor U2529 (N_2529,N_858,N_1325);
nor U2530 (N_2530,N_138,N_840);
xor U2531 (N_2531,N_1973,N_1607);
and U2532 (N_2532,N_769,N_108);
xor U2533 (N_2533,N_1777,N_17);
or U2534 (N_2534,N_557,N_1122);
or U2535 (N_2535,N_732,N_1727);
nor U2536 (N_2536,N_1227,N_741);
xnor U2537 (N_2537,N_1303,N_1675);
xnor U2538 (N_2538,N_698,N_1741);
or U2539 (N_2539,N_278,N_971);
or U2540 (N_2540,N_1474,N_1463);
xor U2541 (N_2541,N_735,N_955);
nand U2542 (N_2542,N_893,N_816);
nor U2543 (N_2543,N_995,N_1659);
nand U2544 (N_2544,N_1840,N_68);
nor U2545 (N_2545,N_1258,N_1071);
nand U2546 (N_2546,N_1522,N_90);
nor U2547 (N_2547,N_1905,N_796);
or U2548 (N_2548,N_103,N_1347);
nor U2549 (N_2549,N_1224,N_1597);
xor U2550 (N_2550,N_1991,N_1748);
nand U2551 (N_2551,N_964,N_443);
xnor U2552 (N_2552,N_512,N_335);
or U2553 (N_2553,N_706,N_963);
xor U2554 (N_2554,N_1524,N_1765);
or U2555 (N_2555,N_169,N_179);
nand U2556 (N_2556,N_729,N_209);
nor U2557 (N_2557,N_574,N_1586);
nand U2558 (N_2558,N_844,N_406);
nor U2559 (N_2559,N_542,N_645);
and U2560 (N_2560,N_531,N_1384);
nor U2561 (N_2561,N_113,N_1860);
xor U2562 (N_2562,N_1426,N_583);
nand U2563 (N_2563,N_38,N_1895);
or U2564 (N_2564,N_1349,N_1265);
or U2565 (N_2565,N_594,N_965);
nor U2566 (N_2566,N_1804,N_1735);
or U2567 (N_2567,N_1211,N_1609);
or U2568 (N_2568,N_718,N_323);
and U2569 (N_2569,N_233,N_1812);
nor U2570 (N_2570,N_242,N_1186);
nand U2571 (N_2571,N_954,N_1077);
nand U2572 (N_2572,N_1618,N_1719);
or U2573 (N_2573,N_1074,N_1893);
or U2574 (N_2574,N_925,N_1139);
nor U2575 (N_2575,N_1775,N_592);
xnor U2576 (N_2576,N_1260,N_1004);
and U2577 (N_2577,N_1706,N_1529);
nand U2578 (N_2578,N_1987,N_362);
nor U2579 (N_2579,N_986,N_1926);
nand U2580 (N_2580,N_798,N_1644);
nor U2581 (N_2581,N_868,N_1673);
and U2582 (N_2582,N_161,N_1711);
nand U2583 (N_2583,N_644,N_109);
and U2584 (N_2584,N_372,N_1526);
or U2585 (N_2585,N_49,N_1021);
or U2586 (N_2586,N_446,N_752);
and U2587 (N_2587,N_608,N_1);
xnor U2588 (N_2588,N_916,N_1768);
nor U2589 (N_2589,N_1236,N_1320);
or U2590 (N_2590,N_142,N_1314);
xnor U2591 (N_2591,N_1481,N_1394);
xor U2592 (N_2592,N_730,N_27);
xor U2593 (N_2593,N_602,N_415);
and U2594 (N_2594,N_361,N_1850);
xor U2595 (N_2595,N_461,N_432);
nor U2596 (N_2596,N_1877,N_684);
xnor U2597 (N_2597,N_1216,N_1556);
nor U2598 (N_2598,N_738,N_688);
or U2599 (N_2599,N_1904,N_699);
xnor U2600 (N_2600,N_1533,N_1981);
and U2601 (N_2601,N_745,N_890);
nand U2602 (N_2602,N_904,N_1671);
or U2603 (N_2603,N_1542,N_157);
and U2604 (N_2604,N_1649,N_930);
or U2605 (N_2605,N_604,N_857);
or U2606 (N_2606,N_620,N_1364);
xor U2607 (N_2607,N_1087,N_439);
or U2608 (N_2608,N_589,N_396);
nand U2609 (N_2609,N_659,N_794);
or U2610 (N_2610,N_928,N_1951);
and U2611 (N_2611,N_501,N_754);
and U2612 (N_2612,N_1715,N_872);
nand U2613 (N_2613,N_1643,N_1444);
and U2614 (N_2614,N_280,N_115);
xor U2615 (N_2615,N_1425,N_457);
and U2616 (N_2616,N_885,N_1890);
and U2617 (N_2617,N_158,N_562);
nand U2618 (N_2618,N_1528,N_1640);
xnor U2619 (N_2619,N_814,N_1769);
nor U2620 (N_2620,N_1120,N_1517);
nand U2621 (N_2621,N_694,N_803);
xor U2622 (N_2622,N_646,N_737);
and U2623 (N_2623,N_1896,N_675);
nor U2624 (N_2624,N_1108,N_633);
and U2625 (N_2625,N_1575,N_80);
and U2626 (N_2626,N_1796,N_1306);
or U2627 (N_2627,N_653,N_472);
and U2628 (N_2628,N_1918,N_1871);
xor U2629 (N_2629,N_1940,N_1257);
or U2630 (N_2630,N_1196,N_265);
xor U2631 (N_2631,N_159,N_952);
xor U2632 (N_2632,N_1791,N_363);
nand U2633 (N_2633,N_1287,N_1477);
nand U2634 (N_2634,N_654,N_1086);
nor U2635 (N_2635,N_244,N_1214);
nand U2636 (N_2636,N_474,N_1276);
nor U2637 (N_2637,N_1195,N_611);
and U2638 (N_2638,N_599,N_825);
nor U2639 (N_2639,N_32,N_465);
or U2640 (N_2640,N_309,N_1316);
and U2641 (N_2641,N_1516,N_843);
nor U2642 (N_2642,N_1949,N_1063);
nor U2643 (N_2643,N_1161,N_757);
nor U2644 (N_2644,N_1159,N_503);
xnor U2645 (N_2645,N_540,N_1745);
nand U2646 (N_2646,N_651,N_1388);
xor U2647 (N_2647,N_710,N_433);
and U2648 (N_2648,N_1574,N_383);
xor U2649 (N_2649,N_1914,N_1263);
and U2650 (N_2650,N_607,N_120);
nor U2651 (N_2651,N_1622,N_548);
nor U2652 (N_2652,N_364,N_199);
nand U2653 (N_2653,N_1240,N_1342);
nor U2654 (N_2654,N_1382,N_786);
or U2655 (N_2655,N_1245,N_325);
and U2656 (N_2656,N_44,N_1808);
or U2657 (N_2657,N_1665,N_1709);
nor U2658 (N_2658,N_1486,N_219);
nand U2659 (N_2659,N_609,N_1755);
nor U2660 (N_2660,N_1538,N_1085);
and U2661 (N_2661,N_1833,N_1612);
and U2662 (N_2662,N_1233,N_828);
or U2663 (N_2663,N_190,N_1434);
nor U2664 (N_2664,N_1160,N_85);
nor U2665 (N_2665,N_0,N_773);
or U2666 (N_2666,N_870,N_1190);
or U2667 (N_2667,N_1083,N_253);
nand U2668 (N_2668,N_919,N_1819);
nand U2669 (N_2669,N_1787,N_1092);
nand U2670 (N_2670,N_1176,N_1064);
nand U2671 (N_2671,N_1213,N_340);
xnor U2672 (N_2672,N_1337,N_1594);
or U2673 (N_2673,N_1795,N_1922);
and U2674 (N_2674,N_587,N_1147);
and U2675 (N_2675,N_269,N_948);
nor U2676 (N_2676,N_1565,N_359);
nand U2677 (N_2677,N_661,N_294);
nand U2678 (N_2678,N_81,N_47);
xor U2679 (N_2679,N_1688,N_1270);
xor U2680 (N_2680,N_256,N_237);
nor U2681 (N_2681,N_739,N_1223);
xnor U2682 (N_2682,N_1798,N_1167);
nor U2683 (N_2683,N_1302,N_1451);
xnor U2684 (N_2684,N_1581,N_1955);
nor U2685 (N_2685,N_974,N_1254);
xnor U2686 (N_2686,N_1469,N_1132);
nor U2687 (N_2687,N_898,N_734);
and U2688 (N_2688,N_172,N_987);
nor U2689 (N_2689,N_1266,N_521);
nand U2690 (N_2690,N_1003,N_1066);
nor U2691 (N_2691,N_920,N_1820);
and U2692 (N_2692,N_378,N_1857);
nor U2693 (N_2693,N_423,N_766);
xnor U2694 (N_2694,N_962,N_1370);
xnor U2695 (N_2695,N_288,N_1573);
and U2696 (N_2696,N_200,N_533);
xor U2697 (N_2697,N_1788,N_1489);
xnor U2698 (N_2698,N_305,N_1345);
or U2699 (N_2699,N_18,N_1123);
and U2700 (N_2700,N_779,N_1326);
or U2701 (N_2701,N_764,N_1596);
and U2702 (N_2702,N_1898,N_590);
and U2703 (N_2703,N_471,N_419);
or U2704 (N_2704,N_572,N_302);
xor U2705 (N_2705,N_173,N_566);
or U2706 (N_2706,N_547,N_1689);
or U2707 (N_2707,N_1631,N_1570);
and U2708 (N_2708,N_65,N_382);
xor U2709 (N_2709,N_197,N_327);
xor U2710 (N_2710,N_310,N_1606);
xor U2711 (N_2711,N_1012,N_1827);
nand U2712 (N_2712,N_1965,N_1019);
or U2713 (N_2713,N_908,N_1331);
and U2714 (N_2714,N_422,N_369);
and U2715 (N_2715,N_1623,N_1647);
nor U2716 (N_2716,N_1359,N_551);
xor U2717 (N_2717,N_1000,N_101);
xnor U2718 (N_2718,N_630,N_1604);
nor U2719 (N_2719,N_224,N_1055);
xnor U2720 (N_2720,N_617,N_829);
or U2721 (N_2721,N_282,N_1127);
xor U2722 (N_2722,N_266,N_353);
and U2723 (N_2723,N_1255,N_231);
nor U2724 (N_2724,N_1495,N_704);
or U2725 (N_2725,N_977,N_398);
xnor U2726 (N_2726,N_1873,N_1806);
and U2727 (N_2727,N_552,N_1358);
and U2728 (N_2728,N_1165,N_1737);
or U2729 (N_2729,N_882,N_631);
nand U2730 (N_2730,N_13,N_626);
and U2731 (N_2731,N_947,N_1392);
nor U2732 (N_2732,N_753,N_166);
nor U2733 (N_2733,N_1323,N_258);
nand U2734 (N_2734,N_727,N_944);
nand U2735 (N_2735,N_272,N_1846);
nor U2736 (N_2736,N_842,N_1936);
nor U2737 (N_2737,N_1921,N_846);
nor U2738 (N_2738,N_1059,N_1913);
xnor U2739 (N_2739,N_48,N_968);
and U2740 (N_2740,N_692,N_1803);
nor U2741 (N_2741,N_573,N_1335);
or U2742 (N_2742,N_720,N_1934);
or U2743 (N_2743,N_203,N_1510);
or U2744 (N_2744,N_386,N_1405);
or U2745 (N_2745,N_522,N_1381);
or U2746 (N_2746,N_1814,N_903);
xnor U2747 (N_2747,N_1150,N_1613);
and U2748 (N_2748,N_1428,N_568);
nand U2749 (N_2749,N_1692,N_519);
nor U2750 (N_2750,N_897,N_1106);
or U2751 (N_2751,N_1870,N_1943);
nand U2752 (N_2752,N_1822,N_1731);
xor U2753 (N_2753,N_1171,N_932);
or U2754 (N_2754,N_259,N_1740);
and U2755 (N_2755,N_410,N_1304);
xor U2756 (N_2756,N_628,N_1336);
nor U2757 (N_2757,N_1813,N_1845);
nor U2758 (N_2758,N_509,N_672);
nor U2759 (N_2759,N_135,N_804);
nor U2760 (N_2760,N_110,N_838);
or U2761 (N_2761,N_395,N_1619);
nand U2762 (N_2762,N_751,N_1441);
nand U2763 (N_2763,N_223,N_1685);
nand U2764 (N_2764,N_76,N_1831);
and U2765 (N_2765,N_1957,N_286);
nand U2766 (N_2766,N_371,N_1420);
xor U2767 (N_2767,N_1746,N_1033);
or U2768 (N_2768,N_517,N_206);
nor U2769 (N_2769,N_86,N_284);
and U2770 (N_2770,N_1917,N_538);
nand U2771 (N_2771,N_1497,N_1156);
nor U2772 (N_2772,N_1826,N_1802);
nor U2773 (N_2773,N_989,N_783);
xor U2774 (N_2774,N_1773,N_621);
nor U2775 (N_2775,N_57,N_1964);
or U2776 (N_2776,N_84,N_639);
and U2777 (N_2777,N_1277,N_682);
and U2778 (N_2778,N_1045,N_53);
xnor U2779 (N_2779,N_1210,N_220);
nand U2780 (N_2780,N_1152,N_214);
xnor U2781 (N_2781,N_1564,N_1010);
nand U2782 (N_2782,N_1111,N_1637);
xnor U2783 (N_2783,N_983,N_1220);
or U2784 (N_2784,N_333,N_1035);
or U2785 (N_2785,N_290,N_1879);
xnor U2786 (N_2786,N_1226,N_516);
nand U2787 (N_2787,N_1705,N_1505);
nor U2788 (N_2788,N_204,N_40);
nor U2789 (N_2789,N_82,N_855);
nor U2790 (N_2790,N_1052,N_494);
xor U2791 (N_2791,N_251,N_586);
nor U2792 (N_2792,N_1327,N_1351);
xor U2793 (N_2793,N_405,N_345);
nand U2794 (N_2794,N_1048,N_23);
or U2795 (N_2795,N_1125,N_487);
and U2796 (N_2796,N_170,N_1043);
nand U2797 (N_2797,N_596,N_1626);
nor U2798 (N_2798,N_1919,N_221);
and U2799 (N_2799,N_712,N_1282);
and U2800 (N_2800,N_167,N_1730);
or U2801 (N_2801,N_1299,N_664);
nand U2802 (N_2802,N_867,N_119);
or U2803 (N_2803,N_1372,N_1834);
nand U2804 (N_2804,N_1177,N_1615);
or U2805 (N_2805,N_1501,N_1143);
or U2806 (N_2806,N_1191,N_1520);
nand U2807 (N_2807,N_1393,N_1946);
xnor U2808 (N_2808,N_1205,N_1761);
and U2809 (N_2809,N_606,N_1807);
xor U2810 (N_2810,N_1151,N_1778);
xor U2811 (N_2811,N_403,N_1118);
nor U2812 (N_2812,N_454,N_1970);
nor U2813 (N_2813,N_1193,N_292);
and U2814 (N_2814,N_331,N_1691);
nor U2815 (N_2815,N_122,N_1075);
nor U2816 (N_2816,N_1368,N_576);
and U2817 (N_2817,N_515,N_1050);
xnor U2818 (N_2818,N_931,N_922);
xor U2819 (N_2819,N_228,N_1219);
nand U2820 (N_2820,N_985,N_125);
xnor U2821 (N_2821,N_1494,N_550);
nor U2822 (N_2822,N_338,N_1912);
nor U2823 (N_2823,N_1031,N_1657);
or U2824 (N_2824,N_1984,N_1350);
nand U2825 (N_2825,N_1283,N_942);
and U2826 (N_2826,N_1442,N_1811);
nor U2827 (N_2827,N_149,N_663);
and U2828 (N_2828,N_1201,N_1617);
nand U2829 (N_2829,N_448,N_1138);
xor U2830 (N_2830,N_1089,N_88);
or U2831 (N_2831,N_1458,N_1264);
and U2832 (N_2832,N_1867,N_900);
and U2833 (N_2833,N_106,N_1894);
nand U2834 (N_2834,N_601,N_1148);
nand U2835 (N_2835,N_1292,N_876);
nand U2836 (N_2836,N_1720,N_174);
and U2837 (N_2837,N_1459,N_782);
xnor U2838 (N_2838,N_697,N_1037);
nand U2839 (N_2839,N_1950,N_1280);
xor U2840 (N_2840,N_658,N_89);
nor U2841 (N_2841,N_1546,N_1759);
nand U2842 (N_2842,N_198,N_124);
and U2843 (N_2843,N_1348,N_1666);
and U2844 (N_2844,N_1126,N_1483);
or U2845 (N_2845,N_1693,N_102);
xnor U2846 (N_2846,N_1854,N_77);
xor U2847 (N_2847,N_1805,N_799);
or U2848 (N_2848,N_1409,N_427);
nand U2849 (N_2849,N_1842,N_246);
and U2850 (N_2850,N_1696,N_523);
and U2851 (N_2851,N_1732,N_811);
and U2852 (N_2852,N_1993,N_1411);
nand U2853 (N_2853,N_273,N_1961);
and U2854 (N_2854,N_892,N_33);
xnor U2855 (N_2855,N_918,N_683);
nand U2856 (N_2856,N_402,N_1355);
nor U2857 (N_2857,N_887,N_1663);
nor U2858 (N_2858,N_768,N_1958);
and U2859 (N_2859,N_330,N_400);
xor U2860 (N_2860,N_1829,N_961);
nor U2861 (N_2861,N_429,N_1550);
nor U2862 (N_2862,N_1416,N_478);
or U2863 (N_2863,N_917,N_716);
and U2864 (N_2864,N_978,N_616);
or U2865 (N_2865,N_610,N_502);
and U2866 (N_2866,N_390,N_1514);
or U2867 (N_2867,N_1543,N_671);
nor U2868 (N_2868,N_1423,N_208);
nand U2869 (N_2869,N_670,N_1952);
and U2870 (N_2870,N_1839,N_873);
nor U2871 (N_2871,N_1960,N_1291);
nor U2872 (N_2872,N_1408,N_1515);
and U2873 (N_2873,N_263,N_1851);
and U2874 (N_2874,N_1722,N_563);
or U2875 (N_2875,N_79,N_1145);
nor U2876 (N_2876,N_1332,N_285);
xor U2877 (N_2877,N_765,N_329);
nand U2878 (N_2878,N_703,N_153);
nand U2879 (N_2879,N_458,N_723);
or U2880 (N_2880,N_817,N_468);
and U2881 (N_2881,N_901,N_1697);
and U2882 (N_2882,N_476,N_1593);
xor U2883 (N_2883,N_466,N_67);
xnor U2884 (N_2884,N_139,N_1942);
nor U2885 (N_2885,N_861,N_1154);
or U2886 (N_2886,N_107,N_1830);
nor U2887 (N_2887,N_762,N_1858);
and U2888 (N_2888,N_685,N_624);
and U2889 (N_2889,N_1790,N_1764);
nor U2890 (N_2890,N_719,N_1823);
or U2891 (N_2891,N_1763,N_1548);
nand U2892 (N_2892,N_856,N_1911);
nor U2893 (N_2893,N_287,N_21);
or U2894 (N_2894,N_34,N_1530);
or U2895 (N_2895,N_1116,N_1624);
nand U2896 (N_2896,N_1256,N_1259);
and U2897 (N_2897,N_1651,N_300);
xor U2898 (N_2898,N_1212,N_787);
nor U2899 (N_2899,N_349,N_31);
or U2900 (N_2900,N_652,N_453);
nand U2901 (N_2901,N_230,N_136);
or U2902 (N_2902,N_1427,N_1856);
xor U2903 (N_2903,N_957,N_1038);
and U2904 (N_2904,N_795,N_721);
nor U2905 (N_2905,N_72,N_307);
xnor U2906 (N_2906,N_8,N_1664);
and U2907 (N_2907,N_1816,N_1962);
nand U2908 (N_2908,N_1868,N_1544);
nor U2909 (N_2909,N_839,N_1672);
nor U2910 (N_2910,N_889,N_1941);
and U2911 (N_2911,N_355,N_1360);
nor U2912 (N_2912,N_14,N_556);
nor U2913 (N_2913,N_1536,N_1747);
and U2914 (N_2914,N_1376,N_749);
nand U2915 (N_2915,N_1396,N_588);
and U2916 (N_2916,N_54,N_789);
nor U2917 (N_2917,N_1513,N_1346);
or U2918 (N_2918,N_647,N_1995);
xnor U2919 (N_2919,N_537,N_1094);
nand U2920 (N_2920,N_1243,N_777);
xor U2921 (N_2921,N_1456,N_1296);
nor U2922 (N_2922,N_1794,N_1726);
nor U2923 (N_2923,N_324,N_845);
or U2924 (N_2924,N_539,N_1656);
or U2925 (N_2925,N_528,N_1690);
and U2926 (N_2926,N_1784,N_1432);
nor U2927 (N_2927,N_486,N_281);
or U2928 (N_2928,N_1527,N_544);
nand U2929 (N_2929,N_1397,N_308);
or U2930 (N_2930,N_1072,N_559);
nor U2931 (N_2931,N_87,N_1357);
nor U2932 (N_2932,N_1321,N_1022);
nand U2933 (N_2933,N_1559,N_191);
xnor U2934 (N_2934,N_264,N_339);
nand U2935 (N_2935,N_1140,N_575);
nand U2936 (N_2936,N_569,N_1284);
nor U2937 (N_2937,N_344,N_1844);
xor U2938 (N_2938,N_1356,N_1751);
and U2939 (N_2939,N_1406,N_613);
nand U2940 (N_2940,N_301,N_350);
nor U2941 (N_2941,N_1333,N_71);
nor U2942 (N_2942,N_850,N_213);
nand U2943 (N_2943,N_1728,N_921);
nor U2944 (N_2944,N_118,N_998);
and U2945 (N_2945,N_713,N_662);
and U2946 (N_2946,N_1929,N_326);
xor U2947 (N_2947,N_1039,N_785);
xnor U2948 (N_2948,N_1774,N_354);
or U2949 (N_2949,N_1248,N_1541);
xnor U2950 (N_2950,N_380,N_1642);
or U2951 (N_2951,N_1976,N_129);
or U2952 (N_2952,N_678,N_1183);
or U2953 (N_2953,N_430,N_180);
or U2954 (N_2954,N_731,N_1237);
nor U2955 (N_2955,N_1025,N_358);
or U2956 (N_2956,N_1032,N_401);
or U2957 (N_2957,N_981,N_1390);
nor U2958 (N_2958,N_1295,N_788);
nand U2959 (N_2959,N_1078,N_1687);
nand U2960 (N_2960,N_747,N_1998);
nand U2961 (N_2961,N_212,N_1185);
nor U2962 (N_2962,N_449,N_1090);
xnor U2963 (N_2963,N_1289,N_366);
nor U2964 (N_2964,N_1837,N_830);
nand U2965 (N_2965,N_1288,N_1076);
xnor U2966 (N_2966,N_373,N_368);
nand U2967 (N_2967,N_1714,N_913);
xor U2968 (N_2968,N_58,N_315);
nor U2969 (N_2969,N_1018,N_1028);
nor U2970 (N_2970,N_1508,N_819);
or U2971 (N_2971,N_1361,N_1318);
nor U2972 (N_2972,N_1065,N_156);
nand U2973 (N_2973,N_217,N_459);
nand U2974 (N_2974,N_1521,N_1244);
xnor U2975 (N_2975,N_909,N_1721);
and U2976 (N_2976,N_1785,N_999);
and U2977 (N_2977,N_1036,N_1084);
nor U2978 (N_2978,N_334,N_834);
and U2979 (N_2979,N_384,N_923);
and U2980 (N_2980,N_1281,N_976);
xnor U2981 (N_2981,N_1978,N_1104);
nor U2982 (N_2982,N_379,N_437);
nor U2983 (N_2983,N_1315,N_1938);
and U2984 (N_2984,N_1251,N_1677);
or U2985 (N_2985,N_1188,N_1208);
xor U2986 (N_2986,N_252,N_3);
and U2987 (N_2987,N_1206,N_1134);
nor U2988 (N_2988,N_1146,N_866);
and U2989 (N_2989,N_529,N_1058);
nor U2990 (N_2990,N_1967,N_25);
or U2991 (N_2991,N_705,N_959);
xor U2992 (N_2992,N_1968,N_126);
and U2993 (N_2993,N_598,N_234);
and U2994 (N_2994,N_812,N_1982);
nand U2995 (N_2995,N_239,N_1989);
nand U2996 (N_2996,N_750,N_257);
xor U2997 (N_2997,N_717,N_1060);
xnor U2998 (N_2998,N_1034,N_1948);
nand U2999 (N_2999,N_1862,N_1041);
nor U3000 (N_3000,N_494,N_371);
xnor U3001 (N_3001,N_763,N_1308);
or U3002 (N_3002,N_630,N_1591);
nor U3003 (N_3003,N_548,N_761);
nand U3004 (N_3004,N_876,N_1144);
and U3005 (N_3005,N_1671,N_764);
xor U3006 (N_3006,N_593,N_295);
nor U3007 (N_3007,N_907,N_1747);
nand U3008 (N_3008,N_1501,N_773);
xnor U3009 (N_3009,N_135,N_80);
and U3010 (N_3010,N_1273,N_1554);
nor U3011 (N_3011,N_1994,N_322);
xor U3012 (N_3012,N_793,N_1612);
or U3013 (N_3013,N_1707,N_1917);
nor U3014 (N_3014,N_702,N_871);
nand U3015 (N_3015,N_182,N_869);
xor U3016 (N_3016,N_117,N_509);
nor U3017 (N_3017,N_75,N_1922);
and U3018 (N_3018,N_1962,N_1843);
or U3019 (N_3019,N_767,N_1637);
nor U3020 (N_3020,N_1866,N_1230);
or U3021 (N_3021,N_449,N_663);
nand U3022 (N_3022,N_1642,N_312);
xor U3023 (N_3023,N_255,N_1918);
nand U3024 (N_3024,N_1448,N_875);
nand U3025 (N_3025,N_1518,N_157);
or U3026 (N_3026,N_1417,N_1831);
nor U3027 (N_3027,N_1611,N_1842);
nand U3028 (N_3028,N_651,N_777);
nand U3029 (N_3029,N_1319,N_1512);
and U3030 (N_3030,N_1500,N_867);
or U3031 (N_3031,N_1315,N_683);
nor U3032 (N_3032,N_479,N_1573);
nor U3033 (N_3033,N_751,N_1920);
and U3034 (N_3034,N_11,N_796);
xor U3035 (N_3035,N_1092,N_1426);
nor U3036 (N_3036,N_1925,N_785);
and U3037 (N_3037,N_164,N_1204);
nor U3038 (N_3038,N_261,N_888);
xor U3039 (N_3039,N_1299,N_1518);
nand U3040 (N_3040,N_121,N_1837);
nor U3041 (N_3041,N_1909,N_209);
xor U3042 (N_3042,N_198,N_932);
or U3043 (N_3043,N_648,N_1217);
or U3044 (N_3044,N_1267,N_190);
xor U3045 (N_3045,N_664,N_50);
or U3046 (N_3046,N_1943,N_860);
nor U3047 (N_3047,N_693,N_1972);
xnor U3048 (N_3048,N_1746,N_1010);
or U3049 (N_3049,N_912,N_1094);
or U3050 (N_3050,N_587,N_484);
or U3051 (N_3051,N_1599,N_1435);
xnor U3052 (N_3052,N_1430,N_382);
and U3053 (N_3053,N_15,N_393);
xnor U3054 (N_3054,N_293,N_375);
nand U3055 (N_3055,N_1069,N_1190);
or U3056 (N_3056,N_394,N_1817);
or U3057 (N_3057,N_805,N_216);
or U3058 (N_3058,N_1449,N_182);
and U3059 (N_3059,N_320,N_991);
nand U3060 (N_3060,N_507,N_1798);
and U3061 (N_3061,N_1768,N_910);
nand U3062 (N_3062,N_1904,N_723);
or U3063 (N_3063,N_928,N_459);
xor U3064 (N_3064,N_225,N_1160);
and U3065 (N_3065,N_869,N_303);
and U3066 (N_3066,N_1802,N_56);
or U3067 (N_3067,N_1162,N_813);
or U3068 (N_3068,N_1878,N_1044);
or U3069 (N_3069,N_633,N_1685);
nor U3070 (N_3070,N_676,N_780);
nand U3071 (N_3071,N_1583,N_75);
nand U3072 (N_3072,N_1919,N_797);
and U3073 (N_3073,N_1477,N_517);
nor U3074 (N_3074,N_1964,N_1786);
and U3075 (N_3075,N_1650,N_1891);
and U3076 (N_3076,N_164,N_700);
nand U3077 (N_3077,N_1009,N_1984);
nor U3078 (N_3078,N_1996,N_612);
and U3079 (N_3079,N_1183,N_1127);
xnor U3080 (N_3080,N_409,N_1811);
xnor U3081 (N_3081,N_151,N_769);
nor U3082 (N_3082,N_586,N_1759);
xnor U3083 (N_3083,N_1050,N_1423);
nand U3084 (N_3084,N_1795,N_984);
nor U3085 (N_3085,N_1675,N_1586);
nand U3086 (N_3086,N_1525,N_1020);
nand U3087 (N_3087,N_1905,N_588);
and U3088 (N_3088,N_1422,N_730);
nor U3089 (N_3089,N_1633,N_171);
xor U3090 (N_3090,N_468,N_1128);
or U3091 (N_3091,N_1814,N_1556);
and U3092 (N_3092,N_1963,N_608);
xnor U3093 (N_3093,N_772,N_1046);
nor U3094 (N_3094,N_647,N_1340);
and U3095 (N_3095,N_1659,N_1279);
xor U3096 (N_3096,N_1240,N_1373);
nor U3097 (N_3097,N_277,N_1192);
nand U3098 (N_3098,N_795,N_1544);
nor U3099 (N_3099,N_1143,N_1403);
nand U3100 (N_3100,N_7,N_1541);
nand U3101 (N_3101,N_737,N_64);
and U3102 (N_3102,N_1892,N_1156);
and U3103 (N_3103,N_1165,N_1320);
nand U3104 (N_3104,N_1213,N_1498);
and U3105 (N_3105,N_581,N_936);
or U3106 (N_3106,N_432,N_1016);
and U3107 (N_3107,N_1799,N_1055);
nor U3108 (N_3108,N_714,N_352);
nor U3109 (N_3109,N_1912,N_1818);
nor U3110 (N_3110,N_489,N_1108);
nor U3111 (N_3111,N_1527,N_796);
nand U3112 (N_3112,N_6,N_1741);
nand U3113 (N_3113,N_928,N_1151);
nand U3114 (N_3114,N_538,N_1088);
nor U3115 (N_3115,N_1493,N_1159);
and U3116 (N_3116,N_4,N_936);
nand U3117 (N_3117,N_1364,N_136);
and U3118 (N_3118,N_579,N_1860);
xor U3119 (N_3119,N_1611,N_604);
nand U3120 (N_3120,N_490,N_1626);
xnor U3121 (N_3121,N_1021,N_42);
nor U3122 (N_3122,N_148,N_814);
nand U3123 (N_3123,N_1072,N_783);
or U3124 (N_3124,N_1157,N_108);
nand U3125 (N_3125,N_1708,N_711);
and U3126 (N_3126,N_1175,N_501);
xnor U3127 (N_3127,N_1173,N_347);
nor U3128 (N_3128,N_977,N_516);
nand U3129 (N_3129,N_47,N_692);
and U3130 (N_3130,N_559,N_977);
and U3131 (N_3131,N_660,N_1194);
nand U3132 (N_3132,N_789,N_1197);
and U3133 (N_3133,N_949,N_192);
nand U3134 (N_3134,N_491,N_1689);
nor U3135 (N_3135,N_1118,N_1866);
and U3136 (N_3136,N_1656,N_1728);
xnor U3137 (N_3137,N_816,N_1727);
nor U3138 (N_3138,N_1498,N_488);
and U3139 (N_3139,N_536,N_1039);
xor U3140 (N_3140,N_263,N_295);
xor U3141 (N_3141,N_1298,N_1371);
xor U3142 (N_3142,N_1293,N_978);
xnor U3143 (N_3143,N_1122,N_526);
nor U3144 (N_3144,N_901,N_811);
or U3145 (N_3145,N_1017,N_1868);
nor U3146 (N_3146,N_13,N_1383);
nand U3147 (N_3147,N_1723,N_1830);
or U3148 (N_3148,N_1885,N_1992);
nor U3149 (N_3149,N_1106,N_845);
and U3150 (N_3150,N_1816,N_925);
or U3151 (N_3151,N_809,N_1120);
nor U3152 (N_3152,N_442,N_621);
or U3153 (N_3153,N_418,N_1426);
xor U3154 (N_3154,N_728,N_84);
and U3155 (N_3155,N_1468,N_1750);
and U3156 (N_3156,N_1404,N_62);
and U3157 (N_3157,N_725,N_844);
xor U3158 (N_3158,N_940,N_1750);
nor U3159 (N_3159,N_351,N_1939);
nor U3160 (N_3160,N_1993,N_1096);
nand U3161 (N_3161,N_734,N_1453);
xor U3162 (N_3162,N_998,N_1416);
nand U3163 (N_3163,N_1538,N_363);
xnor U3164 (N_3164,N_975,N_1943);
and U3165 (N_3165,N_24,N_859);
nor U3166 (N_3166,N_1240,N_671);
nand U3167 (N_3167,N_1613,N_1441);
or U3168 (N_3168,N_1613,N_376);
xor U3169 (N_3169,N_237,N_1360);
nand U3170 (N_3170,N_790,N_158);
xor U3171 (N_3171,N_635,N_155);
nor U3172 (N_3172,N_1961,N_443);
xnor U3173 (N_3173,N_566,N_151);
xor U3174 (N_3174,N_127,N_508);
nor U3175 (N_3175,N_1757,N_1658);
xor U3176 (N_3176,N_1480,N_707);
nand U3177 (N_3177,N_1673,N_930);
xor U3178 (N_3178,N_433,N_1230);
nand U3179 (N_3179,N_1345,N_256);
nand U3180 (N_3180,N_1531,N_1394);
or U3181 (N_3181,N_672,N_1204);
nor U3182 (N_3182,N_1275,N_911);
nand U3183 (N_3183,N_1207,N_1149);
and U3184 (N_3184,N_1054,N_1013);
and U3185 (N_3185,N_1776,N_799);
and U3186 (N_3186,N_1482,N_399);
nor U3187 (N_3187,N_1882,N_131);
and U3188 (N_3188,N_392,N_891);
nand U3189 (N_3189,N_978,N_1985);
nand U3190 (N_3190,N_765,N_896);
and U3191 (N_3191,N_1002,N_1306);
nand U3192 (N_3192,N_1162,N_680);
xor U3193 (N_3193,N_827,N_904);
xor U3194 (N_3194,N_669,N_377);
nor U3195 (N_3195,N_1258,N_130);
nand U3196 (N_3196,N_944,N_1618);
nand U3197 (N_3197,N_1398,N_424);
or U3198 (N_3198,N_1311,N_985);
nor U3199 (N_3199,N_1279,N_692);
nand U3200 (N_3200,N_1953,N_266);
and U3201 (N_3201,N_1793,N_1743);
and U3202 (N_3202,N_960,N_356);
nand U3203 (N_3203,N_682,N_670);
nor U3204 (N_3204,N_1581,N_334);
xor U3205 (N_3205,N_1049,N_1221);
and U3206 (N_3206,N_432,N_1964);
nor U3207 (N_3207,N_971,N_737);
and U3208 (N_3208,N_886,N_109);
nor U3209 (N_3209,N_266,N_542);
nand U3210 (N_3210,N_1850,N_1698);
xor U3211 (N_3211,N_1383,N_330);
nand U3212 (N_3212,N_1573,N_242);
nand U3213 (N_3213,N_999,N_154);
or U3214 (N_3214,N_827,N_859);
and U3215 (N_3215,N_1605,N_1842);
and U3216 (N_3216,N_1548,N_1355);
nand U3217 (N_3217,N_941,N_691);
nor U3218 (N_3218,N_419,N_836);
xor U3219 (N_3219,N_1814,N_1020);
or U3220 (N_3220,N_1778,N_968);
xnor U3221 (N_3221,N_1306,N_401);
or U3222 (N_3222,N_1880,N_1728);
nand U3223 (N_3223,N_1240,N_1664);
xor U3224 (N_3224,N_176,N_784);
and U3225 (N_3225,N_804,N_314);
or U3226 (N_3226,N_1398,N_557);
nor U3227 (N_3227,N_1757,N_1066);
nor U3228 (N_3228,N_992,N_640);
or U3229 (N_3229,N_1667,N_22);
nor U3230 (N_3230,N_1561,N_1595);
or U3231 (N_3231,N_1562,N_1952);
xnor U3232 (N_3232,N_693,N_1470);
and U3233 (N_3233,N_302,N_689);
and U3234 (N_3234,N_1113,N_1054);
nor U3235 (N_3235,N_1704,N_1061);
and U3236 (N_3236,N_1932,N_1838);
nand U3237 (N_3237,N_1081,N_791);
xor U3238 (N_3238,N_256,N_702);
xor U3239 (N_3239,N_1544,N_1390);
nor U3240 (N_3240,N_460,N_1786);
nand U3241 (N_3241,N_786,N_608);
xor U3242 (N_3242,N_1019,N_85);
and U3243 (N_3243,N_959,N_1154);
xor U3244 (N_3244,N_106,N_1153);
nand U3245 (N_3245,N_364,N_1398);
or U3246 (N_3246,N_479,N_57);
nand U3247 (N_3247,N_360,N_231);
or U3248 (N_3248,N_338,N_451);
or U3249 (N_3249,N_74,N_953);
or U3250 (N_3250,N_396,N_1416);
nor U3251 (N_3251,N_1598,N_350);
or U3252 (N_3252,N_799,N_1232);
and U3253 (N_3253,N_1829,N_863);
nand U3254 (N_3254,N_273,N_1754);
xor U3255 (N_3255,N_1616,N_548);
nor U3256 (N_3256,N_988,N_1453);
or U3257 (N_3257,N_1845,N_617);
xnor U3258 (N_3258,N_919,N_1616);
nor U3259 (N_3259,N_1865,N_1708);
nand U3260 (N_3260,N_66,N_1757);
xnor U3261 (N_3261,N_245,N_599);
or U3262 (N_3262,N_1255,N_1586);
xor U3263 (N_3263,N_1768,N_281);
xnor U3264 (N_3264,N_1560,N_1435);
or U3265 (N_3265,N_328,N_835);
and U3266 (N_3266,N_705,N_783);
nand U3267 (N_3267,N_530,N_495);
and U3268 (N_3268,N_1957,N_931);
xor U3269 (N_3269,N_905,N_136);
or U3270 (N_3270,N_670,N_651);
xor U3271 (N_3271,N_528,N_474);
nand U3272 (N_3272,N_750,N_955);
and U3273 (N_3273,N_1071,N_222);
or U3274 (N_3274,N_1017,N_1066);
and U3275 (N_3275,N_1305,N_1115);
or U3276 (N_3276,N_1136,N_1969);
nor U3277 (N_3277,N_957,N_767);
or U3278 (N_3278,N_1582,N_311);
xor U3279 (N_3279,N_957,N_1867);
xnor U3280 (N_3280,N_658,N_239);
or U3281 (N_3281,N_442,N_503);
xor U3282 (N_3282,N_970,N_1075);
nand U3283 (N_3283,N_78,N_1662);
nand U3284 (N_3284,N_391,N_1033);
nand U3285 (N_3285,N_1038,N_1631);
and U3286 (N_3286,N_1023,N_1702);
nor U3287 (N_3287,N_1160,N_1317);
nor U3288 (N_3288,N_939,N_343);
xor U3289 (N_3289,N_954,N_202);
and U3290 (N_3290,N_620,N_1197);
nor U3291 (N_3291,N_1608,N_217);
xnor U3292 (N_3292,N_1943,N_968);
or U3293 (N_3293,N_1638,N_387);
xnor U3294 (N_3294,N_476,N_762);
xnor U3295 (N_3295,N_1469,N_1412);
nor U3296 (N_3296,N_169,N_252);
or U3297 (N_3297,N_485,N_473);
and U3298 (N_3298,N_1716,N_1527);
and U3299 (N_3299,N_1506,N_404);
and U3300 (N_3300,N_334,N_278);
xnor U3301 (N_3301,N_964,N_412);
nor U3302 (N_3302,N_1088,N_1617);
or U3303 (N_3303,N_96,N_1843);
xor U3304 (N_3304,N_1121,N_1836);
xnor U3305 (N_3305,N_1370,N_891);
and U3306 (N_3306,N_333,N_1415);
nand U3307 (N_3307,N_1483,N_318);
xor U3308 (N_3308,N_1064,N_1698);
xnor U3309 (N_3309,N_1786,N_1639);
xor U3310 (N_3310,N_1564,N_694);
xnor U3311 (N_3311,N_1841,N_752);
and U3312 (N_3312,N_951,N_526);
or U3313 (N_3313,N_1192,N_1510);
nand U3314 (N_3314,N_30,N_1501);
nand U3315 (N_3315,N_885,N_1335);
nand U3316 (N_3316,N_542,N_582);
nor U3317 (N_3317,N_612,N_1999);
nand U3318 (N_3318,N_795,N_1083);
nand U3319 (N_3319,N_1955,N_35);
or U3320 (N_3320,N_39,N_1773);
or U3321 (N_3321,N_1478,N_1034);
or U3322 (N_3322,N_599,N_1291);
xnor U3323 (N_3323,N_861,N_1972);
and U3324 (N_3324,N_1536,N_216);
and U3325 (N_3325,N_1166,N_355);
nand U3326 (N_3326,N_420,N_252);
or U3327 (N_3327,N_924,N_1774);
nor U3328 (N_3328,N_263,N_539);
or U3329 (N_3329,N_1710,N_1696);
or U3330 (N_3330,N_1374,N_250);
nand U3331 (N_3331,N_1383,N_133);
nor U3332 (N_3332,N_1364,N_845);
or U3333 (N_3333,N_562,N_518);
nor U3334 (N_3334,N_1991,N_761);
nand U3335 (N_3335,N_1103,N_1213);
and U3336 (N_3336,N_1740,N_104);
nand U3337 (N_3337,N_485,N_1547);
nor U3338 (N_3338,N_1351,N_1015);
nor U3339 (N_3339,N_1061,N_83);
xor U3340 (N_3340,N_1980,N_444);
xnor U3341 (N_3341,N_1458,N_978);
or U3342 (N_3342,N_348,N_1470);
or U3343 (N_3343,N_278,N_1655);
xnor U3344 (N_3344,N_1761,N_955);
xnor U3345 (N_3345,N_1907,N_1109);
nand U3346 (N_3346,N_559,N_1002);
nand U3347 (N_3347,N_1057,N_1511);
and U3348 (N_3348,N_987,N_1539);
nand U3349 (N_3349,N_623,N_676);
nand U3350 (N_3350,N_1984,N_55);
xor U3351 (N_3351,N_717,N_967);
or U3352 (N_3352,N_1304,N_1107);
nand U3353 (N_3353,N_213,N_903);
and U3354 (N_3354,N_37,N_1209);
and U3355 (N_3355,N_378,N_386);
xnor U3356 (N_3356,N_1209,N_683);
nor U3357 (N_3357,N_724,N_139);
nor U3358 (N_3358,N_336,N_1757);
and U3359 (N_3359,N_1991,N_479);
and U3360 (N_3360,N_999,N_420);
nand U3361 (N_3361,N_1318,N_1673);
and U3362 (N_3362,N_940,N_1211);
and U3363 (N_3363,N_744,N_517);
nand U3364 (N_3364,N_1435,N_426);
nor U3365 (N_3365,N_310,N_594);
and U3366 (N_3366,N_505,N_363);
xor U3367 (N_3367,N_911,N_1817);
nand U3368 (N_3368,N_502,N_1971);
or U3369 (N_3369,N_865,N_1574);
nand U3370 (N_3370,N_952,N_561);
nand U3371 (N_3371,N_926,N_1694);
nor U3372 (N_3372,N_592,N_201);
and U3373 (N_3373,N_969,N_707);
xor U3374 (N_3374,N_1663,N_1443);
or U3375 (N_3375,N_434,N_1945);
and U3376 (N_3376,N_1662,N_1289);
nor U3377 (N_3377,N_604,N_755);
or U3378 (N_3378,N_1488,N_702);
nand U3379 (N_3379,N_237,N_946);
or U3380 (N_3380,N_847,N_1657);
nand U3381 (N_3381,N_499,N_1524);
nor U3382 (N_3382,N_1754,N_844);
and U3383 (N_3383,N_1654,N_942);
nand U3384 (N_3384,N_1750,N_1701);
nor U3385 (N_3385,N_1599,N_1766);
and U3386 (N_3386,N_1191,N_746);
or U3387 (N_3387,N_345,N_95);
or U3388 (N_3388,N_1465,N_561);
and U3389 (N_3389,N_1785,N_1056);
nor U3390 (N_3390,N_1514,N_603);
xnor U3391 (N_3391,N_1921,N_1188);
xnor U3392 (N_3392,N_132,N_530);
xnor U3393 (N_3393,N_461,N_883);
xnor U3394 (N_3394,N_1819,N_780);
and U3395 (N_3395,N_1760,N_10);
xor U3396 (N_3396,N_293,N_1166);
and U3397 (N_3397,N_738,N_1833);
and U3398 (N_3398,N_1356,N_13);
nand U3399 (N_3399,N_658,N_1369);
or U3400 (N_3400,N_445,N_1609);
or U3401 (N_3401,N_588,N_378);
xor U3402 (N_3402,N_1152,N_1838);
nor U3403 (N_3403,N_1032,N_1167);
nor U3404 (N_3404,N_1762,N_1385);
xnor U3405 (N_3405,N_379,N_596);
nor U3406 (N_3406,N_1005,N_1228);
nor U3407 (N_3407,N_1708,N_1069);
and U3408 (N_3408,N_1489,N_933);
and U3409 (N_3409,N_1938,N_1738);
and U3410 (N_3410,N_1970,N_1675);
or U3411 (N_3411,N_1225,N_1101);
or U3412 (N_3412,N_99,N_1496);
or U3413 (N_3413,N_1443,N_1217);
and U3414 (N_3414,N_856,N_1496);
nor U3415 (N_3415,N_1683,N_486);
or U3416 (N_3416,N_210,N_358);
nor U3417 (N_3417,N_534,N_715);
and U3418 (N_3418,N_1994,N_491);
nor U3419 (N_3419,N_1289,N_463);
or U3420 (N_3420,N_1682,N_386);
and U3421 (N_3421,N_1111,N_1236);
nor U3422 (N_3422,N_1729,N_985);
and U3423 (N_3423,N_1596,N_900);
nand U3424 (N_3424,N_187,N_743);
nor U3425 (N_3425,N_121,N_372);
nand U3426 (N_3426,N_1013,N_1139);
or U3427 (N_3427,N_687,N_1063);
nand U3428 (N_3428,N_1981,N_1783);
nand U3429 (N_3429,N_1705,N_785);
or U3430 (N_3430,N_275,N_428);
or U3431 (N_3431,N_1526,N_1568);
nor U3432 (N_3432,N_669,N_1226);
or U3433 (N_3433,N_1512,N_523);
nor U3434 (N_3434,N_1334,N_774);
nor U3435 (N_3435,N_346,N_157);
and U3436 (N_3436,N_1877,N_1341);
xor U3437 (N_3437,N_1063,N_812);
and U3438 (N_3438,N_749,N_1681);
and U3439 (N_3439,N_655,N_490);
or U3440 (N_3440,N_1445,N_1226);
nor U3441 (N_3441,N_960,N_953);
nand U3442 (N_3442,N_179,N_98);
nand U3443 (N_3443,N_771,N_544);
or U3444 (N_3444,N_930,N_396);
nor U3445 (N_3445,N_1565,N_1505);
xnor U3446 (N_3446,N_1876,N_1536);
nor U3447 (N_3447,N_1923,N_1319);
xor U3448 (N_3448,N_960,N_708);
nor U3449 (N_3449,N_390,N_12);
nand U3450 (N_3450,N_1244,N_946);
or U3451 (N_3451,N_783,N_50);
nand U3452 (N_3452,N_1249,N_1188);
and U3453 (N_3453,N_458,N_493);
nor U3454 (N_3454,N_1989,N_1188);
and U3455 (N_3455,N_1911,N_578);
or U3456 (N_3456,N_321,N_364);
and U3457 (N_3457,N_1858,N_1731);
or U3458 (N_3458,N_1417,N_1204);
xnor U3459 (N_3459,N_828,N_1102);
or U3460 (N_3460,N_1077,N_1960);
nor U3461 (N_3461,N_1084,N_774);
xnor U3462 (N_3462,N_1012,N_1371);
xor U3463 (N_3463,N_1344,N_1856);
or U3464 (N_3464,N_1408,N_1636);
nand U3465 (N_3465,N_1663,N_1149);
and U3466 (N_3466,N_197,N_439);
and U3467 (N_3467,N_425,N_1469);
and U3468 (N_3468,N_644,N_1136);
nand U3469 (N_3469,N_899,N_180);
or U3470 (N_3470,N_150,N_1562);
nand U3471 (N_3471,N_931,N_1782);
nand U3472 (N_3472,N_1373,N_632);
nand U3473 (N_3473,N_1841,N_1964);
or U3474 (N_3474,N_1129,N_1879);
nand U3475 (N_3475,N_1536,N_977);
or U3476 (N_3476,N_993,N_199);
xnor U3477 (N_3477,N_1144,N_563);
nand U3478 (N_3478,N_1284,N_474);
xor U3479 (N_3479,N_1836,N_204);
or U3480 (N_3480,N_1778,N_1030);
xnor U3481 (N_3481,N_801,N_1729);
xnor U3482 (N_3482,N_919,N_1054);
nor U3483 (N_3483,N_1336,N_477);
and U3484 (N_3484,N_1433,N_942);
nand U3485 (N_3485,N_638,N_856);
or U3486 (N_3486,N_899,N_1732);
and U3487 (N_3487,N_219,N_847);
nand U3488 (N_3488,N_1215,N_1328);
xnor U3489 (N_3489,N_301,N_1259);
nand U3490 (N_3490,N_697,N_858);
xor U3491 (N_3491,N_1384,N_972);
nand U3492 (N_3492,N_1598,N_1625);
nand U3493 (N_3493,N_1774,N_1168);
nor U3494 (N_3494,N_1748,N_38);
or U3495 (N_3495,N_1896,N_186);
xor U3496 (N_3496,N_989,N_305);
nand U3497 (N_3497,N_386,N_1667);
and U3498 (N_3498,N_1777,N_1589);
nand U3499 (N_3499,N_1760,N_286);
nand U3500 (N_3500,N_800,N_1590);
nand U3501 (N_3501,N_374,N_1877);
nand U3502 (N_3502,N_166,N_1019);
or U3503 (N_3503,N_1745,N_513);
nor U3504 (N_3504,N_1206,N_1408);
nand U3505 (N_3505,N_354,N_1610);
nand U3506 (N_3506,N_496,N_26);
or U3507 (N_3507,N_1840,N_1957);
or U3508 (N_3508,N_274,N_1302);
nor U3509 (N_3509,N_1642,N_595);
or U3510 (N_3510,N_303,N_43);
nor U3511 (N_3511,N_172,N_1779);
xnor U3512 (N_3512,N_1624,N_692);
nand U3513 (N_3513,N_1259,N_1419);
xnor U3514 (N_3514,N_949,N_1491);
nand U3515 (N_3515,N_1497,N_202);
and U3516 (N_3516,N_1463,N_1309);
nor U3517 (N_3517,N_1875,N_1420);
or U3518 (N_3518,N_455,N_1711);
xor U3519 (N_3519,N_1873,N_1684);
nor U3520 (N_3520,N_313,N_1796);
nand U3521 (N_3521,N_1322,N_946);
xor U3522 (N_3522,N_1896,N_744);
xnor U3523 (N_3523,N_385,N_1646);
xnor U3524 (N_3524,N_1062,N_940);
nand U3525 (N_3525,N_550,N_598);
and U3526 (N_3526,N_161,N_647);
or U3527 (N_3527,N_1247,N_1939);
nand U3528 (N_3528,N_1529,N_899);
and U3529 (N_3529,N_585,N_1758);
and U3530 (N_3530,N_285,N_597);
xnor U3531 (N_3531,N_1257,N_1218);
nand U3532 (N_3532,N_1786,N_393);
and U3533 (N_3533,N_1980,N_145);
xnor U3534 (N_3534,N_204,N_624);
nor U3535 (N_3535,N_849,N_1279);
xor U3536 (N_3536,N_929,N_893);
xnor U3537 (N_3537,N_413,N_328);
or U3538 (N_3538,N_1795,N_846);
nor U3539 (N_3539,N_155,N_669);
nor U3540 (N_3540,N_1084,N_1853);
and U3541 (N_3541,N_1772,N_1188);
nand U3542 (N_3542,N_1066,N_1809);
nor U3543 (N_3543,N_820,N_1750);
or U3544 (N_3544,N_392,N_814);
xnor U3545 (N_3545,N_1081,N_1553);
or U3546 (N_3546,N_1629,N_1599);
or U3547 (N_3547,N_164,N_1982);
nand U3548 (N_3548,N_56,N_18);
xnor U3549 (N_3549,N_1303,N_1107);
nand U3550 (N_3550,N_281,N_1080);
nor U3551 (N_3551,N_1268,N_1774);
xor U3552 (N_3552,N_404,N_1701);
nor U3553 (N_3553,N_1714,N_810);
and U3554 (N_3554,N_1665,N_686);
nor U3555 (N_3555,N_451,N_1662);
xnor U3556 (N_3556,N_825,N_444);
nor U3557 (N_3557,N_1205,N_942);
xnor U3558 (N_3558,N_1527,N_1206);
and U3559 (N_3559,N_333,N_1991);
or U3560 (N_3560,N_199,N_1127);
nor U3561 (N_3561,N_647,N_417);
and U3562 (N_3562,N_1943,N_1365);
nand U3563 (N_3563,N_1023,N_953);
or U3564 (N_3564,N_1637,N_406);
nand U3565 (N_3565,N_134,N_409);
nand U3566 (N_3566,N_1200,N_1503);
nand U3567 (N_3567,N_812,N_1816);
nand U3568 (N_3568,N_713,N_397);
and U3569 (N_3569,N_1776,N_376);
or U3570 (N_3570,N_1939,N_1799);
nor U3571 (N_3571,N_684,N_442);
nand U3572 (N_3572,N_1767,N_1666);
and U3573 (N_3573,N_170,N_1311);
nor U3574 (N_3574,N_1043,N_317);
xor U3575 (N_3575,N_204,N_267);
and U3576 (N_3576,N_1046,N_1704);
or U3577 (N_3577,N_535,N_195);
and U3578 (N_3578,N_462,N_1596);
nand U3579 (N_3579,N_479,N_70);
or U3580 (N_3580,N_1908,N_1652);
xnor U3581 (N_3581,N_552,N_1770);
nand U3582 (N_3582,N_333,N_1221);
and U3583 (N_3583,N_1252,N_565);
and U3584 (N_3584,N_1566,N_1881);
nand U3585 (N_3585,N_138,N_719);
nand U3586 (N_3586,N_27,N_195);
and U3587 (N_3587,N_34,N_764);
nor U3588 (N_3588,N_1236,N_1133);
xor U3589 (N_3589,N_983,N_1969);
or U3590 (N_3590,N_787,N_1842);
and U3591 (N_3591,N_623,N_198);
nand U3592 (N_3592,N_642,N_1926);
or U3593 (N_3593,N_1456,N_893);
and U3594 (N_3594,N_1341,N_1769);
xnor U3595 (N_3595,N_538,N_1799);
xor U3596 (N_3596,N_521,N_1697);
nand U3597 (N_3597,N_54,N_1955);
nand U3598 (N_3598,N_11,N_461);
and U3599 (N_3599,N_943,N_896);
or U3600 (N_3600,N_1957,N_1602);
nor U3601 (N_3601,N_734,N_1525);
xor U3602 (N_3602,N_1383,N_1726);
or U3603 (N_3603,N_1055,N_356);
nor U3604 (N_3604,N_1372,N_1200);
nand U3605 (N_3605,N_886,N_238);
and U3606 (N_3606,N_106,N_1052);
and U3607 (N_3607,N_725,N_1716);
and U3608 (N_3608,N_1713,N_1783);
or U3609 (N_3609,N_1594,N_165);
xnor U3610 (N_3610,N_1139,N_1882);
nor U3611 (N_3611,N_195,N_878);
nor U3612 (N_3612,N_1240,N_909);
nor U3613 (N_3613,N_726,N_1084);
or U3614 (N_3614,N_606,N_51);
or U3615 (N_3615,N_6,N_16);
nand U3616 (N_3616,N_851,N_1774);
nand U3617 (N_3617,N_1866,N_1227);
or U3618 (N_3618,N_1266,N_39);
xor U3619 (N_3619,N_860,N_1913);
xnor U3620 (N_3620,N_1162,N_740);
xor U3621 (N_3621,N_1344,N_396);
xnor U3622 (N_3622,N_1519,N_239);
nand U3623 (N_3623,N_569,N_1330);
nor U3624 (N_3624,N_501,N_829);
and U3625 (N_3625,N_941,N_875);
and U3626 (N_3626,N_736,N_616);
nor U3627 (N_3627,N_546,N_1993);
and U3628 (N_3628,N_1458,N_786);
nand U3629 (N_3629,N_1318,N_814);
xor U3630 (N_3630,N_1300,N_961);
nand U3631 (N_3631,N_770,N_1091);
nor U3632 (N_3632,N_1015,N_1677);
xnor U3633 (N_3633,N_844,N_481);
nand U3634 (N_3634,N_484,N_1685);
xor U3635 (N_3635,N_1011,N_1190);
nor U3636 (N_3636,N_1821,N_236);
nor U3637 (N_3637,N_1582,N_1111);
and U3638 (N_3638,N_225,N_1672);
xnor U3639 (N_3639,N_1637,N_1089);
nor U3640 (N_3640,N_1465,N_812);
xnor U3641 (N_3641,N_321,N_1945);
or U3642 (N_3642,N_647,N_1035);
or U3643 (N_3643,N_957,N_991);
xor U3644 (N_3644,N_398,N_1263);
nor U3645 (N_3645,N_1800,N_1389);
nor U3646 (N_3646,N_1421,N_1563);
and U3647 (N_3647,N_242,N_218);
or U3648 (N_3648,N_862,N_37);
and U3649 (N_3649,N_453,N_5);
or U3650 (N_3650,N_1038,N_242);
nand U3651 (N_3651,N_210,N_684);
or U3652 (N_3652,N_1988,N_1634);
or U3653 (N_3653,N_120,N_559);
xnor U3654 (N_3654,N_440,N_1788);
or U3655 (N_3655,N_832,N_928);
xor U3656 (N_3656,N_1363,N_1139);
nand U3657 (N_3657,N_1281,N_437);
xnor U3658 (N_3658,N_410,N_821);
nor U3659 (N_3659,N_809,N_111);
nand U3660 (N_3660,N_1576,N_1321);
or U3661 (N_3661,N_997,N_23);
nand U3662 (N_3662,N_1797,N_1074);
or U3663 (N_3663,N_1968,N_698);
nand U3664 (N_3664,N_451,N_1984);
and U3665 (N_3665,N_979,N_1899);
nor U3666 (N_3666,N_188,N_564);
nand U3667 (N_3667,N_34,N_1764);
nand U3668 (N_3668,N_1500,N_1499);
nor U3669 (N_3669,N_1381,N_785);
xor U3670 (N_3670,N_965,N_687);
and U3671 (N_3671,N_1666,N_1796);
or U3672 (N_3672,N_266,N_1731);
nor U3673 (N_3673,N_263,N_825);
nor U3674 (N_3674,N_1346,N_1831);
and U3675 (N_3675,N_227,N_439);
nor U3676 (N_3676,N_1002,N_1189);
nand U3677 (N_3677,N_470,N_1829);
nand U3678 (N_3678,N_905,N_1939);
nor U3679 (N_3679,N_1548,N_501);
nor U3680 (N_3680,N_296,N_1746);
or U3681 (N_3681,N_155,N_1982);
nor U3682 (N_3682,N_1390,N_834);
nor U3683 (N_3683,N_1549,N_1189);
xnor U3684 (N_3684,N_1103,N_495);
xor U3685 (N_3685,N_96,N_1934);
nor U3686 (N_3686,N_174,N_141);
and U3687 (N_3687,N_140,N_432);
and U3688 (N_3688,N_1163,N_180);
nand U3689 (N_3689,N_576,N_847);
and U3690 (N_3690,N_213,N_889);
or U3691 (N_3691,N_1134,N_1382);
nand U3692 (N_3692,N_1021,N_41);
and U3693 (N_3693,N_640,N_491);
nor U3694 (N_3694,N_143,N_1973);
nand U3695 (N_3695,N_913,N_1119);
nor U3696 (N_3696,N_570,N_1000);
nand U3697 (N_3697,N_1099,N_1609);
nand U3698 (N_3698,N_871,N_741);
nand U3699 (N_3699,N_1718,N_1081);
xor U3700 (N_3700,N_568,N_4);
nor U3701 (N_3701,N_1689,N_1626);
or U3702 (N_3702,N_1135,N_611);
nor U3703 (N_3703,N_418,N_710);
or U3704 (N_3704,N_1169,N_859);
and U3705 (N_3705,N_1579,N_882);
or U3706 (N_3706,N_1814,N_1076);
xnor U3707 (N_3707,N_1002,N_589);
and U3708 (N_3708,N_1483,N_1505);
nor U3709 (N_3709,N_578,N_289);
and U3710 (N_3710,N_1060,N_1480);
or U3711 (N_3711,N_388,N_169);
and U3712 (N_3712,N_286,N_334);
nand U3713 (N_3713,N_1066,N_1254);
xor U3714 (N_3714,N_182,N_902);
nand U3715 (N_3715,N_929,N_987);
and U3716 (N_3716,N_1122,N_1773);
nand U3717 (N_3717,N_834,N_1026);
and U3718 (N_3718,N_647,N_629);
xor U3719 (N_3719,N_1839,N_1499);
xor U3720 (N_3720,N_1292,N_640);
xor U3721 (N_3721,N_755,N_1058);
and U3722 (N_3722,N_351,N_977);
or U3723 (N_3723,N_8,N_86);
and U3724 (N_3724,N_1410,N_15);
nor U3725 (N_3725,N_1355,N_317);
nor U3726 (N_3726,N_1466,N_698);
nand U3727 (N_3727,N_569,N_450);
and U3728 (N_3728,N_1437,N_1048);
xor U3729 (N_3729,N_1752,N_1508);
nand U3730 (N_3730,N_248,N_1600);
or U3731 (N_3731,N_74,N_479);
xnor U3732 (N_3732,N_324,N_1441);
and U3733 (N_3733,N_704,N_471);
nand U3734 (N_3734,N_760,N_1457);
nor U3735 (N_3735,N_1673,N_131);
nor U3736 (N_3736,N_1384,N_1682);
or U3737 (N_3737,N_1058,N_453);
xor U3738 (N_3738,N_1149,N_66);
nand U3739 (N_3739,N_477,N_187);
and U3740 (N_3740,N_1854,N_241);
nand U3741 (N_3741,N_612,N_1761);
or U3742 (N_3742,N_1477,N_1007);
xnor U3743 (N_3743,N_1599,N_1961);
or U3744 (N_3744,N_8,N_897);
and U3745 (N_3745,N_1237,N_25);
and U3746 (N_3746,N_1076,N_1831);
and U3747 (N_3747,N_1248,N_1507);
nand U3748 (N_3748,N_999,N_47);
nand U3749 (N_3749,N_949,N_393);
nor U3750 (N_3750,N_871,N_23);
or U3751 (N_3751,N_63,N_462);
xor U3752 (N_3752,N_77,N_969);
or U3753 (N_3753,N_706,N_190);
and U3754 (N_3754,N_1288,N_1672);
xor U3755 (N_3755,N_1598,N_315);
and U3756 (N_3756,N_505,N_7);
nor U3757 (N_3757,N_466,N_1023);
nor U3758 (N_3758,N_177,N_68);
or U3759 (N_3759,N_728,N_334);
or U3760 (N_3760,N_550,N_1286);
or U3761 (N_3761,N_1530,N_268);
or U3762 (N_3762,N_1595,N_1945);
and U3763 (N_3763,N_640,N_1348);
and U3764 (N_3764,N_592,N_1310);
or U3765 (N_3765,N_269,N_1443);
xor U3766 (N_3766,N_643,N_970);
and U3767 (N_3767,N_1723,N_126);
nor U3768 (N_3768,N_3,N_195);
and U3769 (N_3769,N_1684,N_719);
nand U3770 (N_3770,N_1185,N_1549);
nor U3771 (N_3771,N_1371,N_334);
xor U3772 (N_3772,N_1208,N_547);
or U3773 (N_3773,N_1452,N_473);
xnor U3774 (N_3774,N_103,N_251);
xor U3775 (N_3775,N_1508,N_1336);
nand U3776 (N_3776,N_454,N_1656);
xnor U3777 (N_3777,N_1379,N_389);
and U3778 (N_3778,N_1843,N_1796);
or U3779 (N_3779,N_719,N_613);
or U3780 (N_3780,N_994,N_705);
and U3781 (N_3781,N_1636,N_738);
nor U3782 (N_3782,N_1550,N_628);
or U3783 (N_3783,N_470,N_1197);
nor U3784 (N_3784,N_1708,N_1965);
and U3785 (N_3785,N_1609,N_31);
or U3786 (N_3786,N_849,N_650);
xor U3787 (N_3787,N_197,N_1668);
xor U3788 (N_3788,N_779,N_1659);
xor U3789 (N_3789,N_76,N_1420);
and U3790 (N_3790,N_1756,N_1924);
or U3791 (N_3791,N_307,N_863);
or U3792 (N_3792,N_618,N_1478);
or U3793 (N_3793,N_1165,N_404);
and U3794 (N_3794,N_262,N_1385);
nand U3795 (N_3795,N_1080,N_1386);
and U3796 (N_3796,N_1239,N_581);
or U3797 (N_3797,N_198,N_213);
or U3798 (N_3798,N_611,N_703);
or U3799 (N_3799,N_807,N_287);
xnor U3800 (N_3800,N_451,N_217);
nor U3801 (N_3801,N_800,N_416);
nand U3802 (N_3802,N_1289,N_34);
nor U3803 (N_3803,N_1926,N_1248);
or U3804 (N_3804,N_884,N_1734);
nor U3805 (N_3805,N_1593,N_1499);
xor U3806 (N_3806,N_1041,N_772);
xor U3807 (N_3807,N_27,N_457);
xnor U3808 (N_3808,N_712,N_875);
nor U3809 (N_3809,N_210,N_1772);
and U3810 (N_3810,N_206,N_1984);
and U3811 (N_3811,N_1858,N_60);
nor U3812 (N_3812,N_501,N_750);
nor U3813 (N_3813,N_60,N_406);
nand U3814 (N_3814,N_385,N_484);
and U3815 (N_3815,N_1121,N_1161);
nor U3816 (N_3816,N_592,N_1088);
nor U3817 (N_3817,N_57,N_1475);
xor U3818 (N_3818,N_424,N_1263);
nor U3819 (N_3819,N_298,N_1848);
or U3820 (N_3820,N_1870,N_108);
nor U3821 (N_3821,N_1542,N_724);
or U3822 (N_3822,N_106,N_1479);
nand U3823 (N_3823,N_234,N_1521);
and U3824 (N_3824,N_867,N_1712);
and U3825 (N_3825,N_1184,N_1553);
xor U3826 (N_3826,N_1765,N_786);
and U3827 (N_3827,N_1508,N_198);
or U3828 (N_3828,N_1653,N_227);
or U3829 (N_3829,N_1726,N_568);
xor U3830 (N_3830,N_1244,N_0);
and U3831 (N_3831,N_1148,N_1246);
xor U3832 (N_3832,N_387,N_1440);
xor U3833 (N_3833,N_1757,N_156);
or U3834 (N_3834,N_1871,N_1158);
nor U3835 (N_3835,N_917,N_3);
nand U3836 (N_3836,N_731,N_1780);
and U3837 (N_3837,N_1040,N_138);
nand U3838 (N_3838,N_1565,N_1536);
and U3839 (N_3839,N_1118,N_542);
xnor U3840 (N_3840,N_944,N_153);
xor U3841 (N_3841,N_1813,N_536);
nand U3842 (N_3842,N_1916,N_1045);
xnor U3843 (N_3843,N_913,N_2);
xnor U3844 (N_3844,N_599,N_252);
nor U3845 (N_3845,N_1334,N_116);
and U3846 (N_3846,N_844,N_386);
nor U3847 (N_3847,N_237,N_1576);
and U3848 (N_3848,N_308,N_884);
nand U3849 (N_3849,N_1898,N_907);
nand U3850 (N_3850,N_1819,N_301);
nor U3851 (N_3851,N_72,N_163);
and U3852 (N_3852,N_1436,N_1514);
and U3853 (N_3853,N_1949,N_1195);
nand U3854 (N_3854,N_522,N_56);
nor U3855 (N_3855,N_86,N_1746);
xnor U3856 (N_3856,N_1752,N_1799);
or U3857 (N_3857,N_404,N_1107);
nand U3858 (N_3858,N_1011,N_536);
nor U3859 (N_3859,N_614,N_1453);
or U3860 (N_3860,N_1721,N_1793);
xnor U3861 (N_3861,N_377,N_1642);
nor U3862 (N_3862,N_1880,N_1575);
nor U3863 (N_3863,N_1887,N_900);
and U3864 (N_3864,N_408,N_1184);
or U3865 (N_3865,N_1570,N_1191);
and U3866 (N_3866,N_1502,N_568);
or U3867 (N_3867,N_400,N_818);
or U3868 (N_3868,N_1651,N_591);
nand U3869 (N_3869,N_817,N_649);
xnor U3870 (N_3870,N_1120,N_765);
xor U3871 (N_3871,N_265,N_1645);
nor U3872 (N_3872,N_646,N_632);
nand U3873 (N_3873,N_662,N_531);
nor U3874 (N_3874,N_38,N_1066);
nor U3875 (N_3875,N_268,N_1268);
or U3876 (N_3876,N_718,N_1884);
xnor U3877 (N_3877,N_203,N_828);
or U3878 (N_3878,N_354,N_1238);
and U3879 (N_3879,N_1615,N_1106);
nand U3880 (N_3880,N_1214,N_995);
nor U3881 (N_3881,N_1133,N_300);
or U3882 (N_3882,N_1018,N_1330);
nor U3883 (N_3883,N_1532,N_1954);
and U3884 (N_3884,N_562,N_868);
and U3885 (N_3885,N_1181,N_713);
or U3886 (N_3886,N_507,N_634);
nor U3887 (N_3887,N_502,N_1924);
nor U3888 (N_3888,N_1049,N_1406);
xnor U3889 (N_3889,N_304,N_844);
and U3890 (N_3890,N_1183,N_149);
or U3891 (N_3891,N_1915,N_1651);
or U3892 (N_3892,N_346,N_1022);
nor U3893 (N_3893,N_1074,N_150);
and U3894 (N_3894,N_446,N_804);
and U3895 (N_3895,N_561,N_1513);
xor U3896 (N_3896,N_1512,N_1603);
and U3897 (N_3897,N_1619,N_534);
nor U3898 (N_3898,N_510,N_1513);
nor U3899 (N_3899,N_272,N_170);
nor U3900 (N_3900,N_1242,N_833);
or U3901 (N_3901,N_1914,N_1585);
and U3902 (N_3902,N_1061,N_1209);
xnor U3903 (N_3903,N_960,N_1377);
nor U3904 (N_3904,N_180,N_1840);
or U3905 (N_3905,N_1315,N_1574);
nor U3906 (N_3906,N_953,N_725);
xor U3907 (N_3907,N_901,N_876);
nand U3908 (N_3908,N_1960,N_906);
or U3909 (N_3909,N_238,N_1178);
nor U3910 (N_3910,N_3,N_1930);
xor U3911 (N_3911,N_1028,N_1703);
xor U3912 (N_3912,N_832,N_1263);
and U3913 (N_3913,N_1903,N_1682);
nor U3914 (N_3914,N_109,N_279);
nand U3915 (N_3915,N_478,N_1566);
nor U3916 (N_3916,N_310,N_1382);
nor U3917 (N_3917,N_24,N_423);
nor U3918 (N_3918,N_561,N_1766);
and U3919 (N_3919,N_1165,N_1027);
nor U3920 (N_3920,N_598,N_159);
nand U3921 (N_3921,N_1774,N_1249);
nor U3922 (N_3922,N_670,N_1209);
or U3923 (N_3923,N_517,N_85);
nor U3924 (N_3924,N_1794,N_867);
xnor U3925 (N_3925,N_424,N_306);
and U3926 (N_3926,N_1902,N_904);
xor U3927 (N_3927,N_470,N_1721);
nor U3928 (N_3928,N_1360,N_295);
or U3929 (N_3929,N_1398,N_316);
or U3930 (N_3930,N_1221,N_806);
nand U3931 (N_3931,N_1419,N_1667);
nor U3932 (N_3932,N_1086,N_324);
nor U3933 (N_3933,N_398,N_1153);
nor U3934 (N_3934,N_426,N_1022);
and U3935 (N_3935,N_1672,N_1884);
xor U3936 (N_3936,N_1618,N_1584);
nor U3937 (N_3937,N_1836,N_1086);
and U3938 (N_3938,N_425,N_40);
xor U3939 (N_3939,N_1827,N_1798);
nand U3940 (N_3940,N_18,N_1921);
xor U3941 (N_3941,N_190,N_1325);
nor U3942 (N_3942,N_428,N_83);
xor U3943 (N_3943,N_1190,N_1800);
nor U3944 (N_3944,N_868,N_122);
xor U3945 (N_3945,N_1511,N_1714);
nand U3946 (N_3946,N_1290,N_58);
nor U3947 (N_3947,N_873,N_846);
nor U3948 (N_3948,N_561,N_1732);
and U3949 (N_3949,N_1020,N_199);
xor U3950 (N_3950,N_1471,N_539);
nor U3951 (N_3951,N_1898,N_1420);
nor U3952 (N_3952,N_698,N_1444);
or U3953 (N_3953,N_1885,N_247);
xnor U3954 (N_3954,N_1505,N_1798);
and U3955 (N_3955,N_1176,N_1332);
nor U3956 (N_3956,N_663,N_528);
nor U3957 (N_3957,N_704,N_1997);
and U3958 (N_3958,N_1080,N_329);
and U3959 (N_3959,N_269,N_544);
nand U3960 (N_3960,N_131,N_493);
nand U3961 (N_3961,N_1827,N_1325);
and U3962 (N_3962,N_1375,N_674);
nand U3963 (N_3963,N_818,N_836);
xor U3964 (N_3964,N_746,N_1021);
nor U3965 (N_3965,N_910,N_555);
and U3966 (N_3966,N_798,N_1358);
or U3967 (N_3967,N_971,N_666);
nor U3968 (N_3968,N_1653,N_174);
nand U3969 (N_3969,N_633,N_1432);
nand U3970 (N_3970,N_1769,N_889);
xor U3971 (N_3971,N_92,N_1385);
nor U3972 (N_3972,N_465,N_1849);
or U3973 (N_3973,N_1553,N_152);
or U3974 (N_3974,N_246,N_665);
or U3975 (N_3975,N_712,N_317);
nor U3976 (N_3976,N_629,N_440);
and U3977 (N_3977,N_1611,N_1163);
xnor U3978 (N_3978,N_364,N_426);
nor U3979 (N_3979,N_725,N_475);
xor U3980 (N_3980,N_1631,N_461);
nand U3981 (N_3981,N_1820,N_552);
nor U3982 (N_3982,N_1842,N_1304);
or U3983 (N_3983,N_1765,N_236);
and U3984 (N_3984,N_930,N_1414);
nor U3985 (N_3985,N_1072,N_1789);
nor U3986 (N_3986,N_747,N_1121);
xor U3987 (N_3987,N_1717,N_55);
xnor U3988 (N_3988,N_1548,N_581);
xnor U3989 (N_3989,N_302,N_1623);
nand U3990 (N_3990,N_556,N_569);
nand U3991 (N_3991,N_632,N_1875);
xnor U3992 (N_3992,N_1337,N_1955);
nand U3993 (N_3993,N_1218,N_754);
nor U3994 (N_3994,N_1209,N_1367);
xnor U3995 (N_3995,N_1593,N_1097);
or U3996 (N_3996,N_1981,N_1491);
and U3997 (N_3997,N_224,N_300);
nor U3998 (N_3998,N_918,N_1154);
xnor U3999 (N_3999,N_1852,N_1060);
and U4000 (N_4000,N_2323,N_2251);
nor U4001 (N_4001,N_3209,N_2065);
xor U4002 (N_4002,N_2311,N_3767);
nand U4003 (N_4003,N_2166,N_3769);
nand U4004 (N_4004,N_3691,N_3310);
and U4005 (N_4005,N_3839,N_3731);
and U4006 (N_4006,N_2681,N_3408);
and U4007 (N_4007,N_2985,N_2649);
nor U4008 (N_4008,N_2400,N_3817);
or U4009 (N_4009,N_2536,N_3473);
and U4010 (N_4010,N_3646,N_2244);
nand U4011 (N_4011,N_3539,N_3964);
xor U4012 (N_4012,N_2146,N_2566);
and U4013 (N_4013,N_2697,N_2226);
and U4014 (N_4014,N_2891,N_3097);
and U4015 (N_4015,N_3466,N_3459);
nand U4016 (N_4016,N_3859,N_3126);
and U4017 (N_4017,N_2763,N_3193);
xnor U4018 (N_4018,N_3240,N_2627);
or U4019 (N_4019,N_2114,N_2658);
xnor U4020 (N_4020,N_3712,N_3447);
nor U4021 (N_4021,N_2471,N_3454);
nand U4022 (N_4022,N_2593,N_2623);
and U4023 (N_4023,N_3990,N_3878);
nand U4024 (N_4024,N_2437,N_3306);
xor U4025 (N_4025,N_3871,N_3138);
and U4026 (N_4026,N_2125,N_2701);
nand U4027 (N_4027,N_3376,N_3794);
xor U4028 (N_4028,N_2187,N_3321);
nor U4029 (N_4029,N_3457,N_3805);
or U4030 (N_4030,N_2721,N_2603);
xnor U4031 (N_4031,N_2759,N_3012);
xor U4032 (N_4032,N_3139,N_3026);
nand U4033 (N_4033,N_2950,N_3702);
nor U4034 (N_4034,N_2832,N_2825);
nor U4035 (N_4035,N_3673,N_3468);
nor U4036 (N_4036,N_2860,N_3086);
nand U4037 (N_4037,N_2385,N_3977);
xor U4038 (N_4038,N_2271,N_3687);
and U4039 (N_4039,N_2369,N_3505);
nand U4040 (N_4040,N_3207,N_3196);
nand U4041 (N_4041,N_2874,N_3530);
xor U4042 (N_4042,N_2038,N_2227);
nor U4043 (N_4043,N_3172,N_3893);
nor U4044 (N_4044,N_2497,N_3322);
nand U4045 (N_4045,N_2746,N_3287);
xnor U4046 (N_4046,N_2024,N_3594);
xnor U4047 (N_4047,N_3910,N_2961);
nor U4048 (N_4048,N_3617,N_2313);
nand U4049 (N_4049,N_2077,N_3043);
nand U4050 (N_4050,N_3875,N_3075);
and U4051 (N_4051,N_2944,N_3132);
xor U4052 (N_4052,N_3848,N_3865);
and U4053 (N_4053,N_2827,N_3599);
nor U4054 (N_4054,N_2104,N_3582);
xnor U4055 (N_4055,N_3986,N_3658);
nand U4056 (N_4056,N_2039,N_3180);
nor U4057 (N_4057,N_3860,N_2243);
xnor U4058 (N_4058,N_2738,N_2920);
and U4059 (N_4059,N_3532,N_3763);
nor U4060 (N_4060,N_2591,N_2850);
and U4061 (N_4061,N_3863,N_3598);
nor U4062 (N_4062,N_3269,N_2355);
and U4063 (N_4063,N_3359,N_3912);
nor U4064 (N_4064,N_3226,N_3386);
nand U4065 (N_4065,N_3958,N_2690);
or U4066 (N_4066,N_2736,N_2994);
xnor U4067 (N_4067,N_3719,N_2585);
xnor U4068 (N_4068,N_2584,N_2233);
and U4069 (N_4069,N_3162,N_2742);
or U4070 (N_4070,N_3645,N_3411);
and U4071 (N_4071,N_3881,N_3391);
nor U4072 (N_4072,N_2820,N_2667);
or U4073 (N_4073,N_2743,N_3201);
nor U4074 (N_4074,N_3874,N_3784);
or U4075 (N_4075,N_2100,N_3540);
xnor U4076 (N_4076,N_2792,N_3609);
and U4077 (N_4077,N_2021,N_3402);
nand U4078 (N_4078,N_3334,N_2777);
nor U4079 (N_4079,N_2859,N_3738);
xor U4080 (N_4080,N_3786,N_3689);
and U4081 (N_4081,N_3758,N_3536);
xnor U4082 (N_4082,N_2306,N_3818);
or U4083 (N_4083,N_2009,N_3041);
nor U4084 (N_4084,N_2678,N_3394);
xor U4085 (N_4085,N_3724,N_2664);
or U4086 (N_4086,N_2417,N_3980);
or U4087 (N_4087,N_2983,N_2491);
nand U4088 (N_4088,N_2554,N_2693);
xor U4089 (N_4089,N_2749,N_2153);
xor U4090 (N_4090,N_3785,N_3029);
xor U4091 (N_4091,N_2401,N_3605);
or U4092 (N_4092,N_3066,N_2943);
nand U4093 (N_4093,N_2391,N_3134);
nand U4094 (N_4094,N_2800,N_3621);
xnor U4095 (N_4095,N_3660,N_2479);
nor U4096 (N_4096,N_2216,N_3350);
nand U4097 (N_4097,N_3177,N_2117);
nand U4098 (N_4098,N_3975,N_2613);
nor U4099 (N_4099,N_2901,N_3713);
or U4100 (N_4100,N_2068,N_2632);
or U4101 (N_4101,N_2136,N_3850);
nor U4102 (N_4102,N_2949,N_2218);
and U4103 (N_4103,N_2428,N_3613);
xor U4104 (N_4104,N_2299,N_3588);
or U4105 (N_4105,N_3355,N_2045);
xnor U4106 (N_4106,N_2917,N_2288);
and U4107 (N_4107,N_3315,N_3557);
xor U4108 (N_4108,N_3418,N_2062);
nor U4109 (N_4109,N_2982,N_3781);
and U4110 (N_4110,N_3120,N_3119);
nor U4111 (N_4111,N_2550,N_3232);
nor U4112 (N_4112,N_3488,N_2202);
and U4113 (N_4113,N_3141,N_2217);
nand U4114 (N_4114,N_2439,N_3954);
and U4115 (N_4115,N_3427,N_3234);
and U4116 (N_4116,N_2722,N_3314);
or U4117 (N_4117,N_3375,N_2899);
or U4118 (N_4118,N_3511,N_2577);
and U4119 (N_4119,N_3371,N_3096);
nand U4120 (N_4120,N_2250,N_2198);
and U4121 (N_4121,N_3031,N_3789);
nand U4122 (N_4122,N_3705,N_3887);
or U4123 (N_4123,N_3053,N_2779);
xor U4124 (N_4124,N_2958,N_3560);
or U4125 (N_4125,N_2396,N_3534);
xor U4126 (N_4126,N_3111,N_2993);
and U4127 (N_4127,N_2212,N_2752);
and U4128 (N_4128,N_3927,N_2256);
and U4129 (N_4129,N_2641,N_3653);
or U4130 (N_4130,N_3970,N_2530);
nand U4131 (N_4131,N_2302,N_2647);
or U4132 (N_4132,N_3989,N_3243);
and U4133 (N_4133,N_3263,N_3469);
or U4134 (N_4134,N_2141,N_2631);
xor U4135 (N_4135,N_2078,N_3116);
nand U4136 (N_4136,N_2945,N_2972);
and U4137 (N_4137,N_2466,N_3723);
nor U4138 (N_4138,N_3498,N_3823);
or U4139 (N_4139,N_2162,N_3280);
nor U4140 (N_4140,N_2137,N_2711);
nand U4141 (N_4141,N_3065,N_2315);
nand U4142 (N_4142,N_3855,N_2607);
nor U4143 (N_4143,N_3393,N_2524);
nand U4144 (N_4144,N_3347,N_2283);
nor U4145 (N_4145,N_3815,N_3544);
and U4146 (N_4146,N_3746,N_3414);
or U4147 (N_4147,N_2959,N_2149);
xor U4148 (N_4148,N_3857,N_2456);
nor U4149 (N_4149,N_3034,N_2133);
and U4150 (N_4150,N_2535,N_3542);
and U4151 (N_4151,N_3017,N_3639);
or U4152 (N_4152,N_3308,N_2231);
xnor U4153 (N_4153,N_3305,N_3744);
nand U4154 (N_4154,N_3741,N_2526);
and U4155 (N_4155,N_2334,N_2872);
nor U4156 (N_4156,N_2578,N_2817);
or U4157 (N_4157,N_3324,N_2611);
nand U4158 (N_4158,N_2409,N_2942);
or U4159 (N_4159,N_2359,N_2617);
and U4160 (N_4160,N_3399,N_2729);
nand U4161 (N_4161,N_2203,N_3153);
nand U4162 (N_4162,N_2465,N_2925);
or U4163 (N_4163,N_2806,N_3307);
nand U4164 (N_4164,N_3509,N_3077);
or U4165 (N_4165,N_2432,N_2576);
nand U4166 (N_4166,N_2956,N_3128);
and U4167 (N_4167,N_3681,N_3795);
xnor U4168 (N_4168,N_2809,N_3888);
xor U4169 (N_4169,N_3842,N_2328);
xor U4170 (N_4170,N_3776,N_2616);
nor U4171 (N_4171,N_3803,N_2371);
and U4172 (N_4172,N_3819,N_2778);
or U4173 (N_4173,N_2853,N_2142);
nand U4174 (N_4174,N_2989,N_2073);
nand U4175 (N_4175,N_3661,N_2927);
xor U4176 (N_4176,N_3069,N_2067);
or U4177 (N_4177,N_2179,N_3407);
xor U4178 (N_4178,N_2508,N_3461);
nor U4179 (N_4179,N_3486,N_3400);
nor U4180 (N_4180,N_2708,N_3722);
nor U4181 (N_4181,N_2120,N_2544);
xor U4182 (N_4182,N_3650,N_3718);
xor U4183 (N_4183,N_2770,N_3877);
or U4184 (N_4184,N_2357,N_3625);
or U4185 (N_4185,N_2962,N_3677);
nor U4186 (N_4186,N_3514,N_2347);
or U4187 (N_4187,N_2317,N_3166);
and U4188 (N_4188,N_3891,N_3699);
nand U4189 (N_4189,N_3377,N_3965);
or U4190 (N_4190,N_2696,N_3657);
and U4191 (N_4191,N_3747,N_3754);
and U4192 (N_4192,N_2032,N_3853);
xnor U4193 (N_4193,N_3179,N_3429);
or U4194 (N_4194,N_3674,N_2205);
or U4195 (N_4195,N_3659,N_3242);
and U4196 (N_4196,N_3374,N_2050);
and U4197 (N_4197,N_2289,N_3846);
xor U4198 (N_4198,N_2384,N_2116);
or U4199 (N_4199,N_3778,N_2269);
nor U4200 (N_4200,N_2266,N_2420);
xor U4201 (N_4201,N_2837,N_3188);
nor U4202 (N_4202,N_2854,N_3892);
or U4203 (N_4203,N_3301,N_3337);
nand U4204 (N_4204,N_3155,N_3502);
nand U4205 (N_4205,N_2609,N_2265);
or U4206 (N_4206,N_3618,N_3472);
and U4207 (N_4207,N_2522,N_2574);
nand U4208 (N_4208,N_2772,N_2242);
xor U4209 (N_4209,N_2240,N_3279);
or U4210 (N_4210,N_2580,N_3309);
nor U4211 (N_4211,N_2731,N_2795);
and U4212 (N_4212,N_3283,N_2352);
and U4213 (N_4213,N_3707,N_3710);
nor U4214 (N_4214,N_2414,N_3147);
and U4215 (N_4215,N_2545,N_2312);
nor U4216 (N_4216,N_2886,N_2159);
nor U4217 (N_4217,N_2910,N_2127);
nor U4218 (N_4218,N_2913,N_2049);
nor U4219 (N_4219,N_2974,N_3316);
or U4220 (N_4220,N_3206,N_2634);
and U4221 (N_4221,N_2980,N_3071);
or U4222 (N_4222,N_2161,N_2534);
xnor U4223 (N_4223,N_2705,N_2625);
or U4224 (N_4224,N_2002,N_2807);
xnor U4225 (N_4225,N_3090,N_3050);
or U4226 (N_4226,N_2653,N_3431);
and U4227 (N_4227,N_2389,N_3870);
xor U4228 (N_4228,N_2458,N_2871);
nor U4229 (N_4229,N_3148,N_2119);
xnor U4230 (N_4230,N_3230,N_3124);
nand U4231 (N_4231,N_2904,N_2096);
or U4232 (N_4232,N_2619,N_2715);
xnor U4233 (N_4233,N_2200,N_3994);
or U4234 (N_4234,N_3146,N_3938);
and U4235 (N_4235,N_3112,N_3245);
nor U4236 (N_4236,N_2276,N_3336);
xor U4237 (N_4237,N_3083,N_3537);
nand U4238 (N_4238,N_3925,N_2622);
xor U4239 (N_4239,N_2150,N_2408);
and U4240 (N_4240,N_3918,N_2923);
or U4241 (N_4241,N_2745,N_2470);
or U4242 (N_4242,N_2686,N_3821);
and U4243 (N_4243,N_2248,N_3149);
xnor U4244 (N_4244,N_2713,N_3695);
and U4245 (N_4245,N_2586,N_3709);
or U4246 (N_4246,N_2430,N_2140);
nor U4247 (N_4247,N_2838,N_2842);
nor U4248 (N_4248,N_3951,N_2473);
xor U4249 (N_4249,N_2723,N_2571);
or U4250 (N_4250,N_3107,N_2134);
or U4251 (N_4251,N_2953,N_2789);
nor U4252 (N_4252,N_3942,N_3973);
nor U4253 (N_4253,N_2427,N_3231);
nor U4254 (N_4254,N_3142,N_2780);
or U4255 (N_4255,N_3296,N_2981);
or U4256 (N_4256,N_3780,N_2332);
or U4257 (N_4257,N_2630,N_3997);
nand U4258 (N_4258,N_2918,N_2884);
xor U4259 (N_4259,N_2080,N_2551);
xnor U4260 (N_4260,N_3450,N_3793);
and U4261 (N_4261,N_3067,N_2105);
and U4262 (N_4262,N_2033,N_2027);
and U4263 (N_4263,N_3908,N_3797);
or U4264 (N_4264,N_3289,N_2810);
and U4265 (N_4265,N_3042,N_3616);
or U4266 (N_4266,N_3843,N_3638);
or U4267 (N_4267,N_2402,N_3670);
and U4268 (N_4268,N_3932,N_3003);
nand U4269 (N_4269,N_3836,N_3903);
nor U4270 (N_4270,N_3030,N_3637);
and U4271 (N_4271,N_2001,N_3849);
or U4272 (N_4272,N_3759,N_3198);
nor U4273 (N_4273,N_2502,N_2646);
nand U4274 (N_4274,N_2714,N_3317);
nand U4275 (N_4275,N_3647,N_3277);
nor U4276 (N_4276,N_2973,N_3684);
nor U4277 (N_4277,N_2549,N_2675);
xnor U4278 (N_4278,N_2234,N_3612);
xnor U4279 (N_4279,N_2849,N_3313);
nand U4280 (N_4280,N_2000,N_3591);
nand U4281 (N_4281,N_2453,N_2539);
nor U4282 (N_4282,N_2346,N_2298);
nor U4283 (N_4283,N_2669,N_3143);
nand U4284 (N_4284,N_2181,N_2818);
and U4285 (N_4285,N_2195,N_2380);
nand U4286 (N_4286,N_2447,N_2254);
nor U4287 (N_4287,N_2022,N_3861);
xor U4288 (N_4288,N_2761,N_3465);
nand U4289 (N_4289,N_2558,N_3988);
nand U4290 (N_4290,N_3693,N_3607);
nor U4291 (N_4291,N_3113,N_3426);
and U4292 (N_4292,N_3448,N_2422);
xor U4293 (N_4293,N_2184,N_3928);
and U4294 (N_4294,N_2204,N_2025);
xnor U4295 (N_4295,N_2278,N_2037);
or U4296 (N_4296,N_2469,N_3424);
or U4297 (N_4297,N_2012,N_3569);
xnor U4298 (N_4298,N_3444,N_2513);
nor U4299 (N_4299,N_2360,N_3798);
xor U4300 (N_4300,N_2238,N_3257);
xnor U4301 (N_4301,N_2095,N_3222);
nand U4302 (N_4302,N_2434,N_2070);
or U4303 (N_4303,N_2748,N_2520);
or U4304 (N_4304,N_3696,N_2808);
or U4305 (N_4305,N_2433,N_3274);
nand U4306 (N_4306,N_2955,N_3165);
or U4307 (N_4307,N_2329,N_2528);
nor U4308 (N_4308,N_3950,N_3527);
or U4309 (N_4309,N_3868,N_2527);
nand U4310 (N_4310,N_3490,N_3156);
nor U4311 (N_4311,N_3549,N_2767);
nor U4312 (N_4312,N_3227,N_3300);
nand U4313 (N_4313,N_3915,N_3039);
and U4314 (N_4314,N_2351,N_3690);
nor U4315 (N_4315,N_3401,N_2691);
nand U4316 (N_4316,N_2628,N_3183);
and U4317 (N_4317,N_3035,N_3403);
xor U4318 (N_4318,N_3299,N_2031);
nand U4319 (N_4319,N_2660,N_3772);
and U4320 (N_4320,N_3574,N_2754);
and U4321 (N_4321,N_3682,N_2684);
or U4322 (N_4322,N_2887,N_2086);
xor U4323 (N_4323,N_2044,N_2376);
nor U4324 (N_4324,N_2597,N_2556);
nor U4325 (N_4325,N_3896,N_3356);
or U4326 (N_4326,N_2353,N_3409);
nand U4327 (N_4327,N_2518,N_3022);
xor U4328 (N_4328,N_2139,N_3464);
xnor U4329 (N_4329,N_2232,N_2112);
nand U4330 (N_4330,N_3174,N_2774);
xnor U4331 (N_4331,N_3512,N_3940);
nand U4332 (N_4332,N_2052,N_2848);
and U4333 (N_4333,N_2395,N_2998);
nor U4334 (N_4334,N_3028,N_2172);
nand U4335 (N_4335,N_2303,N_2103);
xnor U4336 (N_4336,N_2113,N_3711);
nand U4337 (N_4337,N_2438,N_3771);
nor U4338 (N_4338,N_2907,N_2403);
or U4339 (N_4339,N_2292,N_3291);
and U4340 (N_4340,N_3482,N_3969);
or U4341 (N_4341,N_3191,N_3880);
xor U4342 (N_4342,N_2131,N_3249);
nor U4343 (N_4343,N_3831,N_3665);
xor U4344 (N_4344,N_3905,N_2448);
and U4345 (N_4345,N_3985,N_3876);
or U4346 (N_4346,N_3115,N_2559);
xnor U4347 (N_4347,N_2946,N_3907);
or U4348 (N_4348,N_2514,N_2199);
nor U4349 (N_4349,N_2305,N_3364);
nand U4350 (N_4350,N_2883,N_2503);
nor U4351 (N_4351,N_3862,N_3211);
xor U4352 (N_4352,N_3254,N_2034);
or U4353 (N_4353,N_3742,N_3372);
xnor U4354 (N_4354,N_2567,N_2188);
nand U4355 (N_4355,N_2128,N_2970);
and U4356 (N_4356,N_3700,N_2270);
xnor U4357 (N_4357,N_3370,N_2718);
or U4358 (N_4358,N_2167,N_3501);
or U4359 (N_4359,N_3922,N_2564);
nand U4360 (N_4360,N_3378,N_3072);
or U4361 (N_4361,N_2169,N_3528);
or U4362 (N_4362,N_2379,N_3435);
and U4363 (N_4363,N_2364,N_3239);
and U4364 (N_4364,N_2900,N_2126);
nand U4365 (N_4365,N_2444,N_3290);
nand U4366 (N_4366,N_3353,N_2356);
nor U4367 (N_4367,N_2682,N_2732);
or U4368 (N_4368,N_3416,N_2542);
nor U4369 (N_4369,N_2707,N_2858);
nor U4370 (N_4370,N_3235,N_3396);
nand U4371 (N_4371,N_3456,N_2099);
or U4372 (N_4372,N_3100,N_3799);
or U4373 (N_4373,N_2300,N_3268);
xnor U4374 (N_4374,N_2785,N_3013);
xnor U4375 (N_4375,N_2197,N_2361);
or U4376 (N_4376,N_3643,N_2260);
nand U4377 (N_4377,N_3921,N_3001);
xnor U4378 (N_4378,N_3766,N_3945);
or U4379 (N_4379,N_2796,N_3966);
and U4380 (N_4380,N_2563,N_2835);
nor U4381 (N_4381,N_3672,N_3133);
nor U4382 (N_4382,N_3809,N_3432);
xor U4383 (N_4383,N_3389,N_2781);
or U4384 (N_4384,N_3341,N_3743);
nand U4385 (N_4385,N_2876,N_3587);
and U4386 (N_4386,N_3982,N_3601);
nand U4387 (N_4387,N_3953,N_3824);
or U4388 (N_4388,N_2392,N_2277);
xor U4389 (N_4389,N_3890,N_2857);
nor U4390 (N_4390,N_2787,N_2589);
and U4391 (N_4391,N_3015,N_3236);
or U4392 (N_4392,N_2821,N_2237);
xor U4393 (N_4393,N_3923,N_2336);
and U4394 (N_4394,N_2688,N_2110);
xnor U4395 (N_4395,N_2279,N_2786);
and U4396 (N_4396,N_3487,N_2388);
xor U4397 (N_4397,N_2043,N_2515);
and U4398 (N_4398,N_2063,N_2685);
nor U4399 (N_4399,N_2252,N_2436);
or U4400 (N_4400,N_3900,N_3791);
and U4401 (N_4401,N_3732,N_3760);
and U4402 (N_4402,N_3749,N_3960);
and U4403 (N_4403,N_2865,N_3556);
nand U4404 (N_4404,N_2147,N_3761);
xnor U4405 (N_4405,N_2964,N_2879);
xor U4406 (N_4406,N_3293,N_2957);
nand U4407 (N_4407,N_3292,N_2092);
and U4408 (N_4408,N_3538,N_2138);
xnor U4409 (N_4409,N_2030,N_2247);
nor U4410 (N_4410,N_2794,N_3380);
or U4411 (N_4411,N_2703,N_2291);
nand U4412 (N_4412,N_3641,N_3273);
nand U4413 (N_4413,N_3089,N_2111);
nor U4414 (N_4414,N_2893,N_3417);
and U4415 (N_4415,N_2282,N_3099);
and U4416 (N_4416,N_2737,N_3669);
xor U4417 (N_4417,N_3518,N_3590);
or U4418 (N_4418,N_3550,N_3081);
xnor U4419 (N_4419,N_3276,N_3999);
nand U4420 (N_4420,N_2938,N_2229);
nand U4421 (N_4421,N_3851,N_3131);
and U4422 (N_4422,N_2840,N_3004);
nor U4423 (N_4423,N_3886,N_3820);
xnor U4424 (N_4424,N_3589,N_3879);
or U4425 (N_4425,N_2459,N_2093);
and U4426 (N_4426,N_2969,N_2868);
nor U4427 (N_4427,N_2101,N_2405);
nand U4428 (N_4428,N_2977,N_2867);
xnor U4429 (N_4429,N_3184,N_2057);
or U4430 (N_4430,N_2725,N_2201);
nand U4431 (N_4431,N_2028,N_3398);
and U4432 (N_4432,N_2683,N_2168);
xor U4433 (N_4433,N_3271,N_3118);
xnor U4434 (N_4434,N_2386,N_2863);
nor U4435 (N_4435,N_3369,N_2839);
and U4436 (N_4436,N_2965,N_3439);
nand U4437 (N_4437,N_3847,N_3573);
nor U4438 (N_4438,N_3517,N_3845);
and U4439 (N_4439,N_3603,N_3579);
nor U4440 (N_4440,N_3127,N_3971);
or U4441 (N_4441,N_3552,N_2579);
and U4442 (N_4442,N_3554,N_3320);
or U4443 (N_4443,N_3108,N_3221);
and U4444 (N_4444,N_3093,N_2185);
nand U4445 (N_4445,N_3830,N_3570);
and U4446 (N_4446,N_3508,N_2295);
xnor U4447 (N_4447,N_2370,N_3460);
and U4448 (N_4448,N_2418,N_2933);
and U4449 (N_4449,N_2375,N_2107);
or U4450 (N_4450,N_2618,N_2803);
nor U4451 (N_4451,N_2733,N_2006);
nand U4452 (N_4452,N_3430,N_2449);
nor U4453 (N_4453,N_2213,N_2852);
nor U4454 (N_4454,N_3506,N_3024);
nand U4455 (N_4455,N_2275,N_2354);
or U4456 (N_4456,N_3051,N_2608);
or U4457 (N_4457,N_3628,N_3976);
nor U4458 (N_4458,N_2565,N_3318);
and U4459 (N_4459,N_3858,N_2979);
nand U4460 (N_4460,N_3462,N_2525);
or U4461 (N_4461,N_2489,N_3930);
nand U4462 (N_4462,N_2997,N_2988);
nor U4463 (N_4463,N_3410,N_2239);
nor U4464 (N_4464,N_3828,N_2054);
and U4465 (N_4465,N_3212,N_2454);
nand U4466 (N_4466,N_2679,N_2570);
nor U4467 (N_4467,N_3205,N_3151);
nor U4468 (N_4468,N_2814,N_2186);
xnor U4469 (N_4469,N_3882,N_2478);
and U4470 (N_4470,N_3568,N_2498);
or U4471 (N_4471,N_3802,N_3991);
xor U4472 (N_4472,N_2665,N_2855);
nand U4473 (N_4473,N_2426,N_2079);
nand U4474 (N_4474,N_3622,N_3624);
nand U4475 (N_4475,N_2366,N_3023);
nor U4476 (N_4476,N_3040,N_3841);
or U4477 (N_4477,N_3467,N_2488);
nor U4478 (N_4478,N_2612,N_3685);
nor U4479 (N_4479,N_2562,N_3010);
and U4480 (N_4480,N_3885,N_2460);
xor U4481 (N_4481,N_2557,N_3106);
xor U4482 (N_4482,N_2916,N_2877);
nand U4483 (N_4483,N_3018,N_2783);
or U4484 (N_4484,N_2692,N_2744);
or U4485 (N_4485,N_2183,N_2286);
nor U4486 (N_4486,N_2450,N_2178);
and U4487 (N_4487,N_2776,N_2790);
or U4488 (N_4488,N_2069,N_2727);
nand U4489 (N_4489,N_3957,N_2640);
nand U4490 (N_4490,N_2059,N_3365);
or U4491 (N_4491,N_2419,N_3440);
nand U4492 (N_4492,N_2823,N_2924);
and U4493 (N_4493,N_2098,N_3423);
or U4494 (N_4494,N_2581,N_2784);
nor U4495 (N_4495,N_3395,N_2058);
xnor U4496 (N_4496,N_2143,N_2174);
or U4497 (N_4497,N_2753,N_2151);
nand U4498 (N_4498,N_2245,N_2053);
xor U4499 (N_4499,N_3934,N_2413);
and U4500 (N_4500,N_3158,N_2671);
and U4501 (N_4501,N_3181,N_2163);
nor U4502 (N_4502,N_2674,N_3963);
and U4503 (N_4503,N_3704,N_3543);
xnor U4504 (N_4504,N_3102,N_2091);
nor U4505 (N_4505,N_2225,N_2755);
nor U4506 (N_4506,N_3161,N_2075);
xor U4507 (N_4507,N_2097,N_3475);
xor U4508 (N_4508,N_2728,N_2509);
nand U4509 (N_4509,N_2709,N_2689);
and U4510 (N_4510,N_3248,N_2331);
nor U4511 (N_4511,N_3671,N_3913);
nand U4512 (N_4512,N_3911,N_2843);
nor U4513 (N_4513,N_2533,N_2210);
or U4514 (N_4514,N_2132,N_3074);
nor U4515 (N_4515,N_2464,N_2494);
xnor U4516 (N_4516,N_3178,N_2967);
nor U4517 (N_4517,N_2788,N_3154);
nand U4518 (N_4518,N_2064,N_3379);
xor U4519 (N_4519,N_3854,N_3303);
and U4520 (N_4520,N_3256,N_2804);
nand U4521 (N_4521,N_3260,N_2540);
nand U4522 (N_4522,N_3553,N_3752);
and U4523 (N_4523,N_2510,N_3917);
nand U4524 (N_4524,N_2712,N_2005);
nand U4525 (N_4525,N_2694,N_2934);
nor U4526 (N_4526,N_2056,N_2659);
nand U4527 (N_4527,N_2990,N_3470);
nand U4528 (N_4528,N_2258,N_2164);
nand U4529 (N_4529,N_2764,N_2071);
or U4530 (N_4530,N_2841,N_2845);
and U4531 (N_4531,N_3524,N_2452);
nor U4532 (N_4532,N_3032,N_3826);
nand U4533 (N_4533,N_2768,N_2507);
nor U4534 (N_4534,N_3992,N_3972);
nand U4535 (N_4535,N_3076,N_3576);
nand U4536 (N_4536,N_3054,N_2157);
nor U4537 (N_4537,N_3648,N_3397);
nand U4538 (N_4538,N_3706,N_2398);
or U4539 (N_4539,N_3489,N_2606);
nand U4540 (N_4540,N_2381,N_3748);
nor U4541 (N_4541,N_2257,N_3644);
xor U4542 (N_4542,N_3006,N_2812);
or U4543 (N_4543,N_3002,N_2553);
nor U4544 (N_4544,N_3387,N_2895);
nor U4545 (N_4545,N_3164,N_2090);
nor U4546 (N_4546,N_3816,N_3063);
nor U4547 (N_4547,N_2273,N_3762);
and U4548 (N_4548,N_3463,N_2272);
xnor U4549 (N_4549,N_3103,N_2797);
nand U4550 (N_4550,N_3906,N_3493);
nor U4551 (N_4551,N_2984,N_3941);
and U4552 (N_4552,N_2040,N_3123);
and U4553 (N_4553,N_2477,N_3228);
or U4554 (N_4554,N_2321,N_3135);
xor U4555 (N_4555,N_2948,N_2824);
nor U4556 (N_4556,N_3419,N_2762);
nor U4557 (N_4557,N_2087,N_3325);
and U4558 (N_4558,N_3458,N_2246);
and U4559 (N_4559,N_3244,N_2897);
nor U4560 (N_4560,N_2154,N_3122);
nor U4561 (N_4561,N_2735,N_3340);
xnor U4562 (N_4562,N_2451,N_2831);
nand U4563 (N_4563,N_2223,N_2615);
or U4564 (N_4564,N_2373,N_3297);
or U4565 (N_4565,N_2221,N_2194);
nor U4566 (N_4566,N_2666,N_2122);
nand U4567 (N_4567,N_3087,N_3241);
and U4568 (N_4568,N_3631,N_2211);
or U4569 (N_4569,N_3577,N_2870);
nor U4570 (N_4570,N_2224,N_3642);
nand U4571 (N_4571,N_2176,N_2284);
nand U4572 (N_4572,N_2656,N_2512);
nor U4573 (N_4573,N_2481,N_3262);
xor U4574 (N_4574,N_2844,N_3796);
nor U4575 (N_4575,N_2532,N_3629);
nor U4576 (N_4576,N_3593,N_3105);
nor U4577 (N_4577,N_3171,N_3663);
or U4578 (N_4578,N_3788,N_2757);
and U4579 (N_4579,N_2324,N_2209);
xor U4580 (N_4580,N_3121,N_3753);
nand U4581 (N_4581,N_2911,N_3224);
xnor U4582 (N_4582,N_3392,N_2495);
nor U4583 (N_4583,N_2480,N_2267);
nor U4584 (N_4584,N_2011,N_3483);
nand U4585 (N_4585,N_2878,N_3060);
xor U4586 (N_4586,N_2724,N_3697);
xnor U4587 (N_4587,N_3484,N_2429);
xnor U4588 (N_4588,N_2516,N_3007);
and U4589 (N_4589,N_2548,N_3694);
xor U4590 (N_4590,N_3825,N_3765);
nor U4591 (N_4591,N_2261,N_2773);
nand U4592 (N_4592,N_2875,N_3728);
nand U4593 (N_4593,N_2108,N_2475);
xnor U4594 (N_4594,N_2546,N_2263);
or U4595 (N_4595,N_2416,N_2170);
nand U4596 (N_4596,N_3926,N_2130);
nor U4597 (N_4597,N_2294,N_3252);
and U4598 (N_4598,N_3654,N_2960);
nor U4599 (N_4599,N_3703,N_2274);
and U4600 (N_4600,N_3421,N_3919);
and U4601 (N_4601,N_2932,N_2811);
nor U4602 (N_4602,N_3175,N_2856);
nand U4603 (N_4603,N_3827,N_2072);
or U4604 (N_4604,N_2412,N_2873);
nand U4605 (N_4605,N_2582,N_3323);
or U4606 (N_4606,N_3608,N_3924);
and U4607 (N_4607,N_3838,N_3548);
nand U4608 (N_4608,N_3688,N_2862);
and U4609 (N_4609,N_2782,N_2866);
or U4610 (N_4610,N_3844,N_3288);
or U4611 (N_4611,N_2083,N_2484);
xor U4612 (N_4612,N_3783,N_3413);
or U4613 (N_4613,N_2036,N_3480);
or U4614 (N_4614,N_2106,N_2322);
xnor U4615 (N_4615,N_3445,N_3496);
xnor U4616 (N_4616,N_2493,N_2010);
nand U4617 (N_4617,N_3266,N_2173);
nor U4618 (N_4618,N_2165,N_2588);
or U4619 (N_4619,N_3962,N_3751);
xnor U4620 (N_4620,N_3437,N_3675);
xnor U4621 (N_4621,N_3443,N_2102);
nand U4622 (N_4622,N_2880,N_2791);
xor U4623 (N_4623,N_3987,N_2307);
nor U4624 (N_4624,N_3895,N_3564);
and U4625 (N_4625,N_3500,N_2327);
xnor U4626 (N_4626,N_2644,N_3384);
xnor U4627 (N_4627,N_2023,N_3937);
or U4628 (N_4628,N_3479,N_3258);
xnor U4629 (N_4629,N_3720,N_3555);
nor U4630 (N_4630,N_2082,N_3190);
nor U4631 (N_4631,N_3680,N_2363);
and U4632 (N_4632,N_3967,N_2255);
or U4633 (N_4633,N_2383,N_2042);
xor U4634 (N_4634,N_3770,N_2341);
xor U4635 (N_4635,N_2325,N_3110);
or U4636 (N_4636,N_3412,N_2511);
xnor U4637 (N_4637,N_3202,N_3575);
nor U4638 (N_4638,N_2220,N_3052);
xor U4639 (N_4639,N_3884,N_3664);
nand U4640 (N_4640,N_3057,N_3070);
or U4641 (N_4641,N_2214,N_3078);
nor U4642 (N_4642,N_2730,N_3058);
nor U4643 (N_4643,N_3600,N_2799);
nand U4644 (N_4644,N_3852,N_3894);
nand U4645 (N_4645,N_2485,N_2118);
or U4646 (N_4646,N_2316,N_3551);
nand U4647 (N_4647,N_2645,N_3187);
nand U4648 (N_4648,N_3814,N_2015);
or U4649 (N_4649,N_2968,N_2765);
and U4650 (N_4650,N_2061,N_2741);
and U4651 (N_4651,N_2861,N_3726);
nand U4652 (N_4652,N_3062,N_2995);
or U4653 (N_4653,N_3944,N_2604);
xnor U4654 (N_4654,N_3114,N_3092);
nand U4655 (N_4655,N_2561,N_3633);
xnor U4656 (N_4656,N_2538,N_2521);
nor U4657 (N_4657,N_3329,N_3602);
or U4658 (N_4658,N_3562,N_3091);
nand U4659 (N_4659,N_2483,N_2517);
and U4660 (N_4660,N_3567,N_2293);
nand U4661 (N_4661,N_2643,N_3436);
nand U4662 (N_4662,N_3721,N_2555);
nor U4663 (N_4663,N_3883,N_2020);
and U4664 (N_4664,N_2486,N_3189);
and U4665 (N_4665,N_2706,N_2704);
nor U4666 (N_4666,N_2621,N_2410);
or U4667 (N_4667,N_3104,N_2902);
or U4668 (N_4668,N_3129,N_2287);
or U4669 (N_4669,N_2937,N_2115);
nand U4670 (N_4670,N_2655,N_3130);
xnor U4671 (N_4671,N_2301,N_3757);
and U4672 (N_4672,N_3995,N_3192);
and U4673 (N_4673,N_2672,N_2999);
xor U4674 (N_4674,N_3197,N_3251);
xnor U4675 (N_4675,N_3730,N_2602);
or U4676 (N_4676,N_2531,N_2441);
nand U4677 (N_4677,N_2190,N_3020);
or U4678 (N_4678,N_3352,N_2348);
and U4679 (N_4679,N_3253,N_3952);
nor U4680 (N_4680,N_3729,N_2710);
and U4681 (N_4681,N_2822,N_3813);
xor U4682 (N_4682,N_2805,N_2629);
and U4683 (N_4683,N_3745,N_2716);
xnor U4684 (N_4684,N_3782,N_3056);
and U4685 (N_4685,N_3319,N_3832);
nor U4686 (N_4686,N_3194,N_2626);
and U4687 (N_4687,N_3656,N_3358);
nand U4688 (N_4688,N_2519,N_3904);
or U4689 (N_4689,N_3302,N_2066);
nand U4690 (N_4690,N_3168,N_3088);
nand U4691 (N_4691,N_3929,N_2084);
nand U4692 (N_4692,N_3216,N_2048);
nor U4693 (N_4693,N_3773,N_3453);
nand U4694 (N_4694,N_3014,N_3755);
and U4695 (N_4695,N_3167,N_3596);
and U4696 (N_4696,N_2652,N_3727);
or U4697 (N_4697,N_3219,N_3478);
xor U4698 (N_4698,N_3420,N_2543);
nand U4699 (N_4699,N_2864,N_3516);
nand U4700 (N_4700,N_2560,N_3225);
nand U4701 (N_4701,N_2008,N_3298);
xor U4702 (N_4702,N_3363,N_3565);
xnor U4703 (N_4703,N_3583,N_3085);
nand U4704 (N_4704,N_2129,N_3422);
and U4705 (N_4705,N_3936,N_3047);
and U4706 (N_4706,N_3666,N_2747);
nor U4707 (N_4707,N_3733,N_2007);
nor U4708 (N_4708,N_2881,N_2815);
xor U4709 (N_4709,N_3902,N_3270);
and U4710 (N_4710,N_3474,N_2657);
xor U4711 (N_4711,N_3634,N_2177);
nor U4712 (N_4712,N_2894,N_3275);
nand U4713 (N_4713,N_3630,N_3507);
and U4714 (N_4714,N_2687,N_3611);
nand U4715 (N_4715,N_2775,N_2374);
nor U4716 (N_4716,N_3278,N_2041);
or U4717 (N_4717,N_3351,N_3580);
xor U4718 (N_4718,N_3649,N_2830);
and U4719 (N_4719,N_3898,N_2310);
nand U4720 (N_4720,N_3485,N_2869);
and U4721 (N_4721,N_2156,N_3521);
or U4722 (N_4722,N_2939,N_2547);
xor U4723 (N_4723,N_3790,N_2411);
and U4724 (N_4724,N_3223,N_3717);
nand U4725 (N_4725,N_2222,N_2594);
nor U4726 (N_4726,N_3668,N_2636);
xnor U4727 (N_4727,N_3522,N_3974);
nor U4728 (N_4728,N_2431,N_3592);
nand U4729 (N_4729,N_2651,N_2445);
nand U4730 (N_4730,N_3199,N_3943);
and U4731 (N_4731,N_2846,N_3021);
xnor U4732 (N_4732,N_3504,N_3571);
and U4733 (N_4733,N_3247,N_2991);
xor U4734 (N_4734,N_2462,N_2055);
nand U4735 (N_4735,N_3455,N_2750);
nand U4736 (N_4736,N_3327,N_2638);
nor U4737 (N_4737,N_3652,N_3840);
and U4738 (N_4738,N_2523,N_2793);
xor U4739 (N_4739,N_3833,N_3169);
nand U4740 (N_4740,N_2319,N_2047);
xnor U4741 (N_4741,N_2333,N_2892);
nor U4742 (N_4742,N_3939,N_2828);
xnor U4743 (N_4743,N_3585,N_2717);
or U4744 (N_4744,N_3441,N_3856);
nor U4745 (N_4745,N_3203,N_3737);
xnor U4746 (N_4746,N_3025,N_3740);
and U4747 (N_4747,N_3217,N_2425);
nor U4748 (N_4748,N_2349,N_3332);
nor U4749 (N_4749,N_2587,N_3495);
nor U4750 (N_4750,N_2680,N_2350);
and U4751 (N_4751,N_2144,N_3775);
or U4752 (N_4752,N_2148,N_2378);
xor U4753 (N_4753,N_2152,N_2074);
nor U4754 (N_4754,N_3382,N_2035);
nor U4755 (N_4755,N_3619,N_3811);
xor U4756 (N_4756,N_3812,N_2668);
and U4757 (N_4757,N_2026,N_2898);
and U4758 (N_4758,N_3033,N_3218);
nor U4759 (N_4759,N_2280,N_3446);
nor U4760 (N_4760,N_3210,N_3173);
and U4761 (N_4761,N_3572,N_2909);
or U4762 (N_4762,N_2505,N_3584);
and U4763 (N_4763,N_3993,N_3736);
xnor U4764 (N_4764,N_3438,N_2192);
and U4765 (N_4765,N_2155,N_2387);
nor U4766 (N_4766,N_3405,N_2700);
nand U4767 (N_4767,N_3901,N_2193);
nand U4768 (N_4768,N_3094,N_3547);
xnor U4769 (N_4769,N_3604,N_2281);
nand U4770 (N_4770,N_3343,N_3038);
and U4771 (N_4771,N_3768,N_3360);
nor U4772 (N_4772,N_2051,N_3185);
xor U4773 (N_4773,N_3983,N_2912);
and U4774 (N_4774,N_3933,N_3497);
and U4775 (N_4775,N_3679,N_2829);
and U4776 (N_4776,N_3019,N_3515);
nand U4777 (N_4777,N_2342,N_3061);
and U4778 (N_4778,N_3255,N_3434);
xor U4779 (N_4779,N_2896,N_2605);
nand U4780 (N_4780,N_3238,N_2926);
and U4781 (N_4781,N_3049,N_3715);
nor U4782 (N_4782,N_2230,N_3714);
or U4783 (N_4783,N_3931,N_3792);
xor U4784 (N_4784,N_2596,N_2377);
or U4785 (N_4785,N_2338,N_2541);
xnor U4786 (N_4786,N_2492,N_2259);
nand U4787 (N_4787,N_2882,N_3519);
nor U4788 (N_4788,N_3626,N_2344);
xor U4789 (N_4789,N_3481,N_2235);
or U4790 (N_4790,N_2382,N_3581);
or U4791 (N_4791,N_2739,N_3361);
and U4792 (N_4792,N_2661,N_3079);
xor U4793 (N_4793,N_2847,N_3449);
xor U4794 (N_4794,N_2620,N_2905);
nand U4795 (N_4795,N_2215,N_3959);
nor U4796 (N_4796,N_3304,N_2599);
and U4797 (N_4797,N_2930,N_2330);
nor U4798 (N_4798,N_2552,N_2935);
nor U4799 (N_4799,N_3914,N_3182);
and U4800 (N_4800,N_2941,N_3476);
xor U4801 (N_4801,N_2952,N_3806);
or U4802 (N_4802,N_3281,N_2996);
and U4803 (N_4803,N_2397,N_3916);
nand U4804 (N_4804,N_3683,N_3285);
nor U4805 (N_4805,N_2109,N_3701);
and U4806 (N_4806,N_2992,N_2335);
or U4807 (N_4807,N_2833,N_2583);
nand U4808 (N_4808,N_2504,N_3935);
xor U4809 (N_4809,N_2457,N_3667);
or U4810 (N_4810,N_2637,N_2228);
nand U4811 (N_4811,N_3810,N_3272);
and U4812 (N_4812,N_2455,N_3491);
and U4813 (N_4813,N_2019,N_3494);
or U4814 (N_4814,N_2145,N_3433);
nand U4815 (N_4815,N_2986,N_3899);
nor U4816 (N_4816,N_3259,N_3286);
and U4817 (N_4817,N_2390,N_3345);
or U4818 (N_4818,N_3328,N_2207);
nor U4819 (N_4819,N_2423,N_3578);
nand U4820 (N_4820,N_3009,N_3098);
or U4821 (N_4821,N_3140,N_3708);
xnor U4822 (N_4822,N_3610,N_2487);
and U4823 (N_4823,N_2568,N_2914);
nand U4824 (N_4824,N_3150,N_3981);
nor U4825 (N_4825,N_2971,N_3442);
nand U4826 (N_4826,N_3606,N_3368);
or U4827 (N_4827,N_2472,N_3295);
nor U4828 (N_4828,N_3837,N_2816);
nand U4829 (N_4829,N_3872,N_3330);
and U4830 (N_4830,N_3620,N_2249);
or U4831 (N_4831,N_2798,N_2826);
nand U4832 (N_4832,N_3545,N_2158);
and U4833 (N_4833,N_2695,N_2889);
xnor U4834 (N_4834,N_2766,N_2676);
nor U4835 (N_4835,N_2801,N_2851);
and U4836 (N_4836,N_3208,N_2635);
or U4837 (N_4837,N_2308,N_2819);
and U4838 (N_4838,N_2756,N_3346);
xnor U4839 (N_4839,N_3348,N_3739);
nand U4840 (N_4840,N_2367,N_3632);
xnor U4841 (N_4841,N_3627,N_3160);
xnor U4842 (N_4842,N_2573,N_3068);
xor U4843 (N_4843,N_2677,N_2813);
nor U4844 (N_4844,N_2575,N_3250);
and U4845 (N_4845,N_3586,N_2421);
nor U4846 (N_4846,N_3615,N_3949);
and U4847 (N_4847,N_2662,N_2702);
xor U4848 (N_4848,N_2903,N_3000);
xor U4849 (N_4849,N_2719,N_2253);
nor U4850 (N_4850,N_2337,N_2673);
nand U4851 (N_4851,N_3533,N_3525);
and U4852 (N_4852,N_3008,N_3366);
xor U4853 (N_4853,N_2060,N_3563);
nor U4854 (N_4854,N_3046,N_3559);
xor U4855 (N_4855,N_2309,N_3635);
nor U4856 (N_4856,N_3152,N_3220);
or U4857 (N_4857,N_2393,N_2474);
and U4858 (N_4858,N_3655,N_3835);
and U4859 (N_4859,N_2123,N_3357);
or U4860 (N_4860,N_3233,N_2598);
xor U4861 (N_4861,N_2929,N_3734);
xor U4862 (N_4862,N_3157,N_2440);
nor U4863 (N_4863,N_2171,N_2435);
xnor U4864 (N_4864,N_2921,N_3869);
nor U4865 (N_4865,N_3073,N_3342);
or U4866 (N_4866,N_2501,N_2506);
and U4867 (N_4867,N_3822,N_2182);
nand U4868 (N_4868,N_2769,N_2482);
or U4869 (N_4869,N_3523,N_3640);
or U4870 (N_4870,N_3101,N_2963);
xor U4871 (N_4871,N_3801,N_3037);
or U4872 (N_4872,N_3333,N_2468);
xnor U4873 (N_4873,N_2936,N_3200);
or U4874 (N_4874,N_2415,N_3176);
nand U4875 (N_4875,N_3381,N_2834);
or U4876 (N_4876,N_3349,N_2740);
and U4877 (N_4877,N_3948,N_3452);
or U4878 (N_4878,N_3016,N_2648);
xor U4879 (N_4879,N_2362,N_2219);
nand U4880 (N_4880,N_2296,N_3059);
nand U4881 (N_4881,N_3499,N_2372);
and U4882 (N_4882,N_2358,N_3080);
nand U4883 (N_4883,N_3764,N_2906);
xnor U4884 (N_4884,N_3535,N_3354);
nor U4885 (N_4885,N_2268,N_3623);
nor U4886 (N_4886,N_2610,N_3246);
nor U4887 (N_4887,N_3195,N_3561);
xor U4888 (N_4888,N_3170,N_3390);
and U4889 (N_4889,N_3294,N_2029);
or U4890 (N_4890,N_2339,N_3237);
nor U4891 (N_4891,N_2537,N_3339);
or U4892 (N_4892,N_2624,N_2595);
nor U4893 (N_4893,N_2663,N_2191);
and U4894 (N_4894,N_2529,N_3735);
nor U4895 (N_4895,N_2601,N_2121);
and U4896 (N_4896,N_3055,N_2189);
and U4897 (N_4897,N_3873,N_2264);
xor U4898 (N_4898,N_2915,N_3807);
nor U4899 (N_4899,N_2760,N_2285);
nor U4900 (N_4900,N_3955,N_3676);
or U4901 (N_4901,N_2919,N_2318);
xnor U4902 (N_4902,N_2699,N_2947);
nand U4903 (N_4903,N_2290,N_2404);
nand U4904 (N_4904,N_3558,N_3267);
xor U4905 (N_4905,N_2888,N_2758);
nor U4906 (N_4906,N_2633,N_2196);
or U4907 (N_4907,N_2885,N_2600);
or U4908 (N_4908,N_3546,N_2734);
and U4909 (N_4909,N_2908,N_3686);
nand U4910 (N_4910,N_2124,N_2940);
nor U4911 (N_4911,N_2014,N_3284);
nor U4912 (N_4912,N_3808,N_3503);
nand U4913 (N_4913,N_3264,N_3084);
or U4914 (N_4914,N_2951,N_2208);
and U4915 (N_4915,N_3415,N_2442);
and U4916 (N_4916,N_2443,N_3406);
and U4917 (N_4917,N_3756,N_2046);
xor U4918 (N_4918,N_3213,N_2094);
nand U4919 (N_4919,N_3428,N_3867);
xnor U4920 (N_4920,N_3614,N_3385);
nand U4921 (N_4921,N_3889,N_2297);
xor U4922 (N_4922,N_2890,N_2650);
nand U4923 (N_4923,N_3331,N_2446);
and U4924 (N_4924,N_3048,N_3261);
and U4925 (N_4925,N_2642,N_3159);
xor U4926 (N_4926,N_2590,N_3137);
or U4927 (N_4927,N_3725,N_3777);
and U4928 (N_4928,N_3145,N_3804);
or U4929 (N_4929,N_2931,N_3214);
xnor U4930 (N_4930,N_2476,N_2654);
nand U4931 (N_4931,N_3956,N_3005);
xor U4932 (N_4932,N_3834,N_3774);
nand U4933 (N_4933,N_2320,N_2314);
and U4934 (N_4934,N_3125,N_2467);
xnor U4935 (N_4935,N_2966,N_3344);
nor U4936 (N_4936,N_3866,N_3282);
nor U4937 (N_4937,N_2206,N_3109);
and U4938 (N_4938,N_3692,N_3186);
nor U4939 (N_4939,N_2365,N_2016);
nand U4940 (N_4940,N_2614,N_2340);
and U4941 (N_4941,N_3651,N_3117);
xor U4942 (N_4942,N_3662,N_3404);
and U4943 (N_4943,N_3520,N_3566);
xor U4944 (N_4944,N_3477,N_2569);
nand U4945 (N_4945,N_3961,N_3531);
nor U4946 (N_4946,N_2262,N_2406);
xnor U4947 (N_4947,N_3864,N_2368);
nor U4948 (N_4948,N_3829,N_3044);
and U4949 (N_4949,N_3326,N_2572);
nor U4950 (N_4950,N_3984,N_3144);
or U4951 (N_4951,N_2304,N_3698);
nor U4952 (N_4952,N_3311,N_3526);
or U4953 (N_4953,N_3946,N_3800);
nand U4954 (N_4954,N_3750,N_3996);
nand U4955 (N_4955,N_2720,N_2343);
xor U4956 (N_4956,N_2407,N_2241);
xor U4957 (N_4957,N_2399,N_2802);
xor U4958 (N_4958,N_3215,N_2088);
or U4959 (N_4959,N_2496,N_3947);
and U4960 (N_4960,N_3897,N_3787);
nand U4961 (N_4961,N_2463,N_2751);
and U4962 (N_4962,N_2987,N_3265);
or U4963 (N_4963,N_2976,N_3136);
or U4964 (N_4964,N_2698,N_3335);
nand U4965 (N_4965,N_2670,N_2500);
nor U4966 (N_4966,N_3383,N_2954);
and U4967 (N_4967,N_3492,N_3451);
or U4968 (N_4968,N_2726,N_3011);
or U4969 (N_4969,N_3541,N_2013);
and U4970 (N_4970,N_3064,N_3979);
nor U4971 (N_4971,N_3229,N_2639);
nor U4972 (N_4972,N_2135,N_2771);
nand U4973 (N_4973,N_2018,N_2326);
nor U4974 (N_4974,N_3716,N_3909);
nand U4975 (N_4975,N_3471,N_2004);
and U4976 (N_4976,N_2394,N_3779);
nor U4977 (N_4977,N_2003,N_2499);
nor U4978 (N_4978,N_2160,N_2085);
and U4979 (N_4979,N_3920,N_2017);
nor U4980 (N_4980,N_2175,N_2461);
nor U4981 (N_4981,N_3338,N_2180);
nand U4982 (N_4982,N_3978,N_3367);
nand U4983 (N_4983,N_3529,N_3595);
nand U4984 (N_4984,N_3362,N_2922);
and U4985 (N_4985,N_3998,N_3388);
and U4986 (N_4986,N_2928,N_3204);
and U4987 (N_4987,N_3082,N_2978);
nand U4988 (N_4988,N_2345,N_3027);
nor U4989 (N_4989,N_2089,N_3045);
nor U4990 (N_4990,N_3036,N_2592);
and U4991 (N_4991,N_3373,N_3513);
xor U4992 (N_4992,N_2424,N_3968);
nand U4993 (N_4993,N_2490,N_2975);
nor U4994 (N_4994,N_3636,N_3510);
nor U4995 (N_4995,N_2236,N_3312);
nand U4996 (N_4996,N_3597,N_2836);
nand U4997 (N_4997,N_3425,N_3678);
nor U4998 (N_4998,N_3095,N_3163);
xnor U4999 (N_4999,N_2076,N_2081);
or U5000 (N_5000,N_3043,N_2634);
nand U5001 (N_5001,N_2698,N_3245);
nor U5002 (N_5002,N_3383,N_2597);
nand U5003 (N_5003,N_3514,N_3436);
nor U5004 (N_5004,N_2606,N_2746);
nor U5005 (N_5005,N_2823,N_3121);
nor U5006 (N_5006,N_2807,N_3093);
nor U5007 (N_5007,N_3624,N_3598);
nor U5008 (N_5008,N_2775,N_2501);
xor U5009 (N_5009,N_3368,N_2040);
nor U5010 (N_5010,N_2346,N_2416);
nor U5011 (N_5011,N_2144,N_2154);
nor U5012 (N_5012,N_3200,N_2342);
or U5013 (N_5013,N_3334,N_3786);
xor U5014 (N_5014,N_2882,N_3484);
nand U5015 (N_5015,N_3357,N_2591);
and U5016 (N_5016,N_3856,N_3194);
and U5017 (N_5017,N_2453,N_3778);
or U5018 (N_5018,N_3411,N_2329);
or U5019 (N_5019,N_3709,N_2799);
nand U5020 (N_5020,N_2658,N_3742);
and U5021 (N_5021,N_3663,N_3180);
nand U5022 (N_5022,N_2030,N_3934);
nand U5023 (N_5023,N_3346,N_3295);
or U5024 (N_5024,N_2998,N_2878);
or U5025 (N_5025,N_3872,N_3800);
or U5026 (N_5026,N_2468,N_2256);
nand U5027 (N_5027,N_3699,N_3954);
or U5028 (N_5028,N_2912,N_2345);
or U5029 (N_5029,N_3469,N_2377);
and U5030 (N_5030,N_3345,N_2871);
xnor U5031 (N_5031,N_2757,N_3058);
and U5032 (N_5032,N_2641,N_3222);
or U5033 (N_5033,N_2381,N_2112);
xor U5034 (N_5034,N_2717,N_2321);
or U5035 (N_5035,N_2935,N_2743);
nand U5036 (N_5036,N_2616,N_3200);
nor U5037 (N_5037,N_2983,N_2470);
or U5038 (N_5038,N_3036,N_3369);
and U5039 (N_5039,N_3838,N_2892);
xnor U5040 (N_5040,N_2272,N_3759);
or U5041 (N_5041,N_3025,N_3314);
and U5042 (N_5042,N_3809,N_3492);
and U5043 (N_5043,N_2076,N_3202);
and U5044 (N_5044,N_3348,N_2224);
nand U5045 (N_5045,N_3975,N_2982);
nor U5046 (N_5046,N_3760,N_2838);
nor U5047 (N_5047,N_2447,N_3493);
and U5048 (N_5048,N_3366,N_2377);
xor U5049 (N_5049,N_2814,N_2067);
or U5050 (N_5050,N_3985,N_3322);
xnor U5051 (N_5051,N_3457,N_2839);
nand U5052 (N_5052,N_3008,N_3047);
nand U5053 (N_5053,N_2509,N_2811);
nand U5054 (N_5054,N_3265,N_2539);
nand U5055 (N_5055,N_2369,N_3877);
nand U5056 (N_5056,N_2630,N_3735);
nand U5057 (N_5057,N_3374,N_2453);
nand U5058 (N_5058,N_2280,N_3471);
or U5059 (N_5059,N_3748,N_2351);
nor U5060 (N_5060,N_2040,N_3949);
nand U5061 (N_5061,N_2740,N_2337);
and U5062 (N_5062,N_3861,N_3592);
and U5063 (N_5063,N_3233,N_3064);
nand U5064 (N_5064,N_2674,N_2698);
nor U5065 (N_5065,N_2991,N_3854);
or U5066 (N_5066,N_2936,N_3791);
or U5067 (N_5067,N_3255,N_3887);
or U5068 (N_5068,N_2422,N_2998);
xor U5069 (N_5069,N_3803,N_3165);
xnor U5070 (N_5070,N_3212,N_3783);
and U5071 (N_5071,N_2503,N_2282);
and U5072 (N_5072,N_3352,N_2332);
or U5073 (N_5073,N_3588,N_2392);
nand U5074 (N_5074,N_3293,N_2050);
nor U5075 (N_5075,N_2780,N_3292);
xnor U5076 (N_5076,N_3026,N_3087);
nor U5077 (N_5077,N_3545,N_2562);
nand U5078 (N_5078,N_3726,N_3386);
nand U5079 (N_5079,N_2673,N_2928);
nand U5080 (N_5080,N_2280,N_2012);
or U5081 (N_5081,N_3009,N_3892);
xnor U5082 (N_5082,N_2186,N_2609);
nand U5083 (N_5083,N_2057,N_2192);
xnor U5084 (N_5084,N_3909,N_2494);
or U5085 (N_5085,N_3615,N_3101);
xor U5086 (N_5086,N_2823,N_3997);
xor U5087 (N_5087,N_3334,N_2355);
nor U5088 (N_5088,N_3555,N_3535);
nor U5089 (N_5089,N_2914,N_2582);
and U5090 (N_5090,N_2478,N_2558);
nor U5091 (N_5091,N_3332,N_3719);
xnor U5092 (N_5092,N_3595,N_2737);
and U5093 (N_5093,N_3125,N_2239);
xnor U5094 (N_5094,N_3810,N_3820);
xor U5095 (N_5095,N_3612,N_3963);
or U5096 (N_5096,N_2441,N_2232);
and U5097 (N_5097,N_2011,N_2558);
and U5098 (N_5098,N_3058,N_3658);
nor U5099 (N_5099,N_2840,N_3602);
and U5100 (N_5100,N_3811,N_2210);
xor U5101 (N_5101,N_3694,N_2348);
xnor U5102 (N_5102,N_3401,N_3192);
xor U5103 (N_5103,N_3551,N_3468);
or U5104 (N_5104,N_2741,N_2936);
or U5105 (N_5105,N_3284,N_2474);
and U5106 (N_5106,N_3652,N_2589);
or U5107 (N_5107,N_2596,N_3543);
and U5108 (N_5108,N_3989,N_2714);
or U5109 (N_5109,N_3023,N_3314);
nand U5110 (N_5110,N_3440,N_2411);
nand U5111 (N_5111,N_3132,N_3652);
xor U5112 (N_5112,N_3105,N_2493);
or U5113 (N_5113,N_2226,N_2206);
nand U5114 (N_5114,N_2841,N_3341);
nand U5115 (N_5115,N_2498,N_3767);
or U5116 (N_5116,N_2906,N_3854);
and U5117 (N_5117,N_3835,N_2442);
nand U5118 (N_5118,N_3789,N_2861);
xor U5119 (N_5119,N_2107,N_2969);
or U5120 (N_5120,N_3656,N_3301);
and U5121 (N_5121,N_2289,N_2474);
nor U5122 (N_5122,N_2406,N_3456);
and U5123 (N_5123,N_3033,N_2850);
nand U5124 (N_5124,N_2017,N_3361);
xor U5125 (N_5125,N_2590,N_3159);
nor U5126 (N_5126,N_2458,N_2862);
xor U5127 (N_5127,N_3708,N_2970);
nand U5128 (N_5128,N_3296,N_3515);
or U5129 (N_5129,N_3491,N_3841);
xnor U5130 (N_5130,N_3215,N_2957);
xor U5131 (N_5131,N_2480,N_3880);
or U5132 (N_5132,N_3973,N_2590);
and U5133 (N_5133,N_2616,N_2426);
xor U5134 (N_5134,N_2207,N_2594);
nor U5135 (N_5135,N_2139,N_2300);
and U5136 (N_5136,N_3762,N_3599);
xnor U5137 (N_5137,N_2138,N_3608);
and U5138 (N_5138,N_2329,N_2219);
nor U5139 (N_5139,N_3633,N_3388);
nand U5140 (N_5140,N_3276,N_3106);
xnor U5141 (N_5141,N_2212,N_3197);
or U5142 (N_5142,N_2494,N_2676);
nor U5143 (N_5143,N_2801,N_3569);
xor U5144 (N_5144,N_3294,N_3767);
nor U5145 (N_5145,N_3790,N_3973);
nor U5146 (N_5146,N_2616,N_2601);
nor U5147 (N_5147,N_3182,N_2706);
or U5148 (N_5148,N_2553,N_3077);
xor U5149 (N_5149,N_3742,N_2238);
xor U5150 (N_5150,N_3348,N_2489);
nand U5151 (N_5151,N_2680,N_3408);
and U5152 (N_5152,N_2632,N_3719);
and U5153 (N_5153,N_2474,N_2249);
xor U5154 (N_5154,N_2638,N_2043);
nand U5155 (N_5155,N_3057,N_2946);
nor U5156 (N_5156,N_3748,N_3417);
and U5157 (N_5157,N_2560,N_3710);
xor U5158 (N_5158,N_3778,N_2526);
xnor U5159 (N_5159,N_3364,N_2298);
xor U5160 (N_5160,N_2528,N_3294);
nor U5161 (N_5161,N_2332,N_3818);
nand U5162 (N_5162,N_2962,N_2756);
or U5163 (N_5163,N_3807,N_3767);
nor U5164 (N_5164,N_3159,N_2716);
and U5165 (N_5165,N_2413,N_2398);
nor U5166 (N_5166,N_2047,N_2279);
nor U5167 (N_5167,N_2047,N_3003);
nor U5168 (N_5168,N_3225,N_2278);
xnor U5169 (N_5169,N_3614,N_2882);
or U5170 (N_5170,N_2219,N_3201);
nor U5171 (N_5171,N_3718,N_3207);
xor U5172 (N_5172,N_2050,N_2591);
nor U5173 (N_5173,N_3972,N_2065);
or U5174 (N_5174,N_3985,N_3892);
or U5175 (N_5175,N_3933,N_2551);
nand U5176 (N_5176,N_3032,N_3192);
and U5177 (N_5177,N_2247,N_2362);
and U5178 (N_5178,N_2554,N_3467);
or U5179 (N_5179,N_2922,N_3171);
or U5180 (N_5180,N_2013,N_2706);
and U5181 (N_5181,N_3356,N_2927);
nand U5182 (N_5182,N_2111,N_2127);
nand U5183 (N_5183,N_3442,N_3576);
xor U5184 (N_5184,N_3640,N_3218);
nand U5185 (N_5185,N_3993,N_2544);
or U5186 (N_5186,N_3789,N_2407);
xnor U5187 (N_5187,N_3349,N_3442);
xnor U5188 (N_5188,N_2373,N_3191);
nand U5189 (N_5189,N_3178,N_3488);
nor U5190 (N_5190,N_2180,N_2921);
nor U5191 (N_5191,N_3778,N_2343);
and U5192 (N_5192,N_3906,N_2286);
or U5193 (N_5193,N_2381,N_2967);
nor U5194 (N_5194,N_3088,N_3839);
nand U5195 (N_5195,N_2539,N_2712);
nor U5196 (N_5196,N_2538,N_3165);
nor U5197 (N_5197,N_3192,N_3255);
nand U5198 (N_5198,N_3102,N_2379);
xor U5199 (N_5199,N_2911,N_2424);
or U5200 (N_5200,N_2753,N_3430);
or U5201 (N_5201,N_2666,N_3825);
nand U5202 (N_5202,N_3706,N_3343);
nor U5203 (N_5203,N_3466,N_2744);
nor U5204 (N_5204,N_2361,N_2149);
nand U5205 (N_5205,N_2816,N_2710);
nor U5206 (N_5206,N_2333,N_3488);
nand U5207 (N_5207,N_2218,N_2794);
nand U5208 (N_5208,N_2901,N_2346);
and U5209 (N_5209,N_2799,N_2308);
or U5210 (N_5210,N_2703,N_3085);
nor U5211 (N_5211,N_2538,N_2691);
or U5212 (N_5212,N_2083,N_3761);
xnor U5213 (N_5213,N_3100,N_3109);
and U5214 (N_5214,N_2957,N_3728);
nor U5215 (N_5215,N_3358,N_3339);
nand U5216 (N_5216,N_3962,N_2494);
xnor U5217 (N_5217,N_3787,N_2241);
xor U5218 (N_5218,N_2413,N_3211);
nand U5219 (N_5219,N_3304,N_2899);
xnor U5220 (N_5220,N_2103,N_3684);
or U5221 (N_5221,N_2933,N_3325);
and U5222 (N_5222,N_2641,N_3394);
and U5223 (N_5223,N_3567,N_3407);
or U5224 (N_5224,N_2543,N_2264);
nand U5225 (N_5225,N_2796,N_2424);
nand U5226 (N_5226,N_2683,N_2207);
nand U5227 (N_5227,N_2202,N_2781);
xor U5228 (N_5228,N_2618,N_2430);
or U5229 (N_5229,N_2936,N_2399);
nand U5230 (N_5230,N_3465,N_3142);
xor U5231 (N_5231,N_3641,N_3010);
nand U5232 (N_5232,N_3404,N_3873);
xnor U5233 (N_5233,N_3239,N_2683);
nor U5234 (N_5234,N_3390,N_2626);
or U5235 (N_5235,N_2749,N_3970);
xor U5236 (N_5236,N_2892,N_3683);
xnor U5237 (N_5237,N_3586,N_3300);
nor U5238 (N_5238,N_3037,N_2238);
or U5239 (N_5239,N_3219,N_3176);
or U5240 (N_5240,N_3606,N_2942);
and U5241 (N_5241,N_2453,N_3651);
or U5242 (N_5242,N_3341,N_2056);
nand U5243 (N_5243,N_3352,N_3699);
nor U5244 (N_5244,N_3941,N_3284);
or U5245 (N_5245,N_3397,N_3102);
or U5246 (N_5246,N_3161,N_3544);
and U5247 (N_5247,N_2354,N_3501);
nand U5248 (N_5248,N_3486,N_3148);
nor U5249 (N_5249,N_2188,N_2241);
nand U5250 (N_5250,N_3919,N_2603);
and U5251 (N_5251,N_3902,N_2041);
nand U5252 (N_5252,N_3587,N_2191);
nor U5253 (N_5253,N_3098,N_3440);
xnor U5254 (N_5254,N_3399,N_2991);
nor U5255 (N_5255,N_3079,N_3497);
or U5256 (N_5256,N_3980,N_3526);
or U5257 (N_5257,N_2472,N_2220);
nor U5258 (N_5258,N_3624,N_3806);
nor U5259 (N_5259,N_3277,N_2503);
nor U5260 (N_5260,N_2602,N_3857);
xnor U5261 (N_5261,N_3001,N_2120);
nor U5262 (N_5262,N_3133,N_3550);
and U5263 (N_5263,N_3568,N_2988);
nand U5264 (N_5264,N_3219,N_2661);
nor U5265 (N_5265,N_3556,N_3493);
nand U5266 (N_5266,N_2283,N_2122);
nor U5267 (N_5267,N_3833,N_3261);
nor U5268 (N_5268,N_3941,N_2887);
nand U5269 (N_5269,N_3468,N_3249);
xor U5270 (N_5270,N_2068,N_2552);
nand U5271 (N_5271,N_2124,N_3125);
or U5272 (N_5272,N_3156,N_3837);
nor U5273 (N_5273,N_3087,N_2538);
xnor U5274 (N_5274,N_2913,N_3572);
nor U5275 (N_5275,N_3710,N_3859);
nand U5276 (N_5276,N_2159,N_3162);
nand U5277 (N_5277,N_3320,N_2206);
nor U5278 (N_5278,N_2473,N_3289);
nand U5279 (N_5279,N_2661,N_2775);
xor U5280 (N_5280,N_2271,N_3601);
and U5281 (N_5281,N_3467,N_2012);
and U5282 (N_5282,N_2028,N_3667);
xnor U5283 (N_5283,N_2380,N_3186);
xnor U5284 (N_5284,N_2846,N_2942);
nand U5285 (N_5285,N_3345,N_3629);
xor U5286 (N_5286,N_3223,N_2323);
and U5287 (N_5287,N_2073,N_3932);
nor U5288 (N_5288,N_3125,N_2520);
nor U5289 (N_5289,N_3154,N_3168);
xnor U5290 (N_5290,N_2062,N_2933);
xor U5291 (N_5291,N_3982,N_2378);
nand U5292 (N_5292,N_2013,N_3754);
nand U5293 (N_5293,N_2465,N_2818);
xnor U5294 (N_5294,N_3034,N_3544);
xnor U5295 (N_5295,N_2946,N_3418);
nand U5296 (N_5296,N_3712,N_3876);
nand U5297 (N_5297,N_2847,N_2551);
xnor U5298 (N_5298,N_2079,N_2043);
and U5299 (N_5299,N_2716,N_3097);
nand U5300 (N_5300,N_2689,N_3411);
nand U5301 (N_5301,N_2721,N_2804);
nor U5302 (N_5302,N_2214,N_3773);
and U5303 (N_5303,N_2999,N_2376);
nand U5304 (N_5304,N_3915,N_2704);
nor U5305 (N_5305,N_3486,N_3477);
and U5306 (N_5306,N_2320,N_2787);
nor U5307 (N_5307,N_2609,N_2963);
nor U5308 (N_5308,N_2417,N_2670);
and U5309 (N_5309,N_2112,N_3556);
and U5310 (N_5310,N_2670,N_2712);
xor U5311 (N_5311,N_2487,N_2803);
xnor U5312 (N_5312,N_2343,N_2280);
and U5313 (N_5313,N_3713,N_3319);
or U5314 (N_5314,N_3198,N_2094);
and U5315 (N_5315,N_3620,N_3502);
nand U5316 (N_5316,N_3637,N_3871);
xor U5317 (N_5317,N_3891,N_2193);
xor U5318 (N_5318,N_2394,N_2891);
and U5319 (N_5319,N_2278,N_3922);
or U5320 (N_5320,N_3786,N_3853);
xor U5321 (N_5321,N_2004,N_2022);
nand U5322 (N_5322,N_2540,N_2066);
nor U5323 (N_5323,N_2383,N_2658);
and U5324 (N_5324,N_3474,N_2301);
nand U5325 (N_5325,N_3580,N_3589);
nand U5326 (N_5326,N_3298,N_3539);
or U5327 (N_5327,N_3836,N_3425);
xor U5328 (N_5328,N_3560,N_2438);
and U5329 (N_5329,N_3351,N_2136);
and U5330 (N_5330,N_2066,N_2849);
nand U5331 (N_5331,N_2428,N_3481);
nand U5332 (N_5332,N_2810,N_3809);
and U5333 (N_5333,N_3631,N_2363);
or U5334 (N_5334,N_3605,N_2473);
nor U5335 (N_5335,N_2693,N_2264);
nor U5336 (N_5336,N_3310,N_2728);
or U5337 (N_5337,N_3992,N_2838);
nor U5338 (N_5338,N_3753,N_3136);
xor U5339 (N_5339,N_3704,N_3927);
nor U5340 (N_5340,N_2523,N_2325);
nand U5341 (N_5341,N_2278,N_2451);
nand U5342 (N_5342,N_3250,N_2520);
xor U5343 (N_5343,N_2439,N_2204);
or U5344 (N_5344,N_3755,N_3951);
and U5345 (N_5345,N_2384,N_3599);
or U5346 (N_5346,N_3146,N_2202);
nand U5347 (N_5347,N_3486,N_2795);
and U5348 (N_5348,N_3156,N_2163);
or U5349 (N_5349,N_2806,N_3062);
and U5350 (N_5350,N_2563,N_3937);
nand U5351 (N_5351,N_3878,N_2276);
and U5352 (N_5352,N_3920,N_3131);
and U5353 (N_5353,N_3096,N_3256);
nor U5354 (N_5354,N_3817,N_2553);
or U5355 (N_5355,N_3603,N_2728);
xnor U5356 (N_5356,N_3407,N_2343);
or U5357 (N_5357,N_2946,N_2240);
xor U5358 (N_5358,N_2042,N_3257);
xnor U5359 (N_5359,N_2715,N_2066);
xor U5360 (N_5360,N_2334,N_3765);
or U5361 (N_5361,N_2512,N_2157);
xnor U5362 (N_5362,N_2290,N_2320);
xnor U5363 (N_5363,N_2309,N_2334);
nand U5364 (N_5364,N_3720,N_3031);
and U5365 (N_5365,N_2103,N_3355);
nand U5366 (N_5366,N_3619,N_3115);
or U5367 (N_5367,N_3272,N_3195);
or U5368 (N_5368,N_2198,N_2028);
nor U5369 (N_5369,N_3208,N_3816);
nor U5370 (N_5370,N_3334,N_3975);
xor U5371 (N_5371,N_2908,N_3761);
nor U5372 (N_5372,N_2746,N_3666);
nor U5373 (N_5373,N_2316,N_3057);
xnor U5374 (N_5374,N_3937,N_2322);
nand U5375 (N_5375,N_2500,N_2998);
nand U5376 (N_5376,N_2853,N_2059);
xor U5377 (N_5377,N_2656,N_3642);
nor U5378 (N_5378,N_3230,N_2980);
or U5379 (N_5379,N_3349,N_3005);
nand U5380 (N_5380,N_2821,N_3918);
or U5381 (N_5381,N_3619,N_3209);
nand U5382 (N_5382,N_2712,N_2406);
xnor U5383 (N_5383,N_3934,N_2326);
and U5384 (N_5384,N_3258,N_2933);
xor U5385 (N_5385,N_2412,N_2052);
xor U5386 (N_5386,N_3573,N_3515);
or U5387 (N_5387,N_2561,N_2321);
nand U5388 (N_5388,N_3168,N_2991);
nor U5389 (N_5389,N_2224,N_3867);
and U5390 (N_5390,N_3002,N_3373);
nand U5391 (N_5391,N_2151,N_3565);
and U5392 (N_5392,N_2338,N_2439);
nand U5393 (N_5393,N_2081,N_2357);
and U5394 (N_5394,N_2221,N_2288);
or U5395 (N_5395,N_2746,N_2415);
xor U5396 (N_5396,N_2306,N_2743);
xor U5397 (N_5397,N_3946,N_2048);
or U5398 (N_5398,N_3913,N_2790);
nor U5399 (N_5399,N_3981,N_3714);
or U5400 (N_5400,N_3817,N_2426);
nand U5401 (N_5401,N_3185,N_2123);
nor U5402 (N_5402,N_3763,N_2738);
nor U5403 (N_5403,N_3945,N_2956);
nand U5404 (N_5404,N_2521,N_3882);
nor U5405 (N_5405,N_3308,N_3350);
or U5406 (N_5406,N_2282,N_3695);
or U5407 (N_5407,N_3658,N_3626);
nor U5408 (N_5408,N_3236,N_2941);
nand U5409 (N_5409,N_3307,N_3291);
and U5410 (N_5410,N_3935,N_2596);
nand U5411 (N_5411,N_3653,N_2901);
xnor U5412 (N_5412,N_3933,N_2084);
and U5413 (N_5413,N_2972,N_3948);
or U5414 (N_5414,N_3045,N_3480);
nand U5415 (N_5415,N_2216,N_2661);
or U5416 (N_5416,N_2106,N_2646);
nand U5417 (N_5417,N_2647,N_3489);
nor U5418 (N_5418,N_3840,N_3140);
xnor U5419 (N_5419,N_2049,N_2657);
or U5420 (N_5420,N_2528,N_2098);
xnor U5421 (N_5421,N_2483,N_3734);
and U5422 (N_5422,N_2538,N_3181);
and U5423 (N_5423,N_2938,N_2089);
and U5424 (N_5424,N_3025,N_3967);
nor U5425 (N_5425,N_2712,N_2843);
xor U5426 (N_5426,N_2309,N_3613);
nand U5427 (N_5427,N_2354,N_2821);
xnor U5428 (N_5428,N_2805,N_2522);
nor U5429 (N_5429,N_3465,N_2464);
xnor U5430 (N_5430,N_3555,N_3196);
nand U5431 (N_5431,N_3140,N_2184);
and U5432 (N_5432,N_2103,N_3068);
or U5433 (N_5433,N_2443,N_2426);
or U5434 (N_5434,N_3312,N_3973);
nor U5435 (N_5435,N_2417,N_3054);
nand U5436 (N_5436,N_3792,N_2191);
nand U5437 (N_5437,N_3779,N_3203);
or U5438 (N_5438,N_3416,N_2541);
nand U5439 (N_5439,N_2543,N_3586);
nand U5440 (N_5440,N_3753,N_3807);
xor U5441 (N_5441,N_3528,N_2606);
nand U5442 (N_5442,N_2752,N_3304);
nor U5443 (N_5443,N_3854,N_2705);
nor U5444 (N_5444,N_2086,N_3505);
nor U5445 (N_5445,N_3702,N_3773);
and U5446 (N_5446,N_3363,N_3365);
xor U5447 (N_5447,N_3343,N_2991);
nand U5448 (N_5448,N_2879,N_2119);
or U5449 (N_5449,N_3543,N_3879);
nor U5450 (N_5450,N_3107,N_2385);
or U5451 (N_5451,N_3426,N_3036);
and U5452 (N_5452,N_2723,N_3403);
nand U5453 (N_5453,N_2918,N_3457);
and U5454 (N_5454,N_2367,N_2069);
xnor U5455 (N_5455,N_2821,N_3829);
nand U5456 (N_5456,N_3327,N_2045);
xnor U5457 (N_5457,N_2159,N_3021);
and U5458 (N_5458,N_3535,N_2588);
xor U5459 (N_5459,N_3974,N_3456);
nand U5460 (N_5460,N_2451,N_3114);
or U5461 (N_5461,N_3005,N_3299);
and U5462 (N_5462,N_2814,N_2327);
nand U5463 (N_5463,N_2239,N_3940);
nor U5464 (N_5464,N_3211,N_2309);
nand U5465 (N_5465,N_2971,N_3835);
xnor U5466 (N_5466,N_2341,N_2971);
nor U5467 (N_5467,N_3257,N_2825);
xnor U5468 (N_5468,N_3600,N_2217);
nand U5469 (N_5469,N_3590,N_2479);
nand U5470 (N_5470,N_3223,N_3866);
xnor U5471 (N_5471,N_2663,N_3440);
xor U5472 (N_5472,N_2616,N_2342);
nand U5473 (N_5473,N_2376,N_2776);
or U5474 (N_5474,N_3631,N_2946);
xnor U5475 (N_5475,N_3486,N_3298);
or U5476 (N_5476,N_2897,N_2810);
nand U5477 (N_5477,N_3366,N_2843);
xor U5478 (N_5478,N_2987,N_3435);
nor U5479 (N_5479,N_2693,N_2796);
or U5480 (N_5480,N_3056,N_3522);
or U5481 (N_5481,N_3757,N_3473);
or U5482 (N_5482,N_3276,N_3909);
nor U5483 (N_5483,N_3605,N_2805);
nand U5484 (N_5484,N_2376,N_2852);
and U5485 (N_5485,N_2821,N_2681);
nand U5486 (N_5486,N_2118,N_2452);
nand U5487 (N_5487,N_2659,N_3665);
xnor U5488 (N_5488,N_2911,N_2736);
or U5489 (N_5489,N_3505,N_3433);
nor U5490 (N_5490,N_3394,N_3646);
or U5491 (N_5491,N_3483,N_3053);
and U5492 (N_5492,N_3776,N_2573);
xor U5493 (N_5493,N_3181,N_2055);
and U5494 (N_5494,N_2578,N_3732);
or U5495 (N_5495,N_3011,N_2523);
and U5496 (N_5496,N_2481,N_3470);
and U5497 (N_5497,N_3953,N_2037);
xnor U5498 (N_5498,N_2917,N_3897);
or U5499 (N_5499,N_2607,N_2820);
nor U5500 (N_5500,N_2771,N_2029);
nor U5501 (N_5501,N_2710,N_3731);
nand U5502 (N_5502,N_2981,N_2157);
nand U5503 (N_5503,N_2258,N_2395);
nor U5504 (N_5504,N_3470,N_2014);
nor U5505 (N_5505,N_2548,N_3758);
xor U5506 (N_5506,N_2185,N_3547);
xor U5507 (N_5507,N_2312,N_3677);
or U5508 (N_5508,N_3530,N_3082);
xor U5509 (N_5509,N_3945,N_2887);
or U5510 (N_5510,N_2124,N_3228);
and U5511 (N_5511,N_2992,N_3489);
and U5512 (N_5512,N_2085,N_3137);
and U5513 (N_5513,N_3944,N_2162);
nor U5514 (N_5514,N_3086,N_2355);
nor U5515 (N_5515,N_3261,N_3707);
xnor U5516 (N_5516,N_3903,N_3351);
xnor U5517 (N_5517,N_2206,N_2307);
and U5518 (N_5518,N_3762,N_3535);
nor U5519 (N_5519,N_3660,N_3037);
nand U5520 (N_5520,N_3437,N_2711);
nand U5521 (N_5521,N_2179,N_2819);
or U5522 (N_5522,N_2855,N_2293);
nand U5523 (N_5523,N_3068,N_3752);
and U5524 (N_5524,N_2590,N_2519);
and U5525 (N_5525,N_3192,N_3592);
nand U5526 (N_5526,N_2088,N_2855);
nand U5527 (N_5527,N_3018,N_2127);
nor U5528 (N_5528,N_2414,N_2151);
xor U5529 (N_5529,N_3211,N_3199);
nand U5530 (N_5530,N_2972,N_3100);
nor U5531 (N_5531,N_3865,N_3000);
and U5532 (N_5532,N_2579,N_3218);
nor U5533 (N_5533,N_2394,N_3322);
nor U5534 (N_5534,N_2974,N_3280);
and U5535 (N_5535,N_3083,N_2488);
and U5536 (N_5536,N_3605,N_3483);
nor U5537 (N_5537,N_3215,N_2689);
xor U5538 (N_5538,N_3556,N_2073);
nor U5539 (N_5539,N_2424,N_3908);
xnor U5540 (N_5540,N_3537,N_2776);
xor U5541 (N_5541,N_2334,N_3999);
or U5542 (N_5542,N_2062,N_3500);
and U5543 (N_5543,N_3557,N_3179);
nand U5544 (N_5544,N_2225,N_3034);
nand U5545 (N_5545,N_2234,N_3415);
nor U5546 (N_5546,N_2003,N_2613);
xnor U5547 (N_5547,N_2040,N_2613);
nor U5548 (N_5548,N_2623,N_2510);
nor U5549 (N_5549,N_2211,N_3112);
xnor U5550 (N_5550,N_2217,N_2092);
or U5551 (N_5551,N_2328,N_3847);
and U5552 (N_5552,N_2127,N_2982);
and U5553 (N_5553,N_2063,N_2146);
nor U5554 (N_5554,N_3550,N_2049);
and U5555 (N_5555,N_2290,N_3264);
nor U5556 (N_5556,N_2187,N_3299);
or U5557 (N_5557,N_3274,N_2036);
and U5558 (N_5558,N_3440,N_2077);
nand U5559 (N_5559,N_3730,N_2745);
and U5560 (N_5560,N_2048,N_2964);
and U5561 (N_5561,N_3803,N_3271);
or U5562 (N_5562,N_3674,N_3853);
or U5563 (N_5563,N_3945,N_2001);
and U5564 (N_5564,N_3054,N_3558);
and U5565 (N_5565,N_2613,N_2793);
nand U5566 (N_5566,N_3092,N_2571);
xnor U5567 (N_5567,N_3818,N_3930);
nor U5568 (N_5568,N_2027,N_2818);
and U5569 (N_5569,N_3434,N_2878);
or U5570 (N_5570,N_2152,N_3229);
or U5571 (N_5571,N_3993,N_2234);
or U5572 (N_5572,N_2100,N_2801);
xnor U5573 (N_5573,N_3809,N_3579);
xor U5574 (N_5574,N_2364,N_3878);
or U5575 (N_5575,N_2937,N_3680);
nor U5576 (N_5576,N_2216,N_3585);
or U5577 (N_5577,N_2182,N_2306);
and U5578 (N_5578,N_3786,N_2762);
xnor U5579 (N_5579,N_2218,N_2172);
nor U5580 (N_5580,N_3099,N_2534);
or U5581 (N_5581,N_3296,N_2181);
xnor U5582 (N_5582,N_2017,N_3722);
nand U5583 (N_5583,N_2956,N_2156);
nand U5584 (N_5584,N_2761,N_3250);
nor U5585 (N_5585,N_2223,N_3613);
or U5586 (N_5586,N_2067,N_2612);
and U5587 (N_5587,N_3129,N_2051);
nor U5588 (N_5588,N_2223,N_3162);
and U5589 (N_5589,N_2241,N_3701);
xor U5590 (N_5590,N_3970,N_3445);
nor U5591 (N_5591,N_3488,N_2096);
nor U5592 (N_5592,N_2116,N_3910);
nor U5593 (N_5593,N_3442,N_2503);
xnor U5594 (N_5594,N_3305,N_2604);
or U5595 (N_5595,N_3375,N_3996);
nand U5596 (N_5596,N_3173,N_3228);
nor U5597 (N_5597,N_3589,N_3806);
or U5598 (N_5598,N_2213,N_2171);
and U5599 (N_5599,N_2883,N_3093);
and U5600 (N_5600,N_2778,N_2290);
xnor U5601 (N_5601,N_3795,N_2247);
and U5602 (N_5602,N_3993,N_2108);
and U5603 (N_5603,N_2373,N_3049);
or U5604 (N_5604,N_2589,N_3804);
nor U5605 (N_5605,N_2219,N_3384);
xnor U5606 (N_5606,N_2529,N_3791);
or U5607 (N_5607,N_2437,N_3486);
xnor U5608 (N_5608,N_2120,N_3219);
and U5609 (N_5609,N_3305,N_3458);
xnor U5610 (N_5610,N_2457,N_2429);
nor U5611 (N_5611,N_3913,N_2146);
nand U5612 (N_5612,N_3810,N_3451);
or U5613 (N_5613,N_2416,N_3065);
or U5614 (N_5614,N_3394,N_2940);
or U5615 (N_5615,N_3667,N_2423);
xnor U5616 (N_5616,N_3042,N_2490);
nor U5617 (N_5617,N_2021,N_2925);
and U5618 (N_5618,N_2772,N_3490);
nor U5619 (N_5619,N_3189,N_2564);
or U5620 (N_5620,N_3826,N_2884);
nor U5621 (N_5621,N_2898,N_2396);
or U5622 (N_5622,N_2434,N_2481);
or U5623 (N_5623,N_3551,N_3364);
xnor U5624 (N_5624,N_2240,N_2193);
xnor U5625 (N_5625,N_3647,N_3004);
nor U5626 (N_5626,N_2359,N_2237);
or U5627 (N_5627,N_2355,N_2933);
nand U5628 (N_5628,N_3651,N_3285);
nor U5629 (N_5629,N_2692,N_2008);
nand U5630 (N_5630,N_2625,N_2176);
nor U5631 (N_5631,N_2519,N_3567);
xnor U5632 (N_5632,N_3150,N_2744);
nor U5633 (N_5633,N_3092,N_3299);
nor U5634 (N_5634,N_2930,N_3159);
xnor U5635 (N_5635,N_3064,N_3696);
xor U5636 (N_5636,N_3720,N_3356);
nor U5637 (N_5637,N_2825,N_2081);
and U5638 (N_5638,N_3920,N_2074);
or U5639 (N_5639,N_2835,N_2564);
xor U5640 (N_5640,N_2423,N_2372);
and U5641 (N_5641,N_3773,N_2272);
nand U5642 (N_5642,N_3095,N_2530);
xor U5643 (N_5643,N_2691,N_2311);
and U5644 (N_5644,N_3064,N_3225);
and U5645 (N_5645,N_3738,N_2002);
nand U5646 (N_5646,N_3179,N_2197);
nand U5647 (N_5647,N_2398,N_3268);
xnor U5648 (N_5648,N_3437,N_3109);
or U5649 (N_5649,N_3482,N_3234);
or U5650 (N_5650,N_3005,N_3474);
nand U5651 (N_5651,N_3307,N_3464);
xnor U5652 (N_5652,N_2791,N_3061);
or U5653 (N_5653,N_3638,N_3854);
xnor U5654 (N_5654,N_2008,N_3524);
xor U5655 (N_5655,N_3143,N_3247);
xor U5656 (N_5656,N_3967,N_3886);
xnor U5657 (N_5657,N_2343,N_2872);
nor U5658 (N_5658,N_3635,N_2182);
nand U5659 (N_5659,N_2806,N_3651);
nor U5660 (N_5660,N_3164,N_3312);
nor U5661 (N_5661,N_3567,N_3215);
xnor U5662 (N_5662,N_2099,N_3043);
nand U5663 (N_5663,N_3471,N_2330);
nor U5664 (N_5664,N_3410,N_3777);
nand U5665 (N_5665,N_2857,N_2147);
nand U5666 (N_5666,N_3141,N_3352);
or U5667 (N_5667,N_3980,N_2368);
or U5668 (N_5668,N_3536,N_3017);
and U5669 (N_5669,N_3991,N_2521);
xor U5670 (N_5670,N_3162,N_2213);
nand U5671 (N_5671,N_3956,N_2901);
nand U5672 (N_5672,N_2731,N_3923);
nand U5673 (N_5673,N_3430,N_2505);
xor U5674 (N_5674,N_3680,N_3136);
nor U5675 (N_5675,N_2456,N_3279);
or U5676 (N_5676,N_3227,N_3629);
or U5677 (N_5677,N_2740,N_3000);
xnor U5678 (N_5678,N_2608,N_2346);
nand U5679 (N_5679,N_3683,N_3292);
and U5680 (N_5680,N_2526,N_2905);
or U5681 (N_5681,N_2108,N_3676);
nand U5682 (N_5682,N_2971,N_2412);
xor U5683 (N_5683,N_2698,N_3264);
or U5684 (N_5684,N_3976,N_2961);
and U5685 (N_5685,N_3128,N_2719);
xor U5686 (N_5686,N_3486,N_2452);
nand U5687 (N_5687,N_3771,N_2139);
nand U5688 (N_5688,N_3899,N_3190);
nor U5689 (N_5689,N_3482,N_2800);
nor U5690 (N_5690,N_2861,N_2311);
or U5691 (N_5691,N_3024,N_3699);
xnor U5692 (N_5692,N_3649,N_3737);
and U5693 (N_5693,N_2783,N_2954);
nand U5694 (N_5694,N_2154,N_3114);
or U5695 (N_5695,N_2994,N_3010);
or U5696 (N_5696,N_3651,N_3375);
and U5697 (N_5697,N_3727,N_2590);
nor U5698 (N_5698,N_3795,N_3033);
and U5699 (N_5699,N_3897,N_3712);
nor U5700 (N_5700,N_2303,N_2593);
and U5701 (N_5701,N_2803,N_2373);
and U5702 (N_5702,N_3485,N_2748);
nand U5703 (N_5703,N_3709,N_2288);
xnor U5704 (N_5704,N_2827,N_2141);
xor U5705 (N_5705,N_3965,N_3100);
or U5706 (N_5706,N_3664,N_3799);
nand U5707 (N_5707,N_2354,N_2252);
xor U5708 (N_5708,N_2786,N_3001);
and U5709 (N_5709,N_3270,N_2519);
and U5710 (N_5710,N_3259,N_3207);
or U5711 (N_5711,N_3341,N_2708);
nor U5712 (N_5712,N_3588,N_2149);
and U5713 (N_5713,N_3067,N_2894);
nand U5714 (N_5714,N_3649,N_2261);
xnor U5715 (N_5715,N_3000,N_3426);
nor U5716 (N_5716,N_3798,N_2401);
xor U5717 (N_5717,N_2765,N_2422);
and U5718 (N_5718,N_3480,N_2599);
nor U5719 (N_5719,N_2962,N_2414);
nor U5720 (N_5720,N_2701,N_2769);
nor U5721 (N_5721,N_3869,N_2700);
nand U5722 (N_5722,N_3695,N_2111);
or U5723 (N_5723,N_3965,N_3499);
nand U5724 (N_5724,N_2740,N_2405);
and U5725 (N_5725,N_2758,N_3358);
nand U5726 (N_5726,N_2713,N_2790);
and U5727 (N_5727,N_2554,N_2055);
nor U5728 (N_5728,N_2257,N_2677);
or U5729 (N_5729,N_3617,N_3603);
nand U5730 (N_5730,N_2128,N_3604);
nor U5731 (N_5731,N_2444,N_3163);
xnor U5732 (N_5732,N_2199,N_2432);
xor U5733 (N_5733,N_3134,N_2035);
nor U5734 (N_5734,N_3054,N_3933);
xnor U5735 (N_5735,N_3329,N_2638);
or U5736 (N_5736,N_3339,N_3284);
or U5737 (N_5737,N_2016,N_3507);
or U5738 (N_5738,N_2055,N_2107);
or U5739 (N_5739,N_2490,N_3414);
xnor U5740 (N_5740,N_3715,N_3667);
nor U5741 (N_5741,N_3202,N_2349);
or U5742 (N_5742,N_2270,N_2418);
or U5743 (N_5743,N_2856,N_2045);
nand U5744 (N_5744,N_2800,N_2617);
xnor U5745 (N_5745,N_2119,N_3301);
nor U5746 (N_5746,N_2375,N_2892);
or U5747 (N_5747,N_3319,N_3369);
nand U5748 (N_5748,N_3516,N_3594);
xnor U5749 (N_5749,N_2378,N_3512);
nand U5750 (N_5750,N_2969,N_3470);
or U5751 (N_5751,N_2513,N_3687);
nor U5752 (N_5752,N_2977,N_2927);
nand U5753 (N_5753,N_2272,N_2802);
and U5754 (N_5754,N_3018,N_2890);
or U5755 (N_5755,N_3306,N_3528);
nor U5756 (N_5756,N_2113,N_2762);
xnor U5757 (N_5757,N_3632,N_2152);
xnor U5758 (N_5758,N_3437,N_2662);
and U5759 (N_5759,N_2184,N_3018);
xor U5760 (N_5760,N_2066,N_3748);
xor U5761 (N_5761,N_2198,N_3231);
or U5762 (N_5762,N_2448,N_3794);
xor U5763 (N_5763,N_3094,N_3692);
and U5764 (N_5764,N_3856,N_3958);
or U5765 (N_5765,N_3824,N_2546);
and U5766 (N_5766,N_2429,N_2309);
xnor U5767 (N_5767,N_2707,N_3910);
xor U5768 (N_5768,N_3572,N_3280);
nor U5769 (N_5769,N_2118,N_2634);
nor U5770 (N_5770,N_3291,N_2090);
nand U5771 (N_5771,N_2944,N_2339);
or U5772 (N_5772,N_2503,N_2093);
nand U5773 (N_5773,N_3909,N_2464);
or U5774 (N_5774,N_3643,N_3761);
nand U5775 (N_5775,N_3729,N_2463);
nor U5776 (N_5776,N_3611,N_2128);
nor U5777 (N_5777,N_2379,N_2296);
nand U5778 (N_5778,N_3275,N_3723);
and U5779 (N_5779,N_2738,N_3855);
and U5780 (N_5780,N_3825,N_2508);
and U5781 (N_5781,N_3622,N_3279);
nand U5782 (N_5782,N_3822,N_2249);
and U5783 (N_5783,N_2059,N_3625);
nand U5784 (N_5784,N_3675,N_3961);
and U5785 (N_5785,N_2121,N_3057);
xnor U5786 (N_5786,N_2337,N_2441);
nor U5787 (N_5787,N_2515,N_3328);
or U5788 (N_5788,N_2743,N_3437);
nand U5789 (N_5789,N_2289,N_2761);
and U5790 (N_5790,N_3220,N_3985);
or U5791 (N_5791,N_3115,N_3141);
and U5792 (N_5792,N_2397,N_2497);
nand U5793 (N_5793,N_3411,N_3703);
nor U5794 (N_5794,N_2292,N_2438);
nand U5795 (N_5795,N_3933,N_3382);
xor U5796 (N_5796,N_3982,N_2870);
nor U5797 (N_5797,N_2218,N_3740);
xor U5798 (N_5798,N_3914,N_3909);
or U5799 (N_5799,N_3850,N_2153);
or U5800 (N_5800,N_2347,N_3319);
nor U5801 (N_5801,N_2703,N_3354);
xor U5802 (N_5802,N_2660,N_2513);
and U5803 (N_5803,N_2739,N_2850);
nand U5804 (N_5804,N_2046,N_2031);
or U5805 (N_5805,N_3298,N_3630);
xor U5806 (N_5806,N_2814,N_2731);
nand U5807 (N_5807,N_3048,N_3033);
xnor U5808 (N_5808,N_3968,N_3972);
xor U5809 (N_5809,N_3452,N_3184);
or U5810 (N_5810,N_2642,N_2587);
and U5811 (N_5811,N_3117,N_3347);
xnor U5812 (N_5812,N_2944,N_2573);
or U5813 (N_5813,N_3350,N_2526);
or U5814 (N_5814,N_2029,N_3678);
nor U5815 (N_5815,N_2099,N_3969);
and U5816 (N_5816,N_2251,N_2288);
or U5817 (N_5817,N_3405,N_2223);
nand U5818 (N_5818,N_2061,N_3696);
xor U5819 (N_5819,N_2427,N_2948);
xor U5820 (N_5820,N_2444,N_3382);
or U5821 (N_5821,N_3884,N_3090);
or U5822 (N_5822,N_3244,N_3465);
xnor U5823 (N_5823,N_3744,N_2303);
xnor U5824 (N_5824,N_3146,N_2034);
and U5825 (N_5825,N_3996,N_3258);
nor U5826 (N_5826,N_2416,N_3515);
xnor U5827 (N_5827,N_3954,N_3626);
and U5828 (N_5828,N_2985,N_2610);
or U5829 (N_5829,N_3135,N_2647);
and U5830 (N_5830,N_3902,N_2609);
nand U5831 (N_5831,N_3089,N_2634);
and U5832 (N_5832,N_3754,N_2104);
nand U5833 (N_5833,N_3416,N_2422);
and U5834 (N_5834,N_2419,N_2980);
and U5835 (N_5835,N_2594,N_3783);
and U5836 (N_5836,N_3051,N_2163);
and U5837 (N_5837,N_3119,N_3963);
and U5838 (N_5838,N_3583,N_2139);
xor U5839 (N_5839,N_2371,N_3811);
nor U5840 (N_5840,N_2586,N_3058);
or U5841 (N_5841,N_3337,N_3554);
or U5842 (N_5842,N_3231,N_2749);
or U5843 (N_5843,N_2540,N_3714);
nand U5844 (N_5844,N_2561,N_2078);
and U5845 (N_5845,N_2641,N_2002);
and U5846 (N_5846,N_3963,N_3497);
xor U5847 (N_5847,N_3141,N_2604);
nand U5848 (N_5848,N_2289,N_2781);
or U5849 (N_5849,N_2824,N_3574);
xnor U5850 (N_5850,N_3767,N_3677);
nor U5851 (N_5851,N_3179,N_2978);
or U5852 (N_5852,N_3188,N_3621);
or U5853 (N_5853,N_3430,N_3108);
xor U5854 (N_5854,N_3830,N_3453);
nand U5855 (N_5855,N_2585,N_3055);
nor U5856 (N_5856,N_3572,N_2227);
nand U5857 (N_5857,N_2646,N_2712);
nor U5858 (N_5858,N_2791,N_3015);
or U5859 (N_5859,N_2044,N_3537);
or U5860 (N_5860,N_2345,N_2611);
xnor U5861 (N_5861,N_3047,N_3175);
nor U5862 (N_5862,N_2806,N_2464);
xnor U5863 (N_5863,N_2281,N_3143);
nand U5864 (N_5864,N_3292,N_2480);
and U5865 (N_5865,N_2918,N_2324);
nor U5866 (N_5866,N_2899,N_2890);
xor U5867 (N_5867,N_2931,N_2312);
nor U5868 (N_5868,N_2745,N_3998);
and U5869 (N_5869,N_2505,N_2025);
nor U5870 (N_5870,N_3621,N_2100);
xor U5871 (N_5871,N_3218,N_3198);
nand U5872 (N_5872,N_2043,N_2922);
and U5873 (N_5873,N_2666,N_2318);
nand U5874 (N_5874,N_3163,N_3466);
nand U5875 (N_5875,N_2837,N_3461);
nor U5876 (N_5876,N_2554,N_3073);
or U5877 (N_5877,N_2264,N_2949);
and U5878 (N_5878,N_3429,N_2717);
xor U5879 (N_5879,N_2024,N_2783);
nor U5880 (N_5880,N_2809,N_3374);
xnor U5881 (N_5881,N_2320,N_3140);
or U5882 (N_5882,N_2328,N_3807);
nor U5883 (N_5883,N_2349,N_3544);
nor U5884 (N_5884,N_3488,N_2826);
nand U5885 (N_5885,N_2811,N_3198);
nand U5886 (N_5886,N_3577,N_3644);
nor U5887 (N_5887,N_3395,N_2454);
or U5888 (N_5888,N_2322,N_2228);
and U5889 (N_5889,N_3510,N_2660);
and U5890 (N_5890,N_2469,N_3876);
nand U5891 (N_5891,N_3385,N_2299);
xor U5892 (N_5892,N_3103,N_2442);
nor U5893 (N_5893,N_3125,N_3435);
nand U5894 (N_5894,N_3977,N_2912);
nor U5895 (N_5895,N_2304,N_3655);
nor U5896 (N_5896,N_2939,N_3279);
and U5897 (N_5897,N_3470,N_3924);
and U5898 (N_5898,N_3924,N_3812);
nor U5899 (N_5899,N_3956,N_2422);
or U5900 (N_5900,N_2552,N_3046);
and U5901 (N_5901,N_2757,N_2188);
and U5902 (N_5902,N_2511,N_3925);
or U5903 (N_5903,N_2174,N_2062);
nor U5904 (N_5904,N_2535,N_3159);
nor U5905 (N_5905,N_2651,N_3387);
xnor U5906 (N_5906,N_2770,N_2126);
xor U5907 (N_5907,N_2071,N_3298);
nand U5908 (N_5908,N_3938,N_3871);
and U5909 (N_5909,N_2992,N_3779);
or U5910 (N_5910,N_2009,N_3477);
or U5911 (N_5911,N_3519,N_3700);
nor U5912 (N_5912,N_2750,N_3079);
xnor U5913 (N_5913,N_2031,N_2337);
nand U5914 (N_5914,N_2556,N_2276);
xnor U5915 (N_5915,N_2524,N_3950);
nand U5916 (N_5916,N_2169,N_3473);
or U5917 (N_5917,N_2113,N_3877);
or U5918 (N_5918,N_2549,N_3638);
and U5919 (N_5919,N_2409,N_3995);
and U5920 (N_5920,N_2134,N_2002);
xnor U5921 (N_5921,N_2727,N_2656);
nand U5922 (N_5922,N_2419,N_3991);
and U5923 (N_5923,N_3894,N_3437);
nor U5924 (N_5924,N_3033,N_2349);
xor U5925 (N_5925,N_3423,N_2166);
nand U5926 (N_5926,N_2058,N_2026);
and U5927 (N_5927,N_3922,N_2976);
nand U5928 (N_5928,N_3529,N_2438);
nor U5929 (N_5929,N_2189,N_2265);
nand U5930 (N_5930,N_2453,N_2868);
and U5931 (N_5931,N_3514,N_3948);
nand U5932 (N_5932,N_2569,N_2243);
or U5933 (N_5933,N_2718,N_3670);
nand U5934 (N_5934,N_3617,N_2339);
and U5935 (N_5935,N_3835,N_2003);
nand U5936 (N_5936,N_3611,N_3939);
nand U5937 (N_5937,N_3122,N_2282);
or U5938 (N_5938,N_2144,N_2105);
nor U5939 (N_5939,N_3629,N_2794);
and U5940 (N_5940,N_3093,N_2941);
or U5941 (N_5941,N_3334,N_3058);
nand U5942 (N_5942,N_2460,N_3934);
nand U5943 (N_5943,N_2765,N_2455);
nand U5944 (N_5944,N_2178,N_2448);
and U5945 (N_5945,N_2358,N_3778);
xor U5946 (N_5946,N_2675,N_3447);
nor U5947 (N_5947,N_3039,N_2036);
nor U5948 (N_5948,N_3283,N_2465);
xnor U5949 (N_5949,N_2957,N_2588);
or U5950 (N_5950,N_3265,N_3935);
nor U5951 (N_5951,N_2200,N_3557);
xor U5952 (N_5952,N_2750,N_2958);
or U5953 (N_5953,N_2218,N_3458);
nor U5954 (N_5954,N_3697,N_2942);
or U5955 (N_5955,N_3491,N_2388);
xnor U5956 (N_5956,N_3928,N_2249);
and U5957 (N_5957,N_3795,N_3011);
nand U5958 (N_5958,N_2581,N_2959);
or U5959 (N_5959,N_3089,N_2899);
nor U5960 (N_5960,N_2318,N_2504);
and U5961 (N_5961,N_3976,N_3639);
or U5962 (N_5962,N_3472,N_3997);
nor U5963 (N_5963,N_3490,N_2493);
and U5964 (N_5964,N_3908,N_2486);
xnor U5965 (N_5965,N_3593,N_2392);
or U5966 (N_5966,N_2987,N_2386);
nor U5967 (N_5967,N_2987,N_2950);
and U5968 (N_5968,N_2118,N_2933);
and U5969 (N_5969,N_3878,N_2052);
xor U5970 (N_5970,N_3526,N_2897);
xnor U5971 (N_5971,N_3792,N_3772);
nand U5972 (N_5972,N_2970,N_3009);
and U5973 (N_5973,N_2173,N_3306);
nor U5974 (N_5974,N_3749,N_2028);
nor U5975 (N_5975,N_2067,N_3220);
and U5976 (N_5976,N_3667,N_2671);
or U5977 (N_5977,N_3107,N_2320);
nand U5978 (N_5978,N_2904,N_3408);
or U5979 (N_5979,N_2006,N_2532);
xor U5980 (N_5980,N_2258,N_2205);
or U5981 (N_5981,N_3244,N_2404);
nor U5982 (N_5982,N_2596,N_2058);
or U5983 (N_5983,N_3696,N_2990);
and U5984 (N_5984,N_3511,N_3764);
and U5985 (N_5985,N_3907,N_3574);
xnor U5986 (N_5986,N_3974,N_3955);
nor U5987 (N_5987,N_3341,N_2935);
or U5988 (N_5988,N_3078,N_3486);
nor U5989 (N_5989,N_3889,N_3184);
nor U5990 (N_5990,N_2341,N_2311);
nand U5991 (N_5991,N_3663,N_2516);
or U5992 (N_5992,N_2795,N_2719);
or U5993 (N_5993,N_2343,N_2448);
nor U5994 (N_5994,N_3364,N_3005);
and U5995 (N_5995,N_2799,N_2027);
nand U5996 (N_5996,N_2629,N_3740);
and U5997 (N_5997,N_2913,N_2149);
nor U5998 (N_5998,N_3298,N_2296);
nand U5999 (N_5999,N_3562,N_2823);
or U6000 (N_6000,N_4454,N_5366);
xnor U6001 (N_6001,N_4729,N_5965);
and U6002 (N_6002,N_5192,N_5398);
and U6003 (N_6003,N_5811,N_5312);
nand U6004 (N_6004,N_4558,N_5952);
and U6005 (N_6005,N_4936,N_5852);
and U6006 (N_6006,N_5598,N_4335);
nor U6007 (N_6007,N_4392,N_4032);
or U6008 (N_6008,N_4478,N_5246);
nand U6009 (N_6009,N_5898,N_5086);
or U6010 (N_6010,N_4377,N_4612);
or U6011 (N_6011,N_5487,N_5793);
xnor U6012 (N_6012,N_5834,N_4394);
or U6013 (N_6013,N_4425,N_5334);
nor U6014 (N_6014,N_5039,N_4733);
or U6015 (N_6015,N_4198,N_5482);
nand U6016 (N_6016,N_4974,N_5995);
and U6017 (N_6017,N_5112,N_4338);
xnor U6018 (N_6018,N_4809,N_4743);
nand U6019 (N_6019,N_5236,N_4862);
and U6020 (N_6020,N_4934,N_4426);
nand U6021 (N_6021,N_4928,N_4891);
and U6022 (N_6022,N_4054,N_5743);
nor U6023 (N_6023,N_4705,N_5678);
xor U6024 (N_6024,N_5139,N_5842);
xnor U6025 (N_6025,N_4538,N_4004);
nor U6026 (N_6026,N_5194,N_4080);
and U6027 (N_6027,N_5008,N_5163);
nor U6028 (N_6028,N_5990,N_4189);
and U6029 (N_6029,N_4179,N_5734);
nor U6030 (N_6030,N_5886,N_4503);
nor U6031 (N_6031,N_4146,N_4346);
nand U6032 (N_6032,N_5712,N_5972);
nor U6033 (N_6033,N_4710,N_5189);
or U6034 (N_6034,N_5600,N_4439);
or U6035 (N_6035,N_5009,N_4632);
and U6036 (N_6036,N_4501,N_4232);
or U6037 (N_6037,N_5709,N_4925);
or U6038 (N_6038,N_5862,N_4896);
nor U6039 (N_6039,N_4703,N_5564);
and U6040 (N_6040,N_4473,N_5969);
nor U6041 (N_6041,N_4741,N_5090);
nand U6042 (N_6042,N_5403,N_4332);
nor U6043 (N_6043,N_4460,N_5256);
and U6044 (N_6044,N_5031,N_5446);
or U6045 (N_6045,N_5528,N_4025);
nand U6046 (N_6046,N_4985,N_5715);
nor U6047 (N_6047,N_4587,N_5057);
nor U6048 (N_6048,N_4072,N_4724);
and U6049 (N_6049,N_5079,N_5149);
xnor U6050 (N_6050,N_5107,N_5318);
nand U6051 (N_6051,N_4387,N_4872);
xnor U6052 (N_6052,N_5479,N_4702);
nand U6053 (N_6053,N_5354,N_4154);
xnor U6054 (N_6054,N_5705,N_4611);
and U6055 (N_6055,N_4349,N_5053);
and U6056 (N_6056,N_5098,N_4837);
nand U6057 (N_6057,N_4561,N_4308);
xnor U6058 (N_6058,N_5812,N_4591);
and U6059 (N_6059,N_4968,N_5477);
xnor U6060 (N_6060,N_4415,N_5763);
or U6061 (N_6061,N_4412,N_5359);
or U6062 (N_6062,N_4227,N_4513);
nor U6063 (N_6063,N_5064,N_5530);
and U6064 (N_6064,N_4022,N_5668);
nor U6065 (N_6065,N_5494,N_5252);
or U6066 (N_6066,N_4479,N_4131);
and U6067 (N_6067,N_4776,N_5124);
and U6068 (N_6068,N_5063,N_5830);
and U6069 (N_6069,N_4271,N_4637);
nor U6070 (N_6070,N_4706,N_5178);
nor U6071 (N_6071,N_5373,N_5435);
nand U6072 (N_6072,N_5540,N_4720);
nand U6073 (N_6073,N_5013,N_4677);
nor U6074 (N_6074,N_4083,N_5132);
and U6075 (N_6075,N_4371,N_4246);
xnor U6076 (N_6076,N_4633,N_4844);
and U6077 (N_6077,N_4443,N_5597);
xor U6078 (N_6078,N_5674,N_5946);
or U6079 (N_6079,N_4532,N_4196);
nand U6080 (N_6080,N_4954,N_5999);
nor U6081 (N_6081,N_5263,N_4835);
or U6082 (N_6082,N_5421,N_4116);
nor U6083 (N_6083,N_4038,N_4435);
nand U6084 (N_6084,N_5606,N_5358);
nor U6085 (N_6085,N_4977,N_5719);
nand U6086 (N_6086,N_5877,N_5356);
xnor U6087 (N_6087,N_4222,N_4737);
nor U6088 (N_6088,N_4506,N_5510);
nor U6089 (N_6089,N_4284,N_5786);
nor U6090 (N_6090,N_4530,N_5900);
or U6091 (N_6091,N_5024,N_4327);
nor U6092 (N_6092,N_4715,N_4570);
or U6093 (N_6093,N_4178,N_5945);
and U6094 (N_6094,N_4797,N_4773);
nor U6095 (N_6095,N_4522,N_5046);
xor U6096 (N_6096,N_4785,N_4369);
nand U6097 (N_6097,N_4857,N_4641);
or U6098 (N_6098,N_5440,N_4309);
and U6099 (N_6099,N_4302,N_5805);
and U6100 (N_6100,N_5286,N_4268);
nand U6101 (N_6101,N_5828,N_5397);
and U6102 (N_6102,N_4077,N_5655);
and U6103 (N_6103,N_5514,N_4515);
or U6104 (N_6104,N_5537,N_5534);
nor U6105 (N_6105,N_4593,N_5105);
nor U6106 (N_6106,N_4202,N_4736);
or U6107 (N_6107,N_5382,N_5725);
nand U6108 (N_6108,N_5637,N_5238);
or U6109 (N_6109,N_5422,N_5224);
nor U6110 (N_6110,N_4402,N_4172);
nand U6111 (N_6111,N_4897,N_5295);
or U6112 (N_6112,N_4629,N_5723);
nor U6113 (N_6113,N_4341,N_5428);
xor U6114 (N_6114,N_4043,N_5113);
or U6115 (N_6115,N_4304,N_4483);
nand U6116 (N_6116,N_5760,N_5707);
nor U6117 (N_6117,N_4470,N_4673);
or U6118 (N_6118,N_4517,N_4700);
xor U6119 (N_6119,N_4541,N_4467);
xnor U6120 (N_6120,N_4709,N_4104);
nor U6121 (N_6121,N_5146,N_4003);
and U6122 (N_6122,N_5431,N_5169);
or U6123 (N_6123,N_5036,N_5928);
nand U6124 (N_6124,N_4320,N_4253);
nor U6125 (N_6125,N_4375,N_5621);
nand U6126 (N_6126,N_4815,N_5101);
nand U6127 (N_6127,N_4790,N_5802);
or U6128 (N_6128,N_4667,N_5504);
nand U6129 (N_6129,N_4627,N_4543);
nor U6130 (N_6130,N_4829,N_4868);
and U6131 (N_6131,N_5503,N_4642);
nand U6132 (N_6132,N_5659,N_4544);
and U6133 (N_6133,N_4407,N_5823);
or U6134 (N_6134,N_5242,N_4281);
or U6135 (N_6135,N_5203,N_4449);
xor U6136 (N_6136,N_5200,N_4808);
nor U6137 (N_6137,N_5167,N_5496);
and U6138 (N_6138,N_5187,N_4429);
or U6139 (N_6139,N_5774,N_5075);
and U6140 (N_6140,N_5376,N_4566);
or U6141 (N_6141,N_4067,N_4095);
and U6142 (N_6142,N_4586,N_4123);
nor U6143 (N_6143,N_4786,N_4597);
and U6144 (N_6144,N_4051,N_5015);
or U6145 (N_6145,N_5243,N_5517);
nand U6146 (N_6146,N_4832,N_5237);
and U6147 (N_6147,N_5863,N_5777);
nor U6148 (N_6148,N_5211,N_5249);
nand U6149 (N_6149,N_5392,N_5826);
xnor U6150 (N_6150,N_5924,N_4907);
nand U6151 (N_6151,N_5304,N_4241);
nor U6152 (N_6152,N_4875,N_4171);
nand U6153 (N_6153,N_5415,N_5151);
and U6154 (N_6154,N_4912,N_5557);
nand U6155 (N_6155,N_5752,N_4313);
or U6156 (N_6156,N_5662,N_4895);
xor U6157 (N_6157,N_5984,N_4030);
nand U6158 (N_6158,N_5115,N_5604);
and U6159 (N_6159,N_4184,N_4688);
or U6160 (N_6160,N_5770,N_5335);
nand U6161 (N_6161,N_5615,N_4552);
nand U6162 (N_6162,N_4845,N_4037);
or U6163 (N_6163,N_4055,N_5664);
and U6164 (N_6164,N_5745,N_5677);
and U6165 (N_6165,N_4640,N_4619);
and U6166 (N_6166,N_5569,N_4040);
xor U6167 (N_6167,N_4704,N_4932);
or U6168 (N_6168,N_5257,N_5483);
and U6169 (N_6169,N_4231,N_5448);
and U6170 (N_6170,N_4236,N_5488);
or U6171 (N_6171,N_4063,N_5396);
and U6172 (N_6172,N_5375,N_5410);
xnor U6173 (N_6173,N_5082,N_4383);
or U6174 (N_6174,N_4555,N_5672);
nand U6175 (N_6175,N_5337,N_4824);
and U6176 (N_6176,N_4796,N_4034);
nor U6177 (N_6177,N_4858,N_5866);
nor U6178 (N_6178,N_4628,N_5749);
xor U6179 (N_6179,N_5642,N_5887);
xnor U6180 (N_6180,N_4575,N_5260);
nor U6181 (N_6181,N_5726,N_5616);
and U6182 (N_6182,N_4781,N_5118);
nor U6183 (N_6183,N_4577,N_5294);
xnor U6184 (N_6184,N_5706,N_4249);
nand U6185 (N_6185,N_4605,N_4683);
nand U6186 (N_6186,N_4492,N_5908);
nor U6187 (N_6187,N_4477,N_5650);
nand U6188 (N_6188,N_5176,N_5547);
or U6189 (N_6189,N_4609,N_5476);
nand U6190 (N_6190,N_4825,N_5500);
and U6191 (N_6191,N_5533,N_4442);
and U6192 (N_6192,N_4898,N_4693);
nor U6193 (N_6193,N_4744,N_5188);
nor U6194 (N_6194,N_5948,N_5038);
xnor U6195 (N_6195,N_4242,N_4753);
xnor U6196 (N_6196,N_5136,N_4028);
or U6197 (N_6197,N_5847,N_5379);
nand U6198 (N_6198,N_4441,N_5981);
or U6199 (N_6199,N_4254,N_5808);
or U6200 (N_6200,N_5137,N_5562);
and U6201 (N_6201,N_5751,N_5348);
nor U6202 (N_6202,N_5175,N_5241);
nor U6203 (N_6203,N_5543,N_5929);
or U6204 (N_6204,N_4511,N_4995);
nand U6205 (N_6205,N_5980,N_4959);
and U6206 (N_6206,N_5201,N_4110);
and U6207 (N_6207,N_5754,N_4029);
or U6208 (N_6208,N_5833,N_5579);
nand U6209 (N_6209,N_4811,N_4618);
or U6210 (N_6210,N_4657,N_5322);
xnor U6211 (N_6211,N_5688,N_5895);
xnor U6212 (N_6212,N_5025,N_5787);
xor U6213 (N_6213,N_5587,N_5512);
or U6214 (N_6214,N_4884,N_4939);
nor U6215 (N_6215,N_4488,N_4944);
nand U6216 (N_6216,N_5507,N_4128);
nor U6217 (N_6217,N_5560,N_5595);
or U6218 (N_6218,N_4554,N_4278);
xnor U6219 (N_6219,N_5344,N_4718);
xnor U6220 (N_6220,N_5888,N_5452);
or U6221 (N_6221,N_5791,N_5645);
nand U6222 (N_6222,N_4748,N_4187);
and U6223 (N_6223,N_5350,N_4036);
nand U6224 (N_6224,N_4257,N_5738);
or U6225 (N_6225,N_4181,N_4355);
or U6226 (N_6226,N_4229,N_4307);
or U6227 (N_6227,N_4975,N_5832);
nand U6228 (N_6228,N_5371,N_4011);
and U6229 (N_6229,N_4388,N_5795);
and U6230 (N_6230,N_4420,N_4638);
or U6231 (N_6231,N_4448,N_5316);
nand U6232 (N_6232,N_5071,N_4059);
or U6233 (N_6233,N_4379,N_4604);
xnor U6234 (N_6234,N_4082,N_4913);
xor U6235 (N_6235,N_5610,N_4955);
and U6236 (N_6236,N_5471,N_5352);
and U6237 (N_6237,N_5739,N_5592);
nand U6238 (N_6238,N_4363,N_4670);
or U6239 (N_6239,N_5120,N_5590);
or U6240 (N_6240,N_4337,N_5234);
xor U6241 (N_6241,N_5131,N_5612);
or U6242 (N_6242,N_5906,N_4989);
xnor U6243 (N_6243,N_4947,N_4972);
nor U6244 (N_6244,N_4672,N_5128);
and U6245 (N_6245,N_4070,N_5640);
or U6246 (N_6246,N_5198,N_5497);
xnor U6247 (N_6247,N_4935,N_5976);
nor U6248 (N_6248,N_5170,N_4675);
nand U6249 (N_6249,N_5639,N_5456);
and U6250 (N_6250,N_4205,N_5349);
xnor U6251 (N_6251,N_4789,N_4182);
nor U6252 (N_6252,N_4386,N_5424);
or U6253 (N_6253,N_4911,N_4133);
or U6254 (N_6254,N_5012,N_5219);
or U6255 (N_6255,N_4471,N_4784);
or U6256 (N_6256,N_4060,N_4457);
xnor U6257 (N_6257,N_4926,N_4965);
xnor U6258 (N_6258,N_4049,N_5164);
nor U6259 (N_6259,N_5384,N_4047);
or U6260 (N_6260,N_4991,N_5433);
or U6261 (N_6261,N_5463,N_4264);
or U6262 (N_6262,N_5230,N_4652);
or U6263 (N_6263,N_4462,N_5575);
xnor U6264 (N_6264,N_5561,N_4887);
xor U6265 (N_6265,N_4553,N_5572);
or U6266 (N_6266,N_4804,N_5254);
or U6267 (N_6267,N_4582,N_4261);
nand U6268 (N_6268,N_4957,N_5902);
or U6269 (N_6269,N_4542,N_4916);
and U6270 (N_6270,N_4722,N_5274);
and U6271 (N_6271,N_4144,N_4207);
nand U6272 (N_6272,N_4745,N_5147);
nand U6273 (N_6273,N_4446,N_4382);
nand U6274 (N_6274,N_4026,N_5427);
and U6275 (N_6275,N_4438,N_5625);
nand U6276 (N_6276,N_4486,N_5521);
and U6277 (N_6277,N_4653,N_4016);
nand U6278 (N_6278,N_5554,N_5698);
xor U6279 (N_6279,N_4805,N_5017);
xnor U6280 (N_6280,N_5780,N_4318);
nor U6281 (N_6281,N_4914,N_5810);
nand U6282 (N_6282,N_4342,N_4017);
or U6283 (N_6283,N_4311,N_5045);
and U6284 (N_6284,N_5080,N_5627);
xor U6285 (N_6285,N_5016,N_5042);
nand U6286 (N_6286,N_4573,N_4291);
and U6287 (N_6287,N_5258,N_5034);
and U6288 (N_6288,N_4062,N_5481);
nand U6289 (N_6289,N_5532,N_4772);
or U6290 (N_6290,N_4057,N_4788);
nand U6291 (N_6291,N_5551,N_5935);
xor U6292 (N_6292,N_4258,N_4920);
and U6293 (N_6293,N_5685,N_5617);
or U6294 (N_6294,N_4045,N_4357);
xor U6295 (N_6295,N_4714,N_4177);
xnor U6296 (N_6296,N_4169,N_5958);
and U6297 (N_6297,N_4157,N_4536);
xnor U6298 (N_6298,N_5264,N_4565);
nand U6299 (N_6299,N_5553,N_4643);
and U6300 (N_6300,N_5309,N_5838);
or U6301 (N_6301,N_4340,N_4364);
nand U6302 (N_6302,N_5943,N_5275);
nor U6303 (N_6303,N_4952,N_4817);
nand U6304 (N_6304,N_4399,N_5516);
xnor U6305 (N_6305,N_4801,N_4275);
or U6306 (N_6306,N_4014,N_5216);
nor U6307 (N_6307,N_5412,N_4819);
nor U6308 (N_6308,N_5693,N_4136);
and U6309 (N_6309,N_4750,N_5361);
nand U6310 (N_6310,N_4416,N_4370);
or U6311 (N_6311,N_4663,N_5858);
nand U6312 (N_6312,N_4865,N_4594);
nor U6313 (N_6313,N_5851,N_4738);
and U6314 (N_6314,N_4099,N_5378);
nor U6315 (N_6315,N_4964,N_4233);
or U6316 (N_6316,N_5423,N_4391);
nand U6317 (N_6317,N_4874,N_5629);
nand U6318 (N_6318,N_4607,N_4716);
xor U6319 (N_6319,N_5023,N_4153);
xnor U6320 (N_6320,N_5287,N_4976);
nor U6321 (N_6321,N_5781,N_4101);
xor U6322 (N_6322,N_5975,N_5055);
and U6323 (N_6323,N_5973,N_4319);
xnor U6324 (N_6324,N_5388,N_5209);
nor U6325 (N_6325,N_5957,N_4005);
nor U6326 (N_6326,N_5936,N_5262);
nor U6327 (N_6327,N_5141,N_5297);
and U6328 (N_6328,N_5393,N_5933);
and U6329 (N_6329,N_5631,N_4678);
and U6330 (N_6330,N_5321,N_5223);
xor U6331 (N_6331,N_4185,N_4092);
nor U6332 (N_6332,N_5964,N_4331);
or U6333 (N_6333,N_4218,N_5729);
nand U6334 (N_6334,N_4816,N_4859);
nand U6335 (N_6335,N_5670,N_4197);
and U6336 (N_6336,N_4373,N_4800);
xor U6337 (N_6337,N_5145,N_5613);
nor U6338 (N_6338,N_5315,N_5408);
nor U6339 (N_6339,N_5317,N_5492);
xor U6340 (N_6340,N_5044,N_4353);
and U6341 (N_6341,N_5360,N_4734);
or U6342 (N_6342,N_5550,N_4405);
xnor U6343 (N_6343,N_5699,N_5444);
or U6344 (N_6344,N_5102,N_5985);
or U6345 (N_6345,N_5827,N_5728);
or U6346 (N_6346,N_4746,N_5066);
or U6347 (N_6347,N_5695,N_5380);
xnor U6348 (N_6348,N_5511,N_4108);
nor U6349 (N_6349,N_4882,N_5485);
or U6350 (N_6350,N_5003,N_5893);
nand U6351 (N_6351,N_5915,N_5058);
and U6352 (N_6352,N_4041,N_5202);
and U6353 (N_6353,N_5218,N_5602);
xnor U6354 (N_6354,N_5342,N_4210);
or U6355 (N_6355,N_5156,N_4495);
or U6356 (N_6356,N_4119,N_4073);
nand U6357 (N_6357,N_4287,N_4458);
xor U6358 (N_6358,N_5555,N_5314);
xnor U6359 (N_6359,N_5383,N_5675);
nor U6360 (N_6360,N_4498,N_4430);
xor U6361 (N_6361,N_4105,N_5097);
nor U6362 (N_6362,N_4909,N_5091);
xnor U6363 (N_6363,N_4680,N_4176);
xnor U6364 (N_6364,N_4444,N_4701);
nand U6365 (N_6365,N_5095,N_5667);
xnor U6366 (N_6366,N_4214,N_4322);
and U6367 (N_6367,N_5030,N_4065);
xnor U6368 (N_6368,N_5129,N_4103);
and U6369 (N_6369,N_5620,N_4963);
nor U6370 (N_6370,N_4946,N_5776);
or U6371 (N_6371,N_4306,N_4856);
nand U6372 (N_6372,N_4751,N_5527);
nor U6373 (N_6373,N_5692,N_4598);
nand U6374 (N_6374,N_5596,N_5020);
nand U6375 (N_6375,N_5248,N_4818);
xnor U6376 (N_6376,N_4514,N_4024);
and U6377 (N_6377,N_5462,N_4567);
nand U6378 (N_6378,N_5026,N_5829);
xor U6379 (N_6379,N_5879,N_4767);
nand U6380 (N_6380,N_5855,N_4739);
xnor U6381 (N_6381,N_4234,N_4219);
and U6382 (N_6382,N_5636,N_5859);
and U6383 (N_6383,N_4685,N_5501);
or U6384 (N_6384,N_4948,N_4943);
xnor U6385 (N_6385,N_5819,N_5506);
or U6386 (N_6386,N_5735,N_4831);
xnor U6387 (N_6387,N_5472,N_5979);
or U6388 (N_6388,N_4109,N_4938);
xor U6389 (N_6389,N_5313,N_4668);
and U6390 (N_6390,N_4404,N_5632);
or U6391 (N_6391,N_5329,N_4145);
nor U6392 (N_6392,N_5565,N_5755);
nand U6393 (N_6393,N_5907,N_4549);
xnor U6394 (N_6394,N_4206,N_4669);
xor U6395 (N_6395,N_5062,N_4691);
nor U6396 (N_6396,N_5708,N_5296);
xor U6397 (N_6397,N_5890,N_5803);
nand U6398 (N_6398,N_5000,N_4838);
nor U6399 (N_6399,N_4863,N_4048);
nand U6400 (N_6400,N_4758,N_5765);
nor U6401 (N_6401,N_5566,N_5308);
and U6402 (N_6402,N_4775,N_5404);
and U6403 (N_6403,N_5429,N_4725);
nand U6404 (N_6404,N_5442,N_5988);
and U6405 (N_6405,N_5470,N_5591);
and U6406 (N_6406,N_5614,N_4765);
or U6407 (N_6407,N_4730,N_5368);
and U6408 (N_6408,N_5056,N_5578);
nor U6409 (N_6409,N_5402,N_4682);
nand U6410 (N_6410,N_4323,N_5021);
and U6411 (N_6411,N_5697,N_5007);
xnor U6412 (N_6412,N_4754,N_5439);
nand U6413 (N_6413,N_5239,N_4259);
xor U6414 (N_6414,N_5901,N_4671);
nor U6415 (N_6415,N_5956,N_4707);
or U6416 (N_6416,N_5126,N_4616);
xnor U6417 (N_6417,N_4220,N_5372);
or U6418 (N_6418,N_5520,N_4174);
and U6419 (N_6419,N_5524,N_5857);
xor U6420 (N_6420,N_4225,N_5663);
nor U6421 (N_6421,N_5110,N_5716);
or U6422 (N_6422,N_5815,N_4097);
and U6423 (N_6423,N_4719,N_5119);
nor U6424 (N_6424,N_4200,N_5836);
nand U6425 (N_6425,N_4098,N_4830);
xnor U6426 (N_6426,N_5934,N_4413);
and U6427 (N_6427,N_5338,N_5660);
nor U6428 (N_6428,N_5212,N_5292);
xnor U6429 (N_6429,N_5469,N_5332);
and U6430 (N_6430,N_4440,N_5228);
nor U6431 (N_6431,N_5266,N_4883);
xnor U6432 (N_6432,N_5401,N_4505);
xor U6433 (N_6433,N_4596,N_5775);
nand U6434 (N_6434,N_4251,N_4276);
or U6435 (N_6435,N_5405,N_5331);
xnor U6436 (N_6436,N_5801,N_4828);
xor U6437 (N_6437,N_5109,N_5001);
or U6438 (N_6438,N_4960,N_5099);
nor U6439 (N_6439,N_5267,N_5505);
nand U6440 (N_6440,N_5094,N_5654);
or U6441 (N_6441,N_4623,N_4686);
nand U6442 (N_6442,N_5150,N_5624);
or U6443 (N_6443,N_5293,N_4903);
xor U6444 (N_6444,N_4581,N_5991);
nand U6445 (N_6445,N_5027,N_5122);
xnor U6446 (N_6446,N_5290,N_5796);
and U6447 (N_6447,N_5778,N_4314);
and U6448 (N_6448,N_5861,N_4094);
and U6449 (N_6449,N_4622,N_4813);
or U6450 (N_6450,N_4493,N_5679);
or U6451 (N_6451,N_4138,N_4713);
or U6452 (N_6452,N_4864,N_5319);
nand U6453 (N_6453,N_4915,N_5896);
nand U6454 (N_6454,N_4899,N_5588);
xor U6455 (N_6455,N_5619,N_4615);
nor U6456 (N_6456,N_5545,N_4380);
and U6457 (N_6457,N_4129,N_5445);
nor U6458 (N_6458,N_4820,N_4367);
nor U6459 (N_6459,N_5199,N_5974);
and U6460 (N_6460,N_5400,N_5634);
or U6461 (N_6461,N_4980,N_5193);
or U6462 (N_6462,N_5018,N_4881);
and U6463 (N_6463,N_5894,N_4273);
nand U6464 (N_6464,N_4656,N_5409);
or U6465 (N_6465,N_5741,N_5953);
nand U6466 (N_6466,N_4058,N_4588);
and U6467 (N_6467,N_4624,N_5369);
nand U6468 (N_6468,N_4199,N_4317);
nand U6469 (N_6469,N_5285,N_4132);
nor U6470 (N_6470,N_4600,N_4866);
and U6471 (N_6471,N_5871,N_4676);
nand U6472 (N_6472,N_5468,N_5473);
and U6473 (N_6473,N_5737,N_4984);
xnor U6474 (N_6474,N_5635,N_5869);
xnor U6475 (N_6475,N_4312,N_5100);
xor U6476 (N_6476,N_5977,N_5447);
nor U6477 (N_6477,N_4390,N_4137);
nor U6478 (N_6478,N_4244,N_5970);
or U6479 (N_6479,N_4951,N_5047);
nand U6480 (N_6480,N_4139,N_5594);
nand U6481 (N_6481,N_4918,N_4124);
nor U6482 (N_6482,N_5181,N_4747);
and U6483 (N_6483,N_5824,N_5073);
nand U6484 (N_6484,N_4988,N_5548);
nor U6485 (N_6485,N_5186,N_4580);
xnor U6486 (N_6486,N_5077,N_5443);
or U6487 (N_6487,N_4472,N_5166);
nand U6488 (N_6488,N_5891,N_5922);
nor U6489 (N_6489,N_5766,N_4533);
or U6490 (N_6490,N_4793,N_5700);
and U6491 (N_6491,N_5814,N_5794);
nand U6492 (N_6492,N_5464,N_5395);
or U6493 (N_6493,N_5998,N_5134);
nor U6494 (N_6494,N_5800,N_5905);
nor U6495 (N_6495,N_4823,N_4890);
and U6496 (N_6496,N_4112,N_4089);
nand U6497 (N_6497,N_5067,N_4634);
xor U6498 (N_6498,N_4090,N_5363);
nor U6499 (N_6499,N_5959,N_5982);
or U6500 (N_6500,N_4557,N_4625);
nand U6501 (N_6501,N_4539,N_5454);
xor U6502 (N_6502,N_4931,N_5840);
and U6503 (N_6503,N_4086,N_4126);
nand U6504 (N_6504,N_5740,N_5875);
and U6505 (N_6505,N_4827,N_5160);
xnor U6506 (N_6506,N_5919,N_5955);
nor U6507 (N_6507,N_5327,N_4559);
nand U6508 (N_6508,N_5050,N_4173);
or U6509 (N_6509,N_4135,N_5867);
nor U6510 (N_6510,N_5813,N_4791);
xor U6511 (N_6511,N_4464,N_4595);
nand U6512 (N_6512,N_4161,N_5070);
and U6513 (N_6513,N_4418,N_4344);
nand U6514 (N_6514,N_5381,N_5195);
xor U6515 (N_6515,N_4433,N_5426);
xor U6516 (N_6516,N_5607,N_4252);
nand U6517 (N_6517,N_5168,N_4910);
nand U6518 (N_6518,N_5960,N_4164);
xor U6519 (N_6519,N_5820,N_5284);
nor U6520 (N_6520,N_4902,N_5605);
nor U6521 (N_6521,N_4849,N_5484);
or U6522 (N_6522,N_4620,N_4900);
nand U6523 (N_6523,N_4263,N_4434);
nor U6524 (N_6524,N_4639,N_5940);
nand U6525 (N_6525,N_4238,N_5278);
xor U6526 (N_6526,N_5060,N_5346);
or U6527 (N_6527,N_4469,N_5005);
or U6528 (N_6528,N_5916,N_5457);
xnor U6529 (N_6529,N_4742,N_5526);
or U6530 (N_6530,N_4294,N_4873);
xor U6531 (N_6531,N_4877,N_4520);
nand U6532 (N_6532,N_4217,N_5885);
nor U6533 (N_6533,N_5718,N_5172);
nand U6534 (N_6534,N_4922,N_4451);
nor U6535 (N_6535,N_5116,N_4661);
xor U6536 (N_6536,N_4997,N_4497);
xor U6537 (N_6537,N_5340,N_4301);
nand U6538 (N_6538,N_5938,N_5085);
nor U6539 (N_6539,N_5954,N_5385);
and U6540 (N_6540,N_4613,N_5696);
xnor U6541 (N_6541,N_5153,N_5283);
nor U6542 (N_6542,N_4230,N_5250);
or U6543 (N_6543,N_4050,N_4771);
xnor U6544 (N_6544,N_4726,N_5966);
or U6545 (N_6545,N_4476,N_4962);
or U6546 (N_6546,N_4860,N_5950);
xnor U6547 (N_6547,N_5849,N_5434);
nor U6548 (N_6548,N_4606,N_4708);
and U6549 (N_6549,N_4141,N_5121);
or U6550 (N_6550,N_5920,N_4876);
and U6551 (N_6551,N_4941,N_4846);
and U6552 (N_6552,N_4583,N_4140);
nand U6553 (N_6553,N_4982,N_5618);
nor U6554 (N_6554,N_4998,N_4794);
xnor U6555 (N_6555,N_4983,N_4147);
xor U6556 (N_6556,N_4212,N_4889);
xor U6557 (N_6557,N_5846,N_4159);
nand U6558 (N_6558,N_4428,N_4534);
and U6559 (N_6559,N_5983,N_5762);
nand U6560 (N_6560,N_5686,N_4782);
xnor U6561 (N_6561,N_5208,N_4562);
or U6562 (N_6562,N_4840,N_5182);
and U6563 (N_6563,N_4735,N_5702);
and U6564 (N_6564,N_4762,N_4381);
xor U6565 (N_6565,N_4345,N_4537);
nor U6566 (N_6566,N_5747,N_4152);
and U6567 (N_6567,N_5878,N_4069);
and U6568 (N_6568,N_4423,N_4798);
and U6569 (N_6569,N_4042,N_4118);
or U6570 (N_6570,N_5022,N_5272);
xnor U6571 (N_6571,N_5529,N_5736);
xor U6572 (N_6572,N_5436,N_4906);
xor U6573 (N_6573,N_5364,N_5152);
xnor U6574 (N_6574,N_5748,N_4006);
nand U6575 (N_6575,N_4752,N_4578);
nand U6576 (N_6576,N_4971,N_5582);
and U6577 (N_6577,N_4525,N_4717);
nand U6578 (N_6578,N_5074,N_5549);
nand U6579 (N_6579,N_5214,N_5558);
nand U6580 (N_6580,N_5563,N_4500);
xor U6581 (N_6581,N_4494,N_4919);
or U6582 (N_6582,N_4852,N_4463);
nor U6583 (N_6583,N_5903,N_5713);
nor U6584 (N_6584,N_5779,N_5104);
or U6585 (N_6585,N_5515,N_4066);
and U6586 (N_6586,N_5519,N_4556);
nand U6587 (N_6587,N_4614,N_5028);
or U6588 (N_6588,N_4635,N_4410);
nand U6589 (N_6589,N_5420,N_5430);
or U6590 (N_6590,N_5307,N_5522);
xnor U6591 (N_6591,N_4285,N_4270);
nand U6592 (N_6592,N_5365,N_5559);
nor U6593 (N_6593,N_5673,N_5498);
xnor U6594 (N_6594,N_4348,N_4465);
xnor U6595 (N_6595,N_4969,N_5114);
nand U6596 (N_6596,N_4821,N_4459);
and U6597 (N_6597,N_5014,N_4325);
nor U6598 (N_6598,N_5437,N_4455);
nand U6599 (N_6599,N_4774,N_5854);
xnor U6600 (N_6600,N_4994,N_5389);
nand U6601 (N_6601,N_4321,N_5949);
nand U6602 (N_6602,N_4216,N_5065);
nand U6603 (N_6603,N_5689,N_5490);
xor U6604 (N_6604,N_5608,N_4945);
and U6605 (N_6605,N_4551,N_4940);
and U6606 (N_6606,N_5930,N_4973);
xnor U6607 (N_6607,N_4855,N_4528);
nor U6608 (N_6608,N_5320,N_5889);
xor U6609 (N_6609,N_5465,N_4194);
xor U6610 (N_6610,N_4223,N_4265);
xor U6611 (N_6611,N_5499,N_5721);
and U6612 (N_6612,N_4008,N_4953);
and U6613 (N_6613,N_5874,N_5377);
or U6614 (N_6614,N_5799,N_4088);
and U6615 (N_6615,N_4190,N_5767);
nand U6616 (N_6616,N_4279,N_5544);
nand U6617 (N_6617,N_4681,N_4079);
nand U6618 (N_6618,N_4806,N_5213);
or U6619 (N_6619,N_5730,N_4814);
or U6620 (N_6620,N_4074,N_5932);
nor U6621 (N_6621,N_4524,N_5759);
nand U6622 (N_6622,N_5733,N_5926);
and U6623 (N_6623,N_5425,N_5651);
nor U6624 (N_6624,N_4599,N_5914);
nor U6625 (N_6625,N_4843,N_5536);
xor U6626 (N_6626,N_5148,N_5925);
nor U6627 (N_6627,N_5041,N_4240);
and U6628 (N_6628,N_4778,N_4908);
and U6629 (N_6629,N_5518,N_5652);
nand U6630 (N_6630,N_5704,N_5390);
nor U6631 (N_6631,N_4892,N_5265);
xor U6632 (N_6632,N_4419,N_4487);
xnor U6633 (N_6633,N_4842,N_5996);
xor U6634 (N_6634,N_4761,N_4456);
nor U6635 (N_6635,N_4650,N_4879);
or U6636 (N_6636,N_4356,N_4366);
nand U6637 (N_6637,N_5235,N_4396);
nand U6638 (N_6638,N_4102,N_5051);
nand U6639 (N_6639,N_4621,N_4007);
nor U6640 (N_6640,N_4160,N_4516);
nor U6641 (N_6641,N_4274,N_5449);
nor U6642 (N_6642,N_5269,N_4267);
nand U6643 (N_6643,N_5601,N_4096);
nor U6644 (N_6644,N_4894,N_5860);
xnor U6645 (N_6645,N_4519,N_4266);
nor U6646 (N_6646,N_4917,N_4329);
or U6647 (N_6647,N_5648,N_5788);
or U6648 (N_6648,N_4592,N_5671);
and U6649 (N_6649,N_4880,N_4987);
and U6650 (N_6650,N_5495,N_5180);
or U6651 (N_6651,N_4711,N_4010);
or U6652 (N_6652,N_5912,N_5159);
nand U6653 (N_6653,N_5993,N_4489);
or U6654 (N_6654,N_5764,N_5399);
nor U6655 (N_6655,N_4330,N_5864);
nand U6656 (N_6656,N_5475,N_4411);
and U6657 (N_6657,N_4461,N_4192);
nand U6658 (N_6658,N_5251,N_4361);
nand U6659 (N_6659,N_5576,N_4777);
xor U6660 (N_6660,N_4927,N_5245);
xor U6661 (N_6661,N_4540,N_5087);
nand U6662 (N_6662,N_4631,N_5144);
and U6663 (N_6663,N_4076,N_4490);
or U6664 (N_6664,N_5626,N_4601);
xnor U6665 (N_6665,N_5059,N_4510);
or U6666 (N_6666,N_5474,N_4107);
xnor U6667 (N_6667,N_5822,N_4044);
xor U6668 (N_6668,N_5299,N_5407);
nor U6669 (N_6669,N_5261,N_5328);
xnor U6670 (N_6670,N_5868,N_4723);
nor U6671 (N_6671,N_5220,N_4203);
nand U6672 (N_6672,N_5731,N_5963);
xnor U6673 (N_6673,N_4647,N_4068);
nor U6674 (N_6674,N_4763,N_5391);
nor U6675 (N_6675,N_4052,N_5883);
nor U6676 (N_6676,N_4589,N_4526);
or U6677 (N_6677,N_5782,N_4697);
nor U6678 (N_6678,N_4603,N_5552);
and U6679 (N_6679,N_4966,N_5088);
and U6680 (N_6680,N_5931,N_5450);
and U6681 (N_6681,N_5305,N_5962);
or U6682 (N_6682,N_4289,N_4888);
or U6683 (N_6683,N_5909,N_4151);
nand U6684 (N_6684,N_5690,N_4602);
or U6685 (N_6685,N_4269,N_4847);
and U6686 (N_6686,N_5177,N_5277);
nand U6687 (N_6687,N_4305,N_4694);
or U6688 (N_6688,N_4296,N_4204);
or U6689 (N_6689,N_4300,N_4056);
xnor U6690 (N_6690,N_4630,N_5158);
and U6691 (N_6691,N_5538,N_4360);
nand U6692 (N_6692,N_5418,N_5142);
nor U6693 (N_6693,N_4649,N_4208);
nor U6694 (N_6694,N_4687,N_5806);
or U6695 (N_6695,N_5880,N_5019);
or U6696 (N_6696,N_4158,N_4665);
or U6697 (N_6697,N_5881,N_4728);
and U6698 (N_6698,N_5703,N_5951);
xor U6699 (N_6699,N_5165,N_4277);
or U6700 (N_6700,N_5117,N_4993);
or U6701 (N_6701,N_4822,N_4155);
and U6702 (N_6702,N_5040,N_5054);
xor U6703 (N_6703,N_5746,N_4414);
nor U6704 (N_6704,N_4871,N_5502);
or U6705 (N_6705,N_4585,N_4924);
or U6706 (N_6706,N_5783,N_4749);
or U6707 (N_6707,N_4482,N_5509);
xor U6708 (N_6708,N_4431,N_4523);
xor U6709 (N_6709,N_4013,N_5229);
nand U6710 (N_6710,N_4799,N_4262);
xnor U6711 (N_6711,N_4836,N_4766);
xor U6712 (N_6712,N_5108,N_4002);
and U6713 (N_6713,N_5669,N_4923);
or U6714 (N_6714,N_5831,N_5438);
or U6715 (N_6715,N_4134,N_5413);
nor U6716 (N_6716,N_5419,N_5665);
or U6717 (N_6717,N_5493,N_5843);
xnor U6718 (N_6718,N_4803,N_4576);
and U6719 (N_6719,N_4970,N_4015);
nor U6720 (N_6720,N_4046,N_5761);
xnor U6721 (N_6721,N_4802,N_5682);
or U6722 (N_6722,N_4780,N_5081);
nand U6723 (N_6723,N_4247,N_4215);
and U6724 (N_6724,N_4850,N_4904);
xnor U6725 (N_6725,N_4250,N_5326);
nand U6726 (N_6726,N_5244,N_4408);
xnor U6727 (N_6727,N_5732,N_4445);
and U6728 (N_6728,N_5939,N_4020);
and U6729 (N_6729,N_4759,N_4180);
nand U6730 (N_6730,N_4610,N_4290);
and U6731 (N_6731,N_4757,N_4125);
and U6732 (N_6732,N_4689,N_4664);
and U6733 (N_6733,N_5918,N_5480);
or U6734 (N_6734,N_5310,N_4091);
nand U6735 (N_6735,N_5638,N_4093);
and U6736 (N_6736,N_5571,N_5630);
xor U6737 (N_6737,N_4376,N_4853);
nor U6738 (N_6738,N_4260,N_4674);
nand U6739 (N_6739,N_4861,N_5714);
nor U6740 (N_6740,N_5394,N_4372);
nand U6741 (N_6741,N_4481,N_4690);
or U6742 (N_6742,N_4343,N_4779);
nor U6743 (N_6743,N_4833,N_5458);
or U6744 (N_6744,N_4023,N_4378);
or U6745 (N_6745,N_5270,N_4352);
or U6746 (N_6746,N_5839,N_4755);
and U6747 (N_6747,N_4409,N_4395);
nand U6748 (N_6748,N_5367,N_4039);
xnor U6749 (N_6749,N_5844,N_5546);
nand U6750 (N_6750,N_5856,N_5416);
xor U6751 (N_6751,N_4732,N_4298);
nor U6752 (N_6752,N_4870,N_4545);
or U6753 (N_6753,N_4081,N_5593);
and U6754 (N_6754,N_5004,N_5221);
or U6755 (N_6755,N_5302,N_4397);
xnor U6756 (N_6756,N_4756,N_4351);
and U6757 (N_6757,N_4485,N_5910);
and U6758 (N_6758,N_4167,N_4475);
nand U6759 (N_6759,N_4213,N_5432);
xnor U6760 (N_6760,N_5301,N_5649);
and U6761 (N_6761,N_4400,N_5253);
nand U6762 (N_6762,N_5123,N_4393);
nor U6763 (N_6763,N_5899,N_5486);
xnor U6764 (N_6764,N_5268,N_5154);
nand U6765 (N_6765,N_5644,N_5798);
and U6766 (N_6766,N_4087,N_5577);
and U6767 (N_6767,N_5489,N_4012);
and U6768 (N_6768,N_5386,N_4644);
or U6769 (N_6769,N_5303,N_4949);
nor U6770 (N_6770,N_4033,N_5282);
xor U6771 (N_6771,N_5330,N_5653);
nor U6772 (N_6772,N_5837,N_4368);
or U6773 (N_6773,N_4175,N_4546);
and U6774 (N_6774,N_4841,N_4502);
or U6775 (N_6775,N_4084,N_4114);
nor U6776 (N_6776,N_4111,N_4662);
xor U6777 (N_6777,N_5556,N_4358);
nor U6778 (N_6778,N_5841,N_5773);
or U6779 (N_6779,N_5850,N_4333);
and U6780 (N_6780,N_5942,N_5542);
xor U6781 (N_6781,N_5870,N_5720);
nor U6782 (N_6782,N_5341,N_5647);
xor U6783 (N_6783,N_5130,N_5240);
and U6784 (N_6784,N_5259,N_4768);
and U6785 (N_6785,N_5280,N_5010);
nor U6786 (N_6786,N_4531,N_4942);
xnor U6787 (N_6787,N_5076,N_5414);
and U6788 (N_6788,N_5096,N_4981);
nand U6789 (N_6789,N_5758,N_5611);
or U6790 (N_6790,N_4221,N_5661);
nand U6791 (N_6791,N_4001,N_4149);
and U6792 (N_6792,N_5093,N_5911);
or U6793 (N_6793,N_5111,N_5825);
xnor U6794 (N_6794,N_4326,N_5797);
xor U6795 (N_6795,N_4468,N_5622);
nand U6796 (N_6796,N_5994,N_4075);
nand U6797 (N_6797,N_4245,N_5523);
or U6798 (N_6798,N_5944,N_4295);
nor U6799 (N_6799,N_4535,N_4064);
or U6800 (N_6800,N_4646,N_4826);
nand U6801 (N_6801,N_5513,N_5247);
or U6802 (N_6802,N_4403,N_4142);
xnor U6803 (N_6803,N_4851,N_5184);
xnor U6804 (N_6804,N_5897,N_4496);
nand U6805 (N_6805,N_4201,N_5052);
nand U6806 (N_6806,N_5584,N_4315);
nand U6807 (N_6807,N_4256,N_4990);
and U6808 (N_6808,N_5711,N_4893);
and U6809 (N_6809,N_5006,N_4191);
xor U6810 (N_6810,N_5033,N_5531);
nor U6811 (N_6811,N_5185,N_5232);
nor U6812 (N_6812,N_4795,N_4297);
or U6813 (N_6813,N_4336,N_4193);
xnor U6814 (N_6814,N_4491,N_5061);
nand U6815 (N_6815,N_5771,N_5845);
xor U6816 (N_6816,N_5807,N_5573);
or U6817 (N_6817,N_5710,N_4760);
nor U6818 (N_6818,N_4529,N_4527);
or U6819 (N_6819,N_5683,N_4617);
xnor U6820 (N_6820,N_5947,N_5227);
and U6821 (N_6821,N_5233,N_4474);
and U6822 (N_6822,N_5339,N_4956);
and U6823 (N_6823,N_5271,N_5157);
nand U6824 (N_6824,N_5508,N_5191);
xnor U6825 (N_6825,N_5135,N_4018);
nor U6826 (N_6826,N_5666,N_4783);
xnor U6827 (N_6827,N_5205,N_5276);
nor U6828 (N_6828,N_5460,N_5904);
and U6829 (N_6829,N_4288,N_5992);
nor U6830 (N_6830,N_4299,N_5785);
nor U6831 (N_6831,N_4692,N_5084);
nor U6832 (N_6832,N_4113,N_5978);
and U6833 (N_6833,N_4165,N_4362);
or U6834 (N_6834,N_5769,N_5574);
nand U6835 (N_6835,N_5125,N_4122);
xor U6836 (N_6836,N_4854,N_5362);
xnor U6837 (N_6837,N_5133,N_5173);
xnor U6838 (N_6838,N_4967,N_4572);
nor U6839 (N_6839,N_5048,N_5222);
nand U6840 (N_6840,N_4100,N_5347);
and U6841 (N_6841,N_4186,N_5179);
nand U6842 (N_6842,N_4521,N_4867);
or U6843 (N_6843,N_4401,N_4027);
xor U6844 (N_6844,N_5581,N_5701);
or U6845 (N_6845,N_4807,N_4651);
and U6846 (N_6846,N_5217,N_5853);
xor U6847 (N_6847,N_5750,N_4484);
xnor U6848 (N_6848,N_4106,N_4061);
nor U6849 (N_6849,N_4712,N_5876);
and U6850 (N_6850,N_4170,N_5968);
nand U6851 (N_6851,N_4869,N_5603);
nand U6852 (N_6852,N_4427,N_5068);
xnor U6853 (N_6853,N_4574,N_5190);
xnor U6854 (N_6854,N_5225,N_5816);
nor U6855 (N_6855,N_4499,N_4958);
xnor U6856 (N_6856,N_4769,N_4579);
or U6857 (N_6857,N_4996,N_4009);
xnor U6858 (N_6858,N_4417,N_4292);
xor U6859 (N_6859,N_5628,N_4992);
or U6860 (N_6860,N_5884,N_4564);
nand U6861 (N_6861,N_4239,N_5406);
nor U6862 (N_6862,N_5684,N_5183);
nand U6863 (N_6863,N_5032,N_4283);
xor U6864 (N_6864,N_4354,N_5441);
and U6865 (N_6865,N_4654,N_4655);
and U6866 (N_6866,N_5162,N_5676);
nand U6867 (N_6867,N_5255,N_4571);
xor U6868 (N_6868,N_4560,N_4166);
and U6869 (N_6869,N_5680,N_5539);
or U6870 (N_6870,N_4886,N_5387);
nor U6871 (N_6871,N_4071,N_5937);
nand U6872 (N_6872,N_5491,N_4810);
nand U6873 (N_6873,N_4021,N_5961);
or U6874 (N_6874,N_5453,N_4660);
xor U6875 (N_6875,N_5353,N_5417);
or U6876 (N_6876,N_5037,N_5226);
nand U6877 (N_6877,N_5568,N_4374);
nand U6878 (N_6878,N_5681,N_4930);
or U6879 (N_6879,N_4834,N_5633);
xor U6880 (N_6880,N_4211,N_5525);
nand U6881 (N_6881,N_5722,N_4432);
nor U6882 (N_6882,N_4226,N_4384);
xor U6883 (N_6883,N_4658,N_4406);
nor U6884 (N_6884,N_4421,N_4000);
nor U6885 (N_6885,N_4453,N_5461);
nor U6886 (N_6886,N_4031,N_5821);
nor U6887 (N_6887,N_5043,N_5913);
nand U6888 (N_6888,N_5687,N_4648);
nand U6889 (N_6889,N_5323,N_5411);
nor U6890 (N_6890,N_4626,N_5459);
nor U6891 (N_6891,N_4812,N_4310);
xnor U6892 (N_6892,N_4224,N_4156);
and U6893 (N_6893,N_5997,N_5873);
xnor U6894 (N_6894,N_5049,N_5103);
and U6895 (N_6895,N_4422,N_4929);
and U6896 (N_6896,N_5818,N_4512);
and U6897 (N_6897,N_5161,N_5029);
and U6898 (N_6898,N_4608,N_5772);
nand U6899 (N_6899,N_5155,N_5288);
xor U6900 (N_6900,N_5872,N_4385);
or U6901 (N_6901,N_4563,N_4228);
and U6902 (N_6902,N_5656,N_5757);
nor U6903 (N_6903,N_5196,N_5011);
xnor U6904 (N_6904,N_5343,N_4035);
nand U6905 (N_6905,N_4518,N_5207);
and U6906 (N_6906,N_5987,N_4237);
and U6907 (N_6907,N_4127,N_4590);
or U6908 (N_6908,N_4480,N_5694);
and U6909 (N_6909,N_5967,N_5792);
nor U6910 (N_6910,N_4848,N_5370);
xor U6911 (N_6911,N_4787,N_5311);
xnor U6912 (N_6912,N_5804,N_5923);
xnor U6913 (N_6913,N_4548,N_5069);
nor U6914 (N_6914,N_4508,N_5643);
or U6915 (N_6915,N_5768,N_4921);
nor U6916 (N_6916,N_4424,N_5809);
nor U6917 (N_6917,N_5279,N_5744);
and U6918 (N_6918,N_5589,N_5784);
nand U6919 (N_6919,N_4645,N_4163);
xnor U6920 (N_6920,N_4901,N_5467);
nand U6921 (N_6921,N_4699,N_4243);
nand U6922 (N_6922,N_5072,N_4078);
or U6923 (N_6923,N_5865,N_4053);
nor U6924 (N_6924,N_5231,N_5753);
xnor U6925 (N_6925,N_4280,N_5298);
nand U6926 (N_6926,N_4978,N_5583);
xnor U6927 (N_6927,N_5917,N_5609);
or U6928 (N_6928,N_5541,N_4950);
nor U6929 (N_6929,N_5535,N_4398);
nand U6930 (N_6930,N_4347,N_5127);
or U6931 (N_6931,N_5717,N_5351);
xor U6932 (N_6932,N_5092,N_5691);
and U6933 (N_6933,N_5941,N_4770);
xor U6934 (N_6934,N_4698,N_4195);
xor U6935 (N_6935,N_4339,N_4659);
nand U6936 (N_6936,N_4636,N_4328);
nor U6937 (N_6937,N_5325,N_4120);
or U6938 (N_6938,N_5210,N_5848);
or U6939 (N_6939,N_4447,N_5143);
xor U6940 (N_6940,N_4961,N_4885);
nor U6941 (N_6941,N_4507,N_5089);
nand U6942 (N_6942,N_4740,N_5355);
nand U6943 (N_6943,N_5281,N_4286);
or U6944 (N_6944,N_5451,N_5002);
nand U6945 (N_6945,N_4437,N_5567);
or U6946 (N_6946,N_5333,N_4721);
and U6947 (N_6947,N_4584,N_4117);
and U6948 (N_6948,N_5724,N_5882);
nand U6949 (N_6949,N_4293,N_4666);
or U6950 (N_6950,N_4350,N_5345);
nand U6951 (N_6951,N_4272,N_4466);
or U6952 (N_6952,N_4389,N_5599);
or U6953 (N_6953,N_5171,N_4792);
nor U6954 (N_6954,N_4324,N_4359);
or U6955 (N_6955,N_5174,N_4303);
nor U6956 (N_6956,N_5078,N_4509);
or U6957 (N_6957,N_5466,N_4452);
nor U6958 (N_6958,N_5817,N_5140);
nand U6959 (N_6959,N_5324,N_4979);
xor U6960 (N_6960,N_4764,N_4188);
xnor U6961 (N_6961,N_5204,N_4839);
nand U6962 (N_6962,N_5357,N_4547);
nand U6963 (N_6963,N_4248,N_4986);
nand U6964 (N_6964,N_5756,N_4148);
and U6965 (N_6965,N_4999,N_5986);
nor U6966 (N_6966,N_5927,N_5789);
or U6967 (N_6967,N_4183,N_5306);
nor U6968 (N_6968,N_4504,N_4937);
or U6969 (N_6969,N_5586,N_5646);
xnor U6970 (N_6970,N_5289,N_4905);
or U6971 (N_6971,N_4282,N_4143);
xor U6972 (N_6972,N_5580,N_5106);
xor U6973 (N_6973,N_5215,N_4436);
and U6974 (N_6974,N_4334,N_5197);
and U6975 (N_6975,N_4727,N_4568);
and U6976 (N_6976,N_5206,N_5570);
nor U6977 (N_6977,N_4019,N_5035);
and U6978 (N_6978,N_5138,N_5478);
nor U6979 (N_6979,N_5892,N_5623);
xnor U6980 (N_6980,N_5989,N_4731);
nand U6981 (N_6981,N_5790,N_4150);
or U6982 (N_6982,N_4235,N_4365);
nand U6983 (N_6983,N_4695,N_5641);
nor U6984 (N_6984,N_4450,N_4696);
nand U6985 (N_6985,N_5835,N_4115);
xor U6986 (N_6986,N_4209,N_4121);
nor U6987 (N_6987,N_4550,N_4316);
or U6988 (N_6988,N_5742,N_4130);
nand U6989 (N_6989,N_5273,N_4684);
or U6990 (N_6990,N_5921,N_5083);
xnor U6991 (N_6991,N_4162,N_4569);
xor U6992 (N_6992,N_5585,N_5374);
nand U6993 (N_6993,N_4255,N_5727);
nor U6994 (N_6994,N_5336,N_5657);
xnor U6995 (N_6995,N_4878,N_4168);
and U6996 (N_6996,N_5300,N_5291);
and U6997 (N_6997,N_4085,N_4933);
xnor U6998 (N_6998,N_4679,N_5658);
nand U6999 (N_6999,N_5971,N_5455);
xor U7000 (N_7000,N_4669,N_4667);
nand U7001 (N_7001,N_5468,N_5113);
or U7002 (N_7002,N_5103,N_4643);
nor U7003 (N_7003,N_5712,N_4353);
and U7004 (N_7004,N_5385,N_5017);
nand U7005 (N_7005,N_5346,N_4767);
nand U7006 (N_7006,N_5895,N_5214);
nand U7007 (N_7007,N_5293,N_5422);
or U7008 (N_7008,N_5540,N_5884);
nand U7009 (N_7009,N_4155,N_5347);
nand U7010 (N_7010,N_4038,N_5302);
or U7011 (N_7011,N_4592,N_5129);
or U7012 (N_7012,N_4699,N_4693);
and U7013 (N_7013,N_4733,N_4666);
or U7014 (N_7014,N_4258,N_5474);
or U7015 (N_7015,N_4630,N_4738);
and U7016 (N_7016,N_4136,N_5993);
and U7017 (N_7017,N_4596,N_5292);
and U7018 (N_7018,N_5626,N_4545);
and U7019 (N_7019,N_5432,N_4687);
nand U7020 (N_7020,N_4771,N_5231);
and U7021 (N_7021,N_4480,N_4488);
nand U7022 (N_7022,N_5561,N_5488);
nand U7023 (N_7023,N_4805,N_5679);
nor U7024 (N_7024,N_4071,N_5849);
or U7025 (N_7025,N_4987,N_4509);
nor U7026 (N_7026,N_5154,N_5086);
xnor U7027 (N_7027,N_4473,N_4195);
nor U7028 (N_7028,N_5407,N_5006);
or U7029 (N_7029,N_4510,N_4529);
or U7030 (N_7030,N_5043,N_5875);
nor U7031 (N_7031,N_5094,N_4909);
or U7032 (N_7032,N_4179,N_5715);
or U7033 (N_7033,N_4548,N_5454);
nor U7034 (N_7034,N_5768,N_4623);
or U7035 (N_7035,N_5881,N_4185);
nand U7036 (N_7036,N_4731,N_5037);
and U7037 (N_7037,N_5104,N_4128);
or U7038 (N_7038,N_4953,N_4348);
xnor U7039 (N_7039,N_4624,N_4139);
and U7040 (N_7040,N_5665,N_4364);
nand U7041 (N_7041,N_4943,N_5726);
nand U7042 (N_7042,N_4222,N_5619);
and U7043 (N_7043,N_5569,N_5676);
xor U7044 (N_7044,N_4763,N_5780);
nor U7045 (N_7045,N_5320,N_4589);
or U7046 (N_7046,N_4513,N_4283);
xnor U7047 (N_7047,N_4558,N_5710);
or U7048 (N_7048,N_4346,N_4878);
xnor U7049 (N_7049,N_4790,N_5145);
nand U7050 (N_7050,N_4213,N_5111);
nor U7051 (N_7051,N_4389,N_4294);
and U7052 (N_7052,N_5030,N_4058);
nor U7053 (N_7053,N_5408,N_4574);
or U7054 (N_7054,N_4439,N_4209);
and U7055 (N_7055,N_4530,N_4754);
xnor U7056 (N_7056,N_5831,N_5065);
and U7057 (N_7057,N_5717,N_5704);
and U7058 (N_7058,N_5690,N_4810);
xor U7059 (N_7059,N_4190,N_4800);
or U7060 (N_7060,N_4046,N_4002);
or U7061 (N_7061,N_5056,N_5758);
and U7062 (N_7062,N_4403,N_5619);
and U7063 (N_7063,N_4727,N_5089);
xnor U7064 (N_7064,N_4712,N_4318);
xnor U7065 (N_7065,N_5719,N_5872);
nor U7066 (N_7066,N_4937,N_4491);
nor U7067 (N_7067,N_4007,N_5409);
and U7068 (N_7068,N_5435,N_4980);
or U7069 (N_7069,N_4709,N_4202);
nand U7070 (N_7070,N_4811,N_4358);
and U7071 (N_7071,N_5119,N_4702);
nand U7072 (N_7072,N_4229,N_5492);
nor U7073 (N_7073,N_5214,N_4964);
nand U7074 (N_7074,N_5372,N_4916);
nor U7075 (N_7075,N_5899,N_4810);
xnor U7076 (N_7076,N_5763,N_4709);
nand U7077 (N_7077,N_4277,N_5528);
or U7078 (N_7078,N_4558,N_5974);
nand U7079 (N_7079,N_4018,N_4472);
nand U7080 (N_7080,N_5803,N_4266);
xnor U7081 (N_7081,N_5096,N_5806);
or U7082 (N_7082,N_5238,N_5099);
or U7083 (N_7083,N_4626,N_4629);
and U7084 (N_7084,N_5073,N_4604);
and U7085 (N_7085,N_4020,N_4029);
nor U7086 (N_7086,N_4148,N_5895);
and U7087 (N_7087,N_5284,N_4470);
and U7088 (N_7088,N_5638,N_4904);
nand U7089 (N_7089,N_4172,N_4257);
nor U7090 (N_7090,N_4688,N_4804);
nand U7091 (N_7091,N_5322,N_5548);
nand U7092 (N_7092,N_4743,N_5918);
xor U7093 (N_7093,N_5771,N_4956);
nor U7094 (N_7094,N_5596,N_4570);
nand U7095 (N_7095,N_5527,N_4190);
and U7096 (N_7096,N_4837,N_4148);
xor U7097 (N_7097,N_4878,N_5157);
xor U7098 (N_7098,N_5502,N_5984);
or U7099 (N_7099,N_4379,N_4806);
xor U7100 (N_7100,N_4296,N_4720);
and U7101 (N_7101,N_5101,N_4050);
and U7102 (N_7102,N_4845,N_4826);
or U7103 (N_7103,N_5955,N_4963);
nand U7104 (N_7104,N_4531,N_5217);
nand U7105 (N_7105,N_4544,N_5732);
and U7106 (N_7106,N_5444,N_4197);
and U7107 (N_7107,N_4069,N_4094);
and U7108 (N_7108,N_5149,N_4037);
nor U7109 (N_7109,N_5938,N_4526);
nand U7110 (N_7110,N_4734,N_5415);
and U7111 (N_7111,N_5906,N_4648);
nor U7112 (N_7112,N_5714,N_5753);
and U7113 (N_7113,N_5193,N_4075);
xnor U7114 (N_7114,N_5644,N_4370);
nor U7115 (N_7115,N_5850,N_4119);
or U7116 (N_7116,N_4839,N_5550);
nand U7117 (N_7117,N_4159,N_5702);
xor U7118 (N_7118,N_5802,N_4690);
or U7119 (N_7119,N_5837,N_5852);
nand U7120 (N_7120,N_4158,N_5659);
or U7121 (N_7121,N_4364,N_4915);
and U7122 (N_7122,N_4497,N_4610);
xnor U7123 (N_7123,N_4384,N_4298);
xor U7124 (N_7124,N_4887,N_5539);
and U7125 (N_7125,N_5491,N_4758);
xnor U7126 (N_7126,N_5310,N_5484);
nor U7127 (N_7127,N_4246,N_4583);
xor U7128 (N_7128,N_4321,N_4590);
nand U7129 (N_7129,N_4635,N_4631);
nand U7130 (N_7130,N_5085,N_5784);
xnor U7131 (N_7131,N_5094,N_4789);
xnor U7132 (N_7132,N_5482,N_4605);
xor U7133 (N_7133,N_4943,N_5663);
nor U7134 (N_7134,N_5983,N_5055);
nand U7135 (N_7135,N_4695,N_4371);
and U7136 (N_7136,N_4312,N_5376);
nand U7137 (N_7137,N_5784,N_5095);
and U7138 (N_7138,N_4810,N_4339);
xnor U7139 (N_7139,N_5612,N_4678);
nor U7140 (N_7140,N_4881,N_5285);
and U7141 (N_7141,N_4094,N_4766);
or U7142 (N_7142,N_4474,N_5612);
and U7143 (N_7143,N_4334,N_4990);
xor U7144 (N_7144,N_5085,N_5229);
nand U7145 (N_7145,N_4240,N_5863);
and U7146 (N_7146,N_5966,N_4633);
and U7147 (N_7147,N_4792,N_4187);
nand U7148 (N_7148,N_4313,N_4440);
or U7149 (N_7149,N_4504,N_4490);
xor U7150 (N_7150,N_4733,N_4793);
nor U7151 (N_7151,N_5029,N_4432);
or U7152 (N_7152,N_4924,N_4279);
and U7153 (N_7153,N_4381,N_5323);
nor U7154 (N_7154,N_4925,N_4977);
xor U7155 (N_7155,N_5655,N_4073);
nand U7156 (N_7156,N_4715,N_4684);
xor U7157 (N_7157,N_5855,N_5587);
xor U7158 (N_7158,N_5902,N_4706);
nand U7159 (N_7159,N_4961,N_5727);
xor U7160 (N_7160,N_5132,N_4222);
or U7161 (N_7161,N_5737,N_5880);
xor U7162 (N_7162,N_5120,N_4110);
nor U7163 (N_7163,N_5729,N_5373);
nor U7164 (N_7164,N_4823,N_5464);
and U7165 (N_7165,N_5257,N_4878);
nand U7166 (N_7166,N_4185,N_5681);
nand U7167 (N_7167,N_4929,N_4472);
nor U7168 (N_7168,N_4881,N_5203);
xnor U7169 (N_7169,N_4834,N_4236);
nor U7170 (N_7170,N_5240,N_4431);
and U7171 (N_7171,N_5919,N_5910);
nand U7172 (N_7172,N_5101,N_5945);
nand U7173 (N_7173,N_4809,N_4085);
nor U7174 (N_7174,N_5851,N_4818);
nor U7175 (N_7175,N_5143,N_5571);
and U7176 (N_7176,N_5309,N_5315);
and U7177 (N_7177,N_5942,N_5352);
xor U7178 (N_7178,N_4772,N_5146);
xor U7179 (N_7179,N_4424,N_5402);
xor U7180 (N_7180,N_5468,N_5545);
or U7181 (N_7181,N_4619,N_4519);
and U7182 (N_7182,N_5036,N_5985);
and U7183 (N_7183,N_4101,N_4459);
xor U7184 (N_7184,N_4356,N_4571);
xor U7185 (N_7185,N_5672,N_4772);
and U7186 (N_7186,N_5366,N_4807);
xnor U7187 (N_7187,N_5627,N_5866);
and U7188 (N_7188,N_5507,N_5330);
nor U7189 (N_7189,N_4009,N_5941);
nor U7190 (N_7190,N_5605,N_5542);
and U7191 (N_7191,N_5358,N_5200);
or U7192 (N_7192,N_5456,N_4756);
or U7193 (N_7193,N_5108,N_5735);
nand U7194 (N_7194,N_5241,N_5405);
nand U7195 (N_7195,N_4181,N_5003);
nor U7196 (N_7196,N_4815,N_5345);
and U7197 (N_7197,N_5562,N_4315);
or U7198 (N_7198,N_5552,N_5168);
nor U7199 (N_7199,N_4912,N_4186);
nor U7200 (N_7200,N_4659,N_5988);
and U7201 (N_7201,N_4093,N_5504);
nand U7202 (N_7202,N_5824,N_4667);
nand U7203 (N_7203,N_4463,N_4603);
or U7204 (N_7204,N_5967,N_5612);
nand U7205 (N_7205,N_4286,N_5421);
nor U7206 (N_7206,N_5749,N_4797);
nand U7207 (N_7207,N_4569,N_5525);
xor U7208 (N_7208,N_4865,N_5235);
nand U7209 (N_7209,N_5409,N_5711);
nand U7210 (N_7210,N_4487,N_4763);
or U7211 (N_7211,N_5135,N_5789);
nand U7212 (N_7212,N_5174,N_5441);
xor U7213 (N_7213,N_4127,N_5648);
xor U7214 (N_7214,N_4106,N_5845);
and U7215 (N_7215,N_4718,N_4387);
nand U7216 (N_7216,N_5595,N_5274);
nor U7217 (N_7217,N_5592,N_4724);
and U7218 (N_7218,N_5337,N_5883);
nand U7219 (N_7219,N_4657,N_5064);
and U7220 (N_7220,N_4316,N_5478);
and U7221 (N_7221,N_5445,N_4380);
and U7222 (N_7222,N_5304,N_5231);
and U7223 (N_7223,N_4502,N_5605);
xnor U7224 (N_7224,N_4051,N_4430);
or U7225 (N_7225,N_5893,N_4164);
nor U7226 (N_7226,N_4369,N_5393);
xor U7227 (N_7227,N_4800,N_5224);
xnor U7228 (N_7228,N_4477,N_4078);
xor U7229 (N_7229,N_4689,N_5795);
nor U7230 (N_7230,N_4872,N_4989);
or U7231 (N_7231,N_4128,N_5108);
nor U7232 (N_7232,N_4146,N_4474);
and U7233 (N_7233,N_5135,N_5497);
and U7234 (N_7234,N_5198,N_5591);
nor U7235 (N_7235,N_5589,N_4529);
xnor U7236 (N_7236,N_5376,N_5403);
xor U7237 (N_7237,N_5139,N_5632);
nand U7238 (N_7238,N_4823,N_5915);
nand U7239 (N_7239,N_5653,N_4164);
nand U7240 (N_7240,N_5599,N_5042);
xor U7241 (N_7241,N_4836,N_5719);
xor U7242 (N_7242,N_5746,N_5649);
and U7243 (N_7243,N_4102,N_5661);
nand U7244 (N_7244,N_5462,N_4731);
nor U7245 (N_7245,N_4798,N_4634);
nor U7246 (N_7246,N_5355,N_5236);
and U7247 (N_7247,N_5613,N_5027);
nor U7248 (N_7248,N_4987,N_5141);
xnor U7249 (N_7249,N_5217,N_4929);
and U7250 (N_7250,N_5291,N_4141);
xor U7251 (N_7251,N_5012,N_5033);
nand U7252 (N_7252,N_5440,N_4442);
nor U7253 (N_7253,N_4179,N_4158);
nand U7254 (N_7254,N_5135,N_4416);
nor U7255 (N_7255,N_4073,N_5743);
nand U7256 (N_7256,N_4105,N_5012);
nand U7257 (N_7257,N_4576,N_5116);
or U7258 (N_7258,N_5331,N_5406);
nor U7259 (N_7259,N_5755,N_4097);
xnor U7260 (N_7260,N_4562,N_5317);
nor U7261 (N_7261,N_4083,N_4834);
nor U7262 (N_7262,N_5548,N_5124);
xnor U7263 (N_7263,N_5023,N_4733);
xnor U7264 (N_7264,N_5756,N_4236);
nand U7265 (N_7265,N_4433,N_5619);
nand U7266 (N_7266,N_4417,N_4918);
nor U7267 (N_7267,N_5415,N_4607);
nand U7268 (N_7268,N_4283,N_4681);
and U7269 (N_7269,N_5269,N_4683);
nor U7270 (N_7270,N_4865,N_5262);
or U7271 (N_7271,N_5946,N_5769);
xnor U7272 (N_7272,N_4368,N_4941);
or U7273 (N_7273,N_4388,N_4271);
nand U7274 (N_7274,N_5931,N_5793);
and U7275 (N_7275,N_4205,N_4147);
and U7276 (N_7276,N_5592,N_5827);
nand U7277 (N_7277,N_4525,N_4394);
xor U7278 (N_7278,N_4399,N_4769);
nand U7279 (N_7279,N_4159,N_4205);
nor U7280 (N_7280,N_4792,N_4937);
nor U7281 (N_7281,N_5552,N_4694);
nand U7282 (N_7282,N_4098,N_5911);
nor U7283 (N_7283,N_4560,N_5644);
and U7284 (N_7284,N_5763,N_4656);
and U7285 (N_7285,N_5416,N_5272);
nor U7286 (N_7286,N_4297,N_5245);
and U7287 (N_7287,N_4323,N_4423);
xor U7288 (N_7288,N_5803,N_4386);
nor U7289 (N_7289,N_4620,N_5446);
xor U7290 (N_7290,N_5799,N_5431);
nand U7291 (N_7291,N_5821,N_4566);
nand U7292 (N_7292,N_5265,N_5657);
nor U7293 (N_7293,N_5288,N_4911);
nor U7294 (N_7294,N_4094,N_5043);
and U7295 (N_7295,N_5184,N_4389);
and U7296 (N_7296,N_5403,N_4626);
xor U7297 (N_7297,N_5604,N_4339);
nor U7298 (N_7298,N_5734,N_5722);
or U7299 (N_7299,N_5998,N_4076);
xor U7300 (N_7300,N_5971,N_5270);
and U7301 (N_7301,N_5208,N_4462);
or U7302 (N_7302,N_5834,N_5417);
nor U7303 (N_7303,N_5081,N_5502);
and U7304 (N_7304,N_5888,N_5974);
nor U7305 (N_7305,N_5224,N_4776);
xnor U7306 (N_7306,N_5567,N_5082);
nand U7307 (N_7307,N_4644,N_4280);
or U7308 (N_7308,N_5104,N_4676);
nor U7309 (N_7309,N_5608,N_5531);
or U7310 (N_7310,N_4467,N_4294);
nor U7311 (N_7311,N_4480,N_5309);
nand U7312 (N_7312,N_4943,N_5378);
xnor U7313 (N_7313,N_5308,N_5388);
or U7314 (N_7314,N_5290,N_5088);
nand U7315 (N_7315,N_5982,N_5365);
nor U7316 (N_7316,N_5140,N_4725);
nand U7317 (N_7317,N_5705,N_4248);
or U7318 (N_7318,N_4757,N_4188);
xor U7319 (N_7319,N_5015,N_5120);
or U7320 (N_7320,N_4658,N_5985);
nand U7321 (N_7321,N_4892,N_4773);
and U7322 (N_7322,N_5124,N_5143);
xnor U7323 (N_7323,N_4291,N_5855);
and U7324 (N_7324,N_4777,N_5184);
xnor U7325 (N_7325,N_5577,N_5746);
or U7326 (N_7326,N_5899,N_5631);
nand U7327 (N_7327,N_4225,N_5044);
and U7328 (N_7328,N_5592,N_4498);
xor U7329 (N_7329,N_5184,N_5381);
nor U7330 (N_7330,N_4874,N_5738);
or U7331 (N_7331,N_5712,N_5923);
and U7332 (N_7332,N_4252,N_4319);
xor U7333 (N_7333,N_5995,N_4096);
nand U7334 (N_7334,N_5146,N_4781);
and U7335 (N_7335,N_4532,N_5431);
and U7336 (N_7336,N_4223,N_5771);
nand U7337 (N_7337,N_5437,N_5273);
xor U7338 (N_7338,N_5937,N_4310);
nor U7339 (N_7339,N_4801,N_5693);
and U7340 (N_7340,N_4288,N_4529);
or U7341 (N_7341,N_5707,N_4864);
xor U7342 (N_7342,N_5097,N_4763);
and U7343 (N_7343,N_4676,N_4644);
and U7344 (N_7344,N_5807,N_4010);
and U7345 (N_7345,N_5100,N_5896);
and U7346 (N_7346,N_5453,N_5810);
or U7347 (N_7347,N_5621,N_4458);
nor U7348 (N_7348,N_5505,N_4927);
nand U7349 (N_7349,N_4613,N_5386);
xnor U7350 (N_7350,N_4805,N_5362);
or U7351 (N_7351,N_5207,N_5555);
nand U7352 (N_7352,N_5173,N_4706);
xnor U7353 (N_7353,N_4110,N_5431);
nand U7354 (N_7354,N_4937,N_4865);
nor U7355 (N_7355,N_4648,N_5893);
and U7356 (N_7356,N_5575,N_5595);
xor U7357 (N_7357,N_4246,N_4941);
or U7358 (N_7358,N_5058,N_4198);
xor U7359 (N_7359,N_4823,N_4277);
nand U7360 (N_7360,N_5724,N_5062);
nor U7361 (N_7361,N_5165,N_5119);
xor U7362 (N_7362,N_5623,N_5503);
nor U7363 (N_7363,N_4112,N_5107);
and U7364 (N_7364,N_5363,N_4095);
xnor U7365 (N_7365,N_5492,N_5563);
or U7366 (N_7366,N_4785,N_4033);
nor U7367 (N_7367,N_4368,N_5868);
nand U7368 (N_7368,N_5880,N_4397);
xor U7369 (N_7369,N_4087,N_4327);
and U7370 (N_7370,N_5140,N_4717);
or U7371 (N_7371,N_4740,N_5398);
or U7372 (N_7372,N_4886,N_5795);
nor U7373 (N_7373,N_5224,N_5492);
xnor U7374 (N_7374,N_4380,N_4980);
nor U7375 (N_7375,N_4769,N_4759);
xor U7376 (N_7376,N_5152,N_5999);
xor U7377 (N_7377,N_5351,N_5057);
nor U7378 (N_7378,N_5706,N_4745);
xor U7379 (N_7379,N_5078,N_4288);
nand U7380 (N_7380,N_5555,N_5938);
nor U7381 (N_7381,N_4343,N_4627);
and U7382 (N_7382,N_4855,N_5555);
nand U7383 (N_7383,N_4702,N_4404);
and U7384 (N_7384,N_5330,N_4099);
or U7385 (N_7385,N_4966,N_4777);
and U7386 (N_7386,N_4873,N_4889);
and U7387 (N_7387,N_5124,N_5827);
xor U7388 (N_7388,N_4536,N_4786);
and U7389 (N_7389,N_5478,N_5533);
nand U7390 (N_7390,N_4051,N_5132);
nand U7391 (N_7391,N_4743,N_4016);
and U7392 (N_7392,N_4083,N_4911);
and U7393 (N_7393,N_5963,N_5123);
nand U7394 (N_7394,N_4805,N_4671);
nor U7395 (N_7395,N_5489,N_4096);
nor U7396 (N_7396,N_4174,N_4014);
or U7397 (N_7397,N_4976,N_5427);
nor U7398 (N_7398,N_4445,N_4905);
nand U7399 (N_7399,N_4121,N_5259);
and U7400 (N_7400,N_5244,N_5300);
nand U7401 (N_7401,N_4563,N_5047);
and U7402 (N_7402,N_4798,N_4606);
nor U7403 (N_7403,N_4375,N_4063);
or U7404 (N_7404,N_5828,N_5990);
nand U7405 (N_7405,N_5294,N_4929);
nand U7406 (N_7406,N_4509,N_5797);
nor U7407 (N_7407,N_5983,N_5187);
and U7408 (N_7408,N_5248,N_5710);
xnor U7409 (N_7409,N_5467,N_5886);
nor U7410 (N_7410,N_5445,N_4146);
or U7411 (N_7411,N_5925,N_4605);
xnor U7412 (N_7412,N_4251,N_5357);
or U7413 (N_7413,N_5579,N_4173);
nor U7414 (N_7414,N_5320,N_5125);
nand U7415 (N_7415,N_4892,N_4180);
nor U7416 (N_7416,N_4844,N_4519);
xnor U7417 (N_7417,N_5891,N_4862);
or U7418 (N_7418,N_4393,N_5431);
nor U7419 (N_7419,N_4037,N_4118);
xnor U7420 (N_7420,N_4591,N_5276);
nor U7421 (N_7421,N_4924,N_5202);
nor U7422 (N_7422,N_5642,N_5781);
nor U7423 (N_7423,N_5683,N_4806);
xnor U7424 (N_7424,N_4175,N_4488);
xor U7425 (N_7425,N_4275,N_5834);
nor U7426 (N_7426,N_5737,N_4144);
nand U7427 (N_7427,N_5921,N_4317);
xnor U7428 (N_7428,N_5661,N_5929);
and U7429 (N_7429,N_5695,N_4061);
nand U7430 (N_7430,N_5952,N_5743);
and U7431 (N_7431,N_4626,N_4415);
nor U7432 (N_7432,N_5202,N_4880);
xor U7433 (N_7433,N_4942,N_4443);
and U7434 (N_7434,N_4175,N_5019);
or U7435 (N_7435,N_5398,N_4121);
or U7436 (N_7436,N_4891,N_4178);
nor U7437 (N_7437,N_5465,N_4660);
nand U7438 (N_7438,N_5034,N_5720);
nand U7439 (N_7439,N_4162,N_4136);
xor U7440 (N_7440,N_4465,N_5179);
xor U7441 (N_7441,N_5774,N_5278);
and U7442 (N_7442,N_4677,N_4996);
or U7443 (N_7443,N_5397,N_4965);
nor U7444 (N_7444,N_4449,N_4136);
or U7445 (N_7445,N_5001,N_4873);
and U7446 (N_7446,N_4468,N_5702);
nor U7447 (N_7447,N_4502,N_4124);
and U7448 (N_7448,N_4703,N_4101);
and U7449 (N_7449,N_5913,N_5426);
xnor U7450 (N_7450,N_4258,N_4186);
or U7451 (N_7451,N_5036,N_4630);
nand U7452 (N_7452,N_5424,N_5108);
and U7453 (N_7453,N_4934,N_4281);
or U7454 (N_7454,N_5046,N_5930);
xnor U7455 (N_7455,N_4617,N_4662);
xnor U7456 (N_7456,N_5099,N_4046);
or U7457 (N_7457,N_5383,N_4086);
or U7458 (N_7458,N_5814,N_4162);
nand U7459 (N_7459,N_4835,N_5645);
or U7460 (N_7460,N_5204,N_4157);
xor U7461 (N_7461,N_4251,N_5899);
nor U7462 (N_7462,N_5115,N_5781);
or U7463 (N_7463,N_4169,N_4627);
nor U7464 (N_7464,N_4172,N_5486);
nand U7465 (N_7465,N_4219,N_4630);
nor U7466 (N_7466,N_4957,N_5908);
or U7467 (N_7467,N_5110,N_5778);
and U7468 (N_7468,N_5955,N_4426);
or U7469 (N_7469,N_4638,N_4734);
or U7470 (N_7470,N_5386,N_5514);
or U7471 (N_7471,N_4507,N_5617);
nand U7472 (N_7472,N_5054,N_5340);
nor U7473 (N_7473,N_4375,N_5790);
nor U7474 (N_7474,N_4076,N_5425);
and U7475 (N_7475,N_5862,N_5651);
or U7476 (N_7476,N_4208,N_4803);
xnor U7477 (N_7477,N_4747,N_5690);
nor U7478 (N_7478,N_4792,N_4268);
and U7479 (N_7479,N_5313,N_5662);
nand U7480 (N_7480,N_4705,N_5209);
nand U7481 (N_7481,N_4995,N_5372);
nand U7482 (N_7482,N_4680,N_5456);
xor U7483 (N_7483,N_5883,N_5525);
and U7484 (N_7484,N_4610,N_5278);
nor U7485 (N_7485,N_5240,N_5058);
xnor U7486 (N_7486,N_4827,N_4028);
or U7487 (N_7487,N_4373,N_4013);
nor U7488 (N_7488,N_4460,N_4704);
xor U7489 (N_7489,N_5254,N_4870);
and U7490 (N_7490,N_4299,N_5837);
or U7491 (N_7491,N_5733,N_4563);
nor U7492 (N_7492,N_4498,N_5181);
nand U7493 (N_7493,N_5745,N_4645);
nand U7494 (N_7494,N_5298,N_5459);
or U7495 (N_7495,N_5059,N_4319);
xor U7496 (N_7496,N_4971,N_5823);
xor U7497 (N_7497,N_5370,N_5102);
xor U7498 (N_7498,N_4292,N_4418);
and U7499 (N_7499,N_4562,N_5786);
and U7500 (N_7500,N_4760,N_4333);
nand U7501 (N_7501,N_4065,N_5411);
nor U7502 (N_7502,N_5514,N_5368);
nor U7503 (N_7503,N_5741,N_4518);
or U7504 (N_7504,N_5996,N_5180);
nand U7505 (N_7505,N_5969,N_5858);
and U7506 (N_7506,N_4675,N_5014);
and U7507 (N_7507,N_4979,N_4861);
xor U7508 (N_7508,N_5274,N_5854);
nor U7509 (N_7509,N_4464,N_5174);
nor U7510 (N_7510,N_5787,N_4834);
or U7511 (N_7511,N_4012,N_4404);
or U7512 (N_7512,N_4032,N_4109);
xor U7513 (N_7513,N_5230,N_5768);
and U7514 (N_7514,N_4779,N_5535);
nor U7515 (N_7515,N_4327,N_5285);
nand U7516 (N_7516,N_4529,N_4046);
xnor U7517 (N_7517,N_5975,N_5516);
or U7518 (N_7518,N_4154,N_5453);
or U7519 (N_7519,N_5741,N_5356);
nand U7520 (N_7520,N_4795,N_4568);
nand U7521 (N_7521,N_5616,N_4098);
nor U7522 (N_7522,N_4851,N_4661);
xor U7523 (N_7523,N_5264,N_4812);
nand U7524 (N_7524,N_4554,N_4664);
nor U7525 (N_7525,N_5738,N_5244);
nand U7526 (N_7526,N_4039,N_4450);
nand U7527 (N_7527,N_5304,N_4301);
nor U7528 (N_7528,N_5374,N_4774);
or U7529 (N_7529,N_4447,N_5125);
nand U7530 (N_7530,N_5122,N_4165);
nor U7531 (N_7531,N_4342,N_5589);
xnor U7532 (N_7532,N_5777,N_4141);
nand U7533 (N_7533,N_5247,N_4034);
xnor U7534 (N_7534,N_5975,N_5347);
xor U7535 (N_7535,N_5631,N_5052);
or U7536 (N_7536,N_5671,N_5565);
and U7537 (N_7537,N_5315,N_4691);
and U7538 (N_7538,N_5709,N_5543);
xor U7539 (N_7539,N_5313,N_4971);
and U7540 (N_7540,N_5846,N_5343);
nand U7541 (N_7541,N_4940,N_4761);
nor U7542 (N_7542,N_5683,N_5439);
or U7543 (N_7543,N_4244,N_4938);
nand U7544 (N_7544,N_4757,N_4567);
and U7545 (N_7545,N_4138,N_4038);
and U7546 (N_7546,N_4701,N_5929);
xnor U7547 (N_7547,N_5896,N_5452);
or U7548 (N_7548,N_4215,N_4761);
nor U7549 (N_7549,N_5044,N_4679);
or U7550 (N_7550,N_4159,N_5271);
xor U7551 (N_7551,N_4984,N_5587);
and U7552 (N_7552,N_5576,N_4116);
xnor U7553 (N_7553,N_5242,N_5067);
xor U7554 (N_7554,N_4895,N_5165);
nand U7555 (N_7555,N_4836,N_5063);
or U7556 (N_7556,N_5222,N_5873);
xnor U7557 (N_7557,N_5667,N_4404);
nand U7558 (N_7558,N_4340,N_5132);
nor U7559 (N_7559,N_4690,N_5958);
xnor U7560 (N_7560,N_5584,N_4403);
and U7561 (N_7561,N_5107,N_5340);
nand U7562 (N_7562,N_4744,N_5870);
and U7563 (N_7563,N_5266,N_5540);
nor U7564 (N_7564,N_5743,N_5865);
nor U7565 (N_7565,N_5977,N_4818);
or U7566 (N_7566,N_4314,N_5170);
and U7567 (N_7567,N_5881,N_4399);
nand U7568 (N_7568,N_4298,N_4339);
nand U7569 (N_7569,N_4760,N_5191);
xor U7570 (N_7570,N_5901,N_4699);
nand U7571 (N_7571,N_4386,N_4676);
and U7572 (N_7572,N_4422,N_4935);
or U7573 (N_7573,N_5337,N_4807);
xnor U7574 (N_7574,N_5027,N_4706);
nor U7575 (N_7575,N_4162,N_4120);
xnor U7576 (N_7576,N_4423,N_4829);
xor U7577 (N_7577,N_4883,N_5658);
nor U7578 (N_7578,N_4869,N_5732);
xor U7579 (N_7579,N_4608,N_5958);
xor U7580 (N_7580,N_5811,N_5190);
nor U7581 (N_7581,N_5020,N_5848);
and U7582 (N_7582,N_4663,N_5550);
or U7583 (N_7583,N_5568,N_4013);
xnor U7584 (N_7584,N_5118,N_5739);
xor U7585 (N_7585,N_5178,N_5572);
xor U7586 (N_7586,N_5890,N_5116);
xor U7587 (N_7587,N_4757,N_5931);
and U7588 (N_7588,N_4929,N_4446);
or U7589 (N_7589,N_5638,N_4944);
nand U7590 (N_7590,N_5876,N_4937);
xnor U7591 (N_7591,N_5675,N_4542);
xnor U7592 (N_7592,N_4026,N_4223);
xnor U7593 (N_7593,N_5289,N_5511);
or U7594 (N_7594,N_5741,N_5781);
xnor U7595 (N_7595,N_5104,N_4989);
or U7596 (N_7596,N_5863,N_5037);
nand U7597 (N_7597,N_4417,N_5669);
nor U7598 (N_7598,N_4561,N_4797);
or U7599 (N_7599,N_5452,N_5711);
nor U7600 (N_7600,N_5223,N_5969);
and U7601 (N_7601,N_5839,N_5652);
xnor U7602 (N_7602,N_5643,N_5109);
xor U7603 (N_7603,N_4305,N_4198);
xor U7604 (N_7604,N_4984,N_5616);
and U7605 (N_7605,N_4370,N_4393);
and U7606 (N_7606,N_5332,N_5331);
and U7607 (N_7607,N_5123,N_5654);
nand U7608 (N_7608,N_4329,N_4308);
nor U7609 (N_7609,N_4106,N_4140);
or U7610 (N_7610,N_5516,N_4768);
xor U7611 (N_7611,N_5908,N_4928);
nor U7612 (N_7612,N_4320,N_4026);
xor U7613 (N_7613,N_5727,N_4456);
nor U7614 (N_7614,N_5898,N_4859);
nand U7615 (N_7615,N_4313,N_5632);
nand U7616 (N_7616,N_4757,N_5068);
nand U7617 (N_7617,N_5659,N_5503);
xnor U7618 (N_7618,N_5957,N_4795);
xnor U7619 (N_7619,N_5392,N_4606);
xnor U7620 (N_7620,N_4879,N_4143);
nand U7621 (N_7621,N_5756,N_4364);
xor U7622 (N_7622,N_5570,N_5291);
or U7623 (N_7623,N_4169,N_4244);
nand U7624 (N_7624,N_4878,N_5521);
or U7625 (N_7625,N_5414,N_4590);
nor U7626 (N_7626,N_5486,N_4065);
or U7627 (N_7627,N_5837,N_4487);
nand U7628 (N_7628,N_5150,N_5496);
xor U7629 (N_7629,N_5144,N_5228);
nand U7630 (N_7630,N_4102,N_5624);
or U7631 (N_7631,N_4006,N_4823);
and U7632 (N_7632,N_4720,N_5279);
xnor U7633 (N_7633,N_4060,N_5428);
or U7634 (N_7634,N_5136,N_5939);
nor U7635 (N_7635,N_5881,N_4302);
and U7636 (N_7636,N_5907,N_4951);
xnor U7637 (N_7637,N_4774,N_5281);
nor U7638 (N_7638,N_5999,N_4064);
nor U7639 (N_7639,N_4188,N_4512);
nor U7640 (N_7640,N_5773,N_4789);
xnor U7641 (N_7641,N_5733,N_5425);
xor U7642 (N_7642,N_5141,N_5512);
nor U7643 (N_7643,N_4312,N_5413);
and U7644 (N_7644,N_4237,N_5016);
nor U7645 (N_7645,N_4270,N_5463);
nor U7646 (N_7646,N_5977,N_5444);
xnor U7647 (N_7647,N_5231,N_4761);
nor U7648 (N_7648,N_4827,N_4934);
and U7649 (N_7649,N_5456,N_5237);
xnor U7650 (N_7650,N_4797,N_5904);
or U7651 (N_7651,N_5114,N_4760);
or U7652 (N_7652,N_4554,N_5339);
xor U7653 (N_7653,N_5159,N_5293);
xnor U7654 (N_7654,N_4386,N_4161);
nand U7655 (N_7655,N_4828,N_5148);
xnor U7656 (N_7656,N_5013,N_5869);
nor U7657 (N_7657,N_5447,N_4354);
and U7658 (N_7658,N_4676,N_4206);
xor U7659 (N_7659,N_5048,N_5399);
or U7660 (N_7660,N_4271,N_5616);
nor U7661 (N_7661,N_4337,N_4116);
nand U7662 (N_7662,N_4898,N_4572);
xor U7663 (N_7663,N_4574,N_5043);
and U7664 (N_7664,N_4871,N_4689);
nor U7665 (N_7665,N_4600,N_5933);
xnor U7666 (N_7666,N_4157,N_4356);
and U7667 (N_7667,N_5869,N_4529);
nor U7668 (N_7668,N_5790,N_4968);
or U7669 (N_7669,N_4077,N_5758);
or U7670 (N_7670,N_4690,N_5718);
and U7671 (N_7671,N_4848,N_4438);
nor U7672 (N_7672,N_5005,N_4736);
nand U7673 (N_7673,N_4666,N_5247);
xor U7674 (N_7674,N_5491,N_5906);
or U7675 (N_7675,N_5253,N_5990);
and U7676 (N_7676,N_4210,N_4093);
nand U7677 (N_7677,N_4668,N_5343);
xnor U7678 (N_7678,N_4954,N_5042);
nand U7679 (N_7679,N_5077,N_5935);
nor U7680 (N_7680,N_5288,N_4019);
nor U7681 (N_7681,N_5109,N_4743);
nor U7682 (N_7682,N_4568,N_4297);
xnor U7683 (N_7683,N_4045,N_5386);
nor U7684 (N_7684,N_4744,N_4882);
or U7685 (N_7685,N_4979,N_4834);
and U7686 (N_7686,N_5066,N_5837);
and U7687 (N_7687,N_4452,N_5404);
or U7688 (N_7688,N_4040,N_4631);
and U7689 (N_7689,N_4179,N_4821);
xnor U7690 (N_7690,N_5179,N_5804);
nor U7691 (N_7691,N_4995,N_5450);
xor U7692 (N_7692,N_5555,N_4215);
nor U7693 (N_7693,N_5047,N_4062);
xor U7694 (N_7694,N_5749,N_5924);
xnor U7695 (N_7695,N_5142,N_4444);
or U7696 (N_7696,N_4513,N_4852);
nor U7697 (N_7697,N_5140,N_4053);
or U7698 (N_7698,N_5221,N_5024);
or U7699 (N_7699,N_4671,N_5827);
xor U7700 (N_7700,N_5505,N_5825);
nand U7701 (N_7701,N_4477,N_5302);
nand U7702 (N_7702,N_4010,N_4410);
nand U7703 (N_7703,N_4315,N_5136);
or U7704 (N_7704,N_4577,N_4450);
or U7705 (N_7705,N_5225,N_4578);
nor U7706 (N_7706,N_4531,N_4650);
or U7707 (N_7707,N_5196,N_5033);
xor U7708 (N_7708,N_5071,N_4655);
and U7709 (N_7709,N_5692,N_4659);
nor U7710 (N_7710,N_4325,N_4593);
and U7711 (N_7711,N_5576,N_4852);
nor U7712 (N_7712,N_4858,N_4087);
nand U7713 (N_7713,N_5863,N_5167);
nand U7714 (N_7714,N_4040,N_4471);
nand U7715 (N_7715,N_4482,N_4085);
or U7716 (N_7716,N_5897,N_5543);
nor U7717 (N_7717,N_4066,N_4204);
or U7718 (N_7718,N_4946,N_5548);
or U7719 (N_7719,N_4669,N_4785);
nand U7720 (N_7720,N_4482,N_5525);
xor U7721 (N_7721,N_4481,N_5646);
or U7722 (N_7722,N_4673,N_5099);
nor U7723 (N_7723,N_4444,N_4253);
nand U7724 (N_7724,N_4269,N_5630);
nor U7725 (N_7725,N_5827,N_5385);
nand U7726 (N_7726,N_5660,N_4784);
xnor U7727 (N_7727,N_5086,N_5616);
nor U7728 (N_7728,N_4437,N_5350);
or U7729 (N_7729,N_4598,N_5597);
xor U7730 (N_7730,N_5703,N_4685);
xnor U7731 (N_7731,N_5596,N_5859);
nand U7732 (N_7732,N_5680,N_4274);
and U7733 (N_7733,N_5877,N_5016);
nor U7734 (N_7734,N_4207,N_4661);
and U7735 (N_7735,N_4331,N_4589);
nand U7736 (N_7736,N_5523,N_4134);
or U7737 (N_7737,N_4054,N_4307);
nand U7738 (N_7738,N_5254,N_4896);
nor U7739 (N_7739,N_4170,N_4635);
or U7740 (N_7740,N_5760,N_5393);
or U7741 (N_7741,N_4438,N_5356);
or U7742 (N_7742,N_4122,N_4144);
xor U7743 (N_7743,N_5266,N_4786);
or U7744 (N_7744,N_5354,N_4684);
nor U7745 (N_7745,N_4618,N_4157);
and U7746 (N_7746,N_5532,N_5672);
and U7747 (N_7747,N_4492,N_5096);
and U7748 (N_7748,N_5047,N_5986);
nand U7749 (N_7749,N_4185,N_5618);
or U7750 (N_7750,N_5894,N_5439);
and U7751 (N_7751,N_5351,N_4610);
or U7752 (N_7752,N_5350,N_4759);
nor U7753 (N_7753,N_5899,N_5753);
nand U7754 (N_7754,N_5171,N_5218);
and U7755 (N_7755,N_4965,N_4762);
nand U7756 (N_7756,N_4624,N_5550);
xnor U7757 (N_7757,N_4431,N_4471);
and U7758 (N_7758,N_4338,N_5172);
nor U7759 (N_7759,N_4688,N_4391);
xnor U7760 (N_7760,N_5331,N_5997);
nor U7761 (N_7761,N_4616,N_5261);
xor U7762 (N_7762,N_5198,N_5412);
and U7763 (N_7763,N_4687,N_4781);
nand U7764 (N_7764,N_5038,N_4245);
xnor U7765 (N_7765,N_5990,N_4320);
nor U7766 (N_7766,N_4614,N_4521);
nor U7767 (N_7767,N_5881,N_4325);
nand U7768 (N_7768,N_5634,N_5239);
xor U7769 (N_7769,N_4401,N_5416);
xnor U7770 (N_7770,N_4661,N_5444);
and U7771 (N_7771,N_4583,N_4780);
nor U7772 (N_7772,N_5269,N_4192);
nor U7773 (N_7773,N_4126,N_5209);
nor U7774 (N_7774,N_5228,N_4512);
nand U7775 (N_7775,N_4840,N_4470);
xor U7776 (N_7776,N_5135,N_5145);
xor U7777 (N_7777,N_5284,N_4019);
nand U7778 (N_7778,N_5913,N_5728);
nor U7779 (N_7779,N_4584,N_5050);
xnor U7780 (N_7780,N_4796,N_4307);
xnor U7781 (N_7781,N_4939,N_4710);
nor U7782 (N_7782,N_4039,N_5512);
and U7783 (N_7783,N_4536,N_5674);
nor U7784 (N_7784,N_5870,N_4439);
or U7785 (N_7785,N_5993,N_4300);
and U7786 (N_7786,N_4264,N_4125);
and U7787 (N_7787,N_5103,N_5142);
or U7788 (N_7788,N_4683,N_5653);
xor U7789 (N_7789,N_4928,N_4320);
xnor U7790 (N_7790,N_4774,N_4170);
or U7791 (N_7791,N_5616,N_5258);
or U7792 (N_7792,N_5191,N_4302);
nand U7793 (N_7793,N_4012,N_5103);
nand U7794 (N_7794,N_5291,N_5567);
xnor U7795 (N_7795,N_5190,N_4523);
nor U7796 (N_7796,N_4407,N_5452);
nor U7797 (N_7797,N_5697,N_5437);
or U7798 (N_7798,N_5705,N_4636);
xnor U7799 (N_7799,N_4296,N_4598);
nand U7800 (N_7800,N_4105,N_5809);
nand U7801 (N_7801,N_5310,N_5874);
nand U7802 (N_7802,N_5464,N_4460);
and U7803 (N_7803,N_4323,N_4964);
and U7804 (N_7804,N_5375,N_4331);
and U7805 (N_7805,N_4768,N_4504);
xnor U7806 (N_7806,N_4470,N_4701);
or U7807 (N_7807,N_4742,N_5147);
and U7808 (N_7808,N_5162,N_4356);
xnor U7809 (N_7809,N_4842,N_4073);
xor U7810 (N_7810,N_4869,N_5459);
xnor U7811 (N_7811,N_4971,N_5799);
and U7812 (N_7812,N_4504,N_5801);
nand U7813 (N_7813,N_4698,N_4340);
nor U7814 (N_7814,N_4110,N_4833);
nor U7815 (N_7815,N_4261,N_5684);
and U7816 (N_7816,N_4612,N_5604);
or U7817 (N_7817,N_5342,N_4591);
and U7818 (N_7818,N_5011,N_5970);
and U7819 (N_7819,N_4751,N_4550);
and U7820 (N_7820,N_4093,N_4244);
nor U7821 (N_7821,N_5808,N_5409);
xor U7822 (N_7822,N_4084,N_5537);
or U7823 (N_7823,N_5106,N_5529);
or U7824 (N_7824,N_4724,N_5854);
nand U7825 (N_7825,N_4736,N_4549);
or U7826 (N_7826,N_4461,N_5039);
nand U7827 (N_7827,N_4709,N_4586);
or U7828 (N_7828,N_5753,N_5254);
nor U7829 (N_7829,N_4772,N_4885);
or U7830 (N_7830,N_4941,N_4118);
nand U7831 (N_7831,N_4426,N_4964);
or U7832 (N_7832,N_4518,N_4582);
or U7833 (N_7833,N_5979,N_5288);
or U7834 (N_7834,N_4704,N_4467);
nand U7835 (N_7835,N_4581,N_5258);
and U7836 (N_7836,N_4901,N_4526);
and U7837 (N_7837,N_5060,N_5580);
and U7838 (N_7838,N_5790,N_4415);
or U7839 (N_7839,N_5612,N_4091);
nand U7840 (N_7840,N_5187,N_4794);
nand U7841 (N_7841,N_5150,N_5791);
or U7842 (N_7842,N_5401,N_5480);
nor U7843 (N_7843,N_4676,N_5003);
and U7844 (N_7844,N_4267,N_5967);
nand U7845 (N_7845,N_4208,N_4146);
nand U7846 (N_7846,N_5909,N_5373);
xor U7847 (N_7847,N_5392,N_5725);
xor U7848 (N_7848,N_5903,N_5114);
and U7849 (N_7849,N_4260,N_5739);
and U7850 (N_7850,N_4544,N_4385);
nor U7851 (N_7851,N_5819,N_4925);
xor U7852 (N_7852,N_5865,N_4077);
and U7853 (N_7853,N_5165,N_4189);
nand U7854 (N_7854,N_5925,N_4538);
or U7855 (N_7855,N_5038,N_5507);
and U7856 (N_7856,N_4626,N_4838);
nand U7857 (N_7857,N_5229,N_4896);
or U7858 (N_7858,N_5941,N_4294);
nor U7859 (N_7859,N_5007,N_5601);
nor U7860 (N_7860,N_4388,N_4973);
and U7861 (N_7861,N_4841,N_4489);
and U7862 (N_7862,N_5354,N_5577);
and U7863 (N_7863,N_5443,N_4690);
xnor U7864 (N_7864,N_5813,N_5829);
nor U7865 (N_7865,N_4405,N_5679);
nand U7866 (N_7866,N_5674,N_4078);
xnor U7867 (N_7867,N_4628,N_5291);
nand U7868 (N_7868,N_5787,N_4644);
and U7869 (N_7869,N_5047,N_5247);
xnor U7870 (N_7870,N_5883,N_5011);
xnor U7871 (N_7871,N_4282,N_4956);
nor U7872 (N_7872,N_4853,N_5964);
nand U7873 (N_7873,N_4933,N_4940);
or U7874 (N_7874,N_5784,N_5067);
nand U7875 (N_7875,N_5468,N_4802);
or U7876 (N_7876,N_4220,N_5342);
or U7877 (N_7877,N_4509,N_4376);
nor U7878 (N_7878,N_4495,N_4228);
nor U7879 (N_7879,N_4642,N_5917);
xor U7880 (N_7880,N_4725,N_5273);
or U7881 (N_7881,N_5854,N_5028);
or U7882 (N_7882,N_5097,N_4463);
or U7883 (N_7883,N_4736,N_5044);
nor U7884 (N_7884,N_4082,N_4095);
xnor U7885 (N_7885,N_5142,N_4009);
nor U7886 (N_7886,N_4415,N_5138);
nand U7887 (N_7887,N_5143,N_4321);
nand U7888 (N_7888,N_5719,N_4861);
or U7889 (N_7889,N_5148,N_4886);
nand U7890 (N_7890,N_4479,N_4995);
or U7891 (N_7891,N_4712,N_5351);
nor U7892 (N_7892,N_4050,N_4584);
and U7893 (N_7893,N_4756,N_4171);
or U7894 (N_7894,N_4878,N_5316);
nor U7895 (N_7895,N_5411,N_5173);
nand U7896 (N_7896,N_5315,N_5590);
nor U7897 (N_7897,N_5184,N_4161);
or U7898 (N_7898,N_5758,N_5140);
or U7899 (N_7899,N_4499,N_5640);
and U7900 (N_7900,N_5772,N_4111);
xnor U7901 (N_7901,N_4617,N_5238);
and U7902 (N_7902,N_4586,N_4069);
nand U7903 (N_7903,N_4821,N_4460);
xor U7904 (N_7904,N_5269,N_4443);
nor U7905 (N_7905,N_5525,N_5138);
nand U7906 (N_7906,N_5873,N_5678);
or U7907 (N_7907,N_5989,N_5777);
nand U7908 (N_7908,N_4521,N_4625);
nand U7909 (N_7909,N_5639,N_4380);
nor U7910 (N_7910,N_4558,N_5753);
and U7911 (N_7911,N_4843,N_4365);
nand U7912 (N_7912,N_5253,N_5399);
or U7913 (N_7913,N_5195,N_4625);
xnor U7914 (N_7914,N_4652,N_5976);
nand U7915 (N_7915,N_5058,N_5237);
nor U7916 (N_7916,N_4872,N_4321);
or U7917 (N_7917,N_5991,N_5215);
nor U7918 (N_7918,N_4154,N_4561);
or U7919 (N_7919,N_4184,N_4465);
nor U7920 (N_7920,N_4666,N_4415);
nand U7921 (N_7921,N_4874,N_4693);
and U7922 (N_7922,N_5491,N_5781);
xnor U7923 (N_7923,N_5084,N_4665);
nor U7924 (N_7924,N_4988,N_4665);
nor U7925 (N_7925,N_5411,N_4153);
and U7926 (N_7926,N_4876,N_5181);
xor U7927 (N_7927,N_5670,N_5483);
and U7928 (N_7928,N_5846,N_5600);
nand U7929 (N_7929,N_5373,N_5212);
and U7930 (N_7930,N_4544,N_4554);
nand U7931 (N_7931,N_5683,N_4307);
nand U7932 (N_7932,N_4116,N_5259);
and U7933 (N_7933,N_4444,N_4341);
or U7934 (N_7934,N_5724,N_5056);
xor U7935 (N_7935,N_5855,N_4709);
nand U7936 (N_7936,N_5673,N_5756);
xnor U7937 (N_7937,N_5085,N_4357);
or U7938 (N_7938,N_4182,N_5092);
and U7939 (N_7939,N_4305,N_5928);
nand U7940 (N_7940,N_4015,N_4852);
nand U7941 (N_7941,N_4811,N_5116);
nor U7942 (N_7942,N_5632,N_5668);
nand U7943 (N_7943,N_5253,N_4475);
or U7944 (N_7944,N_4142,N_5745);
xnor U7945 (N_7945,N_4472,N_4853);
or U7946 (N_7946,N_4195,N_5553);
or U7947 (N_7947,N_5994,N_4755);
and U7948 (N_7948,N_4415,N_5438);
nor U7949 (N_7949,N_5759,N_5804);
and U7950 (N_7950,N_5169,N_4629);
and U7951 (N_7951,N_5480,N_4673);
nor U7952 (N_7952,N_4951,N_4071);
xor U7953 (N_7953,N_4574,N_4550);
nand U7954 (N_7954,N_4529,N_4692);
nand U7955 (N_7955,N_5904,N_5600);
and U7956 (N_7956,N_5332,N_4026);
nor U7957 (N_7957,N_4816,N_5324);
or U7958 (N_7958,N_5758,N_4784);
nor U7959 (N_7959,N_5298,N_4714);
nor U7960 (N_7960,N_5844,N_5415);
xor U7961 (N_7961,N_4803,N_4855);
nor U7962 (N_7962,N_5631,N_4058);
or U7963 (N_7963,N_5362,N_5958);
nand U7964 (N_7964,N_5595,N_4043);
or U7965 (N_7965,N_5744,N_4086);
xor U7966 (N_7966,N_5809,N_4401);
and U7967 (N_7967,N_4531,N_5539);
nand U7968 (N_7968,N_4145,N_4776);
xor U7969 (N_7969,N_4570,N_5783);
or U7970 (N_7970,N_5098,N_5962);
or U7971 (N_7971,N_4093,N_4151);
nand U7972 (N_7972,N_4693,N_4379);
nand U7973 (N_7973,N_4051,N_5521);
xor U7974 (N_7974,N_5649,N_5327);
or U7975 (N_7975,N_4114,N_4790);
nor U7976 (N_7976,N_5042,N_4715);
nand U7977 (N_7977,N_4579,N_5056);
and U7978 (N_7978,N_5917,N_5451);
nor U7979 (N_7979,N_5490,N_5642);
or U7980 (N_7980,N_5679,N_4257);
nand U7981 (N_7981,N_4176,N_4040);
nor U7982 (N_7982,N_4767,N_5092);
nand U7983 (N_7983,N_5411,N_4258);
nor U7984 (N_7984,N_4493,N_4204);
nor U7985 (N_7985,N_5602,N_4496);
or U7986 (N_7986,N_4996,N_5881);
nor U7987 (N_7987,N_4122,N_4974);
or U7988 (N_7988,N_5093,N_5539);
and U7989 (N_7989,N_4345,N_5727);
nand U7990 (N_7990,N_5081,N_5828);
nand U7991 (N_7991,N_4511,N_5628);
or U7992 (N_7992,N_4137,N_5701);
and U7993 (N_7993,N_4710,N_4623);
and U7994 (N_7994,N_5315,N_5621);
xor U7995 (N_7995,N_5398,N_5546);
nor U7996 (N_7996,N_4771,N_4255);
nor U7997 (N_7997,N_5289,N_5985);
and U7998 (N_7998,N_5281,N_4140);
and U7999 (N_7999,N_5836,N_5635);
xnor U8000 (N_8000,N_7385,N_6579);
nand U8001 (N_8001,N_6912,N_6176);
and U8002 (N_8002,N_6459,N_6142);
xnor U8003 (N_8003,N_7795,N_6636);
xnor U8004 (N_8004,N_6928,N_7745);
xnor U8005 (N_8005,N_7964,N_6240);
nor U8006 (N_8006,N_6923,N_6591);
and U8007 (N_8007,N_7320,N_7792);
or U8008 (N_8008,N_7999,N_6587);
and U8009 (N_8009,N_7846,N_7835);
xor U8010 (N_8010,N_6227,N_7755);
nand U8011 (N_8011,N_7315,N_6327);
nand U8012 (N_8012,N_7145,N_7699);
nor U8013 (N_8013,N_7251,N_7491);
xnor U8014 (N_8014,N_7129,N_7033);
nor U8015 (N_8015,N_7370,N_6652);
nor U8016 (N_8016,N_7574,N_7741);
xnor U8017 (N_8017,N_6976,N_7006);
or U8018 (N_8018,N_7071,N_6601);
and U8019 (N_8019,N_6299,N_7485);
and U8020 (N_8020,N_7488,N_6233);
and U8021 (N_8021,N_7627,N_6461);
nor U8022 (N_8022,N_7509,N_7447);
nand U8023 (N_8023,N_6085,N_7598);
or U8024 (N_8024,N_7368,N_6692);
nand U8025 (N_8025,N_6651,N_7088);
or U8026 (N_8026,N_7146,N_7990);
nand U8027 (N_8027,N_7101,N_6607);
nand U8028 (N_8028,N_6274,N_6703);
nor U8029 (N_8029,N_7702,N_6048);
xnor U8030 (N_8030,N_7352,N_7142);
and U8031 (N_8031,N_7606,N_6191);
and U8032 (N_8032,N_6401,N_6500);
or U8033 (N_8033,N_6387,N_6945);
or U8034 (N_8034,N_6472,N_7260);
and U8035 (N_8035,N_6850,N_7675);
xor U8036 (N_8036,N_7160,N_6517);
xnor U8037 (N_8037,N_6983,N_6049);
nand U8038 (N_8038,N_6203,N_6292);
xor U8039 (N_8039,N_6244,N_6257);
or U8040 (N_8040,N_6483,N_7858);
or U8041 (N_8041,N_6509,N_6538);
xnor U8042 (N_8042,N_7821,N_7684);
or U8043 (N_8043,N_6305,N_6934);
nand U8044 (N_8044,N_6816,N_6979);
or U8045 (N_8045,N_6139,N_6273);
or U8046 (N_8046,N_6756,N_7378);
xor U8047 (N_8047,N_6732,N_6072);
or U8048 (N_8048,N_6688,N_7324);
xor U8049 (N_8049,N_7109,N_6524);
nor U8050 (N_8050,N_7850,N_6914);
and U8051 (N_8051,N_6569,N_7461);
or U8052 (N_8052,N_7716,N_7818);
nand U8053 (N_8053,N_7736,N_6880);
or U8054 (N_8054,N_6857,N_6539);
nor U8055 (N_8055,N_6130,N_7625);
or U8056 (N_8056,N_7697,N_6451);
or U8057 (N_8057,N_6728,N_7624);
and U8058 (N_8058,N_6553,N_7894);
and U8059 (N_8059,N_6121,N_6836);
xor U8060 (N_8060,N_6403,N_7587);
xnor U8061 (N_8061,N_6852,N_6389);
and U8062 (N_8062,N_6175,N_7877);
or U8063 (N_8063,N_7300,N_7424);
nand U8064 (N_8064,N_6138,N_6847);
and U8065 (N_8065,N_7876,N_7597);
or U8066 (N_8066,N_7502,N_6448);
and U8067 (N_8067,N_7758,N_6061);
or U8068 (N_8068,N_7555,N_7490);
nand U8069 (N_8069,N_7452,N_6382);
xnor U8070 (N_8070,N_7449,N_7861);
or U8071 (N_8071,N_6496,N_7576);
or U8072 (N_8072,N_6102,N_7690);
or U8073 (N_8073,N_7000,N_6047);
nor U8074 (N_8074,N_6222,N_6748);
nor U8075 (N_8075,N_7074,N_7134);
nor U8076 (N_8076,N_6063,N_7395);
nor U8077 (N_8077,N_6626,N_6859);
and U8078 (N_8078,N_7373,N_7920);
or U8079 (N_8079,N_7241,N_6742);
and U8080 (N_8080,N_7568,N_6650);
xor U8081 (N_8081,N_7562,N_7037);
nor U8082 (N_8082,N_6937,N_7215);
nor U8083 (N_8083,N_6902,N_7362);
xnor U8084 (N_8084,N_6842,N_7467);
and U8085 (N_8085,N_6760,N_7454);
xor U8086 (N_8086,N_7356,N_6287);
and U8087 (N_8087,N_6915,N_7805);
and U8088 (N_8088,N_7259,N_6137);
nand U8089 (N_8089,N_6128,N_7904);
or U8090 (N_8090,N_6491,N_6667);
xor U8091 (N_8091,N_7418,N_7830);
nand U8092 (N_8092,N_6062,N_7249);
and U8093 (N_8093,N_6236,N_6625);
or U8094 (N_8094,N_6179,N_6910);
and U8095 (N_8095,N_6457,N_7772);
xor U8096 (N_8096,N_6884,N_7180);
xor U8097 (N_8097,N_6653,N_7820);
nand U8098 (N_8098,N_7198,N_7910);
nor U8099 (N_8099,N_6473,N_7847);
and U8100 (N_8100,N_7206,N_6963);
nor U8101 (N_8101,N_7285,N_7159);
nand U8102 (N_8102,N_6961,N_7984);
xnor U8103 (N_8103,N_6495,N_6219);
nand U8104 (N_8104,N_7882,N_6676);
nand U8105 (N_8105,N_7204,N_6761);
or U8106 (N_8106,N_6886,N_6665);
xor U8107 (N_8107,N_7515,N_7903);
xnor U8108 (N_8108,N_6835,N_6487);
nor U8109 (N_8109,N_7347,N_7610);
xor U8110 (N_8110,N_6317,N_6259);
nor U8111 (N_8111,N_7427,N_7538);
xor U8112 (N_8112,N_6091,N_6116);
nor U8113 (N_8113,N_6250,N_7960);
nor U8114 (N_8114,N_7689,N_7926);
nor U8115 (N_8115,N_7421,N_7015);
nand U8116 (N_8116,N_6547,N_7305);
and U8117 (N_8117,N_7087,N_6699);
or U8118 (N_8118,N_6907,N_7070);
nor U8119 (N_8119,N_7027,N_6195);
or U8120 (N_8120,N_7464,N_6036);
xor U8121 (N_8121,N_6925,N_7954);
nor U8122 (N_8122,N_6573,N_7616);
and U8123 (N_8123,N_6367,N_6194);
and U8124 (N_8124,N_6360,N_7388);
nor U8125 (N_8125,N_7500,N_7340);
nand U8126 (N_8126,N_6391,N_6368);
xnor U8127 (N_8127,N_7687,N_7104);
nand U8128 (N_8128,N_7256,N_7677);
and U8129 (N_8129,N_6935,N_6682);
or U8130 (N_8130,N_6460,N_6098);
or U8131 (N_8131,N_7542,N_7536);
or U8132 (N_8132,N_6431,N_6225);
and U8133 (N_8133,N_7793,N_6507);
and U8134 (N_8134,N_7942,N_6975);
and U8135 (N_8135,N_6437,N_7865);
nor U8136 (N_8136,N_6637,N_7836);
xor U8137 (N_8137,N_7871,N_7510);
and U8138 (N_8138,N_7873,N_7596);
xor U8139 (N_8139,N_6300,N_6870);
nand U8140 (N_8140,N_7039,N_7539);
xor U8141 (N_8141,N_6335,N_7453);
xor U8142 (N_8142,N_6463,N_7280);
or U8143 (N_8143,N_6046,N_7875);
and U8144 (N_8144,N_6697,N_6891);
and U8145 (N_8145,N_6738,N_6634);
or U8146 (N_8146,N_6785,N_6231);
xnor U8147 (N_8147,N_6234,N_7952);
xnor U8148 (N_8148,N_6719,N_7763);
nor U8149 (N_8149,N_7497,N_6316);
xnor U8150 (N_8150,N_7918,N_6205);
nand U8151 (N_8151,N_7679,N_6044);
nand U8152 (N_8152,N_7375,N_7473);
or U8153 (N_8153,N_7535,N_6811);
xnor U8154 (N_8154,N_7270,N_7383);
nor U8155 (N_8155,N_6566,N_7484);
or U8156 (N_8156,N_6708,N_7522);
nand U8157 (N_8157,N_7399,N_6729);
or U8158 (N_8158,N_6221,N_7499);
or U8159 (N_8159,N_6117,N_7199);
xnor U8160 (N_8160,N_7566,N_6603);
nand U8161 (N_8161,N_7807,N_6763);
or U8162 (N_8162,N_6799,N_7468);
xnor U8163 (N_8163,N_7872,N_7661);
xor U8164 (N_8164,N_6548,N_6088);
or U8165 (N_8165,N_7730,N_7672);
xnor U8166 (N_8166,N_7479,N_6320);
and U8167 (N_8167,N_7959,N_7612);
or U8168 (N_8168,N_7989,N_6475);
and U8169 (N_8169,N_7770,N_7781);
and U8170 (N_8170,N_6235,N_6647);
or U8171 (N_8171,N_7981,N_7263);
xor U8172 (N_8172,N_7660,N_6141);
nor U8173 (N_8173,N_6351,N_6201);
nor U8174 (N_8174,N_6642,N_6192);
or U8175 (N_8175,N_6356,N_6693);
nand U8176 (N_8176,N_6096,N_7239);
or U8177 (N_8177,N_6679,N_7042);
or U8178 (N_8178,N_7859,N_7084);
nor U8179 (N_8179,N_7308,N_6947);
xor U8180 (N_8180,N_6997,N_7787);
nand U8181 (N_8181,N_7040,N_7120);
or U8182 (N_8182,N_6602,N_7254);
nor U8183 (N_8183,N_7889,N_6442);
xor U8184 (N_8184,N_6084,N_7611);
nor U8185 (N_8185,N_7851,N_7291);
and U8186 (N_8186,N_6791,N_7666);
xnor U8187 (N_8187,N_6977,N_7316);
nor U8188 (N_8188,N_6993,N_6256);
nor U8189 (N_8189,N_7780,N_7968);
nand U8190 (N_8190,N_7090,N_6798);
nand U8191 (N_8191,N_6707,N_7934);
and U8192 (N_8192,N_6624,N_7132);
xor U8193 (N_8193,N_6359,N_6207);
nor U8194 (N_8194,N_7809,N_6466);
nand U8195 (N_8195,N_7890,N_7481);
xor U8196 (N_8196,N_6804,N_6563);
or U8197 (N_8197,N_7366,N_7585);
nor U8198 (N_8198,N_6125,N_6726);
nand U8199 (N_8199,N_6599,N_7718);
or U8200 (N_8200,N_6932,N_7131);
xor U8201 (N_8201,N_7925,N_7174);
nand U8202 (N_8202,N_7061,N_7543);
nor U8203 (N_8203,N_6497,N_6794);
and U8204 (N_8204,N_6375,N_6861);
and U8205 (N_8205,N_7860,N_6436);
nor U8206 (N_8206,N_7838,N_7746);
nand U8207 (N_8207,N_6833,N_6812);
nand U8208 (N_8208,N_7629,N_7317);
nor U8209 (N_8209,N_7546,N_7083);
xor U8210 (N_8210,N_7067,N_6904);
xor U8211 (N_8211,N_7028,N_7767);
or U8212 (N_8212,N_6095,N_7319);
and U8213 (N_8213,N_6527,N_7682);
xor U8214 (N_8214,N_7032,N_7874);
and U8215 (N_8215,N_6110,N_7178);
xor U8216 (N_8216,N_6357,N_6263);
and U8217 (N_8217,N_7958,N_6004);
xor U8218 (N_8218,N_7163,N_7525);
nor U8219 (N_8219,N_7387,N_7152);
and U8220 (N_8220,N_6877,N_6477);
nor U8221 (N_8221,N_7678,N_7220);
xnor U8222 (N_8222,N_6045,N_7505);
nand U8223 (N_8223,N_6752,N_7680);
nand U8224 (N_8224,N_6696,N_7808);
or U8225 (N_8225,N_6186,N_7100);
xor U8226 (N_8226,N_6988,N_6433);
xnor U8227 (N_8227,N_7092,N_7631);
and U8228 (N_8228,N_7734,N_7407);
nor U8229 (N_8229,N_6890,N_6751);
nand U8230 (N_8230,N_7267,N_6950);
nor U8231 (N_8231,N_7712,N_7940);
nand U8232 (N_8232,N_6585,N_7065);
nand U8233 (N_8233,N_6447,N_7128);
nand U8234 (N_8234,N_7466,N_6388);
nor U8235 (N_8235,N_7516,N_6879);
xor U8236 (N_8236,N_7228,N_7203);
nor U8237 (N_8237,N_6765,N_7759);
and U8238 (N_8238,N_6103,N_7089);
and U8239 (N_8239,N_6485,N_7891);
or U8240 (N_8240,N_6805,N_6020);
and U8241 (N_8241,N_7521,N_7333);
nand U8242 (N_8242,N_6577,N_6899);
or U8243 (N_8243,N_6611,N_6378);
nand U8244 (N_8244,N_7112,N_6820);
nand U8245 (N_8245,N_6887,N_6572);
and U8246 (N_8246,N_7898,N_6536);
nor U8247 (N_8247,N_6479,N_6501);
and U8248 (N_8248,N_7377,N_6689);
and U8249 (N_8249,N_6018,N_7641);
xor U8250 (N_8250,N_6269,N_7642);
nor U8251 (N_8251,N_6126,N_7289);
or U8252 (N_8252,N_6795,N_6167);
nor U8253 (N_8253,N_6092,N_7097);
or U8254 (N_8254,N_6339,N_6373);
and U8255 (N_8255,N_7334,N_7093);
and U8256 (N_8256,N_7049,N_6954);
and U8257 (N_8257,N_6754,N_6808);
and U8258 (N_8258,N_7652,N_7185);
nand U8259 (N_8259,N_7309,N_7966);
and U8260 (N_8260,N_6258,N_7571);
xor U8261 (N_8261,N_7840,N_7116);
and U8262 (N_8262,N_7495,N_6193);
xor U8263 (N_8263,N_6055,N_6372);
xor U8264 (N_8264,N_6106,N_7913);
xnor U8265 (N_8265,N_7676,N_6464);
or U8266 (N_8266,N_7111,N_7279);
xor U8267 (N_8267,N_6776,N_7242);
and U8268 (N_8268,N_6333,N_7945);
or U8269 (N_8269,N_7457,N_7837);
nand U8270 (N_8270,N_6255,N_7800);
and U8271 (N_8271,N_7888,N_7615);
nand U8272 (N_8272,N_6271,N_6054);
nand U8273 (N_8273,N_7965,N_7983);
and U8274 (N_8274,N_6680,N_7237);
nor U8275 (N_8275,N_6797,N_7341);
nand U8276 (N_8276,N_7550,N_6559);
and U8277 (N_8277,N_6281,N_7721);
nand U8278 (N_8278,N_7414,N_6040);
xnor U8279 (N_8279,N_7613,N_7951);
nand U8280 (N_8280,N_7361,N_7292);
or U8281 (N_8281,N_7115,N_7321);
nor U8282 (N_8282,N_7095,N_6122);
nand U8283 (N_8283,N_6198,N_6541);
nand U8284 (N_8284,N_7498,N_7036);
nand U8285 (N_8285,N_6493,N_6987);
nand U8286 (N_8286,N_6077,N_6484);
or U8287 (N_8287,N_7094,N_7899);
or U8288 (N_8288,N_6635,N_7238);
nand U8289 (N_8289,N_7524,N_6218);
or U8290 (N_8290,N_6957,N_7148);
and U8291 (N_8291,N_7360,N_6152);
xor U8292 (N_8292,N_7663,N_7790);
xor U8293 (N_8293,N_7496,N_7953);
nor U8294 (N_8294,N_7085,N_7552);
or U8295 (N_8295,N_6581,N_6383);
nand U8296 (N_8296,N_6921,N_6051);
nand U8297 (N_8297,N_6502,N_6104);
xor U8298 (N_8298,N_7181,N_7798);
nor U8299 (N_8299,N_7191,N_6809);
xor U8300 (N_8300,N_6516,N_6734);
nor U8301 (N_8301,N_6788,N_6350);
nand U8302 (N_8302,N_6731,N_7038);
or U8303 (N_8303,N_6003,N_6366);
nand U8304 (N_8304,N_7886,N_6303);
nor U8305 (N_8305,N_7372,N_7114);
xor U8306 (N_8306,N_6017,N_7478);
xor U8307 (N_8307,N_7063,N_6951);
and U8308 (N_8308,N_6016,N_6955);
and U8309 (N_8309,N_6028,N_6562);
or U8310 (N_8310,N_6124,N_7353);
and U8311 (N_8311,N_7076,N_6414);
nor U8312 (N_8312,N_7578,N_7150);
and U8313 (N_8313,N_7591,N_6489);
nor U8314 (N_8314,N_6528,N_7350);
nor U8315 (N_8315,N_6906,N_6223);
or U8316 (N_8316,N_6858,N_6649);
xnor U8317 (N_8317,N_7136,N_7137);
xor U8318 (N_8318,N_7863,N_7864);
or U8319 (N_8319,N_6329,N_7342);
nor U8320 (N_8320,N_7030,N_7824);
xnor U8321 (N_8321,N_6659,N_6456);
nand U8322 (N_8322,N_6832,N_6163);
or U8323 (N_8323,N_6232,N_7540);
xor U8324 (N_8324,N_6086,N_6006);
nand U8325 (N_8325,N_7769,N_7554);
nand U8326 (N_8326,N_7583,N_7003);
nand U8327 (N_8327,N_7056,N_6400);
nor U8328 (N_8328,N_7575,N_7367);
or U8329 (N_8329,N_7218,N_7658);
or U8330 (N_8330,N_7963,N_6593);
nor U8331 (N_8331,N_7494,N_7102);
and U8332 (N_8332,N_6943,N_7557);
and U8333 (N_8333,N_7825,N_6408);
xnor U8334 (N_8334,N_7726,N_6025);
xnor U8335 (N_8335,N_6019,N_7662);
and U8336 (N_8336,N_7590,N_7079);
nand U8337 (N_8337,N_6766,N_7420);
xor U8338 (N_8338,N_6770,N_7135);
xnor U8339 (N_8339,N_6342,N_6655);
or U8340 (N_8340,N_7523,N_6087);
xnor U8341 (N_8341,N_7429,N_7595);
xor U8342 (N_8342,N_7507,N_6404);
and U8343 (N_8343,N_7197,N_7644);
or U8344 (N_8344,N_6348,N_7747);
nand U8345 (N_8345,N_6038,N_6272);
xnor U8346 (N_8346,N_7879,N_6518);
nand U8347 (N_8347,N_7106,N_6444);
and U8348 (N_8348,N_7533,N_6841);
and U8349 (N_8349,N_7573,N_6545);
and U8350 (N_8350,N_6780,N_7073);
nand U8351 (N_8351,N_7527,N_6161);
nand U8352 (N_8352,N_6249,N_6380);
or U8353 (N_8353,N_6468,N_6825);
nor U8354 (N_8354,N_6893,N_6159);
nand U8355 (N_8355,N_7584,N_6041);
and U8356 (N_8356,N_7916,N_6515);
and U8357 (N_8357,N_7856,N_6453);
xnor U8358 (N_8358,N_6677,N_6114);
nand U8359 (N_8359,N_6714,N_7618);
and U8360 (N_8360,N_7608,N_6481);
xor U8361 (N_8361,N_6177,N_7412);
nand U8362 (N_8362,N_6113,N_6758);
nor U8363 (N_8363,N_7783,N_6009);
or U8364 (N_8364,N_7564,N_6172);
xor U8365 (N_8365,N_7113,N_6133);
nand U8366 (N_8366,N_6962,N_6864);
and U8367 (N_8367,N_6815,N_7950);
and U8368 (N_8368,N_6827,N_7202);
xnor U8369 (N_8369,N_7096,N_6352);
and U8370 (N_8370,N_6648,N_6080);
xnor U8371 (N_8371,N_6343,N_7068);
nand U8372 (N_8372,N_7365,N_6793);
nand U8373 (N_8373,N_7915,N_7883);
nand U8374 (N_8374,N_6662,N_7572);
nand U8375 (N_8375,N_7988,N_6071);
nand U8376 (N_8376,N_7293,N_6349);
nor U8377 (N_8377,N_6911,N_6094);
xnor U8378 (N_8378,N_6100,N_7435);
nand U8379 (N_8379,N_7985,N_7928);
xor U8380 (N_8380,N_6237,N_7169);
or U8381 (N_8381,N_6056,N_7209);
and U8382 (N_8382,N_6318,N_7230);
or U8383 (N_8383,N_6168,N_6023);
or U8384 (N_8384,N_6561,N_7433);
xor U8385 (N_8385,N_7144,N_6633);
and U8386 (N_8386,N_7029,N_6315);
xor U8387 (N_8387,N_6535,N_7483);
or U8388 (N_8388,N_7696,N_6715);
or U8389 (N_8389,N_6313,N_6187);
xor U8390 (N_8390,N_7140,N_7002);
and U8391 (N_8391,N_6613,N_7299);
nor U8392 (N_8392,N_6956,N_6504);
nor U8393 (N_8393,N_6260,N_7796);
xnor U8394 (N_8394,N_7034,N_7601);
and U8395 (N_8395,N_6730,N_7107);
nand U8396 (N_8396,N_6544,N_7994);
and U8397 (N_8397,N_7219,N_6522);
and U8398 (N_8398,N_6610,N_7402);
or U8399 (N_8399,N_7518,N_6423);
nand U8400 (N_8400,N_7729,N_7843);
nand U8401 (N_8401,N_7806,N_7386);
or U8402 (N_8402,N_6644,N_7422);
or U8403 (N_8403,N_7560,N_6638);
nand U8404 (N_8404,N_7804,N_6540);
and U8405 (N_8405,N_6922,N_7171);
nor U8406 (N_8406,N_6369,N_6334);
nand U8407 (N_8407,N_6658,N_7588);
nor U8408 (N_8408,N_7991,N_7921);
and U8409 (N_8409,N_6694,N_6845);
xor U8410 (N_8410,N_7638,N_6716);
or U8411 (N_8411,N_6067,N_6171);
xor U8412 (N_8412,N_6823,N_6576);
or U8413 (N_8413,N_6739,N_7593);
nand U8414 (N_8414,N_7244,N_7448);
or U8415 (N_8415,N_7789,N_7531);
or U8416 (N_8416,N_6482,N_6075);
or U8417 (N_8417,N_7857,N_6546);
or U8418 (N_8418,N_7363,N_7351);
nand U8419 (N_8419,N_6874,N_6446);
or U8420 (N_8420,N_7844,N_6755);
nand U8421 (N_8421,N_7487,N_6412);
and U8422 (N_8422,N_6362,N_7648);
xor U8423 (N_8423,N_7426,N_6953);
nand U8424 (N_8424,N_7348,N_6458);
or U8425 (N_8425,N_7240,N_7226);
and U8426 (N_8426,N_7046,N_6737);
or U8427 (N_8427,N_7938,N_7175);
xor U8428 (N_8428,N_6654,N_7737);
nor U8429 (N_8429,N_7381,N_7719);
and U8430 (N_8430,N_6838,N_6268);
and U8431 (N_8431,N_6079,N_7176);
and U8432 (N_8432,N_6894,N_6147);
nor U8433 (N_8433,N_6415,N_7937);
and U8434 (N_8434,N_7650,N_6490);
nand U8435 (N_8435,N_7547,N_7900);
xor U8436 (N_8436,N_7231,N_6557);
xnor U8437 (N_8437,N_6821,N_6691);
or U8438 (N_8438,N_7799,N_6407);
or U8439 (N_8439,N_6499,N_6355);
xor U8440 (N_8440,N_7567,N_6465);
nor U8441 (N_8441,N_6849,N_6514);
xnor U8442 (N_8442,N_6558,N_6723);
nand U8443 (N_8443,N_6032,N_6439);
nor U8444 (N_8444,N_6285,N_7924);
xnor U8445 (N_8445,N_7337,N_6973);
nor U8446 (N_8446,N_6631,N_7753);
or U8447 (N_8447,N_6488,N_7275);
nand U8448 (N_8448,N_6550,N_6420);
and U8449 (N_8449,N_6289,N_6592);
nand U8450 (N_8450,N_6377,N_6687);
or U8451 (N_8451,N_7025,N_6252);
nand U8452 (N_8452,N_6918,N_7556);
xnor U8453 (N_8453,N_7559,N_7674);
or U8454 (N_8454,N_6209,N_6867);
and U8455 (N_8455,N_6965,N_7413);
and U8456 (N_8456,N_6826,N_6740);
xnor U8457 (N_8457,N_7450,N_7724);
xor U8458 (N_8458,N_7506,N_7651);
or U8459 (N_8459,N_7742,N_7892);
xnor U8460 (N_8460,N_7801,N_7480);
nor U8461 (N_8461,N_7408,N_7819);
and U8462 (N_8462,N_6053,N_7290);
xor U8463 (N_8463,N_6014,N_6609);
nor U8464 (N_8464,N_6646,N_7053);
and U8465 (N_8465,N_7147,N_6083);
nor U8466 (N_8466,N_7743,N_6469);
or U8467 (N_8467,N_7878,N_7996);
nor U8468 (N_8468,N_7234,N_7946);
xor U8469 (N_8469,N_7417,N_7081);
or U8470 (N_8470,N_6486,N_7776);
nor U8471 (N_8471,N_6082,N_6917);
nor U8472 (N_8472,N_7165,N_7155);
or U8473 (N_8473,N_6747,N_6630);
nor U8474 (N_8474,N_7232,N_7961);
nor U8475 (N_8475,N_6948,N_6185);
xor U8476 (N_8476,N_6284,N_7561);
nor U8477 (N_8477,N_7586,N_6628);
xnor U8478 (N_8478,N_7327,N_6265);
nand U8479 (N_8479,N_6969,N_6115);
or U8480 (N_8480,N_7229,N_6429);
nor U8481 (N_8481,N_7437,N_6266);
or U8482 (N_8482,N_6267,N_6551);
nor U8483 (N_8483,N_6312,N_6381);
and U8484 (N_8484,N_6021,N_6898);
xor U8485 (N_8485,N_6744,N_6024);
nor U8486 (N_8486,N_7287,N_7194);
nor U8487 (N_8487,N_7243,N_6081);
xnor U8488 (N_8488,N_6574,N_7045);
or U8489 (N_8489,N_6015,N_7168);
or U8490 (N_8490,N_7108,N_6930);
or U8491 (N_8491,N_6671,N_7649);
and U8492 (N_8492,N_7706,N_7286);
nand U8493 (N_8493,N_7887,N_7941);
nand U8494 (N_8494,N_6011,N_6604);
or U8495 (N_8495,N_7183,N_7848);
nor U8496 (N_8496,N_6787,N_6183);
nand U8497 (N_8497,N_6768,N_6735);
and U8498 (N_8498,N_6230,N_6419);
and U8499 (N_8499,N_6526,N_6190);
nand U8500 (N_8500,N_7276,N_6330);
nor U8501 (N_8501,N_6674,N_7592);
nand U8502 (N_8502,N_6759,N_7326);
nor U8503 (N_8503,N_7973,N_6627);
or U8504 (N_8504,N_7482,N_6480);
xnor U8505 (N_8505,N_7072,N_6717);
or U8506 (N_8506,N_6556,N_7732);
nand U8507 (N_8507,N_7359,N_6498);
nor U8508 (N_8508,N_6332,N_7475);
xor U8509 (N_8509,N_6984,N_6309);
and U8510 (N_8510,N_6402,N_7725);
xnor U8511 (N_8511,N_7978,N_6673);
xnor U8512 (N_8512,N_6008,N_6718);
nor U8513 (N_8513,N_7405,N_6941);
nand U8514 (N_8514,N_7126,N_7817);
nor U8515 (N_8515,N_7423,N_6512);
or U8516 (N_8516,N_6282,N_7250);
nor U8517 (N_8517,N_7224,N_6803);
nand U8518 (N_8518,N_7162,N_6749);
and U8519 (N_8519,N_7749,N_7050);
nand U8520 (N_8520,N_6396,N_7007);
xor U8521 (N_8521,N_7031,N_6279);
xor U8522 (N_8522,N_7274,N_6421);
or U8523 (N_8523,N_6363,N_7604);
nand U8524 (N_8524,N_7344,N_6057);
nor U8525 (N_8525,N_7463,N_6467);
or U8526 (N_8526,N_7594,N_6214);
or U8527 (N_8527,N_6806,N_6361);
nand U8528 (N_8528,N_7103,N_6286);
or U8529 (N_8529,N_7257,N_7969);
xor U8530 (N_8530,N_6345,N_6364);
nand U8531 (N_8531,N_6860,N_7277);
or U8532 (N_8532,N_6411,N_6336);
or U8533 (N_8533,N_6151,N_7972);
and U8534 (N_8534,N_6162,N_7698);
or U8535 (N_8535,N_7929,N_7508);
and U8536 (N_8536,N_7312,N_7664);
xnor U8537 (N_8537,N_6985,N_7911);
xnor U8538 (N_8538,N_7248,N_7816);
nand U8539 (N_8539,N_7520,N_7184);
nor U8540 (N_8540,N_6426,N_6248);
xnor U8541 (N_8541,N_6675,N_6089);
or U8542 (N_8542,N_7167,N_6596);
or U8543 (N_8543,N_6878,N_6606);
nor U8544 (N_8544,N_7703,N_6302);
and U8545 (N_8545,N_7967,N_7579);
nand U8546 (N_8546,N_6099,N_7580);
xnor U8547 (N_8547,N_6532,N_7133);
nand U8548 (N_8548,N_6440,N_7098);
and U8549 (N_8549,N_7306,N_6903);
and U8550 (N_8550,N_6076,N_7459);
xnor U8551 (N_8551,N_7195,N_7047);
or U8552 (N_8552,N_6618,N_6597);
or U8553 (N_8553,N_7831,N_7685);
nor U8554 (N_8554,N_6101,N_7357);
or U8555 (N_8555,N_7634,N_7802);
nand U8556 (N_8556,N_7022,N_6831);
and U8557 (N_8557,N_6964,N_7639);
nand U8558 (N_8558,N_7307,N_6182);
xnor U8559 (N_8559,N_7460,N_7569);
and U8560 (N_8560,N_7811,N_6450);
and U8561 (N_8561,N_6326,N_7503);
nor U8562 (N_8562,N_7217,N_6813);
nand U8563 (N_8563,N_6395,N_6325);
or U8564 (N_8564,N_6270,N_7823);
xor U8565 (N_8565,N_7686,N_7630);
nor U8566 (N_8566,N_7060,N_7766);
nor U8567 (N_8567,N_6229,N_7075);
or U8568 (N_8568,N_7636,N_6112);
and U8569 (N_8569,N_7493,N_7403);
and U8570 (N_8570,N_7691,N_7771);
and U8571 (N_8571,N_6641,N_6246);
nor U8572 (N_8572,N_7779,N_6070);
or U8573 (N_8573,N_6901,N_6854);
or U8574 (N_8574,N_6771,N_6698);
nand U8575 (N_8575,N_6290,N_6288);
nand U8576 (N_8576,N_6875,N_7943);
or U8577 (N_8577,N_7428,N_7271);
or U8578 (N_8578,N_6865,N_6777);
nor U8579 (N_8579,N_6058,N_6210);
or U8580 (N_8580,N_7166,N_6990);
nor U8581 (N_8581,N_6022,N_7694);
nand U8582 (N_8582,N_7208,N_6226);
nand U8583 (N_8583,N_7023,N_7329);
or U8584 (N_8584,N_7325,N_7043);
nand U8585 (N_8585,N_7455,N_7826);
or U8586 (N_8586,N_6129,N_7919);
or U8587 (N_8587,N_6365,N_7659);
and U8588 (N_8588,N_6154,N_6510);
and U8589 (N_8589,N_6424,N_7282);
nand U8590 (N_8590,N_7775,N_7091);
nand U8591 (N_8591,N_6238,N_7563);
or U8592 (N_8592,N_7394,N_6340);
nor U8593 (N_8593,N_6000,N_6936);
nor U8594 (N_8594,N_6829,N_6736);
nand U8595 (N_8595,N_6632,N_7211);
nor U8596 (N_8596,N_6441,N_6394);
or U8597 (N_8597,N_7514,N_6555);
xnor U8598 (N_8598,N_6892,N_6995);
xnor U8599 (N_8599,N_6471,N_6705);
nor U8600 (N_8600,N_6848,N_7471);
or U8601 (N_8601,N_7862,N_7956);
and U8602 (N_8602,N_6066,N_7440);
nand U8603 (N_8603,N_6445,N_6986);
nor U8604 (N_8604,N_7866,N_6856);
xnor U8605 (N_8605,N_7912,N_6503);
and U8606 (N_8606,N_7139,N_7119);
or U8607 (N_8607,N_6119,N_6982);
nor U8608 (N_8608,N_7845,N_7842);
nand U8609 (N_8609,N_7284,N_7410);
or U8610 (N_8610,N_7233,N_6590);
xnor U8611 (N_8611,N_6306,N_7024);
or U8612 (N_8612,N_7297,N_6170);
nor U8613 (N_8613,N_7707,N_7695);
and U8614 (N_8614,N_6344,N_7643);
xor U8615 (N_8615,N_6245,N_6782);
and U8616 (N_8616,N_6681,N_7907);
nand U8617 (N_8617,N_7979,N_7161);
nand U8618 (N_8618,N_7532,N_6417);
nor U8619 (N_8619,N_6727,N_6276);
nor U8620 (N_8620,N_7078,N_6107);
and U8621 (N_8621,N_6118,N_7207);
xor U8622 (N_8622,N_7458,N_7704);
and U8623 (N_8623,N_7349,N_6678);
and U8624 (N_8624,N_6549,N_6090);
xor U8625 (N_8625,N_6817,N_6946);
nand U8626 (N_8626,N_7511,N_6416);
xnor U8627 (N_8627,N_7549,N_7756);
nand U8628 (N_8628,N_7529,N_7051);
nor U8629 (N_8629,N_7693,N_6012);
or U8630 (N_8630,N_7122,N_7462);
nand U8631 (N_8631,N_7472,N_7701);
nor U8632 (N_8632,N_7827,N_6108);
or U8633 (N_8633,N_7617,N_6722);
nor U8634 (N_8634,N_7214,N_7328);
nand U8635 (N_8635,N_7778,N_6967);
or U8636 (N_8636,N_7977,N_7619);
and U8637 (N_8637,N_7582,N_7692);
or U8638 (N_8638,N_6529,N_7118);
or U8639 (N_8639,N_7905,N_7336);
nor U8640 (N_8640,N_6700,N_6996);
nand U8641 (N_8641,N_7192,N_6494);
nor U8642 (N_8642,N_6713,N_6143);
nor U8643 (N_8643,N_6199,N_7935);
or U8644 (N_8644,N_6543,N_6462);
or U8645 (N_8645,N_6866,N_7268);
or U8646 (N_8646,N_6869,N_7717);
nor U8647 (N_8647,N_7832,N_7884);
nand U8648 (N_8648,N_7751,N_6872);
and U8649 (N_8649,N_6721,N_7401);
nand U8650 (N_8650,N_6600,N_6844);
nor U8651 (N_8651,N_6132,N_7442);
nand U8652 (N_8652,N_6989,N_6670);
xor U8653 (N_8653,N_6180,N_6261);
xor U8654 (N_8654,N_6885,N_7179);
nand U8655 (N_8655,N_6889,N_6216);
nor U8656 (N_8656,N_6933,N_7064);
nor U8657 (N_8657,N_7815,N_6301);
nor U8658 (N_8658,N_7671,N_7193);
or U8659 (N_8659,N_7338,N_7995);
xnor U8660 (N_8660,N_7252,N_7812);
xnor U8661 (N_8661,N_6580,N_7013);
and U8662 (N_8662,N_6567,N_6711);
xnor U8663 (N_8663,N_7688,N_6347);
nand U8664 (N_8664,N_6184,N_7752);
nand U8665 (N_8665,N_6775,N_7537);
or U8666 (N_8666,N_7261,N_7902);
nor U8667 (N_8667,N_6204,N_6220);
nand U8668 (N_8668,N_7589,N_7246);
or U8669 (N_8669,N_7869,N_7709);
or U8670 (N_8670,N_6310,N_7265);
and U8671 (N_8671,N_6013,N_7893);
nand U8672 (N_8672,N_7748,N_6616);
nor U8673 (N_8673,N_7489,N_7432);
nand U8674 (N_8674,N_7062,N_6741);
nor U8675 (N_8675,N_6035,N_6905);
or U8676 (N_8676,N_6554,N_7599);
and U8677 (N_8677,N_6971,N_7077);
or U8678 (N_8678,N_6998,N_6153);
nor U8679 (N_8679,N_7216,N_6773);
nand U8680 (N_8680,N_6888,N_7396);
xor U8681 (N_8681,N_7647,N_7298);
xor U8682 (N_8682,N_7897,N_6173);
and U8683 (N_8683,N_6521,N_6005);
or U8684 (N_8684,N_6913,N_6863);
nor U8685 (N_8685,N_7786,N_6200);
or U8686 (N_8686,N_7223,N_7026);
or U8687 (N_8687,N_6784,N_7273);
or U8688 (N_8688,N_7517,N_6959);
nor U8689 (N_8689,N_7258,N_6278);
and U8690 (N_8690,N_6999,N_6896);
nor U8691 (N_8691,N_6586,N_7828);
and U8692 (N_8692,N_7303,N_7731);
xnor U8693 (N_8693,N_6131,N_7264);
nor U8694 (N_8694,N_6612,N_6337);
or U8695 (N_8695,N_6868,N_6422);
nand U8696 (N_8696,N_7001,N_7715);
or U8697 (N_8697,N_6792,N_6243);
or U8698 (N_8698,N_7235,N_6068);
and U8699 (N_8699,N_6322,N_6189);
or U8700 (N_8700,N_7896,N_7295);
or U8701 (N_8701,N_6712,N_7236);
nor U8702 (N_8702,N_7622,N_6974);
nand U8703 (N_8703,N_7545,N_6157);
or U8704 (N_8704,N_7477,N_7656);
xor U8705 (N_8705,N_6702,N_6311);
nor U8706 (N_8706,N_7456,N_6789);
and U8707 (N_8707,N_6614,N_7914);
nand U8708 (N_8708,N_6605,N_6224);
nand U8709 (N_8709,N_6909,N_6840);
or U8710 (N_8710,N_6683,N_6656);
nand U8711 (N_8711,N_7927,N_6851);
nor U8712 (N_8712,N_7957,N_6690);
nor U8713 (N_8713,N_6753,N_6435);
xor U8714 (N_8714,N_6397,N_6568);
or U8715 (N_8715,N_7637,N_6940);
or U8716 (N_8716,N_6657,N_7301);
xor U8717 (N_8717,N_7124,N_7281);
nor U8718 (N_8718,N_7005,N_7553);
xnor U8719 (N_8719,N_7645,N_6296);
nand U8720 (N_8720,N_7376,N_7010);
and U8721 (N_8721,N_6537,N_6215);
nand U8722 (N_8722,N_7397,N_6455);
xnor U8723 (N_8723,N_6007,N_6778);
nor U8724 (N_8724,N_7157,N_6354);
xor U8725 (N_8725,N_7794,N_7931);
xnor U8726 (N_8726,N_6668,N_6060);
xor U8727 (N_8727,N_7017,N_6924);
or U8728 (N_8728,N_6598,N_7980);
and U8729 (N_8729,N_6786,N_7149);
and U8730 (N_8730,N_7711,N_7411);
nand U8731 (N_8731,N_7247,N_7018);
nor U8732 (N_8732,N_6506,N_6582);
nand U8733 (N_8733,N_7976,N_7099);
nor U8734 (N_8734,N_6949,N_6239);
xnor U8735 (N_8735,N_7922,N_6916);
or U8736 (N_8736,N_7519,N_6952);
and U8737 (N_8737,N_7200,N_7400);
xor U8738 (N_8738,N_6968,N_7164);
or U8739 (N_8739,N_7993,N_6392);
xor U8740 (N_8740,N_6120,N_6181);
xor U8741 (N_8741,N_6939,N_6346);
or U8742 (N_8742,N_7901,N_7654);
nand U8743 (N_8743,N_6900,N_7906);
and U8744 (N_8744,N_6944,N_7021);
xnor U8745 (N_8745,N_7255,N_6839);
nor U8746 (N_8746,N_6264,N_6978);
or U8747 (N_8747,N_7713,N_7390);
or U8748 (N_8748,N_6828,N_7158);
nand U8749 (N_8749,N_7012,N_7335);
xor U8750 (N_8750,N_6807,N_6966);
nor U8751 (N_8751,N_6745,N_7880);
xnor U8752 (N_8752,N_6470,N_7544);
nand U8753 (N_8753,N_6217,N_6685);
and U8754 (N_8754,N_6323,N_7186);
or U8755 (N_8755,N_7059,N_7668);
nor U8756 (N_8756,N_6438,N_6307);
xnor U8757 (N_8757,N_7602,N_6123);
and U8758 (N_8758,N_7534,N_7669);
xor U8759 (N_8759,N_7974,N_7853);
nand U8760 (N_8760,N_7153,N_7318);
nand U8761 (N_8761,N_7346,N_7188);
nand U8762 (N_8762,N_6409,N_7558);
and U8763 (N_8763,N_7177,N_7541);
nand U8764 (N_8764,N_7870,N_6733);
xor U8765 (N_8765,N_6684,N_6370);
or U8766 (N_8766,N_7011,N_7443);
nor U8767 (N_8767,N_6992,N_6830);
nand U8768 (N_8768,N_6314,N_6443);
nand U8769 (N_8769,N_6478,N_6664);
and U8770 (N_8770,N_6929,N_7895);
xor U8771 (N_8771,N_7492,N_7512);
or U8772 (N_8772,N_6293,N_7909);
or U8773 (N_8773,N_6818,N_7020);
nor U8774 (N_8774,N_6026,N_7222);
xnor U8775 (N_8775,N_6881,N_6432);
nor U8776 (N_8776,N_7867,N_6073);
or U8777 (N_8777,N_7151,N_6399);
or U8778 (N_8778,N_7354,N_6164);
nor U8779 (N_8779,N_6701,N_7069);
xnor U8780 (N_8780,N_6042,N_6353);
nand U8781 (N_8781,N_6393,N_7392);
nand U8782 (N_8782,N_6837,N_7987);
xnor U8783 (N_8783,N_6994,N_6328);
nor U8784 (N_8784,N_7379,N_7738);
or U8785 (N_8785,N_6615,N_7323);
xor U8786 (N_8786,N_6251,N_7345);
nand U8787 (N_8787,N_7657,N_6324);
nor U8788 (N_8788,N_7415,N_7272);
nand U8789 (N_8789,N_7182,N_6629);
nor U8790 (N_8790,N_6275,N_6338);
or U8791 (N_8791,N_6146,N_6109);
nor U8792 (N_8792,N_7986,N_6031);
and U8793 (N_8793,N_6065,N_7082);
and U8794 (N_8794,N_6105,N_7705);
xnor U8795 (N_8795,N_6981,N_7121);
xnor U8796 (N_8796,N_7646,N_6297);
or U8797 (N_8797,N_6202,N_7304);
xnor U8798 (N_8798,N_7733,N_7501);
xor U8799 (N_8799,N_7829,N_6034);
or U8800 (N_8800,N_6059,N_7570);
xor U8801 (N_8801,N_7470,N_7212);
or U8802 (N_8802,N_7127,N_7035);
nor U8803 (N_8803,N_7190,N_6262);
nor U8804 (N_8804,N_6027,N_6428);
nand U8805 (N_8805,N_6595,N_6779);
nand U8806 (N_8806,N_7486,N_7391);
and U8807 (N_8807,N_6622,N_7735);
and U8808 (N_8808,N_6882,N_6178);
or U8809 (N_8809,N_6796,N_6564);
and U8810 (N_8810,N_6669,N_6476);
nor U8811 (N_8811,N_6376,N_7330);
xor U8812 (N_8812,N_6895,N_7947);
nor U8813 (N_8813,N_6819,N_7196);
or U8814 (N_8814,N_7620,N_7609);
and U8815 (N_8815,N_6750,N_6384);
nor U8816 (N_8816,N_6942,N_6321);
nand U8817 (N_8817,N_7640,N_7655);
or U8818 (N_8818,N_6672,N_7170);
xor U8819 (N_8819,N_7581,N_7154);
and U8820 (N_8820,N_6196,N_6661);
xor U8821 (N_8821,N_7997,N_6150);
and U8822 (N_8822,N_7765,N_6413);
and U8823 (N_8823,N_6295,N_7614);
xnor U8824 (N_8824,N_7369,N_7998);
nand U8825 (N_8825,N_7773,N_6010);
nor U8826 (N_8826,N_7667,N_6097);
xnor U8827 (N_8827,N_7834,N_6254);
xnor U8828 (N_8828,N_7635,N_6149);
and U8829 (N_8829,N_6298,N_6212);
xor U8830 (N_8830,N_6454,N_6873);
nor U8831 (N_8831,N_7266,N_7784);
nand U8832 (N_8832,N_7757,N_6746);
nand U8833 (N_8833,N_7431,N_6643);
nand U8834 (N_8834,N_7322,N_6639);
or U8835 (N_8835,N_7810,N_6247);
or U8836 (N_8836,N_7434,N_7852);
nor U8837 (N_8837,N_6970,N_6127);
xnor U8838 (N_8838,N_7086,N_7080);
xor U8839 (N_8839,N_6757,N_7296);
xor U8840 (N_8840,N_7364,N_6660);
nand U8841 (N_8841,N_6571,N_6897);
nand U8842 (N_8842,N_6926,N_7019);
or U8843 (N_8843,N_6666,N_7294);
nand U8844 (N_8844,N_7813,N_7358);
and U8845 (N_8845,N_6374,N_6033);
nor U8846 (N_8846,N_7839,N_6531);
nand U8847 (N_8847,N_7014,N_7797);
nand U8848 (N_8848,N_6972,N_6706);
nand U8849 (N_8849,N_6379,N_6724);
nor U8850 (N_8850,N_6405,N_6427);
xnor U8851 (N_8851,N_6663,N_6762);
nor U8852 (N_8852,N_7714,N_6720);
nor U8853 (N_8853,N_7398,N_7683);
nor U8854 (N_8854,N_7774,N_6029);
or U8855 (N_8855,N_7868,N_7955);
nand U8856 (N_8856,N_6560,N_7603);
and U8857 (N_8857,N_7444,N_7607);
nor U8858 (N_8858,N_6686,N_7393);
nor U8859 (N_8859,N_6855,N_6449);
or U8860 (N_8860,N_7173,N_7814);
nor U8861 (N_8861,N_6197,N_7632);
nor U8862 (N_8862,N_6619,N_7278);
and U8863 (N_8863,N_6213,N_6136);
xnor U8864 (N_8864,N_6280,N_6960);
or U8865 (N_8865,N_6938,N_6508);
nor U8866 (N_8866,N_7009,N_7205);
nand U8867 (N_8867,N_7105,N_7227);
nand U8868 (N_8868,N_7803,N_7530);
xor U8869 (N_8869,N_6144,N_6228);
and U8870 (N_8870,N_7849,N_7936);
or U8871 (N_8871,N_6843,N_7288);
or U8872 (N_8872,N_7932,N_7058);
and U8873 (N_8873,N_6111,N_6533);
nand U8874 (N_8874,N_6434,N_7822);
xnor U8875 (N_8875,N_7245,N_7908);
nor U8876 (N_8876,N_6608,N_6492);
nor U8877 (N_8877,N_6140,N_7355);
xnor U8878 (N_8878,N_7406,N_6575);
nor U8879 (N_8879,N_6542,N_7841);
xnor U8880 (N_8880,N_7380,N_6704);
xnor U8881 (N_8881,N_7923,N_7885);
and U8882 (N_8882,N_7681,N_7962);
nor U8883 (N_8883,N_7343,N_6277);
nand U8884 (N_8884,N_6166,N_6769);
and U8885 (N_8885,N_7311,N_7526);
and U8886 (N_8886,N_7621,N_7262);
xor U8887 (N_8887,N_6931,N_7110);
nor U8888 (N_8888,N_6519,N_6774);
and U8889 (N_8889,N_6927,N_7446);
nor U8890 (N_8890,N_6135,N_7939);
nand U8891 (N_8891,N_7213,N_6846);
or U8892 (N_8892,N_6919,N_6001);
nand U8893 (N_8893,N_7382,N_6824);
and U8894 (N_8894,N_7404,N_6390);
nand U8895 (N_8895,N_7605,N_6398);
xor U8896 (N_8896,N_7577,N_6474);
nor U8897 (N_8897,N_7416,N_7389);
nor U8898 (N_8898,N_6578,N_6908);
or U8899 (N_8899,N_6418,N_7138);
xnor U8900 (N_8900,N_7881,N_7117);
or U8901 (N_8901,N_6783,N_7744);
and U8902 (N_8902,N_6570,N_7504);
nor U8903 (N_8903,N_7445,N_7441);
xor U8904 (N_8904,N_7782,N_7708);
nand U8905 (N_8905,N_7125,N_7048);
or U8906 (N_8906,N_6452,N_6425);
nand U8907 (N_8907,N_7465,N_7548);
nand U8908 (N_8908,N_7054,N_7762);
nor U8909 (N_8909,N_7310,N_6620);
xor U8910 (N_8910,N_6695,N_6406);
nand U8911 (N_8911,N_7528,N_7436);
xnor U8912 (N_8912,N_7833,N_7949);
xor U8913 (N_8913,N_6208,N_7727);
nand U8914 (N_8914,N_6069,N_6725);
nand U8915 (N_8915,N_7722,N_7371);
and U8916 (N_8916,N_7052,N_7723);
xnor U8917 (N_8917,N_6589,N_6513);
nand U8918 (N_8918,N_6991,N_7210);
nor U8919 (N_8919,N_6211,N_7739);
and U8920 (N_8920,N_7754,N_7764);
nor U8921 (N_8921,N_7513,N_6810);
or U8922 (N_8922,N_6530,N_6134);
and U8923 (N_8923,N_6253,N_7948);
xnor U8924 (N_8924,N_6800,N_7269);
nor U8925 (N_8925,N_7016,N_6283);
nor U8926 (N_8926,N_7930,N_6410);
xnor U8927 (N_8927,N_6623,N_7201);
nor U8928 (N_8928,N_7439,N_6169);
or U8929 (N_8929,N_6030,N_6358);
or U8930 (N_8930,N_6165,N_7189);
xor U8931 (N_8931,N_6743,N_7700);
nand U8932 (N_8932,N_6371,N_7670);
nand U8933 (N_8933,N_7156,N_7225);
nor U8934 (N_8934,N_6188,N_6980);
or U8935 (N_8935,N_6294,N_6802);
and U8936 (N_8936,N_7041,N_6386);
nand U8937 (N_8937,N_7623,N_6617);
xnor U8938 (N_8938,N_7788,N_6525);
and U8939 (N_8939,N_7653,N_7314);
xor U8940 (N_8940,N_7791,N_7172);
nand U8941 (N_8941,N_6341,N_6331);
nand U8942 (N_8942,N_7750,N_7933);
nor U8943 (N_8943,N_6385,N_6594);
or U8944 (N_8944,N_6764,N_6319);
xor U8945 (N_8945,N_7143,N_7332);
nand U8946 (N_8946,N_6523,N_7066);
or U8947 (N_8947,N_7419,N_7283);
nor U8948 (N_8948,N_7740,N_7044);
and U8949 (N_8949,N_7004,N_7409);
or U8950 (N_8950,N_7313,N_7339);
or U8951 (N_8951,N_7425,N_6645);
and U8952 (N_8952,N_6039,N_7785);
or U8953 (N_8953,N_6814,N_7761);
nor U8954 (N_8954,N_7141,N_7992);
or U8955 (N_8955,N_6206,N_6588);
and U8956 (N_8956,N_6052,N_6148);
nor U8957 (N_8957,N_6565,N_6145);
nor U8958 (N_8958,N_7451,N_6781);
xnor U8959 (N_8959,N_7374,N_6534);
nor U8960 (N_8960,N_6002,N_7187);
and U8961 (N_8961,N_6078,N_6155);
or U8962 (N_8962,N_6291,N_6920);
and U8963 (N_8963,N_7855,N_7633);
nor U8964 (N_8964,N_7710,N_6876);
nor U8965 (N_8965,N_6834,N_6822);
or U8966 (N_8966,N_7008,N_7438);
or U8967 (N_8967,N_7551,N_6308);
or U8968 (N_8968,N_6871,N_6583);
and U8969 (N_8969,N_7728,N_6552);
nand U8970 (N_8970,N_7476,N_7760);
or U8971 (N_8971,N_7720,N_6158);
or U8972 (N_8972,N_7971,N_6505);
xnor U8973 (N_8973,N_7854,N_6520);
xnor U8974 (N_8974,N_7665,N_6853);
nor U8975 (N_8975,N_7469,N_7055);
or U8976 (N_8976,N_6958,N_6093);
or U8977 (N_8977,N_6241,N_7944);
or U8978 (N_8978,N_7130,N_7628);
and U8979 (N_8979,N_7123,N_6772);
xor U8980 (N_8980,N_6430,N_6174);
nand U8981 (N_8981,N_7331,N_7430);
xor U8982 (N_8982,N_7384,N_6710);
and U8983 (N_8983,N_7975,N_6709);
and U8984 (N_8984,N_6767,N_6584);
and U8985 (N_8985,N_7673,N_7057);
nand U8986 (N_8986,N_6621,N_6790);
xnor U8987 (N_8987,N_6037,N_6862);
nand U8988 (N_8988,N_6640,N_7970);
nand U8989 (N_8989,N_6050,N_6304);
xor U8990 (N_8990,N_6242,N_6074);
and U8991 (N_8991,N_6883,N_6801);
xnor U8992 (N_8992,N_7302,N_7221);
and U8993 (N_8993,N_6156,N_7917);
or U8994 (N_8994,N_7474,N_6511);
nand U8995 (N_8995,N_6064,N_7982);
or U8996 (N_8996,N_7626,N_7565);
or U8997 (N_8997,N_6043,N_7600);
nor U8998 (N_8998,N_7768,N_7777);
or U8999 (N_8999,N_6160,N_7253);
nor U9000 (N_9000,N_6411,N_6110);
xnor U9001 (N_9001,N_6929,N_7022);
and U9002 (N_9002,N_7958,N_6969);
xnor U9003 (N_9003,N_7955,N_7809);
nor U9004 (N_9004,N_6148,N_7221);
xnor U9005 (N_9005,N_6045,N_7436);
or U9006 (N_9006,N_7179,N_6608);
nor U9007 (N_9007,N_7363,N_7316);
nor U9008 (N_9008,N_7861,N_7817);
nand U9009 (N_9009,N_7110,N_7464);
or U9010 (N_9010,N_7353,N_7081);
or U9011 (N_9011,N_7981,N_6008);
and U9012 (N_9012,N_7033,N_6670);
xnor U9013 (N_9013,N_7642,N_6238);
or U9014 (N_9014,N_6658,N_6488);
nand U9015 (N_9015,N_7574,N_6167);
or U9016 (N_9016,N_7642,N_6226);
nand U9017 (N_9017,N_6962,N_7063);
or U9018 (N_9018,N_6828,N_7114);
xnor U9019 (N_9019,N_7417,N_7756);
nor U9020 (N_9020,N_6823,N_7627);
xor U9021 (N_9021,N_6642,N_7200);
nand U9022 (N_9022,N_6420,N_6069);
nand U9023 (N_9023,N_7824,N_7541);
xor U9024 (N_9024,N_7547,N_6456);
nor U9025 (N_9025,N_6175,N_7373);
xor U9026 (N_9026,N_6300,N_6892);
or U9027 (N_9027,N_7896,N_7858);
or U9028 (N_9028,N_6823,N_6737);
and U9029 (N_9029,N_6496,N_7756);
or U9030 (N_9030,N_7220,N_7497);
xor U9031 (N_9031,N_6832,N_6497);
or U9032 (N_9032,N_7974,N_6711);
or U9033 (N_9033,N_7971,N_7896);
or U9034 (N_9034,N_7106,N_6897);
nor U9035 (N_9035,N_6841,N_6608);
nor U9036 (N_9036,N_7386,N_7256);
nor U9037 (N_9037,N_7458,N_7586);
and U9038 (N_9038,N_6300,N_7298);
xor U9039 (N_9039,N_6778,N_6053);
and U9040 (N_9040,N_6464,N_7729);
and U9041 (N_9041,N_7843,N_6710);
or U9042 (N_9042,N_7275,N_6853);
or U9043 (N_9043,N_6441,N_7647);
nor U9044 (N_9044,N_6559,N_7059);
nor U9045 (N_9045,N_7917,N_6579);
and U9046 (N_9046,N_6066,N_6852);
or U9047 (N_9047,N_6050,N_6131);
nand U9048 (N_9048,N_6201,N_7719);
or U9049 (N_9049,N_7902,N_6087);
nor U9050 (N_9050,N_6512,N_7948);
and U9051 (N_9051,N_7316,N_7998);
and U9052 (N_9052,N_6789,N_6476);
and U9053 (N_9053,N_6487,N_6098);
or U9054 (N_9054,N_6903,N_7715);
nor U9055 (N_9055,N_6709,N_6814);
xor U9056 (N_9056,N_6747,N_6448);
and U9057 (N_9057,N_6406,N_7582);
and U9058 (N_9058,N_6990,N_7284);
nor U9059 (N_9059,N_7858,N_7042);
xor U9060 (N_9060,N_7608,N_6093);
nand U9061 (N_9061,N_7159,N_6112);
and U9062 (N_9062,N_7207,N_7444);
nor U9063 (N_9063,N_7170,N_7830);
nor U9064 (N_9064,N_6865,N_6179);
and U9065 (N_9065,N_6094,N_7284);
and U9066 (N_9066,N_7555,N_7898);
nor U9067 (N_9067,N_7679,N_7479);
nor U9068 (N_9068,N_7486,N_7134);
xor U9069 (N_9069,N_6131,N_7978);
nand U9070 (N_9070,N_7353,N_6080);
xnor U9071 (N_9071,N_7022,N_6829);
xnor U9072 (N_9072,N_7706,N_6552);
or U9073 (N_9073,N_7827,N_6060);
or U9074 (N_9074,N_6232,N_6736);
and U9075 (N_9075,N_6092,N_6756);
xnor U9076 (N_9076,N_7402,N_7774);
and U9077 (N_9077,N_6769,N_6436);
nor U9078 (N_9078,N_7670,N_6707);
xnor U9079 (N_9079,N_6293,N_6344);
and U9080 (N_9080,N_7395,N_6855);
or U9081 (N_9081,N_7613,N_6904);
nor U9082 (N_9082,N_7651,N_6439);
nand U9083 (N_9083,N_7839,N_6824);
and U9084 (N_9084,N_6788,N_7934);
or U9085 (N_9085,N_7683,N_6417);
and U9086 (N_9086,N_6690,N_6716);
nand U9087 (N_9087,N_6585,N_6907);
xor U9088 (N_9088,N_7879,N_7316);
and U9089 (N_9089,N_7739,N_6366);
and U9090 (N_9090,N_6673,N_6323);
or U9091 (N_9091,N_7138,N_6862);
xnor U9092 (N_9092,N_7560,N_6073);
or U9093 (N_9093,N_7699,N_7171);
nand U9094 (N_9094,N_6886,N_7352);
and U9095 (N_9095,N_6096,N_6358);
and U9096 (N_9096,N_6479,N_7420);
or U9097 (N_9097,N_7162,N_7832);
and U9098 (N_9098,N_7335,N_6411);
and U9099 (N_9099,N_7125,N_6684);
and U9100 (N_9100,N_6366,N_6011);
xor U9101 (N_9101,N_6461,N_7648);
nor U9102 (N_9102,N_6874,N_7080);
nand U9103 (N_9103,N_7351,N_6890);
nor U9104 (N_9104,N_7711,N_7415);
xnor U9105 (N_9105,N_6441,N_6801);
and U9106 (N_9106,N_7493,N_6700);
xor U9107 (N_9107,N_6169,N_7487);
nor U9108 (N_9108,N_6963,N_7666);
xnor U9109 (N_9109,N_6431,N_6909);
nand U9110 (N_9110,N_6352,N_6355);
and U9111 (N_9111,N_6206,N_7828);
nor U9112 (N_9112,N_7213,N_7881);
xnor U9113 (N_9113,N_7997,N_6992);
xor U9114 (N_9114,N_7066,N_7864);
xor U9115 (N_9115,N_7714,N_7928);
xnor U9116 (N_9116,N_7983,N_7390);
and U9117 (N_9117,N_7956,N_6341);
nand U9118 (N_9118,N_6363,N_7980);
nand U9119 (N_9119,N_6388,N_7213);
or U9120 (N_9120,N_6699,N_7690);
and U9121 (N_9121,N_7430,N_7542);
xor U9122 (N_9122,N_7729,N_6523);
xor U9123 (N_9123,N_7823,N_7478);
xor U9124 (N_9124,N_6718,N_7436);
and U9125 (N_9125,N_7875,N_6752);
xor U9126 (N_9126,N_7382,N_7702);
and U9127 (N_9127,N_7538,N_6344);
or U9128 (N_9128,N_6539,N_6206);
nand U9129 (N_9129,N_7130,N_7403);
or U9130 (N_9130,N_6182,N_7824);
nand U9131 (N_9131,N_7477,N_6285);
xor U9132 (N_9132,N_6199,N_6668);
and U9133 (N_9133,N_6456,N_7983);
nand U9134 (N_9134,N_7721,N_7242);
nand U9135 (N_9135,N_7856,N_6235);
nand U9136 (N_9136,N_7618,N_7568);
or U9137 (N_9137,N_6511,N_6517);
and U9138 (N_9138,N_7743,N_6454);
xnor U9139 (N_9139,N_7758,N_6216);
or U9140 (N_9140,N_7413,N_6649);
and U9141 (N_9141,N_7350,N_6985);
xor U9142 (N_9142,N_7453,N_6864);
nand U9143 (N_9143,N_7868,N_6612);
or U9144 (N_9144,N_7611,N_6526);
xnor U9145 (N_9145,N_7267,N_7285);
xnor U9146 (N_9146,N_6843,N_7024);
nand U9147 (N_9147,N_7458,N_7378);
nand U9148 (N_9148,N_6321,N_6650);
and U9149 (N_9149,N_6665,N_7844);
xnor U9150 (N_9150,N_6175,N_6608);
nor U9151 (N_9151,N_6256,N_6305);
and U9152 (N_9152,N_6638,N_7941);
nand U9153 (N_9153,N_6526,N_7853);
nand U9154 (N_9154,N_7998,N_7008);
xor U9155 (N_9155,N_7854,N_6469);
nor U9156 (N_9156,N_6820,N_6630);
nor U9157 (N_9157,N_7625,N_6821);
nand U9158 (N_9158,N_7677,N_7094);
nand U9159 (N_9159,N_7628,N_6672);
and U9160 (N_9160,N_6850,N_6463);
and U9161 (N_9161,N_7833,N_7884);
and U9162 (N_9162,N_6127,N_6203);
xnor U9163 (N_9163,N_7864,N_6950);
and U9164 (N_9164,N_7107,N_7614);
and U9165 (N_9165,N_6999,N_6327);
or U9166 (N_9166,N_6714,N_7295);
nor U9167 (N_9167,N_7210,N_7966);
and U9168 (N_9168,N_6267,N_6482);
xor U9169 (N_9169,N_6718,N_6783);
nor U9170 (N_9170,N_6369,N_6278);
or U9171 (N_9171,N_6530,N_6985);
nor U9172 (N_9172,N_7114,N_6478);
and U9173 (N_9173,N_7045,N_7562);
nor U9174 (N_9174,N_6745,N_7099);
and U9175 (N_9175,N_6155,N_7647);
or U9176 (N_9176,N_7610,N_6683);
nor U9177 (N_9177,N_6329,N_7647);
or U9178 (N_9178,N_7140,N_7816);
and U9179 (N_9179,N_7587,N_6954);
nand U9180 (N_9180,N_6264,N_6139);
and U9181 (N_9181,N_6788,N_7169);
nor U9182 (N_9182,N_6818,N_7053);
or U9183 (N_9183,N_6923,N_7474);
nand U9184 (N_9184,N_7763,N_7914);
and U9185 (N_9185,N_6048,N_7962);
and U9186 (N_9186,N_7105,N_7812);
nand U9187 (N_9187,N_6873,N_7532);
xor U9188 (N_9188,N_6786,N_7034);
or U9189 (N_9189,N_6607,N_6229);
nor U9190 (N_9190,N_6361,N_7990);
nor U9191 (N_9191,N_7085,N_7140);
xor U9192 (N_9192,N_7514,N_6619);
nand U9193 (N_9193,N_6021,N_6581);
and U9194 (N_9194,N_6886,N_7438);
or U9195 (N_9195,N_7300,N_7689);
and U9196 (N_9196,N_7839,N_7327);
nand U9197 (N_9197,N_7603,N_6235);
or U9198 (N_9198,N_6118,N_7908);
nor U9199 (N_9199,N_6863,N_7761);
or U9200 (N_9200,N_6749,N_7514);
and U9201 (N_9201,N_6836,N_6141);
xnor U9202 (N_9202,N_6878,N_6083);
and U9203 (N_9203,N_7002,N_7651);
nand U9204 (N_9204,N_6589,N_7411);
nand U9205 (N_9205,N_7740,N_6392);
xor U9206 (N_9206,N_6184,N_7615);
and U9207 (N_9207,N_7332,N_6346);
xnor U9208 (N_9208,N_7063,N_6122);
nand U9209 (N_9209,N_7509,N_6271);
or U9210 (N_9210,N_7001,N_7285);
or U9211 (N_9211,N_7099,N_7346);
or U9212 (N_9212,N_6389,N_6159);
nor U9213 (N_9213,N_6808,N_7092);
and U9214 (N_9214,N_6837,N_7596);
xnor U9215 (N_9215,N_7136,N_7902);
nand U9216 (N_9216,N_6449,N_6620);
nand U9217 (N_9217,N_6990,N_6941);
or U9218 (N_9218,N_7009,N_6603);
xnor U9219 (N_9219,N_7382,N_6399);
nor U9220 (N_9220,N_6364,N_6334);
nand U9221 (N_9221,N_6017,N_6467);
nor U9222 (N_9222,N_6785,N_6402);
nand U9223 (N_9223,N_6451,N_7021);
xnor U9224 (N_9224,N_6072,N_6996);
xnor U9225 (N_9225,N_7979,N_6392);
nand U9226 (N_9226,N_6503,N_6439);
nor U9227 (N_9227,N_6099,N_7890);
xor U9228 (N_9228,N_7517,N_7046);
nand U9229 (N_9229,N_6260,N_7762);
nor U9230 (N_9230,N_7275,N_7369);
xor U9231 (N_9231,N_7876,N_6552);
nor U9232 (N_9232,N_6820,N_7080);
nand U9233 (N_9233,N_6521,N_7562);
nor U9234 (N_9234,N_7625,N_6307);
nand U9235 (N_9235,N_6999,N_6777);
xor U9236 (N_9236,N_6907,N_7358);
nand U9237 (N_9237,N_7156,N_7055);
and U9238 (N_9238,N_6884,N_7439);
nor U9239 (N_9239,N_7095,N_6691);
nor U9240 (N_9240,N_7935,N_7329);
nor U9241 (N_9241,N_6762,N_7892);
or U9242 (N_9242,N_7982,N_7821);
nor U9243 (N_9243,N_7838,N_7618);
and U9244 (N_9244,N_6367,N_6491);
nand U9245 (N_9245,N_6138,N_6117);
or U9246 (N_9246,N_6488,N_6752);
xnor U9247 (N_9247,N_7438,N_6778);
nand U9248 (N_9248,N_7542,N_7809);
nand U9249 (N_9249,N_7321,N_6431);
and U9250 (N_9250,N_6784,N_6758);
and U9251 (N_9251,N_6672,N_7981);
and U9252 (N_9252,N_7202,N_7442);
nor U9253 (N_9253,N_6567,N_6943);
xnor U9254 (N_9254,N_7695,N_6185);
xnor U9255 (N_9255,N_7475,N_6879);
xor U9256 (N_9256,N_6174,N_7050);
and U9257 (N_9257,N_6248,N_6897);
and U9258 (N_9258,N_6262,N_7531);
nand U9259 (N_9259,N_6595,N_7881);
and U9260 (N_9260,N_6734,N_6769);
xnor U9261 (N_9261,N_7354,N_7401);
nand U9262 (N_9262,N_7011,N_6489);
or U9263 (N_9263,N_6951,N_6477);
xor U9264 (N_9264,N_6318,N_7409);
and U9265 (N_9265,N_6380,N_6522);
and U9266 (N_9266,N_7328,N_6829);
xor U9267 (N_9267,N_6825,N_6742);
and U9268 (N_9268,N_7462,N_6391);
and U9269 (N_9269,N_6322,N_6361);
xnor U9270 (N_9270,N_6433,N_6415);
nor U9271 (N_9271,N_6830,N_6414);
nor U9272 (N_9272,N_6804,N_6135);
xnor U9273 (N_9273,N_7983,N_7089);
nand U9274 (N_9274,N_6707,N_6869);
nor U9275 (N_9275,N_6140,N_6785);
nor U9276 (N_9276,N_7539,N_6138);
xor U9277 (N_9277,N_6220,N_7684);
xor U9278 (N_9278,N_6684,N_7766);
xor U9279 (N_9279,N_6285,N_6241);
nand U9280 (N_9280,N_7405,N_7958);
nor U9281 (N_9281,N_7305,N_7529);
nor U9282 (N_9282,N_6629,N_7956);
nand U9283 (N_9283,N_6416,N_7983);
nand U9284 (N_9284,N_7262,N_7003);
and U9285 (N_9285,N_6261,N_7299);
and U9286 (N_9286,N_7674,N_7020);
nor U9287 (N_9287,N_7022,N_7416);
or U9288 (N_9288,N_7055,N_7927);
or U9289 (N_9289,N_6899,N_6816);
nor U9290 (N_9290,N_6696,N_7369);
or U9291 (N_9291,N_6606,N_6334);
xor U9292 (N_9292,N_7785,N_6743);
nand U9293 (N_9293,N_7761,N_6807);
xnor U9294 (N_9294,N_7870,N_6473);
and U9295 (N_9295,N_6523,N_7349);
or U9296 (N_9296,N_7988,N_7970);
xnor U9297 (N_9297,N_6872,N_7022);
xor U9298 (N_9298,N_7343,N_6891);
nor U9299 (N_9299,N_6316,N_6076);
or U9300 (N_9300,N_7491,N_7063);
nor U9301 (N_9301,N_6756,N_7838);
nand U9302 (N_9302,N_6118,N_6311);
or U9303 (N_9303,N_6087,N_7402);
and U9304 (N_9304,N_7396,N_7864);
and U9305 (N_9305,N_6653,N_6275);
nand U9306 (N_9306,N_6728,N_7686);
xor U9307 (N_9307,N_7649,N_6147);
xnor U9308 (N_9308,N_6092,N_7893);
xnor U9309 (N_9309,N_6533,N_6004);
or U9310 (N_9310,N_6733,N_6910);
xnor U9311 (N_9311,N_7313,N_7404);
nor U9312 (N_9312,N_7878,N_6219);
or U9313 (N_9313,N_6152,N_7016);
and U9314 (N_9314,N_7463,N_6130);
nand U9315 (N_9315,N_6185,N_7205);
xor U9316 (N_9316,N_6067,N_6939);
and U9317 (N_9317,N_6115,N_6223);
or U9318 (N_9318,N_7998,N_7075);
and U9319 (N_9319,N_6282,N_7870);
or U9320 (N_9320,N_7190,N_6915);
xnor U9321 (N_9321,N_7078,N_7736);
or U9322 (N_9322,N_6303,N_6065);
nand U9323 (N_9323,N_7224,N_6103);
nor U9324 (N_9324,N_7725,N_7146);
nor U9325 (N_9325,N_7172,N_7057);
or U9326 (N_9326,N_6863,N_7520);
nand U9327 (N_9327,N_7702,N_7371);
nand U9328 (N_9328,N_7847,N_6408);
or U9329 (N_9329,N_7885,N_6666);
or U9330 (N_9330,N_6950,N_7104);
nor U9331 (N_9331,N_7935,N_7499);
nor U9332 (N_9332,N_6871,N_7804);
and U9333 (N_9333,N_7924,N_7082);
nor U9334 (N_9334,N_6325,N_6143);
and U9335 (N_9335,N_7788,N_7348);
xor U9336 (N_9336,N_7588,N_6567);
nor U9337 (N_9337,N_7036,N_6075);
nand U9338 (N_9338,N_7066,N_7136);
xnor U9339 (N_9339,N_6498,N_7521);
xnor U9340 (N_9340,N_7506,N_6432);
xnor U9341 (N_9341,N_7275,N_6884);
or U9342 (N_9342,N_6198,N_6793);
nand U9343 (N_9343,N_6842,N_6278);
xnor U9344 (N_9344,N_7334,N_6645);
nand U9345 (N_9345,N_7092,N_7432);
and U9346 (N_9346,N_7529,N_6767);
nor U9347 (N_9347,N_7430,N_7830);
or U9348 (N_9348,N_7575,N_6218);
and U9349 (N_9349,N_7178,N_6505);
or U9350 (N_9350,N_6408,N_7981);
or U9351 (N_9351,N_7176,N_6757);
nand U9352 (N_9352,N_7409,N_6358);
and U9353 (N_9353,N_7385,N_7242);
nor U9354 (N_9354,N_7383,N_6132);
and U9355 (N_9355,N_6281,N_7900);
nor U9356 (N_9356,N_6181,N_7416);
and U9357 (N_9357,N_6451,N_7484);
and U9358 (N_9358,N_6606,N_6209);
or U9359 (N_9359,N_6014,N_6080);
and U9360 (N_9360,N_6005,N_7078);
or U9361 (N_9361,N_6119,N_7189);
xnor U9362 (N_9362,N_6125,N_7752);
and U9363 (N_9363,N_6692,N_6475);
xnor U9364 (N_9364,N_6570,N_7461);
xnor U9365 (N_9365,N_7250,N_7571);
or U9366 (N_9366,N_6461,N_7673);
nor U9367 (N_9367,N_7655,N_7233);
xor U9368 (N_9368,N_6617,N_7473);
xor U9369 (N_9369,N_6869,N_6646);
nand U9370 (N_9370,N_6725,N_7855);
nor U9371 (N_9371,N_7432,N_7321);
or U9372 (N_9372,N_7552,N_7611);
nand U9373 (N_9373,N_6878,N_6900);
or U9374 (N_9374,N_6981,N_6387);
nor U9375 (N_9375,N_7850,N_7676);
nand U9376 (N_9376,N_6167,N_6996);
nand U9377 (N_9377,N_7036,N_6830);
and U9378 (N_9378,N_6467,N_6432);
xnor U9379 (N_9379,N_7538,N_7373);
nor U9380 (N_9380,N_7980,N_7423);
nand U9381 (N_9381,N_7743,N_6913);
xnor U9382 (N_9382,N_6028,N_6755);
xor U9383 (N_9383,N_7058,N_7855);
or U9384 (N_9384,N_6209,N_6462);
or U9385 (N_9385,N_7018,N_6654);
nor U9386 (N_9386,N_7511,N_7857);
and U9387 (N_9387,N_6348,N_6406);
xor U9388 (N_9388,N_7334,N_7137);
nand U9389 (N_9389,N_6220,N_6785);
xnor U9390 (N_9390,N_6638,N_6766);
nand U9391 (N_9391,N_6185,N_7549);
or U9392 (N_9392,N_7663,N_6989);
nand U9393 (N_9393,N_6988,N_7716);
xnor U9394 (N_9394,N_7344,N_7710);
or U9395 (N_9395,N_7788,N_6415);
xnor U9396 (N_9396,N_6419,N_7960);
nor U9397 (N_9397,N_7947,N_7554);
nand U9398 (N_9398,N_6666,N_7597);
xnor U9399 (N_9399,N_6552,N_6650);
and U9400 (N_9400,N_7863,N_7682);
xor U9401 (N_9401,N_6757,N_6641);
and U9402 (N_9402,N_6137,N_7952);
and U9403 (N_9403,N_7636,N_7366);
nor U9404 (N_9404,N_7818,N_6240);
xnor U9405 (N_9405,N_7825,N_7866);
and U9406 (N_9406,N_7284,N_6074);
or U9407 (N_9407,N_6987,N_7476);
nand U9408 (N_9408,N_7538,N_6607);
xor U9409 (N_9409,N_6441,N_6427);
and U9410 (N_9410,N_6980,N_6124);
and U9411 (N_9411,N_6328,N_7186);
xnor U9412 (N_9412,N_6803,N_7810);
nor U9413 (N_9413,N_6894,N_6009);
nor U9414 (N_9414,N_7746,N_6559);
nand U9415 (N_9415,N_6708,N_6077);
nand U9416 (N_9416,N_7768,N_6724);
nand U9417 (N_9417,N_6290,N_6735);
nand U9418 (N_9418,N_6036,N_7985);
nand U9419 (N_9419,N_7981,N_6209);
xnor U9420 (N_9420,N_6368,N_7282);
and U9421 (N_9421,N_7513,N_7055);
xor U9422 (N_9422,N_7512,N_6141);
and U9423 (N_9423,N_6909,N_6403);
and U9424 (N_9424,N_7259,N_7533);
xor U9425 (N_9425,N_6451,N_6597);
nand U9426 (N_9426,N_6309,N_7443);
nor U9427 (N_9427,N_7112,N_6433);
or U9428 (N_9428,N_6253,N_7652);
nor U9429 (N_9429,N_6634,N_7119);
and U9430 (N_9430,N_7495,N_7999);
xor U9431 (N_9431,N_7927,N_6655);
nand U9432 (N_9432,N_6457,N_7137);
or U9433 (N_9433,N_7972,N_6770);
or U9434 (N_9434,N_6897,N_6734);
and U9435 (N_9435,N_7689,N_7460);
nor U9436 (N_9436,N_6338,N_6498);
and U9437 (N_9437,N_7470,N_6072);
nand U9438 (N_9438,N_6003,N_7734);
and U9439 (N_9439,N_6168,N_6353);
nor U9440 (N_9440,N_6348,N_7910);
or U9441 (N_9441,N_6142,N_7910);
xnor U9442 (N_9442,N_7987,N_7296);
or U9443 (N_9443,N_7310,N_6348);
nand U9444 (N_9444,N_7610,N_6684);
nand U9445 (N_9445,N_6333,N_6110);
and U9446 (N_9446,N_6212,N_6474);
or U9447 (N_9447,N_6333,N_6197);
and U9448 (N_9448,N_7770,N_7568);
xnor U9449 (N_9449,N_7681,N_7726);
nand U9450 (N_9450,N_7121,N_7234);
nand U9451 (N_9451,N_7200,N_7812);
nand U9452 (N_9452,N_7815,N_6829);
nor U9453 (N_9453,N_6395,N_7830);
or U9454 (N_9454,N_6304,N_6242);
nor U9455 (N_9455,N_7446,N_6967);
xnor U9456 (N_9456,N_7578,N_7386);
or U9457 (N_9457,N_7128,N_7535);
and U9458 (N_9458,N_7459,N_6536);
xor U9459 (N_9459,N_7866,N_6350);
xor U9460 (N_9460,N_7888,N_6292);
xor U9461 (N_9461,N_6940,N_6359);
and U9462 (N_9462,N_6426,N_6039);
and U9463 (N_9463,N_6658,N_6330);
nor U9464 (N_9464,N_7990,N_6068);
or U9465 (N_9465,N_6696,N_7414);
xor U9466 (N_9466,N_7872,N_6356);
and U9467 (N_9467,N_7609,N_7918);
or U9468 (N_9468,N_7447,N_7449);
xnor U9469 (N_9469,N_7610,N_6803);
xnor U9470 (N_9470,N_6983,N_6031);
or U9471 (N_9471,N_7966,N_7553);
or U9472 (N_9472,N_7553,N_6488);
nand U9473 (N_9473,N_6193,N_6148);
nand U9474 (N_9474,N_7560,N_6726);
nor U9475 (N_9475,N_6887,N_6117);
nand U9476 (N_9476,N_6601,N_7950);
or U9477 (N_9477,N_6863,N_6137);
and U9478 (N_9478,N_7078,N_6831);
and U9479 (N_9479,N_7038,N_6735);
nand U9480 (N_9480,N_6605,N_7997);
and U9481 (N_9481,N_7468,N_7688);
nand U9482 (N_9482,N_6060,N_7428);
and U9483 (N_9483,N_7827,N_7678);
nor U9484 (N_9484,N_7119,N_6866);
and U9485 (N_9485,N_7754,N_6672);
and U9486 (N_9486,N_6651,N_7506);
nand U9487 (N_9487,N_7806,N_6697);
xor U9488 (N_9488,N_6448,N_7118);
xnor U9489 (N_9489,N_7235,N_6670);
nand U9490 (N_9490,N_7977,N_7316);
xor U9491 (N_9491,N_6471,N_7707);
nor U9492 (N_9492,N_7212,N_7170);
nor U9493 (N_9493,N_7739,N_7835);
nand U9494 (N_9494,N_6928,N_7565);
xor U9495 (N_9495,N_6873,N_7311);
and U9496 (N_9496,N_6219,N_7874);
xor U9497 (N_9497,N_7675,N_6702);
or U9498 (N_9498,N_7545,N_7777);
nand U9499 (N_9499,N_6632,N_7853);
xnor U9500 (N_9500,N_6408,N_6681);
and U9501 (N_9501,N_7915,N_7135);
nor U9502 (N_9502,N_7068,N_6939);
nor U9503 (N_9503,N_7098,N_6694);
nor U9504 (N_9504,N_6741,N_7735);
nor U9505 (N_9505,N_6611,N_6307);
nor U9506 (N_9506,N_6371,N_6825);
or U9507 (N_9507,N_6710,N_7579);
nor U9508 (N_9508,N_7252,N_6591);
xnor U9509 (N_9509,N_7196,N_7441);
or U9510 (N_9510,N_7846,N_6544);
xor U9511 (N_9511,N_6226,N_7231);
and U9512 (N_9512,N_6666,N_7468);
nor U9513 (N_9513,N_7503,N_7596);
and U9514 (N_9514,N_6298,N_7818);
xor U9515 (N_9515,N_6042,N_6465);
and U9516 (N_9516,N_7034,N_7221);
xor U9517 (N_9517,N_7352,N_6647);
nor U9518 (N_9518,N_7951,N_7007);
or U9519 (N_9519,N_6279,N_7398);
and U9520 (N_9520,N_6344,N_6196);
nor U9521 (N_9521,N_7383,N_7983);
nand U9522 (N_9522,N_6834,N_6909);
nor U9523 (N_9523,N_7402,N_6158);
and U9524 (N_9524,N_6573,N_6394);
xnor U9525 (N_9525,N_7529,N_6387);
and U9526 (N_9526,N_7457,N_6261);
and U9527 (N_9527,N_7638,N_6577);
xor U9528 (N_9528,N_6283,N_7042);
nor U9529 (N_9529,N_6315,N_6896);
xnor U9530 (N_9530,N_6026,N_6742);
nor U9531 (N_9531,N_7979,N_7464);
nand U9532 (N_9532,N_7629,N_7435);
nand U9533 (N_9533,N_7335,N_6145);
xor U9534 (N_9534,N_6021,N_6024);
xnor U9535 (N_9535,N_6992,N_6194);
or U9536 (N_9536,N_7566,N_6962);
xor U9537 (N_9537,N_6985,N_7368);
or U9538 (N_9538,N_7790,N_6963);
xnor U9539 (N_9539,N_6296,N_6857);
nand U9540 (N_9540,N_6582,N_7185);
nand U9541 (N_9541,N_6591,N_7658);
nand U9542 (N_9542,N_6355,N_6561);
or U9543 (N_9543,N_6376,N_6339);
xor U9544 (N_9544,N_6633,N_7408);
and U9545 (N_9545,N_6619,N_6040);
or U9546 (N_9546,N_7443,N_7135);
xnor U9547 (N_9547,N_6275,N_7161);
xor U9548 (N_9548,N_7666,N_6208);
nor U9549 (N_9549,N_7845,N_6053);
xor U9550 (N_9550,N_6446,N_6024);
and U9551 (N_9551,N_7205,N_7329);
nand U9552 (N_9552,N_6373,N_6472);
or U9553 (N_9553,N_7337,N_7573);
xor U9554 (N_9554,N_7750,N_6999);
nand U9555 (N_9555,N_6722,N_7328);
or U9556 (N_9556,N_6128,N_7085);
or U9557 (N_9557,N_7173,N_6264);
nand U9558 (N_9558,N_7194,N_6893);
and U9559 (N_9559,N_7789,N_6999);
nor U9560 (N_9560,N_7120,N_6661);
nor U9561 (N_9561,N_6247,N_6067);
xor U9562 (N_9562,N_7037,N_6023);
xnor U9563 (N_9563,N_6707,N_6064);
nor U9564 (N_9564,N_7621,N_6506);
xnor U9565 (N_9565,N_6832,N_6882);
and U9566 (N_9566,N_7540,N_7013);
or U9567 (N_9567,N_6768,N_6854);
and U9568 (N_9568,N_6287,N_7406);
xor U9569 (N_9569,N_7159,N_6878);
nand U9570 (N_9570,N_6163,N_6444);
nand U9571 (N_9571,N_7904,N_7618);
xor U9572 (N_9572,N_7181,N_6909);
or U9573 (N_9573,N_6482,N_7909);
and U9574 (N_9574,N_7840,N_6588);
and U9575 (N_9575,N_6297,N_6695);
nand U9576 (N_9576,N_7874,N_6944);
or U9577 (N_9577,N_6926,N_7639);
nand U9578 (N_9578,N_7934,N_7498);
or U9579 (N_9579,N_7176,N_6515);
and U9580 (N_9580,N_7649,N_7252);
nand U9581 (N_9581,N_6662,N_6913);
or U9582 (N_9582,N_6077,N_6932);
xor U9583 (N_9583,N_7717,N_7755);
or U9584 (N_9584,N_7202,N_7022);
nand U9585 (N_9585,N_7997,N_7137);
xor U9586 (N_9586,N_6595,N_7540);
or U9587 (N_9587,N_7952,N_6542);
nor U9588 (N_9588,N_7296,N_7266);
and U9589 (N_9589,N_6469,N_7806);
nand U9590 (N_9590,N_7912,N_6684);
nand U9591 (N_9591,N_6550,N_6019);
nor U9592 (N_9592,N_6849,N_6701);
nor U9593 (N_9593,N_6188,N_6048);
or U9594 (N_9594,N_7241,N_6903);
nand U9595 (N_9595,N_7333,N_7096);
nand U9596 (N_9596,N_7798,N_7036);
nand U9597 (N_9597,N_6814,N_6543);
and U9598 (N_9598,N_7841,N_6358);
or U9599 (N_9599,N_7244,N_6254);
or U9600 (N_9600,N_6533,N_7569);
or U9601 (N_9601,N_6584,N_6784);
and U9602 (N_9602,N_7006,N_7081);
xor U9603 (N_9603,N_7381,N_6141);
xor U9604 (N_9604,N_7590,N_6490);
or U9605 (N_9605,N_7212,N_6996);
nand U9606 (N_9606,N_7805,N_7230);
nor U9607 (N_9607,N_7051,N_6401);
xor U9608 (N_9608,N_7400,N_6291);
or U9609 (N_9609,N_7505,N_6089);
nor U9610 (N_9610,N_6404,N_6013);
xor U9611 (N_9611,N_7250,N_6323);
xor U9612 (N_9612,N_6365,N_7998);
or U9613 (N_9613,N_6099,N_6477);
or U9614 (N_9614,N_6820,N_7446);
xnor U9615 (N_9615,N_6637,N_6039);
and U9616 (N_9616,N_6345,N_6321);
xor U9617 (N_9617,N_6811,N_7172);
nor U9618 (N_9618,N_7926,N_6209);
and U9619 (N_9619,N_7596,N_6751);
nor U9620 (N_9620,N_6374,N_7352);
or U9621 (N_9621,N_7220,N_6588);
xor U9622 (N_9622,N_6537,N_6186);
xor U9623 (N_9623,N_6866,N_7348);
or U9624 (N_9624,N_7517,N_6948);
nor U9625 (N_9625,N_7224,N_7251);
nand U9626 (N_9626,N_7952,N_6071);
xnor U9627 (N_9627,N_6569,N_6089);
or U9628 (N_9628,N_6411,N_6937);
xnor U9629 (N_9629,N_6290,N_7704);
nand U9630 (N_9630,N_7142,N_7762);
xor U9631 (N_9631,N_7192,N_7500);
or U9632 (N_9632,N_7529,N_6099);
xor U9633 (N_9633,N_7293,N_6619);
and U9634 (N_9634,N_6266,N_6629);
xor U9635 (N_9635,N_7628,N_6456);
or U9636 (N_9636,N_6294,N_7249);
or U9637 (N_9637,N_6618,N_7643);
or U9638 (N_9638,N_7371,N_7747);
nor U9639 (N_9639,N_6547,N_7779);
nand U9640 (N_9640,N_7187,N_7431);
and U9641 (N_9641,N_6804,N_7682);
and U9642 (N_9642,N_7350,N_6642);
or U9643 (N_9643,N_7118,N_6073);
and U9644 (N_9644,N_7011,N_7874);
nand U9645 (N_9645,N_6079,N_7695);
and U9646 (N_9646,N_6028,N_7764);
nand U9647 (N_9647,N_7267,N_7836);
xor U9648 (N_9648,N_6672,N_6507);
nor U9649 (N_9649,N_7928,N_6073);
nor U9650 (N_9650,N_7110,N_6168);
nand U9651 (N_9651,N_7239,N_7899);
and U9652 (N_9652,N_6266,N_7913);
nor U9653 (N_9653,N_6368,N_7341);
nor U9654 (N_9654,N_6914,N_6050);
or U9655 (N_9655,N_6397,N_7977);
nor U9656 (N_9656,N_7597,N_6493);
and U9657 (N_9657,N_6076,N_6577);
or U9658 (N_9658,N_6459,N_6870);
xnor U9659 (N_9659,N_7004,N_6830);
and U9660 (N_9660,N_6402,N_7512);
xor U9661 (N_9661,N_6871,N_7569);
nand U9662 (N_9662,N_6742,N_6559);
and U9663 (N_9663,N_7965,N_7074);
and U9664 (N_9664,N_7442,N_7560);
xor U9665 (N_9665,N_6985,N_6983);
nand U9666 (N_9666,N_7174,N_7194);
xor U9667 (N_9667,N_6562,N_7960);
xnor U9668 (N_9668,N_7606,N_7535);
nand U9669 (N_9669,N_7522,N_6274);
nor U9670 (N_9670,N_7081,N_6089);
nand U9671 (N_9671,N_6842,N_6852);
or U9672 (N_9672,N_7385,N_6890);
and U9673 (N_9673,N_7140,N_7807);
nor U9674 (N_9674,N_6337,N_7737);
or U9675 (N_9675,N_6827,N_7794);
xor U9676 (N_9676,N_6628,N_6771);
or U9677 (N_9677,N_7057,N_6385);
or U9678 (N_9678,N_6381,N_6304);
or U9679 (N_9679,N_7886,N_7874);
and U9680 (N_9680,N_6256,N_7529);
and U9681 (N_9681,N_6592,N_6519);
nand U9682 (N_9682,N_6669,N_6991);
xnor U9683 (N_9683,N_6332,N_6335);
xor U9684 (N_9684,N_7338,N_6037);
nand U9685 (N_9685,N_6326,N_6123);
or U9686 (N_9686,N_7958,N_6545);
or U9687 (N_9687,N_7895,N_7192);
nand U9688 (N_9688,N_7428,N_6227);
nor U9689 (N_9689,N_7985,N_6722);
or U9690 (N_9690,N_7349,N_7692);
nand U9691 (N_9691,N_7579,N_6607);
or U9692 (N_9692,N_6238,N_7830);
and U9693 (N_9693,N_7899,N_7872);
or U9694 (N_9694,N_7438,N_7939);
nor U9695 (N_9695,N_6650,N_7611);
xnor U9696 (N_9696,N_7639,N_7145);
xor U9697 (N_9697,N_7574,N_7561);
nor U9698 (N_9698,N_7971,N_6987);
nand U9699 (N_9699,N_6995,N_6908);
or U9700 (N_9700,N_6504,N_7509);
nand U9701 (N_9701,N_7829,N_6139);
nand U9702 (N_9702,N_7906,N_6575);
nor U9703 (N_9703,N_7615,N_6751);
xnor U9704 (N_9704,N_6351,N_6930);
and U9705 (N_9705,N_6912,N_6909);
nor U9706 (N_9706,N_6550,N_7672);
nor U9707 (N_9707,N_6195,N_6417);
or U9708 (N_9708,N_6767,N_7990);
nor U9709 (N_9709,N_6794,N_7081);
nand U9710 (N_9710,N_6428,N_7056);
nor U9711 (N_9711,N_7788,N_7853);
xor U9712 (N_9712,N_6668,N_6800);
nor U9713 (N_9713,N_7100,N_7844);
and U9714 (N_9714,N_6633,N_6003);
and U9715 (N_9715,N_7139,N_6848);
and U9716 (N_9716,N_7294,N_7750);
xor U9717 (N_9717,N_7639,N_6902);
and U9718 (N_9718,N_7239,N_6817);
xnor U9719 (N_9719,N_7604,N_7091);
nor U9720 (N_9720,N_6970,N_6446);
or U9721 (N_9721,N_6875,N_7269);
and U9722 (N_9722,N_7405,N_6180);
nor U9723 (N_9723,N_6093,N_6282);
nor U9724 (N_9724,N_6785,N_7841);
xnor U9725 (N_9725,N_6128,N_7247);
nand U9726 (N_9726,N_6643,N_7688);
nor U9727 (N_9727,N_7247,N_6847);
nor U9728 (N_9728,N_6266,N_6894);
nor U9729 (N_9729,N_6052,N_6472);
and U9730 (N_9730,N_6672,N_6069);
nand U9731 (N_9731,N_6926,N_6543);
or U9732 (N_9732,N_6936,N_7668);
and U9733 (N_9733,N_7037,N_7521);
xor U9734 (N_9734,N_7213,N_7511);
and U9735 (N_9735,N_6091,N_6486);
or U9736 (N_9736,N_6799,N_6480);
or U9737 (N_9737,N_7664,N_7232);
or U9738 (N_9738,N_6312,N_7454);
and U9739 (N_9739,N_6472,N_6460);
and U9740 (N_9740,N_6454,N_7533);
nor U9741 (N_9741,N_7507,N_6170);
nor U9742 (N_9742,N_7392,N_6606);
nor U9743 (N_9743,N_6876,N_7152);
xnor U9744 (N_9744,N_7049,N_6066);
nand U9745 (N_9745,N_6899,N_7150);
xnor U9746 (N_9746,N_7018,N_7171);
xor U9747 (N_9747,N_7240,N_6790);
or U9748 (N_9748,N_6028,N_7876);
xnor U9749 (N_9749,N_7134,N_7396);
nand U9750 (N_9750,N_6396,N_7174);
nor U9751 (N_9751,N_7970,N_7384);
nand U9752 (N_9752,N_7878,N_7090);
or U9753 (N_9753,N_6646,N_7344);
nand U9754 (N_9754,N_7466,N_6131);
nand U9755 (N_9755,N_7778,N_6987);
nand U9756 (N_9756,N_7120,N_7459);
and U9757 (N_9757,N_7363,N_7093);
nor U9758 (N_9758,N_6670,N_7508);
nand U9759 (N_9759,N_6682,N_6552);
or U9760 (N_9760,N_6236,N_7191);
and U9761 (N_9761,N_7208,N_7637);
nor U9762 (N_9762,N_6391,N_7500);
xor U9763 (N_9763,N_7877,N_6768);
and U9764 (N_9764,N_7039,N_6973);
or U9765 (N_9765,N_7380,N_7102);
and U9766 (N_9766,N_7883,N_6937);
xnor U9767 (N_9767,N_7666,N_7153);
nand U9768 (N_9768,N_6377,N_6270);
or U9769 (N_9769,N_7182,N_7566);
or U9770 (N_9770,N_6009,N_6017);
and U9771 (N_9771,N_7605,N_7670);
nand U9772 (N_9772,N_7477,N_6893);
nand U9773 (N_9773,N_6287,N_6418);
nor U9774 (N_9774,N_7623,N_7231);
and U9775 (N_9775,N_7178,N_6248);
and U9776 (N_9776,N_6249,N_6138);
nand U9777 (N_9777,N_7281,N_6528);
nand U9778 (N_9778,N_6317,N_6071);
and U9779 (N_9779,N_7569,N_6839);
xor U9780 (N_9780,N_7538,N_6746);
or U9781 (N_9781,N_7043,N_6438);
and U9782 (N_9782,N_6198,N_6694);
nand U9783 (N_9783,N_6099,N_7414);
or U9784 (N_9784,N_6165,N_6096);
and U9785 (N_9785,N_7860,N_6781);
and U9786 (N_9786,N_6528,N_7013);
and U9787 (N_9787,N_6263,N_6897);
nand U9788 (N_9788,N_7031,N_7522);
or U9789 (N_9789,N_6351,N_7120);
nand U9790 (N_9790,N_7712,N_6202);
nor U9791 (N_9791,N_7035,N_6077);
and U9792 (N_9792,N_6575,N_6076);
and U9793 (N_9793,N_6354,N_7120);
nor U9794 (N_9794,N_6641,N_6247);
nor U9795 (N_9795,N_7064,N_7631);
and U9796 (N_9796,N_7291,N_7333);
nand U9797 (N_9797,N_7166,N_6287);
nor U9798 (N_9798,N_6300,N_6041);
and U9799 (N_9799,N_6546,N_7764);
nand U9800 (N_9800,N_7567,N_6776);
and U9801 (N_9801,N_6115,N_6952);
and U9802 (N_9802,N_7099,N_7077);
xnor U9803 (N_9803,N_6393,N_6909);
and U9804 (N_9804,N_7650,N_6875);
or U9805 (N_9805,N_6864,N_6913);
xnor U9806 (N_9806,N_7990,N_7263);
or U9807 (N_9807,N_6694,N_7085);
and U9808 (N_9808,N_7410,N_7863);
xor U9809 (N_9809,N_6832,N_7287);
and U9810 (N_9810,N_6807,N_6549);
and U9811 (N_9811,N_6395,N_6839);
xnor U9812 (N_9812,N_7778,N_7107);
nor U9813 (N_9813,N_7041,N_7790);
nor U9814 (N_9814,N_7195,N_7525);
xnor U9815 (N_9815,N_7964,N_7420);
xnor U9816 (N_9816,N_6672,N_7278);
xnor U9817 (N_9817,N_7362,N_6708);
nor U9818 (N_9818,N_7778,N_6086);
xor U9819 (N_9819,N_6959,N_6554);
nor U9820 (N_9820,N_6070,N_7182);
nor U9821 (N_9821,N_7331,N_7787);
or U9822 (N_9822,N_6667,N_7700);
or U9823 (N_9823,N_7808,N_7941);
nand U9824 (N_9824,N_7796,N_7646);
nand U9825 (N_9825,N_6755,N_7826);
nor U9826 (N_9826,N_7253,N_7224);
xor U9827 (N_9827,N_6157,N_7112);
and U9828 (N_9828,N_7185,N_7436);
or U9829 (N_9829,N_7900,N_6195);
nor U9830 (N_9830,N_7298,N_6010);
nand U9831 (N_9831,N_6778,N_6334);
nand U9832 (N_9832,N_6927,N_6181);
or U9833 (N_9833,N_7306,N_6002);
nand U9834 (N_9834,N_7444,N_6613);
nand U9835 (N_9835,N_6556,N_7173);
nor U9836 (N_9836,N_7156,N_7916);
xor U9837 (N_9837,N_7199,N_7791);
xnor U9838 (N_9838,N_7109,N_6132);
xnor U9839 (N_9839,N_7216,N_6303);
nand U9840 (N_9840,N_6242,N_6927);
xnor U9841 (N_9841,N_6117,N_7280);
nand U9842 (N_9842,N_7850,N_7364);
nand U9843 (N_9843,N_7619,N_6445);
nand U9844 (N_9844,N_7026,N_6322);
xor U9845 (N_9845,N_7812,N_6607);
nand U9846 (N_9846,N_6786,N_7738);
or U9847 (N_9847,N_7084,N_7972);
and U9848 (N_9848,N_7165,N_6113);
xnor U9849 (N_9849,N_7340,N_6279);
xor U9850 (N_9850,N_7556,N_6867);
nand U9851 (N_9851,N_7811,N_6776);
nor U9852 (N_9852,N_6656,N_7984);
and U9853 (N_9853,N_6406,N_7285);
nand U9854 (N_9854,N_7197,N_6910);
or U9855 (N_9855,N_6041,N_7147);
or U9856 (N_9856,N_6771,N_7414);
nand U9857 (N_9857,N_6516,N_6455);
or U9858 (N_9858,N_6744,N_7361);
or U9859 (N_9859,N_6231,N_6670);
or U9860 (N_9860,N_6410,N_7307);
or U9861 (N_9861,N_7960,N_6103);
or U9862 (N_9862,N_7177,N_7702);
nor U9863 (N_9863,N_7241,N_6322);
xnor U9864 (N_9864,N_6649,N_7189);
nor U9865 (N_9865,N_6600,N_7121);
or U9866 (N_9866,N_6543,N_6802);
nor U9867 (N_9867,N_7565,N_7911);
nand U9868 (N_9868,N_7730,N_7239);
nand U9869 (N_9869,N_6804,N_7569);
or U9870 (N_9870,N_6783,N_6060);
nor U9871 (N_9871,N_7537,N_7951);
nor U9872 (N_9872,N_7673,N_7202);
nand U9873 (N_9873,N_6276,N_7681);
nor U9874 (N_9874,N_7854,N_6717);
xor U9875 (N_9875,N_7407,N_7753);
xnor U9876 (N_9876,N_6231,N_7360);
and U9877 (N_9877,N_6092,N_6267);
or U9878 (N_9878,N_7094,N_6232);
or U9879 (N_9879,N_7239,N_6380);
or U9880 (N_9880,N_7233,N_7492);
nand U9881 (N_9881,N_6116,N_7493);
and U9882 (N_9882,N_6973,N_7893);
xnor U9883 (N_9883,N_7834,N_6234);
nand U9884 (N_9884,N_6311,N_7979);
nor U9885 (N_9885,N_6058,N_7096);
nor U9886 (N_9886,N_6126,N_6761);
xor U9887 (N_9887,N_6672,N_6816);
and U9888 (N_9888,N_7799,N_6860);
xor U9889 (N_9889,N_6806,N_6162);
nand U9890 (N_9890,N_7853,N_7272);
nand U9891 (N_9891,N_7199,N_6313);
or U9892 (N_9892,N_6539,N_7240);
or U9893 (N_9893,N_6464,N_6050);
nor U9894 (N_9894,N_7474,N_6407);
or U9895 (N_9895,N_7684,N_7832);
nand U9896 (N_9896,N_7438,N_7789);
nor U9897 (N_9897,N_6357,N_6726);
nor U9898 (N_9898,N_6492,N_7902);
xor U9899 (N_9899,N_6619,N_6447);
xor U9900 (N_9900,N_7621,N_7166);
nand U9901 (N_9901,N_6554,N_6875);
nand U9902 (N_9902,N_7842,N_7129);
nor U9903 (N_9903,N_7907,N_7867);
or U9904 (N_9904,N_7893,N_7353);
xor U9905 (N_9905,N_7660,N_6059);
xor U9906 (N_9906,N_7842,N_6436);
nor U9907 (N_9907,N_6443,N_6372);
and U9908 (N_9908,N_6309,N_6938);
and U9909 (N_9909,N_6491,N_6026);
or U9910 (N_9910,N_6727,N_6822);
nor U9911 (N_9911,N_7624,N_7173);
nand U9912 (N_9912,N_7934,N_6583);
nand U9913 (N_9913,N_7500,N_7450);
nand U9914 (N_9914,N_7968,N_7262);
nor U9915 (N_9915,N_7948,N_7002);
nand U9916 (N_9916,N_6506,N_7301);
and U9917 (N_9917,N_7597,N_7813);
xnor U9918 (N_9918,N_6277,N_7977);
xor U9919 (N_9919,N_7369,N_7640);
nand U9920 (N_9920,N_6368,N_7369);
xnor U9921 (N_9921,N_7956,N_7849);
nand U9922 (N_9922,N_6458,N_6137);
xor U9923 (N_9923,N_6303,N_7922);
and U9924 (N_9924,N_6391,N_6172);
or U9925 (N_9925,N_6834,N_7818);
xnor U9926 (N_9926,N_7258,N_7309);
or U9927 (N_9927,N_7056,N_6556);
and U9928 (N_9928,N_6339,N_7008);
xnor U9929 (N_9929,N_7294,N_6382);
or U9930 (N_9930,N_7237,N_7465);
xor U9931 (N_9931,N_6370,N_7506);
nor U9932 (N_9932,N_7356,N_7589);
and U9933 (N_9933,N_6042,N_6350);
or U9934 (N_9934,N_7610,N_6946);
xor U9935 (N_9935,N_7502,N_7896);
xnor U9936 (N_9936,N_7144,N_6967);
nor U9937 (N_9937,N_7039,N_6914);
or U9938 (N_9938,N_7156,N_6988);
nand U9939 (N_9939,N_6412,N_7149);
or U9940 (N_9940,N_7393,N_6554);
and U9941 (N_9941,N_6631,N_7615);
nor U9942 (N_9942,N_7430,N_7955);
or U9943 (N_9943,N_7131,N_6528);
nor U9944 (N_9944,N_7263,N_7624);
and U9945 (N_9945,N_6606,N_6973);
nand U9946 (N_9946,N_6970,N_6262);
nor U9947 (N_9947,N_6129,N_6621);
xnor U9948 (N_9948,N_7887,N_6449);
or U9949 (N_9949,N_7514,N_7043);
and U9950 (N_9950,N_7958,N_6130);
or U9951 (N_9951,N_6126,N_6121);
or U9952 (N_9952,N_7756,N_6881);
xor U9953 (N_9953,N_7054,N_6819);
nor U9954 (N_9954,N_6262,N_7910);
and U9955 (N_9955,N_7957,N_7683);
nor U9956 (N_9956,N_7715,N_7680);
xor U9957 (N_9957,N_6520,N_7292);
nand U9958 (N_9958,N_6470,N_6817);
nand U9959 (N_9959,N_7219,N_7747);
nor U9960 (N_9960,N_7618,N_7616);
or U9961 (N_9961,N_7239,N_7769);
and U9962 (N_9962,N_7325,N_6158);
and U9963 (N_9963,N_7238,N_7112);
nand U9964 (N_9964,N_6581,N_7071);
xnor U9965 (N_9965,N_6093,N_6558);
xnor U9966 (N_9966,N_7015,N_6837);
xnor U9967 (N_9967,N_7727,N_6104);
and U9968 (N_9968,N_7207,N_7396);
nor U9969 (N_9969,N_6890,N_7393);
or U9970 (N_9970,N_7276,N_6622);
nor U9971 (N_9971,N_6556,N_7350);
and U9972 (N_9972,N_6071,N_6982);
and U9973 (N_9973,N_7084,N_6333);
xor U9974 (N_9974,N_7360,N_7853);
nand U9975 (N_9975,N_7987,N_7220);
and U9976 (N_9976,N_7695,N_7379);
nand U9977 (N_9977,N_7572,N_7399);
and U9978 (N_9978,N_7841,N_6633);
or U9979 (N_9979,N_7143,N_7547);
nand U9980 (N_9980,N_6602,N_7326);
and U9981 (N_9981,N_7614,N_7782);
nand U9982 (N_9982,N_6678,N_6735);
or U9983 (N_9983,N_6335,N_7489);
xor U9984 (N_9984,N_6074,N_7219);
and U9985 (N_9985,N_7255,N_7936);
or U9986 (N_9986,N_7227,N_6448);
or U9987 (N_9987,N_7690,N_6741);
or U9988 (N_9988,N_7177,N_7797);
nand U9989 (N_9989,N_7864,N_7980);
xor U9990 (N_9990,N_7042,N_7212);
nand U9991 (N_9991,N_6139,N_7796);
xnor U9992 (N_9992,N_6774,N_7250);
nand U9993 (N_9993,N_6872,N_6619);
xnor U9994 (N_9994,N_7892,N_7065);
nor U9995 (N_9995,N_7653,N_6487);
and U9996 (N_9996,N_7885,N_6159);
and U9997 (N_9997,N_7620,N_6714);
xor U9998 (N_9998,N_6926,N_6587);
nand U9999 (N_9999,N_7508,N_6292);
xnor UO_0 (O_0,N_9210,N_8851);
xor UO_1 (O_1,N_8173,N_8084);
xor UO_2 (O_2,N_9490,N_8672);
nand UO_3 (O_3,N_8552,N_9574);
and UO_4 (O_4,N_9349,N_9216);
nand UO_5 (O_5,N_9658,N_9491);
or UO_6 (O_6,N_8931,N_9243);
xor UO_7 (O_7,N_8031,N_8721);
or UO_8 (O_8,N_9968,N_8965);
nor UO_9 (O_9,N_8560,N_9733);
or UO_10 (O_10,N_8990,N_8348);
xnor UO_11 (O_11,N_8305,N_8509);
and UO_12 (O_12,N_9386,N_9745);
or UO_13 (O_13,N_9563,N_8239);
or UO_14 (O_14,N_8536,N_9127);
or UO_15 (O_15,N_8630,N_9964);
nand UO_16 (O_16,N_8869,N_9242);
and UO_17 (O_17,N_8880,N_8600);
nand UO_18 (O_18,N_9288,N_9058);
nand UO_19 (O_19,N_9041,N_8397);
or UO_20 (O_20,N_9333,N_8043);
or UO_21 (O_21,N_8484,N_8455);
or UO_22 (O_22,N_9638,N_8820);
and UO_23 (O_23,N_9589,N_8944);
nand UO_24 (O_24,N_8710,N_8553);
nor UO_25 (O_25,N_9517,N_8279);
and UO_26 (O_26,N_9321,N_9759);
nand UO_27 (O_27,N_9047,N_9294);
nand UO_28 (O_28,N_8557,N_9291);
nand UO_29 (O_29,N_8467,N_8951);
nor UO_30 (O_30,N_8138,N_9863);
xnor UO_31 (O_31,N_8409,N_8366);
xor UO_32 (O_32,N_8879,N_9796);
and UO_33 (O_33,N_9159,N_9365);
nand UO_34 (O_34,N_8731,N_9032);
nand UO_35 (O_35,N_8642,N_9656);
xor UO_36 (O_36,N_9650,N_8668);
xnor UO_37 (O_37,N_8817,N_9283);
and UO_38 (O_38,N_8741,N_9318);
nand UO_39 (O_39,N_9847,N_9698);
and UO_40 (O_40,N_8493,N_9154);
and UO_41 (O_41,N_9916,N_8812);
nand UO_42 (O_42,N_8690,N_8208);
xor UO_43 (O_43,N_8250,N_8482);
nand UO_44 (O_44,N_8106,N_9609);
nor UO_45 (O_45,N_9225,N_9987);
xor UO_46 (O_46,N_9409,N_9091);
xnor UO_47 (O_47,N_8027,N_8794);
nor UO_48 (O_48,N_9163,N_9534);
and UO_49 (O_49,N_9930,N_9627);
and UO_50 (O_50,N_9815,N_8524);
or UO_51 (O_51,N_9075,N_9498);
xor UO_52 (O_52,N_8995,N_9814);
nor UO_53 (O_53,N_8922,N_8435);
xnor UO_54 (O_54,N_9871,N_8841);
and UO_55 (O_55,N_8087,N_9469);
nor UO_56 (O_56,N_8015,N_8764);
xnor UO_57 (O_57,N_9794,N_9066);
nand UO_58 (O_58,N_9410,N_9633);
xor UO_59 (O_59,N_9382,N_9808);
and UO_60 (O_60,N_9290,N_9778);
and UO_61 (O_61,N_9246,N_8887);
nand UO_62 (O_62,N_9492,N_8573);
xor UO_63 (O_63,N_8161,N_8178);
or UO_64 (O_64,N_9199,N_8976);
xnor UO_65 (O_65,N_8709,N_8751);
xnor UO_66 (O_66,N_8181,N_9104);
and UO_67 (O_67,N_9599,N_9655);
nand UO_68 (O_68,N_8220,N_9695);
nor UO_69 (O_69,N_8582,N_9859);
nor UO_70 (O_70,N_8842,N_8136);
xnor UO_71 (O_71,N_8507,N_9981);
or UO_72 (O_72,N_8074,N_8960);
xnor UO_73 (O_73,N_8018,N_9311);
nor UO_74 (O_74,N_9430,N_8657);
and UO_75 (O_75,N_8702,N_8481);
nand UO_76 (O_76,N_8913,N_9224);
xor UO_77 (O_77,N_9828,N_9348);
xnor UO_78 (O_78,N_9635,N_8412);
xor UO_79 (O_79,N_8432,N_8007);
and UO_80 (O_80,N_8405,N_9717);
or UO_81 (O_81,N_9683,N_8769);
nand UO_82 (O_82,N_9734,N_9843);
and UO_83 (O_83,N_8378,N_8738);
and UO_84 (O_84,N_8190,N_9353);
and UO_85 (O_85,N_8577,N_8754);
nand UO_86 (O_86,N_8896,N_9173);
nor UO_87 (O_87,N_8195,N_8743);
nor UO_88 (O_88,N_8974,N_8933);
xor UO_89 (O_89,N_8639,N_9878);
xnor UO_90 (O_90,N_8608,N_8050);
nand UO_91 (O_91,N_9821,N_8631);
and UO_92 (O_92,N_9639,N_8997);
and UO_93 (O_93,N_9042,N_9113);
nor UO_94 (O_94,N_9699,N_8230);
nand UO_95 (O_95,N_9014,N_8473);
nand UO_96 (O_96,N_9720,N_9152);
xor UO_97 (O_97,N_9258,N_8009);
xnor UO_98 (O_98,N_8616,N_9943);
and UO_99 (O_99,N_8285,N_9284);
or UO_100 (O_100,N_9615,N_8391);
or UO_101 (O_101,N_8717,N_9007);
xor UO_102 (O_102,N_8110,N_9835);
and UO_103 (O_103,N_8541,N_9438);
xor UO_104 (O_104,N_9631,N_8989);
nand UO_105 (O_105,N_8924,N_8908);
nor UO_106 (O_106,N_9562,N_8946);
nor UO_107 (O_107,N_8016,N_8568);
xnor UO_108 (O_108,N_8058,N_8936);
or UO_109 (O_109,N_9372,N_8164);
and UO_110 (O_110,N_8094,N_8329);
nand UO_111 (O_111,N_8749,N_8238);
and UO_112 (O_112,N_9568,N_9391);
nor UO_113 (O_113,N_8450,N_9144);
nor UO_114 (O_114,N_8893,N_8975);
xor UO_115 (O_115,N_9207,N_8677);
nor UO_116 (O_116,N_9221,N_9415);
nor UO_117 (O_117,N_9328,N_9025);
nor UO_118 (O_118,N_9165,N_9545);
nand UO_119 (O_119,N_9933,N_9706);
xor UO_120 (O_120,N_8014,N_9062);
nor UO_121 (O_121,N_9011,N_8440);
or UO_122 (O_122,N_9716,N_8884);
xor UO_123 (O_123,N_8638,N_8872);
nor UO_124 (O_124,N_9952,N_8692);
and UO_125 (O_125,N_8961,N_9023);
nor UO_126 (O_126,N_8765,N_9684);
nand UO_127 (O_127,N_8747,N_9966);
nand UO_128 (O_128,N_8888,N_9806);
and UO_129 (O_129,N_9595,N_9335);
xnor UO_130 (O_130,N_9279,N_9145);
xor UO_131 (O_131,N_8000,N_8904);
nand UO_132 (O_132,N_9974,N_9621);
xor UO_133 (O_133,N_8411,N_8874);
or UO_134 (O_134,N_8514,N_8126);
nor UO_135 (O_135,N_9577,N_9571);
and UO_136 (O_136,N_9485,N_9915);
nand UO_137 (O_137,N_8760,N_8711);
xor UO_138 (O_138,N_9670,N_8495);
xor UO_139 (O_139,N_9949,N_9886);
nor UO_140 (O_140,N_8948,N_8732);
xor UO_141 (O_141,N_9269,N_9676);
nor UO_142 (O_142,N_8092,N_8388);
xnor UO_143 (O_143,N_9422,N_9924);
xnor UO_144 (O_144,N_8984,N_9565);
nor UO_145 (O_145,N_8898,N_9158);
and UO_146 (O_146,N_9929,N_8627);
nand UO_147 (O_147,N_8927,N_9682);
xor UO_148 (O_148,N_9377,N_9728);
nand UO_149 (O_149,N_8648,N_9412);
or UO_150 (O_150,N_8301,N_8459);
nand UO_151 (O_151,N_9687,N_9640);
nor UO_152 (O_152,N_8847,N_8501);
nand UO_153 (O_153,N_9337,N_9746);
and UO_154 (O_154,N_8623,N_9593);
nor UO_155 (O_155,N_8362,N_8371);
xnor UO_156 (O_156,N_8112,N_9866);
nor UO_157 (O_157,N_9921,N_9844);
and UO_158 (O_158,N_8271,N_9555);
and UO_159 (O_159,N_8011,N_8605);
xor UO_160 (O_160,N_8035,N_8601);
nor UO_161 (O_161,N_9157,N_9510);
and UO_162 (O_162,N_8912,N_9895);
or UO_163 (O_163,N_9162,N_8032);
nor UO_164 (O_164,N_8477,N_8263);
or UO_165 (O_165,N_9786,N_8308);
nor UO_166 (O_166,N_9505,N_8671);
xor UO_167 (O_167,N_9250,N_9537);
and UO_168 (O_168,N_8920,N_8347);
xor UO_169 (O_169,N_9692,N_9525);
xnor UO_170 (O_170,N_9230,N_9087);
nand UO_171 (O_171,N_8448,N_9740);
nand UO_172 (O_172,N_8380,N_9013);
or UO_173 (O_173,N_8428,N_8527);
and UO_174 (O_174,N_8996,N_9125);
or UO_175 (O_175,N_8585,N_9553);
nand UO_176 (O_176,N_9742,N_8615);
or UO_177 (O_177,N_9265,N_8039);
nor UO_178 (O_178,N_8590,N_9499);
nand UO_179 (O_179,N_8186,N_9596);
and UO_180 (O_180,N_9834,N_9601);
or UO_181 (O_181,N_8217,N_8352);
nor UO_182 (O_182,N_8068,N_8938);
nand UO_183 (O_183,N_8449,N_9198);
or UO_184 (O_184,N_8252,N_9248);
nand UO_185 (O_185,N_9227,N_9030);
nand UO_186 (O_186,N_8592,N_8024);
and UO_187 (O_187,N_9089,N_9097);
and UO_188 (O_188,N_9592,N_9881);
nor UO_189 (O_189,N_9167,N_9050);
and UO_190 (O_190,N_8158,N_8580);
nand UO_191 (O_191,N_8002,N_8237);
and UO_192 (O_192,N_8107,N_9347);
nand UO_193 (O_193,N_9793,N_8926);
xnor UO_194 (O_194,N_8859,N_8082);
nor UO_195 (O_195,N_8444,N_8656);
xor UO_196 (O_196,N_8205,N_8534);
nand UO_197 (O_197,N_9925,N_9252);
nor UO_198 (O_198,N_9208,N_9186);
nor UO_199 (O_199,N_8101,N_9938);
and UO_200 (O_200,N_8276,N_9940);
and UO_201 (O_201,N_8456,N_8579);
xor UO_202 (O_202,N_8641,N_8515);
and UO_203 (O_203,N_8850,N_9885);
nand UO_204 (O_204,N_8624,N_9824);
nand UO_205 (O_205,N_9332,N_9857);
nor UO_206 (O_206,N_8393,N_8613);
nand UO_207 (O_207,N_8664,N_9823);
or UO_208 (O_208,N_8153,N_9777);
nand UO_209 (O_209,N_8610,N_9033);
and UO_210 (O_210,N_9061,N_9632);
nand UO_211 (O_211,N_8273,N_9253);
or UO_212 (O_212,N_8211,N_9643);
or UO_213 (O_213,N_8375,N_9722);
and UO_214 (O_214,N_8962,N_9953);
nand UO_215 (O_215,N_8376,N_9573);
and UO_216 (O_216,N_8445,N_8742);
or UO_217 (O_217,N_9504,N_9898);
or UO_218 (O_218,N_8785,N_8401);
nor UO_219 (O_219,N_8422,N_8958);
nor UO_220 (O_220,N_8537,N_9416);
nor UO_221 (O_221,N_9705,N_8017);
nor UO_222 (O_222,N_9018,N_9664);
nor UO_223 (O_223,N_9942,N_9889);
nor UO_224 (O_224,N_8360,N_9143);
or UO_225 (O_225,N_8013,N_8629);
nand UO_226 (O_226,N_9045,N_8978);
xor UO_227 (O_227,N_8602,N_8538);
or UO_228 (O_228,N_9111,N_9544);
nand UO_229 (O_229,N_8198,N_8871);
xnor UO_230 (O_230,N_9791,N_8681);
xnor UO_231 (O_231,N_8303,N_8191);
nand UO_232 (O_232,N_9527,N_8703);
and UO_233 (O_233,N_8089,N_9249);
nor UO_234 (O_234,N_8245,N_8950);
nor UO_235 (O_235,N_9182,N_8523);
nand UO_236 (O_236,N_8877,N_8584);
nor UO_237 (O_237,N_8992,N_9865);
or UO_238 (O_238,N_9926,N_8081);
or UO_239 (O_239,N_9972,N_8798);
and UO_240 (O_240,N_8634,N_8522);
or UO_241 (O_241,N_9897,N_8121);
nor UO_242 (O_242,N_9479,N_9219);
or UO_243 (O_243,N_8223,N_8102);
and UO_244 (O_244,N_8932,N_8146);
or UO_245 (O_245,N_9827,N_8241);
xor UO_246 (O_246,N_9368,N_8183);
nor UO_247 (O_247,N_8564,N_9356);
xnor UO_248 (O_248,N_8588,N_9081);
and UO_249 (O_249,N_8963,N_9647);
and UO_250 (O_250,N_8581,N_9489);
or UO_251 (O_251,N_9467,N_8296);
nor UO_252 (O_252,N_9825,N_9059);
nand UO_253 (O_253,N_8790,N_9994);
xnor UO_254 (O_254,N_9095,N_9241);
nand UO_255 (O_255,N_9969,N_8521);
xor UO_256 (O_256,N_9551,N_8511);
or UO_257 (O_257,N_8162,N_9206);
nor UO_258 (O_258,N_8647,N_9472);
nand UO_259 (O_259,N_8465,N_8586);
and UO_260 (O_260,N_9122,N_9400);
xnor UO_261 (O_261,N_8175,N_8057);
or UO_262 (O_262,N_8650,N_8559);
nor UO_263 (O_263,N_9043,N_9932);
or UO_264 (O_264,N_9585,N_9539);
and UO_265 (O_265,N_8715,N_9912);
and UO_266 (O_266,N_8185,N_8189);
xor UO_267 (O_267,N_8621,N_8326);
xor UO_268 (O_268,N_9166,N_8384);
xor UO_269 (O_269,N_8775,N_9550);
nand UO_270 (O_270,N_9285,N_8349);
nand UO_271 (O_271,N_9278,N_8012);
nand UO_272 (O_272,N_8254,N_9121);
xnor UO_273 (O_273,N_8680,N_9255);
nand UO_274 (O_274,N_8818,N_8070);
and UO_275 (O_275,N_8073,N_9329);
or UO_276 (O_276,N_9299,N_8921);
xor UO_277 (O_277,N_8260,N_9024);
nor UO_278 (O_278,N_8076,N_9607);
or UO_279 (O_279,N_9836,N_9986);
or UO_280 (O_280,N_9419,N_8845);
nand UO_281 (O_281,N_9977,N_8314);
nand UO_282 (O_282,N_8519,N_8782);
nor UO_283 (O_283,N_9080,N_9101);
xnor UO_284 (O_284,N_8339,N_9297);
nand UO_285 (O_285,N_8404,N_9567);
xor UO_286 (O_286,N_9098,N_9507);
and UO_287 (O_287,N_8891,N_9137);
or UO_288 (O_288,N_8508,N_8953);
nor UO_289 (O_289,N_9213,N_8735);
and UO_290 (O_290,N_9390,N_8870);
xor UO_291 (O_291,N_8774,N_9894);
xnor UO_292 (O_292,N_8226,N_8460);
and UO_293 (O_293,N_8619,N_8103);
nand UO_294 (O_294,N_9948,N_9106);
and UO_295 (O_295,N_8443,N_8335);
nand UO_296 (O_296,N_9183,N_9939);
xor UO_297 (O_297,N_8159,N_8095);
or UO_298 (O_298,N_9584,N_9135);
nor UO_299 (O_299,N_9523,N_9092);
xor UO_300 (O_300,N_8665,N_9339);
xnor UO_301 (O_301,N_8278,N_9147);
xor UO_302 (O_302,N_8838,N_8750);
nor UO_303 (O_303,N_8867,N_8799);
or UO_304 (O_304,N_8868,N_8202);
and UO_305 (O_305,N_8048,N_9096);
nor UO_306 (O_306,N_9292,N_8340);
xor UO_307 (O_307,N_8122,N_9447);
nand UO_308 (O_308,N_9396,N_9070);
xor UO_309 (O_309,N_9362,N_8029);
and UO_310 (O_310,N_9179,N_8117);
or UO_311 (O_311,N_9341,N_8288);
nor UO_312 (O_312,N_8909,N_9302);
xnor UO_313 (O_313,N_8609,N_8474);
nand UO_314 (O_314,N_9355,N_9375);
and UO_315 (O_315,N_8718,N_9501);
or UO_316 (O_316,N_8398,N_9532);
or UO_317 (O_317,N_8632,N_9945);
and UO_318 (O_318,N_9457,N_9420);
xnor UO_319 (O_319,N_8414,N_9840);
nand UO_320 (O_320,N_8611,N_9558);
nand UO_321 (O_321,N_8430,N_8575);
nand UO_322 (O_322,N_9067,N_8292);
nand UO_323 (O_323,N_8485,N_8020);
nand UO_324 (O_324,N_9211,N_9231);
and UO_325 (O_325,N_9768,N_9579);
and UO_326 (O_326,N_9012,N_9275);
or UO_327 (O_327,N_8172,N_9962);
nand UO_328 (O_328,N_9813,N_9869);
and UO_329 (O_329,N_8895,N_8255);
and UO_330 (O_330,N_8529,N_9784);
xor UO_331 (O_331,N_9244,N_8167);
xor UO_332 (O_332,N_8256,N_9277);
nor UO_333 (O_333,N_9618,N_8476);
and UO_334 (O_334,N_9662,N_8346);
and UO_335 (O_335,N_8821,N_9854);
or UO_336 (O_336,N_8816,N_8767);
and UO_337 (O_337,N_8480,N_8293);
or UO_338 (O_338,N_8688,N_8496);
nor UO_339 (O_339,N_8802,N_8667);
nor UO_340 (O_340,N_9588,N_8780);
and UO_341 (O_341,N_8216,N_8746);
or UO_342 (O_342,N_8287,N_8119);
nor UO_343 (O_343,N_8558,N_8986);
nand UO_344 (O_344,N_8993,N_9956);
and UO_345 (O_345,N_9471,N_9270);
and UO_346 (O_346,N_9910,N_9760);
and UO_347 (O_347,N_8547,N_9016);
nor UO_348 (O_348,N_9659,N_8655);
xor UO_349 (O_349,N_9456,N_9223);
nand UO_350 (O_350,N_8531,N_8377);
and UO_351 (O_351,N_9819,N_9273);
and UO_352 (O_352,N_8885,N_8180);
nor UO_353 (O_353,N_8199,N_9102);
nor UO_354 (O_354,N_8118,N_9373);
xor UO_355 (O_355,N_9606,N_9730);
and UO_356 (O_356,N_9330,N_8160);
or UO_357 (O_357,N_8759,N_8155);
or UO_358 (O_358,N_8135,N_8115);
and UO_359 (O_359,N_9319,N_8298);
nand UO_360 (O_360,N_9963,N_8056);
nand UO_361 (O_361,N_9718,N_9837);
nor UO_362 (O_362,N_8691,N_9913);
nor UO_363 (O_363,N_9392,N_8415);
xor UO_364 (O_364,N_9268,N_9694);
xnor UO_365 (O_365,N_9502,N_9473);
or UO_366 (O_366,N_8442,N_9460);
xnor UO_367 (O_367,N_9315,N_9078);
nor UO_368 (O_368,N_9514,N_8971);
nand UO_369 (O_369,N_9090,N_8807);
and UO_370 (O_370,N_9531,N_8261);
or UO_371 (O_371,N_9641,N_9201);
nand UO_372 (O_372,N_9437,N_9264);
nor UO_373 (O_373,N_9425,N_9947);
nor UO_374 (O_374,N_9801,N_9452);
or UO_375 (O_375,N_8144,N_9237);
nor UO_376 (O_376,N_9406,N_8684);
nand UO_377 (O_377,N_8025,N_8355);
nor UO_378 (O_378,N_8008,N_8518);
and UO_379 (O_379,N_9529,N_8045);
or UO_380 (O_380,N_8637,N_8959);
xor UO_381 (O_381,N_8041,N_9161);
xnor UO_382 (O_382,N_9338,N_9494);
nor UO_383 (O_383,N_9423,N_9436);
nand UO_384 (O_384,N_8436,N_8351);
xnor UO_385 (O_385,N_9669,N_9172);
or UO_386 (O_386,N_8307,N_8096);
nor UO_387 (O_387,N_9623,N_9667);
nor UO_388 (O_388,N_9779,N_8317);
xnor UO_389 (O_389,N_8733,N_9557);
xor UO_390 (O_390,N_9446,N_8291);
xor UO_391 (O_391,N_8756,N_9240);
and UO_392 (O_392,N_9838,N_8367);
or UO_393 (O_393,N_8973,N_8855);
and UO_394 (O_394,N_8725,N_9262);
or UO_395 (O_395,N_9772,N_8427);
and UO_396 (O_396,N_9310,N_8517);
nor UO_397 (O_397,N_8860,N_8801);
and UO_398 (O_398,N_9345,N_8899);
and UO_399 (O_399,N_9766,N_9247);
nand UO_400 (O_400,N_9732,N_8614);
and UO_401 (O_401,N_8707,N_9620);
and UO_402 (O_402,N_9470,N_8979);
nor UO_403 (O_403,N_9927,N_9475);
and UO_404 (O_404,N_9116,N_8528);
nand UO_405 (O_405,N_8942,N_9378);
nor UO_406 (O_406,N_8694,N_8693);
nor UO_407 (O_407,N_8370,N_8535);
nand UO_408 (O_408,N_9578,N_9086);
nand UO_409 (O_409,N_9336,N_8005);
or UO_410 (O_410,N_8257,N_8341);
or UO_411 (O_411,N_8532,N_9903);
nand UO_412 (O_412,N_8969,N_8666);
xor UO_413 (O_413,N_8416,N_9399);
nand UO_414 (O_414,N_8597,N_8643);
nor UO_415 (O_415,N_9902,N_8354);
and UO_416 (O_416,N_8247,N_9281);
and UO_417 (O_417,N_8669,N_8359);
xnor UO_418 (O_418,N_8776,N_8977);
nand UO_419 (O_419,N_8419,N_8569);
or UO_420 (O_420,N_9461,N_9380);
nand UO_421 (O_421,N_9342,N_9996);
or UO_422 (O_422,N_9990,N_9988);
nand UO_423 (O_423,N_8266,N_9203);
or UO_424 (O_424,N_9508,N_8897);
nand UO_425 (O_425,N_9710,N_8026);
xnor UO_426 (O_426,N_9905,N_9833);
xor UO_427 (O_427,N_9123,N_9549);
xnor UO_428 (O_428,N_8830,N_8343);
or UO_429 (O_429,N_9068,N_9830);
and UO_430 (O_430,N_9858,N_9055);
nor UO_431 (O_431,N_9958,N_9919);
nor UO_432 (O_432,N_8406,N_9254);
or UO_433 (O_433,N_8502,N_8574);
or UO_434 (O_434,N_9477,N_8210);
or UO_435 (O_435,N_9747,N_9880);
and UO_436 (O_436,N_8131,N_8678);
xor UO_437 (O_437,N_9598,N_9628);
nor UO_438 (O_438,N_8383,N_8545);
nand UO_439 (O_439,N_8654,N_9130);
xor UO_440 (O_440,N_8964,N_8163);
nor UO_441 (O_441,N_9564,N_8345);
or UO_442 (O_442,N_8636,N_9600);
xor UO_443 (O_443,N_9352,N_8299);
or UO_444 (O_444,N_9992,N_9293);
nand UO_445 (O_445,N_8593,N_9190);
or UO_446 (O_446,N_9999,N_8652);
or UO_447 (O_447,N_8934,N_8395);
or UO_448 (O_448,N_9884,N_8651);
or UO_449 (O_449,N_8300,N_9176);
nand UO_450 (O_450,N_8224,N_8734);
and UO_451 (O_451,N_8396,N_9160);
nor UO_452 (O_452,N_9286,N_8941);
or UO_453 (O_453,N_9364,N_9757);
nand UO_454 (O_454,N_8201,N_9465);
and UO_455 (O_455,N_9637,N_9580);
nor UO_456 (O_456,N_9431,N_9217);
nand UO_457 (O_457,N_9222,N_9171);
nor UO_458 (O_458,N_8748,N_8104);
nand UO_459 (O_459,N_9358,N_9961);
or UO_460 (O_460,N_8374,N_9181);
and UO_461 (O_461,N_9497,N_8188);
nand UO_462 (O_462,N_8753,N_9155);
nor UO_463 (O_463,N_8628,N_9862);
xnor UO_464 (O_464,N_8695,N_8361);
or UO_465 (O_465,N_9448,N_8686);
or UO_466 (O_466,N_8204,N_8849);
or UO_467 (O_467,N_8433,N_8203);
or UO_468 (O_468,N_9308,N_9737);
and UO_469 (O_469,N_8572,N_8272);
xnor UO_470 (O_470,N_9085,N_9401);
and UO_471 (O_471,N_9770,N_8848);
nor UO_472 (O_472,N_8333,N_9424);
nor UO_473 (O_473,N_9094,N_9194);
or UO_474 (O_474,N_9516,N_9148);
nand UO_475 (O_475,N_9538,N_8679);
nand UO_476 (O_476,N_9729,N_9752);
or UO_477 (O_477,N_9707,N_9561);
or UO_478 (O_478,N_8108,N_8730);
nand UO_479 (O_479,N_8399,N_9177);
nand UO_480 (O_480,N_8022,N_8434);
nand UO_481 (O_481,N_9822,N_9530);
nor UO_482 (O_482,N_9381,N_8566);
nand UO_483 (O_483,N_9180,N_8806);
and UO_484 (O_484,N_9887,N_9374);
xor UO_485 (O_485,N_9367,N_9481);
nor UO_486 (O_486,N_8423,N_9139);
nand UO_487 (O_487,N_8808,N_9914);
nand UO_488 (O_488,N_9559,N_9560);
nand UO_489 (O_489,N_8021,N_8353);
and UO_490 (O_490,N_9371,N_8661);
or UO_491 (O_491,N_8833,N_8745);
or UO_492 (O_492,N_9946,N_9957);
and UO_493 (O_493,N_9168,N_9918);
or UO_494 (O_494,N_9389,N_9893);
nor UO_495 (O_495,N_8892,N_9524);
or UO_496 (O_496,N_9883,N_8789);
or UO_497 (O_497,N_9856,N_9326);
nor UO_498 (O_498,N_8525,N_8133);
nor UO_499 (O_499,N_8170,N_9625);
nor UO_500 (O_500,N_9022,N_9556);
nor UO_501 (O_501,N_8994,N_9788);
or UO_502 (O_502,N_8494,N_9877);
nand UO_503 (O_503,N_9074,N_9570);
xor UO_504 (O_504,N_9785,N_9196);
nand UO_505 (O_505,N_9088,N_9802);
and UO_506 (O_506,N_9109,N_9581);
nor UO_507 (O_507,N_8506,N_9280);
and UO_508 (O_508,N_9651,N_9408);
nor UO_509 (O_509,N_8381,N_9636);
nand UO_510 (O_510,N_8334,N_9008);
nand UO_511 (O_511,N_9287,N_9892);
nand UO_512 (O_512,N_8906,N_8386);
and UO_513 (O_513,N_9936,N_8275);
xnor UO_514 (O_514,N_9873,N_8457);
and UO_515 (O_515,N_9804,N_8283);
and UO_516 (O_516,N_9513,N_9758);
xnor UO_517 (O_517,N_8093,N_8675);
nor UO_518 (O_518,N_9439,N_8479);
nor UO_519 (O_519,N_8097,N_8179);
xnor UO_520 (O_520,N_8246,N_8379);
nor UO_521 (O_521,N_8497,N_8947);
nor UO_522 (O_522,N_8327,N_9002);
nor UO_523 (O_523,N_8319,N_9079);
nor UO_524 (O_524,N_9959,N_8949);
or UO_525 (O_525,N_9433,N_8856);
nor UO_526 (O_526,N_8954,N_8392);
and UO_527 (O_527,N_9764,N_8689);
and UO_528 (O_528,N_9259,N_9313);
or UO_529 (O_529,N_8023,N_8171);
or UO_530 (O_530,N_9239,N_8510);
nor UO_531 (O_531,N_9140,N_9672);
nor UO_532 (O_532,N_8622,N_8083);
or UO_533 (O_533,N_8085,N_9001);
nand UO_534 (O_534,N_9861,N_9027);
or UO_535 (O_535,N_8065,N_8649);
or UO_536 (O_536,N_9762,N_9402);
nand UO_537 (O_537,N_8797,N_9039);
nor UO_538 (O_538,N_8864,N_9187);
xnor UO_539 (O_539,N_9282,N_8685);
and UO_540 (O_540,N_9741,N_9646);
nor UO_541 (O_541,N_9346,N_8955);
xor UO_542 (O_542,N_8981,N_8036);
nor UO_543 (O_543,N_9935,N_9769);
nand UO_544 (O_544,N_9920,N_8154);
or UO_545 (O_545,N_9476,N_9681);
nand UO_546 (O_546,N_8736,N_9937);
nor UO_547 (O_547,N_8713,N_9124);
nand UO_548 (O_548,N_9874,N_9693);
xor UO_549 (O_549,N_8727,N_9413);
nand UO_550 (O_550,N_8596,N_9724);
nand UO_551 (O_551,N_9051,N_8533);
or UO_552 (O_552,N_8516,N_9543);
and UO_553 (O_553,N_9626,N_9985);
nor UO_554 (O_554,N_8583,N_9351);
xor UO_555 (O_555,N_9750,N_8321);
nor UO_556 (O_556,N_9115,N_9496);
or UO_557 (O_557,N_8504,N_8242);
and UO_558 (O_558,N_8132,N_8209);
nor UO_559 (O_559,N_8222,N_8090);
and UO_560 (O_560,N_9979,N_8620);
and UO_561 (O_561,N_9468,N_9185);
xor UO_562 (O_562,N_9980,N_9323);
nand UO_563 (O_563,N_8463,N_8796);
or UO_564 (O_564,N_8957,N_8843);
nor UO_565 (O_565,N_9376,N_8852);
xor UO_566 (O_566,N_8324,N_8044);
nor UO_567 (O_567,N_8064,N_8269);
nand UO_568 (O_568,N_9576,N_9711);
nand UO_569 (O_569,N_9083,N_9817);
xor UO_570 (O_570,N_8724,N_9169);
and UO_571 (O_571,N_8792,N_9960);
and UO_572 (O_572,N_8723,N_8387);
nand UO_573 (O_573,N_8439,N_9775);
nand UO_574 (O_574,N_8311,N_9385);
or UO_575 (O_575,N_9810,N_8910);
and UO_576 (O_576,N_8196,N_8441);
or UO_577 (O_577,N_9407,N_8914);
and UO_578 (O_578,N_9427,N_9228);
xnor UO_579 (O_579,N_9663,N_8421);
nand UO_580 (O_580,N_9404,N_8499);
xnor UO_581 (O_581,N_8778,N_9726);
and UO_582 (O_582,N_8111,N_9434);
xor UO_583 (O_583,N_8901,N_8653);
nand UO_584 (O_584,N_9276,N_9798);
nand UO_585 (O_585,N_8229,N_8635);
and UO_586 (O_586,N_9232,N_8739);
and UO_587 (O_587,N_9590,N_9028);
and UO_588 (O_588,N_9005,N_8078);
xnor UO_589 (O_589,N_8069,N_8846);
or UO_590 (O_590,N_8673,N_9369);
and UO_591 (O_591,N_8310,N_9444);
and UO_592 (O_592,N_8309,N_8915);
nor UO_593 (O_593,N_8565,N_8067);
nor UO_594 (O_594,N_8157,N_9675);
xor UO_595 (O_595,N_8490,N_9677);
nand UO_596 (O_596,N_9679,N_8325);
nand UO_597 (O_597,N_8062,N_8322);
xor UO_598 (O_598,N_9809,N_9383);
and UO_599 (O_599,N_9361,N_9755);
nand UO_600 (O_600,N_9509,N_8289);
or UO_601 (O_601,N_9105,N_8251);
or UO_602 (O_602,N_9872,N_9435);
xor UO_603 (O_603,N_8454,N_9701);
and UO_604 (O_604,N_8267,N_9583);
or UO_605 (O_605,N_9660,N_9214);
nor UO_606 (O_606,N_8706,N_9212);
nand UO_607 (O_607,N_9860,N_8489);
or UO_608 (O_608,N_8052,N_9709);
nand UO_609 (O_609,N_8676,N_8207);
or UO_610 (O_610,N_8771,N_9440);
nand UO_611 (O_611,N_8244,N_9831);
nor UO_612 (O_612,N_8972,N_9774);
xnor UO_613 (O_613,N_9845,N_8576);
nand UO_614 (O_614,N_9132,N_8174);
nor UO_615 (O_615,N_8861,N_9998);
nor UO_616 (O_616,N_9056,N_8998);
or UO_617 (O_617,N_8233,N_8814);
nor UO_618 (O_618,N_9046,N_8758);
and UO_619 (O_619,N_8766,N_8281);
xor UO_620 (O_620,N_9944,N_9799);
xor UO_621 (O_621,N_9503,N_8918);
or UO_622 (O_622,N_8822,N_9429);
xnor UO_623 (O_623,N_8687,N_8231);
nand UO_624 (O_624,N_9129,N_8858);
and UO_625 (O_625,N_9907,N_9614);
xnor UO_626 (O_626,N_9756,N_9487);
nand UO_627 (O_627,N_8786,N_8030);
nor UO_628 (O_628,N_9432,N_8755);
nor UO_629 (O_629,N_9515,N_9820);
nand UO_630 (O_630,N_8492,N_9552);
and UO_631 (O_631,N_8645,N_9455);
nand UO_632 (O_632,N_9266,N_9417);
xor UO_633 (O_633,N_9015,N_9783);
and UO_634 (O_634,N_8530,N_9715);
nor UO_635 (O_635,N_8491,N_8249);
nor UO_636 (O_636,N_8332,N_8453);
xor UO_637 (O_637,N_9305,N_8350);
xnor UO_638 (O_638,N_8046,N_9586);
xnor UO_639 (O_639,N_8452,N_9405);
nor UO_640 (O_640,N_8520,N_8033);
or UO_641 (O_641,N_9108,N_9849);
or UO_642 (O_642,N_8834,N_9773);
or UO_643 (O_643,N_8570,N_9688);
nor UO_644 (O_644,N_9941,N_8660);
nor UO_645 (O_645,N_8825,N_8197);
nand UO_646 (O_646,N_8890,N_8149);
or UO_647 (O_647,N_8952,N_9653);
xor UO_648 (O_648,N_9616,N_8342);
or UO_649 (O_649,N_8987,N_8227);
nor UO_650 (O_650,N_8968,N_8280);
nand UO_651 (O_651,N_9119,N_9792);
nor UO_652 (O_652,N_9816,N_8072);
nor UO_653 (O_653,N_8900,N_9781);
nor UO_654 (O_654,N_8988,N_9521);
or UO_655 (O_655,N_8889,N_8318);
nor UO_656 (O_656,N_9993,N_9622);
xor UO_657 (O_657,N_8218,N_8554);
and UO_658 (O_658,N_9118,N_9500);
xnor UO_659 (O_659,N_9909,N_9800);
nand UO_660 (O_660,N_9697,N_9142);
nand UO_661 (O_661,N_8768,N_9582);
and UO_662 (O_662,N_8763,N_8779);
or UO_663 (O_663,N_9754,N_9876);
nor UO_664 (O_664,N_9184,N_8143);
nand UO_665 (O_665,N_8040,N_8147);
and UO_666 (O_666,N_8356,N_9174);
or UO_667 (O_667,N_9057,N_8129);
xnor UO_668 (O_668,N_9360,N_9256);
nand UO_669 (O_669,N_9542,N_8956);
nand UO_670 (O_670,N_9665,N_9065);
or UO_671 (O_671,N_9411,N_8700);
xor UO_672 (O_672,N_9950,N_8930);
xor UO_673 (O_673,N_9736,N_9261);
or UO_674 (O_674,N_8417,N_9767);
nor UO_675 (O_675,N_9236,N_9850);
and UO_676 (O_676,N_9976,N_8983);
nor UO_677 (O_677,N_8705,N_8099);
and UO_678 (O_678,N_9797,N_8823);
nand UO_679 (O_679,N_8865,N_9634);
xor UO_680 (O_680,N_9170,N_9719);
or UO_681 (O_681,N_9188,N_8470);
and UO_682 (O_682,N_8625,N_8633);
nand UO_683 (O_683,N_9234,N_8589);
and UO_684 (O_684,N_8562,N_8028);
nor UO_685 (O_685,N_8809,N_8606);
or UO_686 (O_686,N_8312,N_9393);
xor UO_687 (O_687,N_8402,N_8438);
xor UO_688 (O_688,N_8290,N_8004);
nand UO_689 (O_689,N_9594,N_9686);
xnor UO_690 (O_690,N_8603,N_8148);
and UO_691 (O_691,N_8382,N_9610);
nand UO_692 (O_692,N_9666,N_8425);
nor UO_693 (O_693,N_9989,N_8169);
nor UO_694 (O_694,N_8811,N_8328);
and UO_695 (O_695,N_8461,N_9605);
xor UO_696 (O_696,N_9739,N_8446);
and UO_697 (O_697,N_8001,N_9748);
and UO_698 (O_698,N_8712,N_9548);
nor UO_699 (O_699,N_8253,N_9478);
and UO_700 (O_700,N_8682,N_9309);
or UO_701 (O_701,N_8793,N_8591);
or UO_702 (O_702,N_8683,N_8408);
and UO_703 (O_703,N_8152,N_9604);
xnor UO_704 (O_704,N_8835,N_8800);
xor UO_705 (O_705,N_8182,N_9029);
and UO_706 (O_706,N_8128,N_8478);
nand UO_707 (O_707,N_8815,N_9908);
nand UO_708 (O_708,N_8612,N_8003);
xnor UO_709 (O_709,N_8192,N_8394);
xnor UO_710 (O_710,N_8038,N_9395);
nor UO_711 (O_711,N_9839,N_8221);
and UO_712 (O_712,N_8599,N_9483);
xor UO_713 (O_713,N_9100,N_9536);
or UO_714 (O_714,N_9441,N_9818);
xnor UO_715 (O_715,N_9704,N_8471);
and UO_716 (O_716,N_8086,N_9126);
and UO_717 (O_717,N_9891,N_9303);
and UO_718 (O_718,N_9484,N_9040);
xor UO_719 (O_719,N_9751,N_8546);
and UO_720 (O_720,N_8556,N_9307);
nor UO_721 (O_721,N_9071,N_9324);
xnor UO_722 (O_722,N_8844,N_9649);
nor UO_723 (O_723,N_9480,N_8234);
or UO_724 (O_724,N_8757,N_8966);
xor UO_725 (O_725,N_9612,N_9076);
or UO_726 (O_726,N_9334,N_9826);
and UO_727 (O_727,N_9842,N_8840);
nand UO_728 (O_728,N_8571,N_8331);
or UO_729 (O_729,N_9934,N_8357);
nor UO_730 (O_730,N_9644,N_8943);
and UO_731 (O_731,N_9178,N_9591);
xor UO_732 (O_732,N_9327,N_8140);
nand UO_733 (O_733,N_8166,N_9357);
nor UO_734 (O_734,N_9917,N_9900);
nand UO_735 (O_735,N_8935,N_9107);
nand UO_736 (O_736,N_8124,N_9744);
and UO_737 (O_737,N_8282,N_9398);
xor UO_738 (O_738,N_9403,N_9017);
or UO_739 (O_739,N_8184,N_9229);
and UO_740 (O_740,N_9049,N_8500);
xnor UO_741 (O_741,N_8063,N_9295);
xnor UO_742 (O_742,N_8264,N_8772);
or UO_743 (O_743,N_9370,N_8213);
xnor UO_744 (O_744,N_8219,N_8464);
xor UO_745 (O_745,N_8863,N_9164);
xnor UO_746 (O_746,N_8940,N_8368);
xnor UO_747 (O_747,N_8999,N_8704);
or UO_748 (O_748,N_9205,N_8066);
and UO_749 (O_749,N_8091,N_9267);
nand UO_750 (O_750,N_9156,N_9522);
and UO_751 (O_751,N_8752,N_9073);
nand UO_752 (O_752,N_8400,N_8320);
xor UO_753 (O_753,N_8431,N_9888);
and UO_754 (O_754,N_8626,N_9870);
and UO_755 (O_755,N_8784,N_9696);
or UO_756 (O_756,N_9617,N_8550);
xnor UO_757 (O_757,N_8512,N_9727);
xnor UO_758 (O_758,N_9685,N_9388);
nor UO_759 (O_759,N_8114,N_9708);
nand UO_760 (O_760,N_8640,N_8061);
or UO_761 (O_761,N_8389,N_8130);
nor UO_762 (O_762,N_9359,N_9343);
or UO_763 (O_763,N_9463,N_8125);
xor UO_764 (O_764,N_8826,N_8905);
or UO_765 (O_765,N_8555,N_9597);
and UO_766 (O_766,N_8176,N_9112);
or UO_767 (O_767,N_8075,N_8674);
and UO_768 (O_768,N_9020,N_9077);
and UO_769 (O_769,N_9738,N_9220);
nor UO_770 (O_770,N_8726,N_9965);
nor UO_771 (O_771,N_9466,N_9442);
nand UO_772 (O_772,N_8214,N_9803);
nor UO_773 (O_773,N_9789,N_8127);
nor UO_774 (O_774,N_8315,N_9010);
nor UO_775 (O_775,N_9795,N_8458);
or UO_776 (O_776,N_8472,N_8513);
nand UO_777 (O_777,N_9780,N_8587);
xnor UO_778 (O_778,N_8543,N_8781);
xnor UO_779 (O_779,N_9896,N_9197);
and UO_780 (O_780,N_8447,N_8911);
or UO_781 (O_781,N_9193,N_9771);
nor UO_782 (O_782,N_9991,N_8137);
or UO_783 (O_783,N_9060,N_8466);
nand UO_784 (O_784,N_9006,N_8902);
and UO_785 (O_785,N_8698,N_8701);
xor UO_786 (O_786,N_8803,N_9846);
or UO_787 (O_787,N_8123,N_9238);
xnor UO_788 (O_788,N_8503,N_9811);
nand UO_789 (O_789,N_8873,N_8740);
nand UO_790 (O_790,N_8150,N_8813);
nand UO_791 (O_791,N_8259,N_8827);
nand UO_792 (O_792,N_8945,N_9761);
or UO_793 (O_793,N_8369,N_8049);
xnor UO_794 (O_794,N_8047,N_9973);
xor UO_795 (O_795,N_9251,N_8875);
nor UO_796 (O_796,N_8894,N_8919);
xnor UO_797 (O_797,N_9630,N_9366);
or UO_798 (O_798,N_9978,N_9314);
nand UO_799 (O_799,N_9200,N_9322);
or UO_800 (O_800,N_9245,N_9379);
xnor UO_801 (O_801,N_9691,N_8323);
nor UO_802 (O_802,N_9052,N_9226);
and UO_803 (O_803,N_9462,N_8258);
xnor UO_804 (O_804,N_9611,N_8168);
and UO_805 (O_805,N_9867,N_8853);
nor UO_806 (O_806,N_8295,N_9879);
xnor UO_807 (O_807,N_9131,N_8487);
xnor UO_808 (O_808,N_9864,N_8881);
or UO_809 (O_809,N_9624,N_9084);
and UO_810 (O_810,N_9782,N_8139);
nor UO_811 (O_811,N_8413,N_9004);
or UO_812 (O_812,N_9451,N_9899);
xor UO_813 (O_813,N_8980,N_8854);
nand UO_814 (O_814,N_8907,N_8134);
nor UO_815 (O_815,N_8265,N_8646);
xnor UO_816 (O_816,N_9603,N_8788);
nor UO_817 (O_817,N_8193,N_8363);
nor UO_818 (O_818,N_8561,N_8364);
nand UO_819 (O_819,N_9608,N_9445);
or UO_820 (O_820,N_8228,N_9812);
or UO_821 (O_821,N_8829,N_9805);
or UO_822 (O_822,N_9454,N_8644);
nor UO_823 (O_823,N_9533,N_9271);
nor UO_824 (O_824,N_8051,N_8498);
or UO_825 (O_825,N_8488,N_8658);
and UO_826 (O_826,N_8928,N_8567);
xnor UO_827 (O_827,N_8795,N_9575);
xnor UO_828 (O_828,N_9021,N_8274);
nor UO_829 (O_829,N_9749,N_8212);
xor UO_830 (O_830,N_8916,N_9099);
nor UO_831 (O_831,N_9668,N_9134);
and UO_832 (O_832,N_9317,N_8883);
xor UO_833 (O_833,N_8215,N_9215);
and UO_834 (O_834,N_8316,N_8304);
xor UO_835 (O_835,N_9702,N_9044);
and UO_836 (O_836,N_8708,N_9512);
and UO_837 (O_837,N_9967,N_9547);
xnor UO_838 (O_838,N_9120,N_8783);
or UO_839 (O_839,N_9458,N_8142);
nand UO_840 (O_840,N_8991,N_9260);
nor UO_841 (O_841,N_8549,N_9519);
and UO_842 (O_842,N_9654,N_9753);
nand UO_843 (O_843,N_9674,N_9110);
nor UO_844 (O_844,N_8670,N_8390);
xor UO_845 (O_845,N_8744,N_9063);
or UO_846 (O_846,N_9150,N_8187);
or UO_847 (O_847,N_9235,N_8762);
or UO_848 (O_848,N_9506,N_9453);
and UO_849 (O_849,N_8079,N_9619);
and UO_850 (O_850,N_8595,N_8805);
nand UO_851 (O_851,N_9832,N_8787);
and UO_852 (O_852,N_8330,N_9613);
or UO_853 (O_853,N_8206,N_8373);
nor UO_854 (O_854,N_8403,N_9486);
nand UO_855 (O_855,N_8420,N_9272);
nand UO_856 (O_856,N_9103,N_8120);
or UO_857 (O_857,N_9149,N_8468);
and UO_858 (O_858,N_9141,N_8663);
nand UO_859 (O_859,N_8773,N_8505);
and UO_860 (O_860,N_9629,N_8194);
or UO_861 (O_861,N_9648,N_8720);
xnor UO_862 (O_862,N_9495,N_9731);
and UO_863 (O_863,N_9535,N_9298);
xnor UO_864 (O_864,N_9488,N_8088);
nor UO_865 (O_865,N_8761,N_9450);
or UO_866 (O_866,N_9566,N_8475);
or UO_867 (O_867,N_9645,N_8042);
nand UO_868 (O_868,N_8542,N_8294);
and UO_869 (O_869,N_9572,N_9602);
or UO_870 (O_870,N_9997,N_9852);
or UO_871 (O_871,N_8737,N_9354);
nand UO_872 (O_872,N_9661,N_9723);
nand UO_873 (O_873,N_8662,N_9851);
xor UO_874 (O_874,N_9202,N_8719);
nand UO_875 (O_875,N_8284,N_9725);
and UO_876 (O_876,N_9054,N_9151);
nor UO_877 (O_877,N_8262,N_8240);
xor UO_878 (O_878,N_9984,N_8925);
or UO_879 (O_879,N_9296,N_8037);
xor UO_880 (O_880,N_8985,N_8248);
or UO_881 (O_881,N_9331,N_8714);
nand UO_882 (O_882,N_9072,N_8882);
nand UO_883 (O_883,N_9765,N_8451);
nor UO_884 (O_884,N_8006,N_9133);
nor UO_885 (O_885,N_8165,N_9000);
xor UO_886 (O_886,N_9136,N_8937);
or UO_887 (O_887,N_8151,N_9263);
xnor UO_888 (O_888,N_8697,N_8483);
and UO_889 (O_889,N_9743,N_8540);
nor UO_890 (O_890,N_8486,N_9443);
xor UO_891 (O_891,N_8839,N_9387);
and UO_892 (O_892,N_8607,N_8716);
nand UO_893 (O_893,N_8410,N_8923);
and UO_894 (O_894,N_9678,N_9528);
or UO_895 (O_895,N_8526,N_8080);
nor UO_896 (O_896,N_8113,N_9418);
nand UO_897 (O_897,N_8819,N_8365);
nand UO_898 (O_898,N_9787,N_9680);
and UO_899 (O_899,N_9037,N_8886);
xnor UO_900 (O_900,N_8791,N_9394);
and UO_901 (O_901,N_8578,N_8699);
nor UO_902 (O_902,N_9474,N_9036);
nor UO_903 (O_903,N_9344,N_9713);
nand UO_904 (O_904,N_8232,N_9923);
and UO_905 (O_905,N_9035,N_9587);
nor UO_906 (O_906,N_8967,N_8313);
xnor UO_907 (O_907,N_9189,N_9875);
nor UO_908 (O_908,N_8156,N_8177);
nand UO_909 (O_909,N_8837,N_9138);
xnor UO_910 (O_910,N_9449,N_8225);
and UO_911 (O_911,N_9257,N_8418);
and UO_912 (O_912,N_8939,N_9922);
nor UO_913 (O_913,N_8878,N_9790);
and UO_914 (O_914,N_9890,N_8696);
nand UO_915 (O_915,N_9906,N_9482);
nand UO_916 (O_916,N_9520,N_9995);
and UO_917 (O_917,N_8824,N_8777);
nand UO_918 (O_918,N_9175,N_8836);
nor UO_919 (O_919,N_9384,N_8145);
nand UO_920 (O_920,N_8862,N_9003);
or UO_921 (O_921,N_8544,N_9928);
nand UO_922 (O_922,N_9763,N_8077);
nand UO_923 (O_923,N_9204,N_8539);
xnor UO_924 (O_924,N_8917,N_8141);
and UO_925 (O_925,N_9554,N_9712);
nor UO_926 (O_926,N_9300,N_9882);
xnor UO_927 (O_927,N_9848,N_8437);
xor UO_928 (O_928,N_9289,N_9951);
and UO_929 (O_929,N_8407,N_9114);
and UO_930 (O_930,N_9700,N_9038);
nor UO_931 (O_931,N_9128,N_9048);
nand UO_932 (O_932,N_9970,N_8010);
nand UO_933 (O_933,N_8604,N_9868);
or UO_934 (O_934,N_8302,N_8034);
or UO_935 (O_935,N_9459,N_8804);
and UO_936 (O_936,N_8722,N_9721);
nand UO_937 (O_937,N_9421,N_9829);
or UO_938 (O_938,N_8469,N_8236);
xor UO_939 (O_939,N_8116,N_8876);
or UO_940 (O_940,N_8385,N_8594);
nor UO_941 (O_941,N_9853,N_9931);
and UO_942 (O_942,N_8770,N_9320);
nor UO_943 (O_943,N_9316,N_9153);
nand UO_944 (O_944,N_9350,N_8563);
nor UO_945 (O_945,N_8831,N_9807);
nor UO_946 (O_946,N_8071,N_8286);
nand UO_947 (O_947,N_9312,N_9652);
xnor UO_948 (O_948,N_9689,N_8728);
nor UO_949 (O_949,N_9093,N_8100);
and UO_950 (O_950,N_9735,N_8429);
nand UO_951 (O_951,N_9209,N_8598);
xor UO_952 (O_952,N_9971,N_9340);
and UO_953 (O_953,N_9146,N_9414);
nor UO_954 (O_954,N_8358,N_9511);
nor UO_955 (O_955,N_9026,N_9841);
nor UO_956 (O_956,N_9982,N_9464);
and UO_957 (O_957,N_8098,N_8277);
nor UO_958 (O_958,N_9426,N_9428);
or UO_959 (O_959,N_9901,N_8109);
and UO_960 (O_960,N_9911,N_9904);
xor UO_961 (O_961,N_8105,N_8551);
nand UO_962 (O_962,N_9082,N_9301);
xor UO_963 (O_963,N_9776,N_9955);
or UO_964 (O_964,N_8548,N_8059);
nand UO_965 (O_965,N_9325,N_9671);
nor UO_966 (O_966,N_9526,N_9540);
or UO_967 (O_967,N_8970,N_8336);
nand UO_968 (O_968,N_8337,N_8055);
nand UO_969 (O_969,N_9274,N_9657);
nor UO_970 (O_970,N_9703,N_9304);
nand UO_971 (O_971,N_9493,N_9855);
or UO_972 (O_972,N_8617,N_8297);
nor UO_973 (O_973,N_9518,N_8268);
or UO_974 (O_974,N_9397,N_8060);
nand UO_975 (O_975,N_8903,N_9233);
nor UO_976 (O_976,N_9009,N_8235);
xor UO_977 (O_977,N_8338,N_8832);
nand UO_978 (O_978,N_8243,N_8424);
nand UO_979 (O_979,N_8462,N_8426);
xor UO_980 (O_980,N_8810,N_9192);
nor UO_981 (O_981,N_9569,N_9218);
nor UO_982 (O_982,N_9031,N_9306);
xnor UO_983 (O_983,N_9053,N_9191);
xnor UO_984 (O_984,N_9954,N_9690);
nand UO_985 (O_985,N_8982,N_9975);
xor UO_986 (O_986,N_8306,N_9034);
nand UO_987 (O_987,N_9541,N_9546);
or UO_988 (O_988,N_8857,N_9714);
xor UO_989 (O_989,N_8372,N_9673);
or UO_990 (O_990,N_8828,N_8270);
and UO_991 (O_991,N_8054,N_8659);
xor UO_992 (O_992,N_9983,N_8053);
nand UO_993 (O_993,N_8344,N_9019);
nand UO_994 (O_994,N_8929,N_9642);
or UO_995 (O_995,N_8866,N_8200);
nor UO_996 (O_996,N_8729,N_9195);
nand UO_997 (O_997,N_9064,N_8618);
or UO_998 (O_998,N_9363,N_9117);
and UO_999 (O_999,N_9069,N_8019);
xnor UO_1000 (O_1000,N_8037,N_9953);
and UO_1001 (O_1001,N_8379,N_8754);
xor UO_1002 (O_1002,N_8193,N_8058);
and UO_1003 (O_1003,N_9176,N_9578);
or UO_1004 (O_1004,N_9777,N_9547);
nor UO_1005 (O_1005,N_8009,N_9299);
nor UO_1006 (O_1006,N_9677,N_8824);
or UO_1007 (O_1007,N_9456,N_9637);
xnor UO_1008 (O_1008,N_8341,N_8925);
nand UO_1009 (O_1009,N_8963,N_9491);
nand UO_1010 (O_1010,N_9190,N_9343);
nor UO_1011 (O_1011,N_9894,N_8569);
xnor UO_1012 (O_1012,N_9095,N_8109);
or UO_1013 (O_1013,N_9918,N_9975);
or UO_1014 (O_1014,N_8967,N_8953);
xnor UO_1015 (O_1015,N_8175,N_8347);
nor UO_1016 (O_1016,N_8602,N_8112);
nand UO_1017 (O_1017,N_9064,N_9897);
nand UO_1018 (O_1018,N_9940,N_8545);
nand UO_1019 (O_1019,N_8352,N_9459);
nor UO_1020 (O_1020,N_8683,N_9852);
nand UO_1021 (O_1021,N_8555,N_8022);
nor UO_1022 (O_1022,N_9686,N_9180);
xnor UO_1023 (O_1023,N_9139,N_9310);
xor UO_1024 (O_1024,N_8872,N_8924);
xor UO_1025 (O_1025,N_9922,N_9109);
xor UO_1026 (O_1026,N_9373,N_8181);
xnor UO_1027 (O_1027,N_8803,N_8366);
nor UO_1028 (O_1028,N_8706,N_9749);
xnor UO_1029 (O_1029,N_9445,N_8763);
and UO_1030 (O_1030,N_8711,N_8556);
and UO_1031 (O_1031,N_8870,N_9320);
and UO_1032 (O_1032,N_9142,N_9386);
nor UO_1033 (O_1033,N_8385,N_9653);
and UO_1034 (O_1034,N_8686,N_9086);
nor UO_1035 (O_1035,N_8846,N_8949);
nor UO_1036 (O_1036,N_8289,N_9585);
nor UO_1037 (O_1037,N_9248,N_9110);
or UO_1038 (O_1038,N_8921,N_9233);
nor UO_1039 (O_1039,N_9058,N_8422);
and UO_1040 (O_1040,N_9264,N_8464);
and UO_1041 (O_1041,N_8448,N_8168);
nand UO_1042 (O_1042,N_8580,N_8408);
and UO_1043 (O_1043,N_8900,N_8606);
nand UO_1044 (O_1044,N_8753,N_9678);
nor UO_1045 (O_1045,N_8956,N_8194);
and UO_1046 (O_1046,N_9496,N_8069);
or UO_1047 (O_1047,N_9544,N_8230);
nor UO_1048 (O_1048,N_8288,N_9676);
nand UO_1049 (O_1049,N_9897,N_8732);
or UO_1050 (O_1050,N_9174,N_9741);
or UO_1051 (O_1051,N_8070,N_9376);
nand UO_1052 (O_1052,N_8609,N_8996);
nand UO_1053 (O_1053,N_8769,N_8886);
nand UO_1054 (O_1054,N_9677,N_9271);
or UO_1055 (O_1055,N_8664,N_9394);
nand UO_1056 (O_1056,N_8907,N_9209);
nor UO_1057 (O_1057,N_9623,N_9551);
or UO_1058 (O_1058,N_8513,N_8448);
or UO_1059 (O_1059,N_8144,N_8085);
nor UO_1060 (O_1060,N_9124,N_8073);
or UO_1061 (O_1061,N_8440,N_9642);
or UO_1062 (O_1062,N_9289,N_8496);
or UO_1063 (O_1063,N_9669,N_9346);
and UO_1064 (O_1064,N_9569,N_9784);
and UO_1065 (O_1065,N_8291,N_9272);
or UO_1066 (O_1066,N_9278,N_8817);
or UO_1067 (O_1067,N_8152,N_9515);
and UO_1068 (O_1068,N_9400,N_8293);
nand UO_1069 (O_1069,N_8119,N_9643);
xor UO_1070 (O_1070,N_8600,N_9851);
nand UO_1071 (O_1071,N_9769,N_8288);
xnor UO_1072 (O_1072,N_8996,N_8041);
nand UO_1073 (O_1073,N_8127,N_9421);
nor UO_1074 (O_1074,N_8522,N_9021);
nor UO_1075 (O_1075,N_8346,N_8015);
nor UO_1076 (O_1076,N_8290,N_8489);
or UO_1077 (O_1077,N_8187,N_8186);
xor UO_1078 (O_1078,N_9718,N_9328);
nor UO_1079 (O_1079,N_9206,N_8072);
nand UO_1080 (O_1080,N_9923,N_9848);
nor UO_1081 (O_1081,N_9886,N_9842);
xnor UO_1082 (O_1082,N_9148,N_9342);
or UO_1083 (O_1083,N_9826,N_9930);
and UO_1084 (O_1084,N_9288,N_8360);
nand UO_1085 (O_1085,N_9627,N_9008);
and UO_1086 (O_1086,N_8307,N_9033);
nor UO_1087 (O_1087,N_9712,N_8243);
or UO_1088 (O_1088,N_9318,N_9501);
and UO_1089 (O_1089,N_8298,N_9711);
or UO_1090 (O_1090,N_8433,N_9687);
or UO_1091 (O_1091,N_9512,N_9062);
and UO_1092 (O_1092,N_8511,N_8302);
and UO_1093 (O_1093,N_9695,N_8719);
or UO_1094 (O_1094,N_8869,N_9418);
or UO_1095 (O_1095,N_8117,N_9982);
xor UO_1096 (O_1096,N_8316,N_9716);
nor UO_1097 (O_1097,N_9286,N_9789);
or UO_1098 (O_1098,N_9281,N_8965);
or UO_1099 (O_1099,N_8983,N_9984);
or UO_1100 (O_1100,N_9775,N_8443);
nor UO_1101 (O_1101,N_9290,N_9091);
or UO_1102 (O_1102,N_8662,N_9650);
or UO_1103 (O_1103,N_9611,N_9502);
xor UO_1104 (O_1104,N_8982,N_8578);
xor UO_1105 (O_1105,N_9639,N_8885);
or UO_1106 (O_1106,N_8193,N_9047);
and UO_1107 (O_1107,N_9081,N_9441);
nor UO_1108 (O_1108,N_9774,N_9658);
xnor UO_1109 (O_1109,N_9097,N_8964);
or UO_1110 (O_1110,N_9789,N_8500);
nand UO_1111 (O_1111,N_9753,N_8013);
xnor UO_1112 (O_1112,N_9636,N_9216);
nor UO_1113 (O_1113,N_8048,N_9266);
nor UO_1114 (O_1114,N_8518,N_8363);
nand UO_1115 (O_1115,N_9552,N_9333);
xor UO_1116 (O_1116,N_9840,N_9480);
nand UO_1117 (O_1117,N_9835,N_8514);
nand UO_1118 (O_1118,N_9293,N_9211);
or UO_1119 (O_1119,N_8563,N_8721);
or UO_1120 (O_1120,N_8322,N_9903);
xor UO_1121 (O_1121,N_8761,N_8828);
or UO_1122 (O_1122,N_9860,N_8890);
and UO_1123 (O_1123,N_8228,N_9801);
and UO_1124 (O_1124,N_8220,N_9460);
nand UO_1125 (O_1125,N_8613,N_9215);
or UO_1126 (O_1126,N_9214,N_8312);
nand UO_1127 (O_1127,N_8532,N_9855);
or UO_1128 (O_1128,N_8500,N_8822);
nor UO_1129 (O_1129,N_9678,N_9717);
or UO_1130 (O_1130,N_9116,N_8420);
xnor UO_1131 (O_1131,N_8892,N_8632);
nand UO_1132 (O_1132,N_8557,N_9300);
or UO_1133 (O_1133,N_8200,N_8519);
or UO_1134 (O_1134,N_9652,N_8883);
xor UO_1135 (O_1135,N_8857,N_9017);
nor UO_1136 (O_1136,N_9834,N_8629);
or UO_1137 (O_1137,N_8838,N_8494);
nor UO_1138 (O_1138,N_9082,N_9246);
xor UO_1139 (O_1139,N_8298,N_8367);
or UO_1140 (O_1140,N_9477,N_8014);
nor UO_1141 (O_1141,N_9117,N_9814);
nor UO_1142 (O_1142,N_8936,N_9030);
nand UO_1143 (O_1143,N_8241,N_9088);
nor UO_1144 (O_1144,N_8688,N_8609);
or UO_1145 (O_1145,N_8685,N_9322);
xnor UO_1146 (O_1146,N_9056,N_9894);
nand UO_1147 (O_1147,N_8409,N_8020);
xor UO_1148 (O_1148,N_8936,N_9497);
and UO_1149 (O_1149,N_8903,N_8379);
or UO_1150 (O_1150,N_8896,N_8564);
nor UO_1151 (O_1151,N_9233,N_8165);
or UO_1152 (O_1152,N_8031,N_8544);
or UO_1153 (O_1153,N_8613,N_9421);
nand UO_1154 (O_1154,N_8913,N_9086);
nor UO_1155 (O_1155,N_9456,N_9124);
nand UO_1156 (O_1156,N_9446,N_8520);
and UO_1157 (O_1157,N_8986,N_8602);
and UO_1158 (O_1158,N_9471,N_9863);
and UO_1159 (O_1159,N_9656,N_8621);
or UO_1160 (O_1160,N_8158,N_8915);
or UO_1161 (O_1161,N_8784,N_9013);
or UO_1162 (O_1162,N_9057,N_9625);
xor UO_1163 (O_1163,N_9812,N_8679);
or UO_1164 (O_1164,N_9935,N_8831);
nor UO_1165 (O_1165,N_9581,N_9470);
xor UO_1166 (O_1166,N_9130,N_9562);
nand UO_1167 (O_1167,N_8379,N_8869);
nor UO_1168 (O_1168,N_8248,N_9136);
nand UO_1169 (O_1169,N_8964,N_8053);
xor UO_1170 (O_1170,N_9298,N_8661);
nor UO_1171 (O_1171,N_9969,N_8335);
xnor UO_1172 (O_1172,N_9119,N_9763);
nor UO_1173 (O_1173,N_8514,N_8375);
xor UO_1174 (O_1174,N_8624,N_9926);
or UO_1175 (O_1175,N_9664,N_9597);
or UO_1176 (O_1176,N_8469,N_9373);
and UO_1177 (O_1177,N_8218,N_8599);
nand UO_1178 (O_1178,N_9377,N_8812);
xnor UO_1179 (O_1179,N_9123,N_9593);
or UO_1180 (O_1180,N_8597,N_8625);
nor UO_1181 (O_1181,N_8114,N_9092);
nor UO_1182 (O_1182,N_8274,N_8229);
nor UO_1183 (O_1183,N_8054,N_9115);
xnor UO_1184 (O_1184,N_8466,N_9099);
and UO_1185 (O_1185,N_9828,N_9061);
xnor UO_1186 (O_1186,N_9428,N_8636);
or UO_1187 (O_1187,N_8487,N_9736);
or UO_1188 (O_1188,N_8234,N_9259);
nor UO_1189 (O_1189,N_9127,N_9895);
nor UO_1190 (O_1190,N_9995,N_8764);
and UO_1191 (O_1191,N_8016,N_8981);
nand UO_1192 (O_1192,N_8990,N_8248);
xor UO_1193 (O_1193,N_8101,N_8390);
or UO_1194 (O_1194,N_8586,N_9291);
xor UO_1195 (O_1195,N_9677,N_8498);
nor UO_1196 (O_1196,N_8066,N_8296);
nand UO_1197 (O_1197,N_8175,N_9159);
nand UO_1198 (O_1198,N_9779,N_8031);
nor UO_1199 (O_1199,N_8136,N_9728);
and UO_1200 (O_1200,N_8143,N_9925);
and UO_1201 (O_1201,N_9922,N_9145);
nor UO_1202 (O_1202,N_9351,N_8564);
xor UO_1203 (O_1203,N_9604,N_8629);
or UO_1204 (O_1204,N_9839,N_9362);
xor UO_1205 (O_1205,N_9721,N_8400);
nor UO_1206 (O_1206,N_8754,N_8356);
nor UO_1207 (O_1207,N_8397,N_8978);
xor UO_1208 (O_1208,N_8674,N_8900);
or UO_1209 (O_1209,N_9313,N_8750);
xnor UO_1210 (O_1210,N_8676,N_9314);
nor UO_1211 (O_1211,N_8817,N_9475);
nor UO_1212 (O_1212,N_8877,N_9549);
nand UO_1213 (O_1213,N_9986,N_8800);
xnor UO_1214 (O_1214,N_8923,N_8168);
xor UO_1215 (O_1215,N_8915,N_9855);
or UO_1216 (O_1216,N_9193,N_9311);
nand UO_1217 (O_1217,N_9788,N_9785);
nor UO_1218 (O_1218,N_9402,N_9533);
nor UO_1219 (O_1219,N_8712,N_9068);
or UO_1220 (O_1220,N_9429,N_9059);
and UO_1221 (O_1221,N_9903,N_8542);
nand UO_1222 (O_1222,N_8643,N_8614);
and UO_1223 (O_1223,N_9639,N_9905);
xor UO_1224 (O_1224,N_8745,N_9545);
nand UO_1225 (O_1225,N_8855,N_8091);
nor UO_1226 (O_1226,N_9991,N_8283);
and UO_1227 (O_1227,N_9081,N_8181);
and UO_1228 (O_1228,N_8904,N_9349);
nand UO_1229 (O_1229,N_9794,N_8759);
and UO_1230 (O_1230,N_8249,N_8960);
nor UO_1231 (O_1231,N_9895,N_9493);
and UO_1232 (O_1232,N_9098,N_8931);
nand UO_1233 (O_1233,N_8516,N_9679);
nor UO_1234 (O_1234,N_8242,N_9704);
nand UO_1235 (O_1235,N_9288,N_9987);
and UO_1236 (O_1236,N_8553,N_8589);
nor UO_1237 (O_1237,N_8639,N_9405);
and UO_1238 (O_1238,N_8029,N_9322);
or UO_1239 (O_1239,N_8586,N_9640);
or UO_1240 (O_1240,N_8615,N_8593);
xnor UO_1241 (O_1241,N_9408,N_8427);
and UO_1242 (O_1242,N_8951,N_8949);
xor UO_1243 (O_1243,N_8115,N_9738);
or UO_1244 (O_1244,N_9569,N_9157);
and UO_1245 (O_1245,N_8634,N_9050);
and UO_1246 (O_1246,N_8806,N_8668);
or UO_1247 (O_1247,N_8365,N_8392);
or UO_1248 (O_1248,N_9521,N_9258);
nand UO_1249 (O_1249,N_9924,N_9875);
nor UO_1250 (O_1250,N_8545,N_9458);
xnor UO_1251 (O_1251,N_8519,N_9304);
nand UO_1252 (O_1252,N_9123,N_9087);
or UO_1253 (O_1253,N_9224,N_9953);
nor UO_1254 (O_1254,N_9967,N_9553);
nand UO_1255 (O_1255,N_8115,N_8994);
nand UO_1256 (O_1256,N_8808,N_8051);
nor UO_1257 (O_1257,N_8465,N_9047);
nand UO_1258 (O_1258,N_8211,N_9146);
nand UO_1259 (O_1259,N_9742,N_8391);
nor UO_1260 (O_1260,N_9292,N_8473);
xnor UO_1261 (O_1261,N_8141,N_8542);
and UO_1262 (O_1262,N_9654,N_8544);
nand UO_1263 (O_1263,N_8671,N_9580);
or UO_1264 (O_1264,N_9400,N_9233);
or UO_1265 (O_1265,N_9664,N_9697);
and UO_1266 (O_1266,N_8870,N_8701);
xor UO_1267 (O_1267,N_8237,N_8980);
nand UO_1268 (O_1268,N_8272,N_8790);
nand UO_1269 (O_1269,N_8724,N_9891);
xnor UO_1270 (O_1270,N_9655,N_8511);
or UO_1271 (O_1271,N_9580,N_9108);
nand UO_1272 (O_1272,N_8651,N_9898);
and UO_1273 (O_1273,N_8706,N_9822);
and UO_1274 (O_1274,N_9051,N_9883);
nor UO_1275 (O_1275,N_8919,N_9997);
or UO_1276 (O_1276,N_9381,N_8386);
xnor UO_1277 (O_1277,N_8317,N_9610);
nand UO_1278 (O_1278,N_8971,N_8102);
nand UO_1279 (O_1279,N_8086,N_9011);
and UO_1280 (O_1280,N_9173,N_8844);
or UO_1281 (O_1281,N_9118,N_9162);
xor UO_1282 (O_1282,N_8856,N_9492);
xnor UO_1283 (O_1283,N_8494,N_9623);
nand UO_1284 (O_1284,N_9387,N_9537);
and UO_1285 (O_1285,N_8007,N_9067);
and UO_1286 (O_1286,N_8488,N_9179);
and UO_1287 (O_1287,N_9085,N_8720);
nor UO_1288 (O_1288,N_8827,N_8265);
xor UO_1289 (O_1289,N_9533,N_8975);
or UO_1290 (O_1290,N_8100,N_9829);
or UO_1291 (O_1291,N_8526,N_9294);
nand UO_1292 (O_1292,N_9127,N_8239);
xor UO_1293 (O_1293,N_8357,N_8111);
and UO_1294 (O_1294,N_8845,N_9023);
nor UO_1295 (O_1295,N_8866,N_9743);
or UO_1296 (O_1296,N_8918,N_9664);
or UO_1297 (O_1297,N_9162,N_8249);
and UO_1298 (O_1298,N_9159,N_8413);
and UO_1299 (O_1299,N_8276,N_9716);
and UO_1300 (O_1300,N_9421,N_8372);
and UO_1301 (O_1301,N_8670,N_8402);
and UO_1302 (O_1302,N_9371,N_9104);
or UO_1303 (O_1303,N_8416,N_8463);
or UO_1304 (O_1304,N_9766,N_9620);
or UO_1305 (O_1305,N_8550,N_8907);
nor UO_1306 (O_1306,N_9058,N_9890);
xnor UO_1307 (O_1307,N_9736,N_8867);
nor UO_1308 (O_1308,N_9079,N_8960);
nand UO_1309 (O_1309,N_9536,N_9894);
and UO_1310 (O_1310,N_9716,N_8535);
xnor UO_1311 (O_1311,N_8134,N_8498);
nor UO_1312 (O_1312,N_8316,N_8216);
and UO_1313 (O_1313,N_8529,N_9936);
nand UO_1314 (O_1314,N_9763,N_9449);
nand UO_1315 (O_1315,N_8174,N_8288);
nor UO_1316 (O_1316,N_9312,N_8880);
nor UO_1317 (O_1317,N_8141,N_8964);
or UO_1318 (O_1318,N_8891,N_9875);
nand UO_1319 (O_1319,N_9100,N_9089);
xnor UO_1320 (O_1320,N_8444,N_8343);
nand UO_1321 (O_1321,N_8311,N_9041);
xor UO_1322 (O_1322,N_8273,N_8201);
xor UO_1323 (O_1323,N_9055,N_9206);
xnor UO_1324 (O_1324,N_8895,N_9514);
and UO_1325 (O_1325,N_8187,N_8872);
and UO_1326 (O_1326,N_9967,N_9120);
nor UO_1327 (O_1327,N_8502,N_8504);
nor UO_1328 (O_1328,N_8048,N_8218);
and UO_1329 (O_1329,N_8810,N_9212);
nand UO_1330 (O_1330,N_8478,N_9995);
or UO_1331 (O_1331,N_8005,N_9549);
and UO_1332 (O_1332,N_9223,N_8398);
nor UO_1333 (O_1333,N_9767,N_8048);
nand UO_1334 (O_1334,N_8362,N_9546);
nor UO_1335 (O_1335,N_8242,N_8213);
and UO_1336 (O_1336,N_8569,N_8761);
and UO_1337 (O_1337,N_8492,N_9428);
nand UO_1338 (O_1338,N_8657,N_9688);
or UO_1339 (O_1339,N_8087,N_8584);
or UO_1340 (O_1340,N_8001,N_8572);
nand UO_1341 (O_1341,N_8574,N_9769);
nor UO_1342 (O_1342,N_8059,N_8882);
or UO_1343 (O_1343,N_8140,N_9445);
xnor UO_1344 (O_1344,N_8064,N_9685);
and UO_1345 (O_1345,N_8711,N_8438);
or UO_1346 (O_1346,N_8758,N_9481);
and UO_1347 (O_1347,N_9898,N_9151);
and UO_1348 (O_1348,N_9378,N_8594);
and UO_1349 (O_1349,N_8592,N_9895);
and UO_1350 (O_1350,N_9978,N_9876);
xnor UO_1351 (O_1351,N_8935,N_9947);
nor UO_1352 (O_1352,N_9488,N_9159);
xnor UO_1353 (O_1353,N_9380,N_8338);
nand UO_1354 (O_1354,N_9688,N_8387);
xor UO_1355 (O_1355,N_9800,N_8107);
nand UO_1356 (O_1356,N_9623,N_8316);
or UO_1357 (O_1357,N_9773,N_8285);
nand UO_1358 (O_1358,N_9967,N_9652);
xor UO_1359 (O_1359,N_8694,N_8035);
or UO_1360 (O_1360,N_8439,N_9882);
xnor UO_1361 (O_1361,N_9409,N_8548);
or UO_1362 (O_1362,N_8801,N_9874);
nor UO_1363 (O_1363,N_8570,N_9328);
and UO_1364 (O_1364,N_8997,N_9998);
and UO_1365 (O_1365,N_9286,N_9921);
and UO_1366 (O_1366,N_8546,N_8344);
nor UO_1367 (O_1367,N_8913,N_8587);
or UO_1368 (O_1368,N_9828,N_9187);
and UO_1369 (O_1369,N_8413,N_9246);
or UO_1370 (O_1370,N_9730,N_8373);
and UO_1371 (O_1371,N_8037,N_9220);
xor UO_1372 (O_1372,N_9200,N_8682);
nand UO_1373 (O_1373,N_9939,N_9696);
nor UO_1374 (O_1374,N_9866,N_8355);
or UO_1375 (O_1375,N_8543,N_9167);
nand UO_1376 (O_1376,N_8403,N_8447);
xor UO_1377 (O_1377,N_8300,N_9326);
or UO_1378 (O_1378,N_8964,N_8895);
nor UO_1379 (O_1379,N_8806,N_9607);
xnor UO_1380 (O_1380,N_8668,N_9370);
or UO_1381 (O_1381,N_9255,N_9132);
and UO_1382 (O_1382,N_8822,N_8606);
nand UO_1383 (O_1383,N_8052,N_9089);
xor UO_1384 (O_1384,N_8029,N_9142);
or UO_1385 (O_1385,N_8117,N_8111);
nand UO_1386 (O_1386,N_9159,N_8434);
and UO_1387 (O_1387,N_8810,N_9452);
nand UO_1388 (O_1388,N_8487,N_8572);
and UO_1389 (O_1389,N_8208,N_9590);
nor UO_1390 (O_1390,N_8966,N_8537);
xnor UO_1391 (O_1391,N_8901,N_9432);
or UO_1392 (O_1392,N_9813,N_8929);
or UO_1393 (O_1393,N_9905,N_9845);
nand UO_1394 (O_1394,N_8468,N_9489);
nand UO_1395 (O_1395,N_9703,N_9495);
or UO_1396 (O_1396,N_8924,N_8488);
nand UO_1397 (O_1397,N_8769,N_9057);
or UO_1398 (O_1398,N_8431,N_8403);
and UO_1399 (O_1399,N_8199,N_8554);
nand UO_1400 (O_1400,N_8865,N_8394);
nor UO_1401 (O_1401,N_8855,N_8438);
nand UO_1402 (O_1402,N_9416,N_8977);
nand UO_1403 (O_1403,N_8448,N_8323);
nand UO_1404 (O_1404,N_8819,N_9413);
or UO_1405 (O_1405,N_9622,N_9588);
or UO_1406 (O_1406,N_8503,N_9876);
and UO_1407 (O_1407,N_9486,N_8505);
nand UO_1408 (O_1408,N_9252,N_9708);
nor UO_1409 (O_1409,N_9853,N_9438);
nor UO_1410 (O_1410,N_8741,N_9021);
and UO_1411 (O_1411,N_9516,N_9078);
and UO_1412 (O_1412,N_8560,N_8396);
nand UO_1413 (O_1413,N_8852,N_9580);
xor UO_1414 (O_1414,N_9191,N_8040);
xor UO_1415 (O_1415,N_8371,N_9269);
nand UO_1416 (O_1416,N_9809,N_9285);
xor UO_1417 (O_1417,N_9511,N_8392);
and UO_1418 (O_1418,N_8805,N_8648);
nor UO_1419 (O_1419,N_8978,N_9508);
and UO_1420 (O_1420,N_8257,N_8137);
nand UO_1421 (O_1421,N_8756,N_8880);
and UO_1422 (O_1422,N_9733,N_8810);
xnor UO_1423 (O_1423,N_8303,N_9292);
nor UO_1424 (O_1424,N_8726,N_9481);
nor UO_1425 (O_1425,N_9517,N_8952);
and UO_1426 (O_1426,N_9743,N_8899);
nor UO_1427 (O_1427,N_9564,N_8292);
and UO_1428 (O_1428,N_9248,N_8842);
nor UO_1429 (O_1429,N_9380,N_8259);
or UO_1430 (O_1430,N_8938,N_9117);
and UO_1431 (O_1431,N_9540,N_9331);
or UO_1432 (O_1432,N_9099,N_9370);
nor UO_1433 (O_1433,N_8382,N_9223);
nand UO_1434 (O_1434,N_9237,N_9002);
and UO_1435 (O_1435,N_8870,N_9936);
nand UO_1436 (O_1436,N_8661,N_8095);
nand UO_1437 (O_1437,N_9790,N_9471);
nand UO_1438 (O_1438,N_9299,N_9836);
nand UO_1439 (O_1439,N_8160,N_9089);
or UO_1440 (O_1440,N_9810,N_8017);
nor UO_1441 (O_1441,N_8688,N_9184);
xor UO_1442 (O_1442,N_9989,N_8662);
nand UO_1443 (O_1443,N_8473,N_8349);
or UO_1444 (O_1444,N_8630,N_8291);
nand UO_1445 (O_1445,N_8340,N_9963);
nor UO_1446 (O_1446,N_9564,N_9579);
nor UO_1447 (O_1447,N_9625,N_9120);
or UO_1448 (O_1448,N_8956,N_8516);
xor UO_1449 (O_1449,N_8325,N_8006);
nor UO_1450 (O_1450,N_9339,N_9445);
or UO_1451 (O_1451,N_9894,N_8644);
nand UO_1452 (O_1452,N_8543,N_8029);
nor UO_1453 (O_1453,N_8038,N_8661);
and UO_1454 (O_1454,N_9262,N_9646);
nor UO_1455 (O_1455,N_8032,N_9322);
nor UO_1456 (O_1456,N_8913,N_9470);
xor UO_1457 (O_1457,N_9544,N_8069);
nand UO_1458 (O_1458,N_8574,N_9734);
nor UO_1459 (O_1459,N_8199,N_9558);
xnor UO_1460 (O_1460,N_9495,N_9554);
xor UO_1461 (O_1461,N_8168,N_9374);
and UO_1462 (O_1462,N_8710,N_9948);
nand UO_1463 (O_1463,N_9929,N_9589);
xor UO_1464 (O_1464,N_8667,N_9707);
nand UO_1465 (O_1465,N_8884,N_9665);
nand UO_1466 (O_1466,N_8922,N_8819);
and UO_1467 (O_1467,N_8819,N_9707);
or UO_1468 (O_1468,N_8629,N_8464);
nor UO_1469 (O_1469,N_9261,N_9117);
and UO_1470 (O_1470,N_9194,N_8541);
nor UO_1471 (O_1471,N_8071,N_9326);
nor UO_1472 (O_1472,N_9237,N_9955);
xnor UO_1473 (O_1473,N_8766,N_9584);
nand UO_1474 (O_1474,N_9334,N_8015);
nand UO_1475 (O_1475,N_8260,N_8585);
nand UO_1476 (O_1476,N_8163,N_8495);
or UO_1477 (O_1477,N_8161,N_9446);
nor UO_1478 (O_1478,N_9928,N_9424);
nor UO_1479 (O_1479,N_9145,N_9380);
xnor UO_1480 (O_1480,N_9807,N_8706);
xor UO_1481 (O_1481,N_8392,N_8322);
or UO_1482 (O_1482,N_9284,N_9877);
nand UO_1483 (O_1483,N_9523,N_8638);
nand UO_1484 (O_1484,N_9347,N_8570);
nand UO_1485 (O_1485,N_8493,N_8549);
and UO_1486 (O_1486,N_8759,N_8743);
and UO_1487 (O_1487,N_8890,N_8721);
and UO_1488 (O_1488,N_9557,N_8723);
xor UO_1489 (O_1489,N_9592,N_9933);
and UO_1490 (O_1490,N_8166,N_9579);
or UO_1491 (O_1491,N_9797,N_8709);
nand UO_1492 (O_1492,N_8179,N_9199);
xnor UO_1493 (O_1493,N_9199,N_8395);
or UO_1494 (O_1494,N_8520,N_8625);
and UO_1495 (O_1495,N_9515,N_8623);
xnor UO_1496 (O_1496,N_9591,N_9561);
or UO_1497 (O_1497,N_9989,N_9492);
xnor UO_1498 (O_1498,N_8872,N_9729);
nand UO_1499 (O_1499,N_9840,N_8801);
endmodule