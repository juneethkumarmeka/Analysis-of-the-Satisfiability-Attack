module basic_750_5000_1000_10_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_630,In_726);
and U1 (N_1,In_360,In_730);
nor U2 (N_2,In_50,In_7);
xor U3 (N_3,In_435,In_97);
or U4 (N_4,In_65,In_633);
or U5 (N_5,In_235,In_711);
nor U6 (N_6,In_44,In_584);
or U7 (N_7,In_628,In_308);
nor U8 (N_8,In_452,In_25);
nor U9 (N_9,In_673,In_226);
and U10 (N_10,In_196,In_697);
xnor U11 (N_11,In_8,In_282);
or U12 (N_12,In_285,In_731);
xnor U13 (N_13,In_120,In_131);
xnor U14 (N_14,In_586,In_642);
nor U15 (N_15,In_350,In_221);
nor U16 (N_16,In_68,In_651);
xor U17 (N_17,In_481,In_346);
nand U18 (N_18,In_114,In_229);
nor U19 (N_19,In_557,In_333);
and U20 (N_20,In_189,In_667);
and U21 (N_21,In_301,In_109);
nor U22 (N_22,In_616,In_27);
xnor U23 (N_23,In_553,In_577);
or U24 (N_24,In_603,In_555);
or U25 (N_25,In_256,In_193);
nor U26 (N_26,In_631,In_179);
nor U27 (N_27,In_485,In_211);
nor U28 (N_28,In_100,In_85);
xnor U29 (N_29,In_475,In_99);
xor U30 (N_30,In_454,In_447);
nor U31 (N_31,In_140,In_80);
nor U32 (N_32,In_626,In_228);
or U33 (N_33,In_347,In_232);
and U34 (N_34,In_477,In_71);
nand U35 (N_35,In_184,In_579);
nand U36 (N_36,In_537,In_268);
and U37 (N_37,In_366,In_620);
nor U38 (N_38,In_29,In_458);
xnor U39 (N_39,In_23,In_104);
nand U40 (N_40,In_204,In_135);
or U41 (N_41,In_713,In_265);
nor U42 (N_42,In_385,In_195);
xnor U43 (N_43,In_541,In_147);
and U44 (N_44,In_206,In_736);
xor U45 (N_45,In_469,In_244);
or U46 (N_46,In_66,In_247);
nand U47 (N_47,In_723,In_688);
and U48 (N_48,In_267,In_470);
nor U49 (N_49,In_431,In_327);
and U50 (N_50,In_30,In_672);
and U51 (N_51,In_441,In_559);
nand U52 (N_52,In_406,In_134);
xnor U53 (N_53,In_41,In_510);
xnor U54 (N_54,In_362,In_298);
nand U55 (N_55,In_400,In_177);
xnor U56 (N_56,In_554,In_627);
or U57 (N_57,In_446,In_155);
nor U58 (N_58,In_574,In_450);
and U59 (N_59,In_462,In_205);
xnor U60 (N_60,In_277,In_397);
nor U61 (N_61,In_416,In_329);
xnor U62 (N_62,In_173,In_345);
or U63 (N_63,In_367,In_434);
or U64 (N_64,In_534,In_300);
nand U65 (N_65,In_497,In_84);
and U66 (N_66,In_118,In_359);
or U67 (N_67,In_549,In_523);
nor U68 (N_68,In_461,In_5);
or U69 (N_69,In_575,In_153);
and U70 (N_70,In_210,In_371);
nand U71 (N_71,In_336,In_662);
and U72 (N_72,In_172,In_354);
xor U73 (N_73,In_75,In_207);
xor U74 (N_74,In_401,In_543);
or U75 (N_75,In_91,In_528);
xnor U76 (N_76,In_437,In_525);
xor U77 (N_77,In_505,In_121);
and U78 (N_78,In_746,In_637);
nand U79 (N_79,In_619,In_491);
nor U80 (N_80,In_563,In_604);
xnor U81 (N_81,In_643,In_103);
and U82 (N_82,In_495,In_597);
xor U83 (N_83,In_31,In_258);
nand U84 (N_84,In_58,In_339);
nor U85 (N_85,In_424,In_724);
nand U86 (N_86,In_14,In_666);
nand U87 (N_87,In_227,In_415);
and U88 (N_88,In_79,In_641);
xnor U89 (N_89,In_324,In_378);
or U90 (N_90,In_117,In_388);
nor U91 (N_91,In_356,In_209);
or U92 (N_92,In_669,In_102);
or U93 (N_93,In_421,In_363);
xor U94 (N_94,In_544,In_343);
or U95 (N_95,In_457,In_741);
or U96 (N_96,In_476,In_634);
xor U97 (N_97,In_451,In_183);
xor U98 (N_98,In_583,In_113);
or U99 (N_99,In_352,In_106);
nand U100 (N_100,In_595,In_37);
xor U101 (N_101,In_130,In_623);
and U102 (N_102,In_148,In_368);
or U103 (N_103,In_220,In_53);
and U104 (N_104,In_589,In_518);
nor U105 (N_105,In_279,In_703);
xnor U106 (N_106,In_507,In_18);
or U107 (N_107,In_705,In_464);
xor U108 (N_108,In_384,In_725);
and U109 (N_109,In_291,In_234);
and U110 (N_110,In_9,In_704);
and U111 (N_111,In_677,In_132);
xor U112 (N_112,In_129,In_613);
or U113 (N_113,In_255,In_355);
xnor U114 (N_114,In_22,In_295);
nor U115 (N_115,In_732,In_86);
nand U116 (N_116,In_382,In_311);
or U117 (N_117,In_389,In_548);
nor U118 (N_118,In_214,In_395);
nand U119 (N_119,In_175,In_701);
and U120 (N_120,In_506,In_238);
nor U121 (N_121,In_335,In_373);
or U122 (N_122,In_15,In_47);
nor U123 (N_123,In_167,In_304);
and U124 (N_124,In_453,In_19);
nand U125 (N_125,In_429,In_112);
or U126 (N_126,In_241,In_405);
xnor U127 (N_127,In_200,In_514);
nand U128 (N_128,In_316,In_78);
nor U129 (N_129,In_407,In_152);
or U130 (N_130,In_72,In_739);
nor U131 (N_131,In_264,In_743);
or U132 (N_132,In_208,In_599);
nor U133 (N_133,In_69,In_560);
nor U134 (N_134,In_636,In_108);
and U135 (N_135,In_386,In_487);
nand U136 (N_136,In_133,In_512);
nor U137 (N_137,In_261,In_612);
xnor U138 (N_138,In_656,In_444);
or U139 (N_139,In_521,In_690);
and U140 (N_140,In_710,In_465);
or U141 (N_141,In_517,In_737);
or U142 (N_142,In_82,In_644);
nand U143 (N_143,In_274,In_180);
nor U144 (N_144,In_502,In_542);
xor U145 (N_145,In_522,In_720);
nand U146 (N_146,In_621,In_609);
and U147 (N_147,In_511,In_427);
or U148 (N_148,In_591,In_657);
nand U149 (N_149,In_719,In_90);
xor U150 (N_150,In_92,In_498);
xnor U151 (N_151,In_222,In_276);
and U152 (N_152,In_328,In_556);
or U153 (N_153,In_459,In_376);
xnor U154 (N_154,In_43,In_640);
xnor U155 (N_155,In_281,In_727);
nand U156 (N_156,In_660,In_692);
nand U157 (N_157,In_728,In_394);
nand U158 (N_158,In_249,In_213);
nor U159 (N_159,In_159,In_398);
and U160 (N_160,In_38,In_254);
nand U161 (N_161,In_717,In_449);
xor U162 (N_162,In_588,In_312);
and U163 (N_163,In_381,In_275);
nor U164 (N_164,In_645,In_547);
and U165 (N_165,In_516,In_480);
xnor U166 (N_166,In_478,In_101);
or U167 (N_167,In_145,In_170);
and U168 (N_168,In_94,In_128);
nand U169 (N_169,In_693,In_647);
and U170 (N_170,In_223,In_648);
nor U171 (N_171,In_338,In_411);
or U172 (N_172,In_34,In_578);
or U173 (N_173,In_735,In_608);
or U174 (N_174,In_531,In_163);
and U175 (N_175,In_748,In_219);
nand U176 (N_176,In_323,In_293);
xor U177 (N_177,In_391,In_137);
or U178 (N_178,In_24,In_600);
or U179 (N_179,In_156,In_149);
nand U180 (N_180,In_419,In_593);
or U181 (N_181,In_729,In_315);
nand U182 (N_182,In_251,In_596);
xnor U183 (N_183,In_708,In_598);
and U184 (N_184,In_428,In_606);
xor U185 (N_185,In_224,In_237);
and U186 (N_186,In_269,In_390);
nor U187 (N_187,In_540,In_48);
and U188 (N_188,In_13,In_197);
nor U189 (N_189,In_695,In_320);
or U190 (N_190,In_716,In_83);
and U191 (N_191,In_744,In_337);
nand U192 (N_192,In_64,In_215);
xor U193 (N_193,In_154,In_124);
or U194 (N_194,In_73,In_12);
or U195 (N_195,In_236,In_571);
nand U196 (N_196,In_353,In_722);
nand U197 (N_197,In_545,In_413);
xnor U198 (N_198,In_171,In_54);
nor U199 (N_199,In_423,In_551);
and U200 (N_200,In_576,In_169);
or U201 (N_201,In_515,In_107);
nand U202 (N_202,In_212,In_105);
or U203 (N_203,In_671,In_250);
nor U204 (N_204,In_119,In_365);
and U205 (N_205,In_321,In_466);
nor U206 (N_206,In_661,In_242);
and U207 (N_207,In_202,In_494);
nand U208 (N_208,In_535,In_492);
nand U209 (N_209,In_392,In_404);
or U210 (N_210,In_201,In_687);
xor U211 (N_211,In_294,In_370);
nand U212 (N_212,In_55,In_402);
xor U213 (N_213,In_192,In_721);
and U214 (N_214,In_266,In_62);
xor U215 (N_215,In_259,In_443);
nor U216 (N_216,In_136,In_364);
nor U217 (N_217,In_203,In_610);
and U218 (N_218,In_190,In_162);
nor U219 (N_219,In_292,In_358);
nor U220 (N_220,In_622,In_561);
nand U221 (N_221,In_678,In_745);
nand U222 (N_222,In_527,In_351);
and U223 (N_223,In_436,In_605);
or U224 (N_224,In_60,In_675);
nor U225 (N_225,In_624,In_500);
and U226 (N_226,In_524,In_664);
nand U227 (N_227,In_734,In_519);
nand U228 (N_228,In_262,In_456);
or U229 (N_229,In_573,In_218);
nor U230 (N_230,In_2,In_670);
nor U231 (N_231,In_632,In_143);
nand U232 (N_232,In_322,In_742);
or U233 (N_233,In_414,In_463);
or U234 (N_234,In_654,In_198);
xnor U235 (N_235,In_326,In_26);
and U236 (N_236,In_409,In_747);
nor U237 (N_237,In_490,In_493);
nor U238 (N_238,In_448,In_296);
xnor U239 (N_239,In_349,In_501);
xor U240 (N_240,In_257,In_319);
xor U241 (N_241,In_194,In_77);
nor U242 (N_242,In_460,In_341);
or U243 (N_243,In_417,In_749);
nand U244 (N_244,In_410,In_271);
nor U245 (N_245,In_696,In_594);
nor U246 (N_246,In_684,In_305);
or U247 (N_247,In_74,In_635);
xor U248 (N_248,In_399,In_707);
and U249 (N_249,In_504,In_686);
xor U250 (N_250,In_712,In_3);
xor U251 (N_251,In_699,In_412);
nand U252 (N_252,In_486,In_61);
nand U253 (N_253,In_150,In_303);
nand U254 (N_254,In_655,In_374);
xor U255 (N_255,In_45,In_550);
or U256 (N_256,In_87,In_564);
or U257 (N_257,In_467,In_625);
nand U258 (N_258,In_408,In_420);
nor U259 (N_259,In_6,In_10);
nand U260 (N_260,In_418,In_570);
nand U261 (N_261,In_432,In_538);
xor U262 (N_262,In_284,In_331);
nor U263 (N_263,In_115,In_582);
or U264 (N_264,In_676,In_35);
nand U265 (N_265,In_240,In_611);
or U266 (N_266,In_49,In_174);
xnor U267 (N_267,In_357,In_615);
nand U268 (N_268,In_139,In_617);
or U269 (N_269,In_740,In_658);
nand U270 (N_270,In_473,In_216);
xor U271 (N_271,In_426,In_488);
xnor U272 (N_272,In_715,In_340);
xor U273 (N_273,In_288,In_40);
nand U274 (N_274,In_659,In_587);
xnor U275 (N_275,In_260,In_233);
nor U276 (N_276,In_314,In_652);
nor U277 (N_277,In_93,In_422);
or U278 (N_278,In_629,In_698);
xnor U279 (N_279,In_185,In_127);
nand U280 (N_280,In_20,In_706);
xnor U281 (N_281,In_590,In_88);
xor U282 (N_282,In_51,In_181);
and U283 (N_283,In_110,In_665);
nor U284 (N_284,In_151,In_733);
nor U285 (N_285,In_52,In_96);
xnor U286 (N_286,In_199,In_290);
or U287 (N_287,In_536,In_36);
and U288 (N_288,In_663,In_607);
nand U289 (N_289,In_146,In_243);
and U290 (N_290,In_700,In_361);
and U291 (N_291,In_496,In_325);
nor U292 (N_292,In_569,In_344);
xor U293 (N_293,In_689,In_483);
and U294 (N_294,In_46,In_375);
xor U295 (N_295,In_379,In_520);
and U296 (N_296,In_138,In_161);
nand U297 (N_297,In_714,In_602);
or U298 (N_298,In_484,In_28);
nor U299 (N_299,In_176,In_21);
nor U300 (N_300,In_683,In_318);
and U301 (N_301,In_32,In_187);
nand U302 (N_302,In_168,In_70);
and U303 (N_303,In_442,In_39);
nand U304 (N_304,In_472,In_317);
and U305 (N_305,In_307,In_299);
nand U306 (N_306,In_702,In_489);
and U307 (N_307,In_440,In_278);
nor U308 (N_308,In_141,In_252);
nand U309 (N_309,In_297,In_4);
xor U310 (N_310,In_273,In_95);
or U311 (N_311,In_592,In_508);
nand U312 (N_312,In_618,In_306);
nand U313 (N_313,In_393,In_479);
and U314 (N_314,In_433,In_348);
nand U315 (N_315,In_380,In_680);
nor U316 (N_316,In_217,In_533);
or U317 (N_317,In_302,In_17);
nor U318 (N_318,In_158,In_539);
or U319 (N_319,In_377,In_76);
xor U320 (N_320,In_313,In_33);
nand U321 (N_321,In_144,In_499);
nand U322 (N_322,In_558,In_474);
nor U323 (N_323,In_342,In_468);
or U324 (N_324,In_289,In_125);
xor U325 (N_325,In_270,In_42);
nand U326 (N_326,In_165,In_231);
nand U327 (N_327,In_565,In_694);
nand U328 (N_328,In_639,In_157);
nand U329 (N_329,In_369,In_438);
nor U330 (N_330,In_513,In_567);
or U331 (N_331,In_287,In_122);
or U332 (N_332,In_332,In_191);
nand U333 (N_333,In_585,In_230);
xnor U334 (N_334,In_396,In_580);
and U335 (N_335,In_57,In_403);
nor U336 (N_336,In_682,In_166);
or U337 (N_337,In_164,In_272);
and U338 (N_338,In_111,In_718);
and U339 (N_339,In_239,In_650);
nor U340 (N_340,In_668,In_126);
nand U341 (N_341,In_188,In_89);
nand U342 (N_342,In_546,In_738);
and U343 (N_343,In_387,In_503);
nor U344 (N_344,In_142,In_0);
nand U345 (N_345,In_116,In_372);
nor U346 (N_346,In_246,In_425);
or U347 (N_347,In_482,In_330);
nor U348 (N_348,In_646,In_310);
and U349 (N_349,In_709,In_681);
nand U350 (N_350,In_471,In_1);
nor U351 (N_351,In_286,In_67);
nand U352 (N_352,In_383,In_562);
nor U353 (N_353,In_685,In_178);
xnor U354 (N_354,In_245,In_430);
and U355 (N_355,In_81,In_334);
and U356 (N_356,In_225,In_532);
xnor U357 (N_357,In_679,In_526);
nand U358 (N_358,In_253,In_674);
and U359 (N_359,In_572,In_552);
nand U360 (N_360,In_56,In_309);
and U361 (N_361,In_59,In_649);
nor U362 (N_362,In_509,In_182);
or U363 (N_363,In_614,In_186);
nor U364 (N_364,In_283,In_601);
xnor U365 (N_365,In_98,In_653);
nor U366 (N_366,In_263,In_439);
xor U367 (N_367,In_530,In_566);
or U368 (N_368,In_16,In_691);
and U369 (N_369,In_445,In_529);
nand U370 (N_370,In_160,In_638);
nor U371 (N_371,In_280,In_63);
or U372 (N_372,In_568,In_581);
and U373 (N_373,In_248,In_455);
or U374 (N_374,In_11,In_123);
and U375 (N_375,In_562,In_657);
nor U376 (N_376,In_7,In_330);
nand U377 (N_377,In_428,In_43);
xor U378 (N_378,In_86,In_98);
and U379 (N_379,In_64,In_60);
and U380 (N_380,In_703,In_611);
or U381 (N_381,In_20,In_424);
or U382 (N_382,In_661,In_390);
or U383 (N_383,In_78,In_676);
nor U384 (N_384,In_67,In_582);
nand U385 (N_385,In_69,In_457);
and U386 (N_386,In_493,In_495);
or U387 (N_387,In_82,In_105);
and U388 (N_388,In_592,In_661);
and U389 (N_389,In_389,In_511);
nor U390 (N_390,In_528,In_145);
and U391 (N_391,In_598,In_258);
nand U392 (N_392,In_623,In_220);
nand U393 (N_393,In_109,In_473);
nor U394 (N_394,In_240,In_287);
xnor U395 (N_395,In_130,In_413);
xnor U396 (N_396,In_37,In_217);
xnor U397 (N_397,In_496,In_389);
or U398 (N_398,In_609,In_152);
and U399 (N_399,In_626,In_326);
xor U400 (N_400,In_86,In_667);
nand U401 (N_401,In_74,In_661);
nand U402 (N_402,In_625,In_427);
and U403 (N_403,In_451,In_495);
nor U404 (N_404,In_178,In_186);
nor U405 (N_405,In_468,In_709);
xnor U406 (N_406,In_393,In_728);
nand U407 (N_407,In_79,In_206);
nand U408 (N_408,In_394,In_559);
or U409 (N_409,In_486,In_96);
nand U410 (N_410,In_156,In_638);
xor U411 (N_411,In_159,In_585);
nor U412 (N_412,In_342,In_702);
xor U413 (N_413,In_136,In_384);
xor U414 (N_414,In_453,In_721);
and U415 (N_415,In_742,In_665);
xor U416 (N_416,In_390,In_683);
nor U417 (N_417,In_747,In_359);
xor U418 (N_418,In_397,In_338);
or U419 (N_419,In_26,In_678);
nand U420 (N_420,In_498,In_652);
or U421 (N_421,In_586,In_77);
xnor U422 (N_422,In_333,In_518);
nor U423 (N_423,In_217,In_137);
xor U424 (N_424,In_277,In_70);
and U425 (N_425,In_172,In_494);
nand U426 (N_426,In_302,In_271);
nor U427 (N_427,In_8,In_632);
or U428 (N_428,In_28,In_72);
nor U429 (N_429,In_194,In_276);
and U430 (N_430,In_723,In_506);
xor U431 (N_431,In_134,In_9);
xnor U432 (N_432,In_268,In_674);
or U433 (N_433,In_298,In_568);
nand U434 (N_434,In_202,In_648);
nor U435 (N_435,In_234,In_373);
xor U436 (N_436,In_463,In_608);
nor U437 (N_437,In_580,In_451);
xnor U438 (N_438,In_566,In_725);
or U439 (N_439,In_710,In_413);
and U440 (N_440,In_715,In_368);
nor U441 (N_441,In_366,In_484);
nand U442 (N_442,In_131,In_332);
xnor U443 (N_443,In_542,In_654);
and U444 (N_444,In_522,In_321);
nand U445 (N_445,In_491,In_681);
nor U446 (N_446,In_389,In_450);
nor U447 (N_447,In_221,In_257);
nor U448 (N_448,In_58,In_464);
xnor U449 (N_449,In_214,In_507);
nor U450 (N_450,In_375,In_489);
or U451 (N_451,In_461,In_577);
and U452 (N_452,In_376,In_415);
xor U453 (N_453,In_525,In_154);
xor U454 (N_454,In_192,In_492);
or U455 (N_455,In_578,In_663);
nor U456 (N_456,In_152,In_28);
and U457 (N_457,In_255,In_38);
nor U458 (N_458,In_676,In_355);
nor U459 (N_459,In_502,In_321);
nor U460 (N_460,In_276,In_445);
xor U461 (N_461,In_164,In_45);
and U462 (N_462,In_333,In_47);
or U463 (N_463,In_366,In_590);
and U464 (N_464,In_247,In_599);
nor U465 (N_465,In_242,In_113);
nand U466 (N_466,In_153,In_387);
nand U467 (N_467,In_443,In_10);
or U468 (N_468,In_30,In_572);
nor U469 (N_469,In_580,In_521);
xor U470 (N_470,In_376,In_579);
nor U471 (N_471,In_331,In_348);
nor U472 (N_472,In_111,In_245);
nand U473 (N_473,In_547,In_677);
nor U474 (N_474,In_466,In_454);
or U475 (N_475,In_91,In_612);
or U476 (N_476,In_561,In_91);
xor U477 (N_477,In_159,In_391);
xor U478 (N_478,In_229,In_516);
xor U479 (N_479,In_746,In_693);
and U480 (N_480,In_412,In_508);
xnor U481 (N_481,In_245,In_467);
nor U482 (N_482,In_690,In_142);
nand U483 (N_483,In_46,In_720);
nor U484 (N_484,In_467,In_513);
and U485 (N_485,In_206,In_354);
xor U486 (N_486,In_530,In_349);
xnor U487 (N_487,In_648,In_54);
nand U488 (N_488,In_114,In_605);
xnor U489 (N_489,In_519,In_195);
or U490 (N_490,In_671,In_583);
nor U491 (N_491,In_273,In_602);
or U492 (N_492,In_530,In_631);
or U493 (N_493,In_151,In_282);
or U494 (N_494,In_519,In_664);
xor U495 (N_495,In_399,In_5);
and U496 (N_496,In_296,In_615);
nor U497 (N_497,In_215,In_71);
and U498 (N_498,In_472,In_538);
xnor U499 (N_499,In_627,In_80);
or U500 (N_500,N_193,N_154);
nor U501 (N_501,N_184,N_471);
and U502 (N_502,N_452,N_54);
and U503 (N_503,N_389,N_287);
or U504 (N_504,N_370,N_71);
xnor U505 (N_505,N_31,N_375);
xnor U506 (N_506,N_487,N_464);
xnor U507 (N_507,N_415,N_147);
and U508 (N_508,N_278,N_355);
xor U509 (N_509,N_4,N_8);
nand U510 (N_510,N_148,N_334);
xor U511 (N_511,N_99,N_77);
or U512 (N_512,N_27,N_199);
nand U513 (N_513,N_50,N_35);
nor U514 (N_514,N_243,N_407);
nand U515 (N_515,N_343,N_436);
nor U516 (N_516,N_203,N_476);
and U517 (N_517,N_52,N_222);
or U518 (N_518,N_411,N_107);
xor U519 (N_519,N_49,N_105);
and U520 (N_520,N_316,N_362);
and U521 (N_521,N_311,N_272);
nand U522 (N_522,N_96,N_372);
nor U523 (N_523,N_220,N_44);
and U524 (N_524,N_22,N_92);
xnor U525 (N_525,N_251,N_142);
xnor U526 (N_526,N_84,N_442);
nor U527 (N_527,N_339,N_238);
xnor U528 (N_528,N_26,N_25);
or U529 (N_529,N_421,N_366);
nand U530 (N_530,N_448,N_10);
and U531 (N_531,N_161,N_80);
nor U532 (N_532,N_270,N_379);
or U533 (N_533,N_498,N_133);
xor U534 (N_534,N_43,N_174);
and U535 (N_535,N_100,N_446);
nand U536 (N_536,N_115,N_239);
xor U537 (N_537,N_242,N_479);
and U538 (N_538,N_273,N_202);
xnor U539 (N_539,N_126,N_81);
xor U540 (N_540,N_469,N_201);
xnor U541 (N_541,N_283,N_117);
or U542 (N_542,N_23,N_228);
nand U543 (N_543,N_336,N_56);
xor U544 (N_544,N_300,N_269);
and U545 (N_545,N_268,N_231);
nand U546 (N_546,N_337,N_227);
xor U547 (N_547,N_424,N_91);
nor U548 (N_548,N_419,N_150);
nor U549 (N_549,N_262,N_134);
and U550 (N_550,N_356,N_417);
xnor U551 (N_551,N_474,N_445);
or U552 (N_552,N_408,N_219);
nand U553 (N_553,N_63,N_176);
nor U554 (N_554,N_348,N_431);
nor U555 (N_555,N_40,N_266);
nand U556 (N_556,N_392,N_21);
and U557 (N_557,N_47,N_151);
or U558 (N_558,N_194,N_149);
nor U559 (N_559,N_37,N_158);
and U560 (N_560,N_324,N_102);
xnor U561 (N_561,N_470,N_156);
and U562 (N_562,N_76,N_236);
nor U563 (N_563,N_332,N_214);
nand U564 (N_564,N_490,N_457);
xor U565 (N_565,N_247,N_205);
and U566 (N_566,N_108,N_323);
or U567 (N_567,N_240,N_128);
nor U568 (N_568,N_259,N_489);
nor U569 (N_569,N_265,N_131);
or U570 (N_570,N_24,N_388);
and U571 (N_571,N_465,N_341);
or U572 (N_572,N_17,N_472);
and U573 (N_573,N_123,N_364);
and U574 (N_574,N_101,N_297);
xor U575 (N_575,N_20,N_305);
or U576 (N_576,N_313,N_314);
or U577 (N_577,N_74,N_488);
nor U578 (N_578,N_499,N_182);
or U579 (N_579,N_145,N_136);
xnor U580 (N_580,N_260,N_475);
or U581 (N_581,N_478,N_312);
xnor U582 (N_582,N_274,N_124);
and U583 (N_583,N_138,N_327);
or U584 (N_584,N_98,N_252);
xor U585 (N_585,N_42,N_118);
and U586 (N_586,N_181,N_65);
and U587 (N_587,N_59,N_127);
xor U588 (N_588,N_458,N_144);
xnor U589 (N_589,N_288,N_85);
nor U590 (N_590,N_30,N_468);
or U591 (N_591,N_335,N_432);
or U592 (N_592,N_234,N_284);
nand U593 (N_593,N_382,N_331);
nand U594 (N_594,N_109,N_387);
nor U595 (N_595,N_462,N_319);
nand U596 (N_596,N_394,N_285);
and U597 (N_597,N_157,N_215);
nor U598 (N_598,N_122,N_376);
and U599 (N_599,N_427,N_310);
xnor U600 (N_600,N_32,N_38);
and U601 (N_601,N_106,N_90);
and U602 (N_602,N_33,N_152);
and U603 (N_603,N_422,N_466);
nand U604 (N_604,N_248,N_12);
nand U605 (N_605,N_195,N_481);
nand U606 (N_606,N_164,N_218);
nand U607 (N_607,N_433,N_358);
and U608 (N_608,N_400,N_280);
xnor U609 (N_609,N_19,N_221);
xnor U610 (N_610,N_328,N_253);
xnor U611 (N_611,N_79,N_226);
or U612 (N_612,N_275,N_380);
or U613 (N_613,N_2,N_70);
and U614 (N_614,N_429,N_344);
or U615 (N_615,N_349,N_196);
or U616 (N_616,N_350,N_346);
xor U617 (N_617,N_204,N_453);
or U618 (N_618,N_383,N_290);
nand U619 (N_619,N_111,N_325);
and U620 (N_620,N_423,N_347);
nor U621 (N_621,N_317,N_121);
and U622 (N_622,N_351,N_303);
xor U623 (N_623,N_271,N_82);
or U624 (N_624,N_75,N_493);
and U625 (N_625,N_94,N_291);
nand U626 (N_626,N_463,N_398);
xnor U627 (N_627,N_454,N_345);
or U628 (N_628,N_83,N_413);
xor U629 (N_629,N_57,N_404);
nor U630 (N_630,N_73,N_104);
nand U631 (N_631,N_170,N_449);
or U632 (N_632,N_456,N_267);
xor U633 (N_633,N_360,N_377);
nand U634 (N_634,N_373,N_261);
xor U635 (N_635,N_330,N_307);
nand U636 (N_636,N_321,N_48);
nor U637 (N_637,N_235,N_494);
and U638 (N_638,N_420,N_492);
nor U639 (N_639,N_229,N_318);
nand U640 (N_640,N_301,N_390);
or U641 (N_641,N_14,N_114);
nor U642 (N_642,N_485,N_414);
or U643 (N_643,N_246,N_187);
or U644 (N_644,N_166,N_257);
nand U645 (N_645,N_224,N_61);
or U646 (N_646,N_9,N_13);
xnor U647 (N_647,N_385,N_153);
xnor U648 (N_648,N_233,N_441);
nor U649 (N_649,N_244,N_396);
nand U650 (N_650,N_403,N_120);
nand U651 (N_651,N_207,N_18);
nand U652 (N_652,N_258,N_64);
nor U653 (N_653,N_217,N_125);
or U654 (N_654,N_165,N_338);
or U655 (N_655,N_188,N_369);
nand U656 (N_656,N_173,N_294);
and U657 (N_657,N_254,N_447);
nor U658 (N_658,N_140,N_329);
nor U659 (N_659,N_354,N_16);
or U660 (N_660,N_146,N_1);
nand U661 (N_661,N_46,N_340);
xnor U662 (N_662,N_160,N_298);
nor U663 (N_663,N_11,N_15);
nand U664 (N_664,N_393,N_486);
or U665 (N_665,N_402,N_88);
or U666 (N_666,N_3,N_212);
nand U667 (N_667,N_178,N_384);
nand U668 (N_668,N_304,N_342);
nor U669 (N_669,N_333,N_455);
and U670 (N_670,N_282,N_352);
or U671 (N_671,N_51,N_353);
nor U672 (N_672,N_36,N_289);
xnor U673 (N_673,N_116,N_263);
or U674 (N_674,N_302,N_119);
xor U675 (N_675,N_216,N_34);
nor U676 (N_676,N_418,N_295);
or U677 (N_677,N_6,N_249);
and U678 (N_678,N_361,N_296);
and U679 (N_679,N_60,N_281);
and U680 (N_680,N_484,N_443);
or U681 (N_681,N_168,N_155);
and U682 (N_682,N_135,N_45);
or U683 (N_683,N_477,N_129);
xnor U684 (N_684,N_211,N_172);
nor U685 (N_685,N_132,N_78);
and U686 (N_686,N_286,N_189);
and U687 (N_687,N_409,N_198);
nor U688 (N_688,N_264,N_395);
and U689 (N_689,N_179,N_460);
xor U690 (N_690,N_137,N_496);
nand U691 (N_691,N_190,N_357);
or U692 (N_692,N_112,N_191);
or U693 (N_693,N_175,N_210);
or U694 (N_694,N_276,N_167);
or U695 (N_695,N_497,N_171);
nand U696 (N_696,N_28,N_482);
xor U697 (N_697,N_7,N_237);
nor U698 (N_698,N_438,N_143);
xnor U699 (N_699,N_208,N_322);
and U700 (N_700,N_169,N_130);
or U701 (N_701,N_425,N_401);
nand U702 (N_702,N_39,N_359);
and U703 (N_703,N_292,N_97);
nor U704 (N_704,N_491,N_58);
and U705 (N_705,N_406,N_277);
and U706 (N_706,N_225,N_89);
or U707 (N_707,N_439,N_186);
xor U708 (N_708,N_180,N_86);
xnor U709 (N_709,N_430,N_177);
xor U710 (N_710,N_440,N_426);
nor U711 (N_711,N_223,N_68);
xor U712 (N_712,N_110,N_279);
and U713 (N_713,N_256,N_374);
nor U714 (N_714,N_206,N_435);
nand U715 (N_715,N_192,N_451);
xor U716 (N_716,N_480,N_66);
or U717 (N_717,N_232,N_399);
nor U718 (N_718,N_391,N_209);
and U719 (N_719,N_381,N_363);
nor U720 (N_720,N_473,N_365);
nand U721 (N_721,N_245,N_326);
xnor U722 (N_722,N_241,N_87);
xnor U723 (N_723,N_320,N_162);
or U724 (N_724,N_467,N_299);
xnor U725 (N_725,N_306,N_62);
and U726 (N_726,N_428,N_213);
xor U727 (N_727,N_29,N_5);
xor U728 (N_728,N_67,N_405);
nor U729 (N_729,N_163,N_434);
nor U730 (N_730,N_185,N_410);
nand U731 (N_731,N_412,N_386);
xnor U732 (N_732,N_293,N_437);
or U733 (N_733,N_444,N_141);
and U734 (N_734,N_93,N_309);
nand U735 (N_735,N_368,N_95);
nand U736 (N_736,N_450,N_495);
and U737 (N_737,N_183,N_371);
xnor U738 (N_738,N_139,N_308);
nand U739 (N_739,N_113,N_55);
or U740 (N_740,N_72,N_0);
nand U741 (N_741,N_397,N_378);
xor U742 (N_742,N_459,N_197);
or U743 (N_743,N_250,N_41);
and U744 (N_744,N_200,N_69);
and U745 (N_745,N_255,N_416);
xor U746 (N_746,N_53,N_367);
and U747 (N_747,N_483,N_315);
nand U748 (N_748,N_461,N_230);
or U749 (N_749,N_159,N_103);
nand U750 (N_750,N_312,N_31);
nand U751 (N_751,N_176,N_297);
nand U752 (N_752,N_452,N_496);
and U753 (N_753,N_107,N_401);
nand U754 (N_754,N_169,N_338);
nor U755 (N_755,N_60,N_318);
nand U756 (N_756,N_37,N_305);
nor U757 (N_757,N_30,N_145);
xnor U758 (N_758,N_254,N_367);
xnor U759 (N_759,N_35,N_409);
or U760 (N_760,N_342,N_98);
or U761 (N_761,N_492,N_232);
and U762 (N_762,N_255,N_128);
nand U763 (N_763,N_497,N_123);
nand U764 (N_764,N_313,N_358);
nor U765 (N_765,N_497,N_163);
nand U766 (N_766,N_375,N_48);
and U767 (N_767,N_13,N_314);
nor U768 (N_768,N_37,N_269);
and U769 (N_769,N_210,N_121);
and U770 (N_770,N_38,N_412);
nand U771 (N_771,N_197,N_380);
or U772 (N_772,N_152,N_362);
or U773 (N_773,N_457,N_280);
nand U774 (N_774,N_486,N_189);
nand U775 (N_775,N_431,N_393);
and U776 (N_776,N_469,N_174);
xnor U777 (N_777,N_196,N_404);
or U778 (N_778,N_84,N_52);
nand U779 (N_779,N_112,N_213);
or U780 (N_780,N_56,N_26);
nand U781 (N_781,N_195,N_312);
nand U782 (N_782,N_415,N_12);
xnor U783 (N_783,N_338,N_212);
nor U784 (N_784,N_246,N_404);
or U785 (N_785,N_358,N_131);
and U786 (N_786,N_105,N_482);
or U787 (N_787,N_127,N_164);
and U788 (N_788,N_403,N_303);
xor U789 (N_789,N_315,N_3);
and U790 (N_790,N_196,N_357);
nor U791 (N_791,N_179,N_94);
or U792 (N_792,N_305,N_348);
and U793 (N_793,N_402,N_395);
nand U794 (N_794,N_159,N_24);
xnor U795 (N_795,N_107,N_494);
and U796 (N_796,N_67,N_476);
nor U797 (N_797,N_454,N_255);
and U798 (N_798,N_437,N_390);
and U799 (N_799,N_183,N_458);
and U800 (N_800,N_448,N_147);
nand U801 (N_801,N_469,N_69);
and U802 (N_802,N_39,N_417);
xor U803 (N_803,N_189,N_197);
nor U804 (N_804,N_87,N_52);
nor U805 (N_805,N_25,N_280);
and U806 (N_806,N_400,N_261);
nor U807 (N_807,N_405,N_72);
nand U808 (N_808,N_369,N_398);
or U809 (N_809,N_74,N_499);
nor U810 (N_810,N_209,N_31);
or U811 (N_811,N_50,N_186);
or U812 (N_812,N_276,N_137);
xor U813 (N_813,N_79,N_493);
or U814 (N_814,N_16,N_326);
nor U815 (N_815,N_241,N_263);
xnor U816 (N_816,N_343,N_335);
and U817 (N_817,N_249,N_47);
xnor U818 (N_818,N_37,N_150);
or U819 (N_819,N_157,N_153);
and U820 (N_820,N_32,N_460);
nor U821 (N_821,N_250,N_499);
xor U822 (N_822,N_55,N_197);
and U823 (N_823,N_385,N_482);
or U824 (N_824,N_361,N_367);
nor U825 (N_825,N_333,N_145);
or U826 (N_826,N_433,N_340);
xnor U827 (N_827,N_301,N_77);
nor U828 (N_828,N_178,N_73);
and U829 (N_829,N_153,N_23);
nor U830 (N_830,N_17,N_289);
or U831 (N_831,N_403,N_456);
or U832 (N_832,N_468,N_282);
nand U833 (N_833,N_161,N_490);
nand U834 (N_834,N_328,N_479);
xor U835 (N_835,N_2,N_429);
or U836 (N_836,N_116,N_107);
or U837 (N_837,N_254,N_15);
or U838 (N_838,N_206,N_434);
or U839 (N_839,N_173,N_284);
xor U840 (N_840,N_436,N_167);
nor U841 (N_841,N_379,N_103);
nand U842 (N_842,N_23,N_349);
xor U843 (N_843,N_473,N_461);
or U844 (N_844,N_52,N_246);
and U845 (N_845,N_226,N_259);
and U846 (N_846,N_187,N_81);
nor U847 (N_847,N_186,N_221);
and U848 (N_848,N_312,N_197);
nand U849 (N_849,N_280,N_445);
or U850 (N_850,N_163,N_212);
nand U851 (N_851,N_152,N_326);
nand U852 (N_852,N_446,N_184);
nor U853 (N_853,N_302,N_178);
nand U854 (N_854,N_414,N_296);
or U855 (N_855,N_30,N_265);
xor U856 (N_856,N_29,N_488);
and U857 (N_857,N_365,N_190);
xnor U858 (N_858,N_28,N_103);
nor U859 (N_859,N_437,N_255);
nor U860 (N_860,N_108,N_392);
or U861 (N_861,N_361,N_182);
and U862 (N_862,N_182,N_385);
nor U863 (N_863,N_173,N_299);
nand U864 (N_864,N_213,N_79);
or U865 (N_865,N_61,N_268);
nor U866 (N_866,N_269,N_294);
nor U867 (N_867,N_285,N_244);
or U868 (N_868,N_240,N_70);
or U869 (N_869,N_138,N_228);
xnor U870 (N_870,N_276,N_375);
nand U871 (N_871,N_383,N_254);
and U872 (N_872,N_495,N_242);
and U873 (N_873,N_257,N_17);
nand U874 (N_874,N_313,N_79);
nor U875 (N_875,N_213,N_65);
and U876 (N_876,N_45,N_224);
xnor U877 (N_877,N_240,N_173);
nand U878 (N_878,N_113,N_32);
or U879 (N_879,N_219,N_409);
nand U880 (N_880,N_407,N_441);
nor U881 (N_881,N_54,N_252);
nand U882 (N_882,N_13,N_97);
xor U883 (N_883,N_285,N_67);
and U884 (N_884,N_493,N_221);
nand U885 (N_885,N_266,N_160);
or U886 (N_886,N_140,N_45);
or U887 (N_887,N_343,N_487);
or U888 (N_888,N_51,N_72);
or U889 (N_889,N_328,N_239);
and U890 (N_890,N_159,N_44);
and U891 (N_891,N_20,N_78);
nor U892 (N_892,N_270,N_126);
nor U893 (N_893,N_450,N_229);
or U894 (N_894,N_278,N_362);
nor U895 (N_895,N_275,N_466);
nor U896 (N_896,N_390,N_268);
nand U897 (N_897,N_422,N_1);
nor U898 (N_898,N_350,N_362);
or U899 (N_899,N_289,N_464);
nor U900 (N_900,N_365,N_146);
xor U901 (N_901,N_242,N_432);
nor U902 (N_902,N_499,N_73);
and U903 (N_903,N_191,N_153);
nand U904 (N_904,N_428,N_141);
nand U905 (N_905,N_50,N_80);
or U906 (N_906,N_337,N_452);
nand U907 (N_907,N_444,N_58);
xor U908 (N_908,N_371,N_111);
or U909 (N_909,N_451,N_339);
nand U910 (N_910,N_156,N_64);
and U911 (N_911,N_58,N_214);
xor U912 (N_912,N_247,N_310);
nor U913 (N_913,N_228,N_476);
nand U914 (N_914,N_285,N_308);
or U915 (N_915,N_196,N_191);
and U916 (N_916,N_230,N_304);
nor U917 (N_917,N_430,N_167);
nor U918 (N_918,N_113,N_154);
nor U919 (N_919,N_22,N_352);
xnor U920 (N_920,N_276,N_347);
nor U921 (N_921,N_21,N_120);
xnor U922 (N_922,N_113,N_245);
nand U923 (N_923,N_179,N_102);
xor U924 (N_924,N_35,N_378);
nand U925 (N_925,N_328,N_463);
or U926 (N_926,N_184,N_43);
or U927 (N_927,N_185,N_130);
xor U928 (N_928,N_191,N_471);
nor U929 (N_929,N_419,N_9);
and U930 (N_930,N_154,N_15);
nor U931 (N_931,N_370,N_309);
xnor U932 (N_932,N_277,N_294);
or U933 (N_933,N_200,N_117);
or U934 (N_934,N_297,N_222);
xnor U935 (N_935,N_479,N_154);
nor U936 (N_936,N_325,N_493);
nor U937 (N_937,N_142,N_483);
nor U938 (N_938,N_176,N_324);
nor U939 (N_939,N_326,N_230);
or U940 (N_940,N_138,N_78);
and U941 (N_941,N_251,N_235);
nor U942 (N_942,N_141,N_150);
and U943 (N_943,N_91,N_360);
or U944 (N_944,N_321,N_7);
xor U945 (N_945,N_233,N_13);
xnor U946 (N_946,N_493,N_226);
or U947 (N_947,N_420,N_236);
nor U948 (N_948,N_403,N_461);
nor U949 (N_949,N_6,N_349);
xor U950 (N_950,N_174,N_419);
nor U951 (N_951,N_263,N_35);
or U952 (N_952,N_351,N_83);
and U953 (N_953,N_460,N_3);
or U954 (N_954,N_158,N_150);
nor U955 (N_955,N_417,N_18);
and U956 (N_956,N_214,N_383);
nand U957 (N_957,N_58,N_459);
nand U958 (N_958,N_293,N_140);
nand U959 (N_959,N_483,N_114);
and U960 (N_960,N_482,N_197);
nor U961 (N_961,N_155,N_167);
nor U962 (N_962,N_349,N_45);
nand U963 (N_963,N_375,N_229);
nand U964 (N_964,N_126,N_498);
and U965 (N_965,N_195,N_417);
nand U966 (N_966,N_390,N_348);
or U967 (N_967,N_376,N_217);
or U968 (N_968,N_124,N_337);
nor U969 (N_969,N_401,N_417);
nor U970 (N_970,N_146,N_201);
and U971 (N_971,N_118,N_20);
nor U972 (N_972,N_372,N_93);
or U973 (N_973,N_418,N_57);
xor U974 (N_974,N_266,N_79);
xor U975 (N_975,N_493,N_383);
and U976 (N_976,N_361,N_359);
or U977 (N_977,N_331,N_252);
or U978 (N_978,N_304,N_365);
and U979 (N_979,N_404,N_221);
nor U980 (N_980,N_113,N_226);
nand U981 (N_981,N_329,N_89);
xor U982 (N_982,N_439,N_309);
and U983 (N_983,N_21,N_412);
and U984 (N_984,N_98,N_478);
or U985 (N_985,N_36,N_227);
nand U986 (N_986,N_57,N_246);
or U987 (N_987,N_229,N_476);
and U988 (N_988,N_319,N_278);
nand U989 (N_989,N_80,N_119);
nand U990 (N_990,N_143,N_497);
xor U991 (N_991,N_486,N_165);
nor U992 (N_992,N_452,N_495);
and U993 (N_993,N_230,N_281);
or U994 (N_994,N_89,N_221);
or U995 (N_995,N_44,N_1);
or U996 (N_996,N_471,N_96);
xor U997 (N_997,N_26,N_67);
xnor U998 (N_998,N_173,N_275);
xor U999 (N_999,N_353,N_45);
nor U1000 (N_1000,N_742,N_981);
or U1001 (N_1001,N_892,N_540);
or U1002 (N_1002,N_754,N_854);
nor U1003 (N_1003,N_746,N_618);
and U1004 (N_1004,N_897,N_721);
and U1005 (N_1005,N_913,N_708);
nor U1006 (N_1006,N_557,N_640);
nor U1007 (N_1007,N_703,N_979);
or U1008 (N_1008,N_598,N_907);
or U1009 (N_1009,N_728,N_995);
and U1010 (N_1010,N_926,N_554);
nor U1011 (N_1011,N_610,N_553);
or U1012 (N_1012,N_881,N_857);
nor U1013 (N_1013,N_918,N_645);
or U1014 (N_1014,N_582,N_593);
and U1015 (N_1015,N_562,N_823);
nor U1016 (N_1016,N_501,N_960);
or U1017 (N_1017,N_758,N_595);
and U1018 (N_1018,N_832,N_987);
or U1019 (N_1019,N_513,N_886);
and U1020 (N_1020,N_503,N_500);
nor U1021 (N_1021,N_769,N_580);
and U1022 (N_1022,N_661,N_508);
nor U1023 (N_1023,N_871,N_851);
nand U1024 (N_1024,N_510,N_826);
and U1025 (N_1025,N_620,N_831);
nor U1026 (N_1026,N_938,N_504);
or U1027 (N_1027,N_570,N_560);
or U1028 (N_1028,N_704,N_777);
nor U1029 (N_1029,N_646,N_901);
or U1030 (N_1030,N_741,N_818);
xnor U1031 (N_1031,N_759,N_577);
nor U1032 (N_1032,N_914,N_958);
and U1033 (N_1033,N_942,N_968);
or U1034 (N_1034,N_575,N_633);
nand U1035 (N_1035,N_675,N_530);
nand U1036 (N_1036,N_541,N_651);
and U1037 (N_1037,N_966,N_507);
nand U1038 (N_1038,N_714,N_883);
xnor U1039 (N_1039,N_970,N_853);
or U1040 (N_1040,N_889,N_719);
nor U1041 (N_1041,N_764,N_855);
or U1042 (N_1042,N_794,N_757);
xnor U1043 (N_1043,N_910,N_574);
nand U1044 (N_1044,N_511,N_877);
and U1045 (N_1045,N_864,N_845);
nor U1046 (N_1046,N_969,N_543);
or U1047 (N_1047,N_706,N_967);
or U1048 (N_1048,N_590,N_928);
nor U1049 (N_1049,N_506,N_639);
or U1050 (N_1050,N_898,N_959);
nand U1051 (N_1051,N_996,N_989);
xnor U1052 (N_1052,N_576,N_735);
xnor U1053 (N_1053,N_802,N_890);
nor U1054 (N_1054,N_803,N_626);
nor U1055 (N_1055,N_748,N_895);
xor U1056 (N_1056,N_672,N_584);
and U1057 (N_1057,N_668,N_678);
nor U1058 (N_1058,N_887,N_698);
or U1059 (N_1059,N_791,N_781);
xnor U1060 (N_1060,N_819,N_502);
xor U1061 (N_1061,N_896,N_600);
xor U1062 (N_1062,N_662,N_726);
nand U1063 (N_1063,N_520,N_863);
xor U1064 (N_1064,N_624,N_829);
xor U1065 (N_1065,N_964,N_977);
and U1066 (N_1066,N_788,N_866);
xor U1067 (N_1067,N_786,N_596);
and U1068 (N_1068,N_603,N_933);
or U1069 (N_1069,N_924,N_982);
xor U1070 (N_1070,N_556,N_986);
nor U1071 (N_1071,N_643,N_566);
xnor U1072 (N_1072,N_806,N_800);
and U1073 (N_1073,N_840,N_985);
xor U1074 (N_1074,N_691,N_619);
or U1075 (N_1075,N_974,N_921);
nand U1076 (N_1076,N_711,N_822);
xnor U1077 (N_1077,N_515,N_909);
nor U1078 (N_1078,N_767,N_707);
nor U1079 (N_1079,N_911,N_992);
nor U1080 (N_1080,N_531,N_546);
or U1081 (N_1081,N_874,N_940);
or U1082 (N_1082,N_848,N_903);
nand U1083 (N_1083,N_597,N_649);
and U1084 (N_1084,N_528,N_518);
xor U1085 (N_1085,N_875,N_688);
nand U1086 (N_1086,N_749,N_779);
nor U1087 (N_1087,N_664,N_994);
and U1088 (N_1088,N_984,N_789);
nand U1089 (N_1089,N_718,N_931);
nor U1090 (N_1090,N_569,N_941);
nand U1091 (N_1091,N_867,N_768);
or U1092 (N_1092,N_955,N_542);
nand U1093 (N_1093,N_812,N_573);
nor U1094 (N_1094,N_865,N_923);
or U1095 (N_1095,N_745,N_568);
xor U1096 (N_1096,N_734,N_730);
nand U1097 (N_1097,N_844,N_731);
and U1098 (N_1098,N_551,N_747);
or U1099 (N_1099,N_548,N_642);
or U1100 (N_1100,N_689,N_519);
nand U1101 (N_1101,N_930,N_717);
and U1102 (N_1102,N_801,N_656);
xor U1103 (N_1103,N_771,N_760);
nor U1104 (N_1104,N_808,N_740);
nor U1105 (N_1105,N_505,N_677);
or U1106 (N_1106,N_919,N_699);
xnor U1107 (N_1107,N_686,N_514);
and U1108 (N_1108,N_654,N_715);
or U1109 (N_1109,N_713,N_617);
or U1110 (N_1110,N_849,N_687);
or U1111 (N_1111,N_798,N_536);
nand U1112 (N_1112,N_976,N_807);
and U1113 (N_1113,N_873,N_870);
nor U1114 (N_1114,N_690,N_943);
xor U1115 (N_1115,N_589,N_565);
nor U1116 (N_1116,N_567,N_945);
nor U1117 (N_1117,N_615,N_834);
nand U1118 (N_1118,N_925,N_929);
nand U1119 (N_1119,N_912,N_532);
xnor U1120 (N_1120,N_825,N_533);
nor U1121 (N_1121,N_755,N_663);
or U1122 (N_1122,N_752,N_778);
xnor U1123 (N_1123,N_821,N_916);
nor U1124 (N_1124,N_858,N_632);
and U1125 (N_1125,N_843,N_792);
xor U1126 (N_1126,N_776,N_723);
or U1127 (N_1127,N_744,N_804);
or U1128 (N_1128,N_939,N_962);
nor U1129 (N_1129,N_657,N_634);
xor U1130 (N_1130,N_709,N_888);
and U1131 (N_1131,N_908,N_872);
and U1132 (N_1132,N_836,N_601);
nand U1133 (N_1133,N_529,N_862);
nand U1134 (N_1134,N_838,N_585);
nor U1135 (N_1135,N_522,N_684);
nand U1136 (N_1136,N_681,N_641);
and U1137 (N_1137,N_694,N_673);
or U1138 (N_1138,N_799,N_587);
or U1139 (N_1139,N_559,N_796);
or U1140 (N_1140,N_638,N_751);
nor U1141 (N_1141,N_571,N_535);
or U1142 (N_1142,N_586,N_552);
nand U1143 (N_1143,N_879,N_750);
and U1144 (N_1144,N_846,N_525);
and U1145 (N_1145,N_693,N_629);
or U1146 (N_1146,N_917,N_878);
xnor U1147 (N_1147,N_899,N_692);
or U1148 (N_1148,N_835,N_894);
xnor U1149 (N_1149,N_761,N_630);
nand U1150 (N_1150,N_695,N_782);
and U1151 (N_1151,N_770,N_594);
xor U1152 (N_1152,N_523,N_604);
nand U1153 (N_1153,N_775,N_978);
and U1154 (N_1154,N_763,N_944);
xor U1155 (N_1155,N_653,N_850);
or U1156 (N_1156,N_774,N_859);
xor U1157 (N_1157,N_813,N_647);
and U1158 (N_1158,N_720,N_549);
xnor U1159 (N_1159,N_815,N_737);
nor U1160 (N_1160,N_509,N_700);
nor U1161 (N_1161,N_810,N_716);
nor U1162 (N_1162,N_904,N_581);
or U1163 (N_1163,N_952,N_971);
nand U1164 (N_1164,N_650,N_997);
and U1165 (N_1165,N_550,N_636);
nor U1166 (N_1166,N_797,N_521);
nand U1167 (N_1167,N_790,N_893);
xnor U1168 (N_1168,N_676,N_665);
or U1169 (N_1169,N_833,N_616);
nand U1170 (N_1170,N_793,N_805);
or U1171 (N_1171,N_696,N_674);
nand U1172 (N_1172,N_830,N_667);
and U1173 (N_1173,N_785,N_932);
nand U1174 (N_1174,N_547,N_655);
or U1175 (N_1175,N_900,N_545);
nor U1176 (N_1176,N_784,N_608);
xor U1177 (N_1177,N_606,N_998);
xnor U1178 (N_1178,N_592,N_555);
nor U1179 (N_1179,N_841,N_526);
and U1180 (N_1180,N_599,N_953);
xor U1181 (N_1181,N_660,N_611);
xor U1182 (N_1182,N_621,N_949);
nor U1183 (N_1183,N_683,N_671);
or U1184 (N_1184,N_627,N_876);
or U1185 (N_1185,N_659,N_980);
or U1186 (N_1186,N_666,N_578);
nand U1187 (N_1187,N_884,N_564);
and U1188 (N_1188,N_739,N_652);
and U1189 (N_1189,N_948,N_517);
nor U1190 (N_1190,N_607,N_809);
or U1191 (N_1191,N_612,N_702);
or U1192 (N_1192,N_856,N_538);
xnor U1193 (N_1193,N_965,N_839);
or U1194 (N_1194,N_934,N_685);
and U1195 (N_1195,N_512,N_787);
nand U1196 (N_1196,N_814,N_537);
xor U1197 (N_1197,N_765,N_983);
or U1198 (N_1198,N_902,N_915);
xnor U1199 (N_1199,N_766,N_842);
or U1200 (N_1200,N_816,N_963);
or U1201 (N_1201,N_588,N_756);
xnor U1202 (N_1202,N_563,N_972);
nand U1203 (N_1203,N_975,N_623);
nor U1204 (N_1204,N_712,N_957);
nor U1205 (N_1205,N_644,N_753);
and U1206 (N_1206,N_635,N_946);
and U1207 (N_1207,N_920,N_738);
or U1208 (N_1208,N_780,N_860);
or U1209 (N_1209,N_729,N_935);
nor U1210 (N_1210,N_602,N_954);
nand U1211 (N_1211,N_732,N_772);
and U1212 (N_1212,N_609,N_880);
or U1213 (N_1213,N_937,N_743);
nor U1214 (N_1214,N_572,N_579);
or U1215 (N_1215,N_524,N_628);
nor U1216 (N_1216,N_824,N_847);
nor U1217 (N_1217,N_973,N_885);
and U1218 (N_1218,N_527,N_869);
and U1219 (N_1219,N_727,N_736);
nand U1220 (N_1220,N_827,N_705);
nor U1221 (N_1221,N_828,N_947);
nand U1222 (N_1222,N_795,N_951);
nor U1223 (N_1223,N_697,N_670);
nor U1224 (N_1224,N_837,N_861);
nor U1225 (N_1225,N_648,N_583);
xor U1226 (N_1226,N_710,N_922);
and U1227 (N_1227,N_701,N_906);
and U1228 (N_1228,N_852,N_868);
and U1229 (N_1229,N_625,N_936);
or U1230 (N_1230,N_783,N_561);
xor U1231 (N_1231,N_927,N_993);
nand U1232 (N_1232,N_820,N_956);
nor U1233 (N_1233,N_961,N_637);
nand U1234 (N_1234,N_724,N_733);
or U1235 (N_1235,N_544,N_622);
and U1236 (N_1236,N_539,N_534);
nand U1237 (N_1237,N_631,N_999);
or U1238 (N_1238,N_591,N_614);
nand U1239 (N_1239,N_762,N_558);
nor U1240 (N_1240,N_613,N_658);
or U1241 (N_1241,N_605,N_817);
or U1242 (N_1242,N_725,N_680);
and U1243 (N_1243,N_991,N_950);
nor U1244 (N_1244,N_516,N_988);
nor U1245 (N_1245,N_682,N_905);
nand U1246 (N_1246,N_891,N_990);
nor U1247 (N_1247,N_722,N_679);
and U1248 (N_1248,N_811,N_773);
nor U1249 (N_1249,N_882,N_669);
xnor U1250 (N_1250,N_889,N_723);
and U1251 (N_1251,N_818,N_714);
nand U1252 (N_1252,N_852,N_713);
xnor U1253 (N_1253,N_868,N_773);
nand U1254 (N_1254,N_952,N_510);
nor U1255 (N_1255,N_530,N_728);
nand U1256 (N_1256,N_737,N_862);
nor U1257 (N_1257,N_957,N_544);
nand U1258 (N_1258,N_946,N_659);
and U1259 (N_1259,N_605,N_965);
xnor U1260 (N_1260,N_618,N_709);
nand U1261 (N_1261,N_580,N_641);
xor U1262 (N_1262,N_722,N_885);
or U1263 (N_1263,N_714,N_979);
or U1264 (N_1264,N_743,N_875);
nor U1265 (N_1265,N_970,N_731);
or U1266 (N_1266,N_709,N_528);
nand U1267 (N_1267,N_870,N_625);
and U1268 (N_1268,N_897,N_713);
or U1269 (N_1269,N_525,N_609);
nor U1270 (N_1270,N_854,N_772);
xor U1271 (N_1271,N_797,N_896);
and U1272 (N_1272,N_688,N_867);
xnor U1273 (N_1273,N_621,N_905);
xor U1274 (N_1274,N_607,N_765);
nand U1275 (N_1275,N_923,N_526);
or U1276 (N_1276,N_693,N_574);
or U1277 (N_1277,N_910,N_975);
nor U1278 (N_1278,N_717,N_790);
xor U1279 (N_1279,N_746,N_872);
xor U1280 (N_1280,N_820,N_746);
or U1281 (N_1281,N_642,N_695);
and U1282 (N_1282,N_550,N_818);
xor U1283 (N_1283,N_774,N_730);
or U1284 (N_1284,N_601,N_946);
xor U1285 (N_1285,N_612,N_801);
and U1286 (N_1286,N_948,N_899);
or U1287 (N_1287,N_564,N_630);
or U1288 (N_1288,N_572,N_514);
xnor U1289 (N_1289,N_726,N_941);
or U1290 (N_1290,N_811,N_626);
and U1291 (N_1291,N_528,N_806);
nand U1292 (N_1292,N_790,N_829);
nor U1293 (N_1293,N_579,N_872);
or U1294 (N_1294,N_961,N_657);
nor U1295 (N_1295,N_940,N_599);
and U1296 (N_1296,N_876,N_873);
xnor U1297 (N_1297,N_590,N_815);
or U1298 (N_1298,N_710,N_876);
nor U1299 (N_1299,N_996,N_807);
or U1300 (N_1300,N_991,N_647);
xor U1301 (N_1301,N_637,N_823);
xor U1302 (N_1302,N_701,N_531);
nand U1303 (N_1303,N_606,N_841);
or U1304 (N_1304,N_539,N_560);
nor U1305 (N_1305,N_899,N_944);
or U1306 (N_1306,N_690,N_894);
and U1307 (N_1307,N_814,N_969);
nand U1308 (N_1308,N_976,N_500);
nand U1309 (N_1309,N_616,N_677);
nor U1310 (N_1310,N_898,N_863);
nand U1311 (N_1311,N_882,N_887);
or U1312 (N_1312,N_585,N_641);
and U1313 (N_1313,N_548,N_803);
xor U1314 (N_1314,N_763,N_989);
xor U1315 (N_1315,N_767,N_842);
xor U1316 (N_1316,N_527,N_717);
and U1317 (N_1317,N_862,N_621);
and U1318 (N_1318,N_874,N_917);
nor U1319 (N_1319,N_942,N_583);
nor U1320 (N_1320,N_679,N_976);
nand U1321 (N_1321,N_770,N_817);
or U1322 (N_1322,N_917,N_643);
and U1323 (N_1323,N_894,N_642);
nand U1324 (N_1324,N_503,N_501);
xor U1325 (N_1325,N_870,N_877);
or U1326 (N_1326,N_964,N_642);
nand U1327 (N_1327,N_691,N_873);
or U1328 (N_1328,N_572,N_995);
and U1329 (N_1329,N_801,N_670);
or U1330 (N_1330,N_693,N_972);
or U1331 (N_1331,N_999,N_741);
and U1332 (N_1332,N_976,N_998);
or U1333 (N_1333,N_547,N_663);
xor U1334 (N_1334,N_685,N_913);
xnor U1335 (N_1335,N_730,N_821);
and U1336 (N_1336,N_991,N_727);
nand U1337 (N_1337,N_767,N_530);
or U1338 (N_1338,N_524,N_698);
and U1339 (N_1339,N_701,N_725);
xnor U1340 (N_1340,N_629,N_969);
or U1341 (N_1341,N_766,N_660);
xor U1342 (N_1342,N_995,N_903);
xor U1343 (N_1343,N_789,N_943);
and U1344 (N_1344,N_917,N_709);
and U1345 (N_1345,N_858,N_682);
xor U1346 (N_1346,N_510,N_991);
and U1347 (N_1347,N_905,N_743);
or U1348 (N_1348,N_512,N_748);
and U1349 (N_1349,N_757,N_923);
nand U1350 (N_1350,N_757,N_716);
xnor U1351 (N_1351,N_712,N_576);
nand U1352 (N_1352,N_750,N_818);
xnor U1353 (N_1353,N_888,N_521);
or U1354 (N_1354,N_850,N_664);
and U1355 (N_1355,N_547,N_549);
nor U1356 (N_1356,N_871,N_749);
or U1357 (N_1357,N_851,N_995);
nand U1358 (N_1358,N_860,N_977);
xnor U1359 (N_1359,N_963,N_577);
nand U1360 (N_1360,N_826,N_867);
nor U1361 (N_1361,N_958,N_827);
nor U1362 (N_1362,N_552,N_644);
and U1363 (N_1363,N_926,N_665);
and U1364 (N_1364,N_612,N_934);
or U1365 (N_1365,N_561,N_860);
nand U1366 (N_1366,N_584,N_708);
and U1367 (N_1367,N_642,N_533);
nand U1368 (N_1368,N_655,N_513);
xor U1369 (N_1369,N_890,N_900);
nor U1370 (N_1370,N_773,N_961);
and U1371 (N_1371,N_963,N_871);
or U1372 (N_1372,N_803,N_676);
nand U1373 (N_1373,N_743,N_956);
nor U1374 (N_1374,N_731,N_579);
nor U1375 (N_1375,N_979,N_552);
xnor U1376 (N_1376,N_967,N_940);
or U1377 (N_1377,N_547,N_720);
or U1378 (N_1378,N_816,N_668);
nand U1379 (N_1379,N_512,N_676);
xor U1380 (N_1380,N_514,N_509);
xor U1381 (N_1381,N_880,N_968);
xor U1382 (N_1382,N_789,N_862);
and U1383 (N_1383,N_867,N_765);
and U1384 (N_1384,N_500,N_515);
xor U1385 (N_1385,N_812,N_586);
xnor U1386 (N_1386,N_794,N_535);
and U1387 (N_1387,N_596,N_558);
and U1388 (N_1388,N_727,N_874);
nand U1389 (N_1389,N_511,N_695);
or U1390 (N_1390,N_655,N_935);
nand U1391 (N_1391,N_900,N_806);
nand U1392 (N_1392,N_696,N_663);
nand U1393 (N_1393,N_884,N_630);
nand U1394 (N_1394,N_772,N_880);
xnor U1395 (N_1395,N_888,N_764);
or U1396 (N_1396,N_807,N_825);
or U1397 (N_1397,N_563,N_528);
or U1398 (N_1398,N_776,N_844);
nand U1399 (N_1399,N_771,N_757);
and U1400 (N_1400,N_854,N_601);
and U1401 (N_1401,N_552,N_990);
or U1402 (N_1402,N_817,N_523);
nand U1403 (N_1403,N_853,N_889);
and U1404 (N_1404,N_754,N_824);
nand U1405 (N_1405,N_664,N_876);
nand U1406 (N_1406,N_597,N_592);
nand U1407 (N_1407,N_791,N_689);
and U1408 (N_1408,N_595,N_712);
and U1409 (N_1409,N_547,N_932);
nor U1410 (N_1410,N_665,N_862);
nor U1411 (N_1411,N_961,N_558);
nand U1412 (N_1412,N_953,N_534);
nor U1413 (N_1413,N_732,N_852);
and U1414 (N_1414,N_545,N_952);
nand U1415 (N_1415,N_689,N_857);
nand U1416 (N_1416,N_914,N_984);
and U1417 (N_1417,N_507,N_613);
nand U1418 (N_1418,N_977,N_982);
nand U1419 (N_1419,N_646,N_585);
nor U1420 (N_1420,N_998,N_599);
and U1421 (N_1421,N_738,N_771);
xnor U1422 (N_1422,N_558,N_921);
or U1423 (N_1423,N_621,N_648);
and U1424 (N_1424,N_980,N_614);
nand U1425 (N_1425,N_969,N_684);
xor U1426 (N_1426,N_825,N_811);
nor U1427 (N_1427,N_890,N_821);
xnor U1428 (N_1428,N_819,N_637);
xnor U1429 (N_1429,N_894,N_787);
nor U1430 (N_1430,N_512,N_672);
and U1431 (N_1431,N_673,N_647);
and U1432 (N_1432,N_531,N_821);
or U1433 (N_1433,N_707,N_594);
and U1434 (N_1434,N_631,N_611);
nor U1435 (N_1435,N_948,N_957);
and U1436 (N_1436,N_920,N_845);
and U1437 (N_1437,N_890,N_953);
or U1438 (N_1438,N_594,N_536);
xor U1439 (N_1439,N_947,N_706);
xor U1440 (N_1440,N_950,N_693);
xor U1441 (N_1441,N_654,N_864);
nand U1442 (N_1442,N_964,N_680);
and U1443 (N_1443,N_502,N_538);
and U1444 (N_1444,N_838,N_575);
and U1445 (N_1445,N_929,N_999);
and U1446 (N_1446,N_645,N_618);
nand U1447 (N_1447,N_847,N_762);
nand U1448 (N_1448,N_969,N_789);
or U1449 (N_1449,N_876,N_595);
or U1450 (N_1450,N_999,N_693);
and U1451 (N_1451,N_750,N_741);
or U1452 (N_1452,N_896,N_927);
nand U1453 (N_1453,N_506,N_941);
xor U1454 (N_1454,N_574,N_867);
or U1455 (N_1455,N_734,N_761);
nor U1456 (N_1456,N_974,N_823);
nand U1457 (N_1457,N_902,N_563);
and U1458 (N_1458,N_792,N_651);
xor U1459 (N_1459,N_718,N_852);
xor U1460 (N_1460,N_572,N_694);
nor U1461 (N_1461,N_890,N_993);
or U1462 (N_1462,N_866,N_732);
nor U1463 (N_1463,N_928,N_622);
or U1464 (N_1464,N_730,N_825);
xor U1465 (N_1465,N_869,N_804);
or U1466 (N_1466,N_832,N_513);
nand U1467 (N_1467,N_502,N_954);
and U1468 (N_1468,N_717,N_740);
nand U1469 (N_1469,N_870,N_704);
and U1470 (N_1470,N_708,N_970);
and U1471 (N_1471,N_600,N_555);
and U1472 (N_1472,N_552,N_825);
or U1473 (N_1473,N_998,N_652);
or U1474 (N_1474,N_615,N_978);
nor U1475 (N_1475,N_643,N_577);
xor U1476 (N_1476,N_591,N_757);
and U1477 (N_1477,N_619,N_977);
or U1478 (N_1478,N_543,N_520);
or U1479 (N_1479,N_723,N_970);
and U1480 (N_1480,N_867,N_968);
or U1481 (N_1481,N_694,N_949);
or U1482 (N_1482,N_654,N_614);
nand U1483 (N_1483,N_628,N_668);
or U1484 (N_1484,N_519,N_569);
nand U1485 (N_1485,N_914,N_523);
xor U1486 (N_1486,N_537,N_729);
xor U1487 (N_1487,N_650,N_824);
xor U1488 (N_1488,N_958,N_768);
and U1489 (N_1489,N_665,N_577);
nor U1490 (N_1490,N_673,N_893);
nor U1491 (N_1491,N_981,N_663);
nand U1492 (N_1492,N_680,N_800);
or U1493 (N_1493,N_820,N_730);
nor U1494 (N_1494,N_583,N_831);
nor U1495 (N_1495,N_989,N_708);
and U1496 (N_1496,N_643,N_880);
and U1497 (N_1497,N_759,N_608);
xnor U1498 (N_1498,N_936,N_864);
xor U1499 (N_1499,N_570,N_531);
or U1500 (N_1500,N_1324,N_1266);
and U1501 (N_1501,N_1203,N_1161);
xnor U1502 (N_1502,N_1498,N_1277);
nand U1503 (N_1503,N_1170,N_1241);
or U1504 (N_1504,N_1361,N_1391);
xor U1505 (N_1505,N_1426,N_1292);
nand U1506 (N_1506,N_1191,N_1349);
nor U1507 (N_1507,N_1477,N_1489);
nor U1508 (N_1508,N_1022,N_1054);
xnor U1509 (N_1509,N_1143,N_1459);
nand U1510 (N_1510,N_1204,N_1081);
nor U1511 (N_1511,N_1468,N_1196);
or U1512 (N_1512,N_1096,N_1184);
nand U1513 (N_1513,N_1497,N_1398);
xnor U1514 (N_1514,N_1418,N_1111);
and U1515 (N_1515,N_1420,N_1106);
xnor U1516 (N_1516,N_1058,N_1469);
xor U1517 (N_1517,N_1004,N_1343);
and U1518 (N_1518,N_1453,N_1013);
and U1519 (N_1519,N_1260,N_1166);
xor U1520 (N_1520,N_1094,N_1271);
nand U1521 (N_1521,N_1034,N_1103);
nor U1522 (N_1522,N_1268,N_1086);
or U1523 (N_1523,N_1128,N_1384);
nor U1524 (N_1524,N_1302,N_1172);
or U1525 (N_1525,N_1217,N_1009);
or U1526 (N_1526,N_1187,N_1028);
or U1527 (N_1527,N_1237,N_1262);
nor U1528 (N_1528,N_1338,N_1140);
nor U1529 (N_1529,N_1139,N_1448);
nor U1530 (N_1530,N_1046,N_1104);
xor U1531 (N_1531,N_1296,N_1330);
nor U1532 (N_1532,N_1311,N_1416);
and U1533 (N_1533,N_1363,N_1099);
xnor U1534 (N_1534,N_1201,N_1449);
or U1535 (N_1535,N_1351,N_1354);
xnor U1536 (N_1536,N_1370,N_1098);
nor U1537 (N_1537,N_1215,N_1220);
and U1538 (N_1538,N_1120,N_1236);
and U1539 (N_1539,N_1347,N_1365);
nor U1540 (N_1540,N_1095,N_1454);
and U1541 (N_1541,N_1157,N_1394);
xnor U1542 (N_1542,N_1216,N_1285);
nand U1543 (N_1543,N_1134,N_1035);
xnor U1544 (N_1544,N_1362,N_1005);
or U1545 (N_1545,N_1344,N_1303);
or U1546 (N_1546,N_1155,N_1006);
xnor U1547 (N_1547,N_1414,N_1171);
xnor U1548 (N_1548,N_1345,N_1425);
xnor U1549 (N_1549,N_1480,N_1256);
and U1550 (N_1550,N_1051,N_1481);
nor U1551 (N_1551,N_1091,N_1210);
xnor U1552 (N_1552,N_1325,N_1373);
and U1553 (N_1553,N_1297,N_1309);
xnor U1554 (N_1554,N_1176,N_1401);
or U1555 (N_1555,N_1301,N_1125);
or U1556 (N_1556,N_1494,N_1224);
xor U1557 (N_1557,N_1214,N_1109);
xnor U1558 (N_1558,N_1113,N_1263);
nor U1559 (N_1559,N_1385,N_1499);
or U1560 (N_1560,N_1386,N_1323);
nor U1561 (N_1561,N_1246,N_1240);
xnor U1562 (N_1562,N_1194,N_1319);
xnor U1563 (N_1563,N_1072,N_1410);
xor U1564 (N_1564,N_1366,N_1195);
nor U1565 (N_1565,N_1088,N_1249);
xor U1566 (N_1566,N_1458,N_1174);
and U1567 (N_1567,N_1002,N_1135);
nand U1568 (N_1568,N_1153,N_1295);
and U1569 (N_1569,N_1375,N_1486);
and U1570 (N_1570,N_1478,N_1069);
or U1571 (N_1571,N_1376,N_1071);
nand U1572 (N_1572,N_1016,N_1346);
nor U1573 (N_1573,N_1193,N_1473);
nor U1574 (N_1574,N_1318,N_1211);
xor U1575 (N_1575,N_1333,N_1177);
xor U1576 (N_1576,N_1082,N_1019);
nor U1577 (N_1577,N_1328,N_1092);
and U1578 (N_1578,N_1165,N_1464);
nand U1579 (N_1579,N_1070,N_1329);
nor U1580 (N_1580,N_1223,N_1250);
or U1581 (N_1581,N_1213,N_1050);
and U1582 (N_1582,N_1352,N_1400);
nor U1583 (N_1583,N_1147,N_1015);
or U1584 (N_1584,N_1131,N_1181);
nand U1585 (N_1585,N_1179,N_1253);
nand U1586 (N_1586,N_1380,N_1484);
nor U1587 (N_1587,N_1463,N_1061);
and U1588 (N_1588,N_1017,N_1432);
xor U1589 (N_1589,N_1118,N_1229);
nand U1590 (N_1590,N_1315,N_1462);
and U1591 (N_1591,N_1159,N_1287);
and U1592 (N_1592,N_1383,N_1014);
nor U1593 (N_1593,N_1496,N_1189);
or U1594 (N_1594,N_1258,N_1310);
xnor U1595 (N_1595,N_1259,N_1062);
nor U1596 (N_1596,N_1100,N_1487);
and U1597 (N_1597,N_1105,N_1030);
and U1598 (N_1598,N_1130,N_1122);
xor U1599 (N_1599,N_1076,N_1348);
xnor U1600 (N_1600,N_1374,N_1322);
nor U1601 (N_1601,N_1276,N_1381);
nor U1602 (N_1602,N_1008,N_1320);
or U1603 (N_1603,N_1492,N_1114);
and U1604 (N_1604,N_1197,N_1337);
or U1605 (N_1605,N_1427,N_1447);
and U1606 (N_1606,N_1340,N_1443);
xor U1607 (N_1607,N_1235,N_1412);
nor U1608 (N_1608,N_1080,N_1470);
nor U1609 (N_1609,N_1031,N_1411);
or U1610 (N_1610,N_1299,N_1047);
nand U1611 (N_1611,N_1326,N_1012);
nor U1612 (N_1612,N_1436,N_1112);
and U1613 (N_1613,N_1342,N_1387);
and U1614 (N_1614,N_1180,N_1475);
nand U1615 (N_1615,N_1026,N_1424);
nor U1616 (N_1616,N_1435,N_1298);
and U1617 (N_1617,N_1368,N_1254);
nor U1618 (N_1618,N_1377,N_1207);
xnor U1619 (N_1619,N_1097,N_1212);
and U1620 (N_1620,N_1300,N_1045);
nor U1621 (N_1621,N_1488,N_1456);
xnor U1622 (N_1622,N_1457,N_1409);
xnor U1623 (N_1623,N_1089,N_1378);
and U1624 (N_1624,N_1123,N_1465);
or U1625 (N_1625,N_1186,N_1145);
nand U1626 (N_1626,N_1075,N_1244);
and U1627 (N_1627,N_1039,N_1020);
nand U1628 (N_1628,N_1442,N_1222);
nor U1629 (N_1629,N_1495,N_1079);
xor U1630 (N_1630,N_1049,N_1126);
nor U1631 (N_1631,N_1024,N_1293);
and U1632 (N_1632,N_1044,N_1067);
and U1633 (N_1633,N_1066,N_1138);
xnor U1634 (N_1634,N_1090,N_1068);
xnor U1635 (N_1635,N_1415,N_1150);
nor U1636 (N_1636,N_1036,N_1392);
and U1637 (N_1637,N_1291,N_1431);
or U1638 (N_1638,N_1048,N_1451);
xnor U1639 (N_1639,N_1227,N_1200);
nor U1640 (N_1640,N_1304,N_1314);
or U1641 (N_1641,N_1274,N_1121);
and U1642 (N_1642,N_1476,N_1367);
nor U1643 (N_1643,N_1085,N_1479);
nand U1644 (N_1644,N_1078,N_1230);
and U1645 (N_1645,N_1158,N_1202);
xor U1646 (N_1646,N_1167,N_1225);
nor U1647 (N_1647,N_1149,N_1183);
or U1648 (N_1648,N_1001,N_1219);
xnor U1649 (N_1649,N_1077,N_1041);
xor U1650 (N_1650,N_1434,N_1269);
xnor U1651 (N_1651,N_1185,N_1429);
nor U1652 (N_1652,N_1057,N_1289);
nand U1653 (N_1653,N_1467,N_1408);
nand U1654 (N_1654,N_1152,N_1360);
nand U1655 (N_1655,N_1007,N_1341);
nor U1656 (N_1656,N_1242,N_1209);
and U1657 (N_1657,N_1188,N_1421);
nor U1658 (N_1658,N_1038,N_1115);
nand U1659 (N_1659,N_1052,N_1164);
nor U1660 (N_1660,N_1327,N_1198);
and U1661 (N_1661,N_1192,N_1011);
or U1662 (N_1662,N_1221,N_1405);
xnor U1663 (N_1663,N_1154,N_1107);
nand U1664 (N_1664,N_1472,N_1388);
xor U1665 (N_1665,N_1029,N_1175);
nor U1666 (N_1666,N_1316,N_1151);
xnor U1667 (N_1667,N_1313,N_1422);
or U1668 (N_1668,N_1390,N_1393);
nor U1669 (N_1669,N_1438,N_1372);
nor U1670 (N_1670,N_1137,N_1321);
nand U1671 (N_1671,N_1406,N_1402);
and U1672 (N_1672,N_1307,N_1132);
or U1673 (N_1673,N_1364,N_1334);
xnor U1674 (N_1674,N_1440,N_1124);
and U1675 (N_1675,N_1226,N_1455);
nand U1676 (N_1676,N_1471,N_1141);
nand U1677 (N_1677,N_1437,N_1033);
nand U1678 (N_1678,N_1018,N_1043);
xnor U1679 (N_1679,N_1460,N_1073);
nor U1680 (N_1680,N_1119,N_1208);
nand U1681 (N_1681,N_1397,N_1248);
and U1682 (N_1682,N_1199,N_1239);
nand U1683 (N_1683,N_1445,N_1403);
nand U1684 (N_1684,N_1282,N_1084);
nor U1685 (N_1685,N_1371,N_1419);
or U1686 (N_1686,N_1055,N_1074);
and U1687 (N_1687,N_1452,N_1450);
nand U1688 (N_1688,N_1466,N_1116);
nor U1689 (N_1689,N_1108,N_1228);
xnor U1690 (N_1690,N_1257,N_1286);
and U1691 (N_1691,N_1059,N_1238);
nor U1692 (N_1692,N_1025,N_1396);
or U1693 (N_1693,N_1283,N_1182);
xor U1694 (N_1694,N_1023,N_1336);
nor U1695 (N_1695,N_1133,N_1101);
or U1696 (N_1696,N_1413,N_1358);
or U1697 (N_1697,N_1275,N_1483);
nand U1698 (N_1698,N_1474,N_1003);
nand U1699 (N_1699,N_1273,N_1169);
nor U1700 (N_1700,N_1261,N_1163);
xnor U1701 (N_1701,N_1110,N_1064);
nand U1702 (N_1702,N_1129,N_1162);
xnor U1703 (N_1703,N_1399,N_1308);
nor U1704 (N_1704,N_1270,N_1335);
nor U1705 (N_1705,N_1021,N_1395);
and U1706 (N_1706,N_1190,N_1279);
nand U1707 (N_1707,N_1231,N_1357);
nor U1708 (N_1708,N_1444,N_1280);
and U1709 (N_1709,N_1247,N_1117);
or U1710 (N_1710,N_1265,N_1491);
and U1711 (N_1711,N_1032,N_1355);
nor U1712 (N_1712,N_1056,N_1146);
or U1713 (N_1713,N_1305,N_1000);
and U1714 (N_1714,N_1234,N_1037);
nand U1715 (N_1715,N_1332,N_1168);
nand U1716 (N_1716,N_1290,N_1306);
nand U1717 (N_1717,N_1205,N_1433);
nor U1718 (N_1718,N_1040,N_1312);
or U1719 (N_1719,N_1233,N_1339);
xnor U1720 (N_1720,N_1379,N_1353);
and U1721 (N_1721,N_1417,N_1356);
nor U1722 (N_1722,N_1156,N_1430);
nor U1723 (N_1723,N_1493,N_1252);
xor U1724 (N_1724,N_1218,N_1243);
nor U1725 (N_1725,N_1127,N_1102);
xor U1726 (N_1726,N_1428,N_1294);
and U1727 (N_1727,N_1087,N_1482);
xnor U1728 (N_1728,N_1053,N_1160);
or U1729 (N_1729,N_1173,N_1264);
xnor U1730 (N_1730,N_1423,N_1232);
nor U1731 (N_1731,N_1317,N_1439);
xnor U1732 (N_1732,N_1083,N_1148);
nand U1733 (N_1733,N_1245,N_1404);
nand U1734 (N_1734,N_1027,N_1490);
nand U1735 (N_1735,N_1093,N_1255);
or U1736 (N_1736,N_1382,N_1136);
nor U1737 (N_1737,N_1281,N_1389);
nand U1738 (N_1738,N_1272,N_1407);
and U1739 (N_1739,N_1441,N_1331);
nor U1740 (N_1740,N_1060,N_1284);
or U1741 (N_1741,N_1010,N_1350);
or U1742 (N_1742,N_1278,N_1359);
nor U1743 (N_1743,N_1288,N_1142);
nand U1744 (N_1744,N_1063,N_1178);
or U1745 (N_1745,N_1042,N_1206);
nor U1746 (N_1746,N_1144,N_1251);
nand U1747 (N_1747,N_1065,N_1369);
or U1748 (N_1748,N_1446,N_1267);
or U1749 (N_1749,N_1461,N_1485);
nor U1750 (N_1750,N_1465,N_1195);
or U1751 (N_1751,N_1240,N_1150);
nand U1752 (N_1752,N_1388,N_1176);
nor U1753 (N_1753,N_1080,N_1221);
and U1754 (N_1754,N_1277,N_1077);
xnor U1755 (N_1755,N_1290,N_1217);
nor U1756 (N_1756,N_1443,N_1084);
nor U1757 (N_1757,N_1348,N_1340);
nand U1758 (N_1758,N_1282,N_1305);
nor U1759 (N_1759,N_1156,N_1161);
nand U1760 (N_1760,N_1089,N_1159);
xor U1761 (N_1761,N_1420,N_1067);
nand U1762 (N_1762,N_1359,N_1226);
xor U1763 (N_1763,N_1443,N_1280);
or U1764 (N_1764,N_1307,N_1170);
nand U1765 (N_1765,N_1456,N_1218);
nor U1766 (N_1766,N_1496,N_1053);
and U1767 (N_1767,N_1269,N_1250);
xor U1768 (N_1768,N_1024,N_1260);
nand U1769 (N_1769,N_1163,N_1206);
nand U1770 (N_1770,N_1312,N_1454);
and U1771 (N_1771,N_1127,N_1189);
nand U1772 (N_1772,N_1353,N_1198);
or U1773 (N_1773,N_1399,N_1009);
and U1774 (N_1774,N_1355,N_1287);
and U1775 (N_1775,N_1097,N_1073);
nor U1776 (N_1776,N_1358,N_1135);
nor U1777 (N_1777,N_1198,N_1047);
nor U1778 (N_1778,N_1424,N_1478);
nand U1779 (N_1779,N_1081,N_1428);
and U1780 (N_1780,N_1458,N_1315);
or U1781 (N_1781,N_1282,N_1227);
xor U1782 (N_1782,N_1367,N_1234);
and U1783 (N_1783,N_1056,N_1414);
xor U1784 (N_1784,N_1195,N_1367);
nand U1785 (N_1785,N_1457,N_1151);
or U1786 (N_1786,N_1260,N_1265);
or U1787 (N_1787,N_1084,N_1216);
and U1788 (N_1788,N_1005,N_1326);
nor U1789 (N_1789,N_1234,N_1358);
and U1790 (N_1790,N_1466,N_1407);
or U1791 (N_1791,N_1391,N_1332);
nor U1792 (N_1792,N_1241,N_1060);
nor U1793 (N_1793,N_1418,N_1252);
xnor U1794 (N_1794,N_1093,N_1415);
and U1795 (N_1795,N_1398,N_1366);
nand U1796 (N_1796,N_1124,N_1156);
nand U1797 (N_1797,N_1058,N_1308);
nand U1798 (N_1798,N_1190,N_1480);
xnor U1799 (N_1799,N_1478,N_1303);
nand U1800 (N_1800,N_1382,N_1090);
nand U1801 (N_1801,N_1317,N_1363);
xnor U1802 (N_1802,N_1308,N_1295);
and U1803 (N_1803,N_1100,N_1291);
xor U1804 (N_1804,N_1384,N_1428);
and U1805 (N_1805,N_1423,N_1445);
xnor U1806 (N_1806,N_1440,N_1167);
nor U1807 (N_1807,N_1054,N_1048);
and U1808 (N_1808,N_1080,N_1396);
and U1809 (N_1809,N_1147,N_1138);
and U1810 (N_1810,N_1436,N_1450);
nor U1811 (N_1811,N_1041,N_1150);
nand U1812 (N_1812,N_1191,N_1092);
and U1813 (N_1813,N_1207,N_1114);
nor U1814 (N_1814,N_1360,N_1105);
nand U1815 (N_1815,N_1006,N_1316);
or U1816 (N_1816,N_1454,N_1211);
nand U1817 (N_1817,N_1302,N_1213);
nand U1818 (N_1818,N_1357,N_1110);
xor U1819 (N_1819,N_1146,N_1314);
and U1820 (N_1820,N_1051,N_1277);
and U1821 (N_1821,N_1080,N_1190);
or U1822 (N_1822,N_1072,N_1149);
and U1823 (N_1823,N_1422,N_1477);
and U1824 (N_1824,N_1401,N_1112);
and U1825 (N_1825,N_1022,N_1152);
xor U1826 (N_1826,N_1437,N_1114);
and U1827 (N_1827,N_1456,N_1330);
or U1828 (N_1828,N_1066,N_1083);
and U1829 (N_1829,N_1423,N_1275);
and U1830 (N_1830,N_1336,N_1112);
and U1831 (N_1831,N_1140,N_1485);
or U1832 (N_1832,N_1071,N_1206);
nand U1833 (N_1833,N_1156,N_1262);
or U1834 (N_1834,N_1081,N_1020);
nor U1835 (N_1835,N_1410,N_1446);
nand U1836 (N_1836,N_1027,N_1138);
or U1837 (N_1837,N_1247,N_1195);
xnor U1838 (N_1838,N_1251,N_1485);
or U1839 (N_1839,N_1399,N_1018);
xor U1840 (N_1840,N_1152,N_1431);
xor U1841 (N_1841,N_1030,N_1357);
nor U1842 (N_1842,N_1350,N_1224);
nand U1843 (N_1843,N_1376,N_1235);
xor U1844 (N_1844,N_1429,N_1084);
and U1845 (N_1845,N_1180,N_1304);
and U1846 (N_1846,N_1345,N_1214);
and U1847 (N_1847,N_1475,N_1285);
nand U1848 (N_1848,N_1209,N_1361);
nand U1849 (N_1849,N_1233,N_1196);
nor U1850 (N_1850,N_1448,N_1056);
nor U1851 (N_1851,N_1126,N_1245);
or U1852 (N_1852,N_1127,N_1125);
nand U1853 (N_1853,N_1183,N_1441);
xor U1854 (N_1854,N_1129,N_1173);
nor U1855 (N_1855,N_1418,N_1488);
and U1856 (N_1856,N_1045,N_1119);
nor U1857 (N_1857,N_1285,N_1027);
and U1858 (N_1858,N_1435,N_1160);
nor U1859 (N_1859,N_1074,N_1318);
and U1860 (N_1860,N_1313,N_1245);
nand U1861 (N_1861,N_1323,N_1302);
and U1862 (N_1862,N_1006,N_1116);
or U1863 (N_1863,N_1151,N_1336);
nor U1864 (N_1864,N_1310,N_1154);
nand U1865 (N_1865,N_1409,N_1400);
nand U1866 (N_1866,N_1459,N_1170);
or U1867 (N_1867,N_1207,N_1250);
or U1868 (N_1868,N_1018,N_1223);
or U1869 (N_1869,N_1309,N_1494);
nand U1870 (N_1870,N_1486,N_1438);
nor U1871 (N_1871,N_1492,N_1428);
or U1872 (N_1872,N_1430,N_1169);
nor U1873 (N_1873,N_1342,N_1487);
and U1874 (N_1874,N_1105,N_1439);
or U1875 (N_1875,N_1291,N_1395);
and U1876 (N_1876,N_1156,N_1201);
nor U1877 (N_1877,N_1361,N_1266);
xnor U1878 (N_1878,N_1211,N_1003);
nor U1879 (N_1879,N_1066,N_1348);
nor U1880 (N_1880,N_1122,N_1075);
nor U1881 (N_1881,N_1076,N_1410);
xor U1882 (N_1882,N_1046,N_1053);
xor U1883 (N_1883,N_1314,N_1119);
nand U1884 (N_1884,N_1230,N_1392);
xnor U1885 (N_1885,N_1324,N_1086);
nand U1886 (N_1886,N_1449,N_1327);
nor U1887 (N_1887,N_1188,N_1130);
or U1888 (N_1888,N_1270,N_1411);
nand U1889 (N_1889,N_1381,N_1424);
xnor U1890 (N_1890,N_1210,N_1439);
xnor U1891 (N_1891,N_1128,N_1241);
or U1892 (N_1892,N_1368,N_1303);
nand U1893 (N_1893,N_1395,N_1421);
and U1894 (N_1894,N_1233,N_1079);
nor U1895 (N_1895,N_1091,N_1044);
and U1896 (N_1896,N_1353,N_1275);
nor U1897 (N_1897,N_1470,N_1300);
or U1898 (N_1898,N_1256,N_1263);
nand U1899 (N_1899,N_1121,N_1068);
and U1900 (N_1900,N_1324,N_1454);
or U1901 (N_1901,N_1462,N_1276);
nor U1902 (N_1902,N_1406,N_1374);
xor U1903 (N_1903,N_1229,N_1049);
and U1904 (N_1904,N_1303,N_1062);
nor U1905 (N_1905,N_1046,N_1477);
xnor U1906 (N_1906,N_1147,N_1421);
or U1907 (N_1907,N_1035,N_1447);
and U1908 (N_1908,N_1189,N_1395);
and U1909 (N_1909,N_1336,N_1070);
and U1910 (N_1910,N_1432,N_1116);
nor U1911 (N_1911,N_1125,N_1024);
nor U1912 (N_1912,N_1176,N_1496);
nand U1913 (N_1913,N_1047,N_1375);
nand U1914 (N_1914,N_1465,N_1499);
and U1915 (N_1915,N_1425,N_1338);
or U1916 (N_1916,N_1258,N_1251);
or U1917 (N_1917,N_1090,N_1339);
xnor U1918 (N_1918,N_1195,N_1280);
or U1919 (N_1919,N_1003,N_1455);
or U1920 (N_1920,N_1360,N_1076);
nand U1921 (N_1921,N_1359,N_1426);
and U1922 (N_1922,N_1447,N_1465);
nand U1923 (N_1923,N_1071,N_1139);
or U1924 (N_1924,N_1270,N_1263);
nand U1925 (N_1925,N_1170,N_1048);
or U1926 (N_1926,N_1291,N_1309);
xnor U1927 (N_1927,N_1268,N_1231);
nand U1928 (N_1928,N_1453,N_1123);
nand U1929 (N_1929,N_1066,N_1449);
nor U1930 (N_1930,N_1393,N_1048);
nand U1931 (N_1931,N_1165,N_1159);
and U1932 (N_1932,N_1490,N_1037);
xnor U1933 (N_1933,N_1178,N_1246);
or U1934 (N_1934,N_1205,N_1174);
and U1935 (N_1935,N_1406,N_1320);
nand U1936 (N_1936,N_1081,N_1353);
nor U1937 (N_1937,N_1444,N_1216);
nand U1938 (N_1938,N_1131,N_1362);
and U1939 (N_1939,N_1122,N_1198);
nand U1940 (N_1940,N_1127,N_1060);
xor U1941 (N_1941,N_1422,N_1226);
and U1942 (N_1942,N_1019,N_1446);
and U1943 (N_1943,N_1324,N_1159);
nor U1944 (N_1944,N_1308,N_1350);
xor U1945 (N_1945,N_1212,N_1241);
or U1946 (N_1946,N_1271,N_1466);
and U1947 (N_1947,N_1224,N_1358);
nor U1948 (N_1948,N_1338,N_1357);
nor U1949 (N_1949,N_1200,N_1488);
nor U1950 (N_1950,N_1393,N_1218);
nor U1951 (N_1951,N_1277,N_1130);
xnor U1952 (N_1952,N_1206,N_1444);
nor U1953 (N_1953,N_1082,N_1306);
xor U1954 (N_1954,N_1495,N_1475);
nor U1955 (N_1955,N_1123,N_1387);
xnor U1956 (N_1956,N_1017,N_1245);
and U1957 (N_1957,N_1291,N_1105);
or U1958 (N_1958,N_1314,N_1130);
and U1959 (N_1959,N_1338,N_1074);
or U1960 (N_1960,N_1040,N_1484);
or U1961 (N_1961,N_1128,N_1460);
nor U1962 (N_1962,N_1421,N_1002);
nor U1963 (N_1963,N_1420,N_1006);
and U1964 (N_1964,N_1440,N_1029);
xor U1965 (N_1965,N_1278,N_1203);
nand U1966 (N_1966,N_1052,N_1233);
and U1967 (N_1967,N_1039,N_1324);
nor U1968 (N_1968,N_1318,N_1416);
xor U1969 (N_1969,N_1369,N_1350);
xnor U1970 (N_1970,N_1445,N_1057);
or U1971 (N_1971,N_1368,N_1186);
and U1972 (N_1972,N_1328,N_1291);
nand U1973 (N_1973,N_1208,N_1400);
nor U1974 (N_1974,N_1143,N_1488);
xor U1975 (N_1975,N_1113,N_1230);
nor U1976 (N_1976,N_1258,N_1275);
nor U1977 (N_1977,N_1042,N_1038);
nand U1978 (N_1978,N_1476,N_1493);
nor U1979 (N_1979,N_1081,N_1142);
or U1980 (N_1980,N_1080,N_1435);
nand U1981 (N_1981,N_1499,N_1255);
nand U1982 (N_1982,N_1388,N_1217);
and U1983 (N_1983,N_1483,N_1242);
nor U1984 (N_1984,N_1133,N_1471);
xnor U1985 (N_1985,N_1347,N_1218);
nor U1986 (N_1986,N_1202,N_1041);
or U1987 (N_1987,N_1073,N_1166);
or U1988 (N_1988,N_1350,N_1071);
xnor U1989 (N_1989,N_1118,N_1441);
nand U1990 (N_1990,N_1395,N_1259);
nand U1991 (N_1991,N_1013,N_1153);
xnor U1992 (N_1992,N_1227,N_1060);
xor U1993 (N_1993,N_1472,N_1049);
xor U1994 (N_1994,N_1016,N_1312);
nor U1995 (N_1995,N_1288,N_1384);
nor U1996 (N_1996,N_1374,N_1261);
xor U1997 (N_1997,N_1162,N_1328);
xnor U1998 (N_1998,N_1029,N_1295);
and U1999 (N_1999,N_1065,N_1295);
nand U2000 (N_2000,N_1934,N_1676);
xnor U2001 (N_2001,N_1620,N_1688);
nand U2002 (N_2002,N_1515,N_1501);
and U2003 (N_2003,N_1885,N_1591);
nand U2004 (N_2004,N_1564,N_1912);
nor U2005 (N_2005,N_1702,N_1971);
or U2006 (N_2006,N_1921,N_1899);
nor U2007 (N_2007,N_1861,N_1744);
or U2008 (N_2008,N_1892,N_1815);
or U2009 (N_2009,N_1710,N_1547);
nor U2010 (N_2010,N_1909,N_1545);
or U2011 (N_2011,N_1713,N_1981);
and U2012 (N_2012,N_1877,N_1649);
xor U2013 (N_2013,N_1886,N_1524);
and U2014 (N_2014,N_1999,N_1667);
xnor U2015 (N_2015,N_1946,N_1603);
xnor U2016 (N_2016,N_1629,N_1799);
or U2017 (N_2017,N_1630,N_1532);
nand U2018 (N_2018,N_1735,N_1889);
nor U2019 (N_2019,N_1561,N_1907);
nor U2020 (N_2020,N_1829,N_1928);
or U2021 (N_2021,N_1992,N_1880);
nand U2022 (N_2022,N_1878,N_1840);
xor U2023 (N_2023,N_1917,N_1527);
nor U2024 (N_2024,N_1626,N_1599);
nor U2025 (N_2025,N_1664,N_1567);
and U2026 (N_2026,N_1665,N_1657);
and U2027 (N_2027,N_1595,N_1882);
xor U2028 (N_2028,N_1782,N_1680);
nand U2029 (N_2029,N_1606,N_1555);
xor U2030 (N_2030,N_1890,N_1640);
nor U2031 (N_2031,N_1835,N_1927);
or U2032 (N_2032,N_1834,N_1951);
and U2033 (N_2033,N_1827,N_1997);
nor U2034 (N_2034,N_1760,N_1633);
and U2035 (N_2035,N_1858,N_1594);
nor U2036 (N_2036,N_1718,N_1612);
and U2037 (N_2037,N_1995,N_1706);
nand U2038 (N_2038,N_1778,N_1813);
and U2039 (N_2039,N_1914,N_1699);
and U2040 (N_2040,N_1530,N_1647);
nor U2041 (N_2041,N_1674,N_1582);
nor U2042 (N_2042,N_1940,N_1911);
or U2043 (N_2043,N_1791,N_1500);
xor U2044 (N_2044,N_1919,N_1560);
and U2045 (N_2045,N_1963,N_1952);
nand U2046 (N_2046,N_1823,N_1937);
and U2047 (N_2047,N_1618,N_1558);
nand U2048 (N_2048,N_1766,N_1846);
and U2049 (N_2049,N_1930,N_1721);
nor U2050 (N_2050,N_1502,N_1762);
or U2051 (N_2051,N_1942,N_1571);
nor U2052 (N_2052,N_1893,N_1659);
xor U2053 (N_2053,N_1522,N_1854);
nand U2054 (N_2054,N_1904,N_1774);
or U2055 (N_2055,N_1731,N_1533);
nor U2056 (N_2056,N_1900,N_1538);
nand U2057 (N_2057,N_1518,N_1549);
nand U2058 (N_2058,N_1679,N_1771);
nor U2059 (N_2059,N_1979,N_1580);
xor U2060 (N_2060,N_1777,N_1964);
and U2061 (N_2061,N_1935,N_1913);
nor U2062 (N_2062,N_1802,N_1637);
xor U2063 (N_2063,N_1988,N_1534);
xor U2064 (N_2064,N_1780,N_1644);
nor U2065 (N_2065,N_1642,N_1586);
or U2066 (N_2066,N_1776,N_1821);
or U2067 (N_2067,N_1974,N_1925);
or U2068 (N_2068,N_1770,N_1800);
xnor U2069 (N_2069,N_1695,N_1609);
nand U2070 (N_2070,N_1652,N_1585);
and U2071 (N_2071,N_1830,N_1587);
or U2072 (N_2072,N_1715,N_1970);
xnor U2073 (N_2073,N_1818,N_1751);
nor U2074 (N_2074,N_1897,N_1619);
and U2075 (N_2075,N_1516,N_1903);
or U2076 (N_2076,N_1906,N_1661);
xor U2077 (N_2077,N_1786,N_1572);
nand U2078 (N_2078,N_1519,N_1749);
nor U2079 (N_2079,N_1566,N_1583);
xnor U2080 (N_2080,N_1576,N_1984);
nor U2081 (N_2081,N_1811,N_1738);
nor U2082 (N_2082,N_1570,N_1809);
xor U2083 (N_2083,N_1923,N_1510);
nand U2084 (N_2084,N_1793,N_1926);
and U2085 (N_2085,N_1717,N_1833);
or U2086 (N_2086,N_1938,N_1593);
and U2087 (N_2087,N_1625,N_1607);
and U2088 (N_2088,N_1883,N_1993);
nor U2089 (N_2089,N_1732,N_1658);
nor U2090 (N_2090,N_1977,N_1853);
nor U2091 (N_2091,N_1588,N_1622);
nand U2092 (N_2092,N_1967,N_1565);
or U2093 (N_2093,N_1969,N_1598);
or U2094 (N_2094,N_1756,N_1753);
xnor U2095 (N_2095,N_1960,N_1908);
xnor U2096 (N_2096,N_1767,N_1961);
and U2097 (N_2097,N_1814,N_1696);
xnor U2098 (N_2098,N_1957,N_1563);
xor U2099 (N_2099,N_1863,N_1704);
and U2100 (N_2100,N_1949,N_1804);
or U2101 (N_2101,N_1725,N_1773);
or U2102 (N_2102,N_1507,N_1632);
nor U2103 (N_2103,N_1962,N_1708);
or U2104 (N_2104,N_1698,N_1876);
or U2105 (N_2105,N_1845,N_1611);
nor U2106 (N_2106,N_1888,N_1546);
nor U2107 (N_2107,N_1922,N_1509);
or U2108 (N_2108,N_1584,N_1551);
xnor U2109 (N_2109,N_1850,N_1645);
or U2110 (N_2110,N_1959,N_1990);
xnor U2111 (N_2111,N_1506,N_1727);
nand U2112 (N_2112,N_1529,N_1866);
nor U2113 (N_2113,N_1678,N_1819);
xnor U2114 (N_2114,N_1839,N_1763);
and U2115 (N_2115,N_1662,N_1740);
xor U2116 (N_2116,N_1837,N_1539);
xor U2117 (N_2117,N_1765,N_1875);
and U2118 (N_2118,N_1536,N_1978);
xnor U2119 (N_2119,N_1722,N_1673);
or U2120 (N_2120,N_1958,N_1779);
and U2121 (N_2121,N_1986,N_1944);
and U2122 (N_2122,N_1671,N_1918);
and U2123 (N_2123,N_1734,N_1691);
nor U2124 (N_2124,N_1998,N_1602);
xnor U2125 (N_2125,N_1807,N_1648);
or U2126 (N_2126,N_1817,N_1634);
and U2127 (N_2127,N_1972,N_1871);
or U2128 (N_2128,N_1505,N_1724);
xnor U2129 (N_2129,N_1552,N_1730);
xnor U2130 (N_2130,N_1719,N_1511);
and U2131 (N_2131,N_1631,N_1508);
nand U2132 (N_2132,N_1864,N_1973);
and U2133 (N_2133,N_1550,N_1989);
nor U2134 (N_2134,N_1808,N_1844);
and U2135 (N_2135,N_1683,N_1675);
and U2136 (N_2136,N_1513,N_1761);
xor U2137 (N_2137,N_1701,N_1945);
nand U2138 (N_2138,N_1672,N_1617);
xor U2139 (N_2139,N_1797,N_1504);
nor U2140 (N_2140,N_1976,N_1816);
nand U2141 (N_2141,N_1700,N_1795);
nor U2142 (N_2142,N_1950,N_1947);
xor U2143 (N_2143,N_1954,N_1653);
and U2144 (N_2144,N_1868,N_1798);
or U2145 (N_2145,N_1703,N_1537);
nand U2146 (N_2146,N_1742,N_1826);
or U2147 (N_2147,N_1788,N_1869);
nand U2148 (N_2148,N_1535,N_1843);
nor U2149 (N_2149,N_1677,N_1574);
or U2150 (N_2150,N_1512,N_1982);
or U2151 (N_2151,N_1881,N_1865);
and U2152 (N_2152,N_1568,N_1980);
nor U2153 (N_2153,N_1628,N_1916);
nor U2154 (N_2154,N_1796,N_1641);
nand U2155 (N_2155,N_1623,N_1711);
or U2156 (N_2156,N_1806,N_1707);
xnor U2157 (N_2157,N_1955,N_1663);
xor U2158 (N_2158,N_1604,N_1745);
nor U2159 (N_2159,N_1832,N_1614);
or U2160 (N_2160,N_1983,N_1852);
and U2161 (N_2161,N_1608,N_1859);
and U2162 (N_2162,N_1781,N_1790);
nand U2163 (N_2163,N_1764,N_1553);
and U2164 (N_2164,N_1772,N_1651);
nand U2165 (N_2165,N_1891,N_1820);
or U2166 (N_2166,N_1579,N_1615);
xor U2167 (N_2167,N_1525,N_1842);
nor U2168 (N_2168,N_1822,N_1660);
xnor U2169 (N_2169,N_1685,N_1867);
nor U2170 (N_2170,N_1924,N_1851);
xor U2171 (N_2171,N_1726,N_1856);
xor U2172 (N_2172,N_1520,N_1785);
nand U2173 (N_2173,N_1920,N_1965);
nor U2174 (N_2174,N_1514,N_1936);
and U2175 (N_2175,N_1953,N_1616);
and U2176 (N_2176,N_1682,N_1884);
nand U2177 (N_2177,N_1787,N_1847);
nand U2178 (N_2178,N_1668,N_1646);
nand U2179 (N_2179,N_1810,N_1639);
nor U2180 (N_2180,N_1728,N_1541);
xnor U2181 (N_2181,N_1932,N_1709);
or U2182 (N_2182,N_1543,N_1716);
nand U2183 (N_2183,N_1592,N_1597);
and U2184 (N_2184,N_1870,N_1939);
or U2185 (N_2185,N_1581,N_1650);
xnor U2186 (N_2186,N_1590,N_1966);
nand U2187 (N_2187,N_1905,N_1759);
or U2188 (N_2188,N_1769,N_1720);
and U2189 (N_2189,N_1933,N_1557);
and U2190 (N_2190,N_1758,N_1948);
xnor U2191 (N_2191,N_1783,N_1895);
xnor U2192 (N_2192,N_1669,N_1638);
xnor U2193 (N_2193,N_1575,N_1741);
nand U2194 (N_2194,N_1824,N_1686);
and U2195 (N_2195,N_1887,N_1526);
and U2196 (N_2196,N_1873,N_1956);
and U2197 (N_2197,N_1693,N_1789);
and U2198 (N_2198,N_1712,N_1898);
nor U2199 (N_2199,N_1714,N_1836);
and U2200 (N_2200,N_1775,N_1987);
nand U2201 (N_2201,N_1621,N_1601);
or U2202 (N_2202,N_1848,N_1812);
nor U2203 (N_2203,N_1748,N_1768);
nor U2204 (N_2204,N_1975,N_1896);
nand U2205 (N_2205,N_1801,N_1872);
nor U2206 (N_2206,N_1792,N_1737);
or U2207 (N_2207,N_1841,N_1754);
nand U2208 (N_2208,N_1692,N_1569);
nor U2209 (N_2209,N_1589,N_1996);
xnor U2210 (N_2210,N_1523,N_1517);
nor U2211 (N_2211,N_1559,N_1862);
nor U2212 (N_2212,N_1666,N_1736);
or U2213 (N_2213,N_1743,N_1855);
nor U2214 (N_2214,N_1528,N_1805);
xor U2215 (N_2215,N_1994,N_1849);
xor U2216 (N_2216,N_1931,N_1687);
or U2217 (N_2217,N_1635,N_1689);
and U2218 (N_2218,N_1542,N_1729);
nand U2219 (N_2219,N_1828,N_1752);
nor U2220 (N_2220,N_1910,N_1985);
nand U2221 (N_2221,N_1562,N_1544);
xor U2222 (N_2222,N_1723,N_1739);
xor U2223 (N_2223,N_1784,N_1627);
and U2224 (N_2224,N_1610,N_1531);
or U2225 (N_2225,N_1578,N_1733);
nor U2226 (N_2226,N_1681,N_1503);
or U2227 (N_2227,N_1605,N_1697);
nor U2228 (N_2228,N_1991,N_1831);
nand U2229 (N_2229,N_1643,N_1613);
and U2230 (N_2230,N_1554,N_1915);
or U2231 (N_2231,N_1577,N_1794);
or U2232 (N_2232,N_1901,N_1902);
and U2233 (N_2233,N_1747,N_1825);
xor U2234 (N_2234,N_1838,N_1750);
and U2235 (N_2235,N_1573,N_1755);
or U2236 (N_2236,N_1670,N_1803);
or U2237 (N_2237,N_1694,N_1757);
and U2238 (N_2238,N_1548,N_1874);
xor U2239 (N_2239,N_1746,N_1894);
nor U2240 (N_2240,N_1879,N_1540);
and U2241 (N_2241,N_1943,N_1521);
nor U2242 (N_2242,N_1929,N_1860);
or U2243 (N_2243,N_1654,N_1556);
xnor U2244 (N_2244,N_1857,N_1684);
nor U2245 (N_2245,N_1705,N_1941);
xnor U2246 (N_2246,N_1596,N_1636);
nand U2247 (N_2247,N_1656,N_1690);
nand U2248 (N_2248,N_1655,N_1624);
or U2249 (N_2249,N_1968,N_1600);
nor U2250 (N_2250,N_1525,N_1855);
and U2251 (N_2251,N_1771,N_1920);
nand U2252 (N_2252,N_1927,N_1868);
xnor U2253 (N_2253,N_1911,N_1556);
nand U2254 (N_2254,N_1779,N_1648);
xor U2255 (N_2255,N_1908,N_1938);
nor U2256 (N_2256,N_1639,N_1772);
and U2257 (N_2257,N_1743,N_1609);
nand U2258 (N_2258,N_1574,N_1543);
or U2259 (N_2259,N_1798,N_1988);
and U2260 (N_2260,N_1684,N_1858);
and U2261 (N_2261,N_1813,N_1816);
and U2262 (N_2262,N_1640,N_1846);
or U2263 (N_2263,N_1516,N_1812);
xnor U2264 (N_2264,N_1957,N_1519);
nand U2265 (N_2265,N_1956,N_1783);
xor U2266 (N_2266,N_1789,N_1858);
xnor U2267 (N_2267,N_1764,N_1531);
or U2268 (N_2268,N_1953,N_1801);
nor U2269 (N_2269,N_1882,N_1872);
and U2270 (N_2270,N_1767,N_1978);
or U2271 (N_2271,N_1758,N_1650);
or U2272 (N_2272,N_1753,N_1992);
or U2273 (N_2273,N_1647,N_1832);
nand U2274 (N_2274,N_1615,N_1774);
nand U2275 (N_2275,N_1582,N_1955);
and U2276 (N_2276,N_1874,N_1515);
xor U2277 (N_2277,N_1532,N_1742);
xnor U2278 (N_2278,N_1941,N_1699);
nor U2279 (N_2279,N_1932,N_1853);
nand U2280 (N_2280,N_1799,N_1598);
and U2281 (N_2281,N_1537,N_1849);
nor U2282 (N_2282,N_1882,N_1605);
and U2283 (N_2283,N_1632,N_1694);
xor U2284 (N_2284,N_1939,N_1900);
nand U2285 (N_2285,N_1702,N_1521);
or U2286 (N_2286,N_1571,N_1601);
or U2287 (N_2287,N_1958,N_1534);
nand U2288 (N_2288,N_1651,N_1715);
nor U2289 (N_2289,N_1545,N_1966);
or U2290 (N_2290,N_1659,N_1792);
or U2291 (N_2291,N_1821,N_1807);
or U2292 (N_2292,N_1852,N_1896);
and U2293 (N_2293,N_1615,N_1505);
nand U2294 (N_2294,N_1521,N_1674);
or U2295 (N_2295,N_1734,N_1921);
nand U2296 (N_2296,N_1869,N_1922);
and U2297 (N_2297,N_1854,N_1785);
or U2298 (N_2298,N_1659,N_1953);
xor U2299 (N_2299,N_1637,N_1905);
or U2300 (N_2300,N_1864,N_1685);
xor U2301 (N_2301,N_1907,N_1847);
nand U2302 (N_2302,N_1940,N_1977);
nand U2303 (N_2303,N_1712,N_1635);
nand U2304 (N_2304,N_1555,N_1954);
xor U2305 (N_2305,N_1555,N_1690);
nand U2306 (N_2306,N_1892,N_1795);
nand U2307 (N_2307,N_1773,N_1619);
xor U2308 (N_2308,N_1744,N_1923);
and U2309 (N_2309,N_1682,N_1800);
and U2310 (N_2310,N_1917,N_1939);
nand U2311 (N_2311,N_1688,N_1856);
nor U2312 (N_2312,N_1948,N_1958);
nor U2313 (N_2313,N_1623,N_1911);
or U2314 (N_2314,N_1948,N_1855);
xor U2315 (N_2315,N_1609,N_1694);
xnor U2316 (N_2316,N_1889,N_1675);
nand U2317 (N_2317,N_1903,N_1718);
nand U2318 (N_2318,N_1712,N_1781);
xor U2319 (N_2319,N_1923,N_1534);
nor U2320 (N_2320,N_1650,N_1948);
or U2321 (N_2321,N_1644,N_1820);
xnor U2322 (N_2322,N_1502,N_1609);
and U2323 (N_2323,N_1800,N_1598);
xnor U2324 (N_2324,N_1914,N_1953);
xnor U2325 (N_2325,N_1642,N_1636);
or U2326 (N_2326,N_1743,N_1748);
and U2327 (N_2327,N_1769,N_1829);
and U2328 (N_2328,N_1911,N_1894);
nand U2329 (N_2329,N_1836,N_1815);
nand U2330 (N_2330,N_1724,N_1780);
nand U2331 (N_2331,N_1994,N_1775);
nand U2332 (N_2332,N_1840,N_1514);
or U2333 (N_2333,N_1507,N_1763);
nand U2334 (N_2334,N_1668,N_1638);
nand U2335 (N_2335,N_1753,N_1740);
and U2336 (N_2336,N_1724,N_1567);
or U2337 (N_2337,N_1669,N_1787);
nand U2338 (N_2338,N_1536,N_1551);
nor U2339 (N_2339,N_1872,N_1835);
or U2340 (N_2340,N_1888,N_1708);
nor U2341 (N_2341,N_1925,N_1642);
nand U2342 (N_2342,N_1766,N_1824);
nor U2343 (N_2343,N_1541,N_1653);
nor U2344 (N_2344,N_1555,N_1697);
and U2345 (N_2345,N_1976,N_1536);
xnor U2346 (N_2346,N_1866,N_1585);
nor U2347 (N_2347,N_1984,N_1655);
nand U2348 (N_2348,N_1790,N_1532);
or U2349 (N_2349,N_1562,N_1819);
xor U2350 (N_2350,N_1518,N_1539);
nor U2351 (N_2351,N_1501,N_1638);
xnor U2352 (N_2352,N_1592,N_1663);
xnor U2353 (N_2353,N_1564,N_1558);
and U2354 (N_2354,N_1588,N_1571);
and U2355 (N_2355,N_1882,N_1838);
and U2356 (N_2356,N_1756,N_1831);
or U2357 (N_2357,N_1670,N_1775);
nor U2358 (N_2358,N_1792,N_1506);
or U2359 (N_2359,N_1698,N_1964);
or U2360 (N_2360,N_1985,N_1561);
xnor U2361 (N_2361,N_1917,N_1697);
xor U2362 (N_2362,N_1615,N_1653);
nand U2363 (N_2363,N_1623,N_1857);
or U2364 (N_2364,N_1905,N_1951);
xnor U2365 (N_2365,N_1519,N_1994);
xnor U2366 (N_2366,N_1990,N_1534);
or U2367 (N_2367,N_1652,N_1683);
xnor U2368 (N_2368,N_1906,N_1642);
or U2369 (N_2369,N_1581,N_1585);
xnor U2370 (N_2370,N_1655,N_1909);
nor U2371 (N_2371,N_1791,N_1540);
nor U2372 (N_2372,N_1664,N_1733);
or U2373 (N_2373,N_1584,N_1741);
and U2374 (N_2374,N_1593,N_1765);
and U2375 (N_2375,N_1746,N_1744);
or U2376 (N_2376,N_1525,N_1858);
nor U2377 (N_2377,N_1626,N_1608);
nand U2378 (N_2378,N_1889,N_1821);
or U2379 (N_2379,N_1922,N_1639);
nor U2380 (N_2380,N_1662,N_1741);
nor U2381 (N_2381,N_1999,N_1950);
xor U2382 (N_2382,N_1898,N_1826);
nand U2383 (N_2383,N_1506,N_1962);
nand U2384 (N_2384,N_1808,N_1757);
or U2385 (N_2385,N_1632,N_1578);
nand U2386 (N_2386,N_1887,N_1633);
nand U2387 (N_2387,N_1999,N_1549);
nand U2388 (N_2388,N_1738,N_1728);
and U2389 (N_2389,N_1803,N_1600);
nand U2390 (N_2390,N_1747,N_1836);
xor U2391 (N_2391,N_1858,N_1558);
xor U2392 (N_2392,N_1971,N_1812);
xnor U2393 (N_2393,N_1603,N_1929);
or U2394 (N_2394,N_1990,N_1625);
and U2395 (N_2395,N_1530,N_1582);
or U2396 (N_2396,N_1964,N_1743);
nor U2397 (N_2397,N_1740,N_1937);
nor U2398 (N_2398,N_1517,N_1643);
nand U2399 (N_2399,N_1562,N_1653);
and U2400 (N_2400,N_1724,N_1995);
or U2401 (N_2401,N_1508,N_1592);
nand U2402 (N_2402,N_1652,N_1600);
nand U2403 (N_2403,N_1550,N_1759);
or U2404 (N_2404,N_1854,N_1848);
nor U2405 (N_2405,N_1881,N_1501);
nor U2406 (N_2406,N_1804,N_1926);
or U2407 (N_2407,N_1586,N_1720);
nor U2408 (N_2408,N_1653,N_1675);
or U2409 (N_2409,N_1620,N_1887);
nor U2410 (N_2410,N_1621,N_1860);
or U2411 (N_2411,N_1913,N_1550);
nand U2412 (N_2412,N_1774,N_1696);
nand U2413 (N_2413,N_1737,N_1752);
xnor U2414 (N_2414,N_1795,N_1668);
or U2415 (N_2415,N_1829,N_1586);
nand U2416 (N_2416,N_1719,N_1845);
nor U2417 (N_2417,N_1620,N_1593);
and U2418 (N_2418,N_1603,N_1714);
or U2419 (N_2419,N_1520,N_1848);
xnor U2420 (N_2420,N_1955,N_1763);
xor U2421 (N_2421,N_1733,N_1783);
xnor U2422 (N_2422,N_1583,N_1832);
and U2423 (N_2423,N_1555,N_1930);
and U2424 (N_2424,N_1972,N_1857);
and U2425 (N_2425,N_1577,N_1774);
xor U2426 (N_2426,N_1941,N_1930);
or U2427 (N_2427,N_1587,N_1793);
nor U2428 (N_2428,N_1524,N_1664);
and U2429 (N_2429,N_1733,N_1884);
nand U2430 (N_2430,N_1749,N_1566);
nand U2431 (N_2431,N_1933,N_1726);
nand U2432 (N_2432,N_1608,N_1979);
and U2433 (N_2433,N_1524,N_1788);
and U2434 (N_2434,N_1833,N_1985);
or U2435 (N_2435,N_1688,N_1652);
nor U2436 (N_2436,N_1592,N_1853);
nand U2437 (N_2437,N_1695,N_1989);
xnor U2438 (N_2438,N_1840,N_1703);
nand U2439 (N_2439,N_1502,N_1649);
nand U2440 (N_2440,N_1534,N_1938);
xnor U2441 (N_2441,N_1791,N_1566);
or U2442 (N_2442,N_1725,N_1514);
and U2443 (N_2443,N_1993,N_1931);
or U2444 (N_2444,N_1917,N_1597);
nor U2445 (N_2445,N_1913,N_1758);
nand U2446 (N_2446,N_1709,N_1622);
and U2447 (N_2447,N_1859,N_1705);
nor U2448 (N_2448,N_1840,N_1668);
or U2449 (N_2449,N_1975,N_1971);
and U2450 (N_2450,N_1841,N_1633);
and U2451 (N_2451,N_1585,N_1789);
nor U2452 (N_2452,N_1517,N_1887);
and U2453 (N_2453,N_1582,N_1994);
nor U2454 (N_2454,N_1974,N_1705);
nand U2455 (N_2455,N_1765,N_1839);
nand U2456 (N_2456,N_1783,N_1761);
nor U2457 (N_2457,N_1964,N_1971);
nand U2458 (N_2458,N_1814,N_1580);
or U2459 (N_2459,N_1715,N_1978);
nand U2460 (N_2460,N_1971,N_1695);
xor U2461 (N_2461,N_1889,N_1778);
nor U2462 (N_2462,N_1546,N_1687);
nand U2463 (N_2463,N_1633,N_1912);
and U2464 (N_2464,N_1798,N_1604);
xnor U2465 (N_2465,N_1951,N_1751);
nor U2466 (N_2466,N_1502,N_1935);
and U2467 (N_2467,N_1666,N_1972);
nand U2468 (N_2468,N_1787,N_1503);
nor U2469 (N_2469,N_1573,N_1956);
nand U2470 (N_2470,N_1636,N_1680);
nand U2471 (N_2471,N_1908,N_1945);
nand U2472 (N_2472,N_1958,N_1845);
nand U2473 (N_2473,N_1543,N_1821);
nand U2474 (N_2474,N_1926,N_1747);
nor U2475 (N_2475,N_1811,N_1765);
nor U2476 (N_2476,N_1851,N_1516);
xor U2477 (N_2477,N_1746,N_1855);
nor U2478 (N_2478,N_1643,N_1949);
xor U2479 (N_2479,N_1923,N_1766);
and U2480 (N_2480,N_1601,N_1889);
nand U2481 (N_2481,N_1608,N_1688);
xor U2482 (N_2482,N_1651,N_1574);
or U2483 (N_2483,N_1883,N_1878);
nor U2484 (N_2484,N_1599,N_1800);
nor U2485 (N_2485,N_1738,N_1745);
nor U2486 (N_2486,N_1944,N_1713);
nand U2487 (N_2487,N_1522,N_1816);
nand U2488 (N_2488,N_1606,N_1607);
or U2489 (N_2489,N_1765,N_1891);
or U2490 (N_2490,N_1795,N_1545);
or U2491 (N_2491,N_1792,N_1592);
or U2492 (N_2492,N_1804,N_1940);
xor U2493 (N_2493,N_1668,N_1660);
nand U2494 (N_2494,N_1631,N_1715);
nor U2495 (N_2495,N_1710,N_1544);
nand U2496 (N_2496,N_1874,N_1814);
nand U2497 (N_2497,N_1958,N_1628);
nand U2498 (N_2498,N_1501,N_1768);
or U2499 (N_2499,N_1559,N_1635);
nor U2500 (N_2500,N_2496,N_2060);
or U2501 (N_2501,N_2119,N_2059);
nand U2502 (N_2502,N_2354,N_2222);
nand U2503 (N_2503,N_2282,N_2007);
and U2504 (N_2504,N_2233,N_2068);
and U2505 (N_2505,N_2482,N_2458);
nand U2506 (N_2506,N_2070,N_2263);
nor U2507 (N_2507,N_2046,N_2480);
or U2508 (N_2508,N_2398,N_2189);
or U2509 (N_2509,N_2157,N_2173);
nand U2510 (N_2510,N_2089,N_2112);
xnor U2511 (N_2511,N_2330,N_2341);
xor U2512 (N_2512,N_2388,N_2475);
nand U2513 (N_2513,N_2350,N_2323);
or U2514 (N_2514,N_2013,N_2403);
or U2515 (N_2515,N_2163,N_2250);
or U2516 (N_2516,N_2208,N_2420);
or U2517 (N_2517,N_2061,N_2289);
and U2518 (N_2518,N_2066,N_2078);
nand U2519 (N_2519,N_2453,N_2164);
nor U2520 (N_2520,N_2399,N_2127);
nand U2521 (N_2521,N_2082,N_2045);
nor U2522 (N_2522,N_2073,N_2311);
nor U2523 (N_2523,N_2260,N_2331);
nor U2524 (N_2524,N_2452,N_2246);
nor U2525 (N_2525,N_2322,N_2108);
nand U2526 (N_2526,N_2477,N_2154);
nand U2527 (N_2527,N_2469,N_2143);
nor U2528 (N_2528,N_2237,N_2069);
xor U2529 (N_2529,N_2032,N_2382);
or U2530 (N_2530,N_2367,N_2156);
or U2531 (N_2531,N_2472,N_2318);
xor U2532 (N_2532,N_2002,N_2328);
xor U2533 (N_2533,N_2229,N_2080);
and U2534 (N_2534,N_2215,N_2410);
or U2535 (N_2535,N_2014,N_2280);
or U2536 (N_2536,N_2489,N_2201);
and U2537 (N_2537,N_2174,N_2255);
and U2538 (N_2538,N_2417,N_2168);
nor U2539 (N_2539,N_2374,N_2493);
nor U2540 (N_2540,N_2353,N_2401);
or U2541 (N_2541,N_2220,N_2232);
nor U2542 (N_2542,N_2266,N_2492);
nand U2543 (N_2543,N_2126,N_2451);
xnor U2544 (N_2544,N_2017,N_2104);
nand U2545 (N_2545,N_2314,N_2240);
xor U2546 (N_2546,N_2213,N_2351);
xor U2547 (N_2547,N_2251,N_2212);
or U2548 (N_2548,N_2425,N_2186);
xnor U2549 (N_2549,N_2299,N_2498);
xor U2550 (N_2550,N_2079,N_2057);
or U2551 (N_2551,N_2055,N_2308);
nor U2552 (N_2552,N_2029,N_2359);
nor U2553 (N_2553,N_2144,N_2394);
or U2554 (N_2554,N_2239,N_2333);
nor U2555 (N_2555,N_2204,N_2358);
nor U2556 (N_2556,N_2022,N_2352);
xnor U2557 (N_2557,N_2162,N_2261);
and U2558 (N_2558,N_2443,N_2265);
nand U2559 (N_2559,N_2150,N_2310);
and U2560 (N_2560,N_2490,N_2194);
nor U2561 (N_2561,N_2281,N_2063);
and U2562 (N_2562,N_2210,N_2052);
nand U2563 (N_2563,N_2205,N_2161);
nor U2564 (N_2564,N_2486,N_2244);
or U2565 (N_2565,N_2015,N_2378);
and U2566 (N_2566,N_2437,N_2192);
xor U2567 (N_2567,N_2187,N_2409);
nand U2568 (N_2568,N_2102,N_2040);
and U2569 (N_2569,N_2304,N_2421);
or U2570 (N_2570,N_2054,N_2376);
or U2571 (N_2571,N_2169,N_2277);
nor U2572 (N_2572,N_2305,N_2243);
xnor U2573 (N_2573,N_2468,N_2448);
or U2574 (N_2574,N_2036,N_2396);
nand U2575 (N_2575,N_2444,N_2294);
nor U2576 (N_2576,N_2345,N_2418);
and U2577 (N_2577,N_2268,N_2141);
xnor U2578 (N_2578,N_2198,N_2435);
xnor U2579 (N_2579,N_2130,N_2349);
nand U2580 (N_2580,N_2090,N_2175);
nand U2581 (N_2581,N_2034,N_2447);
nand U2582 (N_2582,N_2365,N_2439);
nor U2583 (N_2583,N_2338,N_2211);
nand U2584 (N_2584,N_2147,N_2180);
nor U2585 (N_2585,N_2491,N_2302);
xnor U2586 (N_2586,N_2326,N_2113);
xor U2587 (N_2587,N_2160,N_2193);
nand U2588 (N_2588,N_2424,N_2231);
xnor U2589 (N_2589,N_2494,N_2320);
xnor U2590 (N_2590,N_2414,N_2171);
xnor U2591 (N_2591,N_2086,N_2380);
and U2592 (N_2592,N_2463,N_2096);
xnor U2593 (N_2593,N_2481,N_2332);
nor U2594 (N_2594,N_2075,N_2190);
or U2595 (N_2595,N_2456,N_2118);
nand U2596 (N_2596,N_2253,N_2436);
or U2597 (N_2597,N_2158,N_2364);
or U2598 (N_2598,N_2392,N_2021);
nor U2599 (N_2599,N_2223,N_2440);
nand U2600 (N_2600,N_2050,N_2362);
or U2601 (N_2601,N_2134,N_2249);
or U2602 (N_2602,N_2296,N_2179);
nor U2603 (N_2603,N_2219,N_2167);
xor U2604 (N_2604,N_2183,N_2001);
or U2605 (N_2605,N_2303,N_2487);
nor U2606 (N_2606,N_2043,N_2321);
nand U2607 (N_2607,N_2360,N_2495);
or U2608 (N_2608,N_2159,N_2081);
xnor U2609 (N_2609,N_2041,N_2407);
nand U2610 (N_2610,N_2467,N_2473);
nor U2611 (N_2611,N_2300,N_2085);
xnor U2612 (N_2612,N_2207,N_2415);
or U2613 (N_2613,N_2419,N_2301);
nand U2614 (N_2614,N_2293,N_2267);
xnor U2615 (N_2615,N_2408,N_2252);
nor U2616 (N_2616,N_2044,N_2372);
xor U2617 (N_2617,N_2076,N_2003);
nand U2618 (N_2618,N_2065,N_2139);
xor U2619 (N_2619,N_2295,N_2151);
nand U2620 (N_2620,N_2049,N_2368);
xor U2621 (N_2621,N_2165,N_2088);
or U2622 (N_2622,N_2384,N_2258);
nor U2623 (N_2623,N_2383,N_2307);
or U2624 (N_2624,N_2274,N_2459);
or U2625 (N_2625,N_2100,N_2020);
nand U2626 (N_2626,N_2325,N_2272);
nor U2627 (N_2627,N_2202,N_2483);
xnor U2628 (N_2628,N_2016,N_2259);
xor U2629 (N_2629,N_2412,N_2371);
or U2630 (N_2630,N_2319,N_2128);
nor U2631 (N_2631,N_2074,N_2117);
nor U2632 (N_2632,N_2099,N_2006);
and U2633 (N_2633,N_2133,N_2288);
nand U2634 (N_2634,N_2111,N_2230);
nor U2635 (N_2635,N_2037,N_2423);
nand U2636 (N_2636,N_2226,N_2460);
xnor U2637 (N_2637,N_2093,N_2428);
nand U2638 (N_2638,N_2142,N_2279);
and U2639 (N_2639,N_2416,N_2047);
or U2640 (N_2640,N_2287,N_2347);
and U2641 (N_2641,N_2071,N_2257);
nor U2642 (N_2642,N_2094,N_2334);
nand U2643 (N_2643,N_2286,N_2324);
nand U2644 (N_2644,N_2309,N_2195);
and U2645 (N_2645,N_2434,N_2373);
and U2646 (N_2646,N_2217,N_2355);
xor U2647 (N_2647,N_2449,N_2234);
xor U2648 (N_2648,N_2038,N_2011);
and U2649 (N_2649,N_2395,N_2077);
xor U2650 (N_2650,N_2339,N_2273);
and U2651 (N_2651,N_2084,N_2209);
xnor U2652 (N_2652,N_2397,N_2177);
xor U2653 (N_2653,N_2402,N_2290);
and U2654 (N_2654,N_2181,N_2457);
nand U2655 (N_2655,N_2297,N_2124);
nand U2656 (N_2656,N_2245,N_2389);
nand U2657 (N_2657,N_2116,N_2363);
and U2658 (N_2658,N_2152,N_2275);
and U2659 (N_2659,N_2433,N_2026);
or U2660 (N_2660,N_2479,N_2067);
and U2661 (N_2661,N_2337,N_2361);
nor U2662 (N_2662,N_2225,N_2441);
nor U2663 (N_2663,N_2466,N_2101);
nand U2664 (N_2664,N_2129,N_2461);
or U2665 (N_2665,N_2499,N_2357);
and U2666 (N_2666,N_2271,N_2283);
and U2667 (N_2667,N_2140,N_2091);
nor U2668 (N_2668,N_2270,N_2474);
nor U2669 (N_2669,N_2053,N_2476);
or U2670 (N_2670,N_2377,N_2125);
nor U2671 (N_2671,N_2199,N_2454);
nor U2672 (N_2672,N_2484,N_2188);
xor U2673 (N_2673,N_2196,N_2122);
nand U2674 (N_2674,N_2284,N_2182);
nor U2675 (N_2675,N_2422,N_2432);
nor U2676 (N_2676,N_2132,N_2012);
xnor U2677 (N_2677,N_2306,N_2107);
nand U2678 (N_2678,N_2115,N_2135);
nor U2679 (N_2679,N_2241,N_2413);
nand U2680 (N_2680,N_2327,N_2455);
and U2681 (N_2681,N_2291,N_2264);
or U2682 (N_2682,N_2411,N_2276);
nor U2683 (N_2683,N_2316,N_2375);
nand U2684 (N_2684,N_2064,N_2004);
and U2685 (N_2685,N_2184,N_2470);
or U2686 (N_2686,N_2200,N_2025);
or U2687 (N_2687,N_2406,N_2248);
nand U2688 (N_2688,N_2442,N_2236);
or U2689 (N_2689,N_2056,N_2247);
or U2690 (N_2690,N_2427,N_2278);
nor U2691 (N_2691,N_2137,N_2042);
and U2692 (N_2692,N_2087,N_2450);
xnor U2693 (N_2693,N_2315,N_2381);
nor U2694 (N_2694,N_2109,N_2391);
and U2695 (N_2695,N_2030,N_2018);
and U2696 (N_2696,N_2404,N_2429);
nor U2697 (N_2697,N_2010,N_2035);
nor U2698 (N_2698,N_2238,N_2340);
xor U2699 (N_2699,N_2095,N_2366);
or U2700 (N_2700,N_2039,N_2138);
xnor U2701 (N_2701,N_2228,N_2446);
or U2702 (N_2702,N_2083,N_2072);
xnor U2703 (N_2703,N_2058,N_2256);
and U2704 (N_2704,N_2336,N_2254);
nand U2705 (N_2705,N_2235,N_2145);
nor U2706 (N_2706,N_2146,N_2464);
nor U2707 (N_2707,N_2062,N_2206);
nor U2708 (N_2708,N_2390,N_2170);
xor U2709 (N_2709,N_2028,N_2123);
or U2710 (N_2710,N_2386,N_2092);
xor U2711 (N_2711,N_2292,N_2033);
and U2712 (N_2712,N_2393,N_2048);
or U2713 (N_2713,N_2098,N_2114);
and U2714 (N_2714,N_2370,N_2426);
or U2715 (N_2715,N_2387,N_2221);
nand U2716 (N_2716,N_2348,N_2385);
xnor U2717 (N_2717,N_2103,N_2329);
xor U2718 (N_2718,N_2262,N_2136);
and U2719 (N_2719,N_2346,N_2166);
xnor U2720 (N_2720,N_2009,N_2148);
nand U2721 (N_2721,N_2488,N_2203);
or U2722 (N_2722,N_2131,N_2120);
or U2723 (N_2723,N_2343,N_2106);
nor U2724 (N_2724,N_2342,N_2379);
nor U2725 (N_2725,N_2405,N_2317);
nand U2726 (N_2726,N_2430,N_2344);
nand U2727 (N_2727,N_2155,N_2121);
nor U2728 (N_2728,N_2185,N_2197);
or U2729 (N_2729,N_2227,N_2031);
and U2730 (N_2730,N_2224,N_2218);
xnor U2731 (N_2731,N_2023,N_2214);
xnor U2732 (N_2732,N_2438,N_2172);
and U2733 (N_2733,N_2153,N_2431);
or U2734 (N_2734,N_2051,N_2176);
or U2735 (N_2735,N_2216,N_2335);
nand U2736 (N_2736,N_2445,N_2313);
nand U2737 (N_2737,N_2285,N_2465);
nor U2738 (N_2738,N_2462,N_2110);
nand U2739 (N_2739,N_2027,N_2008);
xnor U2740 (N_2740,N_2005,N_2178);
and U2741 (N_2741,N_2471,N_2356);
nand U2742 (N_2742,N_2369,N_2485);
nor U2743 (N_2743,N_2097,N_2312);
nand U2744 (N_2744,N_2019,N_2024);
or U2745 (N_2745,N_2105,N_2400);
or U2746 (N_2746,N_2298,N_2191);
nor U2747 (N_2747,N_2242,N_2269);
xnor U2748 (N_2748,N_2149,N_2000);
or U2749 (N_2749,N_2478,N_2497);
and U2750 (N_2750,N_2098,N_2401);
and U2751 (N_2751,N_2328,N_2497);
or U2752 (N_2752,N_2277,N_2225);
xor U2753 (N_2753,N_2085,N_2016);
nor U2754 (N_2754,N_2251,N_2043);
xnor U2755 (N_2755,N_2296,N_2020);
and U2756 (N_2756,N_2091,N_2335);
nand U2757 (N_2757,N_2126,N_2189);
xnor U2758 (N_2758,N_2126,N_2108);
xnor U2759 (N_2759,N_2066,N_2179);
nand U2760 (N_2760,N_2250,N_2276);
nor U2761 (N_2761,N_2459,N_2356);
or U2762 (N_2762,N_2439,N_2098);
or U2763 (N_2763,N_2187,N_2124);
nand U2764 (N_2764,N_2220,N_2279);
xnor U2765 (N_2765,N_2045,N_2317);
nor U2766 (N_2766,N_2315,N_2436);
nand U2767 (N_2767,N_2390,N_2307);
and U2768 (N_2768,N_2486,N_2064);
xnor U2769 (N_2769,N_2482,N_2481);
nor U2770 (N_2770,N_2137,N_2171);
nand U2771 (N_2771,N_2404,N_2146);
or U2772 (N_2772,N_2143,N_2362);
nor U2773 (N_2773,N_2086,N_2393);
and U2774 (N_2774,N_2108,N_2292);
and U2775 (N_2775,N_2374,N_2029);
or U2776 (N_2776,N_2311,N_2250);
and U2777 (N_2777,N_2065,N_2364);
nand U2778 (N_2778,N_2187,N_2039);
nand U2779 (N_2779,N_2085,N_2024);
nor U2780 (N_2780,N_2358,N_2129);
and U2781 (N_2781,N_2363,N_2226);
and U2782 (N_2782,N_2075,N_2379);
or U2783 (N_2783,N_2195,N_2308);
nor U2784 (N_2784,N_2085,N_2342);
and U2785 (N_2785,N_2042,N_2232);
nand U2786 (N_2786,N_2115,N_2432);
nand U2787 (N_2787,N_2228,N_2082);
or U2788 (N_2788,N_2117,N_2238);
xnor U2789 (N_2789,N_2277,N_2286);
or U2790 (N_2790,N_2227,N_2236);
nor U2791 (N_2791,N_2260,N_2392);
nand U2792 (N_2792,N_2210,N_2461);
nand U2793 (N_2793,N_2137,N_2384);
xor U2794 (N_2794,N_2129,N_2100);
and U2795 (N_2795,N_2162,N_2316);
nand U2796 (N_2796,N_2116,N_2383);
nor U2797 (N_2797,N_2105,N_2371);
nand U2798 (N_2798,N_2159,N_2183);
nor U2799 (N_2799,N_2110,N_2451);
nand U2800 (N_2800,N_2141,N_2472);
or U2801 (N_2801,N_2357,N_2436);
nor U2802 (N_2802,N_2387,N_2233);
and U2803 (N_2803,N_2430,N_2101);
nand U2804 (N_2804,N_2003,N_2132);
nand U2805 (N_2805,N_2265,N_2199);
nor U2806 (N_2806,N_2451,N_2415);
or U2807 (N_2807,N_2229,N_2273);
nand U2808 (N_2808,N_2497,N_2031);
or U2809 (N_2809,N_2266,N_2135);
nand U2810 (N_2810,N_2153,N_2368);
or U2811 (N_2811,N_2208,N_2446);
nand U2812 (N_2812,N_2306,N_2069);
and U2813 (N_2813,N_2065,N_2374);
nand U2814 (N_2814,N_2401,N_2115);
or U2815 (N_2815,N_2440,N_2434);
xor U2816 (N_2816,N_2297,N_2271);
xor U2817 (N_2817,N_2481,N_2047);
nand U2818 (N_2818,N_2071,N_2211);
nor U2819 (N_2819,N_2224,N_2213);
nor U2820 (N_2820,N_2139,N_2237);
or U2821 (N_2821,N_2278,N_2239);
or U2822 (N_2822,N_2145,N_2173);
nor U2823 (N_2823,N_2262,N_2431);
or U2824 (N_2824,N_2473,N_2138);
nand U2825 (N_2825,N_2134,N_2286);
or U2826 (N_2826,N_2358,N_2302);
nand U2827 (N_2827,N_2346,N_2194);
and U2828 (N_2828,N_2476,N_2423);
xor U2829 (N_2829,N_2193,N_2416);
nor U2830 (N_2830,N_2185,N_2099);
and U2831 (N_2831,N_2096,N_2338);
xnor U2832 (N_2832,N_2472,N_2406);
nand U2833 (N_2833,N_2152,N_2476);
or U2834 (N_2834,N_2482,N_2231);
nor U2835 (N_2835,N_2411,N_2272);
and U2836 (N_2836,N_2261,N_2068);
and U2837 (N_2837,N_2312,N_2204);
nand U2838 (N_2838,N_2326,N_2313);
or U2839 (N_2839,N_2094,N_2342);
and U2840 (N_2840,N_2150,N_2327);
and U2841 (N_2841,N_2208,N_2060);
or U2842 (N_2842,N_2491,N_2267);
nor U2843 (N_2843,N_2270,N_2367);
nand U2844 (N_2844,N_2084,N_2044);
nand U2845 (N_2845,N_2115,N_2302);
and U2846 (N_2846,N_2102,N_2023);
nor U2847 (N_2847,N_2430,N_2266);
nand U2848 (N_2848,N_2234,N_2260);
nor U2849 (N_2849,N_2052,N_2046);
nor U2850 (N_2850,N_2488,N_2029);
nand U2851 (N_2851,N_2485,N_2097);
nand U2852 (N_2852,N_2064,N_2483);
xnor U2853 (N_2853,N_2057,N_2019);
xnor U2854 (N_2854,N_2298,N_2474);
or U2855 (N_2855,N_2205,N_2470);
and U2856 (N_2856,N_2395,N_2251);
and U2857 (N_2857,N_2394,N_2160);
xor U2858 (N_2858,N_2372,N_2482);
and U2859 (N_2859,N_2111,N_2270);
nand U2860 (N_2860,N_2327,N_2159);
xnor U2861 (N_2861,N_2427,N_2261);
and U2862 (N_2862,N_2489,N_2011);
xor U2863 (N_2863,N_2291,N_2424);
nand U2864 (N_2864,N_2256,N_2499);
and U2865 (N_2865,N_2032,N_2215);
and U2866 (N_2866,N_2011,N_2183);
or U2867 (N_2867,N_2464,N_2273);
nand U2868 (N_2868,N_2337,N_2405);
or U2869 (N_2869,N_2350,N_2336);
xnor U2870 (N_2870,N_2045,N_2043);
xor U2871 (N_2871,N_2411,N_2392);
nor U2872 (N_2872,N_2181,N_2454);
and U2873 (N_2873,N_2441,N_2316);
xnor U2874 (N_2874,N_2120,N_2056);
nand U2875 (N_2875,N_2389,N_2305);
and U2876 (N_2876,N_2275,N_2403);
nand U2877 (N_2877,N_2176,N_2010);
xnor U2878 (N_2878,N_2279,N_2219);
nand U2879 (N_2879,N_2234,N_2249);
nand U2880 (N_2880,N_2260,N_2467);
xor U2881 (N_2881,N_2051,N_2247);
and U2882 (N_2882,N_2440,N_2199);
nor U2883 (N_2883,N_2228,N_2239);
xnor U2884 (N_2884,N_2023,N_2298);
nor U2885 (N_2885,N_2219,N_2094);
nor U2886 (N_2886,N_2421,N_2416);
or U2887 (N_2887,N_2490,N_2223);
or U2888 (N_2888,N_2237,N_2092);
and U2889 (N_2889,N_2192,N_2262);
and U2890 (N_2890,N_2098,N_2015);
xor U2891 (N_2891,N_2486,N_2090);
nand U2892 (N_2892,N_2313,N_2118);
nand U2893 (N_2893,N_2345,N_2228);
nor U2894 (N_2894,N_2289,N_2082);
or U2895 (N_2895,N_2481,N_2411);
nand U2896 (N_2896,N_2421,N_2010);
nor U2897 (N_2897,N_2045,N_2205);
xor U2898 (N_2898,N_2254,N_2472);
nand U2899 (N_2899,N_2419,N_2314);
and U2900 (N_2900,N_2247,N_2305);
and U2901 (N_2901,N_2057,N_2116);
nand U2902 (N_2902,N_2302,N_2477);
and U2903 (N_2903,N_2254,N_2015);
nor U2904 (N_2904,N_2373,N_2461);
xor U2905 (N_2905,N_2147,N_2009);
nor U2906 (N_2906,N_2430,N_2186);
or U2907 (N_2907,N_2266,N_2319);
and U2908 (N_2908,N_2466,N_2353);
xnor U2909 (N_2909,N_2089,N_2050);
xor U2910 (N_2910,N_2054,N_2224);
nor U2911 (N_2911,N_2372,N_2347);
nand U2912 (N_2912,N_2484,N_2394);
or U2913 (N_2913,N_2039,N_2143);
nor U2914 (N_2914,N_2176,N_2458);
or U2915 (N_2915,N_2133,N_2472);
or U2916 (N_2916,N_2345,N_2415);
nor U2917 (N_2917,N_2429,N_2311);
nand U2918 (N_2918,N_2373,N_2221);
nand U2919 (N_2919,N_2251,N_2340);
nor U2920 (N_2920,N_2075,N_2179);
xor U2921 (N_2921,N_2361,N_2370);
nor U2922 (N_2922,N_2055,N_2433);
xnor U2923 (N_2923,N_2061,N_2137);
xor U2924 (N_2924,N_2132,N_2202);
or U2925 (N_2925,N_2105,N_2050);
nand U2926 (N_2926,N_2056,N_2473);
and U2927 (N_2927,N_2253,N_2229);
and U2928 (N_2928,N_2198,N_2102);
xnor U2929 (N_2929,N_2087,N_2406);
and U2930 (N_2930,N_2410,N_2048);
xnor U2931 (N_2931,N_2123,N_2431);
nand U2932 (N_2932,N_2465,N_2434);
nand U2933 (N_2933,N_2386,N_2376);
nand U2934 (N_2934,N_2107,N_2122);
xnor U2935 (N_2935,N_2418,N_2407);
nor U2936 (N_2936,N_2397,N_2206);
nor U2937 (N_2937,N_2269,N_2041);
or U2938 (N_2938,N_2277,N_2189);
and U2939 (N_2939,N_2344,N_2404);
xor U2940 (N_2940,N_2460,N_2283);
and U2941 (N_2941,N_2180,N_2061);
nor U2942 (N_2942,N_2328,N_2436);
nand U2943 (N_2943,N_2473,N_2463);
or U2944 (N_2944,N_2111,N_2316);
xnor U2945 (N_2945,N_2076,N_2382);
and U2946 (N_2946,N_2145,N_2393);
nor U2947 (N_2947,N_2352,N_2066);
and U2948 (N_2948,N_2280,N_2458);
nor U2949 (N_2949,N_2233,N_2225);
xor U2950 (N_2950,N_2264,N_2208);
or U2951 (N_2951,N_2289,N_2464);
xnor U2952 (N_2952,N_2366,N_2378);
xor U2953 (N_2953,N_2083,N_2452);
or U2954 (N_2954,N_2003,N_2291);
or U2955 (N_2955,N_2264,N_2101);
and U2956 (N_2956,N_2074,N_2245);
and U2957 (N_2957,N_2109,N_2362);
nor U2958 (N_2958,N_2079,N_2088);
nand U2959 (N_2959,N_2041,N_2413);
or U2960 (N_2960,N_2146,N_2452);
nand U2961 (N_2961,N_2242,N_2138);
xor U2962 (N_2962,N_2217,N_2023);
or U2963 (N_2963,N_2064,N_2394);
and U2964 (N_2964,N_2254,N_2498);
and U2965 (N_2965,N_2380,N_2066);
or U2966 (N_2966,N_2342,N_2040);
or U2967 (N_2967,N_2496,N_2469);
and U2968 (N_2968,N_2076,N_2183);
nand U2969 (N_2969,N_2181,N_2115);
or U2970 (N_2970,N_2233,N_2385);
nand U2971 (N_2971,N_2163,N_2091);
nand U2972 (N_2972,N_2451,N_2493);
and U2973 (N_2973,N_2205,N_2068);
and U2974 (N_2974,N_2491,N_2046);
nor U2975 (N_2975,N_2011,N_2419);
and U2976 (N_2976,N_2467,N_2137);
or U2977 (N_2977,N_2357,N_2373);
and U2978 (N_2978,N_2472,N_2113);
nand U2979 (N_2979,N_2040,N_2434);
nor U2980 (N_2980,N_2057,N_2076);
nor U2981 (N_2981,N_2444,N_2414);
xor U2982 (N_2982,N_2287,N_2245);
nand U2983 (N_2983,N_2259,N_2481);
nand U2984 (N_2984,N_2389,N_2387);
nor U2985 (N_2985,N_2280,N_2467);
nor U2986 (N_2986,N_2229,N_2002);
nor U2987 (N_2987,N_2197,N_2330);
or U2988 (N_2988,N_2440,N_2453);
nand U2989 (N_2989,N_2416,N_2272);
nor U2990 (N_2990,N_2281,N_2421);
nand U2991 (N_2991,N_2305,N_2146);
nand U2992 (N_2992,N_2381,N_2019);
nor U2993 (N_2993,N_2452,N_2325);
and U2994 (N_2994,N_2474,N_2002);
or U2995 (N_2995,N_2201,N_2270);
and U2996 (N_2996,N_2218,N_2391);
nand U2997 (N_2997,N_2452,N_2223);
nand U2998 (N_2998,N_2221,N_2423);
and U2999 (N_2999,N_2337,N_2078);
or U3000 (N_3000,N_2884,N_2966);
xor U3001 (N_3001,N_2643,N_2736);
nand U3002 (N_3002,N_2975,N_2943);
or U3003 (N_3003,N_2754,N_2729);
xnor U3004 (N_3004,N_2922,N_2624);
nor U3005 (N_3005,N_2569,N_2585);
nand U3006 (N_3006,N_2766,N_2573);
nand U3007 (N_3007,N_2537,N_2633);
nor U3008 (N_3008,N_2807,N_2750);
nand U3009 (N_3009,N_2618,N_2666);
and U3010 (N_3010,N_2731,N_2920);
or U3011 (N_3011,N_2743,N_2518);
and U3012 (N_3012,N_2656,N_2911);
or U3013 (N_3013,N_2741,N_2775);
nand U3014 (N_3014,N_2749,N_2699);
nor U3015 (N_3015,N_2799,N_2578);
nand U3016 (N_3016,N_2780,N_2562);
or U3017 (N_3017,N_2814,N_2613);
nand U3018 (N_3018,N_2925,N_2710);
nand U3019 (N_3019,N_2521,N_2846);
and U3020 (N_3020,N_2730,N_2860);
or U3021 (N_3021,N_2689,N_2813);
and U3022 (N_3022,N_2524,N_2734);
or U3023 (N_3023,N_2529,N_2752);
xor U3024 (N_3024,N_2803,N_2921);
xnor U3025 (N_3025,N_2659,N_2602);
and U3026 (N_3026,N_2984,N_2923);
nand U3027 (N_3027,N_2703,N_2888);
and U3028 (N_3028,N_2548,N_2830);
or U3029 (N_3029,N_2989,N_2856);
nor U3030 (N_3030,N_2982,N_2778);
nand U3031 (N_3031,N_2886,N_2636);
or U3032 (N_3032,N_2959,N_2988);
nor U3033 (N_3033,N_2854,N_2941);
nand U3034 (N_3034,N_2961,N_2620);
xnor U3035 (N_3035,N_2552,N_2576);
and U3036 (N_3036,N_2565,N_2883);
and U3037 (N_3037,N_2842,N_2963);
or U3038 (N_3038,N_2769,N_2616);
nand U3039 (N_3039,N_2822,N_2639);
xnor U3040 (N_3040,N_2628,N_2867);
xnor U3041 (N_3041,N_2833,N_2700);
or U3042 (N_3042,N_2787,N_2800);
nand U3043 (N_3043,N_2789,N_2535);
xnor U3044 (N_3044,N_2516,N_2645);
and U3045 (N_3045,N_2680,N_2508);
or U3046 (N_3046,N_2952,N_2735);
xor U3047 (N_3047,N_2933,N_2834);
or U3048 (N_3048,N_2938,N_2725);
nand U3049 (N_3049,N_2993,N_2575);
nand U3050 (N_3050,N_2983,N_2679);
nor U3051 (N_3051,N_2779,N_2968);
nand U3052 (N_3052,N_2603,N_2517);
nor U3053 (N_3053,N_2642,N_2905);
xor U3054 (N_3054,N_2572,N_2885);
nand U3055 (N_3055,N_2994,N_2976);
xor U3056 (N_3056,N_2733,N_2678);
xnor U3057 (N_3057,N_2969,N_2559);
nand U3058 (N_3058,N_2683,N_2568);
xnor U3059 (N_3059,N_2835,N_2770);
and U3060 (N_3060,N_2870,N_2723);
xor U3061 (N_3061,N_2964,N_2740);
or U3062 (N_3062,N_2672,N_2999);
xor U3063 (N_3063,N_2738,N_2978);
nor U3064 (N_3064,N_2605,N_2687);
xnor U3065 (N_3065,N_2881,N_2717);
nor U3066 (N_3066,N_2808,N_2998);
or U3067 (N_3067,N_2534,N_2853);
and U3068 (N_3068,N_2875,N_2630);
nor U3069 (N_3069,N_2928,N_2893);
xor U3070 (N_3070,N_2691,N_2509);
nand U3071 (N_3071,N_2759,N_2845);
nand U3072 (N_3072,N_2582,N_2797);
nor U3073 (N_3073,N_2614,N_2855);
or U3074 (N_3074,N_2781,N_2598);
and U3075 (N_3075,N_2806,N_2542);
xnor U3076 (N_3076,N_2694,N_2580);
xnor U3077 (N_3077,N_2929,N_2589);
xnor U3078 (N_3078,N_2669,N_2953);
nand U3079 (N_3079,N_2536,N_2757);
nor U3080 (N_3080,N_2866,N_2545);
or U3081 (N_3081,N_2556,N_2748);
and U3082 (N_3082,N_2939,N_2879);
nand U3083 (N_3083,N_2902,N_2530);
nor U3084 (N_3084,N_2810,N_2591);
nor U3085 (N_3085,N_2711,N_2991);
and U3086 (N_3086,N_2593,N_2840);
or U3087 (N_3087,N_2506,N_2995);
or U3088 (N_3088,N_2507,N_2728);
nor U3089 (N_3089,N_2957,N_2702);
nor U3090 (N_3090,N_2617,N_2528);
nand U3091 (N_3091,N_2726,N_2944);
xor U3092 (N_3092,N_2931,N_2651);
and U3093 (N_3093,N_2505,N_2918);
or U3094 (N_3094,N_2632,N_2560);
or U3095 (N_3095,N_2761,N_2502);
xor U3096 (N_3096,N_2954,N_2934);
or U3097 (N_3097,N_2608,N_2732);
and U3098 (N_3098,N_2551,N_2563);
nand U3099 (N_3099,N_2708,N_2772);
or U3100 (N_3100,N_2531,N_2972);
xor U3101 (N_3101,N_2951,N_2892);
and U3102 (N_3102,N_2558,N_2587);
xnor U3103 (N_3103,N_2555,N_2627);
nand U3104 (N_3104,N_2827,N_2841);
and U3105 (N_3105,N_2675,N_2739);
nor U3106 (N_3106,N_2671,N_2705);
nor U3107 (N_3107,N_2626,N_2650);
nand U3108 (N_3108,N_2622,N_2852);
nand U3109 (N_3109,N_2844,N_2997);
nor U3110 (N_3110,N_2566,N_2597);
and U3111 (N_3111,N_2824,N_2936);
nor U3112 (N_3112,N_2512,N_2544);
nor U3113 (N_3113,N_2592,N_2670);
nor U3114 (N_3114,N_2791,N_2977);
nor U3115 (N_3115,N_2801,N_2706);
and U3116 (N_3116,N_2623,N_2527);
and U3117 (N_3117,N_2547,N_2693);
nor U3118 (N_3118,N_2586,N_2831);
and U3119 (N_3119,N_2567,N_2600);
xnor U3120 (N_3120,N_2655,N_2774);
and U3121 (N_3121,N_2912,N_2599);
and U3122 (N_3122,N_2719,N_2677);
xnor U3123 (N_3123,N_2965,N_2784);
and U3124 (N_3124,N_2557,N_2817);
xor U3125 (N_3125,N_2660,N_2596);
nand U3126 (N_3126,N_2909,N_2947);
nand U3127 (N_3127,N_2526,N_2832);
or U3128 (N_3128,N_2756,N_2686);
nand U3129 (N_3129,N_2930,N_2663);
and U3130 (N_3130,N_2980,N_2762);
and U3131 (N_3131,N_2891,N_2768);
nand U3132 (N_3132,N_2744,N_2794);
nand U3133 (N_3133,N_2601,N_2877);
and U3134 (N_3134,N_2776,N_2970);
nor U3135 (N_3135,N_2820,N_2927);
xnor U3136 (N_3136,N_2960,N_2942);
and U3137 (N_3137,N_2788,N_2652);
xnor U3138 (N_3138,N_2570,N_2751);
xor U3139 (N_3139,N_2937,N_2525);
nor U3140 (N_3140,N_2619,N_2747);
nand U3141 (N_3141,N_2900,N_2823);
nand U3142 (N_3142,N_2745,N_2985);
nand U3143 (N_3143,N_2802,N_2815);
and U3144 (N_3144,N_2819,N_2859);
or U3145 (N_3145,N_2588,N_2501);
nand U3146 (N_3146,N_2654,N_2539);
or U3147 (N_3147,N_2812,N_2796);
or U3148 (N_3148,N_2849,N_2707);
xor U3149 (N_3149,N_2722,N_2955);
nor U3150 (N_3150,N_2821,N_2755);
xor U3151 (N_3151,N_2520,N_2661);
and U3152 (N_3152,N_2790,N_2986);
nor U3153 (N_3153,N_2504,N_2716);
xnor U3154 (N_3154,N_2899,N_2514);
nor U3155 (N_3155,N_2667,N_2746);
nor U3156 (N_3156,N_2783,N_2843);
and U3157 (N_3157,N_2742,N_2657);
nor U3158 (N_3158,N_2901,N_2915);
and U3159 (N_3159,N_2887,N_2906);
nor U3160 (N_3160,N_2704,N_2973);
nand U3161 (N_3161,N_2873,N_2763);
nor U3162 (N_3162,N_2904,N_2869);
nand U3163 (N_3163,N_2607,N_2577);
nand U3164 (N_3164,N_2992,N_2647);
nand U3165 (N_3165,N_2919,N_2631);
nor U3166 (N_3166,N_2868,N_2718);
nor U3167 (N_3167,N_2908,N_2910);
nand U3168 (N_3168,N_2753,N_2611);
or U3169 (N_3169,N_2805,N_2851);
nor U3170 (N_3170,N_2981,N_2625);
nor U3171 (N_3171,N_2898,N_2971);
and U3172 (N_3172,N_2554,N_2863);
or U3173 (N_3173,N_2786,N_2850);
xnor U3174 (N_3174,N_2523,N_2701);
xnor U3175 (N_3175,N_2510,N_2727);
or U3176 (N_3176,N_2698,N_2811);
nor U3177 (N_3177,N_2609,N_2816);
xor U3178 (N_3178,N_2945,N_2838);
or U3179 (N_3179,N_2940,N_2950);
nand U3180 (N_3180,N_2914,N_2878);
and U3181 (N_3181,N_2690,N_2764);
nor U3182 (N_3182,N_2546,N_2581);
nand U3183 (N_3183,N_2682,N_2533);
nand U3184 (N_3184,N_2583,N_2635);
nand U3185 (N_3185,N_2584,N_2847);
nor U3186 (N_3186,N_2697,N_2829);
nor U3187 (N_3187,N_2695,N_2681);
nand U3188 (N_3188,N_2662,N_2871);
xor U3189 (N_3189,N_2897,N_2839);
nor U3190 (N_3190,N_2511,N_2604);
or U3191 (N_3191,N_2688,N_2962);
or U3192 (N_3192,N_2709,N_2967);
xor U3193 (N_3193,N_2907,N_2500);
nor U3194 (N_3194,N_2519,N_2595);
nor U3195 (N_3195,N_2612,N_2522);
or U3196 (N_3196,N_2638,N_2550);
or U3197 (N_3197,N_2880,N_2538);
and U3198 (N_3198,N_2996,N_2513);
and U3199 (N_3199,N_2795,N_2858);
and U3200 (N_3200,N_2621,N_2895);
nor U3201 (N_3201,N_2825,N_2692);
nor U3202 (N_3202,N_2714,N_2653);
nand U3203 (N_3203,N_2615,N_2658);
nor U3204 (N_3204,N_2861,N_2958);
xnor U3205 (N_3205,N_2673,N_2646);
xnor U3206 (N_3206,N_2932,N_2674);
nand U3207 (N_3207,N_2553,N_2828);
nand U3208 (N_3208,N_2640,N_2724);
nand U3209 (N_3209,N_2804,N_2579);
or U3210 (N_3210,N_2715,N_2629);
nor U3211 (N_3211,N_2760,N_2862);
xnor U3212 (N_3212,N_2872,N_2903);
and U3213 (N_3213,N_2540,N_2889);
or U3214 (N_3214,N_2890,N_2935);
or U3215 (N_3215,N_2637,N_2956);
nand U3216 (N_3216,N_2590,N_2987);
nor U3217 (N_3217,N_2594,N_2765);
or U3218 (N_3218,N_2515,N_2644);
nand U3219 (N_3219,N_2571,N_2713);
or U3220 (N_3220,N_2668,N_2696);
and U3221 (N_3221,N_2874,N_2649);
nor U3222 (N_3222,N_2773,N_2606);
nand U3223 (N_3223,N_2798,N_2837);
nor U3224 (N_3224,N_2864,N_2946);
and U3225 (N_3225,N_2712,N_2665);
xor U3226 (N_3226,N_2782,N_2541);
nand U3227 (N_3227,N_2503,N_2721);
nand U3228 (N_3228,N_2684,N_2641);
and U3229 (N_3229,N_2826,N_2543);
and U3230 (N_3230,N_2924,N_2882);
and U3231 (N_3231,N_2865,N_2990);
nand U3232 (N_3232,N_2610,N_2926);
nand U3233 (N_3233,N_2792,N_2896);
and U3234 (N_3234,N_2676,N_2777);
xor U3235 (N_3235,N_2974,N_2634);
or U3236 (N_3236,N_2848,N_2532);
xnor U3237 (N_3237,N_2836,N_2771);
nand U3238 (N_3238,N_2574,N_2737);
nand U3239 (N_3239,N_2785,N_2767);
nor U3240 (N_3240,N_2949,N_2793);
and U3241 (N_3241,N_2758,N_2648);
nor U3242 (N_3242,N_2876,N_2809);
and U3243 (N_3243,N_2917,N_2720);
xor U3244 (N_3244,N_2564,N_2948);
and U3245 (N_3245,N_2894,N_2913);
nor U3246 (N_3246,N_2549,N_2561);
and U3247 (N_3247,N_2857,N_2818);
and U3248 (N_3248,N_2979,N_2664);
or U3249 (N_3249,N_2916,N_2685);
nor U3250 (N_3250,N_2687,N_2748);
nand U3251 (N_3251,N_2794,N_2577);
or U3252 (N_3252,N_2635,N_2936);
nor U3253 (N_3253,N_2926,N_2647);
nand U3254 (N_3254,N_2545,N_2649);
nor U3255 (N_3255,N_2946,N_2607);
and U3256 (N_3256,N_2650,N_2837);
nor U3257 (N_3257,N_2942,N_2632);
and U3258 (N_3258,N_2578,N_2519);
or U3259 (N_3259,N_2810,N_2892);
nand U3260 (N_3260,N_2961,N_2879);
xnor U3261 (N_3261,N_2819,N_2843);
xnor U3262 (N_3262,N_2915,N_2638);
and U3263 (N_3263,N_2846,N_2878);
nand U3264 (N_3264,N_2710,N_2939);
nand U3265 (N_3265,N_2592,N_2554);
xnor U3266 (N_3266,N_2984,N_2829);
nand U3267 (N_3267,N_2703,N_2748);
nor U3268 (N_3268,N_2590,N_2514);
xor U3269 (N_3269,N_2568,N_2565);
xor U3270 (N_3270,N_2969,N_2938);
or U3271 (N_3271,N_2677,N_2548);
nand U3272 (N_3272,N_2999,N_2626);
or U3273 (N_3273,N_2565,N_2868);
and U3274 (N_3274,N_2846,N_2550);
or U3275 (N_3275,N_2550,N_2918);
nor U3276 (N_3276,N_2860,N_2711);
nand U3277 (N_3277,N_2896,N_2646);
nor U3278 (N_3278,N_2669,N_2825);
and U3279 (N_3279,N_2513,N_2601);
and U3280 (N_3280,N_2778,N_2515);
xor U3281 (N_3281,N_2998,N_2893);
nand U3282 (N_3282,N_2727,N_2612);
nand U3283 (N_3283,N_2809,N_2700);
nand U3284 (N_3284,N_2953,N_2668);
or U3285 (N_3285,N_2618,N_2893);
nor U3286 (N_3286,N_2706,N_2960);
or U3287 (N_3287,N_2683,N_2977);
nor U3288 (N_3288,N_2655,N_2668);
nand U3289 (N_3289,N_2928,N_2972);
nor U3290 (N_3290,N_2800,N_2938);
nor U3291 (N_3291,N_2898,N_2534);
nor U3292 (N_3292,N_2773,N_2875);
and U3293 (N_3293,N_2617,N_2837);
nor U3294 (N_3294,N_2902,N_2574);
xnor U3295 (N_3295,N_2758,N_2968);
xnor U3296 (N_3296,N_2947,N_2872);
xnor U3297 (N_3297,N_2970,N_2874);
xnor U3298 (N_3298,N_2831,N_2697);
and U3299 (N_3299,N_2525,N_2872);
and U3300 (N_3300,N_2804,N_2920);
or U3301 (N_3301,N_2611,N_2734);
or U3302 (N_3302,N_2520,N_2960);
nor U3303 (N_3303,N_2958,N_2590);
nor U3304 (N_3304,N_2509,N_2987);
and U3305 (N_3305,N_2662,N_2993);
nand U3306 (N_3306,N_2820,N_2864);
or U3307 (N_3307,N_2647,N_2966);
nor U3308 (N_3308,N_2611,N_2732);
or U3309 (N_3309,N_2682,N_2694);
nand U3310 (N_3310,N_2989,N_2732);
and U3311 (N_3311,N_2583,N_2739);
and U3312 (N_3312,N_2930,N_2611);
and U3313 (N_3313,N_2950,N_2750);
nand U3314 (N_3314,N_2875,N_2827);
or U3315 (N_3315,N_2523,N_2948);
xnor U3316 (N_3316,N_2581,N_2976);
or U3317 (N_3317,N_2579,N_2814);
xor U3318 (N_3318,N_2902,N_2845);
xor U3319 (N_3319,N_2707,N_2927);
or U3320 (N_3320,N_2540,N_2825);
xnor U3321 (N_3321,N_2822,N_2779);
and U3322 (N_3322,N_2892,N_2549);
and U3323 (N_3323,N_2742,N_2937);
xnor U3324 (N_3324,N_2569,N_2757);
or U3325 (N_3325,N_2615,N_2996);
or U3326 (N_3326,N_2642,N_2672);
or U3327 (N_3327,N_2933,N_2954);
xor U3328 (N_3328,N_2684,N_2539);
or U3329 (N_3329,N_2739,N_2614);
nor U3330 (N_3330,N_2938,N_2751);
xnor U3331 (N_3331,N_2949,N_2665);
nor U3332 (N_3332,N_2895,N_2617);
nor U3333 (N_3333,N_2743,N_2535);
or U3334 (N_3334,N_2865,N_2884);
nand U3335 (N_3335,N_2663,N_2573);
and U3336 (N_3336,N_2922,N_2572);
nand U3337 (N_3337,N_2614,N_2516);
xor U3338 (N_3338,N_2659,N_2698);
or U3339 (N_3339,N_2852,N_2560);
xor U3340 (N_3340,N_2639,N_2547);
nand U3341 (N_3341,N_2817,N_2927);
and U3342 (N_3342,N_2678,N_2505);
and U3343 (N_3343,N_2897,N_2766);
or U3344 (N_3344,N_2712,N_2970);
nand U3345 (N_3345,N_2774,N_2850);
and U3346 (N_3346,N_2763,N_2619);
xnor U3347 (N_3347,N_2537,N_2984);
and U3348 (N_3348,N_2754,N_2981);
nor U3349 (N_3349,N_2849,N_2950);
nor U3350 (N_3350,N_2772,N_2550);
and U3351 (N_3351,N_2776,N_2808);
nand U3352 (N_3352,N_2995,N_2884);
and U3353 (N_3353,N_2600,N_2634);
and U3354 (N_3354,N_2770,N_2946);
xor U3355 (N_3355,N_2601,N_2564);
or U3356 (N_3356,N_2589,N_2626);
nor U3357 (N_3357,N_2696,N_2974);
and U3358 (N_3358,N_2958,N_2854);
xor U3359 (N_3359,N_2706,N_2916);
or U3360 (N_3360,N_2542,N_2721);
nand U3361 (N_3361,N_2757,N_2552);
nand U3362 (N_3362,N_2588,N_2824);
and U3363 (N_3363,N_2703,N_2629);
xnor U3364 (N_3364,N_2941,N_2647);
nor U3365 (N_3365,N_2958,N_2609);
or U3366 (N_3366,N_2744,N_2762);
or U3367 (N_3367,N_2959,N_2604);
and U3368 (N_3368,N_2707,N_2638);
nor U3369 (N_3369,N_2603,N_2548);
or U3370 (N_3370,N_2884,N_2825);
or U3371 (N_3371,N_2702,N_2584);
nand U3372 (N_3372,N_2942,N_2606);
nor U3373 (N_3373,N_2884,N_2642);
nor U3374 (N_3374,N_2932,N_2995);
or U3375 (N_3375,N_2869,N_2645);
nor U3376 (N_3376,N_2912,N_2931);
and U3377 (N_3377,N_2831,N_2965);
and U3378 (N_3378,N_2879,N_2596);
xnor U3379 (N_3379,N_2941,N_2870);
nor U3380 (N_3380,N_2627,N_2833);
nand U3381 (N_3381,N_2917,N_2503);
and U3382 (N_3382,N_2877,N_2937);
nor U3383 (N_3383,N_2502,N_2587);
nand U3384 (N_3384,N_2651,N_2584);
nand U3385 (N_3385,N_2935,N_2835);
nand U3386 (N_3386,N_2780,N_2563);
and U3387 (N_3387,N_2724,N_2649);
nand U3388 (N_3388,N_2935,N_2978);
xor U3389 (N_3389,N_2916,N_2657);
or U3390 (N_3390,N_2627,N_2908);
or U3391 (N_3391,N_2828,N_2603);
and U3392 (N_3392,N_2583,N_2903);
nand U3393 (N_3393,N_2631,N_2616);
or U3394 (N_3394,N_2827,N_2833);
or U3395 (N_3395,N_2909,N_2801);
or U3396 (N_3396,N_2669,N_2917);
xor U3397 (N_3397,N_2656,N_2825);
nand U3398 (N_3398,N_2530,N_2546);
xnor U3399 (N_3399,N_2888,N_2821);
nor U3400 (N_3400,N_2552,N_2683);
nand U3401 (N_3401,N_2503,N_2725);
and U3402 (N_3402,N_2578,N_2804);
nand U3403 (N_3403,N_2609,N_2933);
nand U3404 (N_3404,N_2511,N_2663);
or U3405 (N_3405,N_2568,N_2673);
xnor U3406 (N_3406,N_2695,N_2913);
nor U3407 (N_3407,N_2527,N_2752);
xor U3408 (N_3408,N_2667,N_2631);
nor U3409 (N_3409,N_2758,N_2676);
nand U3410 (N_3410,N_2721,N_2605);
nor U3411 (N_3411,N_2896,N_2719);
and U3412 (N_3412,N_2817,N_2976);
xor U3413 (N_3413,N_2547,N_2565);
or U3414 (N_3414,N_2630,N_2522);
or U3415 (N_3415,N_2845,N_2574);
xnor U3416 (N_3416,N_2634,N_2937);
and U3417 (N_3417,N_2857,N_2592);
or U3418 (N_3418,N_2813,N_2930);
nand U3419 (N_3419,N_2747,N_2910);
or U3420 (N_3420,N_2504,N_2620);
or U3421 (N_3421,N_2995,N_2776);
or U3422 (N_3422,N_2792,N_2598);
nand U3423 (N_3423,N_2969,N_2828);
nand U3424 (N_3424,N_2701,N_2679);
xnor U3425 (N_3425,N_2533,N_2627);
or U3426 (N_3426,N_2914,N_2663);
nand U3427 (N_3427,N_2758,N_2669);
nor U3428 (N_3428,N_2717,N_2542);
xnor U3429 (N_3429,N_2685,N_2834);
nand U3430 (N_3430,N_2664,N_2545);
xnor U3431 (N_3431,N_2671,N_2879);
nand U3432 (N_3432,N_2848,N_2854);
xor U3433 (N_3433,N_2613,N_2617);
xor U3434 (N_3434,N_2878,N_2720);
nand U3435 (N_3435,N_2565,N_2770);
or U3436 (N_3436,N_2744,N_2837);
nor U3437 (N_3437,N_2531,N_2945);
xnor U3438 (N_3438,N_2736,N_2961);
nand U3439 (N_3439,N_2518,N_2530);
xnor U3440 (N_3440,N_2905,N_2565);
nor U3441 (N_3441,N_2894,N_2512);
nand U3442 (N_3442,N_2886,N_2563);
or U3443 (N_3443,N_2885,N_2645);
xor U3444 (N_3444,N_2758,N_2719);
nor U3445 (N_3445,N_2771,N_2641);
xnor U3446 (N_3446,N_2713,N_2530);
nor U3447 (N_3447,N_2976,N_2927);
nand U3448 (N_3448,N_2582,N_2839);
nor U3449 (N_3449,N_2924,N_2969);
or U3450 (N_3450,N_2979,N_2733);
and U3451 (N_3451,N_2738,N_2778);
nor U3452 (N_3452,N_2891,N_2764);
xnor U3453 (N_3453,N_2995,N_2510);
and U3454 (N_3454,N_2641,N_2617);
or U3455 (N_3455,N_2900,N_2836);
xor U3456 (N_3456,N_2937,N_2614);
or U3457 (N_3457,N_2548,N_2615);
and U3458 (N_3458,N_2831,N_2637);
nor U3459 (N_3459,N_2541,N_2901);
or U3460 (N_3460,N_2677,N_2953);
or U3461 (N_3461,N_2827,N_2806);
or U3462 (N_3462,N_2683,N_2948);
and U3463 (N_3463,N_2640,N_2803);
xnor U3464 (N_3464,N_2847,N_2855);
nand U3465 (N_3465,N_2516,N_2989);
xor U3466 (N_3466,N_2921,N_2649);
and U3467 (N_3467,N_2776,N_2504);
nor U3468 (N_3468,N_2732,N_2560);
nor U3469 (N_3469,N_2599,N_2969);
or U3470 (N_3470,N_2837,N_2778);
nor U3471 (N_3471,N_2987,N_2560);
or U3472 (N_3472,N_2799,N_2984);
xnor U3473 (N_3473,N_2607,N_2818);
and U3474 (N_3474,N_2864,N_2506);
nor U3475 (N_3475,N_2843,N_2870);
xor U3476 (N_3476,N_2714,N_2868);
nand U3477 (N_3477,N_2614,N_2686);
nor U3478 (N_3478,N_2595,N_2959);
nand U3479 (N_3479,N_2734,N_2870);
xnor U3480 (N_3480,N_2899,N_2966);
xor U3481 (N_3481,N_2954,N_2567);
and U3482 (N_3482,N_2816,N_2874);
and U3483 (N_3483,N_2996,N_2664);
xnor U3484 (N_3484,N_2755,N_2551);
nand U3485 (N_3485,N_2842,N_2615);
nand U3486 (N_3486,N_2747,N_2870);
nor U3487 (N_3487,N_2707,N_2947);
xnor U3488 (N_3488,N_2792,N_2778);
or U3489 (N_3489,N_2873,N_2681);
xnor U3490 (N_3490,N_2855,N_2746);
xor U3491 (N_3491,N_2825,N_2801);
and U3492 (N_3492,N_2687,N_2825);
nand U3493 (N_3493,N_2728,N_2699);
xor U3494 (N_3494,N_2833,N_2780);
nand U3495 (N_3495,N_2683,N_2594);
nand U3496 (N_3496,N_2902,N_2852);
and U3497 (N_3497,N_2880,N_2724);
xor U3498 (N_3498,N_2982,N_2691);
or U3499 (N_3499,N_2896,N_2930);
or U3500 (N_3500,N_3345,N_3294);
and U3501 (N_3501,N_3192,N_3271);
nand U3502 (N_3502,N_3057,N_3167);
nor U3503 (N_3503,N_3116,N_3270);
or U3504 (N_3504,N_3257,N_3233);
nand U3505 (N_3505,N_3153,N_3123);
nand U3506 (N_3506,N_3119,N_3203);
nor U3507 (N_3507,N_3364,N_3353);
xor U3508 (N_3508,N_3161,N_3213);
and U3509 (N_3509,N_3019,N_3420);
and U3510 (N_3510,N_3452,N_3384);
nor U3511 (N_3511,N_3075,N_3110);
xnor U3512 (N_3512,N_3306,N_3186);
nand U3513 (N_3513,N_3073,N_3363);
or U3514 (N_3514,N_3050,N_3069);
nor U3515 (N_3515,N_3168,N_3025);
xor U3516 (N_3516,N_3301,N_3284);
xnor U3517 (N_3517,N_3286,N_3037);
nor U3518 (N_3518,N_3296,N_3133);
xor U3519 (N_3519,N_3096,N_3255);
nor U3520 (N_3520,N_3307,N_3425);
nand U3521 (N_3521,N_3132,N_3259);
nand U3522 (N_3522,N_3194,N_3020);
nand U3523 (N_3523,N_3256,N_3409);
or U3524 (N_3524,N_3478,N_3124);
nand U3525 (N_3525,N_3258,N_3042);
nor U3526 (N_3526,N_3154,N_3081);
xor U3527 (N_3527,N_3303,N_3392);
nand U3528 (N_3528,N_3320,N_3144);
nand U3529 (N_3529,N_3369,N_3134);
or U3530 (N_3530,N_3131,N_3018);
xnor U3531 (N_3531,N_3434,N_3224);
nand U3532 (N_3532,N_3054,N_3000);
or U3533 (N_3533,N_3378,N_3190);
nor U3534 (N_3534,N_3059,N_3084);
xor U3535 (N_3535,N_3030,N_3451);
nand U3536 (N_3536,N_3149,N_3055);
nor U3537 (N_3537,N_3298,N_3182);
or U3538 (N_3538,N_3181,N_3129);
or U3539 (N_3539,N_3325,N_3179);
nand U3540 (N_3540,N_3068,N_3048);
or U3541 (N_3541,N_3486,N_3078);
or U3542 (N_3542,N_3022,N_3458);
xnor U3543 (N_3543,N_3099,N_3348);
or U3544 (N_3544,N_3398,N_3397);
and U3545 (N_3545,N_3322,N_3121);
and U3546 (N_3546,N_3017,N_3109);
xor U3547 (N_3547,N_3198,N_3038);
and U3548 (N_3548,N_3231,N_3244);
xnor U3549 (N_3549,N_3360,N_3220);
and U3550 (N_3550,N_3071,N_3074);
nand U3551 (N_3551,N_3235,N_3309);
xor U3552 (N_3552,N_3466,N_3265);
nor U3553 (N_3553,N_3436,N_3379);
or U3554 (N_3554,N_3196,N_3329);
nor U3555 (N_3555,N_3472,N_3261);
and U3556 (N_3556,N_3415,N_3310);
and U3557 (N_3557,N_3305,N_3482);
xnor U3558 (N_3558,N_3498,N_3027);
and U3559 (N_3559,N_3391,N_3247);
and U3560 (N_3560,N_3170,N_3229);
or U3561 (N_3561,N_3063,N_3012);
xor U3562 (N_3562,N_3315,N_3413);
and U3563 (N_3563,N_3439,N_3112);
nand U3564 (N_3564,N_3300,N_3430);
nor U3565 (N_3565,N_3089,N_3135);
nor U3566 (N_3566,N_3281,N_3461);
nand U3567 (N_3567,N_3004,N_3139);
nand U3568 (N_3568,N_3010,N_3032);
or U3569 (N_3569,N_3151,N_3467);
nand U3570 (N_3570,N_3393,N_3240);
xor U3571 (N_3571,N_3023,N_3274);
xor U3572 (N_3572,N_3085,N_3028);
or U3573 (N_3573,N_3263,N_3077);
nor U3574 (N_3574,N_3395,N_3349);
and U3575 (N_3575,N_3404,N_3311);
xnor U3576 (N_3576,N_3444,N_3241);
xnor U3577 (N_3577,N_3491,N_3202);
nand U3578 (N_3578,N_3142,N_3387);
and U3579 (N_3579,N_3282,N_3421);
nor U3580 (N_3580,N_3273,N_3412);
nand U3581 (N_3581,N_3248,N_3001);
xor U3582 (N_3582,N_3172,N_3092);
nor U3583 (N_3583,N_3014,N_3441);
nor U3584 (N_3584,N_3276,N_3357);
or U3585 (N_3585,N_3326,N_3043);
and U3586 (N_3586,N_3480,N_3047);
or U3587 (N_3587,N_3424,N_3386);
nand U3588 (N_3588,N_3489,N_3137);
or U3589 (N_3589,N_3218,N_3100);
or U3590 (N_3590,N_3005,N_3367);
nor U3591 (N_3591,N_3408,N_3332);
and U3592 (N_3592,N_3470,N_3388);
nor U3593 (N_3593,N_3312,N_3150);
or U3594 (N_3594,N_3021,N_3446);
xnor U3595 (N_3595,N_3098,N_3097);
xnor U3596 (N_3596,N_3358,N_3034);
or U3597 (N_3597,N_3374,N_3173);
xnor U3598 (N_3598,N_3447,N_3383);
xnor U3599 (N_3599,N_3013,N_3269);
xor U3600 (N_3600,N_3380,N_3046);
xnor U3601 (N_3601,N_3479,N_3262);
nor U3602 (N_3602,N_3366,N_3403);
or U3603 (N_3603,N_3435,N_3481);
nor U3604 (N_3604,N_3299,N_3477);
nor U3605 (N_3605,N_3108,N_3344);
nand U3606 (N_3606,N_3002,N_3169);
nor U3607 (N_3607,N_3122,N_3476);
and U3608 (N_3608,N_3342,N_3106);
nand U3609 (N_3609,N_3188,N_3015);
nand U3610 (N_3610,N_3459,N_3277);
nand U3611 (N_3611,N_3443,N_3065);
nor U3612 (N_3612,N_3072,N_3471);
xnor U3613 (N_3613,N_3319,N_3211);
nor U3614 (N_3614,N_3234,N_3215);
nor U3615 (N_3615,N_3120,N_3359);
xor U3616 (N_3616,N_3197,N_3204);
and U3617 (N_3617,N_3058,N_3339);
nand U3618 (N_3618,N_3062,N_3102);
or U3619 (N_3619,N_3141,N_3400);
xnor U3620 (N_3620,N_3026,N_3449);
nor U3621 (N_3621,N_3178,N_3343);
and U3622 (N_3622,N_3406,N_3295);
or U3623 (N_3623,N_3183,N_3431);
and U3624 (N_3624,N_3494,N_3440);
or U3625 (N_3625,N_3341,N_3165);
and U3626 (N_3626,N_3289,N_3061);
nor U3627 (N_3627,N_3193,N_3066);
or U3628 (N_3628,N_3352,N_3340);
nand U3629 (N_3629,N_3464,N_3304);
xnor U3630 (N_3630,N_3225,N_3175);
nand U3631 (N_3631,N_3394,N_3487);
xnor U3632 (N_3632,N_3496,N_3492);
nor U3633 (N_3633,N_3128,N_3331);
nor U3634 (N_3634,N_3221,N_3242);
and U3635 (N_3635,N_3474,N_3127);
nor U3636 (N_3636,N_3199,N_3082);
xor U3637 (N_3637,N_3138,N_3375);
xnor U3638 (N_3638,N_3278,N_3254);
nand U3639 (N_3639,N_3070,N_3442);
nand U3640 (N_3640,N_3101,N_3105);
nor U3641 (N_3641,N_3365,N_3453);
and U3642 (N_3642,N_3302,N_3488);
nor U3643 (N_3643,N_3445,N_3158);
and U3644 (N_3644,N_3493,N_3485);
xor U3645 (N_3645,N_3402,N_3268);
xor U3646 (N_3646,N_3163,N_3171);
xnor U3647 (N_3647,N_3407,N_3428);
xor U3648 (N_3648,N_3356,N_3285);
nor U3649 (N_3649,N_3328,N_3297);
nand U3650 (N_3650,N_3126,N_3118);
xor U3651 (N_3651,N_3260,N_3174);
or U3652 (N_3652,N_3450,N_3107);
xnor U3653 (N_3653,N_3433,N_3468);
xnor U3654 (N_3654,N_3080,N_3040);
nor U3655 (N_3655,N_3318,N_3228);
xnor U3656 (N_3656,N_3361,N_3483);
xnor U3657 (N_3657,N_3064,N_3465);
nor U3658 (N_3658,N_3246,N_3288);
and U3659 (N_3659,N_3189,N_3418);
nor U3660 (N_3660,N_3009,N_3016);
xnor U3661 (N_3661,N_3238,N_3390);
xnor U3662 (N_3662,N_3456,N_3094);
nand U3663 (N_3663,N_3372,N_3226);
or U3664 (N_3664,N_3239,N_3206);
nand U3665 (N_3665,N_3399,N_3429);
nor U3666 (N_3666,N_3460,N_3083);
nor U3667 (N_3667,N_3152,N_3024);
nor U3668 (N_3668,N_3267,N_3370);
xnor U3669 (N_3669,N_3416,N_3051);
xor U3670 (N_3670,N_3346,N_3423);
xor U3671 (N_3671,N_3011,N_3266);
nand U3672 (N_3672,N_3053,N_3114);
and U3673 (N_3673,N_3113,N_3373);
nor U3674 (N_3674,N_3362,N_3007);
nor U3675 (N_3675,N_3437,N_3347);
nor U3676 (N_3676,N_3499,N_3210);
xnor U3677 (N_3677,N_3338,N_3003);
nor U3678 (N_3678,N_3475,N_3287);
nand U3679 (N_3679,N_3103,N_3448);
nand U3680 (N_3680,N_3157,N_3291);
nor U3681 (N_3681,N_3350,N_3250);
xnor U3682 (N_3682,N_3243,N_3264);
nor U3683 (N_3683,N_3462,N_3405);
nand U3684 (N_3684,N_3045,N_3130);
or U3685 (N_3685,N_3164,N_3272);
or U3686 (N_3686,N_3316,N_3187);
xor U3687 (N_3687,N_3232,N_3006);
or U3688 (N_3688,N_3185,N_3280);
and U3689 (N_3689,N_3279,N_3200);
nand U3690 (N_3690,N_3290,N_3292);
nor U3691 (N_3691,N_3090,N_3455);
nor U3692 (N_3692,N_3136,N_3029);
nor U3693 (N_3693,N_3463,N_3432);
and U3694 (N_3694,N_3209,N_3438);
or U3695 (N_3695,N_3457,N_3252);
nor U3696 (N_3696,N_3036,N_3079);
nand U3697 (N_3697,N_3166,N_3214);
and U3698 (N_3698,N_3396,N_3039);
nand U3699 (N_3699,N_3159,N_3410);
nor U3700 (N_3700,N_3208,N_3067);
nor U3701 (N_3701,N_3368,N_3143);
or U3702 (N_3702,N_3327,N_3293);
and U3703 (N_3703,N_3355,N_3056);
nand U3704 (N_3704,N_3217,N_3230);
nand U3705 (N_3705,N_3376,N_3146);
or U3706 (N_3706,N_3381,N_3411);
and U3707 (N_3707,N_3495,N_3314);
or U3708 (N_3708,N_3354,N_3180);
and U3709 (N_3709,N_3095,N_3205);
nand U3710 (N_3710,N_3115,N_3401);
xor U3711 (N_3711,N_3426,N_3351);
and U3712 (N_3712,N_3049,N_3333);
nor U3713 (N_3713,N_3052,N_3145);
and U3714 (N_3714,N_3207,N_3033);
or U3715 (N_3715,N_3086,N_3321);
or U3716 (N_3716,N_3160,N_3087);
xor U3717 (N_3717,N_3148,N_3176);
or U3718 (N_3718,N_3125,N_3162);
xnor U3719 (N_3719,N_3473,N_3385);
and U3720 (N_3720,N_3323,N_3336);
nand U3721 (N_3721,N_3245,N_3382);
nand U3722 (N_3722,N_3147,N_3111);
xnor U3723 (N_3723,N_3223,N_3035);
xor U3724 (N_3724,N_3184,N_3117);
and U3725 (N_3725,N_3031,N_3104);
xnor U3726 (N_3726,N_3156,N_3497);
and U3727 (N_3727,N_3155,N_3371);
or U3728 (N_3728,N_3041,N_3417);
or U3729 (N_3729,N_3283,N_3195);
nor U3730 (N_3730,N_3236,N_3330);
nor U3731 (N_3731,N_3222,N_3337);
xnor U3732 (N_3732,N_3140,N_3076);
nand U3733 (N_3733,N_3313,N_3454);
nor U3734 (N_3734,N_3044,N_3253);
nand U3735 (N_3735,N_3490,N_3484);
and U3736 (N_3736,N_3275,N_3469);
nor U3737 (N_3737,N_3191,N_3317);
or U3738 (N_3738,N_3308,N_3249);
or U3739 (N_3739,N_3060,N_3389);
nand U3740 (N_3740,N_3219,N_3414);
nor U3741 (N_3741,N_3177,N_3008);
nand U3742 (N_3742,N_3237,N_3422);
and U3743 (N_3743,N_3093,N_3216);
nand U3744 (N_3744,N_3377,N_3227);
nand U3745 (N_3745,N_3427,N_3212);
nand U3746 (N_3746,N_3251,N_3324);
nand U3747 (N_3747,N_3091,N_3334);
nor U3748 (N_3748,N_3419,N_3201);
nor U3749 (N_3749,N_3088,N_3335);
nor U3750 (N_3750,N_3275,N_3313);
nand U3751 (N_3751,N_3318,N_3389);
xor U3752 (N_3752,N_3286,N_3130);
xnor U3753 (N_3753,N_3148,N_3336);
or U3754 (N_3754,N_3280,N_3397);
nor U3755 (N_3755,N_3133,N_3025);
and U3756 (N_3756,N_3352,N_3358);
nand U3757 (N_3757,N_3301,N_3250);
and U3758 (N_3758,N_3318,N_3191);
xnor U3759 (N_3759,N_3060,N_3453);
nand U3760 (N_3760,N_3447,N_3072);
xor U3761 (N_3761,N_3034,N_3320);
nand U3762 (N_3762,N_3370,N_3376);
xor U3763 (N_3763,N_3045,N_3400);
nor U3764 (N_3764,N_3003,N_3408);
xnor U3765 (N_3765,N_3322,N_3204);
or U3766 (N_3766,N_3288,N_3268);
nor U3767 (N_3767,N_3049,N_3079);
nand U3768 (N_3768,N_3381,N_3469);
nor U3769 (N_3769,N_3027,N_3228);
or U3770 (N_3770,N_3333,N_3497);
xnor U3771 (N_3771,N_3139,N_3358);
or U3772 (N_3772,N_3268,N_3289);
nand U3773 (N_3773,N_3160,N_3449);
nand U3774 (N_3774,N_3111,N_3215);
and U3775 (N_3775,N_3480,N_3372);
or U3776 (N_3776,N_3150,N_3241);
nand U3777 (N_3777,N_3036,N_3264);
and U3778 (N_3778,N_3036,N_3177);
nor U3779 (N_3779,N_3052,N_3125);
nor U3780 (N_3780,N_3347,N_3113);
nor U3781 (N_3781,N_3162,N_3384);
nand U3782 (N_3782,N_3308,N_3059);
xnor U3783 (N_3783,N_3221,N_3453);
nor U3784 (N_3784,N_3417,N_3395);
nand U3785 (N_3785,N_3280,N_3490);
and U3786 (N_3786,N_3227,N_3043);
xor U3787 (N_3787,N_3486,N_3438);
or U3788 (N_3788,N_3370,N_3232);
xor U3789 (N_3789,N_3246,N_3027);
or U3790 (N_3790,N_3366,N_3396);
or U3791 (N_3791,N_3085,N_3451);
xnor U3792 (N_3792,N_3044,N_3108);
and U3793 (N_3793,N_3154,N_3479);
and U3794 (N_3794,N_3363,N_3465);
nand U3795 (N_3795,N_3401,N_3323);
xnor U3796 (N_3796,N_3402,N_3003);
xnor U3797 (N_3797,N_3371,N_3440);
and U3798 (N_3798,N_3235,N_3371);
or U3799 (N_3799,N_3320,N_3139);
or U3800 (N_3800,N_3112,N_3238);
or U3801 (N_3801,N_3351,N_3455);
nor U3802 (N_3802,N_3240,N_3461);
nand U3803 (N_3803,N_3013,N_3471);
nor U3804 (N_3804,N_3405,N_3491);
xor U3805 (N_3805,N_3440,N_3157);
nand U3806 (N_3806,N_3454,N_3451);
xor U3807 (N_3807,N_3425,N_3308);
and U3808 (N_3808,N_3466,N_3418);
nand U3809 (N_3809,N_3448,N_3203);
nor U3810 (N_3810,N_3043,N_3098);
nor U3811 (N_3811,N_3379,N_3499);
and U3812 (N_3812,N_3481,N_3127);
and U3813 (N_3813,N_3322,N_3118);
nand U3814 (N_3814,N_3354,N_3041);
nor U3815 (N_3815,N_3386,N_3082);
xor U3816 (N_3816,N_3036,N_3498);
xor U3817 (N_3817,N_3403,N_3493);
nand U3818 (N_3818,N_3005,N_3400);
nor U3819 (N_3819,N_3401,N_3164);
and U3820 (N_3820,N_3048,N_3385);
nand U3821 (N_3821,N_3048,N_3107);
nand U3822 (N_3822,N_3088,N_3113);
nor U3823 (N_3823,N_3281,N_3106);
or U3824 (N_3824,N_3342,N_3371);
xor U3825 (N_3825,N_3170,N_3418);
or U3826 (N_3826,N_3096,N_3193);
nand U3827 (N_3827,N_3345,N_3437);
nor U3828 (N_3828,N_3332,N_3483);
nand U3829 (N_3829,N_3339,N_3372);
and U3830 (N_3830,N_3345,N_3149);
nand U3831 (N_3831,N_3484,N_3261);
nand U3832 (N_3832,N_3144,N_3377);
nand U3833 (N_3833,N_3118,N_3250);
or U3834 (N_3834,N_3445,N_3497);
nor U3835 (N_3835,N_3200,N_3459);
nor U3836 (N_3836,N_3050,N_3181);
or U3837 (N_3837,N_3272,N_3056);
nand U3838 (N_3838,N_3166,N_3414);
nor U3839 (N_3839,N_3449,N_3218);
or U3840 (N_3840,N_3433,N_3300);
nor U3841 (N_3841,N_3427,N_3418);
nor U3842 (N_3842,N_3104,N_3034);
xor U3843 (N_3843,N_3098,N_3012);
xor U3844 (N_3844,N_3114,N_3287);
xor U3845 (N_3845,N_3051,N_3166);
nor U3846 (N_3846,N_3424,N_3116);
nor U3847 (N_3847,N_3048,N_3033);
or U3848 (N_3848,N_3326,N_3465);
and U3849 (N_3849,N_3361,N_3342);
nand U3850 (N_3850,N_3285,N_3450);
or U3851 (N_3851,N_3175,N_3061);
nand U3852 (N_3852,N_3064,N_3248);
xor U3853 (N_3853,N_3325,N_3453);
xor U3854 (N_3854,N_3043,N_3261);
nor U3855 (N_3855,N_3036,N_3361);
nor U3856 (N_3856,N_3362,N_3245);
nand U3857 (N_3857,N_3294,N_3484);
xor U3858 (N_3858,N_3285,N_3459);
nand U3859 (N_3859,N_3083,N_3001);
nor U3860 (N_3860,N_3254,N_3461);
xor U3861 (N_3861,N_3340,N_3251);
or U3862 (N_3862,N_3495,N_3280);
and U3863 (N_3863,N_3254,N_3486);
xnor U3864 (N_3864,N_3011,N_3432);
and U3865 (N_3865,N_3464,N_3377);
nor U3866 (N_3866,N_3240,N_3028);
nand U3867 (N_3867,N_3058,N_3175);
or U3868 (N_3868,N_3360,N_3218);
or U3869 (N_3869,N_3081,N_3317);
nor U3870 (N_3870,N_3092,N_3461);
nor U3871 (N_3871,N_3140,N_3083);
xor U3872 (N_3872,N_3172,N_3110);
nand U3873 (N_3873,N_3221,N_3052);
xor U3874 (N_3874,N_3001,N_3410);
or U3875 (N_3875,N_3168,N_3154);
nor U3876 (N_3876,N_3007,N_3355);
nand U3877 (N_3877,N_3183,N_3413);
or U3878 (N_3878,N_3059,N_3394);
or U3879 (N_3879,N_3134,N_3276);
nor U3880 (N_3880,N_3330,N_3427);
nor U3881 (N_3881,N_3077,N_3034);
xor U3882 (N_3882,N_3107,N_3473);
xnor U3883 (N_3883,N_3311,N_3153);
nand U3884 (N_3884,N_3060,N_3486);
xor U3885 (N_3885,N_3433,N_3034);
nand U3886 (N_3886,N_3167,N_3451);
and U3887 (N_3887,N_3464,N_3347);
or U3888 (N_3888,N_3436,N_3437);
and U3889 (N_3889,N_3344,N_3383);
nand U3890 (N_3890,N_3347,N_3207);
and U3891 (N_3891,N_3415,N_3089);
and U3892 (N_3892,N_3145,N_3362);
nand U3893 (N_3893,N_3064,N_3240);
xnor U3894 (N_3894,N_3051,N_3095);
or U3895 (N_3895,N_3498,N_3348);
nor U3896 (N_3896,N_3192,N_3203);
nor U3897 (N_3897,N_3214,N_3303);
xnor U3898 (N_3898,N_3440,N_3081);
nand U3899 (N_3899,N_3101,N_3459);
and U3900 (N_3900,N_3023,N_3036);
nand U3901 (N_3901,N_3365,N_3413);
nor U3902 (N_3902,N_3434,N_3179);
or U3903 (N_3903,N_3254,N_3040);
xnor U3904 (N_3904,N_3054,N_3432);
and U3905 (N_3905,N_3248,N_3014);
nor U3906 (N_3906,N_3400,N_3013);
nand U3907 (N_3907,N_3418,N_3143);
nor U3908 (N_3908,N_3409,N_3264);
nor U3909 (N_3909,N_3148,N_3028);
or U3910 (N_3910,N_3359,N_3414);
and U3911 (N_3911,N_3181,N_3440);
or U3912 (N_3912,N_3301,N_3210);
xor U3913 (N_3913,N_3304,N_3254);
nor U3914 (N_3914,N_3322,N_3403);
and U3915 (N_3915,N_3049,N_3196);
nor U3916 (N_3916,N_3430,N_3487);
nand U3917 (N_3917,N_3022,N_3330);
nand U3918 (N_3918,N_3200,N_3495);
and U3919 (N_3919,N_3218,N_3190);
or U3920 (N_3920,N_3012,N_3336);
or U3921 (N_3921,N_3324,N_3286);
nor U3922 (N_3922,N_3197,N_3433);
nand U3923 (N_3923,N_3406,N_3418);
or U3924 (N_3924,N_3103,N_3285);
xor U3925 (N_3925,N_3378,N_3146);
or U3926 (N_3926,N_3220,N_3344);
or U3927 (N_3927,N_3432,N_3395);
nor U3928 (N_3928,N_3036,N_3324);
nor U3929 (N_3929,N_3045,N_3192);
nand U3930 (N_3930,N_3281,N_3248);
and U3931 (N_3931,N_3485,N_3236);
xor U3932 (N_3932,N_3352,N_3311);
xor U3933 (N_3933,N_3376,N_3030);
nor U3934 (N_3934,N_3182,N_3377);
nor U3935 (N_3935,N_3109,N_3421);
nand U3936 (N_3936,N_3415,N_3164);
xnor U3937 (N_3937,N_3017,N_3191);
xnor U3938 (N_3938,N_3238,N_3466);
and U3939 (N_3939,N_3059,N_3071);
nand U3940 (N_3940,N_3321,N_3474);
nand U3941 (N_3941,N_3275,N_3149);
nand U3942 (N_3942,N_3050,N_3422);
or U3943 (N_3943,N_3354,N_3305);
nand U3944 (N_3944,N_3346,N_3392);
and U3945 (N_3945,N_3341,N_3159);
nand U3946 (N_3946,N_3190,N_3088);
nor U3947 (N_3947,N_3060,N_3459);
or U3948 (N_3948,N_3270,N_3275);
and U3949 (N_3949,N_3323,N_3236);
or U3950 (N_3950,N_3391,N_3287);
nand U3951 (N_3951,N_3283,N_3464);
nand U3952 (N_3952,N_3265,N_3390);
nand U3953 (N_3953,N_3085,N_3373);
or U3954 (N_3954,N_3004,N_3220);
and U3955 (N_3955,N_3238,N_3355);
nand U3956 (N_3956,N_3356,N_3390);
and U3957 (N_3957,N_3313,N_3200);
xnor U3958 (N_3958,N_3488,N_3295);
nand U3959 (N_3959,N_3274,N_3149);
nor U3960 (N_3960,N_3490,N_3203);
or U3961 (N_3961,N_3255,N_3133);
and U3962 (N_3962,N_3486,N_3262);
xnor U3963 (N_3963,N_3252,N_3020);
xor U3964 (N_3964,N_3013,N_3460);
or U3965 (N_3965,N_3244,N_3180);
nand U3966 (N_3966,N_3440,N_3191);
nand U3967 (N_3967,N_3088,N_3101);
nand U3968 (N_3968,N_3260,N_3438);
nand U3969 (N_3969,N_3395,N_3285);
xnor U3970 (N_3970,N_3287,N_3260);
xor U3971 (N_3971,N_3063,N_3144);
nor U3972 (N_3972,N_3123,N_3027);
or U3973 (N_3973,N_3160,N_3059);
or U3974 (N_3974,N_3438,N_3073);
xor U3975 (N_3975,N_3266,N_3079);
nor U3976 (N_3976,N_3136,N_3344);
and U3977 (N_3977,N_3491,N_3232);
nand U3978 (N_3978,N_3448,N_3464);
nand U3979 (N_3979,N_3082,N_3282);
and U3980 (N_3980,N_3051,N_3074);
or U3981 (N_3981,N_3152,N_3420);
xor U3982 (N_3982,N_3475,N_3298);
or U3983 (N_3983,N_3269,N_3039);
and U3984 (N_3984,N_3122,N_3302);
xor U3985 (N_3985,N_3235,N_3427);
and U3986 (N_3986,N_3452,N_3304);
nor U3987 (N_3987,N_3301,N_3161);
and U3988 (N_3988,N_3331,N_3103);
xnor U3989 (N_3989,N_3056,N_3333);
nand U3990 (N_3990,N_3462,N_3477);
nand U3991 (N_3991,N_3030,N_3164);
nand U3992 (N_3992,N_3392,N_3070);
and U3993 (N_3993,N_3226,N_3196);
xnor U3994 (N_3994,N_3051,N_3408);
xor U3995 (N_3995,N_3327,N_3404);
and U3996 (N_3996,N_3169,N_3370);
nand U3997 (N_3997,N_3245,N_3422);
xor U3998 (N_3998,N_3366,N_3498);
or U3999 (N_3999,N_3277,N_3292);
nand U4000 (N_4000,N_3706,N_3969);
or U4001 (N_4001,N_3644,N_3749);
nand U4002 (N_4002,N_3899,N_3808);
or U4003 (N_4003,N_3850,N_3782);
and U4004 (N_4004,N_3713,N_3837);
and U4005 (N_4005,N_3809,N_3839);
or U4006 (N_4006,N_3633,N_3638);
nor U4007 (N_4007,N_3885,N_3589);
xor U4008 (N_4008,N_3760,N_3692);
xnor U4009 (N_4009,N_3852,N_3928);
nor U4010 (N_4010,N_3676,N_3798);
nor U4011 (N_4011,N_3636,N_3912);
and U4012 (N_4012,N_3959,N_3549);
and U4013 (N_4013,N_3983,N_3653);
nand U4014 (N_4014,N_3904,N_3550);
nor U4015 (N_4015,N_3687,N_3649);
nor U4016 (N_4016,N_3855,N_3891);
or U4017 (N_4017,N_3859,N_3673);
nor U4018 (N_4018,N_3631,N_3998);
and U4019 (N_4019,N_3917,N_3829);
or U4020 (N_4020,N_3571,N_3920);
nand U4021 (N_4021,N_3783,N_3866);
nand U4022 (N_4022,N_3725,N_3514);
xnor U4023 (N_4023,N_3854,N_3659);
xnor U4024 (N_4024,N_3896,N_3547);
nor U4025 (N_4025,N_3967,N_3728);
xor U4026 (N_4026,N_3968,N_3535);
nand U4027 (N_4027,N_3627,N_3824);
and U4028 (N_4028,N_3606,N_3624);
and U4029 (N_4029,N_3868,N_3874);
or U4030 (N_4030,N_3978,N_3847);
nor U4031 (N_4031,N_3851,N_3913);
or U4032 (N_4032,N_3595,N_3751);
or U4033 (N_4033,N_3816,N_3518);
nor U4034 (N_4034,N_3776,N_3774);
or U4035 (N_4035,N_3598,N_3599);
nand U4036 (N_4036,N_3614,N_3916);
nor U4037 (N_4037,N_3629,N_3648);
xnor U4038 (N_4038,N_3656,N_3863);
and U4039 (N_4039,N_3758,N_3545);
xor U4040 (N_4040,N_3694,N_3801);
nor U4041 (N_4041,N_3792,N_3901);
nor U4042 (N_4042,N_3775,N_3722);
or U4043 (N_4043,N_3554,N_3597);
xnor U4044 (N_4044,N_3752,N_3528);
nand U4045 (N_4045,N_3761,N_3743);
or U4046 (N_4046,N_3861,N_3738);
nand U4047 (N_4047,N_3922,N_3587);
and U4048 (N_4048,N_3684,N_3759);
or U4049 (N_4049,N_3812,N_3583);
xor U4050 (N_4050,N_3556,N_3870);
or U4051 (N_4051,N_3696,N_3892);
or U4052 (N_4052,N_3811,N_3778);
or U4053 (N_4053,N_3947,N_3875);
and U4054 (N_4054,N_3736,N_3585);
or U4055 (N_4055,N_3590,N_3621);
and U4056 (N_4056,N_3560,N_3652);
nor U4057 (N_4057,N_3832,N_3960);
or U4058 (N_4058,N_3680,N_3574);
xor U4059 (N_4059,N_3612,N_3937);
nand U4060 (N_4060,N_3537,N_3867);
or U4061 (N_4061,N_3933,N_3754);
nand U4062 (N_4062,N_3948,N_3987);
nand U4063 (N_4063,N_3577,N_3508);
nand U4064 (N_4064,N_3755,N_3575);
nand U4065 (N_4065,N_3640,N_3646);
nand U4066 (N_4066,N_3525,N_3690);
and U4067 (N_4067,N_3827,N_3720);
nor U4068 (N_4068,N_3503,N_3910);
nor U4069 (N_4069,N_3512,N_3784);
xor U4070 (N_4070,N_3876,N_3552);
nand U4071 (N_4071,N_3989,N_3982);
or U4072 (N_4072,N_3600,N_3840);
xnor U4073 (N_4073,N_3893,N_3538);
nand U4074 (N_4074,N_3958,N_3767);
xor U4075 (N_4075,N_3580,N_3918);
nor U4076 (N_4076,N_3777,N_3838);
nor U4077 (N_4077,N_3693,N_3833);
xor U4078 (N_4078,N_3756,N_3935);
xnor U4079 (N_4079,N_3591,N_3900);
xor U4080 (N_4080,N_3848,N_3679);
xor U4081 (N_4081,N_3524,N_3733);
and U4082 (N_4082,N_3592,N_3611);
xor U4083 (N_4083,N_3729,N_3831);
or U4084 (N_4084,N_3880,N_3740);
xnor U4085 (N_4085,N_3769,N_3651);
nand U4086 (N_4086,N_3544,N_3879);
nor U4087 (N_4087,N_3864,N_3791);
nor U4088 (N_4088,N_3632,N_3963);
xnor U4089 (N_4089,N_3762,N_3539);
nand U4090 (N_4090,N_3888,N_3543);
xor U4091 (N_4091,N_3586,N_3582);
xnor U4092 (N_4092,N_3845,N_3797);
or U4093 (N_4093,N_3700,N_3945);
and U4094 (N_4094,N_3844,N_3976);
or U4095 (N_4095,N_3953,N_3559);
nand U4096 (N_4096,N_3691,N_3618);
or U4097 (N_4097,N_3857,N_3594);
and U4098 (N_4098,N_3871,N_3952);
and U4099 (N_4099,N_3584,N_3787);
nand U4100 (N_4100,N_3942,N_3794);
xor U4101 (N_4101,N_3887,N_3502);
nand U4102 (N_4102,N_3788,N_3661);
xnor U4103 (N_4103,N_3807,N_3746);
nand U4104 (N_4104,N_3737,N_3789);
or U4105 (N_4105,N_3869,N_3919);
nand U4106 (N_4106,N_3639,N_3623);
or U4107 (N_4107,N_3735,N_3997);
and U4108 (N_4108,N_3793,N_3664);
nor U4109 (N_4109,N_3682,N_3955);
nor U4110 (N_4110,N_3883,N_3609);
or U4111 (N_4111,N_3710,N_3516);
or U4112 (N_4112,N_3634,N_3936);
xnor U4113 (N_4113,N_3826,N_3872);
or U4114 (N_4114,N_3568,N_3620);
or U4115 (N_4115,N_3924,N_3841);
nand U4116 (N_4116,N_3810,N_3671);
nor U4117 (N_4117,N_3701,N_3939);
nor U4118 (N_4118,N_3662,N_3938);
nor U4119 (N_4119,N_3772,N_3815);
xor U4120 (N_4120,N_3677,N_3695);
nor U4121 (N_4121,N_3655,N_3820);
or U4122 (N_4122,N_3727,N_3742);
nand U4123 (N_4123,N_3994,N_3570);
or U4124 (N_4124,N_3697,N_3941);
nand U4125 (N_4125,N_3660,N_3940);
nand U4126 (N_4126,N_3925,N_3688);
nor U4127 (N_4127,N_3548,N_3576);
xor U4128 (N_4128,N_3748,N_3800);
nand U4129 (N_4129,N_3519,N_3532);
and U4130 (N_4130,N_3821,N_3814);
and U4131 (N_4131,N_3711,N_3921);
and U4132 (N_4132,N_3526,N_3579);
and U4133 (N_4133,N_3732,N_3616);
nor U4134 (N_4134,N_3895,N_3929);
or U4135 (N_4135,N_3522,N_3617);
nand U4136 (N_4136,N_3906,N_3714);
nand U4137 (N_4137,N_3555,N_3961);
nand U4138 (N_4138,N_3730,N_3951);
or U4139 (N_4139,N_3530,N_3860);
nand U4140 (N_4140,N_3846,N_3641);
nor U4141 (N_4141,N_3603,N_3683);
nand U4142 (N_4142,N_3724,N_3505);
nor U4143 (N_4143,N_3593,N_3964);
or U4144 (N_4144,N_3796,N_3670);
xnor U4145 (N_4145,N_3932,N_3509);
and U4146 (N_4146,N_3914,N_3643);
and U4147 (N_4147,N_3965,N_3581);
or U4148 (N_4148,N_3934,N_3506);
nand U4149 (N_4149,N_3569,N_3578);
nand U4150 (N_4150,N_3842,N_3540);
nor U4151 (N_4151,N_3836,N_3799);
xnor U4152 (N_4152,N_3993,N_3977);
and U4153 (N_4153,N_3626,N_3523);
nor U4154 (N_4154,N_3830,N_3985);
nand U4155 (N_4155,N_3944,N_3981);
nand U4156 (N_4156,N_3889,N_3622);
and U4157 (N_4157,N_3897,N_3658);
nand U4158 (N_4158,N_3877,N_3672);
nand U4159 (N_4159,N_3562,N_3986);
and U4160 (N_4160,N_3962,N_3898);
xor U4161 (N_4161,N_3956,N_3678);
xor U4162 (N_4162,N_3739,N_3610);
nor U4163 (N_4163,N_3957,N_3613);
nor U4164 (N_4164,N_3843,N_3699);
or U4165 (N_4165,N_3647,N_3802);
xnor U4166 (N_4166,N_3665,N_3763);
or U4167 (N_4167,N_3780,N_3753);
and U4168 (N_4168,N_3685,N_3795);
xnor U4169 (N_4169,N_3650,N_3865);
nor U4170 (N_4170,N_3645,N_3573);
nand U4171 (N_4171,N_3954,N_3984);
xnor U4172 (N_4172,N_3943,N_3970);
xor U4173 (N_4173,N_3990,N_3950);
nor U4174 (N_4174,N_3856,N_3806);
xor U4175 (N_4175,N_3533,N_3663);
nor U4176 (N_4176,N_3931,N_3566);
nand U4177 (N_4177,N_3534,N_3723);
or U4178 (N_4178,N_3745,N_3757);
xnor U4179 (N_4179,N_3625,N_3628);
xor U4180 (N_4180,N_3501,N_3803);
and U4181 (N_4181,N_3601,N_3907);
or U4182 (N_4182,N_3712,N_3517);
xor U4183 (N_4183,N_3615,N_3828);
and U4184 (N_4184,N_3719,N_3681);
or U4185 (N_4185,N_3909,N_3911);
nand U4186 (N_4186,N_3619,N_3510);
or U4187 (N_4187,N_3973,N_3642);
and U4188 (N_4188,N_3786,N_3930);
and U4189 (N_4189,N_3708,N_3557);
nand U4190 (N_4190,N_3873,N_3882);
or U4191 (N_4191,N_3520,N_3630);
and U4192 (N_4192,N_3657,N_3823);
or U4193 (N_4193,N_3886,N_3511);
nor U4194 (N_4194,N_3884,N_3988);
or U4195 (N_4195,N_3602,N_3707);
and U4196 (N_4196,N_3654,N_3513);
or U4197 (N_4197,N_3507,N_3531);
nor U4198 (N_4198,N_3995,N_3521);
nand U4199 (N_4199,N_3702,N_3608);
or U4200 (N_4200,N_3881,N_3734);
nand U4201 (N_4201,N_3596,N_3668);
nand U4202 (N_4202,N_3771,N_3561);
xor U4203 (N_4203,N_3768,N_3890);
nand U4204 (N_4204,N_3858,N_3817);
xor U4205 (N_4205,N_3605,N_3996);
xor U4206 (N_4206,N_3980,N_3975);
or U4207 (N_4207,N_3546,N_3527);
nor U4208 (N_4208,N_3849,N_3804);
nor U4209 (N_4209,N_3779,N_3781);
xor U4210 (N_4210,N_3604,N_3731);
or U4211 (N_4211,N_3718,N_3805);
nand U4212 (N_4212,N_3716,N_3529);
nand U4213 (N_4213,N_3974,N_3721);
or U4214 (N_4214,N_3834,N_3819);
nor U4215 (N_4215,N_3741,N_3542);
xnor U4216 (N_4216,N_3926,N_3766);
xnor U4217 (N_4217,N_3750,N_3709);
or U4218 (N_4218,N_3705,N_3607);
nand U4219 (N_4219,N_3905,N_3903);
or U4220 (N_4220,N_3500,N_3747);
xor U4221 (N_4221,N_3785,N_3674);
nor U4222 (N_4222,N_3635,N_3862);
nand U4223 (N_4223,N_3991,N_3698);
xor U4224 (N_4224,N_3992,N_3553);
nor U4225 (N_4225,N_3588,N_3558);
or U4226 (N_4226,N_3946,N_3669);
nand U4227 (N_4227,N_3666,N_3703);
or U4228 (N_4228,N_3790,N_3563);
and U4229 (N_4229,N_3744,N_3894);
nand U4230 (N_4230,N_3822,N_3726);
nand U4231 (N_4231,N_3504,N_3835);
nor U4232 (N_4232,N_3764,N_3818);
xor U4233 (N_4233,N_3966,N_3923);
or U4234 (N_4234,N_3878,N_3515);
nor U4235 (N_4235,N_3541,N_3717);
nor U4236 (N_4236,N_3686,N_3572);
nand U4237 (N_4237,N_3825,N_3770);
and U4238 (N_4238,N_3567,N_3949);
nor U4239 (N_4239,N_3773,N_3564);
nand U4240 (N_4240,N_3972,N_3853);
nand U4241 (N_4241,N_3999,N_3689);
and U4242 (N_4242,N_3715,N_3637);
nand U4243 (N_4243,N_3927,N_3551);
or U4244 (N_4244,N_3675,N_3667);
and U4245 (N_4245,N_3971,N_3915);
or U4246 (N_4246,N_3979,N_3565);
nor U4247 (N_4247,N_3902,N_3813);
or U4248 (N_4248,N_3765,N_3908);
nand U4249 (N_4249,N_3536,N_3704);
nor U4250 (N_4250,N_3542,N_3851);
and U4251 (N_4251,N_3864,N_3676);
or U4252 (N_4252,N_3778,N_3559);
nand U4253 (N_4253,N_3826,N_3960);
nor U4254 (N_4254,N_3832,N_3602);
nand U4255 (N_4255,N_3983,N_3979);
or U4256 (N_4256,N_3824,N_3645);
and U4257 (N_4257,N_3579,N_3916);
xnor U4258 (N_4258,N_3748,N_3847);
nand U4259 (N_4259,N_3726,N_3977);
nand U4260 (N_4260,N_3598,N_3972);
and U4261 (N_4261,N_3885,N_3785);
xor U4262 (N_4262,N_3909,N_3516);
nor U4263 (N_4263,N_3647,N_3925);
or U4264 (N_4264,N_3905,N_3521);
nand U4265 (N_4265,N_3618,N_3967);
nor U4266 (N_4266,N_3556,N_3638);
or U4267 (N_4267,N_3595,N_3628);
or U4268 (N_4268,N_3554,N_3785);
nor U4269 (N_4269,N_3545,N_3630);
and U4270 (N_4270,N_3868,N_3680);
or U4271 (N_4271,N_3924,N_3797);
nor U4272 (N_4272,N_3721,N_3796);
nand U4273 (N_4273,N_3718,N_3955);
nor U4274 (N_4274,N_3844,N_3878);
nor U4275 (N_4275,N_3725,N_3774);
nor U4276 (N_4276,N_3835,N_3967);
nand U4277 (N_4277,N_3861,N_3826);
and U4278 (N_4278,N_3555,N_3964);
nand U4279 (N_4279,N_3520,N_3656);
nand U4280 (N_4280,N_3912,N_3547);
and U4281 (N_4281,N_3917,N_3753);
and U4282 (N_4282,N_3872,N_3619);
xor U4283 (N_4283,N_3959,N_3533);
and U4284 (N_4284,N_3621,N_3671);
and U4285 (N_4285,N_3627,N_3571);
nor U4286 (N_4286,N_3567,N_3897);
xor U4287 (N_4287,N_3839,N_3532);
xnor U4288 (N_4288,N_3932,N_3704);
and U4289 (N_4289,N_3777,N_3790);
xor U4290 (N_4290,N_3540,N_3983);
and U4291 (N_4291,N_3956,N_3623);
or U4292 (N_4292,N_3598,N_3554);
xnor U4293 (N_4293,N_3607,N_3602);
nand U4294 (N_4294,N_3832,N_3692);
and U4295 (N_4295,N_3692,N_3666);
and U4296 (N_4296,N_3958,N_3862);
nand U4297 (N_4297,N_3749,N_3888);
nor U4298 (N_4298,N_3792,N_3929);
xor U4299 (N_4299,N_3691,N_3534);
xnor U4300 (N_4300,N_3610,N_3678);
nand U4301 (N_4301,N_3888,N_3751);
nand U4302 (N_4302,N_3840,N_3842);
and U4303 (N_4303,N_3967,N_3739);
and U4304 (N_4304,N_3524,N_3566);
nand U4305 (N_4305,N_3787,N_3747);
and U4306 (N_4306,N_3734,N_3694);
or U4307 (N_4307,N_3577,N_3925);
nand U4308 (N_4308,N_3633,N_3556);
nand U4309 (N_4309,N_3900,N_3604);
xnor U4310 (N_4310,N_3806,N_3812);
xnor U4311 (N_4311,N_3970,N_3759);
nand U4312 (N_4312,N_3836,N_3922);
nor U4313 (N_4313,N_3798,N_3973);
or U4314 (N_4314,N_3502,N_3618);
nand U4315 (N_4315,N_3773,N_3723);
xnor U4316 (N_4316,N_3864,N_3627);
or U4317 (N_4317,N_3995,N_3752);
nand U4318 (N_4318,N_3648,N_3845);
or U4319 (N_4319,N_3534,N_3770);
nor U4320 (N_4320,N_3529,N_3918);
and U4321 (N_4321,N_3950,N_3786);
and U4322 (N_4322,N_3776,N_3930);
nand U4323 (N_4323,N_3677,N_3894);
nand U4324 (N_4324,N_3635,N_3960);
xnor U4325 (N_4325,N_3597,N_3568);
xor U4326 (N_4326,N_3899,N_3831);
nand U4327 (N_4327,N_3835,N_3723);
nand U4328 (N_4328,N_3758,N_3998);
nand U4329 (N_4329,N_3950,N_3624);
nand U4330 (N_4330,N_3782,N_3925);
or U4331 (N_4331,N_3615,N_3747);
nand U4332 (N_4332,N_3811,N_3548);
nor U4333 (N_4333,N_3857,N_3777);
xnor U4334 (N_4334,N_3736,N_3985);
xnor U4335 (N_4335,N_3765,N_3730);
nand U4336 (N_4336,N_3907,N_3585);
or U4337 (N_4337,N_3596,N_3660);
xnor U4338 (N_4338,N_3913,N_3720);
nor U4339 (N_4339,N_3703,N_3631);
xor U4340 (N_4340,N_3596,N_3620);
and U4341 (N_4341,N_3539,N_3867);
or U4342 (N_4342,N_3765,N_3735);
nand U4343 (N_4343,N_3794,N_3530);
nand U4344 (N_4344,N_3943,N_3707);
nand U4345 (N_4345,N_3946,N_3985);
and U4346 (N_4346,N_3677,N_3593);
nor U4347 (N_4347,N_3961,N_3719);
xnor U4348 (N_4348,N_3866,N_3731);
nand U4349 (N_4349,N_3899,N_3857);
nand U4350 (N_4350,N_3822,N_3923);
and U4351 (N_4351,N_3799,N_3603);
nand U4352 (N_4352,N_3674,N_3833);
nor U4353 (N_4353,N_3794,N_3796);
nand U4354 (N_4354,N_3525,N_3509);
and U4355 (N_4355,N_3719,N_3761);
xor U4356 (N_4356,N_3957,N_3761);
nand U4357 (N_4357,N_3799,N_3821);
and U4358 (N_4358,N_3835,N_3906);
nor U4359 (N_4359,N_3779,N_3563);
nand U4360 (N_4360,N_3775,N_3706);
xnor U4361 (N_4361,N_3784,N_3835);
xor U4362 (N_4362,N_3604,N_3732);
nor U4363 (N_4363,N_3814,N_3679);
and U4364 (N_4364,N_3669,N_3816);
xor U4365 (N_4365,N_3647,N_3740);
and U4366 (N_4366,N_3873,N_3737);
and U4367 (N_4367,N_3585,N_3956);
nand U4368 (N_4368,N_3685,N_3943);
xor U4369 (N_4369,N_3794,N_3564);
and U4370 (N_4370,N_3621,N_3738);
nor U4371 (N_4371,N_3689,N_3739);
nand U4372 (N_4372,N_3883,N_3539);
or U4373 (N_4373,N_3562,N_3795);
and U4374 (N_4374,N_3761,N_3564);
nor U4375 (N_4375,N_3927,N_3672);
xor U4376 (N_4376,N_3789,N_3871);
nand U4377 (N_4377,N_3898,N_3693);
nor U4378 (N_4378,N_3687,N_3964);
or U4379 (N_4379,N_3770,N_3611);
nand U4380 (N_4380,N_3926,N_3743);
and U4381 (N_4381,N_3601,N_3799);
nand U4382 (N_4382,N_3678,N_3851);
xor U4383 (N_4383,N_3835,N_3538);
or U4384 (N_4384,N_3967,N_3670);
or U4385 (N_4385,N_3546,N_3707);
nand U4386 (N_4386,N_3800,N_3919);
nor U4387 (N_4387,N_3978,N_3957);
or U4388 (N_4388,N_3846,N_3983);
xnor U4389 (N_4389,N_3752,N_3788);
nand U4390 (N_4390,N_3554,N_3555);
or U4391 (N_4391,N_3772,N_3795);
or U4392 (N_4392,N_3748,N_3521);
nand U4393 (N_4393,N_3976,N_3685);
nand U4394 (N_4394,N_3579,N_3620);
nand U4395 (N_4395,N_3534,N_3639);
nor U4396 (N_4396,N_3943,N_3503);
nand U4397 (N_4397,N_3784,N_3752);
nand U4398 (N_4398,N_3724,N_3796);
or U4399 (N_4399,N_3719,N_3703);
nor U4400 (N_4400,N_3733,N_3508);
and U4401 (N_4401,N_3511,N_3924);
or U4402 (N_4402,N_3656,N_3973);
nand U4403 (N_4403,N_3874,N_3576);
and U4404 (N_4404,N_3710,N_3791);
or U4405 (N_4405,N_3931,N_3544);
xnor U4406 (N_4406,N_3771,N_3805);
nand U4407 (N_4407,N_3530,N_3690);
nand U4408 (N_4408,N_3884,N_3869);
nor U4409 (N_4409,N_3776,N_3906);
xnor U4410 (N_4410,N_3988,N_3856);
nor U4411 (N_4411,N_3570,N_3698);
and U4412 (N_4412,N_3661,N_3560);
nor U4413 (N_4413,N_3507,N_3757);
or U4414 (N_4414,N_3536,N_3560);
xnor U4415 (N_4415,N_3803,N_3746);
nor U4416 (N_4416,N_3557,N_3715);
xnor U4417 (N_4417,N_3833,N_3929);
and U4418 (N_4418,N_3851,N_3758);
and U4419 (N_4419,N_3789,N_3631);
xnor U4420 (N_4420,N_3648,N_3579);
nor U4421 (N_4421,N_3927,N_3713);
and U4422 (N_4422,N_3966,N_3725);
and U4423 (N_4423,N_3885,N_3529);
nand U4424 (N_4424,N_3909,N_3530);
nand U4425 (N_4425,N_3937,N_3823);
nand U4426 (N_4426,N_3537,N_3568);
nand U4427 (N_4427,N_3715,N_3660);
and U4428 (N_4428,N_3783,N_3724);
or U4429 (N_4429,N_3910,N_3739);
xnor U4430 (N_4430,N_3756,N_3915);
nor U4431 (N_4431,N_3634,N_3783);
xnor U4432 (N_4432,N_3519,N_3534);
or U4433 (N_4433,N_3557,N_3762);
nand U4434 (N_4434,N_3874,N_3668);
nor U4435 (N_4435,N_3640,N_3923);
xor U4436 (N_4436,N_3963,N_3674);
and U4437 (N_4437,N_3535,N_3970);
nand U4438 (N_4438,N_3943,N_3558);
or U4439 (N_4439,N_3626,N_3697);
nand U4440 (N_4440,N_3735,N_3612);
nor U4441 (N_4441,N_3810,N_3893);
nor U4442 (N_4442,N_3629,N_3905);
nor U4443 (N_4443,N_3871,N_3802);
nand U4444 (N_4444,N_3522,N_3779);
nand U4445 (N_4445,N_3809,N_3773);
or U4446 (N_4446,N_3722,N_3571);
or U4447 (N_4447,N_3963,N_3573);
and U4448 (N_4448,N_3974,N_3794);
xnor U4449 (N_4449,N_3908,N_3985);
nor U4450 (N_4450,N_3530,N_3602);
or U4451 (N_4451,N_3942,N_3646);
or U4452 (N_4452,N_3933,N_3527);
nand U4453 (N_4453,N_3958,N_3815);
or U4454 (N_4454,N_3841,N_3945);
nand U4455 (N_4455,N_3879,N_3599);
nor U4456 (N_4456,N_3677,N_3607);
xnor U4457 (N_4457,N_3613,N_3614);
xor U4458 (N_4458,N_3688,N_3860);
and U4459 (N_4459,N_3989,N_3920);
and U4460 (N_4460,N_3750,N_3697);
nor U4461 (N_4461,N_3776,N_3722);
and U4462 (N_4462,N_3908,N_3974);
or U4463 (N_4463,N_3893,N_3571);
and U4464 (N_4464,N_3660,N_3645);
and U4465 (N_4465,N_3636,N_3894);
xor U4466 (N_4466,N_3854,N_3503);
or U4467 (N_4467,N_3761,N_3882);
or U4468 (N_4468,N_3931,N_3832);
nand U4469 (N_4469,N_3802,N_3518);
or U4470 (N_4470,N_3771,N_3504);
nor U4471 (N_4471,N_3960,N_3510);
and U4472 (N_4472,N_3626,N_3782);
and U4473 (N_4473,N_3980,N_3919);
xor U4474 (N_4474,N_3852,N_3853);
or U4475 (N_4475,N_3604,N_3726);
nor U4476 (N_4476,N_3548,N_3802);
or U4477 (N_4477,N_3859,N_3991);
or U4478 (N_4478,N_3569,N_3999);
and U4479 (N_4479,N_3991,N_3828);
xnor U4480 (N_4480,N_3965,N_3720);
xnor U4481 (N_4481,N_3839,N_3999);
xnor U4482 (N_4482,N_3988,N_3707);
and U4483 (N_4483,N_3518,N_3728);
nand U4484 (N_4484,N_3755,N_3696);
or U4485 (N_4485,N_3892,N_3975);
and U4486 (N_4486,N_3539,N_3806);
nor U4487 (N_4487,N_3836,N_3866);
nand U4488 (N_4488,N_3894,N_3967);
nor U4489 (N_4489,N_3990,N_3963);
nand U4490 (N_4490,N_3697,N_3971);
nand U4491 (N_4491,N_3704,N_3944);
xor U4492 (N_4492,N_3511,N_3770);
nor U4493 (N_4493,N_3991,N_3715);
nor U4494 (N_4494,N_3579,N_3874);
nand U4495 (N_4495,N_3515,N_3900);
and U4496 (N_4496,N_3808,N_3678);
nor U4497 (N_4497,N_3603,N_3979);
and U4498 (N_4498,N_3582,N_3926);
and U4499 (N_4499,N_3876,N_3639);
and U4500 (N_4500,N_4267,N_4154);
and U4501 (N_4501,N_4421,N_4079);
xnor U4502 (N_4502,N_4362,N_4031);
nand U4503 (N_4503,N_4100,N_4022);
nand U4504 (N_4504,N_4192,N_4176);
xnor U4505 (N_4505,N_4078,N_4067);
or U4506 (N_4506,N_4372,N_4404);
xnor U4507 (N_4507,N_4481,N_4265);
or U4508 (N_4508,N_4204,N_4315);
nand U4509 (N_4509,N_4274,N_4158);
nor U4510 (N_4510,N_4209,N_4417);
xnor U4511 (N_4511,N_4374,N_4430);
xnor U4512 (N_4512,N_4243,N_4260);
nand U4513 (N_4513,N_4280,N_4049);
or U4514 (N_4514,N_4188,N_4494);
nor U4515 (N_4515,N_4458,N_4488);
nand U4516 (N_4516,N_4091,N_4075);
or U4517 (N_4517,N_4087,N_4097);
or U4518 (N_4518,N_4455,N_4042);
and U4519 (N_4519,N_4223,N_4196);
or U4520 (N_4520,N_4117,N_4189);
xor U4521 (N_4521,N_4376,N_4418);
or U4522 (N_4522,N_4283,N_4318);
and U4523 (N_4523,N_4407,N_4380);
xor U4524 (N_4524,N_4403,N_4433);
and U4525 (N_4525,N_4195,N_4186);
and U4526 (N_4526,N_4304,N_4056);
or U4527 (N_4527,N_4307,N_4227);
nor U4528 (N_4528,N_4353,N_4420);
nor U4529 (N_4529,N_4104,N_4369);
nand U4530 (N_4530,N_4037,N_4301);
nand U4531 (N_4531,N_4244,N_4144);
nand U4532 (N_4532,N_4487,N_4480);
nor U4533 (N_4533,N_4450,N_4469);
nor U4534 (N_4534,N_4239,N_4303);
or U4535 (N_4535,N_4386,N_4090);
nand U4536 (N_4536,N_4083,N_4016);
xor U4537 (N_4537,N_4497,N_4174);
nand U4538 (N_4538,N_4214,N_4366);
and U4539 (N_4539,N_4410,N_4187);
xor U4540 (N_4540,N_4228,N_4483);
and U4541 (N_4541,N_4464,N_4288);
and U4542 (N_4542,N_4477,N_4256);
xor U4543 (N_4543,N_4416,N_4355);
nand U4544 (N_4544,N_4440,N_4019);
xnor U4545 (N_4545,N_4065,N_4479);
and U4546 (N_4546,N_4027,N_4147);
nand U4547 (N_4547,N_4308,N_4368);
or U4548 (N_4548,N_4473,N_4377);
or U4549 (N_4549,N_4086,N_4453);
nor U4550 (N_4550,N_4206,N_4330);
nand U4551 (N_4551,N_4305,N_4391);
nand U4552 (N_4552,N_4482,N_4169);
xnor U4553 (N_4553,N_4264,N_4146);
xor U4554 (N_4554,N_4287,N_4413);
xnor U4555 (N_4555,N_4080,N_4092);
and U4556 (N_4556,N_4339,N_4284);
nand U4557 (N_4557,N_4360,N_4250);
or U4558 (N_4558,N_4061,N_4492);
or U4559 (N_4559,N_4363,N_4498);
and U4560 (N_4560,N_4200,N_4069);
nor U4561 (N_4561,N_4050,N_4249);
nor U4562 (N_4562,N_4382,N_4132);
xor U4563 (N_4563,N_4014,N_4229);
xnor U4564 (N_4564,N_4118,N_4023);
and U4565 (N_4565,N_4460,N_4359);
xor U4566 (N_4566,N_4313,N_4052);
and U4567 (N_4567,N_4438,N_4058);
xor U4568 (N_4568,N_4152,N_4185);
nor U4569 (N_4569,N_4443,N_4322);
nand U4570 (N_4570,N_4142,N_4039);
or U4571 (N_4571,N_4384,N_4066);
and U4572 (N_4572,N_4338,N_4140);
xor U4573 (N_4573,N_4399,N_4074);
or U4574 (N_4574,N_4323,N_4178);
and U4575 (N_4575,N_4105,N_4451);
nand U4576 (N_4576,N_4225,N_4110);
and U4577 (N_4577,N_4115,N_4112);
or U4578 (N_4578,N_4343,N_4390);
or U4579 (N_4579,N_4128,N_4231);
or U4580 (N_4580,N_4414,N_4224);
nand U4581 (N_4581,N_4150,N_4036);
or U4582 (N_4582,N_4300,N_4004);
nand U4583 (N_4583,N_4325,N_4337);
xor U4584 (N_4584,N_4401,N_4435);
nor U4585 (N_4585,N_4070,N_4046);
or U4586 (N_4586,N_4317,N_4254);
xor U4587 (N_4587,N_4261,N_4082);
nand U4588 (N_4588,N_4426,N_4094);
or U4589 (N_4589,N_4273,N_4306);
or U4590 (N_4590,N_4235,N_4099);
or U4591 (N_4591,N_4044,N_4275);
and U4592 (N_4592,N_4020,N_4032);
or U4593 (N_4593,N_4375,N_4166);
nand U4594 (N_4594,N_4373,N_4486);
nand U4595 (N_4595,N_4124,N_4212);
or U4596 (N_4596,N_4262,N_4157);
nand U4597 (N_4597,N_4495,N_4471);
and U4598 (N_4598,N_4015,N_4448);
and U4599 (N_4599,N_4457,N_4321);
nor U4600 (N_4600,N_4397,N_4012);
nor U4601 (N_4601,N_4352,N_4412);
xnor U4602 (N_4602,N_4356,N_4123);
or U4603 (N_4603,N_4029,N_4278);
xor U4604 (N_4604,N_4135,N_4311);
nor U4605 (N_4605,N_4161,N_4345);
and U4606 (N_4606,N_4340,N_4168);
nand U4607 (N_4607,N_4428,N_4470);
nand U4608 (N_4608,N_4038,N_4441);
nor U4609 (N_4609,N_4127,N_4381);
and U4610 (N_4610,N_4259,N_4093);
or U4611 (N_4611,N_4474,N_4002);
nor U4612 (N_4612,N_4272,N_4326);
and U4613 (N_4613,N_4449,N_4263);
nand U4614 (N_4614,N_4172,N_4437);
xnor U4615 (N_4615,N_4021,N_4462);
or U4616 (N_4616,N_4191,N_4130);
xor U4617 (N_4617,N_4309,N_4442);
or U4618 (N_4618,N_4107,N_4496);
and U4619 (N_4619,N_4145,N_4134);
or U4620 (N_4620,N_4162,N_4222);
or U4621 (N_4621,N_4063,N_4490);
or U4622 (N_4622,N_4139,N_4408);
nor U4623 (N_4623,N_4108,N_4351);
or U4624 (N_4624,N_4217,N_4011);
or U4625 (N_4625,N_4076,N_4137);
and U4626 (N_4626,N_4296,N_4276);
nor U4627 (N_4627,N_4255,N_4201);
nor U4628 (N_4628,N_4047,N_4489);
nand U4629 (N_4629,N_4348,N_4153);
or U4630 (N_4630,N_4095,N_4444);
nand U4631 (N_4631,N_4432,N_4336);
nand U4632 (N_4632,N_4247,N_4310);
or U4633 (N_4633,N_4314,N_4060);
or U4634 (N_4634,N_4251,N_4171);
nand U4635 (N_4635,N_4281,N_4024);
nor U4636 (N_4636,N_4294,N_4071);
xor U4637 (N_4637,N_4041,N_4207);
or U4638 (N_4638,N_4165,N_4088);
nor U4639 (N_4639,N_4387,N_4389);
nand U4640 (N_4640,N_4051,N_4111);
nand U4641 (N_4641,N_4151,N_4491);
nand U4642 (N_4642,N_4395,N_4478);
xor U4643 (N_4643,N_4354,N_4447);
nor U4644 (N_4644,N_4148,N_4211);
and U4645 (N_4645,N_4238,N_4269);
or U4646 (N_4646,N_4160,N_4468);
nand U4647 (N_4647,N_4106,N_4102);
nor U4648 (N_4648,N_4003,N_4329);
xor U4649 (N_4649,N_4485,N_4400);
or U4650 (N_4650,N_4033,N_4030);
nand U4651 (N_4651,N_4257,N_4120);
and U4652 (N_4652,N_4316,N_4320);
and U4653 (N_4653,N_4084,N_4053);
nand U4654 (N_4654,N_4006,N_4347);
nor U4655 (N_4655,N_4268,N_4073);
xnor U4656 (N_4656,N_4167,N_4429);
nand U4657 (N_4657,N_4279,N_4341);
and U4658 (N_4658,N_4409,N_4126);
xnor U4659 (N_4659,N_4098,N_4210);
xnor U4660 (N_4660,N_4028,N_4233);
nor U4661 (N_4661,N_4234,N_4427);
nand U4662 (N_4662,N_4057,N_4007);
xnor U4663 (N_4663,N_4245,N_4138);
or U4664 (N_4664,N_4342,N_4371);
or U4665 (N_4665,N_4463,N_4388);
and U4666 (N_4666,N_4452,N_4220);
or U4667 (N_4667,N_4122,N_4180);
nand U4668 (N_4668,N_4045,N_4454);
xnor U4669 (N_4669,N_4163,N_4068);
or U4670 (N_4670,N_4282,N_4131);
nor U4671 (N_4671,N_4005,N_4286);
xnor U4672 (N_4672,N_4445,N_4297);
and U4673 (N_4673,N_4177,N_4232);
nor U4674 (N_4674,N_4393,N_4499);
nor U4675 (N_4675,N_4484,N_4335);
nor U4676 (N_4676,N_4461,N_4103);
and U4677 (N_4677,N_4456,N_4133);
xor U4678 (N_4678,N_4367,N_4230);
xor U4679 (N_4679,N_4170,N_4109);
or U4680 (N_4680,N_4143,N_4493);
xnor U4681 (N_4681,N_4467,N_4277);
nand U4682 (N_4682,N_4182,N_4183);
xnor U4683 (N_4683,N_4034,N_4116);
nor U4684 (N_4684,N_4017,N_4173);
nand U4685 (N_4685,N_4077,N_4018);
and U4686 (N_4686,N_4048,N_4213);
nor U4687 (N_4687,N_4365,N_4156);
or U4688 (N_4688,N_4055,N_4402);
nand U4689 (N_4689,N_4119,N_4364);
and U4690 (N_4690,N_4184,N_4101);
or U4691 (N_4691,N_4149,N_4013);
nor U4692 (N_4692,N_4334,N_4181);
and U4693 (N_4693,N_4197,N_4293);
or U4694 (N_4694,N_4327,N_4298);
nand U4695 (N_4695,N_4346,N_4290);
nand U4696 (N_4696,N_4252,N_4465);
or U4697 (N_4697,N_4246,N_4085);
and U4698 (N_4698,N_4466,N_4240);
nor U4699 (N_4699,N_4072,N_4035);
nor U4700 (N_4700,N_4439,N_4271);
and U4701 (N_4701,N_4385,N_4422);
nor U4702 (N_4702,N_4205,N_4459);
nand U4703 (N_4703,N_4008,N_4241);
xor U4704 (N_4704,N_4202,N_4129);
and U4705 (N_4705,N_4406,N_4199);
and U4706 (N_4706,N_4312,N_4411);
and U4707 (N_4707,N_4324,N_4472);
nor U4708 (N_4708,N_4394,N_4001);
nand U4709 (N_4709,N_4383,N_4319);
xnor U4710 (N_4710,N_4289,N_4136);
xor U4711 (N_4711,N_4328,N_4357);
xnor U4712 (N_4712,N_4446,N_4219);
nor U4713 (N_4713,N_4114,N_4333);
nor U4714 (N_4714,N_4064,N_4424);
xnor U4715 (N_4715,N_4370,N_4242);
or U4716 (N_4716,N_4258,N_4266);
or U4717 (N_4717,N_4436,N_4419);
nor U4718 (N_4718,N_4292,N_4026);
nand U4719 (N_4719,N_4125,N_4216);
xnor U4720 (N_4720,N_4010,N_4331);
or U4721 (N_4721,N_4113,N_4175);
nor U4722 (N_4722,N_4295,N_4203);
and U4723 (N_4723,N_4159,N_4081);
and U4724 (N_4724,N_4164,N_4361);
nor U4725 (N_4725,N_4270,N_4398);
and U4726 (N_4726,N_4194,N_4434);
xor U4727 (N_4727,N_4096,N_4193);
xnor U4728 (N_4728,N_4155,N_4291);
nand U4729 (N_4729,N_4302,N_4226);
nor U4730 (N_4730,N_4344,N_4040);
nand U4731 (N_4731,N_4423,N_4425);
or U4732 (N_4732,N_4236,N_4043);
or U4733 (N_4733,N_4121,N_4221);
or U4734 (N_4734,N_4000,N_4358);
nand U4735 (N_4735,N_4350,N_4431);
and U4736 (N_4736,N_4025,N_4089);
and U4737 (N_4737,N_4179,N_4208);
and U4738 (N_4738,N_4059,N_4332);
nand U4739 (N_4739,N_4253,N_4392);
and U4740 (N_4740,N_4215,N_4396);
xnor U4741 (N_4741,N_4299,N_4054);
xnor U4742 (N_4742,N_4349,N_4379);
or U4743 (N_4743,N_4218,N_4405);
nor U4744 (N_4744,N_4476,N_4141);
nor U4745 (N_4745,N_4415,N_4237);
nand U4746 (N_4746,N_4062,N_4009);
nor U4747 (N_4747,N_4475,N_4198);
nor U4748 (N_4748,N_4248,N_4285);
nand U4749 (N_4749,N_4378,N_4190);
nand U4750 (N_4750,N_4345,N_4319);
nand U4751 (N_4751,N_4196,N_4438);
xnor U4752 (N_4752,N_4275,N_4027);
xnor U4753 (N_4753,N_4451,N_4421);
nor U4754 (N_4754,N_4139,N_4062);
or U4755 (N_4755,N_4284,N_4252);
nor U4756 (N_4756,N_4418,N_4032);
and U4757 (N_4757,N_4453,N_4301);
xor U4758 (N_4758,N_4447,N_4458);
and U4759 (N_4759,N_4394,N_4478);
xor U4760 (N_4760,N_4382,N_4082);
or U4761 (N_4761,N_4276,N_4364);
nor U4762 (N_4762,N_4271,N_4120);
nor U4763 (N_4763,N_4291,N_4432);
or U4764 (N_4764,N_4422,N_4418);
nor U4765 (N_4765,N_4331,N_4400);
nand U4766 (N_4766,N_4030,N_4163);
or U4767 (N_4767,N_4476,N_4046);
and U4768 (N_4768,N_4383,N_4410);
or U4769 (N_4769,N_4479,N_4422);
nand U4770 (N_4770,N_4487,N_4430);
or U4771 (N_4771,N_4046,N_4302);
xnor U4772 (N_4772,N_4445,N_4260);
and U4773 (N_4773,N_4367,N_4266);
or U4774 (N_4774,N_4021,N_4099);
or U4775 (N_4775,N_4214,N_4333);
xor U4776 (N_4776,N_4491,N_4170);
xnor U4777 (N_4777,N_4277,N_4217);
and U4778 (N_4778,N_4064,N_4376);
nor U4779 (N_4779,N_4351,N_4046);
xnor U4780 (N_4780,N_4478,N_4193);
or U4781 (N_4781,N_4317,N_4476);
or U4782 (N_4782,N_4358,N_4403);
and U4783 (N_4783,N_4367,N_4368);
or U4784 (N_4784,N_4470,N_4300);
or U4785 (N_4785,N_4316,N_4374);
nor U4786 (N_4786,N_4191,N_4030);
and U4787 (N_4787,N_4110,N_4403);
nand U4788 (N_4788,N_4081,N_4285);
and U4789 (N_4789,N_4128,N_4030);
or U4790 (N_4790,N_4143,N_4033);
and U4791 (N_4791,N_4173,N_4448);
or U4792 (N_4792,N_4102,N_4094);
or U4793 (N_4793,N_4231,N_4120);
nand U4794 (N_4794,N_4307,N_4260);
or U4795 (N_4795,N_4224,N_4252);
and U4796 (N_4796,N_4460,N_4301);
and U4797 (N_4797,N_4459,N_4386);
nor U4798 (N_4798,N_4302,N_4446);
nor U4799 (N_4799,N_4216,N_4480);
xnor U4800 (N_4800,N_4229,N_4310);
nand U4801 (N_4801,N_4367,N_4006);
nand U4802 (N_4802,N_4154,N_4227);
nor U4803 (N_4803,N_4459,N_4247);
nand U4804 (N_4804,N_4016,N_4155);
and U4805 (N_4805,N_4058,N_4345);
or U4806 (N_4806,N_4201,N_4454);
xnor U4807 (N_4807,N_4028,N_4207);
and U4808 (N_4808,N_4244,N_4021);
and U4809 (N_4809,N_4436,N_4332);
nand U4810 (N_4810,N_4146,N_4265);
or U4811 (N_4811,N_4045,N_4193);
xor U4812 (N_4812,N_4186,N_4469);
nand U4813 (N_4813,N_4381,N_4492);
or U4814 (N_4814,N_4220,N_4154);
nor U4815 (N_4815,N_4171,N_4008);
or U4816 (N_4816,N_4267,N_4454);
nand U4817 (N_4817,N_4233,N_4372);
and U4818 (N_4818,N_4422,N_4073);
and U4819 (N_4819,N_4487,N_4439);
and U4820 (N_4820,N_4078,N_4190);
xnor U4821 (N_4821,N_4189,N_4180);
and U4822 (N_4822,N_4421,N_4373);
nor U4823 (N_4823,N_4431,N_4382);
xnor U4824 (N_4824,N_4198,N_4101);
nor U4825 (N_4825,N_4334,N_4320);
or U4826 (N_4826,N_4053,N_4109);
nand U4827 (N_4827,N_4386,N_4275);
nand U4828 (N_4828,N_4414,N_4161);
nor U4829 (N_4829,N_4474,N_4484);
xor U4830 (N_4830,N_4195,N_4094);
and U4831 (N_4831,N_4428,N_4388);
and U4832 (N_4832,N_4434,N_4338);
nor U4833 (N_4833,N_4011,N_4460);
and U4834 (N_4834,N_4055,N_4447);
and U4835 (N_4835,N_4244,N_4190);
nor U4836 (N_4836,N_4290,N_4113);
nand U4837 (N_4837,N_4170,N_4399);
and U4838 (N_4838,N_4199,N_4258);
xor U4839 (N_4839,N_4147,N_4201);
and U4840 (N_4840,N_4230,N_4229);
nor U4841 (N_4841,N_4064,N_4094);
or U4842 (N_4842,N_4395,N_4497);
xnor U4843 (N_4843,N_4411,N_4313);
and U4844 (N_4844,N_4234,N_4382);
and U4845 (N_4845,N_4301,N_4046);
nor U4846 (N_4846,N_4199,N_4077);
xnor U4847 (N_4847,N_4087,N_4308);
nand U4848 (N_4848,N_4028,N_4428);
or U4849 (N_4849,N_4353,N_4104);
nand U4850 (N_4850,N_4243,N_4027);
nand U4851 (N_4851,N_4409,N_4322);
nor U4852 (N_4852,N_4339,N_4332);
nor U4853 (N_4853,N_4253,N_4044);
nor U4854 (N_4854,N_4384,N_4441);
and U4855 (N_4855,N_4050,N_4408);
xnor U4856 (N_4856,N_4050,N_4064);
and U4857 (N_4857,N_4381,N_4495);
nand U4858 (N_4858,N_4217,N_4226);
nand U4859 (N_4859,N_4025,N_4177);
and U4860 (N_4860,N_4276,N_4398);
nand U4861 (N_4861,N_4158,N_4009);
xor U4862 (N_4862,N_4294,N_4403);
nor U4863 (N_4863,N_4284,N_4143);
nor U4864 (N_4864,N_4266,N_4099);
xnor U4865 (N_4865,N_4289,N_4303);
xor U4866 (N_4866,N_4169,N_4290);
xor U4867 (N_4867,N_4209,N_4161);
nand U4868 (N_4868,N_4367,N_4070);
and U4869 (N_4869,N_4344,N_4196);
and U4870 (N_4870,N_4200,N_4310);
and U4871 (N_4871,N_4401,N_4248);
nor U4872 (N_4872,N_4262,N_4323);
nand U4873 (N_4873,N_4496,N_4300);
nand U4874 (N_4874,N_4044,N_4161);
and U4875 (N_4875,N_4396,N_4102);
nor U4876 (N_4876,N_4378,N_4179);
and U4877 (N_4877,N_4032,N_4017);
xor U4878 (N_4878,N_4057,N_4164);
and U4879 (N_4879,N_4430,N_4088);
nor U4880 (N_4880,N_4482,N_4499);
xnor U4881 (N_4881,N_4418,N_4386);
xor U4882 (N_4882,N_4306,N_4365);
nand U4883 (N_4883,N_4487,N_4242);
nor U4884 (N_4884,N_4384,N_4313);
xnor U4885 (N_4885,N_4328,N_4495);
nor U4886 (N_4886,N_4370,N_4162);
nor U4887 (N_4887,N_4324,N_4131);
nor U4888 (N_4888,N_4280,N_4425);
xnor U4889 (N_4889,N_4002,N_4056);
nand U4890 (N_4890,N_4474,N_4379);
and U4891 (N_4891,N_4150,N_4244);
nand U4892 (N_4892,N_4364,N_4035);
nor U4893 (N_4893,N_4260,N_4098);
nor U4894 (N_4894,N_4030,N_4385);
and U4895 (N_4895,N_4282,N_4101);
nand U4896 (N_4896,N_4313,N_4016);
or U4897 (N_4897,N_4196,N_4117);
nor U4898 (N_4898,N_4469,N_4340);
and U4899 (N_4899,N_4350,N_4115);
and U4900 (N_4900,N_4231,N_4232);
or U4901 (N_4901,N_4113,N_4222);
and U4902 (N_4902,N_4408,N_4410);
xor U4903 (N_4903,N_4143,N_4341);
and U4904 (N_4904,N_4078,N_4266);
xor U4905 (N_4905,N_4350,N_4153);
or U4906 (N_4906,N_4346,N_4275);
or U4907 (N_4907,N_4085,N_4385);
xnor U4908 (N_4908,N_4264,N_4180);
nor U4909 (N_4909,N_4027,N_4297);
or U4910 (N_4910,N_4366,N_4043);
nand U4911 (N_4911,N_4494,N_4448);
nor U4912 (N_4912,N_4100,N_4371);
nand U4913 (N_4913,N_4117,N_4018);
xor U4914 (N_4914,N_4272,N_4205);
nor U4915 (N_4915,N_4157,N_4067);
nand U4916 (N_4916,N_4470,N_4129);
xor U4917 (N_4917,N_4031,N_4204);
and U4918 (N_4918,N_4426,N_4267);
xnor U4919 (N_4919,N_4369,N_4378);
and U4920 (N_4920,N_4385,N_4109);
nand U4921 (N_4921,N_4319,N_4001);
nand U4922 (N_4922,N_4296,N_4212);
and U4923 (N_4923,N_4346,N_4494);
and U4924 (N_4924,N_4219,N_4477);
nor U4925 (N_4925,N_4461,N_4494);
and U4926 (N_4926,N_4424,N_4491);
and U4927 (N_4927,N_4388,N_4093);
or U4928 (N_4928,N_4317,N_4338);
or U4929 (N_4929,N_4136,N_4040);
and U4930 (N_4930,N_4000,N_4127);
nor U4931 (N_4931,N_4196,N_4428);
or U4932 (N_4932,N_4377,N_4266);
and U4933 (N_4933,N_4191,N_4309);
nand U4934 (N_4934,N_4478,N_4057);
xnor U4935 (N_4935,N_4266,N_4313);
nor U4936 (N_4936,N_4116,N_4457);
xnor U4937 (N_4937,N_4316,N_4159);
or U4938 (N_4938,N_4273,N_4136);
nand U4939 (N_4939,N_4340,N_4028);
and U4940 (N_4940,N_4344,N_4290);
nand U4941 (N_4941,N_4116,N_4147);
nor U4942 (N_4942,N_4307,N_4190);
nand U4943 (N_4943,N_4490,N_4080);
nand U4944 (N_4944,N_4075,N_4267);
xnor U4945 (N_4945,N_4127,N_4162);
and U4946 (N_4946,N_4209,N_4447);
or U4947 (N_4947,N_4225,N_4059);
and U4948 (N_4948,N_4237,N_4287);
nor U4949 (N_4949,N_4439,N_4292);
and U4950 (N_4950,N_4168,N_4081);
or U4951 (N_4951,N_4352,N_4091);
or U4952 (N_4952,N_4189,N_4113);
and U4953 (N_4953,N_4436,N_4192);
and U4954 (N_4954,N_4050,N_4111);
xor U4955 (N_4955,N_4436,N_4243);
nor U4956 (N_4956,N_4250,N_4106);
and U4957 (N_4957,N_4101,N_4236);
nand U4958 (N_4958,N_4297,N_4045);
or U4959 (N_4959,N_4349,N_4155);
xor U4960 (N_4960,N_4165,N_4051);
and U4961 (N_4961,N_4231,N_4319);
nand U4962 (N_4962,N_4388,N_4283);
nand U4963 (N_4963,N_4108,N_4254);
nand U4964 (N_4964,N_4471,N_4266);
or U4965 (N_4965,N_4104,N_4456);
or U4966 (N_4966,N_4131,N_4295);
nor U4967 (N_4967,N_4210,N_4180);
xor U4968 (N_4968,N_4489,N_4258);
nand U4969 (N_4969,N_4176,N_4104);
and U4970 (N_4970,N_4190,N_4091);
nand U4971 (N_4971,N_4073,N_4393);
or U4972 (N_4972,N_4128,N_4028);
or U4973 (N_4973,N_4431,N_4117);
or U4974 (N_4974,N_4480,N_4019);
nand U4975 (N_4975,N_4214,N_4178);
nand U4976 (N_4976,N_4050,N_4214);
nor U4977 (N_4977,N_4228,N_4361);
nor U4978 (N_4978,N_4242,N_4275);
or U4979 (N_4979,N_4164,N_4080);
and U4980 (N_4980,N_4022,N_4231);
or U4981 (N_4981,N_4281,N_4184);
or U4982 (N_4982,N_4416,N_4136);
and U4983 (N_4983,N_4028,N_4469);
or U4984 (N_4984,N_4006,N_4230);
and U4985 (N_4985,N_4172,N_4318);
nor U4986 (N_4986,N_4247,N_4370);
or U4987 (N_4987,N_4176,N_4099);
nand U4988 (N_4988,N_4107,N_4223);
nor U4989 (N_4989,N_4037,N_4020);
nand U4990 (N_4990,N_4157,N_4046);
or U4991 (N_4991,N_4049,N_4178);
or U4992 (N_4992,N_4167,N_4271);
nand U4993 (N_4993,N_4469,N_4156);
nand U4994 (N_4994,N_4127,N_4154);
nor U4995 (N_4995,N_4433,N_4373);
xor U4996 (N_4996,N_4235,N_4259);
xor U4997 (N_4997,N_4382,N_4198);
xor U4998 (N_4998,N_4427,N_4307);
or U4999 (N_4999,N_4111,N_4442);
or UO_0 (O_0,N_4571,N_4808);
nand UO_1 (O_1,N_4585,N_4605);
nor UO_2 (O_2,N_4826,N_4617);
xnor UO_3 (O_3,N_4980,N_4880);
or UO_4 (O_4,N_4893,N_4700);
or UO_5 (O_5,N_4950,N_4570);
and UO_6 (O_6,N_4939,N_4833);
xnor UO_7 (O_7,N_4533,N_4793);
or UO_8 (O_8,N_4972,N_4745);
nor UO_9 (O_9,N_4650,N_4866);
or UO_10 (O_10,N_4747,N_4654);
nor UO_11 (O_11,N_4809,N_4759);
and UO_12 (O_12,N_4639,N_4626);
xnor UO_13 (O_13,N_4872,N_4841);
xnor UO_14 (O_14,N_4951,N_4848);
nor UO_15 (O_15,N_4675,N_4858);
and UO_16 (O_16,N_4554,N_4910);
and UO_17 (O_17,N_4727,N_4977);
xor UO_18 (O_18,N_4991,N_4843);
nor UO_19 (O_19,N_4622,N_4688);
nor UO_20 (O_20,N_4876,N_4935);
or UO_21 (O_21,N_4659,N_4800);
xor UO_22 (O_22,N_4803,N_4953);
and UO_23 (O_23,N_4616,N_4899);
and UO_24 (O_24,N_4780,N_4853);
xor UO_25 (O_25,N_4529,N_4805);
nand UO_26 (O_26,N_4658,N_4543);
and UO_27 (O_27,N_4515,N_4721);
or UO_28 (O_28,N_4936,N_4922);
and UO_29 (O_29,N_4924,N_4752);
nand UO_30 (O_30,N_4589,N_4844);
xnor UO_31 (O_31,N_4846,N_4764);
nor UO_32 (O_32,N_4662,N_4535);
or UO_33 (O_33,N_4896,N_4546);
or UO_34 (O_34,N_4537,N_4649);
nand UO_35 (O_35,N_4687,N_4786);
xor UO_36 (O_36,N_4845,N_4566);
or UO_37 (O_37,N_4967,N_4593);
or UO_38 (O_38,N_4864,N_4979);
xor UO_39 (O_39,N_4725,N_4509);
xor UO_40 (O_40,N_4734,N_4847);
xor UO_41 (O_41,N_4520,N_4988);
nand UO_42 (O_42,N_4886,N_4981);
xnor UO_43 (O_43,N_4825,N_4601);
nor UO_44 (O_44,N_4806,N_4708);
or UO_45 (O_45,N_4768,N_4637);
xnor UO_46 (O_46,N_4653,N_4900);
and UO_47 (O_47,N_4770,N_4540);
and UO_48 (O_48,N_4850,N_4565);
nor UO_49 (O_49,N_4606,N_4836);
nor UO_50 (O_50,N_4691,N_4802);
nor UO_51 (O_51,N_4577,N_4792);
nor UO_52 (O_52,N_4871,N_4726);
and UO_53 (O_53,N_4774,N_4735);
xor UO_54 (O_54,N_4832,N_4628);
nand UO_55 (O_55,N_4569,N_4568);
or UO_56 (O_56,N_4859,N_4519);
and UO_57 (O_57,N_4916,N_4968);
xor UO_58 (O_58,N_4706,N_4909);
xor UO_59 (O_59,N_4817,N_4913);
xor UO_60 (O_60,N_4995,N_4647);
nor UO_61 (O_61,N_4771,N_4629);
and UO_62 (O_62,N_4831,N_4711);
nand UO_63 (O_63,N_4563,N_4713);
or UO_64 (O_64,N_4757,N_4633);
or UO_65 (O_65,N_4723,N_4552);
xnor UO_66 (O_66,N_4652,N_4631);
xor UO_67 (O_67,N_4720,N_4765);
xor UO_68 (O_68,N_4962,N_4942);
nand UO_69 (O_69,N_4663,N_4999);
nor UO_70 (O_70,N_4561,N_4505);
xnor UO_71 (O_71,N_4906,N_4709);
nand UO_72 (O_72,N_4615,N_4938);
nand UO_73 (O_73,N_4665,N_4949);
and UO_74 (O_74,N_4672,N_4915);
and UO_75 (O_75,N_4590,N_4702);
xnor UO_76 (O_76,N_4545,N_4588);
or UO_77 (O_77,N_4573,N_4963);
and UO_78 (O_78,N_4661,N_4816);
nand UO_79 (O_79,N_4506,N_4842);
xnor UO_80 (O_80,N_4984,N_4586);
and UO_81 (O_81,N_4576,N_4503);
xor UO_82 (O_82,N_4874,N_4599);
xnor UO_83 (O_83,N_4697,N_4969);
nand UO_84 (O_84,N_4990,N_4591);
and UO_85 (O_85,N_4685,N_4901);
nand UO_86 (O_86,N_4978,N_4557);
or UO_87 (O_87,N_4829,N_4992);
xnor UO_88 (O_88,N_4592,N_4891);
nor UO_89 (O_89,N_4614,N_4609);
nand UO_90 (O_90,N_4987,N_4690);
nor UO_91 (O_91,N_4536,N_4862);
nand UO_92 (O_92,N_4798,N_4676);
nand UO_93 (O_93,N_4716,N_4587);
or UO_94 (O_94,N_4905,N_4553);
nand UO_95 (O_95,N_4550,N_4572);
nor UO_96 (O_96,N_4904,N_4743);
nand UO_97 (O_97,N_4739,N_4917);
or UO_98 (O_98,N_4870,N_4889);
xnor UO_99 (O_99,N_4783,N_4973);
xor UO_100 (O_100,N_4941,N_4983);
nand UO_101 (O_101,N_4584,N_4890);
xnor UO_102 (O_102,N_4753,N_4998);
xor UO_103 (O_103,N_4982,N_4948);
xnor UO_104 (O_104,N_4797,N_4952);
or UO_105 (O_105,N_4641,N_4737);
or UO_106 (O_106,N_4531,N_4878);
nor UO_107 (O_107,N_4994,N_4532);
nand UO_108 (O_108,N_4856,N_4908);
or UO_109 (O_109,N_4501,N_4594);
nand UO_110 (O_110,N_4744,N_4667);
xnor UO_111 (O_111,N_4681,N_4732);
and UO_112 (O_112,N_4863,N_4632);
and UO_113 (O_113,N_4551,N_4898);
nor UO_114 (O_114,N_4789,N_4818);
xnor UO_115 (O_115,N_4640,N_4526);
or UO_116 (O_116,N_4881,N_4674);
and UO_117 (O_117,N_4696,N_4855);
nor UO_118 (O_118,N_4927,N_4758);
nand UO_119 (O_119,N_4760,N_4542);
nor UO_120 (O_120,N_4717,N_4555);
xor UO_121 (O_121,N_4600,N_4656);
and UO_122 (O_122,N_4620,N_4582);
nor UO_123 (O_123,N_4527,N_4779);
and UO_124 (O_124,N_4643,N_4560);
nor UO_125 (O_125,N_4705,N_4903);
or UO_126 (O_126,N_4611,N_4767);
nor UO_127 (O_127,N_4911,N_4812);
or UO_128 (O_128,N_4955,N_4823);
nor UO_129 (O_129,N_4539,N_4677);
and UO_130 (O_130,N_4794,N_4695);
nor UO_131 (O_131,N_4883,N_4714);
xnor UO_132 (O_132,N_4579,N_4921);
or UO_133 (O_133,N_4960,N_4873);
and UO_134 (O_134,N_4651,N_4644);
or UO_135 (O_135,N_4799,N_4508);
nor UO_136 (O_136,N_4610,N_4525);
or UO_137 (O_137,N_4929,N_4678);
xor UO_138 (O_138,N_4940,N_4613);
nor UO_139 (O_139,N_4918,N_4958);
nor UO_140 (O_140,N_4869,N_4985);
xor UO_141 (O_141,N_4887,N_4602);
nor UO_142 (O_142,N_4669,N_4819);
nor UO_143 (O_143,N_4807,N_4504);
or UO_144 (O_144,N_4821,N_4666);
or UO_145 (O_145,N_4738,N_4544);
nor UO_146 (O_146,N_4699,N_4522);
xnor UO_147 (O_147,N_4868,N_4813);
nor UO_148 (O_148,N_4575,N_4603);
or UO_149 (O_149,N_4581,N_4849);
and UO_150 (O_150,N_4693,N_4934);
or UO_151 (O_151,N_4919,N_4523);
and UO_152 (O_152,N_4801,N_4943);
xor UO_153 (O_153,N_4852,N_4635);
nor UO_154 (O_154,N_4976,N_4736);
nand UO_155 (O_155,N_4820,N_4810);
and UO_156 (O_156,N_4882,N_4875);
and UO_157 (O_157,N_4703,N_4507);
xor UO_158 (O_158,N_4785,N_4623);
nor UO_159 (O_159,N_4621,N_4791);
xnor UO_160 (O_160,N_4733,N_4837);
xnor UO_161 (O_161,N_4701,N_4625);
or UO_162 (O_162,N_4974,N_4838);
or UO_163 (O_163,N_4928,N_4558);
and UO_164 (O_164,N_4636,N_4517);
nand UO_165 (O_165,N_4954,N_4634);
xor UO_166 (O_166,N_4930,N_4728);
xnor UO_167 (O_167,N_4993,N_4648);
and UO_168 (O_168,N_4902,N_4567);
or UO_169 (O_169,N_4756,N_4684);
and UO_170 (O_170,N_4989,N_4777);
nand UO_171 (O_171,N_4944,N_4692);
nor UO_172 (O_172,N_4814,N_4740);
or UO_173 (O_173,N_4754,N_4679);
and UO_174 (O_174,N_4719,N_4835);
nand UO_175 (O_175,N_4923,N_4556);
nand UO_176 (O_176,N_4782,N_4961);
xnor UO_177 (O_177,N_4907,N_4524);
nor UO_178 (O_178,N_4502,N_4975);
or UO_179 (O_179,N_4895,N_4996);
and UO_180 (O_180,N_4534,N_4512);
and UO_181 (O_181,N_4748,N_4627);
and UO_182 (O_182,N_4885,N_4965);
and UO_183 (O_183,N_4715,N_4755);
or UO_184 (O_184,N_4957,N_4854);
nand UO_185 (O_185,N_4638,N_4645);
and UO_186 (O_186,N_4604,N_4769);
nand UO_187 (O_187,N_4920,N_4933);
and UO_188 (O_188,N_4742,N_4897);
nor UO_189 (O_189,N_4516,N_4712);
nor UO_190 (O_190,N_4894,N_4722);
xnor UO_191 (O_191,N_4795,N_4761);
xnor UO_192 (O_192,N_4698,N_4578);
or UO_193 (O_193,N_4528,N_4860);
nor UO_194 (O_194,N_4945,N_4784);
and UO_195 (O_195,N_4530,N_4559);
and UO_196 (O_196,N_4877,N_4660);
nand UO_197 (O_197,N_4763,N_4966);
nor UO_198 (O_198,N_4834,N_4619);
nand UO_199 (O_199,N_4959,N_4549);
xnor UO_200 (O_200,N_4773,N_4513);
or UO_201 (O_201,N_4607,N_4657);
nand UO_202 (O_202,N_4861,N_4689);
and UO_203 (O_203,N_4946,N_4564);
nand UO_204 (O_204,N_4932,N_4787);
xor UO_205 (O_205,N_4630,N_4562);
nor UO_206 (O_206,N_4741,N_4704);
or UO_207 (O_207,N_4673,N_4914);
nor UO_208 (O_208,N_4824,N_4680);
or UO_209 (O_209,N_4514,N_4964);
or UO_210 (O_210,N_4931,N_4511);
nand UO_211 (O_211,N_4925,N_4547);
and UO_212 (O_212,N_4912,N_4694);
or UO_213 (O_213,N_4682,N_4781);
xor UO_214 (O_214,N_4762,N_4775);
or UO_215 (O_215,N_4772,N_4598);
nand UO_216 (O_216,N_4751,N_4840);
and UO_217 (O_217,N_4970,N_4750);
xnor UO_218 (O_218,N_4521,N_4865);
nor UO_219 (O_219,N_4608,N_4888);
or UO_220 (O_220,N_4815,N_4851);
or UO_221 (O_221,N_4683,N_4618);
xnor UO_222 (O_222,N_4947,N_4668);
nor UO_223 (O_223,N_4796,N_4729);
xor UO_224 (O_224,N_4671,N_4776);
nand UO_225 (O_225,N_4710,N_4718);
xor UO_226 (O_226,N_4538,N_4822);
xor UO_227 (O_227,N_4956,N_4580);
nand UO_228 (O_228,N_4828,N_4655);
and UO_229 (O_229,N_4686,N_4986);
nor UO_230 (O_230,N_4788,N_4548);
nor UO_231 (O_231,N_4827,N_4597);
xnor UO_232 (O_232,N_4707,N_4884);
nand UO_233 (O_233,N_4778,N_4518);
or UO_234 (O_234,N_4997,N_4804);
or UO_235 (O_235,N_4595,N_4731);
nand UO_236 (O_236,N_4724,N_4857);
nor UO_237 (O_237,N_4790,N_4574);
nor UO_238 (O_238,N_4670,N_4646);
nand UO_239 (O_239,N_4664,N_4811);
nor UO_240 (O_240,N_4937,N_4867);
nand UO_241 (O_241,N_4510,N_4971);
xor UO_242 (O_242,N_4830,N_4766);
and UO_243 (O_243,N_4839,N_4596);
or UO_244 (O_244,N_4926,N_4749);
xor UO_245 (O_245,N_4746,N_4612);
or UO_246 (O_246,N_4500,N_4583);
or UO_247 (O_247,N_4892,N_4730);
xnor UO_248 (O_248,N_4879,N_4541);
xnor UO_249 (O_249,N_4624,N_4642);
nor UO_250 (O_250,N_4677,N_4696);
xor UO_251 (O_251,N_4907,N_4574);
and UO_252 (O_252,N_4582,N_4593);
or UO_253 (O_253,N_4770,N_4544);
xnor UO_254 (O_254,N_4739,N_4600);
xnor UO_255 (O_255,N_4838,N_4644);
and UO_256 (O_256,N_4599,N_4545);
and UO_257 (O_257,N_4505,N_4938);
xor UO_258 (O_258,N_4887,N_4541);
nand UO_259 (O_259,N_4571,N_4854);
nand UO_260 (O_260,N_4668,N_4900);
and UO_261 (O_261,N_4841,N_4581);
nand UO_262 (O_262,N_4884,N_4795);
nand UO_263 (O_263,N_4663,N_4933);
xnor UO_264 (O_264,N_4748,N_4789);
nand UO_265 (O_265,N_4993,N_4678);
nand UO_266 (O_266,N_4812,N_4572);
and UO_267 (O_267,N_4913,N_4765);
or UO_268 (O_268,N_4528,N_4646);
nor UO_269 (O_269,N_4787,N_4542);
xnor UO_270 (O_270,N_4700,N_4500);
xor UO_271 (O_271,N_4769,N_4702);
xor UO_272 (O_272,N_4816,N_4529);
xnor UO_273 (O_273,N_4642,N_4767);
xnor UO_274 (O_274,N_4812,N_4728);
nand UO_275 (O_275,N_4519,N_4664);
xor UO_276 (O_276,N_4761,N_4915);
xnor UO_277 (O_277,N_4584,N_4759);
xor UO_278 (O_278,N_4559,N_4768);
and UO_279 (O_279,N_4944,N_4553);
nand UO_280 (O_280,N_4719,N_4659);
and UO_281 (O_281,N_4763,N_4527);
or UO_282 (O_282,N_4698,N_4914);
and UO_283 (O_283,N_4907,N_4713);
nor UO_284 (O_284,N_4738,N_4832);
and UO_285 (O_285,N_4609,N_4820);
and UO_286 (O_286,N_4767,N_4517);
or UO_287 (O_287,N_4968,N_4736);
or UO_288 (O_288,N_4521,N_4922);
and UO_289 (O_289,N_4886,N_4815);
or UO_290 (O_290,N_4984,N_4614);
nand UO_291 (O_291,N_4581,N_4658);
nor UO_292 (O_292,N_4993,N_4758);
or UO_293 (O_293,N_4910,N_4530);
nor UO_294 (O_294,N_4895,N_4665);
nor UO_295 (O_295,N_4781,N_4777);
nand UO_296 (O_296,N_4822,N_4987);
xor UO_297 (O_297,N_4521,N_4893);
and UO_298 (O_298,N_4862,N_4705);
nand UO_299 (O_299,N_4695,N_4611);
and UO_300 (O_300,N_4671,N_4623);
or UO_301 (O_301,N_4878,N_4931);
xor UO_302 (O_302,N_4948,N_4985);
nor UO_303 (O_303,N_4661,N_4734);
and UO_304 (O_304,N_4511,N_4884);
and UO_305 (O_305,N_4540,N_4678);
nor UO_306 (O_306,N_4705,N_4848);
nand UO_307 (O_307,N_4717,N_4883);
nor UO_308 (O_308,N_4606,N_4947);
nand UO_309 (O_309,N_4743,N_4622);
or UO_310 (O_310,N_4612,N_4783);
or UO_311 (O_311,N_4899,N_4752);
xor UO_312 (O_312,N_4528,N_4671);
xor UO_313 (O_313,N_4527,N_4648);
nand UO_314 (O_314,N_4671,N_4613);
nor UO_315 (O_315,N_4745,N_4741);
and UO_316 (O_316,N_4753,N_4801);
nand UO_317 (O_317,N_4685,N_4506);
nor UO_318 (O_318,N_4691,N_4746);
or UO_319 (O_319,N_4814,N_4594);
and UO_320 (O_320,N_4787,N_4962);
or UO_321 (O_321,N_4714,N_4718);
and UO_322 (O_322,N_4947,N_4636);
nand UO_323 (O_323,N_4813,N_4509);
or UO_324 (O_324,N_4516,N_4611);
nor UO_325 (O_325,N_4724,N_4510);
nand UO_326 (O_326,N_4768,N_4608);
and UO_327 (O_327,N_4711,N_4572);
or UO_328 (O_328,N_4549,N_4565);
nor UO_329 (O_329,N_4968,N_4529);
xnor UO_330 (O_330,N_4864,N_4629);
nand UO_331 (O_331,N_4732,N_4617);
or UO_332 (O_332,N_4948,N_4701);
nor UO_333 (O_333,N_4640,N_4954);
xor UO_334 (O_334,N_4559,N_4504);
nor UO_335 (O_335,N_4918,N_4876);
xor UO_336 (O_336,N_4695,N_4561);
nor UO_337 (O_337,N_4530,N_4790);
nor UO_338 (O_338,N_4918,N_4943);
nor UO_339 (O_339,N_4724,N_4905);
nor UO_340 (O_340,N_4897,N_4732);
nor UO_341 (O_341,N_4755,N_4900);
and UO_342 (O_342,N_4892,N_4519);
nand UO_343 (O_343,N_4890,N_4641);
xnor UO_344 (O_344,N_4746,N_4533);
nor UO_345 (O_345,N_4689,N_4527);
or UO_346 (O_346,N_4613,N_4920);
nand UO_347 (O_347,N_4810,N_4767);
xor UO_348 (O_348,N_4988,N_4622);
or UO_349 (O_349,N_4934,N_4919);
nor UO_350 (O_350,N_4685,N_4719);
nand UO_351 (O_351,N_4844,N_4641);
xnor UO_352 (O_352,N_4960,N_4894);
xnor UO_353 (O_353,N_4748,N_4587);
nor UO_354 (O_354,N_4855,N_4595);
or UO_355 (O_355,N_4787,N_4554);
or UO_356 (O_356,N_4546,N_4680);
xnor UO_357 (O_357,N_4742,N_4883);
and UO_358 (O_358,N_4527,N_4609);
nand UO_359 (O_359,N_4990,N_4598);
and UO_360 (O_360,N_4800,N_4865);
xor UO_361 (O_361,N_4834,N_4747);
or UO_362 (O_362,N_4570,N_4517);
nand UO_363 (O_363,N_4999,N_4974);
and UO_364 (O_364,N_4612,N_4608);
xnor UO_365 (O_365,N_4675,N_4877);
xor UO_366 (O_366,N_4786,N_4804);
xnor UO_367 (O_367,N_4682,N_4604);
and UO_368 (O_368,N_4880,N_4903);
and UO_369 (O_369,N_4876,N_4753);
or UO_370 (O_370,N_4947,N_4734);
or UO_371 (O_371,N_4628,N_4833);
nand UO_372 (O_372,N_4766,N_4772);
nand UO_373 (O_373,N_4532,N_4730);
nor UO_374 (O_374,N_4986,N_4891);
nor UO_375 (O_375,N_4630,N_4574);
nand UO_376 (O_376,N_4753,N_4917);
nor UO_377 (O_377,N_4915,N_4714);
xor UO_378 (O_378,N_4834,N_4977);
xnor UO_379 (O_379,N_4976,N_4654);
nand UO_380 (O_380,N_4670,N_4666);
xnor UO_381 (O_381,N_4590,N_4676);
nor UO_382 (O_382,N_4908,N_4816);
and UO_383 (O_383,N_4688,N_4849);
and UO_384 (O_384,N_4837,N_4556);
xnor UO_385 (O_385,N_4988,N_4943);
nand UO_386 (O_386,N_4681,N_4984);
nor UO_387 (O_387,N_4593,N_4906);
nand UO_388 (O_388,N_4980,N_4767);
and UO_389 (O_389,N_4878,N_4858);
and UO_390 (O_390,N_4775,N_4703);
or UO_391 (O_391,N_4960,N_4967);
nor UO_392 (O_392,N_4949,N_4614);
nor UO_393 (O_393,N_4913,N_4966);
and UO_394 (O_394,N_4636,N_4609);
nand UO_395 (O_395,N_4908,N_4698);
or UO_396 (O_396,N_4907,N_4767);
or UO_397 (O_397,N_4756,N_4893);
xnor UO_398 (O_398,N_4699,N_4921);
nor UO_399 (O_399,N_4661,N_4513);
nor UO_400 (O_400,N_4719,N_4981);
nor UO_401 (O_401,N_4583,N_4993);
nand UO_402 (O_402,N_4657,N_4722);
nor UO_403 (O_403,N_4762,N_4963);
and UO_404 (O_404,N_4831,N_4586);
xnor UO_405 (O_405,N_4504,N_4829);
or UO_406 (O_406,N_4733,N_4699);
xor UO_407 (O_407,N_4635,N_4890);
and UO_408 (O_408,N_4648,N_4636);
and UO_409 (O_409,N_4803,N_4715);
xnor UO_410 (O_410,N_4614,N_4696);
nor UO_411 (O_411,N_4906,N_4682);
nand UO_412 (O_412,N_4668,N_4991);
nand UO_413 (O_413,N_4826,N_4837);
nor UO_414 (O_414,N_4577,N_4909);
nor UO_415 (O_415,N_4533,N_4926);
or UO_416 (O_416,N_4952,N_4525);
nand UO_417 (O_417,N_4722,N_4975);
or UO_418 (O_418,N_4940,N_4759);
xnor UO_419 (O_419,N_4554,N_4599);
and UO_420 (O_420,N_4740,N_4620);
and UO_421 (O_421,N_4571,N_4611);
nand UO_422 (O_422,N_4974,N_4721);
nor UO_423 (O_423,N_4883,N_4964);
nand UO_424 (O_424,N_4754,N_4993);
or UO_425 (O_425,N_4596,N_4737);
nand UO_426 (O_426,N_4838,N_4972);
and UO_427 (O_427,N_4648,N_4684);
or UO_428 (O_428,N_4856,N_4857);
or UO_429 (O_429,N_4751,N_4572);
or UO_430 (O_430,N_4511,N_4590);
nor UO_431 (O_431,N_4946,N_4788);
nand UO_432 (O_432,N_4844,N_4947);
nand UO_433 (O_433,N_4619,N_4717);
nand UO_434 (O_434,N_4967,N_4968);
xor UO_435 (O_435,N_4858,N_4932);
nor UO_436 (O_436,N_4617,N_4674);
xor UO_437 (O_437,N_4968,N_4822);
and UO_438 (O_438,N_4899,N_4522);
or UO_439 (O_439,N_4570,N_4753);
nor UO_440 (O_440,N_4715,N_4645);
nand UO_441 (O_441,N_4944,N_4566);
nand UO_442 (O_442,N_4903,N_4580);
or UO_443 (O_443,N_4792,N_4644);
nand UO_444 (O_444,N_4649,N_4528);
or UO_445 (O_445,N_4660,N_4806);
xor UO_446 (O_446,N_4853,N_4626);
or UO_447 (O_447,N_4554,N_4723);
nand UO_448 (O_448,N_4675,N_4813);
nor UO_449 (O_449,N_4631,N_4861);
xnor UO_450 (O_450,N_4819,N_4991);
nand UO_451 (O_451,N_4764,N_4827);
xor UO_452 (O_452,N_4741,N_4952);
and UO_453 (O_453,N_4695,N_4817);
or UO_454 (O_454,N_4660,N_4599);
xnor UO_455 (O_455,N_4987,N_4502);
or UO_456 (O_456,N_4511,N_4523);
xor UO_457 (O_457,N_4826,N_4608);
nor UO_458 (O_458,N_4796,N_4790);
nor UO_459 (O_459,N_4611,N_4896);
and UO_460 (O_460,N_4928,N_4944);
or UO_461 (O_461,N_4796,N_4673);
and UO_462 (O_462,N_4656,N_4945);
and UO_463 (O_463,N_4569,N_4661);
xor UO_464 (O_464,N_4991,N_4554);
nand UO_465 (O_465,N_4587,N_4574);
and UO_466 (O_466,N_4640,N_4603);
xor UO_467 (O_467,N_4784,N_4980);
and UO_468 (O_468,N_4716,N_4874);
and UO_469 (O_469,N_4507,N_4519);
xor UO_470 (O_470,N_4717,N_4869);
xnor UO_471 (O_471,N_4841,N_4576);
and UO_472 (O_472,N_4919,N_4969);
nand UO_473 (O_473,N_4758,N_4577);
or UO_474 (O_474,N_4536,N_4935);
xnor UO_475 (O_475,N_4611,N_4725);
or UO_476 (O_476,N_4638,N_4829);
and UO_477 (O_477,N_4799,N_4608);
xor UO_478 (O_478,N_4713,N_4616);
or UO_479 (O_479,N_4698,N_4934);
nand UO_480 (O_480,N_4771,N_4584);
xor UO_481 (O_481,N_4746,N_4917);
nand UO_482 (O_482,N_4572,N_4682);
xor UO_483 (O_483,N_4747,N_4839);
or UO_484 (O_484,N_4767,N_4605);
nand UO_485 (O_485,N_4619,N_4620);
xnor UO_486 (O_486,N_4985,N_4649);
nand UO_487 (O_487,N_4994,N_4696);
and UO_488 (O_488,N_4778,N_4914);
xor UO_489 (O_489,N_4835,N_4722);
xnor UO_490 (O_490,N_4925,N_4899);
and UO_491 (O_491,N_4665,N_4662);
and UO_492 (O_492,N_4536,N_4763);
xnor UO_493 (O_493,N_4731,N_4774);
nor UO_494 (O_494,N_4629,N_4890);
nand UO_495 (O_495,N_4780,N_4649);
nand UO_496 (O_496,N_4786,N_4851);
nand UO_497 (O_497,N_4744,N_4684);
nand UO_498 (O_498,N_4713,N_4627);
nand UO_499 (O_499,N_4592,N_4604);
and UO_500 (O_500,N_4625,N_4730);
nor UO_501 (O_501,N_4844,N_4856);
or UO_502 (O_502,N_4644,N_4827);
nand UO_503 (O_503,N_4689,N_4912);
and UO_504 (O_504,N_4935,N_4823);
xor UO_505 (O_505,N_4986,N_4677);
xnor UO_506 (O_506,N_4501,N_4604);
and UO_507 (O_507,N_4618,N_4796);
nor UO_508 (O_508,N_4504,N_4646);
or UO_509 (O_509,N_4521,N_4720);
and UO_510 (O_510,N_4506,N_4525);
and UO_511 (O_511,N_4945,N_4974);
and UO_512 (O_512,N_4933,N_4856);
or UO_513 (O_513,N_4640,N_4762);
nand UO_514 (O_514,N_4989,N_4734);
nand UO_515 (O_515,N_4835,N_4847);
xor UO_516 (O_516,N_4830,N_4921);
and UO_517 (O_517,N_4799,N_4702);
nand UO_518 (O_518,N_4782,N_4694);
and UO_519 (O_519,N_4914,N_4703);
and UO_520 (O_520,N_4727,N_4684);
nor UO_521 (O_521,N_4594,N_4949);
or UO_522 (O_522,N_4859,N_4539);
and UO_523 (O_523,N_4511,N_4690);
and UO_524 (O_524,N_4965,N_4596);
xnor UO_525 (O_525,N_4681,N_4531);
nand UO_526 (O_526,N_4917,N_4832);
and UO_527 (O_527,N_4699,N_4669);
nor UO_528 (O_528,N_4973,N_4862);
nor UO_529 (O_529,N_4547,N_4985);
and UO_530 (O_530,N_4717,N_4736);
and UO_531 (O_531,N_4514,N_4671);
xor UO_532 (O_532,N_4823,N_4793);
nor UO_533 (O_533,N_4671,N_4847);
nand UO_534 (O_534,N_4997,N_4670);
nor UO_535 (O_535,N_4681,N_4933);
or UO_536 (O_536,N_4908,N_4882);
nand UO_537 (O_537,N_4596,N_4766);
nor UO_538 (O_538,N_4556,N_4637);
or UO_539 (O_539,N_4860,N_4877);
nor UO_540 (O_540,N_4948,N_4659);
nor UO_541 (O_541,N_4819,N_4656);
or UO_542 (O_542,N_4656,N_4603);
nor UO_543 (O_543,N_4687,N_4822);
xnor UO_544 (O_544,N_4763,N_4778);
and UO_545 (O_545,N_4979,N_4959);
nor UO_546 (O_546,N_4665,N_4630);
nor UO_547 (O_547,N_4874,N_4977);
nand UO_548 (O_548,N_4897,N_4542);
xnor UO_549 (O_549,N_4506,N_4787);
and UO_550 (O_550,N_4701,N_4623);
nor UO_551 (O_551,N_4569,N_4513);
nand UO_552 (O_552,N_4634,N_4597);
nor UO_553 (O_553,N_4778,N_4691);
xnor UO_554 (O_554,N_4561,N_4569);
nand UO_555 (O_555,N_4999,N_4763);
nand UO_556 (O_556,N_4574,N_4777);
or UO_557 (O_557,N_4665,N_4891);
and UO_558 (O_558,N_4775,N_4757);
nand UO_559 (O_559,N_4952,N_4847);
xor UO_560 (O_560,N_4700,N_4799);
or UO_561 (O_561,N_4571,N_4665);
xnor UO_562 (O_562,N_4546,N_4540);
or UO_563 (O_563,N_4819,N_4993);
or UO_564 (O_564,N_4919,N_4847);
nor UO_565 (O_565,N_4521,N_4762);
nand UO_566 (O_566,N_4869,N_4839);
xnor UO_567 (O_567,N_4999,N_4782);
nand UO_568 (O_568,N_4771,N_4741);
nor UO_569 (O_569,N_4544,N_4910);
nor UO_570 (O_570,N_4807,N_4683);
or UO_571 (O_571,N_4929,N_4956);
xnor UO_572 (O_572,N_4900,N_4646);
and UO_573 (O_573,N_4989,N_4513);
or UO_574 (O_574,N_4922,N_4965);
xnor UO_575 (O_575,N_4960,N_4796);
and UO_576 (O_576,N_4614,N_4960);
and UO_577 (O_577,N_4862,N_4943);
nand UO_578 (O_578,N_4611,N_4888);
or UO_579 (O_579,N_4760,N_4654);
nand UO_580 (O_580,N_4522,N_4583);
xnor UO_581 (O_581,N_4843,N_4580);
or UO_582 (O_582,N_4622,N_4995);
and UO_583 (O_583,N_4583,N_4721);
nor UO_584 (O_584,N_4794,N_4680);
or UO_585 (O_585,N_4586,N_4530);
nand UO_586 (O_586,N_4964,N_4830);
or UO_587 (O_587,N_4679,N_4589);
or UO_588 (O_588,N_4900,N_4621);
xnor UO_589 (O_589,N_4939,N_4543);
nor UO_590 (O_590,N_4716,N_4858);
xor UO_591 (O_591,N_4717,N_4568);
or UO_592 (O_592,N_4990,N_4723);
and UO_593 (O_593,N_4703,N_4919);
nand UO_594 (O_594,N_4589,N_4838);
nor UO_595 (O_595,N_4712,N_4993);
or UO_596 (O_596,N_4608,N_4584);
and UO_597 (O_597,N_4679,N_4594);
and UO_598 (O_598,N_4644,N_4542);
nor UO_599 (O_599,N_4561,N_4816);
xnor UO_600 (O_600,N_4734,N_4936);
or UO_601 (O_601,N_4570,N_4583);
nand UO_602 (O_602,N_4606,N_4692);
or UO_603 (O_603,N_4512,N_4984);
nor UO_604 (O_604,N_4623,N_4612);
and UO_605 (O_605,N_4691,N_4639);
or UO_606 (O_606,N_4806,N_4821);
or UO_607 (O_607,N_4803,N_4740);
nand UO_608 (O_608,N_4590,N_4955);
and UO_609 (O_609,N_4748,N_4983);
nand UO_610 (O_610,N_4903,N_4598);
nor UO_611 (O_611,N_4679,N_4922);
nand UO_612 (O_612,N_4931,N_4671);
nor UO_613 (O_613,N_4572,N_4599);
and UO_614 (O_614,N_4748,N_4980);
xnor UO_615 (O_615,N_4663,N_4619);
nor UO_616 (O_616,N_4688,N_4747);
or UO_617 (O_617,N_4948,N_4824);
and UO_618 (O_618,N_4574,N_4851);
or UO_619 (O_619,N_4737,N_4938);
and UO_620 (O_620,N_4705,N_4797);
xor UO_621 (O_621,N_4641,N_4563);
nand UO_622 (O_622,N_4865,N_4632);
and UO_623 (O_623,N_4781,N_4551);
nor UO_624 (O_624,N_4759,N_4593);
and UO_625 (O_625,N_4668,N_4741);
and UO_626 (O_626,N_4513,N_4898);
xnor UO_627 (O_627,N_4679,N_4841);
nor UO_628 (O_628,N_4677,N_4747);
xnor UO_629 (O_629,N_4868,N_4745);
xnor UO_630 (O_630,N_4505,N_4616);
and UO_631 (O_631,N_4744,N_4738);
and UO_632 (O_632,N_4965,N_4938);
and UO_633 (O_633,N_4604,N_4657);
nand UO_634 (O_634,N_4649,N_4879);
and UO_635 (O_635,N_4867,N_4982);
nor UO_636 (O_636,N_4825,N_4682);
and UO_637 (O_637,N_4826,N_4964);
or UO_638 (O_638,N_4721,N_4706);
and UO_639 (O_639,N_4502,N_4884);
xnor UO_640 (O_640,N_4822,N_4866);
nor UO_641 (O_641,N_4716,N_4651);
xor UO_642 (O_642,N_4553,N_4759);
and UO_643 (O_643,N_4561,N_4759);
xor UO_644 (O_644,N_4549,N_4744);
and UO_645 (O_645,N_4873,N_4783);
nand UO_646 (O_646,N_4519,N_4551);
xor UO_647 (O_647,N_4723,N_4526);
nand UO_648 (O_648,N_4558,N_4934);
nand UO_649 (O_649,N_4812,N_4827);
nand UO_650 (O_650,N_4618,N_4895);
or UO_651 (O_651,N_4929,N_4699);
or UO_652 (O_652,N_4646,N_4977);
nor UO_653 (O_653,N_4787,N_4965);
or UO_654 (O_654,N_4962,N_4521);
or UO_655 (O_655,N_4874,N_4821);
nand UO_656 (O_656,N_4751,N_4933);
or UO_657 (O_657,N_4961,N_4684);
and UO_658 (O_658,N_4620,N_4943);
nand UO_659 (O_659,N_4570,N_4838);
xnor UO_660 (O_660,N_4609,N_4740);
nand UO_661 (O_661,N_4939,N_4716);
xnor UO_662 (O_662,N_4877,N_4759);
and UO_663 (O_663,N_4530,N_4966);
nand UO_664 (O_664,N_4909,N_4584);
xor UO_665 (O_665,N_4539,N_4934);
nor UO_666 (O_666,N_4538,N_4957);
nor UO_667 (O_667,N_4944,N_4963);
nor UO_668 (O_668,N_4523,N_4795);
and UO_669 (O_669,N_4646,N_4946);
nand UO_670 (O_670,N_4678,N_4997);
nand UO_671 (O_671,N_4518,N_4714);
nor UO_672 (O_672,N_4778,N_4694);
and UO_673 (O_673,N_4727,N_4901);
nand UO_674 (O_674,N_4739,N_4599);
xnor UO_675 (O_675,N_4825,N_4967);
and UO_676 (O_676,N_4930,N_4515);
nor UO_677 (O_677,N_4899,N_4633);
nand UO_678 (O_678,N_4907,N_4948);
xor UO_679 (O_679,N_4756,N_4902);
or UO_680 (O_680,N_4556,N_4583);
or UO_681 (O_681,N_4813,N_4585);
nand UO_682 (O_682,N_4673,N_4835);
xnor UO_683 (O_683,N_4912,N_4930);
and UO_684 (O_684,N_4614,N_4580);
nor UO_685 (O_685,N_4561,N_4996);
and UO_686 (O_686,N_4819,N_4693);
nand UO_687 (O_687,N_4672,N_4526);
or UO_688 (O_688,N_4539,N_4922);
nand UO_689 (O_689,N_4867,N_4657);
or UO_690 (O_690,N_4636,N_4794);
and UO_691 (O_691,N_4518,N_4885);
xor UO_692 (O_692,N_4920,N_4763);
nor UO_693 (O_693,N_4577,N_4916);
xor UO_694 (O_694,N_4800,N_4572);
nand UO_695 (O_695,N_4927,N_4723);
and UO_696 (O_696,N_4759,N_4927);
nand UO_697 (O_697,N_4821,N_4556);
or UO_698 (O_698,N_4960,N_4759);
or UO_699 (O_699,N_4775,N_4694);
and UO_700 (O_700,N_4507,N_4576);
and UO_701 (O_701,N_4940,N_4567);
nor UO_702 (O_702,N_4931,N_4741);
nand UO_703 (O_703,N_4661,N_4969);
xor UO_704 (O_704,N_4936,N_4909);
nor UO_705 (O_705,N_4909,N_4841);
xor UO_706 (O_706,N_4881,N_4588);
and UO_707 (O_707,N_4659,N_4568);
xor UO_708 (O_708,N_4980,N_4710);
nor UO_709 (O_709,N_4782,N_4689);
nand UO_710 (O_710,N_4616,N_4983);
or UO_711 (O_711,N_4690,N_4628);
nand UO_712 (O_712,N_4540,N_4936);
and UO_713 (O_713,N_4502,N_4641);
or UO_714 (O_714,N_4919,N_4655);
or UO_715 (O_715,N_4664,N_4965);
and UO_716 (O_716,N_4691,N_4795);
nand UO_717 (O_717,N_4774,N_4600);
nor UO_718 (O_718,N_4922,N_4979);
or UO_719 (O_719,N_4760,N_4955);
nor UO_720 (O_720,N_4650,N_4871);
and UO_721 (O_721,N_4863,N_4815);
nor UO_722 (O_722,N_4510,N_4528);
nand UO_723 (O_723,N_4655,N_4941);
and UO_724 (O_724,N_4571,N_4701);
and UO_725 (O_725,N_4582,N_4857);
and UO_726 (O_726,N_4956,N_4611);
xnor UO_727 (O_727,N_4543,N_4634);
and UO_728 (O_728,N_4526,N_4804);
and UO_729 (O_729,N_4520,N_4731);
or UO_730 (O_730,N_4719,N_4610);
xor UO_731 (O_731,N_4912,N_4514);
nand UO_732 (O_732,N_4715,N_4538);
nor UO_733 (O_733,N_4650,N_4752);
xor UO_734 (O_734,N_4648,N_4941);
nor UO_735 (O_735,N_4906,N_4587);
and UO_736 (O_736,N_4683,N_4558);
nand UO_737 (O_737,N_4651,N_4759);
and UO_738 (O_738,N_4575,N_4507);
nor UO_739 (O_739,N_4869,N_4833);
xnor UO_740 (O_740,N_4622,N_4901);
nand UO_741 (O_741,N_4645,N_4787);
nand UO_742 (O_742,N_4798,N_4908);
or UO_743 (O_743,N_4570,N_4947);
nor UO_744 (O_744,N_4965,N_4509);
nand UO_745 (O_745,N_4995,N_4563);
nand UO_746 (O_746,N_4806,N_4880);
nand UO_747 (O_747,N_4595,N_4847);
and UO_748 (O_748,N_4822,N_4831);
nor UO_749 (O_749,N_4846,N_4785);
nor UO_750 (O_750,N_4507,N_4774);
nor UO_751 (O_751,N_4867,N_4741);
nand UO_752 (O_752,N_4727,N_4825);
nand UO_753 (O_753,N_4624,N_4761);
and UO_754 (O_754,N_4597,N_4969);
nand UO_755 (O_755,N_4605,N_4599);
or UO_756 (O_756,N_4727,N_4920);
or UO_757 (O_757,N_4513,N_4868);
and UO_758 (O_758,N_4525,N_4772);
xor UO_759 (O_759,N_4803,N_4648);
and UO_760 (O_760,N_4623,N_4620);
and UO_761 (O_761,N_4537,N_4943);
nand UO_762 (O_762,N_4645,N_4826);
xor UO_763 (O_763,N_4888,N_4787);
and UO_764 (O_764,N_4587,N_4828);
nor UO_765 (O_765,N_4677,N_4854);
xor UO_766 (O_766,N_4564,N_4695);
and UO_767 (O_767,N_4635,N_4823);
nor UO_768 (O_768,N_4815,N_4526);
or UO_769 (O_769,N_4574,N_4544);
or UO_770 (O_770,N_4611,N_4568);
xor UO_771 (O_771,N_4724,N_4617);
xor UO_772 (O_772,N_4701,N_4593);
or UO_773 (O_773,N_4531,N_4701);
xor UO_774 (O_774,N_4923,N_4686);
nor UO_775 (O_775,N_4871,N_4725);
xnor UO_776 (O_776,N_4775,N_4542);
and UO_777 (O_777,N_4611,N_4599);
and UO_778 (O_778,N_4744,N_4523);
nor UO_779 (O_779,N_4712,N_4500);
or UO_780 (O_780,N_4945,N_4797);
nand UO_781 (O_781,N_4783,N_4666);
xor UO_782 (O_782,N_4961,N_4749);
and UO_783 (O_783,N_4737,N_4788);
or UO_784 (O_784,N_4963,N_4723);
or UO_785 (O_785,N_4653,N_4682);
and UO_786 (O_786,N_4777,N_4562);
xnor UO_787 (O_787,N_4845,N_4534);
and UO_788 (O_788,N_4669,N_4767);
and UO_789 (O_789,N_4982,N_4918);
nor UO_790 (O_790,N_4600,N_4855);
nand UO_791 (O_791,N_4883,N_4833);
or UO_792 (O_792,N_4767,N_4795);
nor UO_793 (O_793,N_4700,N_4715);
and UO_794 (O_794,N_4953,N_4610);
and UO_795 (O_795,N_4705,N_4922);
xnor UO_796 (O_796,N_4611,N_4639);
xnor UO_797 (O_797,N_4858,N_4786);
nor UO_798 (O_798,N_4855,N_4637);
nand UO_799 (O_799,N_4931,N_4575);
nor UO_800 (O_800,N_4874,N_4819);
xor UO_801 (O_801,N_4716,N_4655);
or UO_802 (O_802,N_4527,N_4716);
nor UO_803 (O_803,N_4809,N_4540);
nor UO_804 (O_804,N_4662,N_4671);
nand UO_805 (O_805,N_4862,N_4572);
and UO_806 (O_806,N_4721,N_4700);
nor UO_807 (O_807,N_4835,N_4574);
and UO_808 (O_808,N_4621,N_4824);
and UO_809 (O_809,N_4764,N_4666);
xor UO_810 (O_810,N_4789,N_4685);
nand UO_811 (O_811,N_4930,N_4808);
xor UO_812 (O_812,N_4856,N_4940);
and UO_813 (O_813,N_4604,N_4737);
xnor UO_814 (O_814,N_4600,N_4781);
or UO_815 (O_815,N_4683,N_4889);
or UO_816 (O_816,N_4766,N_4758);
and UO_817 (O_817,N_4673,N_4886);
or UO_818 (O_818,N_4646,N_4986);
nor UO_819 (O_819,N_4631,N_4741);
nor UO_820 (O_820,N_4591,N_4964);
and UO_821 (O_821,N_4549,N_4800);
xnor UO_822 (O_822,N_4577,N_4898);
xor UO_823 (O_823,N_4936,N_4831);
and UO_824 (O_824,N_4532,N_4724);
xor UO_825 (O_825,N_4897,N_4908);
nor UO_826 (O_826,N_4524,N_4960);
or UO_827 (O_827,N_4982,N_4571);
and UO_828 (O_828,N_4980,N_4793);
nand UO_829 (O_829,N_4890,N_4884);
or UO_830 (O_830,N_4844,N_4961);
nand UO_831 (O_831,N_4959,N_4878);
or UO_832 (O_832,N_4968,N_4978);
or UO_833 (O_833,N_4687,N_4620);
nand UO_834 (O_834,N_4580,N_4648);
or UO_835 (O_835,N_4745,N_4915);
nand UO_836 (O_836,N_4529,N_4777);
and UO_837 (O_837,N_4506,N_4592);
xor UO_838 (O_838,N_4532,N_4845);
nand UO_839 (O_839,N_4792,N_4522);
nor UO_840 (O_840,N_4998,N_4754);
or UO_841 (O_841,N_4708,N_4988);
nor UO_842 (O_842,N_4527,N_4790);
nor UO_843 (O_843,N_4820,N_4855);
xnor UO_844 (O_844,N_4708,N_4715);
or UO_845 (O_845,N_4526,N_4915);
and UO_846 (O_846,N_4597,N_4681);
and UO_847 (O_847,N_4682,N_4603);
nand UO_848 (O_848,N_4756,N_4810);
xnor UO_849 (O_849,N_4811,N_4775);
nand UO_850 (O_850,N_4652,N_4749);
and UO_851 (O_851,N_4818,N_4569);
and UO_852 (O_852,N_4883,N_4764);
nand UO_853 (O_853,N_4938,N_4521);
or UO_854 (O_854,N_4521,N_4724);
and UO_855 (O_855,N_4679,N_4856);
or UO_856 (O_856,N_4535,N_4954);
nand UO_857 (O_857,N_4939,N_4907);
or UO_858 (O_858,N_4563,N_4960);
xnor UO_859 (O_859,N_4901,N_4528);
xor UO_860 (O_860,N_4725,N_4850);
and UO_861 (O_861,N_4799,N_4860);
xor UO_862 (O_862,N_4920,N_4818);
and UO_863 (O_863,N_4709,N_4619);
or UO_864 (O_864,N_4752,N_4881);
xnor UO_865 (O_865,N_4516,N_4861);
and UO_866 (O_866,N_4877,N_4843);
or UO_867 (O_867,N_4649,N_4788);
nand UO_868 (O_868,N_4728,N_4527);
nand UO_869 (O_869,N_4882,N_4844);
or UO_870 (O_870,N_4945,N_4899);
nand UO_871 (O_871,N_4810,N_4942);
nand UO_872 (O_872,N_4663,N_4649);
nor UO_873 (O_873,N_4866,N_4752);
nand UO_874 (O_874,N_4863,N_4559);
nor UO_875 (O_875,N_4846,N_4979);
nand UO_876 (O_876,N_4742,N_4748);
or UO_877 (O_877,N_4673,N_4545);
xnor UO_878 (O_878,N_4952,N_4541);
or UO_879 (O_879,N_4600,N_4685);
nand UO_880 (O_880,N_4610,N_4587);
nor UO_881 (O_881,N_4962,N_4828);
and UO_882 (O_882,N_4698,N_4563);
or UO_883 (O_883,N_4577,N_4513);
nor UO_884 (O_884,N_4979,N_4646);
nand UO_885 (O_885,N_4844,N_4920);
or UO_886 (O_886,N_4969,N_4608);
or UO_887 (O_887,N_4776,N_4556);
nor UO_888 (O_888,N_4799,N_4556);
nand UO_889 (O_889,N_4677,N_4998);
and UO_890 (O_890,N_4676,N_4542);
or UO_891 (O_891,N_4707,N_4972);
and UO_892 (O_892,N_4739,N_4987);
and UO_893 (O_893,N_4628,N_4984);
nand UO_894 (O_894,N_4867,N_4827);
nand UO_895 (O_895,N_4698,N_4634);
or UO_896 (O_896,N_4853,N_4880);
nand UO_897 (O_897,N_4876,N_4821);
and UO_898 (O_898,N_4888,N_4944);
xnor UO_899 (O_899,N_4592,N_4723);
nor UO_900 (O_900,N_4981,N_4609);
xnor UO_901 (O_901,N_4860,N_4588);
and UO_902 (O_902,N_4980,N_4663);
xnor UO_903 (O_903,N_4634,N_4941);
nor UO_904 (O_904,N_4692,N_4829);
nor UO_905 (O_905,N_4538,N_4831);
nand UO_906 (O_906,N_4579,N_4589);
nand UO_907 (O_907,N_4849,N_4937);
nor UO_908 (O_908,N_4872,N_4962);
nand UO_909 (O_909,N_4996,N_4649);
nor UO_910 (O_910,N_4983,N_4950);
nand UO_911 (O_911,N_4955,N_4528);
or UO_912 (O_912,N_4536,N_4672);
nand UO_913 (O_913,N_4537,N_4525);
nand UO_914 (O_914,N_4861,N_4757);
xnor UO_915 (O_915,N_4681,N_4502);
or UO_916 (O_916,N_4907,N_4760);
and UO_917 (O_917,N_4599,N_4853);
nand UO_918 (O_918,N_4894,N_4657);
xnor UO_919 (O_919,N_4678,N_4932);
xnor UO_920 (O_920,N_4991,N_4693);
xor UO_921 (O_921,N_4905,N_4786);
nor UO_922 (O_922,N_4682,N_4584);
or UO_923 (O_923,N_4706,N_4814);
or UO_924 (O_924,N_4796,N_4852);
or UO_925 (O_925,N_4673,N_4991);
xnor UO_926 (O_926,N_4682,N_4507);
or UO_927 (O_927,N_4682,N_4609);
nand UO_928 (O_928,N_4881,N_4645);
and UO_929 (O_929,N_4516,N_4877);
or UO_930 (O_930,N_4781,N_4816);
nand UO_931 (O_931,N_4927,N_4513);
nor UO_932 (O_932,N_4676,N_4710);
nand UO_933 (O_933,N_4583,N_4550);
or UO_934 (O_934,N_4638,N_4767);
nand UO_935 (O_935,N_4662,N_4869);
and UO_936 (O_936,N_4842,N_4548);
nor UO_937 (O_937,N_4778,N_4572);
nand UO_938 (O_938,N_4840,N_4809);
xor UO_939 (O_939,N_4853,N_4737);
nand UO_940 (O_940,N_4669,N_4892);
or UO_941 (O_941,N_4542,N_4752);
and UO_942 (O_942,N_4837,N_4799);
or UO_943 (O_943,N_4684,N_4769);
xor UO_944 (O_944,N_4816,N_4622);
or UO_945 (O_945,N_4906,N_4501);
xnor UO_946 (O_946,N_4521,N_4823);
or UO_947 (O_947,N_4852,N_4656);
nor UO_948 (O_948,N_4787,N_4842);
xor UO_949 (O_949,N_4789,N_4813);
and UO_950 (O_950,N_4733,N_4846);
nor UO_951 (O_951,N_4617,N_4884);
xnor UO_952 (O_952,N_4953,N_4688);
nand UO_953 (O_953,N_4876,N_4911);
xnor UO_954 (O_954,N_4910,N_4592);
nor UO_955 (O_955,N_4631,N_4624);
nor UO_956 (O_956,N_4921,N_4865);
and UO_957 (O_957,N_4658,N_4818);
nand UO_958 (O_958,N_4983,N_4714);
nor UO_959 (O_959,N_4833,N_4987);
nor UO_960 (O_960,N_4839,N_4954);
nand UO_961 (O_961,N_4596,N_4522);
and UO_962 (O_962,N_4610,N_4840);
and UO_963 (O_963,N_4956,N_4531);
nor UO_964 (O_964,N_4940,N_4790);
nor UO_965 (O_965,N_4736,N_4942);
and UO_966 (O_966,N_4807,N_4919);
xnor UO_967 (O_967,N_4626,N_4700);
xor UO_968 (O_968,N_4633,N_4612);
xnor UO_969 (O_969,N_4916,N_4636);
and UO_970 (O_970,N_4742,N_4919);
xor UO_971 (O_971,N_4607,N_4810);
nand UO_972 (O_972,N_4526,N_4622);
xor UO_973 (O_973,N_4815,N_4860);
and UO_974 (O_974,N_4562,N_4596);
nand UO_975 (O_975,N_4805,N_4818);
and UO_976 (O_976,N_4839,N_4775);
or UO_977 (O_977,N_4844,N_4944);
xor UO_978 (O_978,N_4716,N_4800);
xnor UO_979 (O_979,N_4749,N_4821);
xnor UO_980 (O_980,N_4798,N_4879);
nand UO_981 (O_981,N_4734,N_4922);
xor UO_982 (O_982,N_4519,N_4790);
nand UO_983 (O_983,N_4858,N_4979);
xnor UO_984 (O_984,N_4911,N_4820);
nor UO_985 (O_985,N_4995,N_4772);
and UO_986 (O_986,N_4987,N_4598);
and UO_987 (O_987,N_4972,N_4830);
or UO_988 (O_988,N_4967,N_4542);
or UO_989 (O_989,N_4896,N_4612);
xor UO_990 (O_990,N_4576,N_4899);
and UO_991 (O_991,N_4712,N_4818);
and UO_992 (O_992,N_4676,N_4721);
and UO_993 (O_993,N_4851,N_4861);
or UO_994 (O_994,N_4805,N_4910);
xor UO_995 (O_995,N_4814,N_4911);
and UO_996 (O_996,N_4515,N_4998);
or UO_997 (O_997,N_4541,N_4705);
xor UO_998 (O_998,N_4985,N_4895);
xor UO_999 (O_999,N_4723,N_4996);
endmodule