module basic_500_3000_500_40_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_166,In_108);
and U1 (N_1,In_268,In_201);
nor U2 (N_2,In_184,In_97);
nand U3 (N_3,In_156,In_98);
or U4 (N_4,In_180,In_139);
and U5 (N_5,In_222,In_418);
nor U6 (N_6,In_181,In_462);
nor U7 (N_7,In_404,In_35);
and U8 (N_8,In_147,In_173);
or U9 (N_9,In_131,In_17);
nor U10 (N_10,In_12,In_431);
or U11 (N_11,In_9,In_351);
xor U12 (N_12,In_46,In_22);
and U13 (N_13,In_286,In_157);
and U14 (N_14,In_423,In_132);
and U15 (N_15,In_379,In_49);
and U16 (N_16,In_323,In_373);
or U17 (N_17,In_187,In_270);
nand U18 (N_18,In_238,In_143);
or U19 (N_19,In_362,In_359);
nor U20 (N_20,In_249,In_440);
nor U21 (N_21,In_101,In_6);
nand U22 (N_22,In_39,In_37);
and U23 (N_23,In_344,In_412);
nand U24 (N_24,In_138,In_493);
nand U25 (N_25,In_290,In_172);
or U26 (N_26,In_305,In_488);
xnor U27 (N_27,In_83,In_482);
and U28 (N_28,In_319,In_189);
or U29 (N_29,In_244,In_289);
and U30 (N_30,In_198,In_356);
nand U31 (N_31,In_260,In_328);
and U32 (N_32,In_297,In_208);
and U33 (N_33,In_70,In_26);
or U34 (N_34,In_273,In_446);
and U35 (N_35,In_455,In_369);
nand U36 (N_36,In_408,In_27);
nand U37 (N_37,In_240,In_5);
nor U38 (N_38,In_76,In_69);
nor U39 (N_39,In_439,In_188);
and U40 (N_40,In_377,In_127);
and U41 (N_41,In_136,In_80);
nor U42 (N_42,In_428,In_56);
nand U43 (N_43,In_41,In_250);
and U44 (N_44,In_470,In_88);
nand U45 (N_45,In_153,In_186);
nor U46 (N_46,In_349,In_331);
or U47 (N_47,In_224,In_129);
nor U48 (N_48,In_341,In_196);
xor U49 (N_49,In_490,In_380);
nor U50 (N_50,In_275,In_242);
nand U51 (N_51,In_474,In_177);
or U52 (N_52,In_21,In_263);
and U53 (N_53,In_383,In_54);
nor U54 (N_54,In_77,In_61);
and U55 (N_55,In_32,In_480);
nand U56 (N_56,In_414,In_140);
or U57 (N_57,In_413,In_403);
nand U58 (N_58,In_481,In_499);
or U59 (N_59,In_287,In_178);
xnor U60 (N_60,In_384,In_265);
and U61 (N_61,In_151,In_416);
nor U62 (N_62,In_357,In_443);
and U63 (N_63,In_479,In_100);
or U64 (N_64,In_473,In_391);
nor U65 (N_65,In_134,In_469);
and U66 (N_66,In_426,In_303);
and U67 (N_67,In_355,In_133);
or U68 (N_68,In_92,In_272);
nor U69 (N_69,In_91,In_176);
or U70 (N_70,In_282,In_497);
or U71 (N_71,In_234,In_398);
nor U72 (N_72,In_407,In_29);
and U73 (N_73,In_336,In_230);
nor U74 (N_74,In_231,In_471);
nor U75 (N_75,In_78,In_121);
nand U76 (N_76,In_459,In_90);
xnor U77 (N_77,In_456,In_329);
and U78 (N_78,In_18,In_194);
xor U79 (N_79,In_294,In_28);
xor U80 (N_80,In_364,N_66);
nand U81 (N_81,In_45,N_36);
nor U82 (N_82,In_93,N_54);
and U83 (N_83,In_269,In_330);
and U84 (N_84,N_57,In_171);
or U85 (N_85,In_13,In_165);
nor U86 (N_86,In_245,In_71);
nand U87 (N_87,N_12,In_406);
and U88 (N_88,In_327,In_252);
nand U89 (N_89,In_55,N_41);
and U90 (N_90,N_50,In_421);
and U91 (N_91,In_74,In_203);
or U92 (N_92,In_333,In_210);
nor U93 (N_93,In_117,N_28);
nand U94 (N_94,In_409,In_448);
nor U95 (N_95,In_216,In_0);
or U96 (N_96,In_2,In_444);
nor U97 (N_97,In_338,In_454);
or U98 (N_98,In_4,In_253);
and U99 (N_99,In_266,In_307);
nor U100 (N_100,In_160,In_169);
nor U101 (N_101,In_126,In_255);
and U102 (N_102,In_25,N_1);
and U103 (N_103,In_343,In_417);
or U104 (N_104,In_42,N_10);
or U105 (N_105,In_113,In_79);
nor U106 (N_106,In_464,In_264);
and U107 (N_107,In_276,N_39);
nor U108 (N_108,In_386,N_60);
or U109 (N_109,In_461,In_144);
xnor U110 (N_110,In_168,In_288);
and U111 (N_111,In_109,In_472);
nor U112 (N_112,N_17,In_419);
nand U113 (N_113,In_450,In_368);
and U114 (N_114,N_27,In_422);
and U115 (N_115,In_484,N_30);
nand U116 (N_116,In_59,In_64);
nor U117 (N_117,In_67,In_382);
nor U118 (N_118,In_306,In_85);
nor U119 (N_119,In_424,In_281);
nor U120 (N_120,In_209,In_346);
and U121 (N_121,In_51,In_34);
and U122 (N_122,In_495,In_105);
nand U123 (N_123,In_436,N_63);
nand U124 (N_124,In_372,N_13);
or U125 (N_125,In_227,N_9);
nor U126 (N_126,In_430,In_309);
nand U127 (N_127,In_192,In_410);
nor U128 (N_128,In_396,N_73);
nand U129 (N_129,N_11,In_259);
nor U130 (N_130,N_22,In_63);
nor U131 (N_131,In_3,N_74);
xor U132 (N_132,In_123,In_58);
nor U133 (N_133,In_318,In_463);
and U134 (N_134,In_291,In_23);
or U135 (N_135,In_15,In_82);
nor U136 (N_136,In_314,In_442);
and U137 (N_137,In_47,In_261);
nand U138 (N_138,In_345,In_52);
xor U139 (N_139,In_256,N_59);
nand U140 (N_140,In_179,In_400);
nor U141 (N_141,In_411,In_283);
nor U142 (N_142,In_1,In_452);
nand U143 (N_143,In_483,In_441);
nor U144 (N_144,In_429,In_279);
nand U145 (N_145,In_44,N_25);
nor U146 (N_146,N_45,In_486);
nand U147 (N_147,N_15,In_228);
nor U148 (N_148,In_311,In_393);
and U149 (N_149,In_211,N_8);
nand U150 (N_150,In_220,In_243);
nor U151 (N_151,N_119,N_48);
nor U152 (N_152,In_326,N_145);
and U153 (N_153,N_42,In_223);
and U154 (N_154,In_280,In_350);
nor U155 (N_155,In_175,In_458);
or U156 (N_156,N_43,N_14);
xor U157 (N_157,In_376,In_233);
xnor U158 (N_158,In_150,In_370);
or U159 (N_159,In_267,In_313);
nor U160 (N_160,N_110,In_122);
and U161 (N_161,In_375,N_49);
and U162 (N_162,In_135,In_381);
nand U163 (N_163,In_30,In_366);
nor U164 (N_164,In_284,N_19);
or U165 (N_165,N_125,In_218);
nor U166 (N_166,N_26,In_427);
or U167 (N_167,In_425,In_207);
xnor U168 (N_168,N_148,In_137);
nor U169 (N_169,In_155,In_116);
or U170 (N_170,In_237,In_378);
xnor U171 (N_171,In_193,In_14);
nor U172 (N_172,In_434,N_94);
nand U173 (N_173,In_374,N_104);
and U174 (N_174,In_213,In_388);
or U175 (N_175,In_130,In_31);
nand U176 (N_176,In_317,In_212);
and U177 (N_177,In_8,In_229);
nand U178 (N_178,In_315,In_354);
and U179 (N_179,N_129,N_131);
nor U180 (N_180,N_118,In_183);
and U181 (N_181,N_114,In_262);
and U182 (N_182,N_52,In_164);
or U183 (N_183,In_361,In_73);
xnor U184 (N_184,N_128,In_225);
nor U185 (N_185,N_56,N_61);
or U186 (N_186,In_219,In_248);
nor U187 (N_187,N_64,N_32);
nand U188 (N_188,In_110,N_98);
nor U189 (N_189,N_72,In_271);
nor U190 (N_190,In_235,In_182);
nor U191 (N_191,In_204,In_112);
nor U192 (N_192,In_316,In_451);
nor U193 (N_193,N_137,N_149);
nand U194 (N_194,In_339,N_139);
or U195 (N_195,N_138,In_302);
nand U196 (N_196,N_134,N_99);
or U197 (N_197,In_390,In_353);
nand U198 (N_198,N_4,In_300);
nor U199 (N_199,N_2,In_399);
nor U200 (N_200,In_394,N_23);
nor U201 (N_201,N_126,In_293);
and U202 (N_202,In_437,In_498);
nor U203 (N_203,In_453,N_29);
or U204 (N_204,In_53,In_199);
and U205 (N_205,In_324,N_81);
or U206 (N_206,In_11,N_111);
nor U207 (N_207,In_205,N_21);
and U208 (N_208,N_3,In_174);
xor U209 (N_209,In_96,N_97);
and U210 (N_210,N_68,N_70);
nand U211 (N_211,In_72,N_55);
and U212 (N_212,In_40,In_371);
or U213 (N_213,In_94,N_143);
or U214 (N_214,In_236,N_16);
nor U215 (N_215,In_124,In_221);
xor U216 (N_216,In_66,N_102);
and U217 (N_217,In_487,N_121);
xor U218 (N_218,In_119,In_10);
nand U219 (N_219,In_494,In_445);
nand U220 (N_220,N_33,In_158);
nand U221 (N_221,N_35,N_46);
and U222 (N_222,In_241,In_114);
or U223 (N_223,In_33,N_130);
nor U224 (N_224,In_397,In_299);
or U225 (N_225,In_365,In_402);
nor U226 (N_226,N_216,N_38);
and U227 (N_227,In_466,In_360);
or U228 (N_228,N_62,In_467);
xor U229 (N_229,N_71,In_202);
nor U230 (N_230,N_193,N_188);
nor U231 (N_231,In_148,N_222);
nand U232 (N_232,In_478,In_87);
or U233 (N_233,In_340,In_460);
nor U234 (N_234,N_209,N_40);
nand U235 (N_235,N_132,N_106);
nand U236 (N_236,N_199,N_162);
and U237 (N_237,N_101,N_215);
nand U238 (N_238,In_57,In_154);
or U239 (N_239,N_163,N_108);
xnor U240 (N_240,N_208,N_167);
and U241 (N_241,In_48,N_88);
nor U242 (N_242,In_301,N_157);
xor U243 (N_243,N_77,N_47);
or U244 (N_244,N_133,N_24);
and U245 (N_245,In_332,N_158);
and U246 (N_246,N_197,N_83);
nor U247 (N_247,N_135,In_274);
or U248 (N_248,In_81,In_247);
nor U249 (N_249,N_58,In_468);
and U250 (N_250,N_85,In_489);
or U251 (N_251,N_142,N_152);
or U252 (N_252,In_239,N_200);
xor U253 (N_253,In_465,N_117);
nand U254 (N_254,N_212,N_224);
and U255 (N_255,N_173,N_184);
nor U256 (N_256,N_172,N_76);
nand U257 (N_257,N_5,N_164);
nand U258 (N_258,In_232,N_100);
or U259 (N_259,In_363,N_210);
and U260 (N_260,In_102,In_254);
or U261 (N_261,In_405,N_223);
nor U262 (N_262,In_62,N_107);
and U263 (N_263,N_204,N_218);
and U264 (N_264,In_167,In_145);
or U265 (N_265,In_257,In_195);
nand U266 (N_266,N_67,N_189);
nand U267 (N_267,In_348,In_107);
nor U268 (N_268,In_334,N_20);
or U269 (N_269,N_6,In_65);
and U270 (N_270,In_128,N_160);
or U271 (N_271,N_124,N_53);
nand U272 (N_272,N_120,In_75);
nand U273 (N_273,N_170,N_146);
xnor U274 (N_274,In_475,In_258);
nand U275 (N_275,N_37,N_206);
or U276 (N_276,In_214,N_79);
xor U277 (N_277,N_140,In_392);
nor U278 (N_278,N_155,N_177);
and U279 (N_279,In_120,N_169);
nor U280 (N_280,In_7,In_449);
nand U281 (N_281,In_352,In_387);
xnor U282 (N_282,N_214,In_99);
or U283 (N_283,In_50,N_191);
and U284 (N_284,In_310,N_51);
nand U285 (N_285,In_152,N_159);
and U286 (N_286,In_278,In_438);
or U287 (N_287,In_401,N_75);
nand U288 (N_288,N_84,In_197);
nand U289 (N_289,In_298,In_163);
nand U290 (N_290,In_335,In_125);
and U291 (N_291,N_203,In_420);
or U292 (N_292,In_367,In_20);
and U293 (N_293,In_86,In_325);
nor U294 (N_294,N_176,In_95);
nor U295 (N_295,In_292,In_476);
nand U296 (N_296,In_308,In_415);
nor U297 (N_297,N_165,In_60);
or U298 (N_298,N_185,N_221);
xnor U299 (N_299,N_90,N_198);
nor U300 (N_300,N_186,N_217);
or U301 (N_301,N_219,In_16);
xor U302 (N_302,N_194,N_274);
nor U303 (N_303,In_103,N_103);
and U304 (N_304,N_282,In_447);
or U305 (N_305,N_292,N_258);
xnor U306 (N_306,N_250,N_181);
or U307 (N_307,In_492,N_291);
nand U308 (N_308,N_231,N_243);
xor U309 (N_309,In_170,N_156);
nor U310 (N_310,N_82,In_496);
and U311 (N_311,N_254,In_43);
nand U312 (N_312,N_256,N_288);
nand U313 (N_313,In_395,N_248);
nand U314 (N_314,N_182,In_190);
and U315 (N_315,In_106,In_141);
xor U316 (N_316,N_205,N_244);
and U317 (N_317,N_272,N_211);
nor U318 (N_318,In_246,N_174);
nor U319 (N_319,N_78,In_24);
or U320 (N_320,N_136,N_230);
nor U321 (N_321,In_226,N_295);
nor U322 (N_322,N_150,N_252);
nor U323 (N_323,N_92,N_233);
nand U324 (N_324,N_275,N_96);
and U325 (N_325,In_36,N_290);
or U326 (N_326,In_491,N_262);
xor U327 (N_327,N_180,N_293);
xnor U328 (N_328,N_298,N_112);
nand U329 (N_329,N_178,In_84);
or U330 (N_330,N_69,N_80);
xnor U331 (N_331,N_278,N_123);
or U332 (N_332,N_257,In_295);
or U333 (N_333,N_227,In_191);
nor U334 (N_334,In_277,N_109);
or U335 (N_335,N_255,In_251);
nor U336 (N_336,N_179,In_477);
nand U337 (N_337,N_171,N_226);
or U338 (N_338,N_115,N_285);
nand U339 (N_339,N_277,N_202);
nand U340 (N_340,N_296,N_259);
and U341 (N_341,In_215,N_265);
nor U342 (N_342,N_213,N_151);
and U343 (N_343,In_389,In_457);
xor U344 (N_344,In_385,N_260);
and U345 (N_345,N_166,In_206);
nand U346 (N_346,N_236,In_217);
nor U347 (N_347,N_192,N_269);
or U348 (N_348,N_239,In_185);
nand U349 (N_349,N_105,N_116);
xor U350 (N_350,N_207,In_159);
or U351 (N_351,N_229,N_34);
or U352 (N_352,In_347,N_91);
nand U353 (N_353,In_111,N_65);
nor U354 (N_354,In_485,N_44);
or U355 (N_355,N_153,N_287);
xor U356 (N_356,N_232,N_201);
xor U357 (N_357,N_168,N_7);
xor U358 (N_358,N_113,N_261);
nand U359 (N_359,N_270,N_220);
or U360 (N_360,N_86,In_296);
and U361 (N_361,N_190,N_234);
nand U362 (N_362,N_228,N_299);
or U363 (N_363,N_18,N_183);
or U364 (N_364,In_200,In_285);
nor U365 (N_365,N_245,N_235);
and U366 (N_366,N_175,N_141);
xor U367 (N_367,In_162,In_358);
nor U368 (N_368,N_253,In_118);
nor U369 (N_369,In_322,In_142);
or U370 (N_370,N_284,N_246);
and U371 (N_371,N_283,In_115);
or U372 (N_372,N_297,In_68);
nand U373 (N_373,In_89,In_342);
xnor U374 (N_374,In_435,N_93);
nor U375 (N_375,In_146,N_353);
nor U376 (N_376,N_294,N_144);
nand U377 (N_377,N_360,N_334);
and U378 (N_378,N_331,N_315);
and U379 (N_379,N_301,N_325);
nand U380 (N_380,N_330,In_104);
and U381 (N_381,N_369,N_351);
nand U382 (N_382,N_271,In_432);
nor U383 (N_383,N_247,N_359);
xor U384 (N_384,N_361,N_241);
and U385 (N_385,N_238,N_347);
nand U386 (N_386,N_346,In_312);
and U387 (N_387,N_312,N_349);
or U388 (N_388,N_267,N_195);
and U389 (N_389,N_310,N_311);
and U390 (N_390,N_314,N_305);
nand U391 (N_391,N_161,N_249);
or U392 (N_392,N_280,N_87);
or U393 (N_393,N_340,N_300);
and U394 (N_394,N_317,N_342);
nor U395 (N_395,In_321,N_371);
or U396 (N_396,In_433,N_302);
nor U397 (N_397,N_276,N_313);
and U398 (N_398,N_316,N_122);
nand U399 (N_399,N_304,N_345);
nand U400 (N_400,N_89,N_251);
nor U401 (N_401,N_364,N_373);
nand U402 (N_402,N_95,In_304);
or U403 (N_403,In_337,N_268);
xor U404 (N_404,N_362,N_338);
xor U405 (N_405,N_273,N_327);
or U406 (N_406,N_367,N_365);
xor U407 (N_407,N_329,N_319);
or U408 (N_408,In_38,N_237);
nand U409 (N_409,N_242,N_321);
and U410 (N_410,N_154,N_147);
and U411 (N_411,N_324,N_343);
or U412 (N_412,N_368,N_320);
or U413 (N_413,N_344,N_350);
nor U414 (N_414,N_225,N_0);
nand U415 (N_415,N_348,N_354);
nor U416 (N_416,N_357,N_323);
nor U417 (N_417,N_341,N_322);
and U418 (N_418,N_303,N_374);
nand U419 (N_419,N_127,N_187);
and U420 (N_420,N_328,N_279);
nor U421 (N_421,N_196,N_264);
nand U422 (N_422,N_31,N_281);
or U423 (N_423,N_339,N_358);
nand U424 (N_424,In_161,N_240);
nor U425 (N_425,N_355,N_263);
or U426 (N_426,In_19,N_336);
nand U427 (N_427,N_370,N_366);
nand U428 (N_428,N_309,N_318);
nand U429 (N_429,N_372,N_335);
nand U430 (N_430,N_306,N_289);
nor U431 (N_431,N_266,N_326);
nand U432 (N_432,N_308,N_352);
nand U433 (N_433,N_337,N_332);
and U434 (N_434,In_320,N_286);
nor U435 (N_435,N_356,N_363);
nor U436 (N_436,In_149,N_307);
nand U437 (N_437,N_333,In_38);
or U438 (N_438,N_301,N_338);
or U439 (N_439,N_268,N_346);
and U440 (N_440,N_286,N_294);
xnor U441 (N_441,N_326,N_89);
and U442 (N_442,N_311,N_356);
xnor U443 (N_443,N_338,N_341);
nor U444 (N_444,N_249,N_374);
and U445 (N_445,In_433,N_307);
or U446 (N_446,In_19,N_266);
nand U447 (N_447,N_271,N_302);
and U448 (N_448,N_301,In_312);
nor U449 (N_449,N_322,N_373);
nor U450 (N_450,N_433,N_418);
xnor U451 (N_451,N_403,N_420);
or U452 (N_452,N_409,N_386);
nand U453 (N_453,N_377,N_427);
nand U454 (N_454,N_425,N_388);
nor U455 (N_455,N_439,N_379);
nand U456 (N_456,N_410,N_422);
xor U457 (N_457,N_405,N_390);
nor U458 (N_458,N_446,N_407);
nor U459 (N_459,N_441,N_429);
or U460 (N_460,N_414,N_415);
nand U461 (N_461,N_404,N_443);
nor U462 (N_462,N_445,N_381);
and U463 (N_463,N_448,N_394);
nor U464 (N_464,N_449,N_432);
and U465 (N_465,N_416,N_384);
nor U466 (N_466,N_376,N_401);
nand U467 (N_467,N_426,N_387);
or U468 (N_468,N_375,N_389);
and U469 (N_469,N_436,N_423);
nand U470 (N_470,N_391,N_392);
nand U471 (N_471,N_385,N_399);
xor U472 (N_472,N_434,N_442);
xnor U473 (N_473,N_419,N_437);
xor U474 (N_474,N_440,N_382);
or U475 (N_475,N_400,N_396);
nand U476 (N_476,N_424,N_395);
nor U477 (N_477,N_402,N_411);
and U478 (N_478,N_413,N_408);
or U479 (N_479,N_383,N_444);
xor U480 (N_480,N_431,N_435);
nor U481 (N_481,N_447,N_430);
and U482 (N_482,N_398,N_406);
nor U483 (N_483,N_378,N_412);
xor U484 (N_484,N_438,N_393);
or U485 (N_485,N_428,N_421);
nor U486 (N_486,N_397,N_380);
and U487 (N_487,N_417,N_449);
or U488 (N_488,N_447,N_444);
or U489 (N_489,N_388,N_395);
and U490 (N_490,N_389,N_434);
nor U491 (N_491,N_414,N_447);
xor U492 (N_492,N_436,N_406);
xor U493 (N_493,N_376,N_408);
or U494 (N_494,N_391,N_403);
or U495 (N_495,N_439,N_418);
and U496 (N_496,N_375,N_419);
or U497 (N_497,N_414,N_430);
nor U498 (N_498,N_418,N_386);
or U499 (N_499,N_420,N_395);
and U500 (N_500,N_419,N_382);
nor U501 (N_501,N_398,N_437);
nor U502 (N_502,N_424,N_430);
or U503 (N_503,N_413,N_400);
xnor U504 (N_504,N_447,N_393);
and U505 (N_505,N_383,N_395);
and U506 (N_506,N_380,N_409);
nand U507 (N_507,N_441,N_426);
and U508 (N_508,N_446,N_430);
or U509 (N_509,N_405,N_375);
nand U510 (N_510,N_399,N_448);
nand U511 (N_511,N_433,N_421);
and U512 (N_512,N_390,N_380);
nor U513 (N_513,N_418,N_399);
nor U514 (N_514,N_427,N_398);
nor U515 (N_515,N_377,N_392);
xnor U516 (N_516,N_392,N_400);
xor U517 (N_517,N_421,N_402);
and U518 (N_518,N_448,N_389);
nand U519 (N_519,N_384,N_381);
nor U520 (N_520,N_437,N_392);
nand U521 (N_521,N_420,N_394);
and U522 (N_522,N_442,N_415);
nand U523 (N_523,N_411,N_406);
nand U524 (N_524,N_378,N_441);
nand U525 (N_525,N_463,N_453);
nand U526 (N_526,N_501,N_510);
or U527 (N_527,N_496,N_483);
and U528 (N_528,N_475,N_450);
nor U529 (N_529,N_519,N_478);
or U530 (N_530,N_469,N_459);
and U531 (N_531,N_502,N_476);
nor U532 (N_532,N_461,N_488);
or U533 (N_533,N_456,N_486);
nor U534 (N_534,N_523,N_470);
xor U535 (N_535,N_507,N_451);
nand U536 (N_536,N_506,N_460);
or U537 (N_537,N_489,N_513);
and U538 (N_538,N_514,N_458);
nand U539 (N_539,N_467,N_454);
and U540 (N_540,N_521,N_484);
and U541 (N_541,N_493,N_500);
nor U542 (N_542,N_487,N_464);
or U543 (N_543,N_495,N_452);
and U544 (N_544,N_499,N_472);
nand U545 (N_545,N_474,N_512);
and U546 (N_546,N_462,N_522);
and U547 (N_547,N_508,N_511);
nor U548 (N_548,N_457,N_491);
nor U549 (N_549,N_492,N_517);
and U550 (N_550,N_490,N_479);
nand U551 (N_551,N_515,N_455);
and U552 (N_552,N_473,N_481);
nor U553 (N_553,N_509,N_516);
nand U554 (N_554,N_503,N_518);
nor U555 (N_555,N_498,N_466);
and U556 (N_556,N_477,N_505);
nor U557 (N_557,N_482,N_524);
nand U558 (N_558,N_468,N_480);
and U559 (N_559,N_497,N_494);
nand U560 (N_560,N_465,N_471);
xor U561 (N_561,N_504,N_520);
or U562 (N_562,N_485,N_495);
and U563 (N_563,N_491,N_514);
or U564 (N_564,N_500,N_522);
nand U565 (N_565,N_495,N_450);
or U566 (N_566,N_451,N_498);
nor U567 (N_567,N_499,N_515);
or U568 (N_568,N_468,N_496);
or U569 (N_569,N_477,N_494);
and U570 (N_570,N_514,N_464);
nor U571 (N_571,N_457,N_465);
and U572 (N_572,N_508,N_510);
nor U573 (N_573,N_479,N_519);
or U574 (N_574,N_495,N_497);
and U575 (N_575,N_483,N_452);
nand U576 (N_576,N_470,N_498);
nand U577 (N_577,N_516,N_453);
or U578 (N_578,N_458,N_493);
and U579 (N_579,N_464,N_513);
or U580 (N_580,N_501,N_478);
or U581 (N_581,N_459,N_519);
nand U582 (N_582,N_483,N_509);
or U583 (N_583,N_450,N_488);
nor U584 (N_584,N_489,N_500);
and U585 (N_585,N_514,N_452);
or U586 (N_586,N_462,N_466);
nor U587 (N_587,N_479,N_476);
or U588 (N_588,N_464,N_484);
nor U589 (N_589,N_462,N_451);
nor U590 (N_590,N_497,N_460);
or U591 (N_591,N_498,N_501);
and U592 (N_592,N_488,N_456);
or U593 (N_593,N_521,N_469);
nor U594 (N_594,N_476,N_467);
nand U595 (N_595,N_509,N_510);
nor U596 (N_596,N_467,N_453);
nand U597 (N_597,N_466,N_501);
and U598 (N_598,N_494,N_500);
nor U599 (N_599,N_507,N_489);
nand U600 (N_600,N_599,N_567);
xor U601 (N_601,N_533,N_595);
nor U602 (N_602,N_525,N_553);
nand U603 (N_603,N_527,N_584);
and U604 (N_604,N_528,N_540);
and U605 (N_605,N_530,N_559);
xnor U606 (N_606,N_562,N_588);
nor U607 (N_607,N_556,N_591);
nand U608 (N_608,N_538,N_572);
or U609 (N_609,N_593,N_543);
and U610 (N_610,N_571,N_592);
nand U611 (N_611,N_585,N_526);
or U612 (N_612,N_575,N_544);
nand U613 (N_613,N_576,N_581);
xor U614 (N_614,N_555,N_549);
nand U615 (N_615,N_577,N_596);
and U616 (N_616,N_594,N_529);
nand U617 (N_617,N_552,N_563);
nand U618 (N_618,N_574,N_548);
nor U619 (N_619,N_546,N_586);
xnor U620 (N_620,N_551,N_557);
or U621 (N_621,N_598,N_582);
or U622 (N_622,N_535,N_573);
xnor U623 (N_623,N_554,N_589);
or U624 (N_624,N_565,N_560);
nor U625 (N_625,N_570,N_541);
nor U626 (N_626,N_587,N_583);
nand U627 (N_627,N_568,N_545);
xnor U628 (N_628,N_534,N_537);
nand U629 (N_629,N_542,N_536);
and U630 (N_630,N_579,N_569);
and U631 (N_631,N_547,N_564);
or U632 (N_632,N_561,N_590);
nor U633 (N_633,N_566,N_580);
xor U634 (N_634,N_531,N_539);
nor U635 (N_635,N_597,N_532);
nor U636 (N_636,N_558,N_578);
or U637 (N_637,N_550,N_594);
or U638 (N_638,N_594,N_599);
and U639 (N_639,N_528,N_574);
nor U640 (N_640,N_528,N_568);
nor U641 (N_641,N_586,N_570);
or U642 (N_642,N_531,N_526);
xnor U643 (N_643,N_588,N_540);
nand U644 (N_644,N_555,N_594);
or U645 (N_645,N_596,N_590);
or U646 (N_646,N_564,N_561);
nand U647 (N_647,N_535,N_527);
nor U648 (N_648,N_565,N_538);
or U649 (N_649,N_550,N_595);
xor U650 (N_650,N_530,N_528);
and U651 (N_651,N_533,N_543);
or U652 (N_652,N_536,N_580);
and U653 (N_653,N_568,N_576);
and U654 (N_654,N_554,N_566);
nand U655 (N_655,N_540,N_577);
and U656 (N_656,N_554,N_526);
or U657 (N_657,N_598,N_540);
nor U658 (N_658,N_557,N_534);
or U659 (N_659,N_593,N_528);
nor U660 (N_660,N_589,N_541);
and U661 (N_661,N_578,N_572);
xnor U662 (N_662,N_534,N_577);
or U663 (N_663,N_581,N_556);
and U664 (N_664,N_534,N_595);
and U665 (N_665,N_593,N_557);
and U666 (N_666,N_575,N_545);
or U667 (N_667,N_587,N_564);
nand U668 (N_668,N_543,N_564);
nor U669 (N_669,N_580,N_585);
or U670 (N_670,N_526,N_596);
xor U671 (N_671,N_526,N_542);
xor U672 (N_672,N_588,N_539);
nor U673 (N_673,N_542,N_580);
and U674 (N_674,N_528,N_565);
and U675 (N_675,N_652,N_643);
and U676 (N_676,N_668,N_632);
or U677 (N_677,N_631,N_618);
nand U678 (N_678,N_674,N_663);
nor U679 (N_679,N_612,N_650);
or U680 (N_680,N_667,N_646);
or U681 (N_681,N_623,N_655);
nor U682 (N_682,N_624,N_651);
and U683 (N_683,N_630,N_607);
nand U684 (N_684,N_640,N_641);
or U685 (N_685,N_638,N_659);
nor U686 (N_686,N_637,N_614);
nor U687 (N_687,N_647,N_610);
and U688 (N_688,N_657,N_629);
nand U689 (N_689,N_639,N_673);
nor U690 (N_690,N_665,N_661);
or U691 (N_691,N_649,N_625);
or U692 (N_692,N_669,N_613);
and U693 (N_693,N_648,N_662);
nor U694 (N_694,N_670,N_616);
or U695 (N_695,N_666,N_656);
xnor U696 (N_696,N_654,N_615);
and U697 (N_697,N_617,N_627);
nand U698 (N_698,N_626,N_619);
or U699 (N_699,N_609,N_644);
xnor U700 (N_700,N_622,N_634);
nand U701 (N_701,N_608,N_606);
and U702 (N_702,N_602,N_645);
xnor U703 (N_703,N_611,N_664);
xor U704 (N_704,N_600,N_633);
nand U705 (N_705,N_603,N_636);
nand U706 (N_706,N_672,N_660);
or U707 (N_707,N_635,N_621);
nor U708 (N_708,N_642,N_671);
nor U709 (N_709,N_620,N_604);
and U710 (N_710,N_628,N_601);
nand U711 (N_711,N_605,N_658);
nand U712 (N_712,N_653,N_672);
nand U713 (N_713,N_618,N_647);
and U714 (N_714,N_606,N_612);
and U715 (N_715,N_625,N_634);
or U716 (N_716,N_610,N_644);
nor U717 (N_717,N_661,N_663);
nor U718 (N_718,N_645,N_611);
nand U719 (N_719,N_605,N_611);
nand U720 (N_720,N_640,N_648);
and U721 (N_721,N_635,N_663);
and U722 (N_722,N_611,N_673);
xor U723 (N_723,N_632,N_639);
nor U724 (N_724,N_609,N_646);
nor U725 (N_725,N_600,N_617);
nor U726 (N_726,N_639,N_614);
xor U727 (N_727,N_672,N_602);
nor U728 (N_728,N_638,N_655);
and U729 (N_729,N_634,N_645);
and U730 (N_730,N_626,N_662);
or U731 (N_731,N_606,N_613);
nor U732 (N_732,N_626,N_630);
nand U733 (N_733,N_623,N_604);
and U734 (N_734,N_608,N_640);
and U735 (N_735,N_661,N_664);
and U736 (N_736,N_629,N_612);
or U737 (N_737,N_642,N_622);
or U738 (N_738,N_665,N_647);
nand U739 (N_739,N_641,N_630);
and U740 (N_740,N_670,N_629);
nor U741 (N_741,N_636,N_673);
nor U742 (N_742,N_611,N_665);
nor U743 (N_743,N_655,N_659);
nand U744 (N_744,N_661,N_609);
or U745 (N_745,N_600,N_631);
nand U746 (N_746,N_624,N_671);
nor U747 (N_747,N_672,N_667);
nor U748 (N_748,N_613,N_665);
or U749 (N_749,N_658,N_645);
nor U750 (N_750,N_680,N_683);
and U751 (N_751,N_738,N_720);
or U752 (N_752,N_719,N_749);
nand U753 (N_753,N_731,N_684);
and U754 (N_754,N_708,N_705);
or U755 (N_755,N_743,N_695);
nor U756 (N_756,N_682,N_677);
nor U757 (N_757,N_740,N_716);
nor U758 (N_758,N_748,N_676);
nand U759 (N_759,N_739,N_694);
or U760 (N_760,N_706,N_686);
and U761 (N_761,N_692,N_712);
and U762 (N_762,N_744,N_687);
or U763 (N_763,N_729,N_734);
or U764 (N_764,N_714,N_723);
and U765 (N_765,N_698,N_715);
nand U766 (N_766,N_681,N_691);
and U767 (N_767,N_747,N_710);
nor U768 (N_768,N_718,N_726);
nand U769 (N_769,N_737,N_697);
xor U770 (N_770,N_733,N_713);
and U771 (N_771,N_741,N_688);
or U772 (N_772,N_730,N_717);
and U773 (N_773,N_735,N_742);
nand U774 (N_774,N_722,N_703);
nor U775 (N_775,N_693,N_701);
nor U776 (N_776,N_699,N_707);
nand U777 (N_777,N_702,N_704);
or U778 (N_778,N_727,N_685);
xnor U779 (N_779,N_678,N_746);
or U780 (N_780,N_732,N_689);
nand U781 (N_781,N_711,N_725);
xnor U782 (N_782,N_724,N_709);
or U783 (N_783,N_728,N_696);
nor U784 (N_784,N_745,N_679);
nor U785 (N_785,N_700,N_690);
and U786 (N_786,N_736,N_675);
nor U787 (N_787,N_721,N_693);
nor U788 (N_788,N_690,N_724);
or U789 (N_789,N_727,N_747);
and U790 (N_790,N_729,N_689);
nand U791 (N_791,N_744,N_730);
or U792 (N_792,N_699,N_735);
or U793 (N_793,N_685,N_706);
or U794 (N_794,N_733,N_690);
nor U795 (N_795,N_677,N_693);
and U796 (N_796,N_703,N_715);
nand U797 (N_797,N_698,N_690);
and U798 (N_798,N_728,N_733);
nand U799 (N_799,N_720,N_702);
and U800 (N_800,N_739,N_727);
nand U801 (N_801,N_739,N_692);
and U802 (N_802,N_737,N_695);
nand U803 (N_803,N_736,N_725);
and U804 (N_804,N_726,N_678);
nor U805 (N_805,N_737,N_717);
nor U806 (N_806,N_700,N_677);
or U807 (N_807,N_706,N_682);
or U808 (N_808,N_703,N_692);
or U809 (N_809,N_679,N_719);
nand U810 (N_810,N_708,N_702);
or U811 (N_811,N_709,N_723);
and U812 (N_812,N_712,N_720);
and U813 (N_813,N_714,N_685);
and U814 (N_814,N_684,N_739);
nand U815 (N_815,N_701,N_733);
and U816 (N_816,N_747,N_741);
and U817 (N_817,N_683,N_728);
nand U818 (N_818,N_703,N_729);
nor U819 (N_819,N_696,N_683);
nor U820 (N_820,N_679,N_689);
and U821 (N_821,N_730,N_686);
nor U822 (N_822,N_737,N_675);
xor U823 (N_823,N_693,N_746);
or U824 (N_824,N_716,N_691);
nor U825 (N_825,N_807,N_763);
xor U826 (N_826,N_823,N_773);
or U827 (N_827,N_755,N_810);
and U828 (N_828,N_776,N_811);
nand U829 (N_829,N_791,N_790);
nand U830 (N_830,N_818,N_789);
nor U831 (N_831,N_782,N_822);
nor U832 (N_832,N_805,N_774);
nor U833 (N_833,N_783,N_767);
nand U834 (N_834,N_754,N_815);
nand U835 (N_835,N_799,N_778);
nor U836 (N_836,N_766,N_784);
nand U837 (N_837,N_806,N_813);
nand U838 (N_838,N_758,N_824);
nand U839 (N_839,N_801,N_772);
or U840 (N_840,N_779,N_777);
nand U841 (N_841,N_808,N_794);
nor U842 (N_842,N_765,N_786);
nand U843 (N_843,N_800,N_792);
nand U844 (N_844,N_787,N_757);
and U845 (N_845,N_788,N_753);
nand U846 (N_846,N_769,N_798);
nor U847 (N_847,N_804,N_796);
xor U848 (N_848,N_759,N_816);
and U849 (N_849,N_817,N_780);
nand U850 (N_850,N_761,N_814);
nor U851 (N_851,N_751,N_762);
and U852 (N_852,N_793,N_821);
nand U853 (N_853,N_768,N_764);
nand U854 (N_854,N_812,N_775);
or U855 (N_855,N_819,N_785);
or U856 (N_856,N_809,N_771);
xnor U857 (N_857,N_803,N_756);
or U858 (N_858,N_797,N_795);
and U859 (N_859,N_760,N_802);
nor U860 (N_860,N_820,N_770);
nand U861 (N_861,N_752,N_781);
nand U862 (N_862,N_750,N_800);
nor U863 (N_863,N_794,N_757);
nand U864 (N_864,N_817,N_818);
or U865 (N_865,N_782,N_781);
nor U866 (N_866,N_758,N_764);
nand U867 (N_867,N_756,N_813);
or U868 (N_868,N_763,N_794);
or U869 (N_869,N_807,N_781);
and U870 (N_870,N_752,N_816);
or U871 (N_871,N_752,N_803);
or U872 (N_872,N_811,N_805);
nor U873 (N_873,N_767,N_751);
and U874 (N_874,N_798,N_771);
or U875 (N_875,N_792,N_816);
and U876 (N_876,N_820,N_786);
or U877 (N_877,N_803,N_783);
nor U878 (N_878,N_817,N_808);
or U879 (N_879,N_824,N_794);
nor U880 (N_880,N_763,N_796);
or U881 (N_881,N_801,N_787);
or U882 (N_882,N_820,N_785);
nor U883 (N_883,N_770,N_794);
and U884 (N_884,N_772,N_812);
nor U885 (N_885,N_806,N_809);
or U886 (N_886,N_815,N_773);
nand U887 (N_887,N_753,N_759);
xnor U888 (N_888,N_813,N_761);
nand U889 (N_889,N_812,N_782);
nand U890 (N_890,N_820,N_783);
xnor U891 (N_891,N_798,N_804);
nand U892 (N_892,N_781,N_817);
nand U893 (N_893,N_767,N_752);
xnor U894 (N_894,N_788,N_771);
and U895 (N_895,N_759,N_812);
nor U896 (N_896,N_762,N_780);
nand U897 (N_897,N_789,N_777);
and U898 (N_898,N_762,N_764);
nor U899 (N_899,N_769,N_772);
nand U900 (N_900,N_854,N_836);
nand U901 (N_901,N_842,N_864);
nor U902 (N_902,N_858,N_862);
and U903 (N_903,N_868,N_885);
or U904 (N_904,N_889,N_883);
and U905 (N_905,N_869,N_870);
and U906 (N_906,N_857,N_832);
or U907 (N_907,N_880,N_899);
nand U908 (N_908,N_837,N_866);
and U909 (N_909,N_888,N_873);
nand U910 (N_910,N_860,N_881);
nand U911 (N_911,N_846,N_859);
or U912 (N_912,N_896,N_827);
and U913 (N_913,N_876,N_871);
nor U914 (N_914,N_845,N_894);
nor U915 (N_915,N_825,N_863);
or U916 (N_916,N_892,N_848);
and U917 (N_917,N_872,N_831);
nor U918 (N_918,N_877,N_884);
or U919 (N_919,N_826,N_887);
or U920 (N_920,N_879,N_838);
xnor U921 (N_921,N_875,N_841);
or U922 (N_922,N_893,N_829);
or U923 (N_923,N_897,N_874);
or U924 (N_924,N_853,N_886);
and U925 (N_925,N_891,N_851);
nor U926 (N_926,N_834,N_833);
or U927 (N_927,N_839,N_856);
and U928 (N_928,N_852,N_890);
nand U929 (N_929,N_855,N_850);
nor U930 (N_930,N_849,N_895);
or U931 (N_931,N_843,N_882);
nand U932 (N_932,N_867,N_878);
nand U933 (N_933,N_830,N_865);
nand U934 (N_934,N_844,N_835);
and U935 (N_935,N_898,N_847);
and U936 (N_936,N_828,N_840);
nand U937 (N_937,N_861,N_850);
and U938 (N_938,N_890,N_858);
nor U939 (N_939,N_869,N_873);
nor U940 (N_940,N_845,N_852);
or U941 (N_941,N_841,N_894);
and U942 (N_942,N_861,N_897);
xnor U943 (N_943,N_838,N_833);
nor U944 (N_944,N_887,N_880);
and U945 (N_945,N_895,N_872);
or U946 (N_946,N_869,N_896);
nor U947 (N_947,N_883,N_859);
nand U948 (N_948,N_861,N_867);
and U949 (N_949,N_894,N_860);
nor U950 (N_950,N_890,N_869);
nand U951 (N_951,N_838,N_887);
xor U952 (N_952,N_869,N_876);
nand U953 (N_953,N_870,N_868);
and U954 (N_954,N_855,N_889);
nand U955 (N_955,N_847,N_846);
and U956 (N_956,N_861,N_869);
xnor U957 (N_957,N_837,N_845);
nor U958 (N_958,N_861,N_827);
nand U959 (N_959,N_880,N_893);
nor U960 (N_960,N_866,N_826);
and U961 (N_961,N_885,N_846);
nor U962 (N_962,N_839,N_847);
and U963 (N_963,N_873,N_871);
or U964 (N_964,N_846,N_843);
nand U965 (N_965,N_875,N_867);
nand U966 (N_966,N_845,N_879);
and U967 (N_967,N_891,N_880);
and U968 (N_968,N_882,N_835);
nand U969 (N_969,N_863,N_856);
or U970 (N_970,N_881,N_846);
and U971 (N_971,N_831,N_898);
and U972 (N_972,N_851,N_831);
or U973 (N_973,N_893,N_877);
and U974 (N_974,N_872,N_843);
or U975 (N_975,N_917,N_910);
and U976 (N_976,N_924,N_947);
or U977 (N_977,N_931,N_938);
or U978 (N_978,N_957,N_961);
and U979 (N_979,N_912,N_939);
nor U980 (N_980,N_902,N_950);
nand U981 (N_981,N_905,N_964);
nor U982 (N_982,N_965,N_941);
nor U983 (N_983,N_937,N_942);
or U984 (N_984,N_955,N_932);
or U985 (N_985,N_935,N_946);
or U986 (N_986,N_956,N_900);
or U987 (N_987,N_913,N_968);
nor U988 (N_988,N_934,N_908);
nand U989 (N_989,N_901,N_970);
nand U990 (N_990,N_930,N_945);
and U991 (N_991,N_943,N_922);
nor U992 (N_992,N_958,N_918);
and U993 (N_993,N_944,N_904);
or U994 (N_994,N_966,N_909);
or U995 (N_995,N_952,N_903);
and U996 (N_996,N_925,N_907);
nor U997 (N_997,N_921,N_940);
nand U998 (N_998,N_928,N_916);
nor U999 (N_999,N_963,N_919);
nand U1000 (N_1000,N_927,N_972);
or U1001 (N_1001,N_920,N_936);
nand U1002 (N_1002,N_969,N_960);
and U1003 (N_1003,N_929,N_949);
nand U1004 (N_1004,N_962,N_923);
or U1005 (N_1005,N_954,N_926);
or U1006 (N_1006,N_951,N_906);
nor U1007 (N_1007,N_914,N_974);
xnor U1008 (N_1008,N_915,N_911);
or U1009 (N_1009,N_973,N_959);
or U1010 (N_1010,N_933,N_967);
nor U1011 (N_1011,N_948,N_971);
nor U1012 (N_1012,N_953,N_911);
nor U1013 (N_1013,N_929,N_931);
nand U1014 (N_1014,N_938,N_958);
and U1015 (N_1015,N_904,N_960);
and U1016 (N_1016,N_932,N_971);
or U1017 (N_1017,N_906,N_902);
nand U1018 (N_1018,N_922,N_934);
or U1019 (N_1019,N_949,N_939);
nor U1020 (N_1020,N_973,N_944);
nand U1021 (N_1021,N_916,N_941);
and U1022 (N_1022,N_970,N_929);
xnor U1023 (N_1023,N_926,N_953);
or U1024 (N_1024,N_955,N_909);
or U1025 (N_1025,N_951,N_910);
or U1026 (N_1026,N_958,N_914);
nor U1027 (N_1027,N_954,N_965);
xor U1028 (N_1028,N_968,N_972);
xor U1029 (N_1029,N_964,N_917);
nand U1030 (N_1030,N_958,N_972);
nand U1031 (N_1031,N_922,N_939);
or U1032 (N_1032,N_961,N_938);
and U1033 (N_1033,N_905,N_902);
and U1034 (N_1034,N_946,N_937);
and U1035 (N_1035,N_943,N_963);
nand U1036 (N_1036,N_900,N_906);
nand U1037 (N_1037,N_943,N_927);
and U1038 (N_1038,N_937,N_972);
or U1039 (N_1039,N_967,N_973);
nor U1040 (N_1040,N_945,N_915);
nand U1041 (N_1041,N_933,N_901);
nand U1042 (N_1042,N_925,N_957);
and U1043 (N_1043,N_953,N_900);
nor U1044 (N_1044,N_940,N_938);
xor U1045 (N_1045,N_921,N_938);
nor U1046 (N_1046,N_900,N_950);
nand U1047 (N_1047,N_952,N_936);
nor U1048 (N_1048,N_924,N_956);
or U1049 (N_1049,N_901,N_946);
nor U1050 (N_1050,N_998,N_983);
xnor U1051 (N_1051,N_1048,N_991);
or U1052 (N_1052,N_1013,N_1021);
nand U1053 (N_1053,N_997,N_1004);
nand U1054 (N_1054,N_989,N_1027);
nand U1055 (N_1055,N_1025,N_1000);
and U1056 (N_1056,N_1035,N_1003);
or U1057 (N_1057,N_1045,N_978);
nor U1058 (N_1058,N_981,N_1010);
or U1059 (N_1059,N_1023,N_1037);
nand U1060 (N_1060,N_1002,N_977);
nor U1061 (N_1061,N_988,N_994);
nor U1062 (N_1062,N_1047,N_1028);
and U1063 (N_1063,N_1014,N_1030);
nand U1064 (N_1064,N_975,N_992);
and U1065 (N_1065,N_1009,N_1017);
nor U1066 (N_1066,N_1032,N_1006);
nor U1067 (N_1067,N_980,N_984);
or U1068 (N_1068,N_1036,N_987);
and U1069 (N_1069,N_1007,N_1034);
and U1070 (N_1070,N_1031,N_1044);
and U1071 (N_1071,N_1040,N_979);
nand U1072 (N_1072,N_1016,N_1042);
nor U1073 (N_1073,N_1005,N_1026);
xor U1074 (N_1074,N_995,N_993);
or U1075 (N_1075,N_976,N_1019);
nand U1076 (N_1076,N_1015,N_1043);
or U1077 (N_1077,N_1039,N_1033);
xor U1078 (N_1078,N_1046,N_1029);
nor U1079 (N_1079,N_990,N_1049);
nand U1080 (N_1080,N_996,N_1041);
nor U1081 (N_1081,N_982,N_985);
and U1082 (N_1082,N_1020,N_1024);
and U1083 (N_1083,N_1008,N_1012);
or U1084 (N_1084,N_1018,N_986);
nor U1085 (N_1085,N_999,N_1038);
nand U1086 (N_1086,N_1011,N_1001);
and U1087 (N_1087,N_1022,N_996);
or U1088 (N_1088,N_1031,N_984);
or U1089 (N_1089,N_1028,N_1005);
nand U1090 (N_1090,N_1022,N_987);
and U1091 (N_1091,N_1044,N_991);
or U1092 (N_1092,N_1020,N_1030);
nand U1093 (N_1093,N_987,N_994);
nand U1094 (N_1094,N_1036,N_1009);
or U1095 (N_1095,N_1016,N_977);
and U1096 (N_1096,N_1017,N_997);
nor U1097 (N_1097,N_1007,N_1042);
nor U1098 (N_1098,N_1023,N_1029);
or U1099 (N_1099,N_1031,N_996);
nand U1100 (N_1100,N_989,N_998);
or U1101 (N_1101,N_1007,N_1036);
or U1102 (N_1102,N_1037,N_1045);
nand U1103 (N_1103,N_1013,N_1036);
or U1104 (N_1104,N_1002,N_1012);
or U1105 (N_1105,N_978,N_1037);
and U1106 (N_1106,N_1020,N_1008);
nor U1107 (N_1107,N_1042,N_994);
nand U1108 (N_1108,N_1047,N_1030);
nand U1109 (N_1109,N_1011,N_1040);
or U1110 (N_1110,N_988,N_1025);
and U1111 (N_1111,N_1033,N_1043);
and U1112 (N_1112,N_1002,N_1014);
and U1113 (N_1113,N_1005,N_1036);
nor U1114 (N_1114,N_977,N_1029);
nand U1115 (N_1115,N_1040,N_988);
nor U1116 (N_1116,N_1000,N_1041);
nor U1117 (N_1117,N_986,N_978);
or U1118 (N_1118,N_1001,N_999);
or U1119 (N_1119,N_1007,N_1048);
nand U1120 (N_1120,N_980,N_1020);
and U1121 (N_1121,N_1046,N_1028);
nor U1122 (N_1122,N_1046,N_1031);
or U1123 (N_1123,N_1013,N_985);
nor U1124 (N_1124,N_1015,N_1000);
xor U1125 (N_1125,N_1058,N_1069);
or U1126 (N_1126,N_1111,N_1050);
nand U1127 (N_1127,N_1118,N_1068);
xor U1128 (N_1128,N_1053,N_1075);
or U1129 (N_1129,N_1101,N_1113);
and U1130 (N_1130,N_1107,N_1054);
or U1131 (N_1131,N_1108,N_1070);
and U1132 (N_1132,N_1088,N_1116);
or U1133 (N_1133,N_1055,N_1098);
xor U1134 (N_1134,N_1067,N_1074);
nor U1135 (N_1135,N_1120,N_1096);
and U1136 (N_1136,N_1106,N_1078);
nor U1137 (N_1137,N_1110,N_1086);
or U1138 (N_1138,N_1082,N_1051);
nand U1139 (N_1139,N_1089,N_1064);
nor U1140 (N_1140,N_1062,N_1079);
or U1141 (N_1141,N_1066,N_1052);
nand U1142 (N_1142,N_1117,N_1114);
and U1143 (N_1143,N_1112,N_1061);
nand U1144 (N_1144,N_1083,N_1071);
or U1145 (N_1145,N_1100,N_1059);
nor U1146 (N_1146,N_1072,N_1077);
or U1147 (N_1147,N_1097,N_1109);
and U1148 (N_1148,N_1081,N_1094);
nand U1149 (N_1149,N_1057,N_1099);
nor U1150 (N_1150,N_1102,N_1104);
nand U1151 (N_1151,N_1103,N_1122);
and U1152 (N_1152,N_1056,N_1065);
nor U1153 (N_1153,N_1124,N_1095);
and U1154 (N_1154,N_1063,N_1076);
or U1155 (N_1155,N_1092,N_1121);
and U1156 (N_1156,N_1093,N_1090);
nor U1157 (N_1157,N_1091,N_1087);
nor U1158 (N_1158,N_1119,N_1123);
or U1159 (N_1159,N_1085,N_1060);
or U1160 (N_1160,N_1115,N_1105);
and U1161 (N_1161,N_1080,N_1073);
xor U1162 (N_1162,N_1084,N_1072);
or U1163 (N_1163,N_1056,N_1074);
nand U1164 (N_1164,N_1109,N_1081);
or U1165 (N_1165,N_1067,N_1091);
xor U1166 (N_1166,N_1057,N_1072);
nor U1167 (N_1167,N_1107,N_1079);
nand U1168 (N_1168,N_1078,N_1053);
nor U1169 (N_1169,N_1085,N_1083);
and U1170 (N_1170,N_1057,N_1069);
nand U1171 (N_1171,N_1061,N_1096);
and U1172 (N_1172,N_1061,N_1110);
and U1173 (N_1173,N_1122,N_1108);
and U1174 (N_1174,N_1057,N_1098);
and U1175 (N_1175,N_1122,N_1074);
nand U1176 (N_1176,N_1066,N_1109);
and U1177 (N_1177,N_1076,N_1075);
or U1178 (N_1178,N_1091,N_1052);
or U1179 (N_1179,N_1077,N_1085);
or U1180 (N_1180,N_1112,N_1106);
or U1181 (N_1181,N_1064,N_1076);
and U1182 (N_1182,N_1123,N_1120);
or U1183 (N_1183,N_1092,N_1062);
and U1184 (N_1184,N_1096,N_1072);
and U1185 (N_1185,N_1076,N_1060);
and U1186 (N_1186,N_1105,N_1110);
nand U1187 (N_1187,N_1100,N_1098);
or U1188 (N_1188,N_1069,N_1061);
nor U1189 (N_1189,N_1115,N_1109);
nand U1190 (N_1190,N_1081,N_1098);
nor U1191 (N_1191,N_1087,N_1102);
nand U1192 (N_1192,N_1118,N_1073);
nor U1193 (N_1193,N_1092,N_1053);
nand U1194 (N_1194,N_1073,N_1089);
or U1195 (N_1195,N_1102,N_1078);
or U1196 (N_1196,N_1057,N_1090);
nand U1197 (N_1197,N_1077,N_1074);
or U1198 (N_1198,N_1076,N_1081);
or U1199 (N_1199,N_1101,N_1057);
or U1200 (N_1200,N_1152,N_1189);
nand U1201 (N_1201,N_1160,N_1135);
nand U1202 (N_1202,N_1126,N_1155);
nand U1203 (N_1203,N_1170,N_1185);
or U1204 (N_1204,N_1165,N_1176);
or U1205 (N_1205,N_1175,N_1182);
nor U1206 (N_1206,N_1125,N_1144);
or U1207 (N_1207,N_1180,N_1177);
and U1208 (N_1208,N_1197,N_1137);
or U1209 (N_1209,N_1184,N_1191);
and U1210 (N_1210,N_1190,N_1136);
and U1211 (N_1211,N_1141,N_1194);
or U1212 (N_1212,N_1129,N_1196);
nor U1213 (N_1213,N_1130,N_1173);
or U1214 (N_1214,N_1174,N_1146);
and U1215 (N_1215,N_1143,N_1198);
nor U1216 (N_1216,N_1172,N_1183);
and U1217 (N_1217,N_1134,N_1150);
nor U1218 (N_1218,N_1181,N_1133);
nor U1219 (N_1219,N_1142,N_1167);
xor U1220 (N_1220,N_1145,N_1193);
or U1221 (N_1221,N_1154,N_1161);
nand U1222 (N_1222,N_1179,N_1140);
and U1223 (N_1223,N_1139,N_1132);
or U1224 (N_1224,N_1149,N_1192);
nand U1225 (N_1225,N_1131,N_1166);
nand U1226 (N_1226,N_1187,N_1163);
nor U1227 (N_1227,N_1156,N_1128);
nand U1228 (N_1228,N_1169,N_1195);
nor U1229 (N_1229,N_1162,N_1199);
nand U1230 (N_1230,N_1147,N_1159);
or U1231 (N_1231,N_1127,N_1153);
nand U1232 (N_1232,N_1178,N_1157);
nand U1233 (N_1233,N_1164,N_1188);
or U1234 (N_1234,N_1171,N_1151);
and U1235 (N_1235,N_1186,N_1148);
or U1236 (N_1236,N_1158,N_1138);
nand U1237 (N_1237,N_1168,N_1140);
or U1238 (N_1238,N_1130,N_1183);
or U1239 (N_1239,N_1137,N_1190);
nor U1240 (N_1240,N_1178,N_1161);
and U1241 (N_1241,N_1167,N_1187);
or U1242 (N_1242,N_1132,N_1153);
or U1243 (N_1243,N_1129,N_1193);
or U1244 (N_1244,N_1152,N_1163);
nand U1245 (N_1245,N_1125,N_1174);
nand U1246 (N_1246,N_1145,N_1160);
and U1247 (N_1247,N_1179,N_1164);
and U1248 (N_1248,N_1166,N_1137);
or U1249 (N_1249,N_1128,N_1198);
and U1250 (N_1250,N_1133,N_1166);
and U1251 (N_1251,N_1195,N_1198);
nand U1252 (N_1252,N_1152,N_1136);
and U1253 (N_1253,N_1191,N_1140);
nand U1254 (N_1254,N_1148,N_1155);
nor U1255 (N_1255,N_1194,N_1186);
or U1256 (N_1256,N_1173,N_1140);
nor U1257 (N_1257,N_1143,N_1173);
nor U1258 (N_1258,N_1152,N_1150);
nor U1259 (N_1259,N_1166,N_1154);
and U1260 (N_1260,N_1197,N_1187);
or U1261 (N_1261,N_1154,N_1176);
and U1262 (N_1262,N_1175,N_1157);
nor U1263 (N_1263,N_1155,N_1128);
or U1264 (N_1264,N_1157,N_1125);
nor U1265 (N_1265,N_1149,N_1198);
nor U1266 (N_1266,N_1127,N_1150);
nand U1267 (N_1267,N_1131,N_1128);
or U1268 (N_1268,N_1193,N_1185);
nor U1269 (N_1269,N_1146,N_1173);
or U1270 (N_1270,N_1172,N_1154);
xor U1271 (N_1271,N_1191,N_1182);
nand U1272 (N_1272,N_1126,N_1140);
nor U1273 (N_1273,N_1168,N_1139);
xor U1274 (N_1274,N_1172,N_1180);
nand U1275 (N_1275,N_1270,N_1250);
and U1276 (N_1276,N_1209,N_1259);
and U1277 (N_1277,N_1205,N_1242);
xor U1278 (N_1278,N_1264,N_1220);
and U1279 (N_1279,N_1254,N_1239);
nor U1280 (N_1280,N_1271,N_1269);
nand U1281 (N_1281,N_1221,N_1206);
nor U1282 (N_1282,N_1256,N_1203);
or U1283 (N_1283,N_1268,N_1207);
nand U1284 (N_1284,N_1257,N_1249);
xor U1285 (N_1285,N_1202,N_1214);
and U1286 (N_1286,N_1274,N_1248);
and U1287 (N_1287,N_1216,N_1226);
nor U1288 (N_1288,N_1265,N_1210);
and U1289 (N_1289,N_1245,N_1223);
or U1290 (N_1290,N_1260,N_1222);
nor U1291 (N_1291,N_1244,N_1213);
nand U1292 (N_1292,N_1204,N_1258);
and U1293 (N_1293,N_1237,N_1243);
nor U1294 (N_1294,N_1263,N_1211);
or U1295 (N_1295,N_1232,N_1262);
or U1296 (N_1296,N_1251,N_1234);
xnor U1297 (N_1297,N_1238,N_1247);
nand U1298 (N_1298,N_1227,N_1233);
xnor U1299 (N_1299,N_1235,N_1267);
and U1300 (N_1300,N_1208,N_1225);
nor U1301 (N_1301,N_1229,N_1273);
nor U1302 (N_1302,N_1224,N_1218);
nor U1303 (N_1303,N_1253,N_1215);
nand U1304 (N_1304,N_1261,N_1246);
nand U1305 (N_1305,N_1230,N_1231);
nand U1306 (N_1306,N_1200,N_1228);
and U1307 (N_1307,N_1217,N_1212);
and U1308 (N_1308,N_1255,N_1266);
nor U1309 (N_1309,N_1219,N_1236);
or U1310 (N_1310,N_1240,N_1272);
xnor U1311 (N_1311,N_1252,N_1241);
or U1312 (N_1312,N_1201,N_1243);
or U1313 (N_1313,N_1211,N_1201);
nand U1314 (N_1314,N_1200,N_1220);
nor U1315 (N_1315,N_1243,N_1267);
and U1316 (N_1316,N_1238,N_1270);
and U1317 (N_1317,N_1274,N_1209);
nor U1318 (N_1318,N_1237,N_1254);
or U1319 (N_1319,N_1205,N_1212);
nand U1320 (N_1320,N_1271,N_1200);
xnor U1321 (N_1321,N_1257,N_1252);
or U1322 (N_1322,N_1260,N_1232);
or U1323 (N_1323,N_1261,N_1274);
nand U1324 (N_1324,N_1244,N_1270);
and U1325 (N_1325,N_1216,N_1258);
or U1326 (N_1326,N_1240,N_1262);
nor U1327 (N_1327,N_1247,N_1226);
or U1328 (N_1328,N_1237,N_1266);
nor U1329 (N_1329,N_1268,N_1239);
nand U1330 (N_1330,N_1202,N_1259);
or U1331 (N_1331,N_1273,N_1266);
and U1332 (N_1332,N_1224,N_1242);
and U1333 (N_1333,N_1217,N_1239);
and U1334 (N_1334,N_1231,N_1272);
xor U1335 (N_1335,N_1248,N_1211);
nand U1336 (N_1336,N_1219,N_1238);
and U1337 (N_1337,N_1263,N_1252);
nand U1338 (N_1338,N_1205,N_1215);
and U1339 (N_1339,N_1222,N_1204);
or U1340 (N_1340,N_1272,N_1234);
nor U1341 (N_1341,N_1202,N_1273);
nand U1342 (N_1342,N_1236,N_1213);
xor U1343 (N_1343,N_1245,N_1227);
nor U1344 (N_1344,N_1222,N_1256);
nand U1345 (N_1345,N_1237,N_1214);
nor U1346 (N_1346,N_1209,N_1220);
or U1347 (N_1347,N_1271,N_1252);
or U1348 (N_1348,N_1263,N_1229);
nand U1349 (N_1349,N_1252,N_1240);
xnor U1350 (N_1350,N_1313,N_1314);
nor U1351 (N_1351,N_1286,N_1322);
nand U1352 (N_1352,N_1289,N_1285);
nand U1353 (N_1353,N_1334,N_1336);
and U1354 (N_1354,N_1343,N_1279);
nand U1355 (N_1355,N_1333,N_1315);
nand U1356 (N_1356,N_1307,N_1301);
or U1357 (N_1357,N_1281,N_1312);
and U1358 (N_1358,N_1288,N_1319);
xor U1359 (N_1359,N_1349,N_1316);
nand U1360 (N_1360,N_1346,N_1293);
nor U1361 (N_1361,N_1325,N_1341);
nand U1362 (N_1362,N_1277,N_1284);
nor U1363 (N_1363,N_1332,N_1308);
or U1364 (N_1364,N_1309,N_1297);
nand U1365 (N_1365,N_1331,N_1311);
nor U1366 (N_1366,N_1337,N_1276);
nand U1367 (N_1367,N_1299,N_1295);
nand U1368 (N_1368,N_1282,N_1304);
or U1369 (N_1369,N_1310,N_1329);
nand U1370 (N_1370,N_1320,N_1348);
or U1371 (N_1371,N_1338,N_1302);
and U1372 (N_1372,N_1275,N_1347);
nand U1373 (N_1373,N_1330,N_1292);
or U1374 (N_1374,N_1298,N_1340);
and U1375 (N_1375,N_1306,N_1287);
and U1376 (N_1376,N_1324,N_1328);
nor U1377 (N_1377,N_1291,N_1342);
nor U1378 (N_1378,N_1345,N_1344);
nand U1379 (N_1379,N_1326,N_1323);
or U1380 (N_1380,N_1321,N_1303);
or U1381 (N_1381,N_1335,N_1283);
nand U1382 (N_1382,N_1305,N_1318);
and U1383 (N_1383,N_1317,N_1296);
xnor U1384 (N_1384,N_1290,N_1280);
xor U1385 (N_1385,N_1294,N_1278);
or U1386 (N_1386,N_1327,N_1339);
or U1387 (N_1387,N_1300,N_1308);
nor U1388 (N_1388,N_1343,N_1281);
nand U1389 (N_1389,N_1317,N_1284);
nand U1390 (N_1390,N_1275,N_1289);
or U1391 (N_1391,N_1310,N_1285);
or U1392 (N_1392,N_1291,N_1325);
nand U1393 (N_1393,N_1325,N_1283);
or U1394 (N_1394,N_1283,N_1320);
or U1395 (N_1395,N_1280,N_1291);
nor U1396 (N_1396,N_1320,N_1346);
and U1397 (N_1397,N_1331,N_1293);
nand U1398 (N_1398,N_1312,N_1341);
and U1399 (N_1399,N_1302,N_1311);
nor U1400 (N_1400,N_1345,N_1297);
nand U1401 (N_1401,N_1305,N_1340);
and U1402 (N_1402,N_1295,N_1298);
nor U1403 (N_1403,N_1329,N_1282);
and U1404 (N_1404,N_1288,N_1292);
and U1405 (N_1405,N_1324,N_1308);
or U1406 (N_1406,N_1285,N_1308);
nand U1407 (N_1407,N_1326,N_1290);
and U1408 (N_1408,N_1304,N_1347);
and U1409 (N_1409,N_1285,N_1278);
nor U1410 (N_1410,N_1305,N_1341);
nor U1411 (N_1411,N_1283,N_1277);
nand U1412 (N_1412,N_1293,N_1316);
and U1413 (N_1413,N_1316,N_1319);
or U1414 (N_1414,N_1345,N_1314);
or U1415 (N_1415,N_1290,N_1314);
or U1416 (N_1416,N_1290,N_1324);
nor U1417 (N_1417,N_1291,N_1284);
and U1418 (N_1418,N_1341,N_1330);
nand U1419 (N_1419,N_1298,N_1344);
nor U1420 (N_1420,N_1280,N_1293);
nor U1421 (N_1421,N_1321,N_1301);
or U1422 (N_1422,N_1328,N_1290);
or U1423 (N_1423,N_1349,N_1346);
or U1424 (N_1424,N_1321,N_1320);
nor U1425 (N_1425,N_1417,N_1397);
nand U1426 (N_1426,N_1388,N_1405);
xnor U1427 (N_1427,N_1366,N_1363);
nand U1428 (N_1428,N_1364,N_1353);
and U1429 (N_1429,N_1402,N_1406);
or U1430 (N_1430,N_1400,N_1386);
nor U1431 (N_1431,N_1384,N_1371);
or U1432 (N_1432,N_1394,N_1380);
nand U1433 (N_1433,N_1350,N_1395);
nand U1434 (N_1434,N_1379,N_1418);
nor U1435 (N_1435,N_1393,N_1407);
and U1436 (N_1436,N_1381,N_1374);
and U1437 (N_1437,N_1370,N_1387);
nand U1438 (N_1438,N_1421,N_1369);
nor U1439 (N_1439,N_1413,N_1360);
and U1440 (N_1440,N_1420,N_1412);
nor U1441 (N_1441,N_1396,N_1373);
and U1442 (N_1442,N_1382,N_1355);
or U1443 (N_1443,N_1389,N_1376);
xnor U1444 (N_1444,N_1378,N_1367);
nor U1445 (N_1445,N_1351,N_1383);
and U1446 (N_1446,N_1385,N_1424);
nand U1447 (N_1447,N_1377,N_1375);
nor U1448 (N_1448,N_1399,N_1423);
nor U1449 (N_1449,N_1398,N_1414);
nor U1450 (N_1450,N_1352,N_1368);
or U1451 (N_1451,N_1410,N_1403);
nand U1452 (N_1452,N_1415,N_1401);
and U1453 (N_1453,N_1416,N_1411);
or U1454 (N_1454,N_1404,N_1358);
or U1455 (N_1455,N_1359,N_1365);
xnor U1456 (N_1456,N_1408,N_1390);
xnor U1457 (N_1457,N_1362,N_1354);
nor U1458 (N_1458,N_1357,N_1391);
and U1459 (N_1459,N_1419,N_1422);
nor U1460 (N_1460,N_1372,N_1409);
and U1461 (N_1461,N_1392,N_1356);
nand U1462 (N_1462,N_1361,N_1389);
xor U1463 (N_1463,N_1395,N_1400);
nor U1464 (N_1464,N_1376,N_1370);
nor U1465 (N_1465,N_1423,N_1404);
or U1466 (N_1466,N_1367,N_1376);
or U1467 (N_1467,N_1414,N_1391);
or U1468 (N_1468,N_1353,N_1384);
and U1469 (N_1469,N_1358,N_1395);
or U1470 (N_1470,N_1418,N_1366);
nor U1471 (N_1471,N_1379,N_1352);
or U1472 (N_1472,N_1401,N_1374);
nand U1473 (N_1473,N_1407,N_1396);
and U1474 (N_1474,N_1363,N_1365);
or U1475 (N_1475,N_1405,N_1404);
nand U1476 (N_1476,N_1365,N_1373);
or U1477 (N_1477,N_1362,N_1424);
or U1478 (N_1478,N_1423,N_1386);
and U1479 (N_1479,N_1424,N_1395);
xor U1480 (N_1480,N_1396,N_1368);
nand U1481 (N_1481,N_1383,N_1421);
and U1482 (N_1482,N_1411,N_1368);
nand U1483 (N_1483,N_1355,N_1423);
nand U1484 (N_1484,N_1366,N_1415);
xnor U1485 (N_1485,N_1359,N_1399);
nor U1486 (N_1486,N_1393,N_1411);
or U1487 (N_1487,N_1358,N_1369);
or U1488 (N_1488,N_1387,N_1409);
and U1489 (N_1489,N_1354,N_1373);
or U1490 (N_1490,N_1380,N_1362);
nand U1491 (N_1491,N_1389,N_1380);
and U1492 (N_1492,N_1411,N_1390);
nand U1493 (N_1493,N_1388,N_1377);
nor U1494 (N_1494,N_1390,N_1361);
nor U1495 (N_1495,N_1377,N_1386);
xor U1496 (N_1496,N_1394,N_1369);
nand U1497 (N_1497,N_1404,N_1407);
and U1498 (N_1498,N_1384,N_1376);
or U1499 (N_1499,N_1361,N_1355);
xor U1500 (N_1500,N_1462,N_1498);
nor U1501 (N_1501,N_1430,N_1446);
nand U1502 (N_1502,N_1463,N_1436);
xnor U1503 (N_1503,N_1433,N_1434);
or U1504 (N_1504,N_1470,N_1454);
and U1505 (N_1505,N_1431,N_1465);
nand U1506 (N_1506,N_1448,N_1490);
and U1507 (N_1507,N_1492,N_1440);
nor U1508 (N_1508,N_1495,N_1437);
and U1509 (N_1509,N_1429,N_1496);
or U1510 (N_1510,N_1473,N_1450);
or U1511 (N_1511,N_1485,N_1499);
nor U1512 (N_1512,N_1460,N_1425);
and U1513 (N_1513,N_1488,N_1481);
and U1514 (N_1514,N_1482,N_1476);
nor U1515 (N_1515,N_1456,N_1467);
nor U1516 (N_1516,N_1469,N_1468);
nand U1517 (N_1517,N_1455,N_1444);
or U1518 (N_1518,N_1491,N_1487);
and U1519 (N_1519,N_1494,N_1438);
nor U1520 (N_1520,N_1432,N_1466);
xor U1521 (N_1521,N_1474,N_1477);
and U1522 (N_1522,N_1483,N_1461);
or U1523 (N_1523,N_1484,N_1497);
or U1524 (N_1524,N_1458,N_1445);
and U1525 (N_1525,N_1443,N_1464);
nor U1526 (N_1526,N_1435,N_1457);
and U1527 (N_1527,N_1478,N_1493);
nor U1528 (N_1528,N_1459,N_1439);
and U1529 (N_1529,N_1471,N_1475);
and U1530 (N_1530,N_1441,N_1451);
and U1531 (N_1531,N_1489,N_1428);
or U1532 (N_1532,N_1447,N_1472);
or U1533 (N_1533,N_1486,N_1427);
nand U1534 (N_1534,N_1479,N_1442);
or U1535 (N_1535,N_1426,N_1453);
or U1536 (N_1536,N_1452,N_1449);
xor U1537 (N_1537,N_1480,N_1452);
nand U1538 (N_1538,N_1462,N_1474);
or U1539 (N_1539,N_1446,N_1464);
nor U1540 (N_1540,N_1437,N_1454);
nor U1541 (N_1541,N_1426,N_1466);
nand U1542 (N_1542,N_1497,N_1461);
xor U1543 (N_1543,N_1475,N_1447);
nand U1544 (N_1544,N_1429,N_1462);
or U1545 (N_1545,N_1450,N_1429);
nand U1546 (N_1546,N_1468,N_1437);
xor U1547 (N_1547,N_1479,N_1443);
nand U1548 (N_1548,N_1437,N_1489);
or U1549 (N_1549,N_1453,N_1439);
or U1550 (N_1550,N_1431,N_1478);
nand U1551 (N_1551,N_1456,N_1460);
or U1552 (N_1552,N_1462,N_1493);
or U1553 (N_1553,N_1465,N_1443);
xor U1554 (N_1554,N_1467,N_1479);
xor U1555 (N_1555,N_1444,N_1482);
xnor U1556 (N_1556,N_1493,N_1443);
nand U1557 (N_1557,N_1447,N_1431);
nor U1558 (N_1558,N_1458,N_1461);
and U1559 (N_1559,N_1488,N_1436);
nand U1560 (N_1560,N_1442,N_1434);
xor U1561 (N_1561,N_1469,N_1496);
xnor U1562 (N_1562,N_1466,N_1463);
or U1563 (N_1563,N_1483,N_1439);
xnor U1564 (N_1564,N_1451,N_1452);
or U1565 (N_1565,N_1455,N_1477);
nand U1566 (N_1566,N_1481,N_1466);
nand U1567 (N_1567,N_1468,N_1434);
or U1568 (N_1568,N_1468,N_1439);
xor U1569 (N_1569,N_1431,N_1425);
nand U1570 (N_1570,N_1430,N_1439);
or U1571 (N_1571,N_1453,N_1499);
and U1572 (N_1572,N_1487,N_1484);
nand U1573 (N_1573,N_1470,N_1441);
nor U1574 (N_1574,N_1441,N_1472);
or U1575 (N_1575,N_1544,N_1523);
and U1576 (N_1576,N_1534,N_1509);
xor U1577 (N_1577,N_1565,N_1527);
nand U1578 (N_1578,N_1570,N_1554);
nor U1579 (N_1579,N_1531,N_1539);
xor U1580 (N_1580,N_1528,N_1543);
or U1581 (N_1581,N_1571,N_1541);
or U1582 (N_1582,N_1550,N_1553);
and U1583 (N_1583,N_1559,N_1566);
or U1584 (N_1584,N_1503,N_1535);
or U1585 (N_1585,N_1524,N_1540);
xor U1586 (N_1586,N_1525,N_1574);
and U1587 (N_1587,N_1506,N_1551);
nand U1588 (N_1588,N_1573,N_1552);
and U1589 (N_1589,N_1518,N_1569);
nand U1590 (N_1590,N_1561,N_1516);
or U1591 (N_1591,N_1515,N_1556);
nor U1592 (N_1592,N_1549,N_1558);
and U1593 (N_1593,N_1568,N_1508);
nor U1594 (N_1594,N_1504,N_1507);
or U1595 (N_1595,N_1547,N_1562);
xnor U1596 (N_1596,N_1537,N_1520);
and U1597 (N_1597,N_1567,N_1545);
or U1598 (N_1598,N_1529,N_1542);
xor U1599 (N_1599,N_1526,N_1538);
nand U1600 (N_1600,N_1564,N_1500);
nor U1601 (N_1601,N_1519,N_1512);
or U1602 (N_1602,N_1560,N_1548);
or U1603 (N_1603,N_1514,N_1517);
nand U1604 (N_1604,N_1513,N_1546);
or U1605 (N_1605,N_1555,N_1563);
nand U1606 (N_1606,N_1557,N_1501);
nor U1607 (N_1607,N_1536,N_1533);
nand U1608 (N_1608,N_1522,N_1510);
and U1609 (N_1609,N_1530,N_1521);
or U1610 (N_1610,N_1532,N_1505);
nor U1611 (N_1611,N_1502,N_1511);
and U1612 (N_1612,N_1572,N_1515);
nor U1613 (N_1613,N_1505,N_1542);
nand U1614 (N_1614,N_1540,N_1545);
nor U1615 (N_1615,N_1564,N_1557);
nor U1616 (N_1616,N_1551,N_1543);
nand U1617 (N_1617,N_1558,N_1571);
nor U1618 (N_1618,N_1553,N_1502);
nor U1619 (N_1619,N_1513,N_1562);
and U1620 (N_1620,N_1521,N_1528);
or U1621 (N_1621,N_1551,N_1552);
nor U1622 (N_1622,N_1543,N_1546);
and U1623 (N_1623,N_1527,N_1560);
nor U1624 (N_1624,N_1538,N_1547);
nor U1625 (N_1625,N_1534,N_1536);
nor U1626 (N_1626,N_1514,N_1519);
nand U1627 (N_1627,N_1543,N_1561);
nor U1628 (N_1628,N_1559,N_1523);
or U1629 (N_1629,N_1524,N_1531);
nor U1630 (N_1630,N_1512,N_1571);
or U1631 (N_1631,N_1509,N_1513);
nand U1632 (N_1632,N_1522,N_1534);
nand U1633 (N_1633,N_1555,N_1560);
or U1634 (N_1634,N_1550,N_1513);
and U1635 (N_1635,N_1535,N_1527);
and U1636 (N_1636,N_1508,N_1547);
nor U1637 (N_1637,N_1559,N_1521);
or U1638 (N_1638,N_1546,N_1566);
and U1639 (N_1639,N_1548,N_1519);
and U1640 (N_1640,N_1520,N_1553);
nor U1641 (N_1641,N_1547,N_1511);
or U1642 (N_1642,N_1511,N_1560);
or U1643 (N_1643,N_1527,N_1518);
or U1644 (N_1644,N_1539,N_1552);
nor U1645 (N_1645,N_1564,N_1574);
nor U1646 (N_1646,N_1563,N_1561);
nand U1647 (N_1647,N_1544,N_1564);
and U1648 (N_1648,N_1508,N_1558);
or U1649 (N_1649,N_1524,N_1519);
nand U1650 (N_1650,N_1597,N_1645);
xor U1651 (N_1651,N_1646,N_1642);
or U1652 (N_1652,N_1605,N_1616);
and U1653 (N_1653,N_1586,N_1599);
or U1654 (N_1654,N_1619,N_1610);
nor U1655 (N_1655,N_1603,N_1636);
or U1656 (N_1656,N_1631,N_1643);
or U1657 (N_1657,N_1622,N_1578);
nor U1658 (N_1658,N_1588,N_1601);
or U1659 (N_1659,N_1608,N_1648);
nor U1660 (N_1660,N_1580,N_1579);
nand U1661 (N_1661,N_1598,N_1625);
and U1662 (N_1662,N_1595,N_1623);
or U1663 (N_1663,N_1600,N_1607);
nand U1664 (N_1664,N_1615,N_1593);
nor U1665 (N_1665,N_1592,N_1594);
and U1666 (N_1666,N_1637,N_1596);
nor U1667 (N_1667,N_1647,N_1635);
or U1668 (N_1668,N_1618,N_1626);
or U1669 (N_1669,N_1617,N_1639);
and U1670 (N_1670,N_1577,N_1576);
nand U1671 (N_1671,N_1585,N_1575);
or U1672 (N_1672,N_1602,N_1624);
nand U1673 (N_1673,N_1629,N_1584);
nor U1674 (N_1674,N_1633,N_1620);
nand U1675 (N_1675,N_1638,N_1611);
nor U1676 (N_1676,N_1614,N_1613);
nand U1677 (N_1677,N_1628,N_1589);
or U1678 (N_1678,N_1581,N_1606);
and U1679 (N_1679,N_1630,N_1649);
nor U1680 (N_1680,N_1609,N_1583);
or U1681 (N_1681,N_1632,N_1590);
or U1682 (N_1682,N_1627,N_1621);
nand U1683 (N_1683,N_1587,N_1644);
nor U1684 (N_1684,N_1641,N_1640);
nand U1685 (N_1685,N_1591,N_1604);
xor U1686 (N_1686,N_1582,N_1612);
nand U1687 (N_1687,N_1634,N_1638);
nor U1688 (N_1688,N_1637,N_1618);
nand U1689 (N_1689,N_1577,N_1595);
or U1690 (N_1690,N_1604,N_1648);
nor U1691 (N_1691,N_1579,N_1593);
or U1692 (N_1692,N_1600,N_1594);
or U1693 (N_1693,N_1646,N_1595);
and U1694 (N_1694,N_1575,N_1623);
and U1695 (N_1695,N_1641,N_1601);
nand U1696 (N_1696,N_1581,N_1630);
or U1697 (N_1697,N_1582,N_1593);
and U1698 (N_1698,N_1608,N_1646);
or U1699 (N_1699,N_1587,N_1624);
nor U1700 (N_1700,N_1611,N_1630);
and U1701 (N_1701,N_1582,N_1644);
nor U1702 (N_1702,N_1579,N_1623);
and U1703 (N_1703,N_1610,N_1602);
nand U1704 (N_1704,N_1613,N_1609);
nor U1705 (N_1705,N_1615,N_1592);
nor U1706 (N_1706,N_1636,N_1625);
nor U1707 (N_1707,N_1646,N_1636);
nand U1708 (N_1708,N_1614,N_1635);
nand U1709 (N_1709,N_1647,N_1634);
or U1710 (N_1710,N_1602,N_1648);
nand U1711 (N_1711,N_1575,N_1646);
nand U1712 (N_1712,N_1640,N_1596);
nor U1713 (N_1713,N_1627,N_1601);
nor U1714 (N_1714,N_1610,N_1595);
xnor U1715 (N_1715,N_1619,N_1593);
nor U1716 (N_1716,N_1615,N_1646);
and U1717 (N_1717,N_1598,N_1637);
nand U1718 (N_1718,N_1610,N_1622);
and U1719 (N_1719,N_1627,N_1585);
and U1720 (N_1720,N_1620,N_1637);
xnor U1721 (N_1721,N_1576,N_1609);
nor U1722 (N_1722,N_1593,N_1626);
nand U1723 (N_1723,N_1637,N_1589);
and U1724 (N_1724,N_1599,N_1581);
and U1725 (N_1725,N_1654,N_1684);
and U1726 (N_1726,N_1719,N_1658);
xor U1727 (N_1727,N_1697,N_1701);
nand U1728 (N_1728,N_1716,N_1718);
or U1729 (N_1729,N_1706,N_1665);
and U1730 (N_1730,N_1689,N_1660);
or U1731 (N_1731,N_1651,N_1683);
and U1732 (N_1732,N_1700,N_1674);
nor U1733 (N_1733,N_1722,N_1707);
nand U1734 (N_1734,N_1709,N_1657);
or U1735 (N_1735,N_1667,N_1685);
nor U1736 (N_1736,N_1680,N_1677);
or U1737 (N_1737,N_1678,N_1672);
and U1738 (N_1738,N_1666,N_1659);
or U1739 (N_1739,N_1686,N_1662);
nand U1740 (N_1740,N_1713,N_1708);
or U1741 (N_1741,N_1679,N_1675);
nor U1742 (N_1742,N_1668,N_1670);
and U1743 (N_1743,N_1705,N_1724);
nor U1744 (N_1744,N_1698,N_1704);
or U1745 (N_1745,N_1695,N_1687);
xor U1746 (N_1746,N_1692,N_1693);
nor U1747 (N_1747,N_1712,N_1681);
nor U1748 (N_1748,N_1676,N_1669);
nand U1749 (N_1749,N_1653,N_1652);
nand U1750 (N_1750,N_1661,N_1720);
nor U1751 (N_1751,N_1694,N_1721);
nand U1752 (N_1752,N_1715,N_1656);
nor U1753 (N_1753,N_1688,N_1702);
nor U1754 (N_1754,N_1671,N_1714);
nand U1755 (N_1755,N_1723,N_1699);
and U1756 (N_1756,N_1717,N_1663);
and U1757 (N_1757,N_1655,N_1664);
xnor U1758 (N_1758,N_1650,N_1710);
nor U1759 (N_1759,N_1696,N_1673);
xnor U1760 (N_1760,N_1711,N_1703);
or U1761 (N_1761,N_1690,N_1682);
or U1762 (N_1762,N_1691,N_1698);
or U1763 (N_1763,N_1663,N_1723);
nand U1764 (N_1764,N_1682,N_1715);
or U1765 (N_1765,N_1687,N_1713);
nor U1766 (N_1766,N_1672,N_1651);
and U1767 (N_1767,N_1712,N_1652);
or U1768 (N_1768,N_1675,N_1706);
or U1769 (N_1769,N_1682,N_1704);
nand U1770 (N_1770,N_1683,N_1691);
nand U1771 (N_1771,N_1710,N_1694);
nand U1772 (N_1772,N_1677,N_1712);
nor U1773 (N_1773,N_1722,N_1671);
or U1774 (N_1774,N_1723,N_1697);
nand U1775 (N_1775,N_1653,N_1659);
nor U1776 (N_1776,N_1656,N_1706);
and U1777 (N_1777,N_1708,N_1677);
nor U1778 (N_1778,N_1685,N_1722);
xor U1779 (N_1779,N_1656,N_1720);
nand U1780 (N_1780,N_1662,N_1710);
nand U1781 (N_1781,N_1721,N_1715);
nand U1782 (N_1782,N_1707,N_1702);
and U1783 (N_1783,N_1698,N_1720);
and U1784 (N_1784,N_1676,N_1715);
nor U1785 (N_1785,N_1721,N_1700);
nor U1786 (N_1786,N_1650,N_1677);
or U1787 (N_1787,N_1715,N_1691);
nand U1788 (N_1788,N_1675,N_1715);
or U1789 (N_1789,N_1713,N_1702);
or U1790 (N_1790,N_1696,N_1675);
and U1791 (N_1791,N_1658,N_1690);
nand U1792 (N_1792,N_1716,N_1686);
and U1793 (N_1793,N_1673,N_1693);
or U1794 (N_1794,N_1682,N_1670);
nor U1795 (N_1795,N_1669,N_1679);
or U1796 (N_1796,N_1721,N_1670);
or U1797 (N_1797,N_1655,N_1689);
xor U1798 (N_1798,N_1701,N_1679);
or U1799 (N_1799,N_1664,N_1663);
nand U1800 (N_1800,N_1788,N_1727);
and U1801 (N_1801,N_1782,N_1795);
nor U1802 (N_1802,N_1761,N_1740);
xnor U1803 (N_1803,N_1763,N_1726);
or U1804 (N_1804,N_1789,N_1765);
nor U1805 (N_1805,N_1786,N_1751);
nand U1806 (N_1806,N_1749,N_1769);
and U1807 (N_1807,N_1734,N_1758);
or U1808 (N_1808,N_1757,N_1794);
or U1809 (N_1809,N_1752,N_1750);
or U1810 (N_1810,N_1775,N_1730);
and U1811 (N_1811,N_1762,N_1729);
nor U1812 (N_1812,N_1728,N_1777);
nor U1813 (N_1813,N_1731,N_1747);
or U1814 (N_1814,N_1739,N_1736);
nand U1815 (N_1815,N_1759,N_1796);
nor U1816 (N_1816,N_1780,N_1793);
and U1817 (N_1817,N_1776,N_1781);
nand U1818 (N_1818,N_1746,N_1741);
nor U1819 (N_1819,N_1766,N_1772);
and U1820 (N_1820,N_1735,N_1767);
nand U1821 (N_1821,N_1732,N_1764);
and U1822 (N_1822,N_1787,N_1778);
and U1823 (N_1823,N_1733,N_1797);
nor U1824 (N_1824,N_1798,N_1784);
or U1825 (N_1825,N_1770,N_1753);
or U1826 (N_1826,N_1744,N_1790);
nand U1827 (N_1827,N_1791,N_1738);
and U1828 (N_1828,N_1768,N_1743);
xor U1829 (N_1829,N_1760,N_1799);
nand U1830 (N_1830,N_1783,N_1756);
xor U1831 (N_1831,N_1725,N_1771);
or U1832 (N_1832,N_1754,N_1785);
nand U1833 (N_1833,N_1748,N_1779);
nand U1834 (N_1834,N_1774,N_1773);
or U1835 (N_1835,N_1737,N_1755);
and U1836 (N_1836,N_1742,N_1745);
and U1837 (N_1837,N_1792,N_1796);
xor U1838 (N_1838,N_1741,N_1735);
nor U1839 (N_1839,N_1780,N_1778);
and U1840 (N_1840,N_1752,N_1785);
and U1841 (N_1841,N_1743,N_1785);
nor U1842 (N_1842,N_1759,N_1778);
nor U1843 (N_1843,N_1798,N_1777);
nand U1844 (N_1844,N_1764,N_1796);
or U1845 (N_1845,N_1796,N_1745);
and U1846 (N_1846,N_1783,N_1766);
or U1847 (N_1847,N_1739,N_1738);
or U1848 (N_1848,N_1779,N_1790);
and U1849 (N_1849,N_1799,N_1749);
xor U1850 (N_1850,N_1747,N_1765);
nand U1851 (N_1851,N_1748,N_1737);
xor U1852 (N_1852,N_1754,N_1780);
or U1853 (N_1853,N_1792,N_1742);
nor U1854 (N_1854,N_1753,N_1734);
xor U1855 (N_1855,N_1792,N_1788);
nor U1856 (N_1856,N_1727,N_1795);
or U1857 (N_1857,N_1779,N_1752);
nand U1858 (N_1858,N_1759,N_1762);
nor U1859 (N_1859,N_1739,N_1741);
nor U1860 (N_1860,N_1742,N_1758);
nor U1861 (N_1861,N_1765,N_1748);
nand U1862 (N_1862,N_1748,N_1726);
nand U1863 (N_1863,N_1748,N_1768);
or U1864 (N_1864,N_1757,N_1792);
and U1865 (N_1865,N_1776,N_1744);
nand U1866 (N_1866,N_1743,N_1794);
nand U1867 (N_1867,N_1789,N_1798);
nand U1868 (N_1868,N_1798,N_1795);
or U1869 (N_1869,N_1781,N_1763);
and U1870 (N_1870,N_1782,N_1749);
nand U1871 (N_1871,N_1781,N_1777);
nor U1872 (N_1872,N_1786,N_1767);
and U1873 (N_1873,N_1792,N_1762);
and U1874 (N_1874,N_1737,N_1746);
nor U1875 (N_1875,N_1827,N_1860);
or U1876 (N_1876,N_1864,N_1857);
or U1877 (N_1877,N_1806,N_1833);
nand U1878 (N_1878,N_1844,N_1854);
nand U1879 (N_1879,N_1811,N_1822);
nand U1880 (N_1880,N_1850,N_1843);
or U1881 (N_1881,N_1814,N_1817);
and U1882 (N_1882,N_1839,N_1826);
nor U1883 (N_1883,N_1871,N_1859);
nor U1884 (N_1884,N_1807,N_1815);
and U1885 (N_1885,N_1856,N_1862);
nor U1886 (N_1886,N_1851,N_1830);
or U1887 (N_1887,N_1816,N_1813);
and U1888 (N_1888,N_1825,N_1848);
nand U1889 (N_1889,N_1829,N_1828);
nor U1890 (N_1890,N_1819,N_1804);
and U1891 (N_1891,N_1870,N_1820);
and U1892 (N_1892,N_1874,N_1861);
nor U1893 (N_1893,N_1868,N_1855);
nand U1894 (N_1894,N_1802,N_1818);
or U1895 (N_1895,N_1803,N_1863);
nand U1896 (N_1896,N_1849,N_1869);
xnor U1897 (N_1897,N_1837,N_1810);
and U1898 (N_1898,N_1834,N_1867);
and U1899 (N_1899,N_1835,N_1841);
or U1900 (N_1900,N_1872,N_1836);
nand U1901 (N_1901,N_1838,N_1865);
and U1902 (N_1902,N_1812,N_1831);
xnor U1903 (N_1903,N_1823,N_1808);
or U1904 (N_1904,N_1821,N_1824);
nor U1905 (N_1905,N_1805,N_1840);
and U1906 (N_1906,N_1801,N_1800);
nand U1907 (N_1907,N_1832,N_1853);
nor U1908 (N_1908,N_1873,N_1866);
or U1909 (N_1909,N_1845,N_1852);
nand U1910 (N_1910,N_1809,N_1846);
nand U1911 (N_1911,N_1858,N_1847);
or U1912 (N_1912,N_1842,N_1807);
and U1913 (N_1913,N_1837,N_1841);
and U1914 (N_1914,N_1809,N_1811);
or U1915 (N_1915,N_1859,N_1824);
or U1916 (N_1916,N_1868,N_1813);
nor U1917 (N_1917,N_1805,N_1826);
and U1918 (N_1918,N_1865,N_1839);
or U1919 (N_1919,N_1828,N_1865);
xor U1920 (N_1920,N_1873,N_1832);
or U1921 (N_1921,N_1801,N_1811);
nor U1922 (N_1922,N_1802,N_1850);
nand U1923 (N_1923,N_1872,N_1859);
or U1924 (N_1924,N_1841,N_1854);
or U1925 (N_1925,N_1829,N_1806);
and U1926 (N_1926,N_1840,N_1806);
and U1927 (N_1927,N_1800,N_1853);
or U1928 (N_1928,N_1810,N_1848);
nor U1929 (N_1929,N_1821,N_1855);
nand U1930 (N_1930,N_1859,N_1804);
and U1931 (N_1931,N_1856,N_1803);
nand U1932 (N_1932,N_1831,N_1800);
nor U1933 (N_1933,N_1874,N_1842);
and U1934 (N_1934,N_1809,N_1860);
or U1935 (N_1935,N_1810,N_1867);
nor U1936 (N_1936,N_1818,N_1858);
nand U1937 (N_1937,N_1852,N_1817);
nor U1938 (N_1938,N_1816,N_1830);
or U1939 (N_1939,N_1836,N_1848);
xnor U1940 (N_1940,N_1830,N_1809);
xor U1941 (N_1941,N_1864,N_1868);
nor U1942 (N_1942,N_1808,N_1826);
or U1943 (N_1943,N_1828,N_1839);
or U1944 (N_1944,N_1828,N_1802);
and U1945 (N_1945,N_1857,N_1809);
and U1946 (N_1946,N_1866,N_1806);
nor U1947 (N_1947,N_1805,N_1806);
nand U1948 (N_1948,N_1833,N_1819);
and U1949 (N_1949,N_1836,N_1831);
nand U1950 (N_1950,N_1934,N_1914);
nor U1951 (N_1951,N_1939,N_1876);
and U1952 (N_1952,N_1938,N_1885);
nor U1953 (N_1953,N_1923,N_1903);
or U1954 (N_1954,N_1907,N_1904);
nor U1955 (N_1955,N_1887,N_1883);
xnor U1956 (N_1956,N_1913,N_1881);
nor U1957 (N_1957,N_1944,N_1932);
nor U1958 (N_1958,N_1926,N_1930);
nor U1959 (N_1959,N_1902,N_1924);
and U1960 (N_1960,N_1919,N_1921);
and U1961 (N_1961,N_1943,N_1909);
and U1962 (N_1962,N_1884,N_1893);
nand U1963 (N_1963,N_1895,N_1889);
or U1964 (N_1964,N_1935,N_1918);
or U1965 (N_1965,N_1928,N_1947);
nor U1966 (N_1966,N_1949,N_1901);
xor U1967 (N_1967,N_1898,N_1896);
or U1968 (N_1968,N_1882,N_1891);
nand U1969 (N_1969,N_1886,N_1875);
or U1970 (N_1970,N_1897,N_1877);
nand U1971 (N_1971,N_1933,N_1888);
nand U1972 (N_1972,N_1892,N_1936);
and U1973 (N_1973,N_1879,N_1948);
nand U1974 (N_1974,N_1912,N_1906);
nor U1975 (N_1975,N_1908,N_1946);
and U1976 (N_1976,N_1905,N_1899);
or U1977 (N_1977,N_1929,N_1910);
or U1978 (N_1978,N_1942,N_1880);
nor U1979 (N_1979,N_1890,N_1931);
xnor U1980 (N_1980,N_1894,N_1937);
nor U1981 (N_1981,N_1900,N_1925);
or U1982 (N_1982,N_1917,N_1920);
nand U1983 (N_1983,N_1945,N_1915);
or U1984 (N_1984,N_1878,N_1940);
nor U1985 (N_1985,N_1916,N_1922);
nand U1986 (N_1986,N_1927,N_1911);
nand U1987 (N_1987,N_1941,N_1925);
xnor U1988 (N_1988,N_1883,N_1916);
nor U1989 (N_1989,N_1885,N_1894);
or U1990 (N_1990,N_1901,N_1948);
and U1991 (N_1991,N_1907,N_1920);
nor U1992 (N_1992,N_1890,N_1884);
or U1993 (N_1993,N_1897,N_1930);
and U1994 (N_1994,N_1899,N_1946);
nand U1995 (N_1995,N_1948,N_1940);
and U1996 (N_1996,N_1877,N_1909);
or U1997 (N_1997,N_1909,N_1878);
nor U1998 (N_1998,N_1940,N_1949);
and U1999 (N_1999,N_1936,N_1917);
and U2000 (N_2000,N_1927,N_1944);
nand U2001 (N_2001,N_1935,N_1936);
nand U2002 (N_2002,N_1940,N_1928);
nand U2003 (N_2003,N_1941,N_1943);
nand U2004 (N_2004,N_1900,N_1947);
or U2005 (N_2005,N_1922,N_1911);
or U2006 (N_2006,N_1895,N_1905);
nor U2007 (N_2007,N_1878,N_1886);
nand U2008 (N_2008,N_1948,N_1941);
and U2009 (N_2009,N_1891,N_1942);
nor U2010 (N_2010,N_1947,N_1892);
or U2011 (N_2011,N_1896,N_1932);
nor U2012 (N_2012,N_1942,N_1890);
nor U2013 (N_2013,N_1880,N_1913);
nor U2014 (N_2014,N_1935,N_1893);
or U2015 (N_2015,N_1909,N_1902);
nand U2016 (N_2016,N_1927,N_1887);
nor U2017 (N_2017,N_1891,N_1947);
or U2018 (N_2018,N_1888,N_1948);
nor U2019 (N_2019,N_1941,N_1936);
nor U2020 (N_2020,N_1901,N_1907);
and U2021 (N_2021,N_1891,N_1876);
nor U2022 (N_2022,N_1890,N_1880);
and U2023 (N_2023,N_1894,N_1931);
or U2024 (N_2024,N_1884,N_1897);
nand U2025 (N_2025,N_2003,N_1979);
nor U2026 (N_2026,N_1957,N_1998);
and U2027 (N_2027,N_1980,N_1972);
nor U2028 (N_2028,N_1965,N_1984);
nand U2029 (N_2029,N_2009,N_2007);
or U2030 (N_2030,N_2016,N_1981);
nor U2031 (N_2031,N_2024,N_2018);
or U2032 (N_2032,N_1992,N_2013);
or U2033 (N_2033,N_1970,N_1950);
nand U2034 (N_2034,N_1990,N_2000);
nand U2035 (N_2035,N_1954,N_2005);
xor U2036 (N_2036,N_2011,N_1975);
nand U2037 (N_2037,N_2004,N_1988);
or U2038 (N_2038,N_1997,N_1960);
xnor U2039 (N_2039,N_1964,N_2014);
nor U2040 (N_2040,N_2006,N_1971);
nand U2041 (N_2041,N_1974,N_1982);
nor U2042 (N_2042,N_1962,N_1967);
nor U2043 (N_2043,N_1961,N_1958);
or U2044 (N_2044,N_1968,N_1996);
xnor U2045 (N_2045,N_2023,N_1966);
or U2046 (N_2046,N_1983,N_1999);
nor U2047 (N_2047,N_1952,N_1993);
xnor U2048 (N_2048,N_1953,N_1963);
or U2049 (N_2049,N_2022,N_1951);
nand U2050 (N_2050,N_1986,N_2017);
nor U2051 (N_2051,N_2008,N_2010);
nand U2052 (N_2052,N_1977,N_1959);
nand U2053 (N_2053,N_1955,N_1987);
nor U2054 (N_2054,N_1989,N_1976);
nand U2055 (N_2055,N_1956,N_2002);
and U2056 (N_2056,N_1973,N_2021);
and U2057 (N_2057,N_2012,N_2001);
nor U2058 (N_2058,N_1978,N_1995);
and U2059 (N_2059,N_2019,N_1985);
nand U2060 (N_2060,N_2020,N_1969);
and U2061 (N_2061,N_1994,N_2015);
xor U2062 (N_2062,N_1991,N_1962);
and U2063 (N_2063,N_1960,N_1982);
or U2064 (N_2064,N_1960,N_2010);
nand U2065 (N_2065,N_2005,N_1973);
nand U2066 (N_2066,N_1977,N_1962);
and U2067 (N_2067,N_2013,N_1980);
nand U2068 (N_2068,N_2000,N_2005);
nor U2069 (N_2069,N_1968,N_2006);
xnor U2070 (N_2070,N_1955,N_1989);
nor U2071 (N_2071,N_2004,N_1951);
and U2072 (N_2072,N_1976,N_1985);
nor U2073 (N_2073,N_2015,N_1955);
nor U2074 (N_2074,N_2006,N_1959);
and U2075 (N_2075,N_1975,N_2006);
nor U2076 (N_2076,N_1991,N_1979);
or U2077 (N_2077,N_2017,N_2006);
and U2078 (N_2078,N_1998,N_1986);
or U2079 (N_2079,N_1991,N_2004);
nand U2080 (N_2080,N_2021,N_2011);
nand U2081 (N_2081,N_1960,N_1974);
and U2082 (N_2082,N_1965,N_1975);
xor U2083 (N_2083,N_1985,N_1970);
xnor U2084 (N_2084,N_1989,N_1975);
and U2085 (N_2085,N_2016,N_1964);
nand U2086 (N_2086,N_1972,N_2020);
and U2087 (N_2087,N_1986,N_1959);
nand U2088 (N_2088,N_1988,N_1954);
nor U2089 (N_2089,N_1962,N_1963);
or U2090 (N_2090,N_1995,N_1994);
nand U2091 (N_2091,N_1964,N_1962);
xor U2092 (N_2092,N_2024,N_2021);
and U2093 (N_2093,N_1991,N_1960);
nand U2094 (N_2094,N_2011,N_2006);
nand U2095 (N_2095,N_2017,N_1953);
or U2096 (N_2096,N_2003,N_1953);
nand U2097 (N_2097,N_2020,N_1951);
xor U2098 (N_2098,N_1983,N_1991);
and U2099 (N_2099,N_1973,N_1951);
nor U2100 (N_2100,N_2057,N_2033);
and U2101 (N_2101,N_2071,N_2086);
and U2102 (N_2102,N_2065,N_2030);
nor U2103 (N_2103,N_2038,N_2081);
or U2104 (N_2104,N_2090,N_2043);
nor U2105 (N_2105,N_2062,N_2068);
and U2106 (N_2106,N_2082,N_2088);
and U2107 (N_2107,N_2069,N_2056);
or U2108 (N_2108,N_2046,N_2036);
and U2109 (N_2109,N_2059,N_2075);
or U2110 (N_2110,N_2095,N_2042);
or U2111 (N_2111,N_2049,N_2058);
nor U2112 (N_2112,N_2031,N_2091);
and U2113 (N_2113,N_2048,N_2040);
nand U2114 (N_2114,N_2029,N_2098);
xor U2115 (N_2115,N_2074,N_2050);
or U2116 (N_2116,N_2076,N_2063);
nor U2117 (N_2117,N_2099,N_2039);
nand U2118 (N_2118,N_2064,N_2089);
or U2119 (N_2119,N_2079,N_2055);
xor U2120 (N_2120,N_2053,N_2073);
nand U2121 (N_2121,N_2035,N_2034);
nor U2122 (N_2122,N_2026,N_2078);
and U2123 (N_2123,N_2077,N_2051);
xnor U2124 (N_2124,N_2096,N_2060);
nor U2125 (N_2125,N_2052,N_2066);
xor U2126 (N_2126,N_2032,N_2087);
and U2127 (N_2127,N_2044,N_2097);
or U2128 (N_2128,N_2027,N_2054);
xnor U2129 (N_2129,N_2045,N_2072);
nor U2130 (N_2130,N_2061,N_2025);
or U2131 (N_2131,N_2080,N_2028);
nand U2132 (N_2132,N_2094,N_2084);
and U2133 (N_2133,N_2093,N_2070);
and U2134 (N_2134,N_2085,N_2041);
nor U2135 (N_2135,N_2083,N_2092);
or U2136 (N_2136,N_2037,N_2047);
and U2137 (N_2137,N_2067,N_2044);
nor U2138 (N_2138,N_2029,N_2084);
nor U2139 (N_2139,N_2087,N_2084);
nor U2140 (N_2140,N_2038,N_2061);
nor U2141 (N_2141,N_2081,N_2047);
xor U2142 (N_2142,N_2067,N_2087);
nand U2143 (N_2143,N_2082,N_2064);
and U2144 (N_2144,N_2029,N_2050);
or U2145 (N_2145,N_2077,N_2031);
and U2146 (N_2146,N_2041,N_2049);
nor U2147 (N_2147,N_2028,N_2038);
nand U2148 (N_2148,N_2074,N_2036);
nand U2149 (N_2149,N_2036,N_2035);
xor U2150 (N_2150,N_2044,N_2051);
or U2151 (N_2151,N_2087,N_2088);
nand U2152 (N_2152,N_2026,N_2068);
nor U2153 (N_2153,N_2050,N_2066);
and U2154 (N_2154,N_2042,N_2040);
or U2155 (N_2155,N_2056,N_2089);
and U2156 (N_2156,N_2060,N_2081);
nor U2157 (N_2157,N_2067,N_2074);
or U2158 (N_2158,N_2053,N_2042);
nand U2159 (N_2159,N_2073,N_2038);
nand U2160 (N_2160,N_2037,N_2048);
nand U2161 (N_2161,N_2094,N_2054);
nand U2162 (N_2162,N_2047,N_2093);
or U2163 (N_2163,N_2039,N_2088);
nor U2164 (N_2164,N_2093,N_2079);
or U2165 (N_2165,N_2057,N_2088);
nor U2166 (N_2166,N_2069,N_2049);
and U2167 (N_2167,N_2056,N_2062);
xnor U2168 (N_2168,N_2027,N_2082);
and U2169 (N_2169,N_2064,N_2069);
nor U2170 (N_2170,N_2082,N_2080);
and U2171 (N_2171,N_2040,N_2064);
nand U2172 (N_2172,N_2052,N_2036);
or U2173 (N_2173,N_2036,N_2094);
nor U2174 (N_2174,N_2035,N_2081);
nand U2175 (N_2175,N_2112,N_2172);
or U2176 (N_2176,N_2159,N_2131);
or U2177 (N_2177,N_2117,N_2168);
and U2178 (N_2178,N_2106,N_2149);
and U2179 (N_2179,N_2122,N_2136);
nand U2180 (N_2180,N_2110,N_2165);
nor U2181 (N_2181,N_2114,N_2120);
and U2182 (N_2182,N_2143,N_2160);
or U2183 (N_2183,N_2140,N_2156);
or U2184 (N_2184,N_2130,N_2151);
nand U2185 (N_2185,N_2174,N_2128);
or U2186 (N_2186,N_2126,N_2105);
and U2187 (N_2187,N_2119,N_2161);
xor U2188 (N_2188,N_2148,N_2163);
xnor U2189 (N_2189,N_2135,N_2129);
and U2190 (N_2190,N_2102,N_2103);
nand U2191 (N_2191,N_2123,N_2173);
nor U2192 (N_2192,N_2157,N_2154);
nor U2193 (N_2193,N_2132,N_2153);
or U2194 (N_2194,N_2158,N_2118);
nor U2195 (N_2195,N_2167,N_2152);
nand U2196 (N_2196,N_2134,N_2164);
or U2197 (N_2197,N_2127,N_2124);
xor U2198 (N_2198,N_2145,N_2101);
and U2199 (N_2199,N_2150,N_2139);
nand U2200 (N_2200,N_2133,N_2111);
and U2201 (N_2201,N_2104,N_2155);
and U2202 (N_2202,N_2137,N_2115);
or U2203 (N_2203,N_2109,N_2125);
nor U2204 (N_2204,N_2171,N_2116);
and U2205 (N_2205,N_2147,N_2107);
nand U2206 (N_2206,N_2142,N_2141);
or U2207 (N_2207,N_2108,N_2146);
and U2208 (N_2208,N_2121,N_2170);
nor U2209 (N_2209,N_2138,N_2144);
and U2210 (N_2210,N_2166,N_2162);
nand U2211 (N_2211,N_2100,N_2113);
nor U2212 (N_2212,N_2169,N_2156);
nand U2213 (N_2213,N_2124,N_2125);
nand U2214 (N_2214,N_2140,N_2136);
or U2215 (N_2215,N_2127,N_2141);
or U2216 (N_2216,N_2149,N_2159);
and U2217 (N_2217,N_2112,N_2155);
and U2218 (N_2218,N_2166,N_2149);
nand U2219 (N_2219,N_2157,N_2140);
nor U2220 (N_2220,N_2150,N_2102);
nor U2221 (N_2221,N_2169,N_2122);
or U2222 (N_2222,N_2142,N_2151);
nand U2223 (N_2223,N_2144,N_2148);
nand U2224 (N_2224,N_2162,N_2160);
or U2225 (N_2225,N_2144,N_2160);
xnor U2226 (N_2226,N_2157,N_2114);
nor U2227 (N_2227,N_2173,N_2109);
and U2228 (N_2228,N_2153,N_2119);
xor U2229 (N_2229,N_2139,N_2157);
and U2230 (N_2230,N_2109,N_2174);
and U2231 (N_2231,N_2152,N_2109);
or U2232 (N_2232,N_2157,N_2106);
nand U2233 (N_2233,N_2122,N_2110);
nor U2234 (N_2234,N_2117,N_2103);
nand U2235 (N_2235,N_2103,N_2154);
xnor U2236 (N_2236,N_2121,N_2158);
and U2237 (N_2237,N_2130,N_2122);
and U2238 (N_2238,N_2174,N_2160);
or U2239 (N_2239,N_2102,N_2155);
and U2240 (N_2240,N_2160,N_2170);
and U2241 (N_2241,N_2144,N_2121);
nand U2242 (N_2242,N_2159,N_2166);
nor U2243 (N_2243,N_2150,N_2132);
or U2244 (N_2244,N_2138,N_2124);
xor U2245 (N_2245,N_2130,N_2174);
nor U2246 (N_2246,N_2169,N_2117);
nor U2247 (N_2247,N_2145,N_2104);
nand U2248 (N_2248,N_2138,N_2109);
and U2249 (N_2249,N_2106,N_2164);
or U2250 (N_2250,N_2224,N_2182);
or U2251 (N_2251,N_2235,N_2201);
nor U2252 (N_2252,N_2198,N_2188);
nor U2253 (N_2253,N_2227,N_2223);
or U2254 (N_2254,N_2246,N_2208);
xor U2255 (N_2255,N_2180,N_2195);
xnor U2256 (N_2256,N_2225,N_2221);
nand U2257 (N_2257,N_2215,N_2186);
nand U2258 (N_2258,N_2178,N_2245);
nand U2259 (N_2259,N_2176,N_2202);
or U2260 (N_2260,N_2241,N_2184);
or U2261 (N_2261,N_2203,N_2187);
nor U2262 (N_2262,N_2234,N_2214);
and U2263 (N_2263,N_2217,N_2238);
xnor U2264 (N_2264,N_2196,N_2213);
xnor U2265 (N_2265,N_2209,N_2249);
nor U2266 (N_2266,N_2183,N_2204);
or U2267 (N_2267,N_2248,N_2191);
nor U2268 (N_2268,N_2232,N_2226);
nand U2269 (N_2269,N_2228,N_2216);
nor U2270 (N_2270,N_2218,N_2197);
or U2271 (N_2271,N_2239,N_2212);
and U2272 (N_2272,N_2175,N_2189);
and U2273 (N_2273,N_2247,N_2236);
nor U2274 (N_2274,N_2177,N_2205);
nor U2275 (N_2275,N_2230,N_2242);
nor U2276 (N_2276,N_2233,N_2192);
nand U2277 (N_2277,N_2181,N_2244);
nand U2278 (N_2278,N_2185,N_2229);
nand U2279 (N_2279,N_2237,N_2222);
nand U2280 (N_2280,N_2219,N_2206);
and U2281 (N_2281,N_2179,N_2243);
nand U2282 (N_2282,N_2210,N_2220);
and U2283 (N_2283,N_2211,N_2194);
or U2284 (N_2284,N_2231,N_2199);
or U2285 (N_2285,N_2193,N_2207);
nor U2286 (N_2286,N_2200,N_2240);
or U2287 (N_2287,N_2190,N_2213);
and U2288 (N_2288,N_2188,N_2194);
xor U2289 (N_2289,N_2236,N_2209);
and U2290 (N_2290,N_2210,N_2204);
and U2291 (N_2291,N_2240,N_2248);
xor U2292 (N_2292,N_2239,N_2187);
nand U2293 (N_2293,N_2212,N_2238);
nand U2294 (N_2294,N_2187,N_2222);
or U2295 (N_2295,N_2243,N_2237);
nor U2296 (N_2296,N_2248,N_2224);
xor U2297 (N_2297,N_2220,N_2222);
or U2298 (N_2298,N_2230,N_2204);
and U2299 (N_2299,N_2199,N_2226);
or U2300 (N_2300,N_2217,N_2243);
and U2301 (N_2301,N_2179,N_2183);
nor U2302 (N_2302,N_2183,N_2234);
nor U2303 (N_2303,N_2201,N_2236);
nor U2304 (N_2304,N_2219,N_2240);
nor U2305 (N_2305,N_2222,N_2180);
nand U2306 (N_2306,N_2213,N_2238);
or U2307 (N_2307,N_2226,N_2204);
nand U2308 (N_2308,N_2217,N_2189);
and U2309 (N_2309,N_2188,N_2218);
and U2310 (N_2310,N_2176,N_2196);
nor U2311 (N_2311,N_2181,N_2213);
or U2312 (N_2312,N_2215,N_2178);
and U2313 (N_2313,N_2244,N_2218);
or U2314 (N_2314,N_2177,N_2248);
xnor U2315 (N_2315,N_2205,N_2216);
xnor U2316 (N_2316,N_2191,N_2192);
or U2317 (N_2317,N_2243,N_2195);
or U2318 (N_2318,N_2187,N_2179);
nand U2319 (N_2319,N_2175,N_2219);
nand U2320 (N_2320,N_2182,N_2194);
nand U2321 (N_2321,N_2198,N_2233);
or U2322 (N_2322,N_2234,N_2198);
or U2323 (N_2323,N_2220,N_2216);
nand U2324 (N_2324,N_2245,N_2244);
xor U2325 (N_2325,N_2260,N_2304);
or U2326 (N_2326,N_2297,N_2314);
nand U2327 (N_2327,N_2263,N_2295);
or U2328 (N_2328,N_2250,N_2323);
nor U2329 (N_2329,N_2266,N_2310);
or U2330 (N_2330,N_2285,N_2268);
and U2331 (N_2331,N_2267,N_2277);
xnor U2332 (N_2332,N_2256,N_2289);
or U2333 (N_2333,N_2254,N_2272);
and U2334 (N_2334,N_2296,N_2251);
and U2335 (N_2335,N_2313,N_2316);
or U2336 (N_2336,N_2273,N_2288);
xnor U2337 (N_2337,N_2294,N_2262);
nand U2338 (N_2338,N_2307,N_2286);
and U2339 (N_2339,N_2275,N_2287);
nor U2340 (N_2340,N_2322,N_2309);
and U2341 (N_2341,N_2324,N_2319);
xnor U2342 (N_2342,N_2303,N_2315);
and U2343 (N_2343,N_2305,N_2284);
xor U2344 (N_2344,N_2252,N_2261);
and U2345 (N_2345,N_2293,N_2301);
or U2346 (N_2346,N_2300,N_2258);
or U2347 (N_2347,N_2257,N_2302);
nand U2348 (N_2348,N_2255,N_2269);
nor U2349 (N_2349,N_2290,N_2274);
and U2350 (N_2350,N_2283,N_2279);
nor U2351 (N_2351,N_2271,N_2299);
and U2352 (N_2352,N_2259,N_2282);
nand U2353 (N_2353,N_2321,N_2317);
xor U2354 (N_2354,N_2281,N_2265);
nand U2355 (N_2355,N_2298,N_2320);
nand U2356 (N_2356,N_2291,N_2278);
or U2357 (N_2357,N_2292,N_2312);
and U2358 (N_2358,N_2280,N_2308);
and U2359 (N_2359,N_2318,N_2276);
or U2360 (N_2360,N_2253,N_2311);
or U2361 (N_2361,N_2306,N_2264);
or U2362 (N_2362,N_2270,N_2283);
or U2363 (N_2363,N_2290,N_2322);
or U2364 (N_2364,N_2267,N_2254);
nor U2365 (N_2365,N_2256,N_2300);
xor U2366 (N_2366,N_2255,N_2251);
or U2367 (N_2367,N_2283,N_2264);
and U2368 (N_2368,N_2275,N_2322);
nor U2369 (N_2369,N_2264,N_2260);
and U2370 (N_2370,N_2272,N_2320);
xnor U2371 (N_2371,N_2287,N_2322);
or U2372 (N_2372,N_2276,N_2308);
and U2373 (N_2373,N_2314,N_2322);
nand U2374 (N_2374,N_2279,N_2311);
xor U2375 (N_2375,N_2283,N_2306);
xor U2376 (N_2376,N_2290,N_2300);
and U2377 (N_2377,N_2278,N_2254);
and U2378 (N_2378,N_2316,N_2272);
nand U2379 (N_2379,N_2310,N_2317);
and U2380 (N_2380,N_2268,N_2278);
nand U2381 (N_2381,N_2277,N_2253);
and U2382 (N_2382,N_2266,N_2318);
nor U2383 (N_2383,N_2315,N_2257);
nor U2384 (N_2384,N_2310,N_2299);
xor U2385 (N_2385,N_2322,N_2251);
nor U2386 (N_2386,N_2306,N_2284);
and U2387 (N_2387,N_2275,N_2255);
nor U2388 (N_2388,N_2319,N_2272);
xor U2389 (N_2389,N_2308,N_2252);
xnor U2390 (N_2390,N_2294,N_2312);
and U2391 (N_2391,N_2262,N_2290);
nand U2392 (N_2392,N_2311,N_2250);
xor U2393 (N_2393,N_2257,N_2250);
and U2394 (N_2394,N_2281,N_2253);
or U2395 (N_2395,N_2303,N_2260);
and U2396 (N_2396,N_2291,N_2276);
nor U2397 (N_2397,N_2305,N_2256);
or U2398 (N_2398,N_2289,N_2275);
nor U2399 (N_2399,N_2316,N_2296);
and U2400 (N_2400,N_2332,N_2343);
or U2401 (N_2401,N_2392,N_2325);
and U2402 (N_2402,N_2349,N_2378);
xor U2403 (N_2403,N_2341,N_2394);
or U2404 (N_2404,N_2360,N_2348);
nand U2405 (N_2405,N_2331,N_2357);
and U2406 (N_2406,N_2396,N_2390);
nand U2407 (N_2407,N_2397,N_2386);
nor U2408 (N_2408,N_2372,N_2338);
xnor U2409 (N_2409,N_2369,N_2342);
or U2410 (N_2410,N_2374,N_2376);
and U2411 (N_2411,N_2379,N_2370);
or U2412 (N_2412,N_2358,N_2363);
or U2413 (N_2413,N_2365,N_2368);
xor U2414 (N_2414,N_2328,N_2337);
nand U2415 (N_2415,N_2362,N_2371);
nand U2416 (N_2416,N_2334,N_2347);
or U2417 (N_2417,N_2327,N_2329);
nand U2418 (N_2418,N_2393,N_2391);
nand U2419 (N_2419,N_2377,N_2335);
or U2420 (N_2420,N_2350,N_2336);
and U2421 (N_2421,N_2398,N_2381);
and U2422 (N_2422,N_2359,N_2354);
nor U2423 (N_2423,N_2389,N_2351);
nor U2424 (N_2424,N_2344,N_2387);
xor U2425 (N_2425,N_2333,N_2375);
nand U2426 (N_2426,N_2395,N_2361);
and U2427 (N_2427,N_2367,N_2330);
and U2428 (N_2428,N_2340,N_2346);
nor U2429 (N_2429,N_2380,N_2384);
and U2430 (N_2430,N_2339,N_2352);
nor U2431 (N_2431,N_2356,N_2399);
and U2432 (N_2432,N_2366,N_2385);
nor U2433 (N_2433,N_2388,N_2353);
and U2434 (N_2434,N_2383,N_2345);
nand U2435 (N_2435,N_2355,N_2364);
and U2436 (N_2436,N_2373,N_2382);
or U2437 (N_2437,N_2326,N_2387);
nor U2438 (N_2438,N_2358,N_2361);
and U2439 (N_2439,N_2363,N_2351);
or U2440 (N_2440,N_2398,N_2331);
or U2441 (N_2441,N_2337,N_2370);
nand U2442 (N_2442,N_2397,N_2329);
nand U2443 (N_2443,N_2392,N_2359);
or U2444 (N_2444,N_2366,N_2356);
nand U2445 (N_2445,N_2394,N_2384);
or U2446 (N_2446,N_2333,N_2369);
or U2447 (N_2447,N_2325,N_2339);
nand U2448 (N_2448,N_2325,N_2386);
xnor U2449 (N_2449,N_2382,N_2361);
and U2450 (N_2450,N_2377,N_2347);
and U2451 (N_2451,N_2383,N_2391);
and U2452 (N_2452,N_2339,N_2377);
nand U2453 (N_2453,N_2346,N_2347);
nand U2454 (N_2454,N_2383,N_2359);
or U2455 (N_2455,N_2351,N_2329);
nor U2456 (N_2456,N_2348,N_2328);
and U2457 (N_2457,N_2329,N_2356);
nor U2458 (N_2458,N_2390,N_2340);
nor U2459 (N_2459,N_2377,N_2389);
nor U2460 (N_2460,N_2349,N_2368);
or U2461 (N_2461,N_2348,N_2356);
nor U2462 (N_2462,N_2373,N_2341);
or U2463 (N_2463,N_2351,N_2343);
and U2464 (N_2464,N_2355,N_2346);
nand U2465 (N_2465,N_2396,N_2379);
nor U2466 (N_2466,N_2336,N_2388);
nand U2467 (N_2467,N_2398,N_2378);
and U2468 (N_2468,N_2371,N_2345);
and U2469 (N_2469,N_2366,N_2359);
nor U2470 (N_2470,N_2384,N_2381);
xor U2471 (N_2471,N_2399,N_2387);
nor U2472 (N_2472,N_2353,N_2334);
or U2473 (N_2473,N_2335,N_2343);
and U2474 (N_2474,N_2348,N_2350);
nor U2475 (N_2475,N_2413,N_2453);
or U2476 (N_2476,N_2406,N_2415);
and U2477 (N_2477,N_2464,N_2436);
nand U2478 (N_2478,N_2401,N_2429);
or U2479 (N_2479,N_2431,N_2434);
xnor U2480 (N_2480,N_2422,N_2457);
or U2481 (N_2481,N_2412,N_2410);
nor U2482 (N_2482,N_2441,N_2465);
nor U2483 (N_2483,N_2402,N_2435);
and U2484 (N_2484,N_2459,N_2430);
nor U2485 (N_2485,N_2473,N_2421);
nor U2486 (N_2486,N_2446,N_2428);
nor U2487 (N_2487,N_2400,N_2471);
and U2488 (N_2488,N_2423,N_2425);
nand U2489 (N_2489,N_2420,N_2449);
and U2490 (N_2490,N_2454,N_2462);
and U2491 (N_2491,N_2404,N_2463);
or U2492 (N_2492,N_2467,N_2445);
and U2493 (N_2493,N_2411,N_2414);
or U2494 (N_2494,N_2468,N_2443);
nor U2495 (N_2495,N_2437,N_2439);
or U2496 (N_2496,N_2417,N_2456);
xnor U2497 (N_2497,N_2444,N_2466);
or U2498 (N_2498,N_2427,N_2424);
xor U2499 (N_2499,N_2432,N_2450);
or U2500 (N_2500,N_2469,N_2438);
and U2501 (N_2501,N_2447,N_2416);
nor U2502 (N_2502,N_2405,N_2451);
and U2503 (N_2503,N_2408,N_2455);
xor U2504 (N_2504,N_2470,N_2409);
nand U2505 (N_2505,N_2418,N_2426);
nor U2506 (N_2506,N_2452,N_2458);
and U2507 (N_2507,N_2448,N_2407);
nand U2508 (N_2508,N_2472,N_2419);
nor U2509 (N_2509,N_2440,N_2460);
or U2510 (N_2510,N_2442,N_2403);
xnor U2511 (N_2511,N_2474,N_2461);
or U2512 (N_2512,N_2433,N_2438);
or U2513 (N_2513,N_2406,N_2404);
and U2514 (N_2514,N_2424,N_2469);
and U2515 (N_2515,N_2470,N_2472);
nor U2516 (N_2516,N_2431,N_2423);
or U2517 (N_2517,N_2469,N_2440);
nand U2518 (N_2518,N_2417,N_2444);
nor U2519 (N_2519,N_2400,N_2431);
and U2520 (N_2520,N_2424,N_2417);
or U2521 (N_2521,N_2467,N_2406);
nor U2522 (N_2522,N_2433,N_2435);
and U2523 (N_2523,N_2410,N_2417);
nand U2524 (N_2524,N_2466,N_2419);
xor U2525 (N_2525,N_2428,N_2426);
or U2526 (N_2526,N_2474,N_2469);
or U2527 (N_2527,N_2446,N_2432);
nor U2528 (N_2528,N_2452,N_2468);
nand U2529 (N_2529,N_2449,N_2448);
and U2530 (N_2530,N_2429,N_2444);
or U2531 (N_2531,N_2421,N_2457);
nor U2532 (N_2532,N_2425,N_2434);
nor U2533 (N_2533,N_2471,N_2473);
and U2534 (N_2534,N_2453,N_2469);
xor U2535 (N_2535,N_2453,N_2422);
nand U2536 (N_2536,N_2469,N_2407);
and U2537 (N_2537,N_2465,N_2424);
nand U2538 (N_2538,N_2444,N_2402);
and U2539 (N_2539,N_2467,N_2434);
nor U2540 (N_2540,N_2402,N_2422);
or U2541 (N_2541,N_2466,N_2457);
and U2542 (N_2542,N_2452,N_2428);
nor U2543 (N_2543,N_2424,N_2468);
xnor U2544 (N_2544,N_2405,N_2474);
nand U2545 (N_2545,N_2437,N_2416);
and U2546 (N_2546,N_2465,N_2438);
and U2547 (N_2547,N_2417,N_2454);
xnor U2548 (N_2548,N_2460,N_2412);
nand U2549 (N_2549,N_2448,N_2436);
and U2550 (N_2550,N_2548,N_2479);
or U2551 (N_2551,N_2516,N_2523);
nand U2552 (N_2552,N_2513,N_2543);
nor U2553 (N_2553,N_2505,N_2485);
or U2554 (N_2554,N_2480,N_2511);
nand U2555 (N_2555,N_2497,N_2507);
nand U2556 (N_2556,N_2486,N_2518);
or U2557 (N_2557,N_2489,N_2490);
xnor U2558 (N_2558,N_2476,N_2541);
nand U2559 (N_2559,N_2534,N_2501);
nand U2560 (N_2560,N_2539,N_2492);
nand U2561 (N_2561,N_2531,N_2494);
nand U2562 (N_2562,N_2524,N_2510);
nand U2563 (N_2563,N_2515,N_2483);
or U2564 (N_2564,N_2522,N_2508);
nand U2565 (N_2565,N_2509,N_2475);
or U2566 (N_2566,N_2498,N_2512);
and U2567 (N_2567,N_2477,N_2536);
nor U2568 (N_2568,N_2538,N_2530);
xnor U2569 (N_2569,N_2529,N_2482);
or U2570 (N_2570,N_2528,N_2495);
and U2571 (N_2571,N_2496,N_2514);
nor U2572 (N_2572,N_2519,N_2502);
nand U2573 (N_2573,N_2547,N_2532);
or U2574 (N_2574,N_2525,N_2527);
nor U2575 (N_2575,N_2487,N_2520);
nand U2576 (N_2576,N_2488,N_2545);
or U2577 (N_2577,N_2481,N_2526);
nand U2578 (N_2578,N_2540,N_2504);
nor U2579 (N_2579,N_2491,N_2546);
and U2580 (N_2580,N_2499,N_2533);
or U2581 (N_2581,N_2493,N_2537);
or U2582 (N_2582,N_2542,N_2549);
or U2583 (N_2583,N_2517,N_2506);
nor U2584 (N_2584,N_2521,N_2544);
nor U2585 (N_2585,N_2503,N_2484);
nor U2586 (N_2586,N_2478,N_2535);
or U2587 (N_2587,N_2500,N_2508);
or U2588 (N_2588,N_2510,N_2490);
or U2589 (N_2589,N_2479,N_2539);
nand U2590 (N_2590,N_2515,N_2507);
xor U2591 (N_2591,N_2496,N_2483);
nor U2592 (N_2592,N_2525,N_2513);
xor U2593 (N_2593,N_2509,N_2496);
nand U2594 (N_2594,N_2510,N_2484);
xor U2595 (N_2595,N_2519,N_2507);
and U2596 (N_2596,N_2506,N_2524);
or U2597 (N_2597,N_2477,N_2502);
nor U2598 (N_2598,N_2525,N_2544);
nand U2599 (N_2599,N_2484,N_2486);
nand U2600 (N_2600,N_2545,N_2530);
nand U2601 (N_2601,N_2542,N_2510);
or U2602 (N_2602,N_2514,N_2504);
and U2603 (N_2603,N_2482,N_2487);
nor U2604 (N_2604,N_2510,N_2485);
nor U2605 (N_2605,N_2499,N_2484);
or U2606 (N_2606,N_2495,N_2547);
and U2607 (N_2607,N_2522,N_2544);
or U2608 (N_2608,N_2543,N_2495);
or U2609 (N_2609,N_2541,N_2510);
xor U2610 (N_2610,N_2485,N_2496);
xnor U2611 (N_2611,N_2527,N_2516);
nor U2612 (N_2612,N_2528,N_2539);
or U2613 (N_2613,N_2527,N_2478);
or U2614 (N_2614,N_2531,N_2537);
nor U2615 (N_2615,N_2491,N_2514);
nand U2616 (N_2616,N_2516,N_2540);
xor U2617 (N_2617,N_2502,N_2523);
and U2618 (N_2618,N_2528,N_2502);
or U2619 (N_2619,N_2488,N_2515);
and U2620 (N_2620,N_2503,N_2516);
or U2621 (N_2621,N_2539,N_2503);
or U2622 (N_2622,N_2509,N_2494);
and U2623 (N_2623,N_2525,N_2549);
and U2624 (N_2624,N_2542,N_2530);
and U2625 (N_2625,N_2564,N_2596);
or U2626 (N_2626,N_2584,N_2560);
nor U2627 (N_2627,N_2594,N_2570);
or U2628 (N_2628,N_2600,N_2557);
nor U2629 (N_2629,N_2583,N_2622);
and U2630 (N_2630,N_2601,N_2613);
nand U2631 (N_2631,N_2577,N_2606);
and U2632 (N_2632,N_2565,N_2567);
and U2633 (N_2633,N_2624,N_2587);
nand U2634 (N_2634,N_2608,N_2575);
and U2635 (N_2635,N_2551,N_2597);
and U2636 (N_2636,N_2585,N_2595);
and U2637 (N_2637,N_2568,N_2593);
and U2638 (N_2638,N_2574,N_2571);
nand U2639 (N_2639,N_2604,N_2566);
nand U2640 (N_2640,N_2580,N_2623);
xnor U2641 (N_2641,N_2603,N_2619);
or U2642 (N_2642,N_2592,N_2588);
and U2643 (N_2643,N_2572,N_2569);
nor U2644 (N_2644,N_2561,N_2582);
nand U2645 (N_2645,N_2615,N_2602);
and U2646 (N_2646,N_2590,N_2618);
nand U2647 (N_2647,N_2559,N_2552);
nand U2648 (N_2648,N_2617,N_2576);
nand U2649 (N_2649,N_2578,N_2610);
and U2650 (N_2650,N_2599,N_2591);
nand U2651 (N_2651,N_2612,N_2598);
and U2652 (N_2652,N_2614,N_2553);
or U2653 (N_2653,N_2563,N_2607);
or U2654 (N_2654,N_2581,N_2620);
or U2655 (N_2655,N_2621,N_2586);
nand U2656 (N_2656,N_2554,N_2562);
nor U2657 (N_2657,N_2550,N_2611);
nor U2658 (N_2658,N_2609,N_2573);
and U2659 (N_2659,N_2556,N_2579);
nand U2660 (N_2660,N_2558,N_2555);
nand U2661 (N_2661,N_2616,N_2605);
nand U2662 (N_2662,N_2589,N_2572);
and U2663 (N_2663,N_2565,N_2623);
nand U2664 (N_2664,N_2601,N_2550);
nand U2665 (N_2665,N_2594,N_2551);
nor U2666 (N_2666,N_2590,N_2601);
nor U2667 (N_2667,N_2607,N_2570);
nor U2668 (N_2668,N_2559,N_2554);
nor U2669 (N_2669,N_2597,N_2585);
nor U2670 (N_2670,N_2550,N_2618);
or U2671 (N_2671,N_2616,N_2608);
nor U2672 (N_2672,N_2598,N_2601);
or U2673 (N_2673,N_2616,N_2590);
or U2674 (N_2674,N_2616,N_2598);
nor U2675 (N_2675,N_2601,N_2603);
nand U2676 (N_2676,N_2615,N_2555);
and U2677 (N_2677,N_2553,N_2558);
and U2678 (N_2678,N_2560,N_2618);
nor U2679 (N_2679,N_2559,N_2560);
nor U2680 (N_2680,N_2572,N_2581);
nand U2681 (N_2681,N_2591,N_2566);
nand U2682 (N_2682,N_2619,N_2602);
or U2683 (N_2683,N_2610,N_2619);
or U2684 (N_2684,N_2553,N_2578);
or U2685 (N_2685,N_2619,N_2557);
nand U2686 (N_2686,N_2624,N_2591);
and U2687 (N_2687,N_2608,N_2568);
and U2688 (N_2688,N_2553,N_2619);
and U2689 (N_2689,N_2577,N_2599);
nand U2690 (N_2690,N_2595,N_2608);
or U2691 (N_2691,N_2597,N_2577);
and U2692 (N_2692,N_2584,N_2600);
and U2693 (N_2693,N_2564,N_2610);
nand U2694 (N_2694,N_2587,N_2564);
nor U2695 (N_2695,N_2585,N_2562);
nand U2696 (N_2696,N_2603,N_2559);
nand U2697 (N_2697,N_2619,N_2617);
or U2698 (N_2698,N_2610,N_2623);
xor U2699 (N_2699,N_2616,N_2572);
nand U2700 (N_2700,N_2686,N_2631);
nor U2701 (N_2701,N_2694,N_2699);
nand U2702 (N_2702,N_2640,N_2685);
nand U2703 (N_2703,N_2677,N_2627);
and U2704 (N_2704,N_2637,N_2642);
nor U2705 (N_2705,N_2661,N_2668);
nand U2706 (N_2706,N_2643,N_2693);
or U2707 (N_2707,N_2667,N_2676);
and U2708 (N_2708,N_2690,N_2680);
nor U2709 (N_2709,N_2692,N_2626);
nand U2710 (N_2710,N_2660,N_2665);
or U2711 (N_2711,N_2664,N_2682);
and U2712 (N_2712,N_2695,N_2634);
xor U2713 (N_2713,N_2657,N_2653);
nand U2714 (N_2714,N_2641,N_2674);
nand U2715 (N_2715,N_2639,N_2673);
or U2716 (N_2716,N_2654,N_2688);
and U2717 (N_2717,N_2689,N_2629);
or U2718 (N_2718,N_2628,N_2666);
or U2719 (N_2719,N_2648,N_2652);
xnor U2720 (N_2720,N_2646,N_2679);
nand U2721 (N_2721,N_2658,N_2684);
xor U2722 (N_2722,N_2663,N_2625);
xnor U2723 (N_2723,N_2662,N_2644);
nand U2724 (N_2724,N_2696,N_2675);
nand U2725 (N_2725,N_2683,N_2638);
and U2726 (N_2726,N_2647,N_2645);
xnor U2727 (N_2727,N_2697,N_2632);
or U2728 (N_2728,N_2659,N_2672);
or U2729 (N_2729,N_2650,N_2656);
and U2730 (N_2730,N_2687,N_2681);
xnor U2731 (N_2731,N_2691,N_2651);
nand U2732 (N_2732,N_2655,N_2670);
nand U2733 (N_2733,N_2649,N_2635);
or U2734 (N_2734,N_2633,N_2630);
nand U2735 (N_2735,N_2678,N_2636);
or U2736 (N_2736,N_2669,N_2698);
nor U2737 (N_2737,N_2671,N_2658);
xor U2738 (N_2738,N_2655,N_2637);
nand U2739 (N_2739,N_2632,N_2672);
and U2740 (N_2740,N_2632,N_2690);
and U2741 (N_2741,N_2693,N_2681);
nand U2742 (N_2742,N_2691,N_2634);
xor U2743 (N_2743,N_2646,N_2677);
and U2744 (N_2744,N_2670,N_2637);
nand U2745 (N_2745,N_2685,N_2649);
nand U2746 (N_2746,N_2645,N_2633);
nand U2747 (N_2747,N_2653,N_2683);
nand U2748 (N_2748,N_2684,N_2679);
or U2749 (N_2749,N_2666,N_2691);
xnor U2750 (N_2750,N_2650,N_2699);
nor U2751 (N_2751,N_2692,N_2655);
and U2752 (N_2752,N_2675,N_2649);
and U2753 (N_2753,N_2698,N_2687);
nand U2754 (N_2754,N_2666,N_2659);
nor U2755 (N_2755,N_2694,N_2686);
nand U2756 (N_2756,N_2639,N_2653);
and U2757 (N_2757,N_2652,N_2670);
and U2758 (N_2758,N_2645,N_2673);
or U2759 (N_2759,N_2640,N_2660);
xnor U2760 (N_2760,N_2651,N_2646);
nand U2761 (N_2761,N_2645,N_2699);
nor U2762 (N_2762,N_2664,N_2689);
or U2763 (N_2763,N_2651,N_2667);
and U2764 (N_2764,N_2653,N_2681);
nand U2765 (N_2765,N_2675,N_2633);
and U2766 (N_2766,N_2699,N_2648);
nand U2767 (N_2767,N_2652,N_2688);
or U2768 (N_2768,N_2687,N_2666);
and U2769 (N_2769,N_2657,N_2673);
nand U2770 (N_2770,N_2666,N_2675);
or U2771 (N_2771,N_2699,N_2635);
xnor U2772 (N_2772,N_2645,N_2649);
or U2773 (N_2773,N_2639,N_2625);
or U2774 (N_2774,N_2629,N_2688);
or U2775 (N_2775,N_2701,N_2741);
or U2776 (N_2776,N_2756,N_2733);
nand U2777 (N_2777,N_2763,N_2712);
or U2778 (N_2778,N_2705,N_2723);
or U2779 (N_2779,N_2758,N_2702);
nor U2780 (N_2780,N_2713,N_2750);
nand U2781 (N_2781,N_2703,N_2747);
and U2782 (N_2782,N_2774,N_2765);
and U2783 (N_2783,N_2706,N_2737);
or U2784 (N_2784,N_2760,N_2743);
or U2785 (N_2785,N_2736,N_2746);
or U2786 (N_2786,N_2745,N_2764);
or U2787 (N_2787,N_2766,N_2773);
nand U2788 (N_2788,N_2748,N_2753);
nand U2789 (N_2789,N_2761,N_2725);
and U2790 (N_2790,N_2709,N_2728);
and U2791 (N_2791,N_2749,N_2731);
nor U2792 (N_2792,N_2754,N_2769);
nand U2793 (N_2793,N_2744,N_2762);
or U2794 (N_2794,N_2770,N_2704);
and U2795 (N_2795,N_2732,N_2738);
and U2796 (N_2796,N_2700,N_2716);
nor U2797 (N_2797,N_2714,N_2710);
and U2798 (N_2798,N_2771,N_2717);
and U2799 (N_2799,N_2767,N_2711);
nand U2800 (N_2800,N_2721,N_2751);
or U2801 (N_2801,N_2740,N_2734);
nor U2802 (N_2802,N_2755,N_2708);
nor U2803 (N_2803,N_2718,N_2729);
nor U2804 (N_2804,N_2757,N_2735);
nor U2805 (N_2805,N_2727,N_2722);
nand U2806 (N_2806,N_2752,N_2772);
or U2807 (N_2807,N_2707,N_2720);
or U2808 (N_2808,N_2715,N_2742);
and U2809 (N_2809,N_2724,N_2759);
xnor U2810 (N_2810,N_2768,N_2726);
nand U2811 (N_2811,N_2719,N_2739);
nor U2812 (N_2812,N_2730,N_2744);
and U2813 (N_2813,N_2701,N_2750);
nand U2814 (N_2814,N_2761,N_2759);
or U2815 (N_2815,N_2715,N_2723);
and U2816 (N_2816,N_2718,N_2736);
nor U2817 (N_2817,N_2751,N_2715);
nor U2818 (N_2818,N_2772,N_2769);
nor U2819 (N_2819,N_2755,N_2702);
nand U2820 (N_2820,N_2741,N_2714);
nor U2821 (N_2821,N_2738,N_2719);
nand U2822 (N_2822,N_2766,N_2719);
or U2823 (N_2823,N_2719,N_2714);
nor U2824 (N_2824,N_2741,N_2768);
or U2825 (N_2825,N_2748,N_2713);
nor U2826 (N_2826,N_2761,N_2703);
or U2827 (N_2827,N_2744,N_2752);
nor U2828 (N_2828,N_2730,N_2741);
nor U2829 (N_2829,N_2709,N_2713);
or U2830 (N_2830,N_2700,N_2731);
nor U2831 (N_2831,N_2731,N_2769);
and U2832 (N_2832,N_2712,N_2748);
nor U2833 (N_2833,N_2712,N_2753);
nor U2834 (N_2834,N_2754,N_2752);
xor U2835 (N_2835,N_2734,N_2771);
nor U2836 (N_2836,N_2700,N_2711);
or U2837 (N_2837,N_2759,N_2733);
nand U2838 (N_2838,N_2738,N_2757);
nor U2839 (N_2839,N_2768,N_2745);
xnor U2840 (N_2840,N_2743,N_2717);
or U2841 (N_2841,N_2703,N_2740);
xor U2842 (N_2842,N_2728,N_2733);
nand U2843 (N_2843,N_2718,N_2762);
or U2844 (N_2844,N_2773,N_2725);
or U2845 (N_2845,N_2742,N_2747);
and U2846 (N_2846,N_2767,N_2721);
nand U2847 (N_2847,N_2710,N_2718);
nor U2848 (N_2848,N_2746,N_2758);
or U2849 (N_2849,N_2740,N_2754);
or U2850 (N_2850,N_2841,N_2779);
nand U2851 (N_2851,N_2825,N_2828);
nor U2852 (N_2852,N_2846,N_2840);
or U2853 (N_2853,N_2835,N_2783);
nor U2854 (N_2854,N_2826,N_2777);
and U2855 (N_2855,N_2813,N_2847);
or U2856 (N_2856,N_2849,N_2782);
nor U2857 (N_2857,N_2792,N_2842);
and U2858 (N_2858,N_2822,N_2827);
or U2859 (N_2859,N_2816,N_2834);
xnor U2860 (N_2860,N_2839,N_2796);
and U2861 (N_2861,N_2778,N_2829);
nor U2862 (N_2862,N_2844,N_2802);
or U2863 (N_2863,N_2819,N_2807);
and U2864 (N_2864,N_2812,N_2780);
xnor U2865 (N_2865,N_2806,N_2795);
nand U2866 (N_2866,N_2784,N_2811);
or U2867 (N_2867,N_2785,N_2820);
or U2868 (N_2868,N_2838,N_2794);
nor U2869 (N_2869,N_2833,N_2824);
nor U2870 (N_2870,N_2843,N_2809);
nand U2871 (N_2871,N_2791,N_2797);
nor U2872 (N_2872,N_2800,N_2803);
and U2873 (N_2873,N_2801,N_2817);
nand U2874 (N_2874,N_2798,N_2776);
and U2875 (N_2875,N_2815,N_2799);
and U2876 (N_2876,N_2786,N_2832);
nand U2877 (N_2877,N_2830,N_2845);
nor U2878 (N_2878,N_2788,N_2789);
and U2879 (N_2879,N_2781,N_2848);
and U2880 (N_2880,N_2821,N_2787);
or U2881 (N_2881,N_2837,N_2808);
nand U2882 (N_2882,N_2775,N_2814);
and U2883 (N_2883,N_2804,N_2831);
and U2884 (N_2884,N_2823,N_2805);
nor U2885 (N_2885,N_2810,N_2836);
or U2886 (N_2886,N_2790,N_2793);
or U2887 (N_2887,N_2818,N_2779);
or U2888 (N_2888,N_2801,N_2803);
nand U2889 (N_2889,N_2818,N_2821);
and U2890 (N_2890,N_2814,N_2827);
or U2891 (N_2891,N_2808,N_2823);
nand U2892 (N_2892,N_2786,N_2829);
or U2893 (N_2893,N_2806,N_2817);
and U2894 (N_2894,N_2820,N_2788);
nor U2895 (N_2895,N_2809,N_2800);
xnor U2896 (N_2896,N_2831,N_2841);
nand U2897 (N_2897,N_2833,N_2791);
nor U2898 (N_2898,N_2780,N_2816);
nor U2899 (N_2899,N_2821,N_2829);
or U2900 (N_2900,N_2785,N_2787);
xnor U2901 (N_2901,N_2829,N_2796);
and U2902 (N_2902,N_2831,N_2778);
nand U2903 (N_2903,N_2787,N_2782);
and U2904 (N_2904,N_2814,N_2847);
nor U2905 (N_2905,N_2815,N_2813);
and U2906 (N_2906,N_2840,N_2839);
nor U2907 (N_2907,N_2843,N_2815);
nand U2908 (N_2908,N_2784,N_2814);
or U2909 (N_2909,N_2824,N_2843);
nand U2910 (N_2910,N_2846,N_2778);
and U2911 (N_2911,N_2827,N_2802);
and U2912 (N_2912,N_2798,N_2793);
and U2913 (N_2913,N_2792,N_2833);
or U2914 (N_2914,N_2848,N_2785);
and U2915 (N_2915,N_2801,N_2789);
and U2916 (N_2916,N_2818,N_2808);
and U2917 (N_2917,N_2827,N_2816);
and U2918 (N_2918,N_2848,N_2821);
nor U2919 (N_2919,N_2807,N_2827);
and U2920 (N_2920,N_2778,N_2802);
or U2921 (N_2921,N_2840,N_2825);
xnor U2922 (N_2922,N_2820,N_2799);
nor U2923 (N_2923,N_2828,N_2824);
nand U2924 (N_2924,N_2806,N_2808);
nor U2925 (N_2925,N_2888,N_2873);
nand U2926 (N_2926,N_2883,N_2870);
nor U2927 (N_2927,N_2917,N_2853);
nand U2928 (N_2928,N_2866,N_2869);
or U2929 (N_2929,N_2911,N_2913);
xor U2930 (N_2930,N_2912,N_2902);
or U2931 (N_2931,N_2905,N_2909);
xnor U2932 (N_2932,N_2879,N_2924);
xnor U2933 (N_2933,N_2858,N_2859);
or U2934 (N_2934,N_2890,N_2887);
or U2935 (N_2935,N_2881,N_2865);
and U2936 (N_2936,N_2880,N_2854);
or U2937 (N_2937,N_2907,N_2852);
and U2938 (N_2938,N_2919,N_2898);
nor U2939 (N_2939,N_2894,N_2904);
nand U2940 (N_2940,N_2860,N_2856);
nor U2941 (N_2941,N_2851,N_2885);
and U2942 (N_2942,N_2857,N_2861);
or U2943 (N_2943,N_2921,N_2906);
xnor U2944 (N_2944,N_2908,N_2876);
xor U2945 (N_2945,N_2867,N_2855);
or U2946 (N_2946,N_2886,N_2914);
nor U2947 (N_2947,N_2915,N_2862);
and U2948 (N_2948,N_2899,N_2893);
or U2949 (N_2949,N_2889,N_2920);
xnor U2950 (N_2950,N_2896,N_2850);
or U2951 (N_2951,N_2864,N_2918);
nand U2952 (N_2952,N_2877,N_2882);
and U2953 (N_2953,N_2897,N_2923);
nand U2954 (N_2954,N_2916,N_2878);
nor U2955 (N_2955,N_2874,N_2922);
nor U2956 (N_2956,N_2892,N_2901);
nor U2957 (N_2957,N_2900,N_2863);
or U2958 (N_2958,N_2895,N_2891);
nand U2959 (N_2959,N_2910,N_2868);
xor U2960 (N_2960,N_2875,N_2871);
and U2961 (N_2961,N_2903,N_2884);
and U2962 (N_2962,N_2872,N_2922);
and U2963 (N_2963,N_2855,N_2915);
and U2964 (N_2964,N_2878,N_2857);
or U2965 (N_2965,N_2886,N_2901);
nand U2966 (N_2966,N_2860,N_2853);
or U2967 (N_2967,N_2882,N_2876);
or U2968 (N_2968,N_2916,N_2914);
or U2969 (N_2969,N_2910,N_2859);
nor U2970 (N_2970,N_2866,N_2884);
or U2971 (N_2971,N_2865,N_2874);
nor U2972 (N_2972,N_2859,N_2902);
and U2973 (N_2973,N_2901,N_2867);
nand U2974 (N_2974,N_2884,N_2850);
or U2975 (N_2975,N_2898,N_2881);
nand U2976 (N_2976,N_2891,N_2892);
and U2977 (N_2977,N_2890,N_2913);
nor U2978 (N_2978,N_2904,N_2920);
nand U2979 (N_2979,N_2873,N_2900);
and U2980 (N_2980,N_2880,N_2894);
xnor U2981 (N_2981,N_2878,N_2923);
nor U2982 (N_2982,N_2909,N_2864);
nand U2983 (N_2983,N_2890,N_2875);
nand U2984 (N_2984,N_2874,N_2897);
and U2985 (N_2985,N_2863,N_2868);
nor U2986 (N_2986,N_2860,N_2876);
and U2987 (N_2987,N_2909,N_2852);
nor U2988 (N_2988,N_2909,N_2911);
or U2989 (N_2989,N_2924,N_2862);
and U2990 (N_2990,N_2888,N_2860);
or U2991 (N_2991,N_2854,N_2855);
or U2992 (N_2992,N_2880,N_2852);
nand U2993 (N_2993,N_2908,N_2915);
nor U2994 (N_2994,N_2898,N_2913);
nand U2995 (N_2995,N_2862,N_2873);
or U2996 (N_2996,N_2871,N_2907);
and U2997 (N_2997,N_2851,N_2875);
nor U2998 (N_2998,N_2902,N_2884);
nand U2999 (N_2999,N_2869,N_2862);
nor UO_0 (O_0,N_2987,N_2995);
xnor UO_1 (O_1,N_2941,N_2933);
nor UO_2 (O_2,N_2925,N_2952);
nand UO_3 (O_3,N_2955,N_2953);
nor UO_4 (O_4,N_2977,N_2956);
xnor UO_5 (O_5,N_2958,N_2939);
or UO_6 (O_6,N_2997,N_2926);
or UO_7 (O_7,N_2972,N_2982);
nor UO_8 (O_8,N_2971,N_2947);
or UO_9 (O_9,N_2936,N_2979);
and UO_10 (O_10,N_2950,N_2963);
or UO_11 (O_11,N_2994,N_2991);
nand UO_12 (O_12,N_2998,N_2988);
nand UO_13 (O_13,N_2962,N_2993);
and UO_14 (O_14,N_2992,N_2937);
nand UO_15 (O_15,N_2951,N_2996);
nand UO_16 (O_16,N_2967,N_2970);
nor UO_17 (O_17,N_2940,N_2957);
nand UO_18 (O_18,N_2976,N_2990);
and UO_19 (O_19,N_2966,N_2983);
nor UO_20 (O_20,N_2949,N_2999);
nand UO_21 (O_21,N_2969,N_2964);
nor UO_22 (O_22,N_2927,N_2980);
xnor UO_23 (O_23,N_2965,N_2961);
or UO_24 (O_24,N_2981,N_2942);
nand UO_25 (O_25,N_2948,N_2986);
nand UO_26 (O_26,N_2929,N_2978);
nand UO_27 (O_27,N_2975,N_2932);
nand UO_28 (O_28,N_2974,N_2938);
xor UO_29 (O_29,N_2935,N_2960);
or UO_30 (O_30,N_2945,N_2984);
xor UO_31 (O_31,N_2930,N_2931);
xor UO_32 (O_32,N_2934,N_2946);
nor UO_33 (O_33,N_2973,N_2944);
or UO_34 (O_34,N_2959,N_2954);
xnor UO_35 (O_35,N_2985,N_2928);
nor UO_36 (O_36,N_2989,N_2943);
nand UO_37 (O_37,N_2968,N_2948);
nor UO_38 (O_38,N_2952,N_2989);
nor UO_39 (O_39,N_2927,N_2995);
nand UO_40 (O_40,N_2959,N_2958);
or UO_41 (O_41,N_2946,N_2992);
nand UO_42 (O_42,N_2983,N_2998);
nor UO_43 (O_43,N_2977,N_2967);
nor UO_44 (O_44,N_2954,N_2952);
or UO_45 (O_45,N_2976,N_2968);
or UO_46 (O_46,N_2957,N_2928);
xor UO_47 (O_47,N_2959,N_2974);
and UO_48 (O_48,N_2953,N_2958);
or UO_49 (O_49,N_2956,N_2948);
xor UO_50 (O_50,N_2930,N_2993);
xor UO_51 (O_51,N_2974,N_2994);
nand UO_52 (O_52,N_2948,N_2959);
and UO_53 (O_53,N_2977,N_2976);
nand UO_54 (O_54,N_2997,N_2973);
nand UO_55 (O_55,N_2943,N_2961);
and UO_56 (O_56,N_2939,N_2926);
and UO_57 (O_57,N_2925,N_2926);
and UO_58 (O_58,N_2951,N_2988);
xnor UO_59 (O_59,N_2938,N_2989);
and UO_60 (O_60,N_2966,N_2948);
or UO_61 (O_61,N_2968,N_2987);
and UO_62 (O_62,N_2965,N_2981);
nor UO_63 (O_63,N_2936,N_2955);
nor UO_64 (O_64,N_2928,N_2961);
xor UO_65 (O_65,N_2988,N_2977);
nor UO_66 (O_66,N_2974,N_2929);
and UO_67 (O_67,N_2947,N_2933);
xnor UO_68 (O_68,N_2993,N_2961);
nand UO_69 (O_69,N_2926,N_2974);
or UO_70 (O_70,N_2986,N_2959);
and UO_71 (O_71,N_2928,N_2956);
nand UO_72 (O_72,N_2952,N_2926);
nor UO_73 (O_73,N_2943,N_2968);
and UO_74 (O_74,N_2942,N_2935);
or UO_75 (O_75,N_2964,N_2973);
nor UO_76 (O_76,N_2930,N_2929);
nor UO_77 (O_77,N_2950,N_2959);
and UO_78 (O_78,N_2940,N_2973);
nor UO_79 (O_79,N_2982,N_2939);
nor UO_80 (O_80,N_2968,N_2956);
and UO_81 (O_81,N_2964,N_2948);
or UO_82 (O_82,N_2984,N_2950);
xor UO_83 (O_83,N_2955,N_2927);
and UO_84 (O_84,N_2975,N_2988);
or UO_85 (O_85,N_2929,N_2953);
xor UO_86 (O_86,N_2970,N_2939);
or UO_87 (O_87,N_2944,N_2975);
nor UO_88 (O_88,N_2981,N_2991);
or UO_89 (O_89,N_2945,N_2994);
nor UO_90 (O_90,N_2964,N_2994);
nor UO_91 (O_91,N_2955,N_2994);
nor UO_92 (O_92,N_2933,N_2932);
nor UO_93 (O_93,N_2971,N_2998);
nor UO_94 (O_94,N_2972,N_2958);
and UO_95 (O_95,N_2994,N_2969);
nand UO_96 (O_96,N_2949,N_2956);
nor UO_97 (O_97,N_2987,N_2994);
and UO_98 (O_98,N_2934,N_2977);
nand UO_99 (O_99,N_2947,N_2961);
and UO_100 (O_100,N_2965,N_2983);
or UO_101 (O_101,N_2982,N_2985);
xnor UO_102 (O_102,N_2933,N_2949);
or UO_103 (O_103,N_2946,N_2977);
nor UO_104 (O_104,N_2960,N_2976);
nor UO_105 (O_105,N_2927,N_2962);
xnor UO_106 (O_106,N_2935,N_2986);
nor UO_107 (O_107,N_2942,N_2993);
nor UO_108 (O_108,N_2995,N_2929);
xor UO_109 (O_109,N_2992,N_2976);
or UO_110 (O_110,N_2950,N_2999);
nand UO_111 (O_111,N_2937,N_2932);
nand UO_112 (O_112,N_2987,N_2979);
nor UO_113 (O_113,N_2967,N_2941);
nor UO_114 (O_114,N_2931,N_2934);
and UO_115 (O_115,N_2977,N_2968);
xnor UO_116 (O_116,N_2977,N_2964);
or UO_117 (O_117,N_2970,N_2954);
or UO_118 (O_118,N_2968,N_2974);
and UO_119 (O_119,N_2963,N_2964);
or UO_120 (O_120,N_2931,N_2973);
xnor UO_121 (O_121,N_2926,N_2930);
nand UO_122 (O_122,N_2982,N_2927);
nor UO_123 (O_123,N_2946,N_2961);
nand UO_124 (O_124,N_2954,N_2971);
or UO_125 (O_125,N_2949,N_2931);
or UO_126 (O_126,N_2985,N_2953);
and UO_127 (O_127,N_2995,N_2932);
nand UO_128 (O_128,N_2990,N_2963);
and UO_129 (O_129,N_2957,N_2955);
nor UO_130 (O_130,N_2954,N_2949);
or UO_131 (O_131,N_2946,N_2966);
and UO_132 (O_132,N_2988,N_2980);
and UO_133 (O_133,N_2974,N_2935);
nor UO_134 (O_134,N_2979,N_2954);
or UO_135 (O_135,N_2956,N_2950);
and UO_136 (O_136,N_2950,N_2987);
or UO_137 (O_137,N_2957,N_2979);
nor UO_138 (O_138,N_2956,N_2974);
and UO_139 (O_139,N_2949,N_2939);
nand UO_140 (O_140,N_2933,N_2953);
or UO_141 (O_141,N_2981,N_2957);
nand UO_142 (O_142,N_2936,N_2952);
nor UO_143 (O_143,N_2964,N_2970);
or UO_144 (O_144,N_2930,N_2994);
and UO_145 (O_145,N_2941,N_2976);
and UO_146 (O_146,N_2960,N_2965);
nand UO_147 (O_147,N_2981,N_2954);
or UO_148 (O_148,N_2969,N_2987);
and UO_149 (O_149,N_2937,N_2941);
and UO_150 (O_150,N_2990,N_2977);
and UO_151 (O_151,N_2939,N_2954);
nor UO_152 (O_152,N_2965,N_2963);
and UO_153 (O_153,N_2982,N_2956);
nor UO_154 (O_154,N_2947,N_2925);
nor UO_155 (O_155,N_2999,N_2961);
or UO_156 (O_156,N_2964,N_2939);
and UO_157 (O_157,N_2954,N_2976);
nor UO_158 (O_158,N_2949,N_2986);
xnor UO_159 (O_159,N_2994,N_2925);
and UO_160 (O_160,N_2962,N_2928);
and UO_161 (O_161,N_2951,N_2971);
nand UO_162 (O_162,N_2980,N_2936);
nand UO_163 (O_163,N_2942,N_2971);
and UO_164 (O_164,N_2964,N_2983);
nand UO_165 (O_165,N_2937,N_2978);
and UO_166 (O_166,N_2976,N_2934);
nand UO_167 (O_167,N_2994,N_2977);
nand UO_168 (O_168,N_2950,N_2939);
or UO_169 (O_169,N_2959,N_2968);
nand UO_170 (O_170,N_2927,N_2971);
and UO_171 (O_171,N_2967,N_2992);
and UO_172 (O_172,N_2928,N_2952);
nand UO_173 (O_173,N_2938,N_2939);
nor UO_174 (O_174,N_2982,N_2953);
and UO_175 (O_175,N_2974,N_2936);
or UO_176 (O_176,N_2934,N_2991);
nand UO_177 (O_177,N_2964,N_2979);
or UO_178 (O_178,N_2939,N_2927);
nand UO_179 (O_179,N_2971,N_2991);
nand UO_180 (O_180,N_2951,N_2967);
xor UO_181 (O_181,N_2967,N_2999);
nor UO_182 (O_182,N_2935,N_2964);
or UO_183 (O_183,N_2931,N_2992);
or UO_184 (O_184,N_2946,N_2980);
or UO_185 (O_185,N_2943,N_2948);
nor UO_186 (O_186,N_2996,N_2971);
nand UO_187 (O_187,N_2978,N_2936);
and UO_188 (O_188,N_2927,N_2992);
nor UO_189 (O_189,N_2956,N_2976);
and UO_190 (O_190,N_2961,N_2949);
or UO_191 (O_191,N_2961,N_2931);
or UO_192 (O_192,N_2969,N_2946);
or UO_193 (O_193,N_2925,N_2976);
and UO_194 (O_194,N_2950,N_2962);
and UO_195 (O_195,N_2995,N_2947);
and UO_196 (O_196,N_2952,N_2972);
nor UO_197 (O_197,N_2937,N_2961);
nor UO_198 (O_198,N_2985,N_2954);
nand UO_199 (O_199,N_2988,N_2961);
or UO_200 (O_200,N_2985,N_2976);
and UO_201 (O_201,N_2989,N_2941);
nand UO_202 (O_202,N_2981,N_2973);
xor UO_203 (O_203,N_2951,N_2931);
or UO_204 (O_204,N_2928,N_2947);
xor UO_205 (O_205,N_2971,N_2931);
or UO_206 (O_206,N_2981,N_2987);
nand UO_207 (O_207,N_2984,N_2955);
nor UO_208 (O_208,N_2964,N_2965);
nand UO_209 (O_209,N_2927,N_2949);
nand UO_210 (O_210,N_2964,N_2986);
and UO_211 (O_211,N_2956,N_2972);
and UO_212 (O_212,N_2930,N_2945);
and UO_213 (O_213,N_2960,N_2952);
and UO_214 (O_214,N_2959,N_2973);
nand UO_215 (O_215,N_2992,N_2981);
or UO_216 (O_216,N_2992,N_2962);
nand UO_217 (O_217,N_2949,N_2938);
nand UO_218 (O_218,N_2989,N_2950);
nand UO_219 (O_219,N_2962,N_2983);
nand UO_220 (O_220,N_2947,N_2967);
nor UO_221 (O_221,N_2926,N_2988);
and UO_222 (O_222,N_2964,N_2968);
or UO_223 (O_223,N_2972,N_2980);
nor UO_224 (O_224,N_2977,N_2959);
and UO_225 (O_225,N_2989,N_2954);
nand UO_226 (O_226,N_2982,N_2994);
or UO_227 (O_227,N_2965,N_2954);
nor UO_228 (O_228,N_2925,N_2990);
or UO_229 (O_229,N_2997,N_2965);
or UO_230 (O_230,N_2957,N_2970);
or UO_231 (O_231,N_2984,N_2960);
and UO_232 (O_232,N_2945,N_2975);
xnor UO_233 (O_233,N_2972,N_2962);
nand UO_234 (O_234,N_2948,N_2945);
nor UO_235 (O_235,N_2952,N_2982);
xor UO_236 (O_236,N_2932,N_2934);
nand UO_237 (O_237,N_2941,N_2994);
and UO_238 (O_238,N_2944,N_2995);
nor UO_239 (O_239,N_2980,N_2954);
or UO_240 (O_240,N_2944,N_2996);
or UO_241 (O_241,N_2992,N_2930);
nor UO_242 (O_242,N_2976,N_2937);
nor UO_243 (O_243,N_2982,N_2962);
or UO_244 (O_244,N_2982,N_2980);
and UO_245 (O_245,N_2959,N_2938);
nor UO_246 (O_246,N_2972,N_2977);
and UO_247 (O_247,N_2999,N_2947);
xor UO_248 (O_248,N_2937,N_2984);
nor UO_249 (O_249,N_2940,N_2963);
nor UO_250 (O_250,N_2994,N_2950);
nor UO_251 (O_251,N_2990,N_2926);
nor UO_252 (O_252,N_2953,N_2932);
xor UO_253 (O_253,N_2963,N_2996);
or UO_254 (O_254,N_2944,N_2926);
and UO_255 (O_255,N_2981,N_2970);
nand UO_256 (O_256,N_2966,N_2931);
nor UO_257 (O_257,N_2966,N_2984);
xor UO_258 (O_258,N_2955,N_2944);
xor UO_259 (O_259,N_2989,N_2986);
or UO_260 (O_260,N_2992,N_2989);
and UO_261 (O_261,N_2940,N_2925);
nand UO_262 (O_262,N_2935,N_2998);
nor UO_263 (O_263,N_2967,N_2968);
nand UO_264 (O_264,N_2934,N_2959);
nand UO_265 (O_265,N_2946,N_2929);
nand UO_266 (O_266,N_2990,N_2973);
nor UO_267 (O_267,N_2939,N_2946);
nor UO_268 (O_268,N_2990,N_2997);
or UO_269 (O_269,N_2931,N_2938);
and UO_270 (O_270,N_2987,N_2925);
xor UO_271 (O_271,N_2961,N_2953);
nand UO_272 (O_272,N_2929,N_2933);
or UO_273 (O_273,N_2974,N_2943);
nor UO_274 (O_274,N_2978,N_2982);
nand UO_275 (O_275,N_2992,N_2936);
nand UO_276 (O_276,N_2978,N_2925);
nor UO_277 (O_277,N_2997,N_2933);
xor UO_278 (O_278,N_2956,N_2988);
nor UO_279 (O_279,N_2994,N_2996);
or UO_280 (O_280,N_2998,N_2930);
nand UO_281 (O_281,N_2999,N_2992);
nor UO_282 (O_282,N_2959,N_2978);
nor UO_283 (O_283,N_2977,N_2958);
and UO_284 (O_284,N_2937,N_2948);
or UO_285 (O_285,N_2982,N_2947);
xnor UO_286 (O_286,N_2982,N_2988);
and UO_287 (O_287,N_2998,N_2991);
and UO_288 (O_288,N_2931,N_2935);
and UO_289 (O_289,N_2983,N_2956);
or UO_290 (O_290,N_2988,N_2954);
nand UO_291 (O_291,N_2950,N_2932);
nand UO_292 (O_292,N_2940,N_2986);
nand UO_293 (O_293,N_2972,N_2995);
or UO_294 (O_294,N_2931,N_2970);
and UO_295 (O_295,N_2943,N_2977);
and UO_296 (O_296,N_2991,N_2941);
xor UO_297 (O_297,N_2959,N_2928);
or UO_298 (O_298,N_2997,N_2970);
and UO_299 (O_299,N_2991,N_2972);
nand UO_300 (O_300,N_2937,N_2983);
nor UO_301 (O_301,N_2956,N_2964);
xor UO_302 (O_302,N_2956,N_2929);
nor UO_303 (O_303,N_2958,N_2996);
and UO_304 (O_304,N_2980,N_2948);
or UO_305 (O_305,N_2997,N_2957);
nor UO_306 (O_306,N_2963,N_2981);
and UO_307 (O_307,N_2958,N_2941);
nand UO_308 (O_308,N_2953,N_2981);
and UO_309 (O_309,N_2944,N_2949);
nand UO_310 (O_310,N_2980,N_2928);
and UO_311 (O_311,N_2978,N_2975);
xor UO_312 (O_312,N_2966,N_2991);
xnor UO_313 (O_313,N_2936,N_2977);
and UO_314 (O_314,N_2989,N_2942);
nor UO_315 (O_315,N_2980,N_2981);
and UO_316 (O_316,N_2934,N_2954);
and UO_317 (O_317,N_2960,N_2943);
xor UO_318 (O_318,N_2965,N_2944);
xnor UO_319 (O_319,N_2967,N_2932);
and UO_320 (O_320,N_2980,N_2997);
or UO_321 (O_321,N_2952,N_2953);
nand UO_322 (O_322,N_2993,N_2980);
or UO_323 (O_323,N_2934,N_2972);
or UO_324 (O_324,N_2986,N_2934);
and UO_325 (O_325,N_2992,N_2934);
and UO_326 (O_326,N_2976,N_2943);
nand UO_327 (O_327,N_2931,N_2985);
or UO_328 (O_328,N_2946,N_2952);
nand UO_329 (O_329,N_2951,N_2930);
and UO_330 (O_330,N_2927,N_2952);
and UO_331 (O_331,N_2928,N_2974);
nor UO_332 (O_332,N_2931,N_2998);
nand UO_333 (O_333,N_2975,N_2957);
nand UO_334 (O_334,N_2925,N_2937);
and UO_335 (O_335,N_2981,N_2947);
or UO_336 (O_336,N_2987,N_2966);
nor UO_337 (O_337,N_2948,N_2979);
nor UO_338 (O_338,N_2928,N_2990);
or UO_339 (O_339,N_2934,N_2952);
nor UO_340 (O_340,N_2944,N_2980);
nand UO_341 (O_341,N_2955,N_2971);
nor UO_342 (O_342,N_2965,N_2938);
nand UO_343 (O_343,N_2962,N_2940);
or UO_344 (O_344,N_2997,N_2928);
nand UO_345 (O_345,N_2971,N_2980);
and UO_346 (O_346,N_2982,N_2983);
and UO_347 (O_347,N_2997,N_2945);
nand UO_348 (O_348,N_2980,N_2986);
or UO_349 (O_349,N_2965,N_2933);
or UO_350 (O_350,N_2944,N_2945);
or UO_351 (O_351,N_2951,N_2943);
and UO_352 (O_352,N_2969,N_2998);
and UO_353 (O_353,N_2966,N_2952);
or UO_354 (O_354,N_2986,N_2960);
nor UO_355 (O_355,N_2958,N_2999);
and UO_356 (O_356,N_2939,N_2956);
nor UO_357 (O_357,N_2936,N_2944);
and UO_358 (O_358,N_2961,N_2972);
nand UO_359 (O_359,N_2941,N_2959);
or UO_360 (O_360,N_2953,N_2991);
or UO_361 (O_361,N_2955,N_2985);
nor UO_362 (O_362,N_2929,N_2990);
and UO_363 (O_363,N_2938,N_2996);
nand UO_364 (O_364,N_2946,N_2958);
and UO_365 (O_365,N_2933,N_2989);
and UO_366 (O_366,N_2939,N_2955);
or UO_367 (O_367,N_2973,N_2999);
nor UO_368 (O_368,N_2927,N_2968);
nand UO_369 (O_369,N_2976,N_2975);
and UO_370 (O_370,N_2988,N_2952);
or UO_371 (O_371,N_2938,N_2935);
nand UO_372 (O_372,N_2929,N_2979);
or UO_373 (O_373,N_2925,N_2972);
or UO_374 (O_374,N_2989,N_2971);
nor UO_375 (O_375,N_2989,N_2928);
and UO_376 (O_376,N_2927,N_2976);
and UO_377 (O_377,N_2960,N_2945);
nand UO_378 (O_378,N_2990,N_2979);
nand UO_379 (O_379,N_2970,N_2978);
or UO_380 (O_380,N_2989,N_2934);
nand UO_381 (O_381,N_2999,N_2977);
xnor UO_382 (O_382,N_2964,N_2958);
or UO_383 (O_383,N_2975,N_2956);
nor UO_384 (O_384,N_2938,N_2937);
or UO_385 (O_385,N_2999,N_2966);
xnor UO_386 (O_386,N_2940,N_2966);
or UO_387 (O_387,N_2988,N_2949);
or UO_388 (O_388,N_2983,N_2970);
nor UO_389 (O_389,N_2956,N_2947);
nor UO_390 (O_390,N_2987,N_2951);
and UO_391 (O_391,N_2948,N_2941);
and UO_392 (O_392,N_2979,N_2956);
xor UO_393 (O_393,N_2962,N_2970);
nand UO_394 (O_394,N_2952,N_2941);
or UO_395 (O_395,N_2993,N_2971);
and UO_396 (O_396,N_2948,N_2946);
xor UO_397 (O_397,N_2932,N_2939);
and UO_398 (O_398,N_2956,N_2945);
nand UO_399 (O_399,N_2956,N_2980);
and UO_400 (O_400,N_2933,N_2945);
and UO_401 (O_401,N_2939,N_2951);
and UO_402 (O_402,N_2966,N_2980);
or UO_403 (O_403,N_2930,N_2948);
and UO_404 (O_404,N_2937,N_2965);
or UO_405 (O_405,N_2930,N_2966);
or UO_406 (O_406,N_2970,N_2968);
and UO_407 (O_407,N_2961,N_2976);
and UO_408 (O_408,N_2947,N_2969);
nor UO_409 (O_409,N_2973,N_2937);
or UO_410 (O_410,N_2940,N_2993);
and UO_411 (O_411,N_2925,N_2930);
nand UO_412 (O_412,N_2998,N_2987);
nand UO_413 (O_413,N_2962,N_2981);
or UO_414 (O_414,N_2958,N_2987);
and UO_415 (O_415,N_2928,N_2936);
nand UO_416 (O_416,N_2970,N_2953);
and UO_417 (O_417,N_2975,N_2968);
or UO_418 (O_418,N_2936,N_2993);
and UO_419 (O_419,N_2984,N_2939);
nor UO_420 (O_420,N_2995,N_2973);
or UO_421 (O_421,N_2990,N_2947);
nand UO_422 (O_422,N_2946,N_2976);
and UO_423 (O_423,N_2983,N_2925);
xor UO_424 (O_424,N_2933,N_2942);
nand UO_425 (O_425,N_2970,N_2932);
nor UO_426 (O_426,N_2925,N_2938);
nor UO_427 (O_427,N_2963,N_2926);
or UO_428 (O_428,N_2936,N_2956);
and UO_429 (O_429,N_2950,N_2946);
xnor UO_430 (O_430,N_2951,N_2955);
nand UO_431 (O_431,N_2940,N_2991);
and UO_432 (O_432,N_2925,N_2929);
or UO_433 (O_433,N_2967,N_2990);
nand UO_434 (O_434,N_2947,N_2948);
nand UO_435 (O_435,N_2950,N_2992);
nor UO_436 (O_436,N_2956,N_2951);
nor UO_437 (O_437,N_2929,N_2955);
nor UO_438 (O_438,N_2956,N_2944);
nor UO_439 (O_439,N_2961,N_2973);
nor UO_440 (O_440,N_2954,N_2942);
nand UO_441 (O_441,N_2985,N_2999);
nor UO_442 (O_442,N_2961,N_2958);
nand UO_443 (O_443,N_2998,N_2960);
nand UO_444 (O_444,N_2985,N_2944);
and UO_445 (O_445,N_2971,N_2964);
nor UO_446 (O_446,N_2955,N_2973);
and UO_447 (O_447,N_2998,N_2973);
nor UO_448 (O_448,N_2986,N_2947);
nand UO_449 (O_449,N_2932,N_2981);
xnor UO_450 (O_450,N_2990,N_2971);
xnor UO_451 (O_451,N_2977,N_2938);
nand UO_452 (O_452,N_2963,N_2994);
nor UO_453 (O_453,N_2964,N_2944);
or UO_454 (O_454,N_2976,N_2986);
nor UO_455 (O_455,N_2977,N_2945);
nand UO_456 (O_456,N_2969,N_2929);
and UO_457 (O_457,N_2990,N_2933);
nor UO_458 (O_458,N_2947,N_2985);
nor UO_459 (O_459,N_2967,N_2975);
or UO_460 (O_460,N_2935,N_2958);
nor UO_461 (O_461,N_2998,N_2989);
and UO_462 (O_462,N_2988,N_2962);
nor UO_463 (O_463,N_2936,N_2991);
xnor UO_464 (O_464,N_2974,N_2984);
or UO_465 (O_465,N_2927,N_2961);
nor UO_466 (O_466,N_2957,N_2992);
and UO_467 (O_467,N_2926,N_2941);
and UO_468 (O_468,N_2925,N_2946);
or UO_469 (O_469,N_2946,N_2986);
and UO_470 (O_470,N_2943,N_2965);
nor UO_471 (O_471,N_2953,N_2930);
nand UO_472 (O_472,N_2941,N_2995);
nand UO_473 (O_473,N_2936,N_2994);
nor UO_474 (O_474,N_2963,N_2984);
or UO_475 (O_475,N_2947,N_2994);
nand UO_476 (O_476,N_2954,N_2926);
or UO_477 (O_477,N_2926,N_2977);
and UO_478 (O_478,N_2978,N_2949);
nor UO_479 (O_479,N_2952,N_2991);
or UO_480 (O_480,N_2964,N_2942);
nor UO_481 (O_481,N_2962,N_2974);
xnor UO_482 (O_482,N_2969,N_2934);
nand UO_483 (O_483,N_2967,N_2942);
or UO_484 (O_484,N_2932,N_2948);
xor UO_485 (O_485,N_2981,N_2952);
or UO_486 (O_486,N_2938,N_2963);
nand UO_487 (O_487,N_2932,N_2980);
nor UO_488 (O_488,N_2934,N_2942);
nor UO_489 (O_489,N_2951,N_2936);
and UO_490 (O_490,N_2978,N_2928);
nand UO_491 (O_491,N_2994,N_2926);
nand UO_492 (O_492,N_2932,N_2965);
or UO_493 (O_493,N_2937,N_2951);
nor UO_494 (O_494,N_2978,N_2987);
and UO_495 (O_495,N_2943,N_2985);
nor UO_496 (O_496,N_2935,N_2944);
nand UO_497 (O_497,N_2984,N_2998);
nand UO_498 (O_498,N_2999,N_2978);
or UO_499 (O_499,N_2993,N_2975);
endmodule