module basic_750_5000_1000_50_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_595,In_540);
or U1 (N_1,In_182,In_127);
or U2 (N_2,In_747,In_273);
nand U3 (N_3,In_106,In_296);
xnor U4 (N_4,In_435,In_52);
or U5 (N_5,In_268,In_159);
and U6 (N_6,In_627,In_316);
or U7 (N_7,In_277,In_537);
xor U8 (N_8,In_594,In_348);
nand U9 (N_9,In_513,In_489);
nor U10 (N_10,In_254,In_449);
or U11 (N_11,In_333,In_572);
nand U12 (N_12,In_620,In_745);
nand U13 (N_13,In_560,In_45);
nor U14 (N_14,In_351,In_675);
xor U15 (N_15,In_553,In_37);
or U16 (N_16,In_591,In_456);
or U17 (N_17,In_686,In_77);
nand U18 (N_18,In_68,In_547);
and U19 (N_19,In_415,In_196);
and U20 (N_20,In_364,In_311);
or U21 (N_21,In_232,In_154);
nand U22 (N_22,In_377,In_243);
or U23 (N_23,In_372,In_567);
and U24 (N_24,In_429,In_169);
nor U25 (N_25,In_42,In_62);
or U26 (N_26,In_26,In_242);
and U27 (N_27,In_302,In_576);
nor U28 (N_28,In_163,In_423);
nor U29 (N_29,In_331,In_667);
nand U30 (N_30,In_198,In_214);
and U31 (N_31,In_624,In_186);
or U32 (N_32,In_500,In_707);
and U33 (N_33,In_211,In_293);
nand U34 (N_34,In_12,In_610);
xor U35 (N_35,In_663,In_561);
or U36 (N_36,In_5,In_225);
nand U37 (N_37,In_230,In_668);
or U38 (N_38,In_693,In_278);
or U39 (N_39,In_286,In_116);
nand U40 (N_40,In_137,In_358);
xor U41 (N_41,In_460,In_57);
and U42 (N_42,In_29,In_521);
nand U43 (N_43,In_212,In_501);
xnor U44 (N_44,In_111,In_734);
or U45 (N_45,In_644,In_19);
xor U46 (N_46,In_607,In_606);
nand U47 (N_47,In_365,In_704);
nand U48 (N_48,In_340,In_475);
nand U49 (N_49,In_265,In_120);
or U50 (N_50,In_447,In_541);
or U51 (N_51,In_643,In_147);
and U52 (N_52,In_307,In_162);
and U53 (N_53,In_164,In_24);
nand U54 (N_54,In_744,In_430);
xnor U55 (N_55,In_176,In_95);
nand U56 (N_56,In_432,In_71);
or U57 (N_57,In_258,In_319);
and U58 (N_58,In_695,In_35);
or U59 (N_59,In_395,In_46);
nor U60 (N_60,In_532,In_203);
and U61 (N_61,In_584,In_596);
or U62 (N_62,In_244,In_464);
or U63 (N_63,In_231,In_51);
nor U64 (N_64,In_226,In_574);
xor U65 (N_65,In_27,In_115);
or U66 (N_66,In_701,In_603);
nand U67 (N_67,In_128,In_180);
xor U68 (N_68,In_93,In_674);
nor U69 (N_69,In_132,In_403);
nand U70 (N_70,In_321,In_343);
and U71 (N_71,In_65,In_17);
and U72 (N_72,In_253,In_538);
nand U73 (N_73,In_641,In_251);
and U74 (N_74,In_405,In_376);
and U75 (N_75,In_109,In_91);
or U76 (N_76,In_285,In_488);
nor U77 (N_77,In_290,In_313);
or U78 (N_78,In_737,In_310);
nand U79 (N_79,In_6,In_505);
xor U80 (N_80,In_483,In_563);
nor U81 (N_81,In_528,In_61);
and U82 (N_82,In_201,In_548);
nand U83 (N_83,In_558,In_660);
nand U84 (N_84,In_438,In_288);
nor U85 (N_85,In_329,In_729);
nand U86 (N_86,In_472,In_213);
or U87 (N_87,In_291,In_525);
nand U88 (N_88,In_347,In_205);
nand U89 (N_89,In_317,In_129);
or U90 (N_90,In_4,In_36);
nand U91 (N_91,In_298,In_718);
or U92 (N_92,In_499,In_90);
nand U93 (N_93,In_714,In_535);
and U94 (N_94,In_283,In_112);
nor U95 (N_95,In_239,In_397);
nand U96 (N_96,In_455,In_178);
or U97 (N_97,In_247,In_301);
and U98 (N_98,In_312,In_206);
nand U99 (N_99,In_739,In_349);
xor U100 (N_100,N_11,In_386);
xnor U101 (N_101,In_605,In_192);
nor U102 (N_102,In_742,In_101);
nor U103 (N_103,In_86,In_749);
and U104 (N_104,In_299,In_613);
or U105 (N_105,N_80,In_122);
or U106 (N_106,In_124,In_385);
and U107 (N_107,In_216,In_140);
nand U108 (N_108,In_496,In_346);
and U109 (N_109,In_698,N_18);
xor U110 (N_110,In_690,N_4);
and U111 (N_111,N_93,In_590);
nand U112 (N_112,In_609,In_661);
nand U113 (N_113,In_381,N_36);
nand U114 (N_114,In_49,In_659);
nand U115 (N_115,N_19,In_515);
nand U116 (N_116,In_166,In_631);
or U117 (N_117,In_134,In_531);
nand U118 (N_118,In_480,In_527);
or U119 (N_119,In_696,In_300);
or U120 (N_120,In_325,In_421);
nand U121 (N_121,In_238,In_82);
or U122 (N_122,In_662,In_599);
nand U123 (N_123,In_411,In_56);
and U124 (N_124,N_45,N_2);
and U125 (N_125,In_53,In_269);
or U126 (N_126,In_491,In_534);
or U127 (N_127,In_632,In_139);
and U128 (N_128,In_133,In_15);
and U129 (N_129,In_387,In_373);
nor U130 (N_130,In_565,In_451);
or U131 (N_131,In_478,In_9);
and U132 (N_132,N_44,In_619);
or U133 (N_133,In_170,In_740);
xor U134 (N_134,In_568,In_604);
nand U135 (N_135,In_399,In_363);
nand U136 (N_136,N_92,In_585);
or U137 (N_137,In_741,In_517);
or U138 (N_138,In_559,N_24);
xor U139 (N_139,In_303,In_694);
and U140 (N_140,In_458,In_621);
or U141 (N_141,In_723,In_727);
or U142 (N_142,In_433,In_691);
or U143 (N_143,In_352,In_508);
and U144 (N_144,In_215,In_160);
nand U145 (N_145,N_6,In_366);
nand U146 (N_146,In_282,In_502);
nor U147 (N_147,In_407,In_197);
nor U148 (N_148,In_380,N_28);
nand U149 (N_149,N_89,In_717);
and U150 (N_150,In_81,In_284);
nand U151 (N_151,In_697,In_382);
and U152 (N_152,In_681,N_21);
nor U153 (N_153,In_246,In_204);
or U154 (N_154,In_582,N_87);
nor U155 (N_155,In_390,In_406);
or U156 (N_156,In_67,In_367);
and U157 (N_157,In_107,N_40);
and U158 (N_158,In_362,In_509);
and U159 (N_159,N_26,N_23);
nor U160 (N_160,In_324,N_34);
or U161 (N_161,In_87,In_700);
nand U162 (N_162,In_119,In_673);
and U163 (N_163,In_544,In_172);
nor U164 (N_164,In_38,In_448);
nor U165 (N_165,In_743,In_233);
or U166 (N_166,In_34,In_279);
or U167 (N_167,N_16,In_396);
nand U168 (N_168,In_275,In_550);
and U169 (N_169,In_511,In_633);
or U170 (N_170,In_654,N_47);
nand U171 (N_171,In_184,In_257);
and U172 (N_172,In_642,In_419);
xor U173 (N_173,In_100,In_477);
nor U174 (N_174,In_398,In_434);
or U175 (N_175,In_195,In_431);
nor U176 (N_176,In_80,In_187);
nand U177 (N_177,N_5,In_721);
or U178 (N_178,In_506,In_735);
nand U179 (N_179,In_70,In_493);
or U180 (N_180,N_1,In_649);
nand U181 (N_181,In_144,In_191);
and U182 (N_182,In_40,N_96);
nand U183 (N_183,In_648,In_148);
nor U184 (N_184,In_193,In_188);
and U185 (N_185,In_8,N_65);
nor U186 (N_186,N_25,In_549);
or U187 (N_187,In_504,In_337);
nor U188 (N_188,In_401,In_731);
nor U189 (N_189,N_62,In_646);
xnor U190 (N_190,In_185,N_69);
and U191 (N_191,In_672,In_692);
or U192 (N_192,In_645,In_43);
and U193 (N_193,In_445,In_171);
nor U194 (N_194,In_520,In_618);
or U195 (N_195,N_56,In_274);
and U196 (N_196,In_468,In_248);
and U197 (N_197,N_76,In_581);
xor U198 (N_198,In_485,In_309);
nand U199 (N_199,In_30,In_183);
and U200 (N_200,In_223,N_46);
or U201 (N_201,In_157,N_104);
and U202 (N_202,N_118,In_552);
xnor U203 (N_203,N_188,N_165);
nand U204 (N_204,In_138,In_682);
nor U205 (N_205,In_227,N_112);
nand U206 (N_206,N_99,In_76);
and U207 (N_207,N_116,In_292);
or U208 (N_208,In_25,N_161);
or U209 (N_209,In_593,In_135);
nand U210 (N_210,In_623,N_134);
nand U211 (N_211,N_168,In_424);
xnor U212 (N_212,In_653,N_191);
nand U213 (N_213,In_587,In_571);
nand U214 (N_214,In_444,In_261);
and U215 (N_215,In_462,In_114);
and U216 (N_216,In_240,N_111);
and U217 (N_217,In_168,In_711);
or U218 (N_218,In_569,In_450);
nand U219 (N_219,N_73,N_181);
nor U220 (N_220,N_84,In_327);
nor U221 (N_221,N_180,In_689);
and U222 (N_222,In_592,N_148);
and U223 (N_223,In_494,In_440);
and U224 (N_224,In_542,In_469);
xnor U225 (N_225,In_276,In_566);
nand U226 (N_226,In_75,In_259);
nor U227 (N_227,N_50,In_85);
or U228 (N_228,In_173,In_720);
nand U229 (N_229,In_687,In_416);
xnor U230 (N_230,In_158,In_79);
nand U231 (N_231,In_738,N_121);
nand U232 (N_232,In_18,In_482);
xor U233 (N_233,In_486,In_570);
or U234 (N_234,In_601,N_157);
or U235 (N_235,In_131,N_90);
xnor U236 (N_236,In_437,In_145);
or U237 (N_237,In_650,In_252);
and U238 (N_238,In_245,N_88);
or U239 (N_239,N_189,In_467);
and U240 (N_240,In_235,In_355);
and U241 (N_241,In_516,In_219);
or U242 (N_242,In_208,N_77);
nor U243 (N_243,N_137,In_457);
and U244 (N_244,In_249,In_562);
or U245 (N_245,In_530,In_330);
nor U246 (N_246,In_512,In_639);
or U247 (N_247,In_539,In_522);
or U248 (N_248,N_193,N_178);
and U249 (N_249,In_224,In_479);
or U250 (N_250,N_37,In_418);
nand U251 (N_251,In_161,In_589);
or U252 (N_252,N_182,In_626);
nand U253 (N_253,In_617,In_94);
or U254 (N_254,N_61,In_492);
nand U255 (N_255,In_410,In_146);
and U256 (N_256,N_163,In_150);
or U257 (N_257,In_375,In_629);
or U258 (N_258,In_688,N_156);
xnor U259 (N_259,N_185,In_99);
xor U260 (N_260,In_326,In_652);
nor U261 (N_261,N_67,N_81);
nor U262 (N_262,In_294,In_130);
nor U263 (N_263,In_495,In_446);
xor U264 (N_264,N_43,In_63);
or U265 (N_265,N_125,In_556);
nor U266 (N_266,In_533,In_526);
xor U267 (N_267,N_141,In_706);
and U268 (N_268,N_195,In_497);
or U269 (N_269,N_198,N_98);
xor U270 (N_270,In_108,In_58);
xor U271 (N_271,N_33,In_655);
or U272 (N_272,N_159,In_616);
or U273 (N_273,N_41,N_68);
or U274 (N_274,In_578,In_402);
and U275 (N_275,N_58,In_60);
xnor U276 (N_276,In_289,In_608);
and U277 (N_277,In_167,In_474);
or U278 (N_278,N_133,In_428);
nand U279 (N_279,In_280,N_97);
or U280 (N_280,In_318,In_84);
or U281 (N_281,In_408,In_452);
nand U282 (N_282,In_121,In_625);
nor U283 (N_283,In_425,N_196);
nand U284 (N_284,In_666,In_600);
nor U285 (N_285,In_156,In_676);
nand U286 (N_286,N_55,In_722);
or U287 (N_287,In_262,In_234);
nor U288 (N_288,In_315,In_22);
nand U289 (N_289,In_23,In_177);
or U290 (N_290,N_75,In_11);
xor U291 (N_291,In_404,In_336);
nand U292 (N_292,In_357,In_524);
xnor U293 (N_293,In_189,In_360);
and U294 (N_294,In_417,In_155);
nand U295 (N_295,In_41,In_677);
nor U296 (N_296,In_409,In_217);
xor U297 (N_297,In_647,In_536);
and U298 (N_298,In_586,N_110);
nand U299 (N_299,In_391,N_155);
xnor U300 (N_300,N_177,In_703);
xnor U301 (N_301,In_142,In_436);
xor U302 (N_302,In_712,In_523);
nand U303 (N_303,N_227,In_199);
or U304 (N_304,In_484,In_710);
or U305 (N_305,N_114,In_684);
or U306 (N_306,In_218,N_240);
nand U307 (N_307,In_579,N_49);
or U308 (N_308,In_481,N_285);
nand U309 (N_309,In_614,In_384);
and U310 (N_310,N_59,In_3);
and U311 (N_311,In_476,In_266);
and U312 (N_312,In_635,N_63);
and U313 (N_313,In_388,In_229);
or U314 (N_314,In_636,N_292);
nor U315 (N_315,N_239,In_110);
nand U316 (N_316,In_490,In_88);
nand U317 (N_317,In_728,In_389);
or U318 (N_318,N_48,N_0);
and U319 (N_319,N_128,In_514);
and U320 (N_320,In_174,In_32);
nor U321 (N_321,In_264,In_394);
or U322 (N_322,In_175,N_70);
and U323 (N_323,In_612,N_179);
or U324 (N_324,N_247,N_275);
nor U325 (N_325,In_344,In_136);
nand U326 (N_326,In_305,N_205);
nand U327 (N_327,In_118,In_439);
xor U328 (N_328,In_699,N_297);
or U329 (N_329,In_359,N_144);
nor U330 (N_330,N_140,In_339);
or U331 (N_331,N_214,In_611);
or U332 (N_332,N_153,N_254);
nand U333 (N_333,In_66,N_271);
xnor U334 (N_334,In_724,In_422);
and U335 (N_335,In_125,N_30);
nand U336 (N_336,N_197,In_21);
nor U337 (N_337,In_369,In_39);
xnor U338 (N_338,In_510,In_306);
nor U339 (N_339,In_202,N_79);
nand U340 (N_340,In_441,In_338);
and U341 (N_341,N_31,N_129);
nand U342 (N_342,In_165,In_637);
nand U343 (N_343,In_665,N_252);
and U344 (N_344,N_123,In_236);
nor U345 (N_345,N_64,In_255);
or U346 (N_346,In_320,N_22);
xor U347 (N_347,In_345,N_105);
and U348 (N_348,In_263,In_241);
nand U349 (N_349,N_219,In_732);
or U350 (N_350,In_55,N_250);
nand U351 (N_351,N_35,In_498);
or U352 (N_352,In_702,In_210);
nor U353 (N_353,In_726,In_638);
xnor U354 (N_354,In_220,In_1);
or U355 (N_355,In_72,In_117);
or U356 (N_356,In_209,In_250);
and U357 (N_357,In_602,N_127);
or U358 (N_358,In_413,In_678);
or U359 (N_359,In_664,In_465);
and U360 (N_360,N_138,N_139);
and U361 (N_361,In_736,In_78);
nand U362 (N_362,N_283,In_335);
and U363 (N_363,In_105,N_101);
or U364 (N_364,N_42,N_203);
nand U365 (N_365,N_208,N_117);
nor U366 (N_366,In_153,In_48);
nor U367 (N_367,In_634,N_233);
nor U368 (N_368,In_304,In_683);
or U369 (N_369,N_299,In_374);
nand U370 (N_370,N_268,In_141);
nand U371 (N_371,N_207,N_251);
nand U372 (N_372,N_145,N_7);
or U373 (N_373,N_290,In_378);
nor U374 (N_374,N_199,In_713);
or U375 (N_375,In_83,N_217);
nand U376 (N_376,N_162,In_658);
nor U377 (N_377,N_126,N_10);
and U378 (N_378,In_332,In_651);
xor U379 (N_379,N_225,In_287);
nand U380 (N_380,In_126,N_12);
nor U381 (N_381,N_170,In_370);
nor U382 (N_382,N_85,N_284);
nor U383 (N_383,N_289,N_32);
and U384 (N_384,In_143,In_237);
xnor U385 (N_385,N_131,N_94);
nor U386 (N_386,N_288,In_281);
and U387 (N_387,N_206,N_210);
nand U388 (N_388,In_519,N_192);
or U389 (N_389,N_160,N_201);
and U390 (N_390,N_54,In_529);
nand U391 (N_391,N_270,N_27);
nor U392 (N_392,In_588,In_383);
nor U393 (N_393,N_119,In_716);
or U394 (N_394,N_102,In_152);
nor U395 (N_395,In_575,In_393);
or U396 (N_396,N_187,N_20);
and U397 (N_397,N_78,In_442);
nand U398 (N_398,In_507,N_216);
xnor U399 (N_399,N_71,In_33);
or U400 (N_400,In_151,In_733);
nor U401 (N_401,In_427,N_74);
and U402 (N_402,N_388,N_362);
and U403 (N_403,In_354,In_13);
nand U404 (N_404,In_2,In_470);
and U405 (N_405,In_123,N_228);
or U406 (N_406,N_147,N_261);
nor U407 (N_407,N_374,N_135);
xor U408 (N_408,N_150,N_301);
nor U409 (N_409,In_314,In_459);
nand U410 (N_410,N_399,N_113);
nand U411 (N_411,N_255,N_108);
nor U412 (N_412,N_130,N_296);
xor U413 (N_413,N_396,In_580);
nand U414 (N_414,In_503,N_330);
nor U415 (N_415,N_324,N_258);
and U416 (N_416,N_354,In_356);
nand U417 (N_417,In_368,N_238);
and U418 (N_418,N_259,N_107);
or U419 (N_419,N_83,N_332);
xnor U420 (N_420,In_670,N_293);
nor U421 (N_421,N_277,N_204);
xnor U422 (N_422,N_236,N_222);
or U423 (N_423,N_124,N_343);
nand U424 (N_424,N_387,N_224);
nor U425 (N_425,N_174,In_270);
nand U426 (N_426,In_487,In_228);
nor U427 (N_427,In_420,N_245);
or U428 (N_428,In_104,In_322);
nand U429 (N_429,N_257,N_278);
xnor U430 (N_430,N_360,In_543);
nand U431 (N_431,N_392,N_152);
or U432 (N_432,N_281,N_350);
nand U433 (N_433,In_725,N_158);
nor U434 (N_434,In_461,In_577);
or U435 (N_435,N_363,N_262);
nand U436 (N_436,N_218,N_395);
and U437 (N_437,In_295,In_557);
nor U438 (N_438,N_307,N_349);
or U439 (N_439,N_132,N_246);
nor U440 (N_440,N_352,In_97);
nor U441 (N_441,N_232,In_103);
nor U442 (N_442,N_241,In_598);
nand U443 (N_443,In_463,In_392);
or U444 (N_444,In_473,N_368);
nor U445 (N_445,N_287,N_231);
and U446 (N_446,In_190,N_220);
nand U447 (N_447,N_235,In_679);
nand U448 (N_448,In_297,In_551);
nand U449 (N_449,N_172,N_154);
or U450 (N_450,N_305,N_353);
nor U451 (N_451,In_615,N_376);
nand U452 (N_452,In_89,N_369);
nand U453 (N_453,N_164,N_213);
and U454 (N_454,N_242,N_311);
and U455 (N_455,In_656,N_82);
nor U456 (N_456,In_256,N_272);
nand U457 (N_457,N_381,N_398);
nand U458 (N_458,N_314,In_353);
nand U459 (N_459,N_319,N_356);
nand U460 (N_460,N_279,N_310);
or U461 (N_461,N_302,N_115);
and U462 (N_462,N_66,N_345);
and U463 (N_463,N_209,N_234);
nand U464 (N_464,N_91,N_375);
xnor U465 (N_465,N_339,N_327);
nand U466 (N_466,In_719,In_207);
and U467 (N_467,In_379,In_680);
or U468 (N_468,In_454,In_453);
nor U469 (N_469,In_371,In_73);
or U470 (N_470,N_265,N_304);
xor U471 (N_471,In_748,N_318);
or U472 (N_472,In_573,N_184);
nand U473 (N_473,N_72,In_179);
nand U474 (N_474,N_171,In_583);
and U475 (N_475,N_280,N_136);
or U476 (N_476,N_176,N_323);
and U477 (N_477,N_29,N_122);
nand U478 (N_478,N_229,N_291);
nor U479 (N_479,N_249,N_378);
nand U480 (N_480,N_276,N_267);
nor U481 (N_481,N_322,N_230);
or U482 (N_482,N_370,In_709);
or U483 (N_483,In_260,N_100);
nor U484 (N_484,N_169,In_715);
nor U485 (N_485,N_321,In_640);
nand U486 (N_486,In_705,In_341);
xor U487 (N_487,N_274,N_194);
nor U488 (N_488,N_340,N_282);
nor U489 (N_489,In_59,N_103);
xor U490 (N_490,N_202,N_364);
nor U491 (N_491,N_151,In_271);
nor U492 (N_492,In_746,N_357);
and U493 (N_493,N_337,N_260);
nor U494 (N_494,In_7,N_8);
or U495 (N_495,In_546,N_14);
and U496 (N_496,N_221,N_333);
or U497 (N_497,In_74,N_317);
nand U498 (N_498,N_38,N_226);
nor U499 (N_499,N_39,In_414);
and U500 (N_500,N_86,In_0);
nand U501 (N_501,In_222,N_380);
and U502 (N_502,N_361,N_498);
xor U503 (N_503,N_390,N_467);
and U504 (N_504,N_313,N_372);
and U505 (N_505,N_477,N_57);
and U506 (N_506,N_473,N_386);
nor U507 (N_507,N_384,In_149);
or U508 (N_508,In_671,N_294);
nor U509 (N_509,N_433,N_53);
xnor U510 (N_510,N_425,N_303);
or U511 (N_511,N_413,N_435);
and U512 (N_512,In_64,N_461);
and U513 (N_513,In_564,N_52);
or U514 (N_514,In_323,In_328);
xor U515 (N_515,N_458,N_373);
and U516 (N_516,N_456,N_454);
xor U517 (N_517,In_50,N_253);
and U518 (N_518,N_149,N_465);
nor U519 (N_519,N_397,N_328);
or U520 (N_520,N_17,N_410);
and U521 (N_521,N_186,N_400);
or U522 (N_522,In_31,N_462);
nor U523 (N_523,N_423,In_28);
and U524 (N_524,N_223,N_15);
nand U525 (N_525,N_446,N_351);
nand U526 (N_526,N_211,N_403);
or U527 (N_527,N_478,N_436);
nand U528 (N_528,N_326,N_445);
and U529 (N_529,N_334,N_371);
xor U530 (N_530,N_382,In_471);
or U531 (N_531,In_628,N_348);
or U532 (N_532,N_331,In_92);
and U533 (N_533,N_309,N_359);
nor U534 (N_534,N_9,In_44);
nand U535 (N_535,N_295,N_60);
nor U536 (N_536,N_488,N_109);
nor U537 (N_537,N_167,N_441);
or U538 (N_538,In_272,In_267);
nand U539 (N_539,N_393,N_447);
nand U540 (N_540,In_200,N_476);
xnor U541 (N_541,N_451,N_444);
nand U542 (N_542,N_355,N_450);
or U543 (N_543,In_730,N_449);
nor U544 (N_544,N_341,N_406);
nand U545 (N_545,N_312,N_448);
and U546 (N_546,N_237,In_102);
or U547 (N_547,N_298,N_407);
and U548 (N_548,N_190,N_489);
nor U549 (N_549,N_379,N_365);
nor U550 (N_550,N_437,N_338);
and U551 (N_551,In_597,N_439);
and U552 (N_552,N_346,N_325);
nand U553 (N_553,N_412,N_469);
and U554 (N_554,N_420,N_175);
nand U555 (N_555,N_463,In_54);
nor U556 (N_556,N_389,N_409);
xnor U557 (N_557,In_669,In_400);
nor U558 (N_558,N_453,N_429);
and U559 (N_559,N_430,N_142);
nor U560 (N_560,N_248,N_411);
or U561 (N_561,N_417,In_98);
xnor U562 (N_562,N_344,N_434);
nand U563 (N_563,N_306,N_497);
and U564 (N_564,N_95,N_336);
nand U565 (N_565,N_394,N_13);
and U566 (N_566,In_545,N_472);
or U567 (N_567,In_113,In_96);
or U568 (N_568,N_269,In_443);
nor U569 (N_569,N_401,N_315);
nor U570 (N_570,N_263,N_487);
nor U571 (N_571,In_10,N_329);
and U572 (N_572,N_166,In_342);
nor U573 (N_573,N_431,In_16);
nor U574 (N_574,N_424,N_418);
nor U575 (N_575,In_350,N_215);
nor U576 (N_576,N_377,N_416);
nor U577 (N_577,N_256,N_466);
nor U578 (N_578,N_474,N_422);
nand U579 (N_579,N_273,N_316);
nand U580 (N_580,N_402,In_657);
nor U581 (N_581,N_358,N_494);
nand U582 (N_582,N_408,N_481);
nor U583 (N_583,In_20,N_146);
nor U584 (N_584,N_342,N_264);
xor U585 (N_585,N_440,N_496);
and U586 (N_586,N_493,In_334);
nand U587 (N_587,N_475,N_470);
nor U588 (N_588,N_106,In_630);
or U589 (N_589,N_212,N_490);
nand U590 (N_590,N_391,N_486);
and U591 (N_591,N_455,N_3);
and U592 (N_592,N_385,N_452);
nand U593 (N_593,N_404,N_438);
nor U594 (N_594,N_482,N_143);
nand U595 (N_595,N_120,N_442);
and U596 (N_596,N_183,In_181);
nor U597 (N_597,In_685,In_194);
nand U598 (N_598,N_414,N_173);
or U599 (N_599,N_320,N_308);
nor U600 (N_600,N_580,N_432);
xnor U601 (N_601,N_512,N_554);
nand U602 (N_602,In_361,N_579);
and U603 (N_603,N_566,N_525);
nand U604 (N_604,N_541,N_563);
nand U605 (N_605,N_51,N_243);
nor U606 (N_606,N_593,N_300);
or U607 (N_607,N_562,N_558);
or U608 (N_608,N_514,N_528);
or U609 (N_609,In_412,N_539);
and U610 (N_610,N_532,N_383);
nor U611 (N_611,N_200,N_492);
or U612 (N_612,N_546,N_495);
and U613 (N_613,N_500,N_535);
xor U614 (N_614,N_484,N_536);
nand U615 (N_615,In_69,N_459);
and U616 (N_616,N_586,N_427);
and U617 (N_617,N_499,In_622);
nand U618 (N_618,N_457,N_560);
or U619 (N_619,N_524,N_244);
or U620 (N_620,N_286,N_585);
or U621 (N_621,N_502,N_533);
nand U622 (N_622,N_567,N_483);
nand U623 (N_623,N_491,N_556);
or U624 (N_624,N_531,In_466);
nand U625 (N_625,N_573,N_506);
or U626 (N_626,N_509,N_594);
or U627 (N_627,N_589,N_367);
nand U628 (N_628,N_568,N_479);
or U629 (N_629,N_564,N_571);
nor U630 (N_630,In_47,N_523);
and U631 (N_631,N_591,N_542);
nor U632 (N_632,N_520,N_511);
nor U633 (N_633,N_553,N_572);
and U634 (N_634,N_428,N_574);
and U635 (N_635,N_508,In_308);
nand U636 (N_636,N_501,In_554);
and U637 (N_637,N_569,N_522);
nor U638 (N_638,N_521,N_597);
xor U639 (N_639,N_405,N_415);
nand U640 (N_640,N_565,N_587);
nand U641 (N_641,N_519,N_530);
and U642 (N_642,N_538,N_460);
or U643 (N_643,N_480,N_583);
and U644 (N_644,N_598,N_504);
or U645 (N_645,N_578,N_550);
nor U646 (N_646,N_549,N_576);
nand U647 (N_647,N_559,In_221);
nand U648 (N_648,N_545,N_347);
nand U649 (N_649,N_515,N_529);
and U650 (N_650,N_582,N_419);
and U651 (N_651,N_468,N_507);
nand U652 (N_652,N_534,N_526);
nor U653 (N_653,In_555,N_443);
or U654 (N_654,N_505,N_518);
xor U655 (N_655,N_584,N_266);
xnor U656 (N_656,N_517,N_577);
nor U657 (N_657,N_548,N_588);
or U658 (N_658,N_599,In_426);
or U659 (N_659,N_421,N_547);
nor U660 (N_660,N_552,N_366);
nand U661 (N_661,N_516,N_596);
xor U662 (N_662,N_551,N_471);
nand U663 (N_663,N_426,N_513);
or U664 (N_664,N_544,N_581);
nor U665 (N_665,N_575,N_543);
or U666 (N_666,N_595,N_561);
or U667 (N_667,N_590,In_14);
nand U668 (N_668,N_510,N_555);
nor U669 (N_669,N_503,In_518);
and U670 (N_670,In_708,N_592);
and U671 (N_671,N_335,N_570);
nand U672 (N_672,N_557,N_527);
nor U673 (N_673,N_537,N_485);
nor U674 (N_674,N_464,N_540);
nand U675 (N_675,N_564,In_221);
nand U676 (N_676,N_508,N_415);
and U677 (N_677,N_566,N_503);
and U678 (N_678,N_538,N_527);
and U679 (N_679,N_518,N_300);
nand U680 (N_680,N_556,N_534);
or U681 (N_681,N_570,N_536);
nor U682 (N_682,N_243,N_585);
xor U683 (N_683,N_535,N_521);
and U684 (N_684,N_266,N_366);
nor U685 (N_685,N_464,N_500);
or U686 (N_686,N_560,N_505);
and U687 (N_687,N_529,In_14);
or U688 (N_688,N_51,N_556);
or U689 (N_689,N_554,In_555);
nor U690 (N_690,N_574,N_565);
nand U691 (N_691,N_589,N_575);
or U692 (N_692,In_308,N_558);
xnor U693 (N_693,N_502,N_510);
and U694 (N_694,N_578,N_243);
nor U695 (N_695,N_588,N_566);
nor U696 (N_696,In_14,N_483);
and U697 (N_697,N_501,N_506);
nand U698 (N_698,N_515,N_574);
or U699 (N_699,N_534,In_412);
and U700 (N_700,N_688,N_677);
or U701 (N_701,N_624,N_662);
xor U702 (N_702,N_630,N_607);
nand U703 (N_703,N_683,N_673);
nor U704 (N_704,N_645,N_664);
and U705 (N_705,N_682,N_656);
and U706 (N_706,N_665,N_609);
or U707 (N_707,N_696,N_612);
nand U708 (N_708,N_657,N_684);
or U709 (N_709,N_618,N_666);
xnor U710 (N_710,N_629,N_641);
nand U711 (N_711,N_614,N_636);
or U712 (N_712,N_642,N_690);
or U713 (N_713,N_628,N_679);
and U714 (N_714,N_632,N_610);
nand U715 (N_715,N_623,N_654);
xnor U716 (N_716,N_675,N_667);
xor U717 (N_717,N_613,N_695);
and U718 (N_718,N_699,N_697);
and U719 (N_719,N_603,N_652);
nand U720 (N_720,N_620,N_601);
nand U721 (N_721,N_626,N_680);
xor U722 (N_722,N_663,N_681);
or U723 (N_723,N_634,N_655);
nor U724 (N_724,N_648,N_692);
or U725 (N_725,N_693,N_658);
nand U726 (N_726,N_640,N_659);
nand U727 (N_727,N_605,N_644);
nor U728 (N_728,N_691,N_611);
nor U729 (N_729,N_686,N_674);
xor U730 (N_730,N_635,N_622);
and U731 (N_731,N_694,N_606);
or U732 (N_732,N_685,N_638);
nor U733 (N_733,N_676,N_647);
nor U734 (N_734,N_671,N_669);
nor U735 (N_735,N_650,N_678);
nand U736 (N_736,N_619,N_689);
nand U737 (N_737,N_672,N_651);
nand U738 (N_738,N_646,N_698);
and U739 (N_739,N_608,N_602);
nand U740 (N_740,N_625,N_615);
or U741 (N_741,N_600,N_660);
nand U742 (N_742,N_639,N_649);
or U743 (N_743,N_643,N_670);
nor U744 (N_744,N_653,N_627);
and U745 (N_745,N_616,N_631);
or U746 (N_746,N_668,N_604);
and U747 (N_747,N_661,N_621);
and U748 (N_748,N_617,N_687);
and U749 (N_749,N_633,N_637);
or U750 (N_750,N_655,N_636);
nand U751 (N_751,N_670,N_609);
nand U752 (N_752,N_604,N_633);
and U753 (N_753,N_687,N_606);
and U754 (N_754,N_623,N_666);
or U755 (N_755,N_630,N_601);
or U756 (N_756,N_683,N_625);
nor U757 (N_757,N_681,N_642);
nor U758 (N_758,N_649,N_673);
nor U759 (N_759,N_693,N_646);
and U760 (N_760,N_682,N_690);
nand U761 (N_761,N_681,N_643);
and U762 (N_762,N_661,N_619);
nor U763 (N_763,N_689,N_632);
nor U764 (N_764,N_699,N_640);
nor U765 (N_765,N_686,N_662);
or U766 (N_766,N_663,N_656);
xor U767 (N_767,N_661,N_604);
nand U768 (N_768,N_605,N_604);
nor U769 (N_769,N_619,N_681);
nand U770 (N_770,N_624,N_668);
or U771 (N_771,N_607,N_654);
nor U772 (N_772,N_627,N_667);
xor U773 (N_773,N_618,N_604);
and U774 (N_774,N_693,N_630);
nand U775 (N_775,N_680,N_640);
nor U776 (N_776,N_627,N_675);
nand U777 (N_777,N_698,N_651);
and U778 (N_778,N_678,N_612);
nand U779 (N_779,N_650,N_648);
nor U780 (N_780,N_619,N_633);
nor U781 (N_781,N_617,N_650);
or U782 (N_782,N_667,N_616);
or U783 (N_783,N_682,N_674);
and U784 (N_784,N_679,N_634);
nand U785 (N_785,N_665,N_620);
or U786 (N_786,N_644,N_673);
and U787 (N_787,N_676,N_636);
and U788 (N_788,N_659,N_633);
nand U789 (N_789,N_671,N_613);
nand U790 (N_790,N_663,N_686);
nor U791 (N_791,N_654,N_651);
and U792 (N_792,N_617,N_626);
nand U793 (N_793,N_612,N_617);
xor U794 (N_794,N_614,N_638);
nor U795 (N_795,N_615,N_606);
nand U796 (N_796,N_690,N_606);
xnor U797 (N_797,N_603,N_666);
and U798 (N_798,N_670,N_682);
nor U799 (N_799,N_643,N_646);
nor U800 (N_800,N_707,N_762);
or U801 (N_801,N_774,N_755);
nor U802 (N_802,N_797,N_757);
nor U803 (N_803,N_734,N_717);
xor U804 (N_804,N_701,N_739);
or U805 (N_805,N_783,N_706);
nand U806 (N_806,N_791,N_733);
nor U807 (N_807,N_720,N_788);
nand U808 (N_808,N_776,N_723);
nor U809 (N_809,N_721,N_725);
nand U810 (N_810,N_715,N_708);
nand U811 (N_811,N_786,N_789);
xor U812 (N_812,N_718,N_724);
or U813 (N_813,N_747,N_740);
nor U814 (N_814,N_738,N_756);
nor U815 (N_815,N_749,N_761);
nand U816 (N_816,N_711,N_770);
xor U817 (N_817,N_704,N_730);
or U818 (N_818,N_779,N_778);
or U819 (N_819,N_767,N_742);
nand U820 (N_820,N_784,N_799);
nand U821 (N_821,N_790,N_782);
nor U822 (N_822,N_785,N_766);
nor U823 (N_823,N_780,N_713);
nor U824 (N_824,N_792,N_743);
nand U825 (N_825,N_748,N_735);
or U826 (N_826,N_798,N_753);
or U827 (N_827,N_781,N_710);
or U828 (N_828,N_777,N_719);
or U829 (N_829,N_794,N_746);
xnor U830 (N_830,N_727,N_793);
and U831 (N_831,N_744,N_714);
nor U832 (N_832,N_773,N_750);
or U833 (N_833,N_703,N_754);
nor U834 (N_834,N_722,N_771);
nand U835 (N_835,N_795,N_705);
nor U836 (N_836,N_741,N_731);
and U837 (N_837,N_728,N_752);
nand U838 (N_838,N_769,N_732);
or U839 (N_839,N_764,N_765);
nor U840 (N_840,N_737,N_775);
nand U841 (N_841,N_736,N_787);
and U842 (N_842,N_763,N_758);
and U843 (N_843,N_712,N_745);
nor U844 (N_844,N_768,N_716);
nand U845 (N_845,N_751,N_702);
and U846 (N_846,N_772,N_759);
xnor U847 (N_847,N_700,N_729);
or U848 (N_848,N_726,N_709);
and U849 (N_849,N_796,N_760);
or U850 (N_850,N_784,N_706);
nor U851 (N_851,N_723,N_748);
nand U852 (N_852,N_709,N_778);
nand U853 (N_853,N_786,N_728);
nor U854 (N_854,N_774,N_797);
and U855 (N_855,N_798,N_795);
nand U856 (N_856,N_755,N_710);
xor U857 (N_857,N_737,N_795);
and U858 (N_858,N_782,N_705);
or U859 (N_859,N_780,N_736);
nor U860 (N_860,N_720,N_708);
nand U861 (N_861,N_777,N_701);
or U862 (N_862,N_733,N_732);
and U863 (N_863,N_705,N_725);
xnor U864 (N_864,N_717,N_790);
nor U865 (N_865,N_764,N_751);
nand U866 (N_866,N_779,N_755);
xnor U867 (N_867,N_731,N_734);
nand U868 (N_868,N_762,N_738);
xor U869 (N_869,N_769,N_782);
and U870 (N_870,N_719,N_766);
and U871 (N_871,N_758,N_707);
or U872 (N_872,N_704,N_725);
and U873 (N_873,N_758,N_752);
and U874 (N_874,N_765,N_771);
or U875 (N_875,N_730,N_707);
nor U876 (N_876,N_751,N_711);
xor U877 (N_877,N_736,N_722);
and U878 (N_878,N_720,N_791);
or U879 (N_879,N_776,N_712);
nand U880 (N_880,N_732,N_737);
xnor U881 (N_881,N_713,N_791);
and U882 (N_882,N_729,N_740);
nor U883 (N_883,N_754,N_738);
nand U884 (N_884,N_745,N_785);
and U885 (N_885,N_771,N_745);
and U886 (N_886,N_783,N_747);
or U887 (N_887,N_706,N_760);
nor U888 (N_888,N_701,N_718);
nor U889 (N_889,N_782,N_748);
and U890 (N_890,N_709,N_773);
nand U891 (N_891,N_751,N_710);
nand U892 (N_892,N_777,N_769);
nor U893 (N_893,N_740,N_722);
nor U894 (N_894,N_707,N_712);
and U895 (N_895,N_769,N_774);
nor U896 (N_896,N_734,N_783);
and U897 (N_897,N_728,N_713);
or U898 (N_898,N_741,N_720);
and U899 (N_899,N_764,N_722);
or U900 (N_900,N_828,N_891);
nand U901 (N_901,N_859,N_880);
and U902 (N_902,N_840,N_847);
and U903 (N_903,N_823,N_831);
nor U904 (N_904,N_821,N_845);
xnor U905 (N_905,N_895,N_843);
xnor U906 (N_906,N_844,N_829);
and U907 (N_907,N_869,N_856);
nand U908 (N_908,N_872,N_833);
xor U909 (N_909,N_813,N_808);
nand U910 (N_910,N_883,N_852);
nand U911 (N_911,N_816,N_851);
nand U912 (N_912,N_855,N_815);
xnor U913 (N_913,N_874,N_882);
or U914 (N_914,N_841,N_826);
or U915 (N_915,N_835,N_825);
and U916 (N_916,N_810,N_819);
xor U917 (N_917,N_827,N_893);
nor U918 (N_918,N_857,N_839);
nor U919 (N_919,N_824,N_807);
and U920 (N_920,N_850,N_802);
nor U921 (N_921,N_848,N_865);
or U922 (N_922,N_854,N_811);
or U923 (N_923,N_862,N_800);
xor U924 (N_924,N_846,N_876);
xnor U925 (N_925,N_894,N_887);
nand U926 (N_926,N_898,N_803);
and U927 (N_927,N_860,N_834);
xnor U928 (N_928,N_897,N_842);
nor U929 (N_929,N_866,N_884);
or U930 (N_930,N_812,N_836);
nand U931 (N_931,N_881,N_830);
and U932 (N_932,N_864,N_817);
and U933 (N_933,N_822,N_801);
nand U934 (N_934,N_877,N_896);
xnor U935 (N_935,N_832,N_885);
nor U936 (N_936,N_879,N_838);
nor U937 (N_937,N_892,N_867);
nor U938 (N_938,N_837,N_890);
nor U939 (N_939,N_868,N_818);
nand U940 (N_940,N_809,N_899);
nand U941 (N_941,N_820,N_805);
and U942 (N_942,N_878,N_853);
and U943 (N_943,N_873,N_888);
or U944 (N_944,N_814,N_875);
and U945 (N_945,N_804,N_870);
and U946 (N_946,N_863,N_849);
or U947 (N_947,N_871,N_806);
xnor U948 (N_948,N_886,N_858);
or U949 (N_949,N_861,N_889);
and U950 (N_950,N_876,N_812);
xnor U951 (N_951,N_873,N_872);
and U952 (N_952,N_849,N_874);
nor U953 (N_953,N_853,N_857);
or U954 (N_954,N_889,N_887);
nand U955 (N_955,N_899,N_868);
and U956 (N_956,N_818,N_855);
nor U957 (N_957,N_842,N_819);
xor U958 (N_958,N_808,N_821);
or U959 (N_959,N_872,N_894);
nand U960 (N_960,N_870,N_866);
nand U961 (N_961,N_826,N_846);
or U962 (N_962,N_866,N_871);
and U963 (N_963,N_828,N_869);
or U964 (N_964,N_804,N_839);
nor U965 (N_965,N_829,N_809);
or U966 (N_966,N_879,N_869);
or U967 (N_967,N_836,N_822);
and U968 (N_968,N_822,N_842);
and U969 (N_969,N_809,N_842);
or U970 (N_970,N_829,N_863);
or U971 (N_971,N_863,N_835);
xor U972 (N_972,N_870,N_897);
and U973 (N_973,N_875,N_802);
or U974 (N_974,N_821,N_863);
and U975 (N_975,N_844,N_853);
or U976 (N_976,N_851,N_841);
or U977 (N_977,N_898,N_877);
xnor U978 (N_978,N_859,N_846);
and U979 (N_979,N_866,N_877);
and U980 (N_980,N_856,N_846);
nor U981 (N_981,N_803,N_881);
xor U982 (N_982,N_899,N_833);
nand U983 (N_983,N_857,N_823);
nor U984 (N_984,N_898,N_817);
nor U985 (N_985,N_825,N_831);
or U986 (N_986,N_886,N_882);
or U987 (N_987,N_823,N_822);
and U988 (N_988,N_879,N_803);
or U989 (N_989,N_870,N_858);
nand U990 (N_990,N_860,N_862);
and U991 (N_991,N_843,N_808);
nand U992 (N_992,N_851,N_862);
nor U993 (N_993,N_800,N_839);
or U994 (N_994,N_833,N_835);
and U995 (N_995,N_827,N_833);
or U996 (N_996,N_825,N_851);
or U997 (N_997,N_824,N_845);
nand U998 (N_998,N_845,N_855);
and U999 (N_999,N_871,N_877);
and U1000 (N_1000,N_933,N_972);
or U1001 (N_1001,N_940,N_995);
nor U1002 (N_1002,N_938,N_948);
xor U1003 (N_1003,N_955,N_917);
nand U1004 (N_1004,N_983,N_946);
nor U1005 (N_1005,N_905,N_976);
nand U1006 (N_1006,N_965,N_919);
or U1007 (N_1007,N_949,N_926);
xnor U1008 (N_1008,N_984,N_992);
nor U1009 (N_1009,N_959,N_969);
nand U1010 (N_1010,N_960,N_937);
nand U1011 (N_1011,N_957,N_978);
nand U1012 (N_1012,N_925,N_975);
or U1013 (N_1013,N_939,N_915);
nand U1014 (N_1014,N_932,N_914);
or U1015 (N_1015,N_999,N_996);
nor U1016 (N_1016,N_953,N_918);
nand U1017 (N_1017,N_954,N_988);
xor U1018 (N_1018,N_942,N_991);
nor U1019 (N_1019,N_922,N_935);
and U1020 (N_1020,N_916,N_906);
nor U1021 (N_1021,N_997,N_967);
nand U1022 (N_1022,N_963,N_970);
or U1023 (N_1023,N_931,N_964);
and U1024 (N_1024,N_900,N_968);
nand U1025 (N_1025,N_961,N_980);
nand U1026 (N_1026,N_943,N_901);
nand U1027 (N_1027,N_962,N_930);
or U1028 (N_1028,N_974,N_977);
and U1029 (N_1029,N_998,N_982);
or U1030 (N_1030,N_907,N_971);
or U1031 (N_1031,N_902,N_994);
xor U1032 (N_1032,N_923,N_979);
and U1033 (N_1033,N_934,N_910);
or U1034 (N_1034,N_928,N_985);
nand U1035 (N_1035,N_956,N_936);
and U1036 (N_1036,N_913,N_989);
nand U1037 (N_1037,N_908,N_920);
nor U1038 (N_1038,N_924,N_981);
nand U1039 (N_1039,N_990,N_921);
nand U1040 (N_1040,N_941,N_958);
nand U1041 (N_1041,N_986,N_911);
and U1042 (N_1042,N_944,N_927);
nand U1043 (N_1043,N_945,N_966);
and U1044 (N_1044,N_993,N_912);
or U1045 (N_1045,N_929,N_973);
or U1046 (N_1046,N_952,N_951);
or U1047 (N_1047,N_909,N_903);
nor U1048 (N_1048,N_950,N_947);
and U1049 (N_1049,N_904,N_987);
nand U1050 (N_1050,N_973,N_927);
nand U1051 (N_1051,N_982,N_922);
nor U1052 (N_1052,N_913,N_970);
and U1053 (N_1053,N_964,N_900);
nand U1054 (N_1054,N_909,N_917);
nor U1055 (N_1055,N_944,N_995);
nor U1056 (N_1056,N_903,N_963);
nand U1057 (N_1057,N_924,N_949);
nand U1058 (N_1058,N_976,N_910);
nand U1059 (N_1059,N_963,N_905);
nor U1060 (N_1060,N_964,N_917);
or U1061 (N_1061,N_977,N_950);
and U1062 (N_1062,N_909,N_938);
or U1063 (N_1063,N_942,N_926);
or U1064 (N_1064,N_969,N_921);
or U1065 (N_1065,N_917,N_985);
or U1066 (N_1066,N_969,N_989);
and U1067 (N_1067,N_980,N_976);
and U1068 (N_1068,N_964,N_995);
nand U1069 (N_1069,N_920,N_960);
or U1070 (N_1070,N_979,N_905);
nand U1071 (N_1071,N_904,N_931);
nor U1072 (N_1072,N_935,N_957);
nand U1073 (N_1073,N_956,N_952);
or U1074 (N_1074,N_939,N_913);
nor U1075 (N_1075,N_921,N_963);
and U1076 (N_1076,N_986,N_923);
and U1077 (N_1077,N_969,N_902);
and U1078 (N_1078,N_982,N_980);
nand U1079 (N_1079,N_937,N_923);
or U1080 (N_1080,N_929,N_956);
nand U1081 (N_1081,N_914,N_968);
nand U1082 (N_1082,N_930,N_922);
and U1083 (N_1083,N_999,N_943);
nand U1084 (N_1084,N_971,N_903);
nor U1085 (N_1085,N_979,N_924);
xor U1086 (N_1086,N_999,N_927);
nor U1087 (N_1087,N_982,N_942);
nand U1088 (N_1088,N_956,N_960);
and U1089 (N_1089,N_952,N_999);
and U1090 (N_1090,N_952,N_946);
or U1091 (N_1091,N_924,N_917);
nor U1092 (N_1092,N_947,N_945);
nor U1093 (N_1093,N_906,N_988);
or U1094 (N_1094,N_959,N_976);
and U1095 (N_1095,N_939,N_918);
and U1096 (N_1096,N_911,N_984);
and U1097 (N_1097,N_990,N_984);
and U1098 (N_1098,N_903,N_933);
or U1099 (N_1099,N_938,N_956);
and U1100 (N_1100,N_1091,N_1095);
nor U1101 (N_1101,N_1056,N_1041);
nand U1102 (N_1102,N_1083,N_1063);
or U1103 (N_1103,N_1068,N_1021);
and U1104 (N_1104,N_1060,N_1017);
nor U1105 (N_1105,N_1054,N_1046);
nand U1106 (N_1106,N_1097,N_1057);
nor U1107 (N_1107,N_1045,N_1080);
and U1108 (N_1108,N_1050,N_1022);
or U1109 (N_1109,N_1025,N_1090);
nand U1110 (N_1110,N_1086,N_1006);
xor U1111 (N_1111,N_1040,N_1074);
nand U1112 (N_1112,N_1002,N_1007);
nand U1113 (N_1113,N_1015,N_1069);
xor U1114 (N_1114,N_1093,N_1055);
nor U1115 (N_1115,N_1084,N_1077);
and U1116 (N_1116,N_1053,N_1061);
or U1117 (N_1117,N_1037,N_1009);
or U1118 (N_1118,N_1010,N_1003);
and U1119 (N_1119,N_1026,N_1064);
nor U1120 (N_1120,N_1078,N_1092);
or U1121 (N_1121,N_1008,N_1071);
nand U1122 (N_1122,N_1047,N_1023);
xnor U1123 (N_1123,N_1076,N_1059);
or U1124 (N_1124,N_1024,N_1019);
xnor U1125 (N_1125,N_1081,N_1058);
nand U1126 (N_1126,N_1030,N_1096);
nand U1127 (N_1127,N_1085,N_1098);
nand U1128 (N_1128,N_1035,N_1036);
and U1129 (N_1129,N_1062,N_1070);
nor U1130 (N_1130,N_1033,N_1043);
or U1131 (N_1131,N_1032,N_1044);
and U1132 (N_1132,N_1013,N_1067);
xnor U1133 (N_1133,N_1099,N_1079);
nand U1134 (N_1134,N_1004,N_1020);
and U1135 (N_1135,N_1011,N_1016);
nand U1136 (N_1136,N_1005,N_1088);
or U1137 (N_1137,N_1031,N_1029);
nand U1138 (N_1138,N_1075,N_1018);
or U1139 (N_1139,N_1027,N_1072);
nor U1140 (N_1140,N_1089,N_1052);
nand U1141 (N_1141,N_1038,N_1001);
nor U1142 (N_1142,N_1049,N_1028);
and U1143 (N_1143,N_1034,N_1094);
and U1144 (N_1144,N_1039,N_1082);
and U1145 (N_1145,N_1087,N_1073);
nand U1146 (N_1146,N_1014,N_1065);
or U1147 (N_1147,N_1000,N_1051);
nand U1148 (N_1148,N_1042,N_1066);
and U1149 (N_1149,N_1012,N_1048);
nand U1150 (N_1150,N_1022,N_1082);
nand U1151 (N_1151,N_1098,N_1071);
nor U1152 (N_1152,N_1018,N_1036);
nand U1153 (N_1153,N_1075,N_1087);
and U1154 (N_1154,N_1022,N_1099);
nand U1155 (N_1155,N_1055,N_1044);
nand U1156 (N_1156,N_1091,N_1072);
and U1157 (N_1157,N_1082,N_1045);
xnor U1158 (N_1158,N_1057,N_1011);
or U1159 (N_1159,N_1016,N_1062);
and U1160 (N_1160,N_1035,N_1048);
nand U1161 (N_1161,N_1055,N_1048);
and U1162 (N_1162,N_1086,N_1052);
and U1163 (N_1163,N_1092,N_1013);
and U1164 (N_1164,N_1008,N_1005);
or U1165 (N_1165,N_1001,N_1011);
nor U1166 (N_1166,N_1039,N_1063);
or U1167 (N_1167,N_1084,N_1027);
xor U1168 (N_1168,N_1025,N_1091);
nand U1169 (N_1169,N_1029,N_1095);
and U1170 (N_1170,N_1047,N_1058);
or U1171 (N_1171,N_1017,N_1092);
and U1172 (N_1172,N_1068,N_1039);
and U1173 (N_1173,N_1010,N_1032);
nand U1174 (N_1174,N_1063,N_1022);
nor U1175 (N_1175,N_1041,N_1031);
and U1176 (N_1176,N_1062,N_1053);
nor U1177 (N_1177,N_1065,N_1032);
and U1178 (N_1178,N_1023,N_1016);
xor U1179 (N_1179,N_1091,N_1010);
xor U1180 (N_1180,N_1064,N_1039);
and U1181 (N_1181,N_1090,N_1023);
nor U1182 (N_1182,N_1061,N_1008);
and U1183 (N_1183,N_1041,N_1024);
or U1184 (N_1184,N_1027,N_1093);
and U1185 (N_1185,N_1080,N_1075);
and U1186 (N_1186,N_1029,N_1009);
nor U1187 (N_1187,N_1063,N_1065);
nor U1188 (N_1188,N_1004,N_1080);
nand U1189 (N_1189,N_1058,N_1011);
and U1190 (N_1190,N_1058,N_1086);
or U1191 (N_1191,N_1001,N_1095);
nor U1192 (N_1192,N_1084,N_1060);
nand U1193 (N_1193,N_1016,N_1065);
and U1194 (N_1194,N_1040,N_1054);
and U1195 (N_1195,N_1022,N_1020);
xnor U1196 (N_1196,N_1023,N_1048);
nor U1197 (N_1197,N_1016,N_1043);
and U1198 (N_1198,N_1087,N_1054);
or U1199 (N_1199,N_1096,N_1056);
and U1200 (N_1200,N_1178,N_1198);
nand U1201 (N_1201,N_1123,N_1171);
and U1202 (N_1202,N_1190,N_1135);
nand U1203 (N_1203,N_1186,N_1125);
xor U1204 (N_1204,N_1159,N_1158);
and U1205 (N_1205,N_1196,N_1129);
nor U1206 (N_1206,N_1170,N_1173);
and U1207 (N_1207,N_1197,N_1118);
or U1208 (N_1208,N_1136,N_1105);
nor U1209 (N_1209,N_1110,N_1144);
and U1210 (N_1210,N_1104,N_1127);
and U1211 (N_1211,N_1193,N_1130);
nor U1212 (N_1212,N_1179,N_1142);
and U1213 (N_1213,N_1140,N_1141);
or U1214 (N_1214,N_1148,N_1164);
or U1215 (N_1215,N_1124,N_1120);
and U1216 (N_1216,N_1181,N_1150);
nor U1217 (N_1217,N_1195,N_1114);
and U1218 (N_1218,N_1161,N_1162);
nor U1219 (N_1219,N_1132,N_1157);
nor U1220 (N_1220,N_1167,N_1126);
nand U1221 (N_1221,N_1108,N_1185);
or U1222 (N_1222,N_1189,N_1160);
nand U1223 (N_1223,N_1184,N_1191);
and U1224 (N_1224,N_1145,N_1109);
nor U1225 (N_1225,N_1122,N_1180);
nand U1226 (N_1226,N_1143,N_1176);
nand U1227 (N_1227,N_1131,N_1154);
or U1228 (N_1228,N_1168,N_1133);
nand U1229 (N_1229,N_1137,N_1172);
nor U1230 (N_1230,N_1156,N_1119);
or U1231 (N_1231,N_1187,N_1169);
nand U1232 (N_1232,N_1106,N_1117);
and U1233 (N_1233,N_1153,N_1146);
or U1234 (N_1234,N_1174,N_1166);
or U1235 (N_1235,N_1111,N_1194);
nor U1236 (N_1236,N_1183,N_1152);
xor U1237 (N_1237,N_1101,N_1192);
nand U1238 (N_1238,N_1149,N_1128);
nor U1239 (N_1239,N_1134,N_1188);
nor U1240 (N_1240,N_1116,N_1121);
or U1241 (N_1241,N_1147,N_1113);
and U1242 (N_1242,N_1155,N_1115);
or U1243 (N_1243,N_1103,N_1163);
nor U1244 (N_1244,N_1138,N_1165);
or U1245 (N_1245,N_1182,N_1175);
and U1246 (N_1246,N_1100,N_1112);
nor U1247 (N_1247,N_1102,N_1177);
and U1248 (N_1248,N_1199,N_1151);
xnor U1249 (N_1249,N_1107,N_1139);
nand U1250 (N_1250,N_1104,N_1192);
nand U1251 (N_1251,N_1124,N_1140);
or U1252 (N_1252,N_1114,N_1155);
xnor U1253 (N_1253,N_1157,N_1119);
nand U1254 (N_1254,N_1173,N_1112);
nor U1255 (N_1255,N_1116,N_1176);
or U1256 (N_1256,N_1116,N_1170);
nand U1257 (N_1257,N_1198,N_1146);
or U1258 (N_1258,N_1109,N_1158);
nor U1259 (N_1259,N_1149,N_1132);
nor U1260 (N_1260,N_1148,N_1124);
nor U1261 (N_1261,N_1152,N_1163);
nor U1262 (N_1262,N_1188,N_1174);
nor U1263 (N_1263,N_1149,N_1175);
or U1264 (N_1264,N_1116,N_1138);
or U1265 (N_1265,N_1159,N_1151);
xnor U1266 (N_1266,N_1145,N_1176);
or U1267 (N_1267,N_1109,N_1132);
nand U1268 (N_1268,N_1124,N_1198);
nor U1269 (N_1269,N_1166,N_1165);
nand U1270 (N_1270,N_1110,N_1128);
or U1271 (N_1271,N_1159,N_1134);
nand U1272 (N_1272,N_1101,N_1183);
nand U1273 (N_1273,N_1149,N_1126);
and U1274 (N_1274,N_1150,N_1135);
nand U1275 (N_1275,N_1171,N_1114);
or U1276 (N_1276,N_1160,N_1199);
and U1277 (N_1277,N_1171,N_1145);
and U1278 (N_1278,N_1168,N_1169);
xor U1279 (N_1279,N_1180,N_1184);
xnor U1280 (N_1280,N_1116,N_1119);
xnor U1281 (N_1281,N_1192,N_1120);
nor U1282 (N_1282,N_1132,N_1129);
nand U1283 (N_1283,N_1144,N_1132);
nand U1284 (N_1284,N_1137,N_1135);
and U1285 (N_1285,N_1146,N_1101);
or U1286 (N_1286,N_1114,N_1123);
xnor U1287 (N_1287,N_1130,N_1156);
nor U1288 (N_1288,N_1144,N_1169);
or U1289 (N_1289,N_1104,N_1198);
and U1290 (N_1290,N_1100,N_1139);
nor U1291 (N_1291,N_1124,N_1108);
xor U1292 (N_1292,N_1140,N_1127);
and U1293 (N_1293,N_1127,N_1193);
nand U1294 (N_1294,N_1132,N_1176);
or U1295 (N_1295,N_1122,N_1148);
and U1296 (N_1296,N_1163,N_1102);
nor U1297 (N_1297,N_1122,N_1144);
nor U1298 (N_1298,N_1165,N_1159);
nand U1299 (N_1299,N_1133,N_1109);
and U1300 (N_1300,N_1202,N_1224);
or U1301 (N_1301,N_1256,N_1239);
nor U1302 (N_1302,N_1240,N_1269);
nor U1303 (N_1303,N_1260,N_1212);
and U1304 (N_1304,N_1245,N_1205);
nor U1305 (N_1305,N_1222,N_1261);
nand U1306 (N_1306,N_1219,N_1216);
and U1307 (N_1307,N_1211,N_1292);
or U1308 (N_1308,N_1296,N_1251);
nand U1309 (N_1309,N_1236,N_1235);
or U1310 (N_1310,N_1226,N_1290);
nand U1311 (N_1311,N_1242,N_1228);
nor U1312 (N_1312,N_1267,N_1203);
or U1313 (N_1313,N_1232,N_1247);
nand U1314 (N_1314,N_1250,N_1214);
and U1315 (N_1315,N_1273,N_1254);
and U1316 (N_1316,N_1208,N_1248);
xor U1317 (N_1317,N_1234,N_1293);
or U1318 (N_1318,N_1243,N_1271);
xnor U1319 (N_1319,N_1287,N_1299);
and U1320 (N_1320,N_1283,N_1238);
and U1321 (N_1321,N_1262,N_1215);
nor U1322 (N_1322,N_1268,N_1233);
and U1323 (N_1323,N_1282,N_1249);
or U1324 (N_1324,N_1229,N_1210);
nor U1325 (N_1325,N_1241,N_1279);
and U1326 (N_1326,N_1207,N_1277);
xor U1327 (N_1327,N_1206,N_1231);
or U1328 (N_1328,N_1274,N_1264);
nand U1329 (N_1329,N_1278,N_1200);
and U1330 (N_1330,N_1201,N_1285);
nor U1331 (N_1331,N_1246,N_1272);
and U1332 (N_1332,N_1263,N_1253);
or U1333 (N_1333,N_1266,N_1281);
and U1334 (N_1334,N_1275,N_1259);
and U1335 (N_1335,N_1244,N_1286);
nor U1336 (N_1336,N_1288,N_1225);
or U1337 (N_1337,N_1217,N_1230);
or U1338 (N_1338,N_1220,N_1291);
and U1339 (N_1339,N_1221,N_1289);
and U1340 (N_1340,N_1270,N_1258);
nor U1341 (N_1341,N_1276,N_1218);
nor U1342 (N_1342,N_1237,N_1294);
nand U1343 (N_1343,N_1280,N_1213);
and U1344 (N_1344,N_1265,N_1209);
nor U1345 (N_1345,N_1252,N_1223);
nand U1346 (N_1346,N_1227,N_1255);
or U1347 (N_1347,N_1295,N_1257);
nor U1348 (N_1348,N_1297,N_1204);
and U1349 (N_1349,N_1284,N_1298);
or U1350 (N_1350,N_1278,N_1243);
nor U1351 (N_1351,N_1229,N_1205);
nor U1352 (N_1352,N_1299,N_1297);
nand U1353 (N_1353,N_1200,N_1262);
nand U1354 (N_1354,N_1283,N_1261);
or U1355 (N_1355,N_1261,N_1256);
or U1356 (N_1356,N_1227,N_1267);
xor U1357 (N_1357,N_1298,N_1201);
and U1358 (N_1358,N_1249,N_1200);
or U1359 (N_1359,N_1256,N_1218);
or U1360 (N_1360,N_1254,N_1261);
nor U1361 (N_1361,N_1283,N_1210);
nand U1362 (N_1362,N_1201,N_1271);
nand U1363 (N_1363,N_1204,N_1222);
nand U1364 (N_1364,N_1284,N_1201);
xor U1365 (N_1365,N_1237,N_1255);
and U1366 (N_1366,N_1206,N_1213);
xnor U1367 (N_1367,N_1241,N_1257);
nand U1368 (N_1368,N_1288,N_1205);
nand U1369 (N_1369,N_1222,N_1205);
or U1370 (N_1370,N_1238,N_1286);
nor U1371 (N_1371,N_1266,N_1288);
or U1372 (N_1372,N_1225,N_1298);
nor U1373 (N_1373,N_1261,N_1293);
and U1374 (N_1374,N_1277,N_1271);
and U1375 (N_1375,N_1260,N_1233);
nor U1376 (N_1376,N_1208,N_1206);
xnor U1377 (N_1377,N_1220,N_1289);
xor U1378 (N_1378,N_1287,N_1286);
xor U1379 (N_1379,N_1241,N_1289);
xor U1380 (N_1380,N_1205,N_1218);
nor U1381 (N_1381,N_1271,N_1280);
nand U1382 (N_1382,N_1210,N_1227);
nor U1383 (N_1383,N_1299,N_1217);
nor U1384 (N_1384,N_1273,N_1243);
or U1385 (N_1385,N_1281,N_1221);
and U1386 (N_1386,N_1216,N_1257);
nand U1387 (N_1387,N_1290,N_1284);
and U1388 (N_1388,N_1226,N_1261);
nor U1389 (N_1389,N_1275,N_1249);
or U1390 (N_1390,N_1265,N_1295);
nor U1391 (N_1391,N_1236,N_1267);
or U1392 (N_1392,N_1245,N_1239);
and U1393 (N_1393,N_1299,N_1263);
nor U1394 (N_1394,N_1228,N_1265);
and U1395 (N_1395,N_1274,N_1277);
or U1396 (N_1396,N_1238,N_1250);
nand U1397 (N_1397,N_1212,N_1267);
and U1398 (N_1398,N_1245,N_1290);
nand U1399 (N_1399,N_1249,N_1287);
and U1400 (N_1400,N_1382,N_1375);
nand U1401 (N_1401,N_1385,N_1362);
xnor U1402 (N_1402,N_1338,N_1391);
nand U1403 (N_1403,N_1325,N_1304);
nor U1404 (N_1404,N_1357,N_1315);
nand U1405 (N_1405,N_1358,N_1318);
and U1406 (N_1406,N_1368,N_1372);
and U1407 (N_1407,N_1332,N_1367);
nand U1408 (N_1408,N_1398,N_1305);
nor U1409 (N_1409,N_1389,N_1335);
nor U1410 (N_1410,N_1381,N_1347);
and U1411 (N_1411,N_1333,N_1393);
nor U1412 (N_1412,N_1340,N_1309);
nor U1413 (N_1413,N_1317,N_1300);
and U1414 (N_1414,N_1380,N_1308);
nand U1415 (N_1415,N_1339,N_1306);
or U1416 (N_1416,N_1388,N_1345);
and U1417 (N_1417,N_1334,N_1322);
nand U1418 (N_1418,N_1361,N_1319);
nand U1419 (N_1419,N_1363,N_1350);
and U1420 (N_1420,N_1371,N_1330);
and U1421 (N_1421,N_1312,N_1352);
nand U1422 (N_1422,N_1310,N_1360);
xnor U1423 (N_1423,N_1311,N_1324);
and U1424 (N_1424,N_1314,N_1307);
nand U1425 (N_1425,N_1346,N_1377);
or U1426 (N_1426,N_1369,N_1355);
or U1427 (N_1427,N_1342,N_1366);
nor U1428 (N_1428,N_1301,N_1397);
or U1429 (N_1429,N_1353,N_1341);
nand U1430 (N_1430,N_1313,N_1378);
or U1431 (N_1431,N_1387,N_1364);
nand U1432 (N_1432,N_1376,N_1331);
nor U1433 (N_1433,N_1302,N_1327);
nor U1434 (N_1434,N_1336,N_1390);
or U1435 (N_1435,N_1365,N_1349);
or U1436 (N_1436,N_1386,N_1316);
nor U1437 (N_1437,N_1383,N_1326);
or U1438 (N_1438,N_1396,N_1323);
and U1439 (N_1439,N_1348,N_1399);
nand U1440 (N_1440,N_1328,N_1329);
and U1441 (N_1441,N_1303,N_1359);
or U1442 (N_1442,N_1395,N_1392);
nor U1443 (N_1443,N_1320,N_1379);
and U1444 (N_1444,N_1370,N_1394);
or U1445 (N_1445,N_1337,N_1354);
xor U1446 (N_1446,N_1373,N_1384);
nor U1447 (N_1447,N_1356,N_1344);
nor U1448 (N_1448,N_1374,N_1321);
and U1449 (N_1449,N_1343,N_1351);
and U1450 (N_1450,N_1315,N_1362);
or U1451 (N_1451,N_1327,N_1314);
and U1452 (N_1452,N_1302,N_1314);
nand U1453 (N_1453,N_1333,N_1396);
nor U1454 (N_1454,N_1377,N_1309);
nor U1455 (N_1455,N_1380,N_1376);
nand U1456 (N_1456,N_1316,N_1331);
nor U1457 (N_1457,N_1316,N_1304);
nand U1458 (N_1458,N_1394,N_1382);
and U1459 (N_1459,N_1375,N_1384);
nand U1460 (N_1460,N_1368,N_1393);
nand U1461 (N_1461,N_1317,N_1348);
nand U1462 (N_1462,N_1339,N_1325);
nand U1463 (N_1463,N_1369,N_1318);
and U1464 (N_1464,N_1313,N_1333);
nor U1465 (N_1465,N_1398,N_1337);
or U1466 (N_1466,N_1326,N_1338);
nand U1467 (N_1467,N_1305,N_1315);
or U1468 (N_1468,N_1337,N_1300);
nor U1469 (N_1469,N_1338,N_1385);
or U1470 (N_1470,N_1337,N_1340);
nor U1471 (N_1471,N_1359,N_1373);
and U1472 (N_1472,N_1346,N_1363);
nand U1473 (N_1473,N_1349,N_1386);
nor U1474 (N_1474,N_1367,N_1349);
nor U1475 (N_1475,N_1300,N_1313);
and U1476 (N_1476,N_1399,N_1377);
and U1477 (N_1477,N_1347,N_1317);
nor U1478 (N_1478,N_1397,N_1387);
or U1479 (N_1479,N_1379,N_1340);
or U1480 (N_1480,N_1311,N_1349);
nand U1481 (N_1481,N_1322,N_1347);
and U1482 (N_1482,N_1346,N_1306);
nand U1483 (N_1483,N_1392,N_1339);
and U1484 (N_1484,N_1328,N_1315);
nand U1485 (N_1485,N_1349,N_1378);
nor U1486 (N_1486,N_1382,N_1348);
or U1487 (N_1487,N_1301,N_1355);
or U1488 (N_1488,N_1305,N_1362);
xnor U1489 (N_1489,N_1330,N_1314);
nor U1490 (N_1490,N_1310,N_1356);
or U1491 (N_1491,N_1348,N_1398);
or U1492 (N_1492,N_1343,N_1361);
and U1493 (N_1493,N_1336,N_1392);
nor U1494 (N_1494,N_1337,N_1364);
nand U1495 (N_1495,N_1336,N_1398);
xnor U1496 (N_1496,N_1303,N_1372);
and U1497 (N_1497,N_1399,N_1385);
or U1498 (N_1498,N_1302,N_1315);
nand U1499 (N_1499,N_1302,N_1359);
nand U1500 (N_1500,N_1465,N_1442);
nor U1501 (N_1501,N_1463,N_1444);
nor U1502 (N_1502,N_1472,N_1490);
and U1503 (N_1503,N_1432,N_1448);
xnor U1504 (N_1504,N_1483,N_1457);
nor U1505 (N_1505,N_1458,N_1409);
and U1506 (N_1506,N_1438,N_1494);
nand U1507 (N_1507,N_1424,N_1491);
and U1508 (N_1508,N_1462,N_1489);
xnor U1509 (N_1509,N_1456,N_1436);
xor U1510 (N_1510,N_1477,N_1427);
and U1511 (N_1511,N_1499,N_1474);
and U1512 (N_1512,N_1446,N_1497);
nor U1513 (N_1513,N_1404,N_1417);
or U1514 (N_1514,N_1445,N_1471);
nor U1515 (N_1515,N_1476,N_1473);
nand U1516 (N_1516,N_1482,N_1441);
and U1517 (N_1517,N_1437,N_1493);
nor U1518 (N_1518,N_1484,N_1433);
nor U1519 (N_1519,N_1469,N_1495);
and U1520 (N_1520,N_1410,N_1418);
or U1521 (N_1521,N_1468,N_1478);
nor U1522 (N_1522,N_1440,N_1439);
nand U1523 (N_1523,N_1479,N_1461);
nand U1524 (N_1524,N_1420,N_1460);
nand U1525 (N_1525,N_1487,N_1459);
or U1526 (N_1526,N_1454,N_1492);
nor U1527 (N_1527,N_1426,N_1488);
nand U1528 (N_1528,N_1452,N_1447);
nand U1529 (N_1529,N_1421,N_1403);
and U1530 (N_1530,N_1413,N_1451);
and U1531 (N_1531,N_1466,N_1401);
or U1532 (N_1532,N_1496,N_1480);
xnor U1533 (N_1533,N_1443,N_1467);
and U1534 (N_1534,N_1415,N_1402);
and U1535 (N_1535,N_1475,N_1406);
nand U1536 (N_1536,N_1405,N_1425);
and U1537 (N_1537,N_1464,N_1411);
or U1538 (N_1538,N_1434,N_1428);
and U1539 (N_1539,N_1414,N_1485);
or U1540 (N_1540,N_1430,N_1400);
or U1541 (N_1541,N_1455,N_1470);
and U1542 (N_1542,N_1423,N_1412);
and U1543 (N_1543,N_1453,N_1435);
and U1544 (N_1544,N_1416,N_1449);
or U1545 (N_1545,N_1408,N_1481);
or U1546 (N_1546,N_1498,N_1429);
xnor U1547 (N_1547,N_1407,N_1431);
nand U1548 (N_1548,N_1422,N_1450);
nor U1549 (N_1549,N_1486,N_1419);
nor U1550 (N_1550,N_1473,N_1428);
nor U1551 (N_1551,N_1486,N_1428);
or U1552 (N_1552,N_1472,N_1452);
and U1553 (N_1553,N_1402,N_1425);
nand U1554 (N_1554,N_1463,N_1401);
and U1555 (N_1555,N_1476,N_1432);
nand U1556 (N_1556,N_1418,N_1499);
xnor U1557 (N_1557,N_1457,N_1430);
or U1558 (N_1558,N_1493,N_1402);
or U1559 (N_1559,N_1481,N_1407);
nor U1560 (N_1560,N_1429,N_1453);
nand U1561 (N_1561,N_1495,N_1486);
or U1562 (N_1562,N_1437,N_1452);
and U1563 (N_1563,N_1478,N_1474);
or U1564 (N_1564,N_1455,N_1465);
xnor U1565 (N_1565,N_1463,N_1471);
nor U1566 (N_1566,N_1404,N_1473);
or U1567 (N_1567,N_1495,N_1404);
or U1568 (N_1568,N_1439,N_1422);
nand U1569 (N_1569,N_1401,N_1443);
or U1570 (N_1570,N_1483,N_1403);
and U1571 (N_1571,N_1436,N_1459);
nand U1572 (N_1572,N_1416,N_1444);
or U1573 (N_1573,N_1479,N_1403);
nor U1574 (N_1574,N_1474,N_1493);
or U1575 (N_1575,N_1499,N_1475);
and U1576 (N_1576,N_1451,N_1470);
and U1577 (N_1577,N_1450,N_1461);
or U1578 (N_1578,N_1487,N_1470);
and U1579 (N_1579,N_1469,N_1416);
nand U1580 (N_1580,N_1421,N_1401);
nor U1581 (N_1581,N_1413,N_1443);
xnor U1582 (N_1582,N_1431,N_1430);
xor U1583 (N_1583,N_1418,N_1446);
and U1584 (N_1584,N_1465,N_1412);
nor U1585 (N_1585,N_1400,N_1415);
xnor U1586 (N_1586,N_1411,N_1432);
nand U1587 (N_1587,N_1458,N_1477);
or U1588 (N_1588,N_1457,N_1406);
or U1589 (N_1589,N_1443,N_1416);
nand U1590 (N_1590,N_1415,N_1418);
and U1591 (N_1591,N_1426,N_1474);
or U1592 (N_1592,N_1446,N_1449);
nor U1593 (N_1593,N_1430,N_1471);
nand U1594 (N_1594,N_1419,N_1420);
and U1595 (N_1595,N_1466,N_1490);
and U1596 (N_1596,N_1476,N_1463);
xor U1597 (N_1597,N_1425,N_1407);
or U1598 (N_1598,N_1421,N_1431);
or U1599 (N_1599,N_1434,N_1431);
xnor U1600 (N_1600,N_1533,N_1557);
nand U1601 (N_1601,N_1584,N_1513);
nor U1602 (N_1602,N_1587,N_1575);
xnor U1603 (N_1603,N_1592,N_1585);
nand U1604 (N_1604,N_1554,N_1560);
and U1605 (N_1605,N_1543,N_1586);
nor U1606 (N_1606,N_1590,N_1540);
or U1607 (N_1607,N_1527,N_1598);
or U1608 (N_1608,N_1582,N_1503);
and U1609 (N_1609,N_1546,N_1530);
xnor U1610 (N_1610,N_1580,N_1550);
or U1611 (N_1611,N_1552,N_1571);
or U1612 (N_1612,N_1593,N_1594);
nor U1613 (N_1613,N_1531,N_1507);
nand U1614 (N_1614,N_1526,N_1538);
and U1615 (N_1615,N_1588,N_1569);
and U1616 (N_1616,N_1559,N_1561);
or U1617 (N_1617,N_1547,N_1570);
and U1618 (N_1618,N_1555,N_1548);
nand U1619 (N_1619,N_1562,N_1577);
or U1620 (N_1620,N_1520,N_1535);
or U1621 (N_1621,N_1558,N_1565);
and U1622 (N_1622,N_1532,N_1511);
or U1623 (N_1623,N_1524,N_1505);
nand U1624 (N_1624,N_1504,N_1502);
xnor U1625 (N_1625,N_1572,N_1508);
nor U1626 (N_1626,N_1545,N_1541);
nand U1627 (N_1627,N_1512,N_1551);
nor U1628 (N_1628,N_1506,N_1578);
and U1629 (N_1629,N_1581,N_1516);
nor U1630 (N_1630,N_1500,N_1549);
or U1631 (N_1631,N_1556,N_1514);
nor U1632 (N_1632,N_1544,N_1539);
or U1633 (N_1633,N_1521,N_1510);
nor U1634 (N_1634,N_1597,N_1525);
or U1635 (N_1635,N_1519,N_1595);
nor U1636 (N_1636,N_1564,N_1583);
or U1637 (N_1637,N_1509,N_1528);
xnor U1638 (N_1638,N_1563,N_1596);
or U1639 (N_1639,N_1591,N_1566);
nor U1640 (N_1640,N_1536,N_1515);
and U1641 (N_1641,N_1518,N_1574);
nand U1642 (N_1642,N_1534,N_1589);
or U1643 (N_1643,N_1576,N_1529);
xor U1644 (N_1644,N_1567,N_1517);
nor U1645 (N_1645,N_1542,N_1522);
and U1646 (N_1646,N_1501,N_1523);
and U1647 (N_1647,N_1573,N_1568);
xor U1648 (N_1648,N_1599,N_1579);
nand U1649 (N_1649,N_1553,N_1537);
nor U1650 (N_1650,N_1532,N_1516);
xor U1651 (N_1651,N_1587,N_1562);
xor U1652 (N_1652,N_1542,N_1569);
and U1653 (N_1653,N_1529,N_1511);
and U1654 (N_1654,N_1540,N_1568);
nor U1655 (N_1655,N_1588,N_1514);
and U1656 (N_1656,N_1567,N_1573);
xnor U1657 (N_1657,N_1575,N_1570);
and U1658 (N_1658,N_1549,N_1522);
nand U1659 (N_1659,N_1563,N_1507);
nand U1660 (N_1660,N_1538,N_1530);
nor U1661 (N_1661,N_1557,N_1536);
nor U1662 (N_1662,N_1528,N_1562);
nand U1663 (N_1663,N_1584,N_1573);
or U1664 (N_1664,N_1549,N_1599);
nor U1665 (N_1665,N_1592,N_1574);
nor U1666 (N_1666,N_1545,N_1519);
or U1667 (N_1667,N_1562,N_1510);
xnor U1668 (N_1668,N_1599,N_1564);
nor U1669 (N_1669,N_1543,N_1565);
xor U1670 (N_1670,N_1544,N_1549);
or U1671 (N_1671,N_1581,N_1597);
and U1672 (N_1672,N_1515,N_1540);
nand U1673 (N_1673,N_1534,N_1578);
nand U1674 (N_1674,N_1540,N_1531);
nand U1675 (N_1675,N_1511,N_1531);
nand U1676 (N_1676,N_1560,N_1573);
nor U1677 (N_1677,N_1577,N_1567);
nor U1678 (N_1678,N_1504,N_1561);
nand U1679 (N_1679,N_1560,N_1537);
and U1680 (N_1680,N_1534,N_1575);
xor U1681 (N_1681,N_1599,N_1515);
xor U1682 (N_1682,N_1564,N_1546);
or U1683 (N_1683,N_1537,N_1566);
nor U1684 (N_1684,N_1549,N_1561);
nor U1685 (N_1685,N_1592,N_1572);
nor U1686 (N_1686,N_1597,N_1596);
nand U1687 (N_1687,N_1517,N_1588);
nand U1688 (N_1688,N_1567,N_1572);
nand U1689 (N_1689,N_1531,N_1506);
nand U1690 (N_1690,N_1525,N_1557);
or U1691 (N_1691,N_1520,N_1586);
nor U1692 (N_1692,N_1517,N_1560);
xor U1693 (N_1693,N_1515,N_1577);
nor U1694 (N_1694,N_1595,N_1542);
xor U1695 (N_1695,N_1580,N_1508);
nor U1696 (N_1696,N_1515,N_1569);
nor U1697 (N_1697,N_1575,N_1571);
or U1698 (N_1698,N_1549,N_1591);
xor U1699 (N_1699,N_1500,N_1505);
nor U1700 (N_1700,N_1655,N_1662);
nand U1701 (N_1701,N_1604,N_1638);
and U1702 (N_1702,N_1676,N_1620);
nand U1703 (N_1703,N_1666,N_1643);
xor U1704 (N_1704,N_1652,N_1653);
xnor U1705 (N_1705,N_1665,N_1635);
xnor U1706 (N_1706,N_1630,N_1657);
nand U1707 (N_1707,N_1696,N_1632);
and U1708 (N_1708,N_1681,N_1646);
or U1709 (N_1709,N_1627,N_1661);
nand U1710 (N_1710,N_1602,N_1624);
and U1711 (N_1711,N_1685,N_1656);
and U1712 (N_1712,N_1617,N_1687);
nand U1713 (N_1713,N_1671,N_1697);
nor U1714 (N_1714,N_1629,N_1667);
or U1715 (N_1715,N_1686,N_1699);
nand U1716 (N_1716,N_1669,N_1619);
nand U1717 (N_1717,N_1695,N_1616);
nand U1718 (N_1718,N_1664,N_1672);
nand U1719 (N_1719,N_1626,N_1621);
or U1720 (N_1720,N_1654,N_1623);
nor U1721 (N_1721,N_1608,N_1609);
or U1722 (N_1722,N_1633,N_1613);
and U1723 (N_1723,N_1688,N_1674);
nor U1724 (N_1724,N_1658,N_1600);
nor U1725 (N_1725,N_1615,N_1678);
or U1726 (N_1726,N_1650,N_1648);
nor U1727 (N_1727,N_1628,N_1689);
nand U1728 (N_1728,N_1673,N_1668);
and U1729 (N_1729,N_1603,N_1618);
nand U1730 (N_1730,N_1607,N_1684);
nand U1731 (N_1731,N_1641,N_1631);
nor U1732 (N_1732,N_1636,N_1683);
or U1733 (N_1733,N_1670,N_1677);
nand U1734 (N_1734,N_1691,N_1614);
nor U1735 (N_1735,N_1644,N_1606);
nand U1736 (N_1736,N_1692,N_1612);
nor U1737 (N_1737,N_1610,N_1611);
or U1738 (N_1738,N_1651,N_1682);
nand U1739 (N_1739,N_1698,N_1640);
and U1740 (N_1740,N_1675,N_1642);
nor U1741 (N_1741,N_1637,N_1663);
or U1742 (N_1742,N_1605,N_1625);
nor U1743 (N_1743,N_1622,N_1601);
xnor U1744 (N_1744,N_1645,N_1647);
nor U1745 (N_1745,N_1690,N_1659);
nand U1746 (N_1746,N_1649,N_1679);
and U1747 (N_1747,N_1693,N_1680);
nand U1748 (N_1748,N_1694,N_1634);
nor U1749 (N_1749,N_1660,N_1639);
nor U1750 (N_1750,N_1686,N_1677);
or U1751 (N_1751,N_1625,N_1649);
nand U1752 (N_1752,N_1677,N_1694);
or U1753 (N_1753,N_1698,N_1663);
or U1754 (N_1754,N_1652,N_1630);
xor U1755 (N_1755,N_1627,N_1674);
xor U1756 (N_1756,N_1696,N_1671);
xnor U1757 (N_1757,N_1639,N_1679);
nand U1758 (N_1758,N_1611,N_1670);
nand U1759 (N_1759,N_1670,N_1686);
and U1760 (N_1760,N_1604,N_1673);
nand U1761 (N_1761,N_1685,N_1648);
or U1762 (N_1762,N_1601,N_1693);
or U1763 (N_1763,N_1653,N_1622);
nand U1764 (N_1764,N_1671,N_1611);
or U1765 (N_1765,N_1690,N_1602);
nand U1766 (N_1766,N_1681,N_1699);
nand U1767 (N_1767,N_1628,N_1650);
nor U1768 (N_1768,N_1684,N_1613);
nor U1769 (N_1769,N_1619,N_1695);
nand U1770 (N_1770,N_1657,N_1614);
nand U1771 (N_1771,N_1698,N_1643);
nor U1772 (N_1772,N_1675,N_1639);
and U1773 (N_1773,N_1697,N_1699);
nand U1774 (N_1774,N_1663,N_1617);
or U1775 (N_1775,N_1694,N_1620);
or U1776 (N_1776,N_1634,N_1685);
xnor U1777 (N_1777,N_1697,N_1637);
or U1778 (N_1778,N_1699,N_1693);
or U1779 (N_1779,N_1625,N_1604);
nor U1780 (N_1780,N_1648,N_1658);
or U1781 (N_1781,N_1635,N_1680);
nor U1782 (N_1782,N_1657,N_1698);
xor U1783 (N_1783,N_1641,N_1658);
nand U1784 (N_1784,N_1613,N_1652);
nand U1785 (N_1785,N_1684,N_1639);
or U1786 (N_1786,N_1642,N_1611);
nor U1787 (N_1787,N_1613,N_1645);
nor U1788 (N_1788,N_1629,N_1696);
xor U1789 (N_1789,N_1610,N_1659);
and U1790 (N_1790,N_1688,N_1653);
and U1791 (N_1791,N_1643,N_1676);
and U1792 (N_1792,N_1666,N_1625);
or U1793 (N_1793,N_1616,N_1600);
or U1794 (N_1794,N_1661,N_1679);
nand U1795 (N_1795,N_1620,N_1686);
nor U1796 (N_1796,N_1657,N_1691);
and U1797 (N_1797,N_1681,N_1622);
nand U1798 (N_1798,N_1619,N_1689);
or U1799 (N_1799,N_1687,N_1626);
and U1800 (N_1800,N_1730,N_1705);
nor U1801 (N_1801,N_1726,N_1782);
nor U1802 (N_1802,N_1783,N_1703);
or U1803 (N_1803,N_1752,N_1733);
and U1804 (N_1804,N_1785,N_1713);
nand U1805 (N_1805,N_1711,N_1773);
nor U1806 (N_1806,N_1731,N_1774);
xnor U1807 (N_1807,N_1793,N_1780);
and U1808 (N_1808,N_1717,N_1707);
and U1809 (N_1809,N_1790,N_1712);
or U1810 (N_1810,N_1746,N_1744);
nand U1811 (N_1811,N_1702,N_1714);
or U1812 (N_1812,N_1796,N_1745);
nor U1813 (N_1813,N_1753,N_1722);
or U1814 (N_1814,N_1768,N_1741);
nand U1815 (N_1815,N_1750,N_1797);
nand U1816 (N_1816,N_1781,N_1716);
and U1817 (N_1817,N_1736,N_1789);
nand U1818 (N_1818,N_1786,N_1791);
nor U1819 (N_1819,N_1777,N_1764);
and U1820 (N_1820,N_1735,N_1765);
or U1821 (N_1821,N_1719,N_1792);
or U1822 (N_1822,N_1779,N_1776);
xor U1823 (N_1823,N_1759,N_1739);
nand U1824 (N_1824,N_1729,N_1706);
nand U1825 (N_1825,N_1799,N_1798);
or U1826 (N_1826,N_1701,N_1721);
nor U1827 (N_1827,N_1715,N_1727);
nor U1828 (N_1828,N_1700,N_1740);
nand U1829 (N_1829,N_1761,N_1755);
nor U1830 (N_1830,N_1732,N_1751);
xnor U1831 (N_1831,N_1762,N_1794);
or U1832 (N_1832,N_1756,N_1766);
nand U1833 (N_1833,N_1760,N_1742);
nor U1834 (N_1834,N_1738,N_1704);
nor U1835 (N_1835,N_1795,N_1770);
or U1836 (N_1836,N_1754,N_1772);
nand U1837 (N_1837,N_1743,N_1725);
and U1838 (N_1838,N_1718,N_1771);
and U1839 (N_1839,N_1710,N_1767);
or U1840 (N_1840,N_1757,N_1763);
nand U1841 (N_1841,N_1787,N_1758);
or U1842 (N_1842,N_1723,N_1788);
or U1843 (N_1843,N_1749,N_1734);
nor U1844 (N_1844,N_1709,N_1724);
and U1845 (N_1845,N_1708,N_1737);
nand U1846 (N_1846,N_1775,N_1748);
and U1847 (N_1847,N_1720,N_1784);
nand U1848 (N_1848,N_1769,N_1778);
or U1849 (N_1849,N_1728,N_1747);
nor U1850 (N_1850,N_1789,N_1775);
nor U1851 (N_1851,N_1777,N_1727);
or U1852 (N_1852,N_1777,N_1760);
and U1853 (N_1853,N_1703,N_1749);
or U1854 (N_1854,N_1737,N_1711);
and U1855 (N_1855,N_1749,N_1782);
xnor U1856 (N_1856,N_1741,N_1710);
or U1857 (N_1857,N_1753,N_1721);
xnor U1858 (N_1858,N_1790,N_1729);
and U1859 (N_1859,N_1736,N_1743);
or U1860 (N_1860,N_1783,N_1763);
nor U1861 (N_1861,N_1752,N_1705);
nand U1862 (N_1862,N_1710,N_1724);
nor U1863 (N_1863,N_1777,N_1785);
nand U1864 (N_1864,N_1730,N_1740);
nor U1865 (N_1865,N_1788,N_1771);
nor U1866 (N_1866,N_1736,N_1777);
nand U1867 (N_1867,N_1780,N_1785);
and U1868 (N_1868,N_1752,N_1740);
nor U1869 (N_1869,N_1764,N_1709);
and U1870 (N_1870,N_1763,N_1768);
nand U1871 (N_1871,N_1786,N_1724);
xnor U1872 (N_1872,N_1748,N_1764);
nand U1873 (N_1873,N_1779,N_1743);
or U1874 (N_1874,N_1786,N_1753);
nor U1875 (N_1875,N_1779,N_1706);
nor U1876 (N_1876,N_1736,N_1756);
or U1877 (N_1877,N_1712,N_1734);
or U1878 (N_1878,N_1774,N_1741);
or U1879 (N_1879,N_1763,N_1785);
or U1880 (N_1880,N_1763,N_1777);
nor U1881 (N_1881,N_1730,N_1781);
nand U1882 (N_1882,N_1719,N_1738);
and U1883 (N_1883,N_1765,N_1764);
nor U1884 (N_1884,N_1762,N_1769);
and U1885 (N_1885,N_1797,N_1753);
nor U1886 (N_1886,N_1788,N_1757);
nor U1887 (N_1887,N_1792,N_1755);
nor U1888 (N_1888,N_1733,N_1719);
or U1889 (N_1889,N_1790,N_1719);
nand U1890 (N_1890,N_1724,N_1747);
nor U1891 (N_1891,N_1737,N_1742);
nand U1892 (N_1892,N_1708,N_1733);
and U1893 (N_1893,N_1761,N_1787);
nor U1894 (N_1894,N_1741,N_1724);
xnor U1895 (N_1895,N_1767,N_1729);
or U1896 (N_1896,N_1775,N_1767);
or U1897 (N_1897,N_1723,N_1787);
xnor U1898 (N_1898,N_1704,N_1774);
nor U1899 (N_1899,N_1712,N_1737);
nor U1900 (N_1900,N_1871,N_1845);
or U1901 (N_1901,N_1814,N_1875);
nand U1902 (N_1902,N_1857,N_1873);
or U1903 (N_1903,N_1829,N_1892);
and U1904 (N_1904,N_1835,N_1839);
nor U1905 (N_1905,N_1885,N_1819);
nor U1906 (N_1906,N_1836,N_1821);
or U1907 (N_1907,N_1846,N_1801);
and U1908 (N_1908,N_1897,N_1812);
or U1909 (N_1909,N_1802,N_1820);
or U1910 (N_1910,N_1877,N_1848);
nand U1911 (N_1911,N_1809,N_1816);
nor U1912 (N_1912,N_1842,N_1825);
and U1913 (N_1913,N_1804,N_1840);
or U1914 (N_1914,N_1890,N_1863);
nand U1915 (N_1915,N_1869,N_1843);
nand U1916 (N_1916,N_1859,N_1824);
or U1917 (N_1917,N_1889,N_1817);
nor U1918 (N_1918,N_1883,N_1876);
nor U1919 (N_1919,N_1822,N_1818);
and U1920 (N_1920,N_1841,N_1853);
nor U1921 (N_1921,N_1828,N_1838);
and U1922 (N_1922,N_1815,N_1803);
and U1923 (N_1923,N_1896,N_1830);
or U1924 (N_1924,N_1806,N_1811);
nand U1925 (N_1925,N_1854,N_1847);
or U1926 (N_1926,N_1810,N_1881);
nand U1927 (N_1927,N_1831,N_1850);
and U1928 (N_1928,N_1837,N_1882);
or U1929 (N_1929,N_1844,N_1895);
xnor U1930 (N_1930,N_1833,N_1805);
or U1931 (N_1931,N_1827,N_1880);
nor U1932 (N_1932,N_1856,N_1823);
nand U1933 (N_1933,N_1878,N_1868);
or U1934 (N_1934,N_1813,N_1884);
nor U1935 (N_1935,N_1894,N_1861);
nand U1936 (N_1936,N_1826,N_1891);
or U1937 (N_1937,N_1865,N_1807);
or U1938 (N_1938,N_1832,N_1852);
nor U1939 (N_1939,N_1898,N_1834);
and U1940 (N_1940,N_1849,N_1800);
nand U1941 (N_1941,N_1864,N_1888);
nand U1942 (N_1942,N_1893,N_1866);
and U1943 (N_1943,N_1851,N_1862);
or U1944 (N_1944,N_1858,N_1899);
and U1945 (N_1945,N_1887,N_1855);
or U1946 (N_1946,N_1860,N_1879);
nand U1947 (N_1947,N_1872,N_1808);
and U1948 (N_1948,N_1874,N_1870);
or U1949 (N_1949,N_1886,N_1867);
xor U1950 (N_1950,N_1840,N_1860);
or U1951 (N_1951,N_1871,N_1824);
or U1952 (N_1952,N_1897,N_1849);
or U1953 (N_1953,N_1878,N_1847);
xor U1954 (N_1954,N_1850,N_1889);
nor U1955 (N_1955,N_1888,N_1810);
or U1956 (N_1956,N_1868,N_1875);
nand U1957 (N_1957,N_1827,N_1809);
and U1958 (N_1958,N_1816,N_1881);
nand U1959 (N_1959,N_1868,N_1870);
nand U1960 (N_1960,N_1889,N_1860);
nand U1961 (N_1961,N_1836,N_1846);
and U1962 (N_1962,N_1872,N_1855);
and U1963 (N_1963,N_1875,N_1883);
xnor U1964 (N_1964,N_1863,N_1806);
nor U1965 (N_1965,N_1859,N_1823);
or U1966 (N_1966,N_1803,N_1830);
xnor U1967 (N_1967,N_1818,N_1842);
nor U1968 (N_1968,N_1856,N_1850);
nand U1969 (N_1969,N_1853,N_1871);
or U1970 (N_1970,N_1827,N_1832);
and U1971 (N_1971,N_1888,N_1827);
and U1972 (N_1972,N_1806,N_1843);
nand U1973 (N_1973,N_1810,N_1843);
and U1974 (N_1974,N_1857,N_1861);
nand U1975 (N_1975,N_1880,N_1898);
nand U1976 (N_1976,N_1828,N_1806);
nand U1977 (N_1977,N_1852,N_1844);
or U1978 (N_1978,N_1828,N_1865);
nor U1979 (N_1979,N_1866,N_1865);
and U1980 (N_1980,N_1860,N_1863);
or U1981 (N_1981,N_1876,N_1893);
and U1982 (N_1982,N_1889,N_1851);
nor U1983 (N_1983,N_1887,N_1808);
nor U1984 (N_1984,N_1858,N_1872);
xor U1985 (N_1985,N_1846,N_1889);
and U1986 (N_1986,N_1819,N_1823);
or U1987 (N_1987,N_1872,N_1807);
and U1988 (N_1988,N_1880,N_1825);
or U1989 (N_1989,N_1810,N_1856);
and U1990 (N_1990,N_1898,N_1831);
nand U1991 (N_1991,N_1869,N_1804);
nor U1992 (N_1992,N_1869,N_1831);
and U1993 (N_1993,N_1847,N_1823);
and U1994 (N_1994,N_1823,N_1872);
nand U1995 (N_1995,N_1879,N_1881);
or U1996 (N_1996,N_1847,N_1866);
or U1997 (N_1997,N_1829,N_1802);
nand U1998 (N_1998,N_1866,N_1894);
nand U1999 (N_1999,N_1887,N_1823);
or U2000 (N_2000,N_1929,N_1998);
nor U2001 (N_2001,N_1957,N_1904);
nor U2002 (N_2002,N_1902,N_1983);
or U2003 (N_2003,N_1913,N_1905);
or U2004 (N_2004,N_1926,N_1985);
and U2005 (N_2005,N_1987,N_1934);
nor U2006 (N_2006,N_1996,N_1971);
nand U2007 (N_2007,N_1901,N_1940);
nand U2008 (N_2008,N_1915,N_1943);
and U2009 (N_2009,N_1922,N_1962);
nand U2010 (N_2010,N_1997,N_1936);
nor U2011 (N_2011,N_1908,N_1993);
nor U2012 (N_2012,N_1927,N_1925);
and U2013 (N_2013,N_1961,N_1963);
nand U2014 (N_2014,N_1960,N_1965);
and U2015 (N_2015,N_1931,N_1939);
nand U2016 (N_2016,N_1919,N_1967);
and U2017 (N_2017,N_1968,N_1935);
xor U2018 (N_2018,N_1914,N_1944);
and U2019 (N_2019,N_1949,N_1991);
nor U2020 (N_2020,N_1953,N_1992);
and U2021 (N_2021,N_1972,N_1903);
nand U2022 (N_2022,N_1938,N_1964);
nand U2023 (N_2023,N_1924,N_1916);
nor U2024 (N_2024,N_1973,N_1969);
nand U2025 (N_2025,N_1970,N_1946);
nand U2026 (N_2026,N_1910,N_1945);
nor U2027 (N_2027,N_1977,N_1900);
nor U2028 (N_2028,N_1933,N_1999);
nand U2029 (N_2029,N_1952,N_1941);
and U2030 (N_2030,N_1958,N_1989);
or U2031 (N_2031,N_1986,N_1909);
and U2032 (N_2032,N_1912,N_1917);
and U2033 (N_2033,N_1930,N_1918);
nand U2034 (N_2034,N_1982,N_1956);
nor U2035 (N_2035,N_1948,N_1955);
or U2036 (N_2036,N_1950,N_1942);
nor U2037 (N_2037,N_1920,N_1954);
or U2038 (N_2038,N_1981,N_1923);
or U2039 (N_2039,N_1978,N_1932);
xnor U2040 (N_2040,N_1951,N_1906);
nand U2041 (N_2041,N_1975,N_1966);
or U2042 (N_2042,N_1980,N_1928);
nand U2043 (N_2043,N_1911,N_1979);
nand U2044 (N_2044,N_1974,N_1984);
and U2045 (N_2045,N_1959,N_1976);
nor U2046 (N_2046,N_1995,N_1921);
nor U2047 (N_2047,N_1988,N_1947);
xnor U2048 (N_2048,N_1990,N_1994);
nor U2049 (N_2049,N_1907,N_1937);
nor U2050 (N_2050,N_1997,N_1908);
nand U2051 (N_2051,N_1993,N_1900);
and U2052 (N_2052,N_1985,N_1907);
nand U2053 (N_2053,N_1992,N_1946);
or U2054 (N_2054,N_1957,N_1902);
and U2055 (N_2055,N_1966,N_1945);
or U2056 (N_2056,N_1964,N_1998);
and U2057 (N_2057,N_1971,N_1970);
nor U2058 (N_2058,N_1983,N_1982);
nor U2059 (N_2059,N_1994,N_1909);
nor U2060 (N_2060,N_1982,N_1913);
nor U2061 (N_2061,N_1991,N_1988);
or U2062 (N_2062,N_1965,N_1913);
or U2063 (N_2063,N_1936,N_1973);
nor U2064 (N_2064,N_1941,N_1988);
or U2065 (N_2065,N_1906,N_1930);
and U2066 (N_2066,N_1992,N_1926);
or U2067 (N_2067,N_1933,N_1939);
nand U2068 (N_2068,N_1930,N_1940);
nand U2069 (N_2069,N_1975,N_1907);
or U2070 (N_2070,N_1915,N_1900);
nand U2071 (N_2071,N_1908,N_1906);
nor U2072 (N_2072,N_1920,N_1946);
or U2073 (N_2073,N_1985,N_1994);
nor U2074 (N_2074,N_1920,N_1971);
nand U2075 (N_2075,N_1938,N_1915);
nor U2076 (N_2076,N_1926,N_1982);
and U2077 (N_2077,N_1963,N_1925);
and U2078 (N_2078,N_1917,N_1941);
or U2079 (N_2079,N_1920,N_1962);
and U2080 (N_2080,N_1907,N_1922);
or U2081 (N_2081,N_1981,N_1942);
xor U2082 (N_2082,N_1934,N_1989);
nor U2083 (N_2083,N_1946,N_1940);
and U2084 (N_2084,N_1930,N_1948);
xnor U2085 (N_2085,N_1937,N_1905);
nand U2086 (N_2086,N_1975,N_1950);
or U2087 (N_2087,N_1913,N_1999);
nand U2088 (N_2088,N_1960,N_1972);
xnor U2089 (N_2089,N_1996,N_1912);
and U2090 (N_2090,N_1985,N_1906);
and U2091 (N_2091,N_1915,N_1988);
nand U2092 (N_2092,N_1998,N_1926);
and U2093 (N_2093,N_1979,N_1960);
xnor U2094 (N_2094,N_1977,N_1916);
nor U2095 (N_2095,N_1994,N_1956);
and U2096 (N_2096,N_1908,N_1952);
nand U2097 (N_2097,N_1927,N_1990);
or U2098 (N_2098,N_1989,N_1904);
nor U2099 (N_2099,N_1970,N_1950);
or U2100 (N_2100,N_2095,N_2046);
nor U2101 (N_2101,N_2080,N_2072);
and U2102 (N_2102,N_2082,N_2028);
nor U2103 (N_2103,N_2074,N_2056);
nor U2104 (N_2104,N_2088,N_2050);
nand U2105 (N_2105,N_2043,N_2065);
xor U2106 (N_2106,N_2003,N_2020);
nor U2107 (N_2107,N_2045,N_2034);
nand U2108 (N_2108,N_2039,N_2077);
nand U2109 (N_2109,N_2002,N_2029);
and U2110 (N_2110,N_2083,N_2016);
nor U2111 (N_2111,N_2036,N_2025);
nand U2112 (N_2112,N_2057,N_2093);
nor U2113 (N_2113,N_2076,N_2086);
nand U2114 (N_2114,N_2049,N_2097);
or U2115 (N_2115,N_2098,N_2079);
nand U2116 (N_2116,N_2087,N_2011);
and U2117 (N_2117,N_2038,N_2075);
or U2118 (N_2118,N_2084,N_2009);
nand U2119 (N_2119,N_2019,N_2042);
nand U2120 (N_2120,N_2015,N_2067);
nand U2121 (N_2121,N_2012,N_2017);
and U2122 (N_2122,N_2051,N_2001);
nor U2123 (N_2123,N_2047,N_2078);
xnor U2124 (N_2124,N_2091,N_2007);
nor U2125 (N_2125,N_2030,N_2069);
and U2126 (N_2126,N_2018,N_2035);
nand U2127 (N_2127,N_2032,N_2037);
and U2128 (N_2128,N_2089,N_2006);
nand U2129 (N_2129,N_2099,N_2070);
nand U2130 (N_2130,N_2033,N_2063);
nand U2131 (N_2131,N_2053,N_2021);
xnor U2132 (N_2132,N_2048,N_2062);
and U2133 (N_2133,N_2054,N_2026);
xnor U2134 (N_2134,N_2014,N_2092);
nand U2135 (N_2135,N_2068,N_2041);
nand U2136 (N_2136,N_2013,N_2000);
or U2137 (N_2137,N_2096,N_2073);
and U2138 (N_2138,N_2060,N_2024);
nand U2139 (N_2139,N_2090,N_2066);
and U2140 (N_2140,N_2008,N_2044);
and U2141 (N_2141,N_2031,N_2010);
nand U2142 (N_2142,N_2052,N_2058);
or U2143 (N_2143,N_2055,N_2023);
and U2144 (N_2144,N_2081,N_2004);
nor U2145 (N_2145,N_2022,N_2027);
nand U2146 (N_2146,N_2005,N_2064);
or U2147 (N_2147,N_2061,N_2040);
nand U2148 (N_2148,N_2071,N_2059);
nor U2149 (N_2149,N_2085,N_2094);
nand U2150 (N_2150,N_2095,N_2042);
nor U2151 (N_2151,N_2038,N_2051);
xnor U2152 (N_2152,N_2054,N_2036);
nand U2153 (N_2153,N_2002,N_2036);
and U2154 (N_2154,N_2037,N_2042);
and U2155 (N_2155,N_2005,N_2075);
nand U2156 (N_2156,N_2023,N_2059);
or U2157 (N_2157,N_2090,N_2037);
xor U2158 (N_2158,N_2045,N_2066);
and U2159 (N_2159,N_2025,N_2043);
nand U2160 (N_2160,N_2005,N_2024);
or U2161 (N_2161,N_2072,N_2040);
and U2162 (N_2162,N_2084,N_2051);
and U2163 (N_2163,N_2072,N_2069);
or U2164 (N_2164,N_2088,N_2026);
and U2165 (N_2165,N_2003,N_2082);
nor U2166 (N_2166,N_2077,N_2049);
or U2167 (N_2167,N_2073,N_2045);
or U2168 (N_2168,N_2039,N_2081);
nor U2169 (N_2169,N_2024,N_2083);
or U2170 (N_2170,N_2079,N_2077);
nor U2171 (N_2171,N_2066,N_2080);
nand U2172 (N_2172,N_2066,N_2020);
or U2173 (N_2173,N_2022,N_2039);
or U2174 (N_2174,N_2007,N_2066);
or U2175 (N_2175,N_2097,N_2079);
or U2176 (N_2176,N_2021,N_2007);
or U2177 (N_2177,N_2066,N_2091);
and U2178 (N_2178,N_2047,N_2009);
or U2179 (N_2179,N_2000,N_2042);
nand U2180 (N_2180,N_2069,N_2059);
nor U2181 (N_2181,N_2057,N_2052);
xor U2182 (N_2182,N_2051,N_2064);
nand U2183 (N_2183,N_2089,N_2024);
or U2184 (N_2184,N_2008,N_2027);
nand U2185 (N_2185,N_2017,N_2040);
xor U2186 (N_2186,N_2098,N_2001);
nor U2187 (N_2187,N_2078,N_2056);
or U2188 (N_2188,N_2061,N_2081);
nand U2189 (N_2189,N_2025,N_2074);
and U2190 (N_2190,N_2047,N_2023);
nor U2191 (N_2191,N_2057,N_2082);
nand U2192 (N_2192,N_2008,N_2099);
nand U2193 (N_2193,N_2004,N_2023);
nand U2194 (N_2194,N_2072,N_2085);
or U2195 (N_2195,N_2062,N_2052);
and U2196 (N_2196,N_2021,N_2012);
or U2197 (N_2197,N_2038,N_2087);
nor U2198 (N_2198,N_2014,N_2017);
or U2199 (N_2199,N_2057,N_2019);
or U2200 (N_2200,N_2175,N_2154);
nand U2201 (N_2201,N_2173,N_2110);
nand U2202 (N_2202,N_2106,N_2189);
nor U2203 (N_2203,N_2119,N_2179);
and U2204 (N_2204,N_2123,N_2109);
xor U2205 (N_2205,N_2118,N_2127);
and U2206 (N_2206,N_2131,N_2139);
or U2207 (N_2207,N_2187,N_2149);
nor U2208 (N_2208,N_2143,N_2103);
or U2209 (N_2209,N_2152,N_2181);
and U2210 (N_2210,N_2141,N_2162);
nor U2211 (N_2211,N_2120,N_2177);
and U2212 (N_2212,N_2137,N_2196);
or U2213 (N_2213,N_2182,N_2155);
nor U2214 (N_2214,N_2134,N_2164);
and U2215 (N_2215,N_2153,N_2113);
or U2216 (N_2216,N_2133,N_2115);
or U2217 (N_2217,N_2107,N_2197);
and U2218 (N_2218,N_2171,N_2104);
nor U2219 (N_2219,N_2100,N_2136);
and U2220 (N_2220,N_2193,N_2101);
xor U2221 (N_2221,N_2116,N_2159);
nor U2222 (N_2222,N_2169,N_2126);
nand U2223 (N_2223,N_2130,N_2135);
nand U2224 (N_2224,N_2122,N_2172);
or U2225 (N_2225,N_2147,N_2102);
nand U2226 (N_2226,N_2186,N_2156);
nor U2227 (N_2227,N_2121,N_2158);
nand U2228 (N_2228,N_2178,N_2114);
and U2229 (N_2229,N_2163,N_2170);
xnor U2230 (N_2230,N_2132,N_2176);
xor U2231 (N_2231,N_2192,N_2112);
or U2232 (N_2232,N_2125,N_2195);
xor U2233 (N_2233,N_2145,N_2183);
or U2234 (N_2234,N_2146,N_2150);
nor U2235 (N_2235,N_2142,N_2151);
nand U2236 (N_2236,N_2144,N_2129);
and U2237 (N_2237,N_2111,N_2165);
nor U2238 (N_2238,N_2166,N_2108);
nor U2239 (N_2239,N_2174,N_2117);
or U2240 (N_2240,N_2199,N_2160);
and U2241 (N_2241,N_2161,N_2124);
nor U2242 (N_2242,N_2194,N_2167);
nand U2243 (N_2243,N_2148,N_2185);
nand U2244 (N_2244,N_2184,N_2168);
xor U2245 (N_2245,N_2128,N_2140);
and U2246 (N_2246,N_2157,N_2180);
or U2247 (N_2247,N_2138,N_2188);
and U2248 (N_2248,N_2198,N_2105);
nor U2249 (N_2249,N_2190,N_2191);
nor U2250 (N_2250,N_2137,N_2131);
nand U2251 (N_2251,N_2148,N_2100);
and U2252 (N_2252,N_2143,N_2129);
xnor U2253 (N_2253,N_2135,N_2175);
nor U2254 (N_2254,N_2104,N_2173);
and U2255 (N_2255,N_2130,N_2158);
nand U2256 (N_2256,N_2167,N_2195);
nand U2257 (N_2257,N_2133,N_2154);
nor U2258 (N_2258,N_2122,N_2132);
and U2259 (N_2259,N_2104,N_2122);
nand U2260 (N_2260,N_2120,N_2115);
nor U2261 (N_2261,N_2158,N_2159);
nor U2262 (N_2262,N_2181,N_2123);
and U2263 (N_2263,N_2192,N_2113);
or U2264 (N_2264,N_2151,N_2137);
nand U2265 (N_2265,N_2102,N_2134);
nor U2266 (N_2266,N_2191,N_2111);
nor U2267 (N_2267,N_2116,N_2153);
or U2268 (N_2268,N_2142,N_2105);
nand U2269 (N_2269,N_2105,N_2131);
nor U2270 (N_2270,N_2186,N_2175);
or U2271 (N_2271,N_2184,N_2102);
or U2272 (N_2272,N_2194,N_2102);
nor U2273 (N_2273,N_2127,N_2163);
and U2274 (N_2274,N_2127,N_2168);
nand U2275 (N_2275,N_2128,N_2144);
nand U2276 (N_2276,N_2165,N_2104);
or U2277 (N_2277,N_2142,N_2197);
nand U2278 (N_2278,N_2180,N_2115);
and U2279 (N_2279,N_2155,N_2186);
or U2280 (N_2280,N_2184,N_2133);
and U2281 (N_2281,N_2188,N_2155);
or U2282 (N_2282,N_2100,N_2167);
nand U2283 (N_2283,N_2174,N_2171);
nor U2284 (N_2284,N_2187,N_2141);
xor U2285 (N_2285,N_2146,N_2137);
nor U2286 (N_2286,N_2147,N_2140);
nor U2287 (N_2287,N_2103,N_2189);
or U2288 (N_2288,N_2153,N_2162);
nand U2289 (N_2289,N_2193,N_2137);
xnor U2290 (N_2290,N_2145,N_2120);
xnor U2291 (N_2291,N_2154,N_2115);
and U2292 (N_2292,N_2142,N_2180);
or U2293 (N_2293,N_2148,N_2141);
nand U2294 (N_2294,N_2144,N_2195);
or U2295 (N_2295,N_2123,N_2136);
or U2296 (N_2296,N_2106,N_2118);
nand U2297 (N_2297,N_2103,N_2105);
and U2298 (N_2298,N_2149,N_2183);
xnor U2299 (N_2299,N_2192,N_2165);
and U2300 (N_2300,N_2237,N_2228);
nand U2301 (N_2301,N_2233,N_2272);
nor U2302 (N_2302,N_2202,N_2264);
nor U2303 (N_2303,N_2291,N_2238);
or U2304 (N_2304,N_2295,N_2222);
or U2305 (N_2305,N_2262,N_2288);
or U2306 (N_2306,N_2232,N_2277);
nor U2307 (N_2307,N_2253,N_2269);
or U2308 (N_2308,N_2281,N_2271);
nand U2309 (N_2309,N_2205,N_2275);
and U2310 (N_2310,N_2244,N_2284);
nor U2311 (N_2311,N_2259,N_2256);
nand U2312 (N_2312,N_2261,N_2212);
xnor U2313 (N_2313,N_2260,N_2219);
and U2314 (N_2314,N_2221,N_2246);
nand U2315 (N_2315,N_2251,N_2283);
or U2316 (N_2316,N_2289,N_2223);
and U2317 (N_2317,N_2294,N_2278);
and U2318 (N_2318,N_2287,N_2267);
and U2319 (N_2319,N_2257,N_2229);
nor U2320 (N_2320,N_2241,N_2210);
nand U2321 (N_2321,N_2225,N_2201);
or U2322 (N_2322,N_2245,N_2209);
nand U2323 (N_2323,N_2296,N_2274);
nor U2324 (N_2324,N_2206,N_2254);
nor U2325 (N_2325,N_2230,N_2208);
or U2326 (N_2326,N_2285,N_2200);
nand U2327 (N_2327,N_2236,N_2282);
or U2328 (N_2328,N_2293,N_2299);
and U2329 (N_2329,N_2276,N_2258);
or U2330 (N_2330,N_2250,N_2249);
or U2331 (N_2331,N_2231,N_2252);
xor U2332 (N_2332,N_2240,N_2297);
or U2333 (N_2333,N_2216,N_2211);
nor U2334 (N_2334,N_2217,N_2273);
nor U2335 (N_2335,N_2290,N_2204);
nand U2336 (N_2336,N_2242,N_2215);
or U2337 (N_2337,N_2270,N_2248);
nor U2338 (N_2338,N_2268,N_2234);
or U2339 (N_2339,N_2203,N_2207);
or U2340 (N_2340,N_2243,N_2214);
nand U2341 (N_2341,N_2224,N_2213);
and U2342 (N_2342,N_2218,N_2239);
nand U2343 (N_2343,N_2255,N_2298);
and U2344 (N_2344,N_2265,N_2279);
and U2345 (N_2345,N_2263,N_2227);
nor U2346 (N_2346,N_2220,N_2292);
nor U2347 (N_2347,N_2280,N_2247);
and U2348 (N_2348,N_2286,N_2235);
nand U2349 (N_2349,N_2226,N_2266);
nand U2350 (N_2350,N_2271,N_2260);
and U2351 (N_2351,N_2223,N_2216);
xor U2352 (N_2352,N_2243,N_2255);
nor U2353 (N_2353,N_2252,N_2265);
or U2354 (N_2354,N_2207,N_2205);
nor U2355 (N_2355,N_2262,N_2280);
and U2356 (N_2356,N_2255,N_2217);
or U2357 (N_2357,N_2211,N_2200);
or U2358 (N_2358,N_2255,N_2273);
nand U2359 (N_2359,N_2276,N_2264);
and U2360 (N_2360,N_2229,N_2295);
and U2361 (N_2361,N_2227,N_2291);
nand U2362 (N_2362,N_2210,N_2205);
nand U2363 (N_2363,N_2225,N_2280);
xnor U2364 (N_2364,N_2274,N_2205);
nor U2365 (N_2365,N_2214,N_2285);
nor U2366 (N_2366,N_2288,N_2233);
or U2367 (N_2367,N_2207,N_2217);
nor U2368 (N_2368,N_2262,N_2267);
nand U2369 (N_2369,N_2256,N_2293);
and U2370 (N_2370,N_2260,N_2224);
or U2371 (N_2371,N_2242,N_2264);
and U2372 (N_2372,N_2204,N_2205);
nand U2373 (N_2373,N_2261,N_2266);
or U2374 (N_2374,N_2200,N_2257);
and U2375 (N_2375,N_2265,N_2210);
or U2376 (N_2376,N_2296,N_2203);
and U2377 (N_2377,N_2252,N_2275);
nand U2378 (N_2378,N_2202,N_2275);
xor U2379 (N_2379,N_2210,N_2289);
nand U2380 (N_2380,N_2212,N_2283);
nand U2381 (N_2381,N_2215,N_2214);
nand U2382 (N_2382,N_2293,N_2228);
nand U2383 (N_2383,N_2231,N_2264);
nor U2384 (N_2384,N_2268,N_2215);
nand U2385 (N_2385,N_2263,N_2287);
and U2386 (N_2386,N_2229,N_2249);
and U2387 (N_2387,N_2225,N_2271);
and U2388 (N_2388,N_2216,N_2283);
and U2389 (N_2389,N_2200,N_2231);
or U2390 (N_2390,N_2205,N_2253);
nor U2391 (N_2391,N_2271,N_2276);
or U2392 (N_2392,N_2241,N_2288);
and U2393 (N_2393,N_2224,N_2293);
nor U2394 (N_2394,N_2218,N_2212);
nor U2395 (N_2395,N_2242,N_2214);
or U2396 (N_2396,N_2248,N_2272);
and U2397 (N_2397,N_2209,N_2265);
or U2398 (N_2398,N_2252,N_2290);
nor U2399 (N_2399,N_2229,N_2296);
or U2400 (N_2400,N_2339,N_2357);
nor U2401 (N_2401,N_2328,N_2336);
nor U2402 (N_2402,N_2378,N_2340);
or U2403 (N_2403,N_2377,N_2318);
or U2404 (N_2404,N_2366,N_2332);
nand U2405 (N_2405,N_2365,N_2394);
nand U2406 (N_2406,N_2362,N_2380);
xor U2407 (N_2407,N_2370,N_2313);
nand U2408 (N_2408,N_2363,N_2330);
or U2409 (N_2409,N_2345,N_2383);
and U2410 (N_2410,N_2312,N_2304);
nor U2411 (N_2411,N_2355,N_2309);
and U2412 (N_2412,N_2347,N_2342);
xnor U2413 (N_2413,N_2358,N_2335);
nor U2414 (N_2414,N_2371,N_2334);
nand U2415 (N_2415,N_2396,N_2361);
and U2416 (N_2416,N_2352,N_2386);
and U2417 (N_2417,N_2300,N_2399);
nand U2418 (N_2418,N_2301,N_2323);
xnor U2419 (N_2419,N_2325,N_2322);
or U2420 (N_2420,N_2368,N_2398);
nor U2421 (N_2421,N_2326,N_2395);
or U2422 (N_2422,N_2392,N_2319);
and U2423 (N_2423,N_2348,N_2364);
or U2424 (N_2424,N_2308,N_2373);
and U2425 (N_2425,N_2333,N_2344);
nor U2426 (N_2426,N_2350,N_2341);
nand U2427 (N_2427,N_2307,N_2317);
nor U2428 (N_2428,N_2353,N_2385);
nand U2429 (N_2429,N_2374,N_2388);
and U2430 (N_2430,N_2310,N_2349);
or U2431 (N_2431,N_2376,N_2359);
nand U2432 (N_2432,N_2321,N_2391);
nand U2433 (N_2433,N_2311,N_2303);
or U2434 (N_2434,N_2346,N_2327);
nor U2435 (N_2435,N_2381,N_2379);
and U2436 (N_2436,N_2329,N_2372);
or U2437 (N_2437,N_2324,N_2389);
nor U2438 (N_2438,N_2306,N_2302);
and U2439 (N_2439,N_2375,N_2351);
and U2440 (N_2440,N_2369,N_2356);
or U2441 (N_2441,N_2397,N_2354);
and U2442 (N_2442,N_2387,N_2360);
nor U2443 (N_2443,N_2314,N_2331);
or U2444 (N_2444,N_2384,N_2320);
nor U2445 (N_2445,N_2343,N_2305);
xnor U2446 (N_2446,N_2390,N_2382);
or U2447 (N_2447,N_2367,N_2337);
and U2448 (N_2448,N_2316,N_2393);
or U2449 (N_2449,N_2338,N_2315);
nand U2450 (N_2450,N_2309,N_2387);
nand U2451 (N_2451,N_2374,N_2330);
xor U2452 (N_2452,N_2336,N_2348);
nand U2453 (N_2453,N_2347,N_2312);
nor U2454 (N_2454,N_2384,N_2398);
nor U2455 (N_2455,N_2368,N_2301);
and U2456 (N_2456,N_2370,N_2388);
nor U2457 (N_2457,N_2341,N_2390);
or U2458 (N_2458,N_2380,N_2312);
or U2459 (N_2459,N_2338,N_2350);
or U2460 (N_2460,N_2390,N_2396);
and U2461 (N_2461,N_2314,N_2360);
or U2462 (N_2462,N_2361,N_2314);
and U2463 (N_2463,N_2315,N_2349);
or U2464 (N_2464,N_2353,N_2351);
nor U2465 (N_2465,N_2373,N_2394);
nor U2466 (N_2466,N_2330,N_2398);
nand U2467 (N_2467,N_2344,N_2331);
and U2468 (N_2468,N_2374,N_2323);
and U2469 (N_2469,N_2376,N_2319);
and U2470 (N_2470,N_2323,N_2353);
and U2471 (N_2471,N_2320,N_2337);
and U2472 (N_2472,N_2309,N_2314);
xor U2473 (N_2473,N_2366,N_2321);
nand U2474 (N_2474,N_2343,N_2306);
nand U2475 (N_2475,N_2315,N_2380);
nor U2476 (N_2476,N_2346,N_2365);
nand U2477 (N_2477,N_2385,N_2360);
nand U2478 (N_2478,N_2355,N_2328);
nor U2479 (N_2479,N_2351,N_2379);
nor U2480 (N_2480,N_2365,N_2388);
nor U2481 (N_2481,N_2382,N_2318);
nand U2482 (N_2482,N_2366,N_2339);
and U2483 (N_2483,N_2341,N_2352);
nor U2484 (N_2484,N_2373,N_2367);
and U2485 (N_2485,N_2362,N_2335);
nor U2486 (N_2486,N_2381,N_2315);
and U2487 (N_2487,N_2349,N_2319);
and U2488 (N_2488,N_2356,N_2351);
nor U2489 (N_2489,N_2307,N_2394);
and U2490 (N_2490,N_2388,N_2344);
and U2491 (N_2491,N_2361,N_2352);
nor U2492 (N_2492,N_2305,N_2347);
nor U2493 (N_2493,N_2354,N_2349);
nand U2494 (N_2494,N_2366,N_2345);
nor U2495 (N_2495,N_2303,N_2376);
and U2496 (N_2496,N_2369,N_2354);
or U2497 (N_2497,N_2314,N_2387);
and U2498 (N_2498,N_2392,N_2386);
xor U2499 (N_2499,N_2353,N_2375);
or U2500 (N_2500,N_2493,N_2415);
nand U2501 (N_2501,N_2401,N_2444);
nor U2502 (N_2502,N_2406,N_2432);
nand U2503 (N_2503,N_2498,N_2423);
or U2504 (N_2504,N_2484,N_2491);
nand U2505 (N_2505,N_2453,N_2428);
nand U2506 (N_2506,N_2430,N_2420);
xnor U2507 (N_2507,N_2457,N_2439);
nand U2508 (N_2508,N_2477,N_2476);
or U2509 (N_2509,N_2429,N_2467);
nor U2510 (N_2510,N_2487,N_2424);
nor U2511 (N_2511,N_2456,N_2495);
and U2512 (N_2512,N_2494,N_2416);
and U2513 (N_2513,N_2419,N_2460);
or U2514 (N_2514,N_2469,N_2400);
and U2515 (N_2515,N_2473,N_2440);
or U2516 (N_2516,N_2486,N_2417);
or U2517 (N_2517,N_2450,N_2402);
nand U2518 (N_2518,N_2418,N_2442);
nor U2519 (N_2519,N_2475,N_2431);
nand U2520 (N_2520,N_2449,N_2472);
nand U2521 (N_2521,N_2447,N_2451);
nand U2522 (N_2522,N_2426,N_2425);
or U2523 (N_2523,N_2421,N_2438);
nor U2524 (N_2524,N_2485,N_2483);
nor U2525 (N_2525,N_2403,N_2470);
and U2526 (N_2526,N_2448,N_2490);
nor U2527 (N_2527,N_2454,N_2412);
and U2528 (N_2528,N_2434,N_2408);
nand U2529 (N_2529,N_2465,N_2481);
nand U2530 (N_2530,N_2499,N_2488);
or U2531 (N_2531,N_2404,N_2455);
nand U2532 (N_2532,N_2443,N_2471);
xor U2533 (N_2533,N_2474,N_2405);
or U2534 (N_2534,N_2497,N_2496);
xor U2535 (N_2535,N_2414,N_2436);
and U2536 (N_2536,N_2479,N_2409);
or U2537 (N_2537,N_2445,N_2492);
nor U2538 (N_2538,N_2489,N_2435);
or U2539 (N_2539,N_2462,N_2452);
nand U2540 (N_2540,N_2480,N_2437);
or U2541 (N_2541,N_2463,N_2441);
nand U2542 (N_2542,N_2468,N_2422);
and U2543 (N_2543,N_2478,N_2413);
nor U2544 (N_2544,N_2427,N_2411);
and U2545 (N_2545,N_2410,N_2459);
nand U2546 (N_2546,N_2482,N_2458);
or U2547 (N_2547,N_2466,N_2446);
or U2548 (N_2548,N_2464,N_2461);
and U2549 (N_2549,N_2433,N_2407);
nand U2550 (N_2550,N_2476,N_2436);
nand U2551 (N_2551,N_2421,N_2493);
and U2552 (N_2552,N_2487,N_2416);
nand U2553 (N_2553,N_2486,N_2457);
or U2554 (N_2554,N_2419,N_2485);
nor U2555 (N_2555,N_2442,N_2484);
and U2556 (N_2556,N_2468,N_2418);
or U2557 (N_2557,N_2473,N_2441);
nor U2558 (N_2558,N_2410,N_2421);
nor U2559 (N_2559,N_2416,N_2438);
nand U2560 (N_2560,N_2422,N_2461);
and U2561 (N_2561,N_2473,N_2404);
nand U2562 (N_2562,N_2405,N_2469);
nor U2563 (N_2563,N_2428,N_2423);
nand U2564 (N_2564,N_2455,N_2498);
nor U2565 (N_2565,N_2476,N_2457);
nand U2566 (N_2566,N_2419,N_2482);
and U2567 (N_2567,N_2469,N_2481);
xor U2568 (N_2568,N_2477,N_2415);
nor U2569 (N_2569,N_2437,N_2448);
and U2570 (N_2570,N_2488,N_2456);
xnor U2571 (N_2571,N_2455,N_2440);
nor U2572 (N_2572,N_2453,N_2423);
nor U2573 (N_2573,N_2471,N_2423);
or U2574 (N_2574,N_2413,N_2421);
nand U2575 (N_2575,N_2422,N_2414);
and U2576 (N_2576,N_2459,N_2477);
nor U2577 (N_2577,N_2421,N_2476);
and U2578 (N_2578,N_2438,N_2456);
nand U2579 (N_2579,N_2487,N_2436);
and U2580 (N_2580,N_2498,N_2473);
nor U2581 (N_2581,N_2424,N_2455);
or U2582 (N_2582,N_2466,N_2402);
and U2583 (N_2583,N_2439,N_2443);
or U2584 (N_2584,N_2419,N_2496);
xnor U2585 (N_2585,N_2400,N_2445);
or U2586 (N_2586,N_2438,N_2457);
nor U2587 (N_2587,N_2402,N_2474);
and U2588 (N_2588,N_2435,N_2459);
nand U2589 (N_2589,N_2428,N_2433);
nor U2590 (N_2590,N_2450,N_2482);
nor U2591 (N_2591,N_2409,N_2463);
nand U2592 (N_2592,N_2472,N_2467);
nor U2593 (N_2593,N_2459,N_2461);
nand U2594 (N_2594,N_2441,N_2497);
xnor U2595 (N_2595,N_2499,N_2413);
xor U2596 (N_2596,N_2499,N_2480);
or U2597 (N_2597,N_2498,N_2483);
or U2598 (N_2598,N_2460,N_2476);
or U2599 (N_2599,N_2432,N_2494);
nand U2600 (N_2600,N_2500,N_2544);
nand U2601 (N_2601,N_2573,N_2553);
or U2602 (N_2602,N_2516,N_2503);
and U2603 (N_2603,N_2522,N_2576);
nor U2604 (N_2604,N_2588,N_2551);
xnor U2605 (N_2605,N_2552,N_2578);
or U2606 (N_2606,N_2547,N_2584);
nand U2607 (N_2607,N_2535,N_2558);
nand U2608 (N_2608,N_2579,N_2562);
nand U2609 (N_2609,N_2528,N_2507);
nor U2610 (N_2610,N_2564,N_2581);
and U2611 (N_2611,N_2533,N_2560);
and U2612 (N_2612,N_2574,N_2519);
and U2613 (N_2613,N_2523,N_2536);
and U2614 (N_2614,N_2571,N_2543);
nor U2615 (N_2615,N_2556,N_2572);
xnor U2616 (N_2616,N_2510,N_2525);
nand U2617 (N_2617,N_2549,N_2591);
nand U2618 (N_2618,N_2597,N_2502);
nor U2619 (N_2619,N_2540,N_2546);
nor U2620 (N_2620,N_2598,N_2587);
or U2621 (N_2621,N_2563,N_2529);
nand U2622 (N_2622,N_2582,N_2534);
and U2623 (N_2623,N_2555,N_2583);
nor U2624 (N_2624,N_2569,N_2520);
and U2625 (N_2625,N_2538,N_2570);
or U2626 (N_2626,N_2514,N_2593);
nand U2627 (N_2627,N_2565,N_2511);
nor U2628 (N_2628,N_2537,N_2589);
and U2629 (N_2629,N_2577,N_2580);
nand U2630 (N_2630,N_2513,N_2517);
nand U2631 (N_2631,N_2590,N_2531);
nand U2632 (N_2632,N_2521,N_2561);
nand U2633 (N_2633,N_2585,N_2515);
nand U2634 (N_2634,N_2548,N_2509);
nor U2635 (N_2635,N_2527,N_2539);
nor U2636 (N_2636,N_2596,N_2504);
nor U2637 (N_2637,N_2501,N_2541);
xor U2638 (N_2638,N_2575,N_2592);
nor U2639 (N_2639,N_2586,N_2568);
or U2640 (N_2640,N_2599,N_2508);
nand U2641 (N_2641,N_2506,N_2594);
and U2642 (N_2642,N_2567,N_2545);
and U2643 (N_2643,N_2554,N_2550);
and U2644 (N_2644,N_2530,N_2518);
nor U2645 (N_2645,N_2559,N_2557);
nand U2646 (N_2646,N_2566,N_2524);
xnor U2647 (N_2647,N_2542,N_2526);
nor U2648 (N_2648,N_2505,N_2512);
or U2649 (N_2649,N_2532,N_2595);
or U2650 (N_2650,N_2581,N_2574);
and U2651 (N_2651,N_2572,N_2533);
nor U2652 (N_2652,N_2522,N_2549);
nand U2653 (N_2653,N_2521,N_2540);
nor U2654 (N_2654,N_2534,N_2510);
xnor U2655 (N_2655,N_2528,N_2529);
nand U2656 (N_2656,N_2584,N_2582);
nor U2657 (N_2657,N_2503,N_2502);
nand U2658 (N_2658,N_2538,N_2572);
and U2659 (N_2659,N_2512,N_2521);
nand U2660 (N_2660,N_2588,N_2576);
nand U2661 (N_2661,N_2544,N_2505);
nand U2662 (N_2662,N_2534,N_2512);
nor U2663 (N_2663,N_2577,N_2506);
nand U2664 (N_2664,N_2583,N_2598);
or U2665 (N_2665,N_2563,N_2562);
and U2666 (N_2666,N_2573,N_2510);
nor U2667 (N_2667,N_2557,N_2554);
nor U2668 (N_2668,N_2560,N_2516);
nand U2669 (N_2669,N_2552,N_2569);
nor U2670 (N_2670,N_2574,N_2568);
or U2671 (N_2671,N_2508,N_2521);
and U2672 (N_2672,N_2579,N_2599);
nor U2673 (N_2673,N_2552,N_2535);
and U2674 (N_2674,N_2543,N_2562);
or U2675 (N_2675,N_2518,N_2535);
or U2676 (N_2676,N_2578,N_2573);
or U2677 (N_2677,N_2542,N_2509);
nand U2678 (N_2678,N_2519,N_2536);
nand U2679 (N_2679,N_2516,N_2579);
nor U2680 (N_2680,N_2562,N_2559);
or U2681 (N_2681,N_2575,N_2506);
nor U2682 (N_2682,N_2501,N_2519);
nand U2683 (N_2683,N_2589,N_2516);
nor U2684 (N_2684,N_2521,N_2545);
or U2685 (N_2685,N_2514,N_2582);
nor U2686 (N_2686,N_2513,N_2504);
nor U2687 (N_2687,N_2566,N_2532);
or U2688 (N_2688,N_2583,N_2514);
or U2689 (N_2689,N_2564,N_2548);
nand U2690 (N_2690,N_2557,N_2502);
xnor U2691 (N_2691,N_2549,N_2532);
nor U2692 (N_2692,N_2576,N_2584);
nor U2693 (N_2693,N_2579,N_2534);
and U2694 (N_2694,N_2514,N_2568);
nor U2695 (N_2695,N_2525,N_2595);
nand U2696 (N_2696,N_2521,N_2505);
nand U2697 (N_2697,N_2548,N_2591);
nand U2698 (N_2698,N_2593,N_2528);
or U2699 (N_2699,N_2594,N_2584);
nor U2700 (N_2700,N_2633,N_2682);
nor U2701 (N_2701,N_2638,N_2617);
or U2702 (N_2702,N_2663,N_2666);
nand U2703 (N_2703,N_2621,N_2680);
nand U2704 (N_2704,N_2695,N_2688);
and U2705 (N_2705,N_2643,N_2620);
and U2706 (N_2706,N_2676,N_2694);
nand U2707 (N_2707,N_2644,N_2619);
and U2708 (N_2708,N_2684,N_2679);
nand U2709 (N_2709,N_2685,N_2665);
or U2710 (N_2710,N_2626,N_2634);
and U2711 (N_2711,N_2611,N_2689);
or U2712 (N_2712,N_2603,N_2645);
xor U2713 (N_2713,N_2647,N_2683);
or U2714 (N_2714,N_2613,N_2678);
and U2715 (N_2715,N_2631,N_2655);
nand U2716 (N_2716,N_2636,N_2653);
and U2717 (N_2717,N_2609,N_2654);
and U2718 (N_2718,N_2693,N_2601);
or U2719 (N_2719,N_2607,N_2615);
or U2720 (N_2720,N_2616,N_2691);
nor U2721 (N_2721,N_2670,N_2681);
nand U2722 (N_2722,N_2632,N_2664);
or U2723 (N_2723,N_2629,N_2657);
nor U2724 (N_2724,N_2672,N_2635);
nor U2725 (N_2725,N_2651,N_2630);
nor U2726 (N_2726,N_2659,N_2612);
nor U2727 (N_2727,N_2618,N_2667);
or U2728 (N_2728,N_2692,N_2686);
and U2729 (N_2729,N_2677,N_2646);
nand U2730 (N_2730,N_2641,N_2602);
nand U2731 (N_2731,N_2639,N_2669);
and U2732 (N_2732,N_2660,N_2698);
nor U2733 (N_2733,N_2637,N_2627);
nand U2734 (N_2734,N_2608,N_2696);
and U2735 (N_2735,N_2642,N_2656);
and U2736 (N_2736,N_2640,N_2697);
nor U2737 (N_2737,N_2662,N_2623);
nor U2738 (N_2738,N_2674,N_2625);
xnor U2739 (N_2739,N_2604,N_2610);
nor U2740 (N_2740,N_2605,N_2614);
and U2741 (N_2741,N_2652,N_2649);
nor U2742 (N_2742,N_2661,N_2687);
or U2743 (N_2743,N_2600,N_2622);
and U2744 (N_2744,N_2671,N_2675);
or U2745 (N_2745,N_2648,N_2673);
nand U2746 (N_2746,N_2650,N_2606);
or U2747 (N_2747,N_2624,N_2658);
and U2748 (N_2748,N_2628,N_2699);
nand U2749 (N_2749,N_2668,N_2690);
xnor U2750 (N_2750,N_2620,N_2699);
or U2751 (N_2751,N_2698,N_2606);
xnor U2752 (N_2752,N_2680,N_2682);
nor U2753 (N_2753,N_2656,N_2602);
or U2754 (N_2754,N_2653,N_2606);
nand U2755 (N_2755,N_2619,N_2696);
nand U2756 (N_2756,N_2647,N_2603);
or U2757 (N_2757,N_2635,N_2684);
and U2758 (N_2758,N_2682,N_2660);
nand U2759 (N_2759,N_2635,N_2607);
nand U2760 (N_2760,N_2694,N_2629);
nand U2761 (N_2761,N_2614,N_2613);
nand U2762 (N_2762,N_2630,N_2631);
and U2763 (N_2763,N_2661,N_2641);
nand U2764 (N_2764,N_2637,N_2661);
and U2765 (N_2765,N_2620,N_2625);
nor U2766 (N_2766,N_2621,N_2632);
nand U2767 (N_2767,N_2634,N_2693);
and U2768 (N_2768,N_2628,N_2679);
and U2769 (N_2769,N_2675,N_2683);
nor U2770 (N_2770,N_2611,N_2655);
nor U2771 (N_2771,N_2688,N_2602);
nand U2772 (N_2772,N_2640,N_2664);
nor U2773 (N_2773,N_2689,N_2617);
and U2774 (N_2774,N_2657,N_2638);
nor U2775 (N_2775,N_2608,N_2639);
nand U2776 (N_2776,N_2664,N_2645);
and U2777 (N_2777,N_2652,N_2665);
or U2778 (N_2778,N_2698,N_2640);
and U2779 (N_2779,N_2632,N_2691);
and U2780 (N_2780,N_2651,N_2646);
and U2781 (N_2781,N_2670,N_2656);
or U2782 (N_2782,N_2654,N_2663);
or U2783 (N_2783,N_2682,N_2624);
xor U2784 (N_2784,N_2605,N_2672);
or U2785 (N_2785,N_2633,N_2696);
nand U2786 (N_2786,N_2643,N_2624);
nand U2787 (N_2787,N_2609,N_2621);
or U2788 (N_2788,N_2640,N_2635);
nor U2789 (N_2789,N_2627,N_2654);
nor U2790 (N_2790,N_2638,N_2680);
xor U2791 (N_2791,N_2605,N_2600);
nor U2792 (N_2792,N_2647,N_2622);
nand U2793 (N_2793,N_2696,N_2614);
and U2794 (N_2794,N_2613,N_2642);
or U2795 (N_2795,N_2660,N_2648);
nand U2796 (N_2796,N_2610,N_2627);
or U2797 (N_2797,N_2667,N_2603);
nor U2798 (N_2798,N_2624,N_2625);
nor U2799 (N_2799,N_2612,N_2618);
nor U2800 (N_2800,N_2785,N_2755);
nand U2801 (N_2801,N_2712,N_2765);
nand U2802 (N_2802,N_2735,N_2789);
nor U2803 (N_2803,N_2705,N_2749);
and U2804 (N_2804,N_2788,N_2714);
nor U2805 (N_2805,N_2798,N_2731);
xor U2806 (N_2806,N_2767,N_2776);
and U2807 (N_2807,N_2784,N_2752);
or U2808 (N_2808,N_2710,N_2723);
and U2809 (N_2809,N_2758,N_2780);
and U2810 (N_2810,N_2783,N_2737);
xor U2811 (N_2811,N_2732,N_2774);
and U2812 (N_2812,N_2702,N_2721);
or U2813 (N_2813,N_2704,N_2738);
and U2814 (N_2814,N_2762,N_2716);
and U2815 (N_2815,N_2787,N_2799);
nand U2816 (N_2816,N_2742,N_2761);
nand U2817 (N_2817,N_2756,N_2779);
nand U2818 (N_2818,N_2764,N_2791);
or U2819 (N_2819,N_2718,N_2782);
or U2820 (N_2820,N_2744,N_2769);
nor U2821 (N_2821,N_2720,N_2778);
and U2822 (N_2822,N_2707,N_2727);
and U2823 (N_2823,N_2773,N_2701);
nor U2824 (N_2824,N_2709,N_2760);
nand U2825 (N_2825,N_2708,N_2713);
xor U2826 (N_2826,N_2703,N_2757);
and U2827 (N_2827,N_2729,N_2763);
or U2828 (N_2828,N_2795,N_2711);
xor U2829 (N_2829,N_2794,N_2777);
and U2830 (N_2830,N_2747,N_2796);
and U2831 (N_2831,N_2786,N_2754);
xor U2832 (N_2832,N_2740,N_2724);
and U2833 (N_2833,N_2700,N_2745);
and U2834 (N_2834,N_2730,N_2775);
and U2835 (N_2835,N_2728,N_2741);
or U2836 (N_2836,N_2793,N_2750);
or U2837 (N_2837,N_2751,N_2743);
and U2838 (N_2838,N_2768,N_2748);
xor U2839 (N_2839,N_2736,N_2766);
nand U2840 (N_2840,N_2722,N_2706);
xnor U2841 (N_2841,N_2781,N_2746);
and U2842 (N_2842,N_2797,N_2725);
or U2843 (N_2843,N_2771,N_2753);
nor U2844 (N_2844,N_2759,N_2726);
and U2845 (N_2845,N_2790,N_2772);
nand U2846 (N_2846,N_2734,N_2770);
nor U2847 (N_2847,N_2739,N_2719);
and U2848 (N_2848,N_2715,N_2792);
or U2849 (N_2849,N_2733,N_2717);
xnor U2850 (N_2850,N_2708,N_2795);
nor U2851 (N_2851,N_2763,N_2760);
xnor U2852 (N_2852,N_2769,N_2775);
xor U2853 (N_2853,N_2700,N_2729);
nor U2854 (N_2854,N_2762,N_2775);
nor U2855 (N_2855,N_2756,N_2718);
nor U2856 (N_2856,N_2727,N_2792);
nor U2857 (N_2857,N_2712,N_2753);
or U2858 (N_2858,N_2734,N_2786);
or U2859 (N_2859,N_2727,N_2760);
or U2860 (N_2860,N_2733,N_2734);
or U2861 (N_2861,N_2793,N_2748);
nor U2862 (N_2862,N_2782,N_2716);
and U2863 (N_2863,N_2746,N_2716);
nand U2864 (N_2864,N_2754,N_2743);
nand U2865 (N_2865,N_2717,N_2705);
or U2866 (N_2866,N_2768,N_2773);
nor U2867 (N_2867,N_2793,N_2738);
nand U2868 (N_2868,N_2750,N_2753);
nand U2869 (N_2869,N_2752,N_2719);
nand U2870 (N_2870,N_2754,N_2768);
nor U2871 (N_2871,N_2730,N_2798);
nor U2872 (N_2872,N_2714,N_2701);
or U2873 (N_2873,N_2757,N_2764);
or U2874 (N_2874,N_2710,N_2724);
nand U2875 (N_2875,N_2734,N_2747);
or U2876 (N_2876,N_2785,N_2727);
or U2877 (N_2877,N_2702,N_2755);
nor U2878 (N_2878,N_2709,N_2784);
or U2879 (N_2879,N_2765,N_2741);
nor U2880 (N_2880,N_2784,N_2767);
nor U2881 (N_2881,N_2775,N_2783);
and U2882 (N_2882,N_2747,N_2730);
nand U2883 (N_2883,N_2777,N_2769);
or U2884 (N_2884,N_2747,N_2703);
and U2885 (N_2885,N_2797,N_2772);
nand U2886 (N_2886,N_2749,N_2701);
nand U2887 (N_2887,N_2784,N_2798);
nor U2888 (N_2888,N_2705,N_2723);
xnor U2889 (N_2889,N_2752,N_2739);
nor U2890 (N_2890,N_2733,N_2745);
xor U2891 (N_2891,N_2709,N_2775);
or U2892 (N_2892,N_2776,N_2725);
nor U2893 (N_2893,N_2742,N_2707);
xnor U2894 (N_2894,N_2761,N_2719);
or U2895 (N_2895,N_2746,N_2793);
nor U2896 (N_2896,N_2708,N_2797);
nand U2897 (N_2897,N_2790,N_2708);
nand U2898 (N_2898,N_2776,N_2748);
or U2899 (N_2899,N_2718,N_2724);
nand U2900 (N_2900,N_2869,N_2800);
nor U2901 (N_2901,N_2865,N_2830);
nand U2902 (N_2902,N_2841,N_2884);
nor U2903 (N_2903,N_2881,N_2870);
and U2904 (N_2904,N_2879,N_2883);
nor U2905 (N_2905,N_2840,N_2896);
and U2906 (N_2906,N_2878,N_2859);
nor U2907 (N_2907,N_2872,N_2860);
nand U2908 (N_2908,N_2834,N_2816);
nand U2909 (N_2909,N_2864,N_2867);
nor U2910 (N_2910,N_2863,N_2802);
and U2911 (N_2911,N_2852,N_2853);
or U2912 (N_2912,N_2871,N_2805);
and U2913 (N_2913,N_2846,N_2838);
nand U2914 (N_2914,N_2845,N_2803);
nand U2915 (N_2915,N_2831,N_2877);
and U2916 (N_2916,N_2837,N_2857);
or U2917 (N_2917,N_2880,N_2829);
and U2918 (N_2918,N_2849,N_2855);
and U2919 (N_2919,N_2839,N_2894);
nor U2920 (N_2920,N_2836,N_2873);
or U2921 (N_2921,N_2827,N_2843);
or U2922 (N_2922,N_2807,N_2804);
and U2923 (N_2923,N_2888,N_2850);
or U2924 (N_2924,N_2817,N_2856);
nand U2925 (N_2925,N_2893,N_2828);
nor U2926 (N_2926,N_2825,N_2874);
nand U2927 (N_2927,N_2897,N_2861);
nand U2928 (N_2928,N_2833,N_2842);
or U2929 (N_2929,N_2875,N_2882);
nor U2930 (N_2930,N_2887,N_2847);
xor U2931 (N_2931,N_2818,N_2806);
nor U2932 (N_2932,N_2826,N_2811);
nor U2933 (N_2933,N_2851,N_2823);
nor U2934 (N_2934,N_2862,N_2814);
and U2935 (N_2935,N_2810,N_2899);
and U2936 (N_2936,N_2892,N_2808);
or U2937 (N_2937,N_2858,N_2885);
xor U2938 (N_2938,N_2898,N_2889);
and U2939 (N_2939,N_2891,N_2832);
and U2940 (N_2940,N_2815,N_2835);
nand U2941 (N_2941,N_2868,N_2876);
or U2942 (N_2942,N_2801,N_2819);
nand U2943 (N_2943,N_2809,N_2895);
nand U2944 (N_2944,N_2886,N_2866);
nand U2945 (N_2945,N_2822,N_2820);
xnor U2946 (N_2946,N_2844,N_2890);
xor U2947 (N_2947,N_2854,N_2824);
nor U2948 (N_2948,N_2821,N_2812);
or U2949 (N_2949,N_2813,N_2848);
nor U2950 (N_2950,N_2836,N_2880);
and U2951 (N_2951,N_2812,N_2809);
nor U2952 (N_2952,N_2859,N_2850);
or U2953 (N_2953,N_2832,N_2864);
xnor U2954 (N_2954,N_2814,N_2877);
nand U2955 (N_2955,N_2805,N_2880);
and U2956 (N_2956,N_2894,N_2800);
or U2957 (N_2957,N_2812,N_2899);
nand U2958 (N_2958,N_2815,N_2822);
nand U2959 (N_2959,N_2876,N_2824);
nand U2960 (N_2960,N_2846,N_2857);
xor U2961 (N_2961,N_2802,N_2805);
and U2962 (N_2962,N_2879,N_2895);
nor U2963 (N_2963,N_2801,N_2811);
or U2964 (N_2964,N_2849,N_2890);
nand U2965 (N_2965,N_2877,N_2857);
nor U2966 (N_2966,N_2816,N_2868);
nand U2967 (N_2967,N_2887,N_2892);
xnor U2968 (N_2968,N_2803,N_2813);
nand U2969 (N_2969,N_2822,N_2892);
and U2970 (N_2970,N_2866,N_2840);
nand U2971 (N_2971,N_2847,N_2846);
xnor U2972 (N_2972,N_2858,N_2854);
or U2973 (N_2973,N_2888,N_2824);
xnor U2974 (N_2974,N_2839,N_2808);
xnor U2975 (N_2975,N_2873,N_2867);
or U2976 (N_2976,N_2826,N_2874);
nor U2977 (N_2977,N_2826,N_2890);
or U2978 (N_2978,N_2866,N_2873);
and U2979 (N_2979,N_2857,N_2859);
or U2980 (N_2980,N_2861,N_2804);
or U2981 (N_2981,N_2850,N_2817);
nor U2982 (N_2982,N_2853,N_2888);
and U2983 (N_2983,N_2827,N_2838);
nor U2984 (N_2984,N_2880,N_2888);
nand U2985 (N_2985,N_2832,N_2833);
nand U2986 (N_2986,N_2881,N_2852);
or U2987 (N_2987,N_2834,N_2800);
nor U2988 (N_2988,N_2867,N_2821);
nand U2989 (N_2989,N_2848,N_2823);
and U2990 (N_2990,N_2802,N_2835);
xor U2991 (N_2991,N_2889,N_2816);
nand U2992 (N_2992,N_2877,N_2895);
nand U2993 (N_2993,N_2866,N_2800);
and U2994 (N_2994,N_2837,N_2899);
nor U2995 (N_2995,N_2897,N_2888);
nor U2996 (N_2996,N_2884,N_2861);
nor U2997 (N_2997,N_2869,N_2858);
nor U2998 (N_2998,N_2849,N_2820);
nor U2999 (N_2999,N_2856,N_2891);
xnor U3000 (N_3000,N_2947,N_2930);
nand U3001 (N_3001,N_2996,N_2986);
or U3002 (N_3002,N_2962,N_2923);
and U3003 (N_3003,N_2942,N_2965);
nand U3004 (N_3004,N_2926,N_2939);
nor U3005 (N_3005,N_2963,N_2929);
xnor U3006 (N_3006,N_2975,N_2989);
nor U3007 (N_3007,N_2924,N_2950);
or U3008 (N_3008,N_2901,N_2938);
or U3009 (N_3009,N_2976,N_2957);
or U3010 (N_3010,N_2952,N_2928);
nor U3011 (N_3011,N_2945,N_2980);
nor U3012 (N_3012,N_2921,N_2967);
or U3013 (N_3013,N_2964,N_2933);
or U3014 (N_3014,N_2994,N_2993);
or U3015 (N_3015,N_2982,N_2912);
nand U3016 (N_3016,N_2934,N_2927);
or U3017 (N_3017,N_2988,N_2978);
nor U3018 (N_3018,N_2999,N_2913);
nor U3019 (N_3019,N_2997,N_2958);
and U3020 (N_3020,N_2949,N_2944);
and U3021 (N_3021,N_2948,N_2992);
nor U3022 (N_3022,N_2900,N_2911);
or U3023 (N_3023,N_2940,N_2931);
or U3024 (N_3024,N_2932,N_2907);
or U3025 (N_3025,N_2920,N_2995);
and U3026 (N_3026,N_2935,N_2916);
or U3027 (N_3027,N_2943,N_2904);
nand U3028 (N_3028,N_2968,N_2998);
nand U3029 (N_3029,N_2903,N_2936);
xor U3030 (N_3030,N_2981,N_2984);
nor U3031 (N_3031,N_2979,N_2953);
and U3032 (N_3032,N_2971,N_2917);
and U3033 (N_3033,N_2960,N_2987);
nand U3034 (N_3034,N_2905,N_2910);
nor U3035 (N_3035,N_2941,N_2966);
nor U3036 (N_3036,N_2970,N_2946);
and U3037 (N_3037,N_2918,N_2955);
or U3038 (N_3038,N_2991,N_2990);
and U3039 (N_3039,N_2909,N_2961);
nor U3040 (N_3040,N_2902,N_2959);
nor U3041 (N_3041,N_2954,N_2983);
xnor U3042 (N_3042,N_2956,N_2937);
nor U3043 (N_3043,N_2914,N_2972);
or U3044 (N_3044,N_2969,N_2973);
xnor U3045 (N_3045,N_2985,N_2919);
nand U3046 (N_3046,N_2925,N_2915);
nor U3047 (N_3047,N_2974,N_2922);
xnor U3048 (N_3048,N_2951,N_2908);
xnor U3049 (N_3049,N_2906,N_2977);
or U3050 (N_3050,N_2937,N_2965);
and U3051 (N_3051,N_2904,N_2936);
and U3052 (N_3052,N_2992,N_2972);
nand U3053 (N_3053,N_2948,N_2943);
nor U3054 (N_3054,N_2966,N_2949);
nor U3055 (N_3055,N_2943,N_2954);
nor U3056 (N_3056,N_2902,N_2980);
nand U3057 (N_3057,N_2922,N_2930);
nor U3058 (N_3058,N_2994,N_2931);
nor U3059 (N_3059,N_2988,N_2906);
or U3060 (N_3060,N_2912,N_2946);
or U3061 (N_3061,N_2989,N_2945);
or U3062 (N_3062,N_2960,N_2967);
nand U3063 (N_3063,N_2924,N_2917);
nand U3064 (N_3064,N_2928,N_2957);
nor U3065 (N_3065,N_2935,N_2956);
and U3066 (N_3066,N_2921,N_2925);
nor U3067 (N_3067,N_2962,N_2991);
or U3068 (N_3068,N_2923,N_2950);
xnor U3069 (N_3069,N_2983,N_2924);
or U3070 (N_3070,N_2906,N_2974);
or U3071 (N_3071,N_2907,N_2955);
nor U3072 (N_3072,N_2935,N_2965);
or U3073 (N_3073,N_2985,N_2925);
and U3074 (N_3074,N_2950,N_2994);
xnor U3075 (N_3075,N_2927,N_2993);
or U3076 (N_3076,N_2979,N_2943);
nor U3077 (N_3077,N_2967,N_2997);
or U3078 (N_3078,N_2996,N_2920);
nand U3079 (N_3079,N_2995,N_2935);
and U3080 (N_3080,N_2951,N_2967);
or U3081 (N_3081,N_2907,N_2964);
xor U3082 (N_3082,N_2933,N_2939);
nor U3083 (N_3083,N_2995,N_2979);
or U3084 (N_3084,N_2936,N_2954);
nand U3085 (N_3085,N_2959,N_2990);
nand U3086 (N_3086,N_2945,N_2919);
nor U3087 (N_3087,N_2977,N_2974);
and U3088 (N_3088,N_2957,N_2915);
or U3089 (N_3089,N_2904,N_2965);
nand U3090 (N_3090,N_2970,N_2922);
or U3091 (N_3091,N_2928,N_2962);
nor U3092 (N_3092,N_2978,N_2920);
nor U3093 (N_3093,N_2944,N_2988);
nand U3094 (N_3094,N_2900,N_2985);
or U3095 (N_3095,N_2900,N_2953);
nor U3096 (N_3096,N_2968,N_2952);
xnor U3097 (N_3097,N_2952,N_2974);
or U3098 (N_3098,N_2922,N_2931);
and U3099 (N_3099,N_2948,N_2962);
and U3100 (N_3100,N_3049,N_3035);
and U3101 (N_3101,N_3086,N_3057);
nand U3102 (N_3102,N_3091,N_3017);
xnor U3103 (N_3103,N_3077,N_3081);
nand U3104 (N_3104,N_3093,N_3039);
nor U3105 (N_3105,N_3090,N_3084);
and U3106 (N_3106,N_3046,N_3011);
and U3107 (N_3107,N_3016,N_3094);
nor U3108 (N_3108,N_3003,N_3031);
and U3109 (N_3109,N_3002,N_3079);
or U3110 (N_3110,N_3092,N_3082);
or U3111 (N_3111,N_3010,N_3099);
and U3112 (N_3112,N_3063,N_3000);
nand U3113 (N_3113,N_3040,N_3051);
nand U3114 (N_3114,N_3018,N_3020);
and U3115 (N_3115,N_3050,N_3068);
nor U3116 (N_3116,N_3043,N_3048);
nor U3117 (N_3117,N_3088,N_3062);
nor U3118 (N_3118,N_3041,N_3034);
or U3119 (N_3119,N_3023,N_3076);
or U3120 (N_3120,N_3095,N_3075);
nor U3121 (N_3121,N_3004,N_3059);
nand U3122 (N_3122,N_3074,N_3025);
xnor U3123 (N_3123,N_3089,N_3058);
or U3124 (N_3124,N_3044,N_3080);
nand U3125 (N_3125,N_3061,N_3085);
nor U3126 (N_3126,N_3045,N_3047);
nand U3127 (N_3127,N_3054,N_3012);
or U3128 (N_3128,N_3064,N_3069);
and U3129 (N_3129,N_3026,N_3042);
nor U3130 (N_3130,N_3070,N_3007);
nor U3131 (N_3131,N_3053,N_3037);
nor U3132 (N_3132,N_3028,N_3005);
or U3133 (N_3133,N_3032,N_3067);
and U3134 (N_3134,N_3072,N_3060);
nor U3135 (N_3135,N_3019,N_3027);
nand U3136 (N_3136,N_3097,N_3001);
xor U3137 (N_3137,N_3056,N_3015);
or U3138 (N_3138,N_3065,N_3055);
nor U3139 (N_3139,N_3008,N_3024);
nor U3140 (N_3140,N_3014,N_3087);
nor U3141 (N_3141,N_3078,N_3036);
nor U3142 (N_3142,N_3052,N_3083);
nor U3143 (N_3143,N_3021,N_3038);
nand U3144 (N_3144,N_3022,N_3029);
nor U3145 (N_3145,N_3030,N_3009);
nor U3146 (N_3146,N_3096,N_3071);
and U3147 (N_3147,N_3066,N_3033);
nor U3148 (N_3148,N_3073,N_3098);
or U3149 (N_3149,N_3013,N_3006);
nand U3150 (N_3150,N_3073,N_3059);
and U3151 (N_3151,N_3065,N_3072);
nor U3152 (N_3152,N_3035,N_3033);
and U3153 (N_3153,N_3041,N_3039);
or U3154 (N_3154,N_3020,N_3034);
nand U3155 (N_3155,N_3097,N_3056);
or U3156 (N_3156,N_3002,N_3058);
nand U3157 (N_3157,N_3031,N_3045);
nor U3158 (N_3158,N_3013,N_3070);
nor U3159 (N_3159,N_3044,N_3082);
or U3160 (N_3160,N_3093,N_3058);
xnor U3161 (N_3161,N_3014,N_3057);
nor U3162 (N_3162,N_3004,N_3007);
and U3163 (N_3163,N_3095,N_3050);
nor U3164 (N_3164,N_3081,N_3038);
nor U3165 (N_3165,N_3078,N_3032);
or U3166 (N_3166,N_3080,N_3058);
and U3167 (N_3167,N_3070,N_3022);
xor U3168 (N_3168,N_3057,N_3019);
or U3169 (N_3169,N_3088,N_3002);
nor U3170 (N_3170,N_3091,N_3012);
or U3171 (N_3171,N_3075,N_3048);
and U3172 (N_3172,N_3036,N_3069);
nor U3173 (N_3173,N_3001,N_3044);
or U3174 (N_3174,N_3083,N_3089);
xnor U3175 (N_3175,N_3085,N_3086);
xnor U3176 (N_3176,N_3056,N_3090);
nor U3177 (N_3177,N_3061,N_3036);
and U3178 (N_3178,N_3077,N_3072);
nor U3179 (N_3179,N_3028,N_3067);
or U3180 (N_3180,N_3057,N_3081);
nor U3181 (N_3181,N_3015,N_3032);
or U3182 (N_3182,N_3047,N_3052);
nand U3183 (N_3183,N_3044,N_3038);
and U3184 (N_3184,N_3040,N_3008);
nor U3185 (N_3185,N_3098,N_3056);
or U3186 (N_3186,N_3039,N_3070);
and U3187 (N_3187,N_3095,N_3014);
nor U3188 (N_3188,N_3047,N_3040);
nand U3189 (N_3189,N_3073,N_3075);
or U3190 (N_3190,N_3094,N_3010);
nand U3191 (N_3191,N_3070,N_3064);
nand U3192 (N_3192,N_3077,N_3099);
and U3193 (N_3193,N_3045,N_3098);
xor U3194 (N_3194,N_3097,N_3092);
and U3195 (N_3195,N_3090,N_3051);
nand U3196 (N_3196,N_3005,N_3052);
or U3197 (N_3197,N_3059,N_3054);
nand U3198 (N_3198,N_3002,N_3030);
nand U3199 (N_3199,N_3052,N_3040);
and U3200 (N_3200,N_3189,N_3143);
and U3201 (N_3201,N_3145,N_3107);
or U3202 (N_3202,N_3114,N_3121);
xor U3203 (N_3203,N_3177,N_3169);
or U3204 (N_3204,N_3105,N_3112);
nand U3205 (N_3205,N_3125,N_3150);
nand U3206 (N_3206,N_3162,N_3106);
xnor U3207 (N_3207,N_3135,N_3149);
or U3208 (N_3208,N_3140,N_3156);
and U3209 (N_3209,N_3110,N_3128);
nor U3210 (N_3210,N_3144,N_3136);
or U3211 (N_3211,N_3153,N_3183);
or U3212 (N_3212,N_3100,N_3115);
or U3213 (N_3213,N_3101,N_3141);
nor U3214 (N_3214,N_3160,N_3194);
or U3215 (N_3215,N_3157,N_3134);
nand U3216 (N_3216,N_3111,N_3198);
and U3217 (N_3217,N_3196,N_3127);
and U3218 (N_3218,N_3137,N_3129);
and U3219 (N_3219,N_3124,N_3132);
nor U3220 (N_3220,N_3199,N_3185);
nor U3221 (N_3221,N_3123,N_3188);
and U3222 (N_3222,N_3113,N_3155);
nor U3223 (N_3223,N_3159,N_3116);
nand U3224 (N_3224,N_3138,N_3171);
nand U3225 (N_3225,N_3118,N_3191);
and U3226 (N_3226,N_3192,N_3130);
nor U3227 (N_3227,N_3180,N_3102);
and U3228 (N_3228,N_3152,N_3186);
and U3229 (N_3229,N_3120,N_3104);
nand U3230 (N_3230,N_3146,N_3163);
nor U3231 (N_3231,N_3176,N_3154);
nor U3232 (N_3232,N_3195,N_3109);
xnor U3233 (N_3233,N_3197,N_3167);
xnor U3234 (N_3234,N_3158,N_3166);
or U3235 (N_3235,N_3103,N_3117);
nor U3236 (N_3236,N_3182,N_3190);
nor U3237 (N_3237,N_3181,N_3168);
xor U3238 (N_3238,N_3131,N_3108);
or U3239 (N_3239,N_3175,N_3133);
and U3240 (N_3240,N_3126,N_3142);
nand U3241 (N_3241,N_3174,N_3184);
or U3242 (N_3242,N_3170,N_3187);
nand U3243 (N_3243,N_3122,N_3139);
nor U3244 (N_3244,N_3119,N_3173);
and U3245 (N_3245,N_3161,N_3148);
nand U3246 (N_3246,N_3164,N_3193);
or U3247 (N_3247,N_3172,N_3178);
or U3248 (N_3248,N_3179,N_3165);
nand U3249 (N_3249,N_3151,N_3147);
nor U3250 (N_3250,N_3130,N_3143);
xor U3251 (N_3251,N_3120,N_3130);
nand U3252 (N_3252,N_3119,N_3101);
nand U3253 (N_3253,N_3172,N_3133);
or U3254 (N_3254,N_3183,N_3106);
nand U3255 (N_3255,N_3199,N_3116);
nor U3256 (N_3256,N_3113,N_3175);
and U3257 (N_3257,N_3145,N_3127);
or U3258 (N_3258,N_3102,N_3181);
nor U3259 (N_3259,N_3181,N_3190);
nor U3260 (N_3260,N_3178,N_3149);
and U3261 (N_3261,N_3146,N_3159);
nor U3262 (N_3262,N_3152,N_3195);
nor U3263 (N_3263,N_3131,N_3103);
and U3264 (N_3264,N_3135,N_3171);
nand U3265 (N_3265,N_3183,N_3131);
or U3266 (N_3266,N_3151,N_3181);
nor U3267 (N_3267,N_3191,N_3178);
and U3268 (N_3268,N_3114,N_3132);
nand U3269 (N_3269,N_3108,N_3169);
or U3270 (N_3270,N_3151,N_3157);
nand U3271 (N_3271,N_3195,N_3113);
nand U3272 (N_3272,N_3127,N_3122);
nand U3273 (N_3273,N_3160,N_3174);
or U3274 (N_3274,N_3157,N_3119);
and U3275 (N_3275,N_3189,N_3177);
xnor U3276 (N_3276,N_3100,N_3177);
or U3277 (N_3277,N_3131,N_3187);
nand U3278 (N_3278,N_3129,N_3160);
and U3279 (N_3279,N_3161,N_3113);
or U3280 (N_3280,N_3109,N_3184);
or U3281 (N_3281,N_3188,N_3149);
nor U3282 (N_3282,N_3105,N_3123);
or U3283 (N_3283,N_3189,N_3148);
and U3284 (N_3284,N_3135,N_3122);
nor U3285 (N_3285,N_3163,N_3177);
nand U3286 (N_3286,N_3119,N_3197);
and U3287 (N_3287,N_3134,N_3124);
nand U3288 (N_3288,N_3113,N_3166);
or U3289 (N_3289,N_3169,N_3189);
or U3290 (N_3290,N_3151,N_3121);
nand U3291 (N_3291,N_3177,N_3125);
and U3292 (N_3292,N_3160,N_3136);
nand U3293 (N_3293,N_3103,N_3137);
and U3294 (N_3294,N_3105,N_3188);
nand U3295 (N_3295,N_3161,N_3149);
nand U3296 (N_3296,N_3164,N_3166);
xor U3297 (N_3297,N_3130,N_3137);
nor U3298 (N_3298,N_3149,N_3176);
nand U3299 (N_3299,N_3101,N_3189);
xor U3300 (N_3300,N_3276,N_3237);
or U3301 (N_3301,N_3241,N_3219);
nand U3302 (N_3302,N_3268,N_3240);
or U3303 (N_3303,N_3274,N_3295);
and U3304 (N_3304,N_3258,N_3281);
nor U3305 (N_3305,N_3212,N_3255);
nor U3306 (N_3306,N_3204,N_3290);
xnor U3307 (N_3307,N_3248,N_3251);
or U3308 (N_3308,N_3233,N_3298);
xnor U3309 (N_3309,N_3236,N_3263);
nand U3310 (N_3310,N_3259,N_3282);
nand U3311 (N_3311,N_3252,N_3288);
nor U3312 (N_3312,N_3223,N_3222);
nor U3313 (N_3313,N_3247,N_3243);
and U3314 (N_3314,N_3228,N_3253);
nand U3315 (N_3315,N_3264,N_3227);
or U3316 (N_3316,N_3234,N_3265);
or U3317 (N_3317,N_3260,N_3296);
nand U3318 (N_3318,N_3283,N_3206);
or U3319 (N_3319,N_3272,N_3286);
nand U3320 (N_3320,N_3249,N_3213);
nand U3321 (N_3321,N_3230,N_3218);
nor U3322 (N_3322,N_3291,N_3279);
and U3323 (N_3323,N_3232,N_3254);
xnor U3324 (N_3324,N_3246,N_3266);
xnor U3325 (N_3325,N_3225,N_3242);
or U3326 (N_3326,N_3209,N_3256);
nor U3327 (N_3327,N_3220,N_3207);
or U3328 (N_3328,N_3297,N_3257);
and U3329 (N_3329,N_3294,N_3210);
nand U3330 (N_3330,N_3285,N_3208);
nor U3331 (N_3331,N_3261,N_3269);
nor U3332 (N_3332,N_3250,N_3262);
nand U3333 (N_3333,N_3215,N_3200);
nand U3334 (N_3334,N_3292,N_3289);
nor U3335 (N_3335,N_3299,N_3275);
or U3336 (N_3336,N_3229,N_3216);
nor U3337 (N_3337,N_3278,N_3280);
xor U3338 (N_3338,N_3284,N_3245);
xor U3339 (N_3339,N_3287,N_3201);
nor U3340 (N_3340,N_3221,N_3238);
nor U3341 (N_3341,N_3239,N_3277);
xnor U3342 (N_3342,N_3226,N_3293);
and U3343 (N_3343,N_3205,N_3244);
xnor U3344 (N_3344,N_3270,N_3271);
or U3345 (N_3345,N_3273,N_3235);
nand U3346 (N_3346,N_3224,N_3211);
and U3347 (N_3347,N_3202,N_3214);
xnor U3348 (N_3348,N_3231,N_3203);
nand U3349 (N_3349,N_3217,N_3267);
or U3350 (N_3350,N_3226,N_3257);
nand U3351 (N_3351,N_3251,N_3235);
and U3352 (N_3352,N_3270,N_3229);
and U3353 (N_3353,N_3201,N_3237);
and U3354 (N_3354,N_3260,N_3293);
and U3355 (N_3355,N_3251,N_3263);
nand U3356 (N_3356,N_3206,N_3240);
nand U3357 (N_3357,N_3228,N_3264);
nor U3358 (N_3358,N_3284,N_3203);
nand U3359 (N_3359,N_3280,N_3293);
and U3360 (N_3360,N_3267,N_3270);
nand U3361 (N_3361,N_3208,N_3263);
and U3362 (N_3362,N_3230,N_3203);
or U3363 (N_3363,N_3237,N_3222);
nor U3364 (N_3364,N_3204,N_3267);
and U3365 (N_3365,N_3252,N_3276);
or U3366 (N_3366,N_3262,N_3261);
nor U3367 (N_3367,N_3227,N_3240);
or U3368 (N_3368,N_3292,N_3280);
or U3369 (N_3369,N_3276,N_3242);
xor U3370 (N_3370,N_3231,N_3243);
nand U3371 (N_3371,N_3241,N_3247);
nand U3372 (N_3372,N_3207,N_3295);
and U3373 (N_3373,N_3203,N_3277);
xor U3374 (N_3374,N_3211,N_3225);
or U3375 (N_3375,N_3254,N_3212);
nand U3376 (N_3376,N_3276,N_3228);
and U3377 (N_3377,N_3270,N_3289);
and U3378 (N_3378,N_3204,N_3256);
and U3379 (N_3379,N_3214,N_3208);
or U3380 (N_3380,N_3210,N_3291);
or U3381 (N_3381,N_3211,N_3239);
or U3382 (N_3382,N_3245,N_3231);
and U3383 (N_3383,N_3276,N_3290);
xor U3384 (N_3384,N_3233,N_3284);
xnor U3385 (N_3385,N_3238,N_3276);
xnor U3386 (N_3386,N_3261,N_3288);
nor U3387 (N_3387,N_3251,N_3259);
or U3388 (N_3388,N_3297,N_3268);
and U3389 (N_3389,N_3234,N_3216);
nor U3390 (N_3390,N_3205,N_3208);
and U3391 (N_3391,N_3259,N_3242);
or U3392 (N_3392,N_3268,N_3239);
and U3393 (N_3393,N_3208,N_3256);
nand U3394 (N_3394,N_3217,N_3259);
xnor U3395 (N_3395,N_3211,N_3223);
and U3396 (N_3396,N_3297,N_3205);
nand U3397 (N_3397,N_3230,N_3253);
nand U3398 (N_3398,N_3258,N_3247);
nand U3399 (N_3399,N_3269,N_3215);
nand U3400 (N_3400,N_3359,N_3343);
nor U3401 (N_3401,N_3318,N_3398);
or U3402 (N_3402,N_3351,N_3303);
xor U3403 (N_3403,N_3310,N_3326);
xnor U3404 (N_3404,N_3306,N_3355);
and U3405 (N_3405,N_3338,N_3319);
and U3406 (N_3406,N_3388,N_3376);
or U3407 (N_3407,N_3312,N_3387);
xor U3408 (N_3408,N_3329,N_3366);
nand U3409 (N_3409,N_3362,N_3328);
nor U3410 (N_3410,N_3380,N_3399);
nand U3411 (N_3411,N_3322,N_3368);
nand U3412 (N_3412,N_3367,N_3377);
or U3413 (N_3413,N_3308,N_3342);
nand U3414 (N_3414,N_3337,N_3372);
nand U3415 (N_3415,N_3384,N_3393);
and U3416 (N_3416,N_3320,N_3360);
and U3417 (N_3417,N_3327,N_3321);
nor U3418 (N_3418,N_3374,N_3379);
nand U3419 (N_3419,N_3370,N_3301);
nor U3420 (N_3420,N_3389,N_3344);
and U3421 (N_3421,N_3363,N_3345);
and U3422 (N_3422,N_3390,N_3302);
or U3423 (N_3423,N_3365,N_3331);
nor U3424 (N_3424,N_3324,N_3314);
and U3425 (N_3425,N_3349,N_3332);
nor U3426 (N_3426,N_3313,N_3357);
nand U3427 (N_3427,N_3341,N_3382);
and U3428 (N_3428,N_3373,N_3333);
nor U3429 (N_3429,N_3307,N_3381);
nand U3430 (N_3430,N_3300,N_3347);
and U3431 (N_3431,N_3325,N_3354);
nor U3432 (N_3432,N_3330,N_3346);
or U3433 (N_3433,N_3350,N_3339);
nor U3434 (N_3434,N_3353,N_3356);
or U3435 (N_3435,N_3311,N_3348);
nor U3436 (N_3436,N_3396,N_3334);
and U3437 (N_3437,N_3375,N_3385);
or U3438 (N_3438,N_3394,N_3352);
xor U3439 (N_3439,N_3386,N_3335);
nor U3440 (N_3440,N_3340,N_3304);
nor U3441 (N_3441,N_3323,N_3316);
xor U3442 (N_3442,N_3397,N_3305);
or U3443 (N_3443,N_3358,N_3395);
and U3444 (N_3444,N_3369,N_3383);
or U3445 (N_3445,N_3371,N_3317);
or U3446 (N_3446,N_3361,N_3392);
and U3447 (N_3447,N_3309,N_3336);
and U3448 (N_3448,N_3391,N_3315);
nand U3449 (N_3449,N_3378,N_3364);
and U3450 (N_3450,N_3335,N_3379);
nand U3451 (N_3451,N_3324,N_3353);
xnor U3452 (N_3452,N_3323,N_3350);
or U3453 (N_3453,N_3322,N_3330);
and U3454 (N_3454,N_3333,N_3319);
nand U3455 (N_3455,N_3361,N_3350);
nand U3456 (N_3456,N_3385,N_3313);
or U3457 (N_3457,N_3372,N_3341);
nor U3458 (N_3458,N_3345,N_3349);
and U3459 (N_3459,N_3399,N_3326);
and U3460 (N_3460,N_3364,N_3355);
nand U3461 (N_3461,N_3356,N_3398);
nor U3462 (N_3462,N_3394,N_3385);
or U3463 (N_3463,N_3399,N_3386);
and U3464 (N_3464,N_3325,N_3351);
and U3465 (N_3465,N_3387,N_3366);
nor U3466 (N_3466,N_3367,N_3398);
or U3467 (N_3467,N_3352,N_3324);
nand U3468 (N_3468,N_3361,N_3360);
or U3469 (N_3469,N_3321,N_3382);
xnor U3470 (N_3470,N_3399,N_3374);
or U3471 (N_3471,N_3303,N_3386);
nand U3472 (N_3472,N_3363,N_3322);
xor U3473 (N_3473,N_3304,N_3325);
and U3474 (N_3474,N_3367,N_3307);
and U3475 (N_3475,N_3316,N_3330);
xnor U3476 (N_3476,N_3391,N_3320);
xor U3477 (N_3477,N_3326,N_3384);
or U3478 (N_3478,N_3363,N_3337);
nand U3479 (N_3479,N_3320,N_3398);
xnor U3480 (N_3480,N_3354,N_3318);
nand U3481 (N_3481,N_3304,N_3384);
and U3482 (N_3482,N_3339,N_3334);
nor U3483 (N_3483,N_3347,N_3338);
nand U3484 (N_3484,N_3334,N_3363);
nand U3485 (N_3485,N_3307,N_3305);
or U3486 (N_3486,N_3317,N_3301);
or U3487 (N_3487,N_3374,N_3309);
nor U3488 (N_3488,N_3315,N_3363);
or U3489 (N_3489,N_3310,N_3324);
or U3490 (N_3490,N_3353,N_3357);
nand U3491 (N_3491,N_3342,N_3325);
nand U3492 (N_3492,N_3374,N_3378);
nor U3493 (N_3493,N_3329,N_3350);
nand U3494 (N_3494,N_3315,N_3385);
nand U3495 (N_3495,N_3378,N_3300);
nor U3496 (N_3496,N_3382,N_3398);
xor U3497 (N_3497,N_3314,N_3360);
xnor U3498 (N_3498,N_3331,N_3327);
nor U3499 (N_3499,N_3394,N_3389);
xnor U3500 (N_3500,N_3476,N_3432);
nor U3501 (N_3501,N_3496,N_3403);
nor U3502 (N_3502,N_3467,N_3413);
xnor U3503 (N_3503,N_3453,N_3404);
nand U3504 (N_3504,N_3429,N_3414);
or U3505 (N_3505,N_3495,N_3479);
nand U3506 (N_3506,N_3472,N_3465);
nand U3507 (N_3507,N_3489,N_3422);
xnor U3508 (N_3508,N_3400,N_3477);
nand U3509 (N_3509,N_3481,N_3427);
and U3510 (N_3510,N_3433,N_3487);
nor U3511 (N_3511,N_3450,N_3462);
or U3512 (N_3512,N_3470,N_3485);
and U3513 (N_3513,N_3452,N_3445);
and U3514 (N_3514,N_3446,N_3475);
nand U3515 (N_3515,N_3461,N_3439);
and U3516 (N_3516,N_3402,N_3420);
nand U3517 (N_3517,N_3469,N_3442);
or U3518 (N_3518,N_3490,N_3494);
xnor U3519 (N_3519,N_3415,N_3497);
nor U3520 (N_3520,N_3410,N_3449);
or U3521 (N_3521,N_3438,N_3457);
and U3522 (N_3522,N_3498,N_3468);
xor U3523 (N_3523,N_3491,N_3412);
xor U3524 (N_3524,N_3411,N_3488);
and U3525 (N_3525,N_3408,N_3440);
or U3526 (N_3526,N_3493,N_3464);
and U3527 (N_3527,N_3405,N_3417);
nand U3528 (N_3528,N_3480,N_3434);
or U3529 (N_3529,N_3409,N_3406);
or U3530 (N_3530,N_3478,N_3471);
nor U3531 (N_3531,N_3483,N_3423);
nor U3532 (N_3532,N_3418,N_3474);
nor U3533 (N_3533,N_3421,N_3419);
nor U3534 (N_3534,N_3451,N_3425);
and U3535 (N_3535,N_3435,N_3444);
or U3536 (N_3536,N_3437,N_3486);
or U3537 (N_3537,N_3441,N_3443);
nand U3538 (N_3538,N_3407,N_3458);
xor U3539 (N_3539,N_3428,N_3460);
nor U3540 (N_3540,N_3447,N_3431);
nand U3541 (N_3541,N_3492,N_3424);
or U3542 (N_3542,N_3430,N_3499);
nor U3543 (N_3543,N_3482,N_3416);
or U3544 (N_3544,N_3484,N_3466);
or U3545 (N_3545,N_3448,N_3463);
and U3546 (N_3546,N_3454,N_3473);
nand U3547 (N_3547,N_3455,N_3426);
or U3548 (N_3548,N_3456,N_3459);
or U3549 (N_3549,N_3436,N_3401);
nand U3550 (N_3550,N_3469,N_3445);
and U3551 (N_3551,N_3490,N_3436);
or U3552 (N_3552,N_3409,N_3459);
and U3553 (N_3553,N_3427,N_3486);
nor U3554 (N_3554,N_3467,N_3434);
nand U3555 (N_3555,N_3464,N_3488);
nor U3556 (N_3556,N_3469,N_3485);
nor U3557 (N_3557,N_3420,N_3425);
and U3558 (N_3558,N_3479,N_3488);
nor U3559 (N_3559,N_3477,N_3464);
xnor U3560 (N_3560,N_3459,N_3429);
nand U3561 (N_3561,N_3404,N_3450);
xor U3562 (N_3562,N_3428,N_3456);
and U3563 (N_3563,N_3422,N_3488);
nand U3564 (N_3564,N_3440,N_3492);
nand U3565 (N_3565,N_3417,N_3434);
or U3566 (N_3566,N_3407,N_3405);
or U3567 (N_3567,N_3494,N_3486);
or U3568 (N_3568,N_3464,N_3481);
nand U3569 (N_3569,N_3407,N_3438);
nor U3570 (N_3570,N_3414,N_3492);
and U3571 (N_3571,N_3410,N_3460);
and U3572 (N_3572,N_3493,N_3475);
nor U3573 (N_3573,N_3416,N_3449);
nor U3574 (N_3574,N_3466,N_3441);
nor U3575 (N_3575,N_3423,N_3403);
nor U3576 (N_3576,N_3441,N_3454);
nand U3577 (N_3577,N_3411,N_3485);
and U3578 (N_3578,N_3450,N_3465);
or U3579 (N_3579,N_3491,N_3472);
xor U3580 (N_3580,N_3473,N_3489);
xnor U3581 (N_3581,N_3495,N_3405);
and U3582 (N_3582,N_3408,N_3483);
or U3583 (N_3583,N_3403,N_3469);
or U3584 (N_3584,N_3437,N_3456);
or U3585 (N_3585,N_3401,N_3409);
or U3586 (N_3586,N_3456,N_3473);
or U3587 (N_3587,N_3466,N_3496);
and U3588 (N_3588,N_3423,N_3405);
nand U3589 (N_3589,N_3414,N_3411);
nand U3590 (N_3590,N_3469,N_3450);
or U3591 (N_3591,N_3459,N_3476);
and U3592 (N_3592,N_3409,N_3460);
nor U3593 (N_3593,N_3468,N_3467);
nand U3594 (N_3594,N_3434,N_3411);
nor U3595 (N_3595,N_3411,N_3407);
nand U3596 (N_3596,N_3499,N_3418);
or U3597 (N_3597,N_3427,N_3442);
and U3598 (N_3598,N_3496,N_3476);
xor U3599 (N_3599,N_3467,N_3496);
nand U3600 (N_3600,N_3584,N_3521);
xnor U3601 (N_3601,N_3546,N_3519);
nand U3602 (N_3602,N_3573,N_3568);
or U3603 (N_3603,N_3555,N_3542);
and U3604 (N_3604,N_3502,N_3539);
and U3605 (N_3605,N_3569,N_3545);
nor U3606 (N_3606,N_3572,N_3591);
or U3607 (N_3607,N_3505,N_3523);
nand U3608 (N_3608,N_3578,N_3500);
nor U3609 (N_3609,N_3597,N_3552);
nor U3610 (N_3610,N_3535,N_3501);
or U3611 (N_3611,N_3565,N_3508);
xnor U3612 (N_3612,N_3560,N_3512);
or U3613 (N_3613,N_3503,N_3564);
and U3614 (N_3614,N_3596,N_3557);
nor U3615 (N_3615,N_3507,N_3524);
xor U3616 (N_3616,N_3561,N_3588);
or U3617 (N_3617,N_3549,N_3506);
xnor U3618 (N_3618,N_3558,N_3554);
xor U3619 (N_3619,N_3515,N_3528);
or U3620 (N_3620,N_3598,N_3571);
or U3621 (N_3621,N_3579,N_3594);
or U3622 (N_3622,N_3536,N_3525);
and U3623 (N_3623,N_3581,N_3595);
and U3624 (N_3624,N_3537,N_3513);
or U3625 (N_3625,N_3530,N_3593);
and U3626 (N_3626,N_3587,N_3551);
and U3627 (N_3627,N_3526,N_3544);
nand U3628 (N_3628,N_3580,N_3520);
nor U3629 (N_3629,N_3559,N_3563);
nor U3630 (N_3630,N_3531,N_3514);
xor U3631 (N_3631,N_3582,N_3550);
xnor U3632 (N_3632,N_3547,N_3548);
nand U3633 (N_3633,N_3533,N_3583);
nor U3634 (N_3634,N_3570,N_3576);
nand U3635 (N_3635,N_3504,N_3574);
or U3636 (N_3636,N_3586,N_3577);
nor U3637 (N_3637,N_3517,N_3510);
and U3638 (N_3638,N_3590,N_3566);
nand U3639 (N_3639,N_3553,N_3575);
nand U3640 (N_3640,N_3516,N_3522);
xnor U3641 (N_3641,N_3541,N_3585);
or U3642 (N_3642,N_3543,N_3592);
nor U3643 (N_3643,N_3540,N_3511);
or U3644 (N_3644,N_3599,N_3527);
or U3645 (N_3645,N_3518,N_3532);
or U3646 (N_3646,N_3562,N_3534);
nor U3647 (N_3647,N_3556,N_3538);
nand U3648 (N_3648,N_3509,N_3567);
and U3649 (N_3649,N_3589,N_3529);
nor U3650 (N_3650,N_3519,N_3581);
nor U3651 (N_3651,N_3521,N_3588);
or U3652 (N_3652,N_3505,N_3520);
nor U3653 (N_3653,N_3527,N_3542);
and U3654 (N_3654,N_3514,N_3547);
nand U3655 (N_3655,N_3540,N_3534);
or U3656 (N_3656,N_3557,N_3501);
or U3657 (N_3657,N_3558,N_3579);
and U3658 (N_3658,N_3543,N_3578);
nor U3659 (N_3659,N_3571,N_3599);
nor U3660 (N_3660,N_3570,N_3566);
nor U3661 (N_3661,N_3505,N_3518);
xor U3662 (N_3662,N_3502,N_3530);
xor U3663 (N_3663,N_3583,N_3526);
nor U3664 (N_3664,N_3557,N_3502);
xnor U3665 (N_3665,N_3580,N_3532);
xor U3666 (N_3666,N_3502,N_3513);
nand U3667 (N_3667,N_3517,N_3501);
xnor U3668 (N_3668,N_3594,N_3557);
nor U3669 (N_3669,N_3571,N_3520);
and U3670 (N_3670,N_3587,N_3512);
nor U3671 (N_3671,N_3500,N_3581);
xnor U3672 (N_3672,N_3593,N_3521);
nand U3673 (N_3673,N_3510,N_3574);
or U3674 (N_3674,N_3519,N_3542);
nor U3675 (N_3675,N_3500,N_3538);
nor U3676 (N_3676,N_3587,N_3520);
or U3677 (N_3677,N_3508,N_3548);
nor U3678 (N_3678,N_3528,N_3506);
nand U3679 (N_3679,N_3587,N_3568);
and U3680 (N_3680,N_3561,N_3596);
nor U3681 (N_3681,N_3558,N_3549);
nor U3682 (N_3682,N_3533,N_3555);
nor U3683 (N_3683,N_3572,N_3573);
and U3684 (N_3684,N_3551,N_3544);
and U3685 (N_3685,N_3510,N_3590);
and U3686 (N_3686,N_3554,N_3565);
xor U3687 (N_3687,N_3576,N_3565);
nor U3688 (N_3688,N_3555,N_3526);
or U3689 (N_3689,N_3541,N_3529);
or U3690 (N_3690,N_3544,N_3523);
nor U3691 (N_3691,N_3521,N_3555);
or U3692 (N_3692,N_3588,N_3509);
nor U3693 (N_3693,N_3521,N_3570);
and U3694 (N_3694,N_3515,N_3558);
or U3695 (N_3695,N_3527,N_3552);
and U3696 (N_3696,N_3538,N_3501);
nand U3697 (N_3697,N_3507,N_3510);
or U3698 (N_3698,N_3553,N_3516);
nand U3699 (N_3699,N_3523,N_3502);
and U3700 (N_3700,N_3667,N_3659);
xor U3701 (N_3701,N_3683,N_3650);
or U3702 (N_3702,N_3625,N_3609);
or U3703 (N_3703,N_3696,N_3699);
or U3704 (N_3704,N_3642,N_3635);
and U3705 (N_3705,N_3620,N_3673);
and U3706 (N_3706,N_3627,N_3658);
and U3707 (N_3707,N_3665,N_3628);
or U3708 (N_3708,N_3653,N_3669);
or U3709 (N_3709,N_3685,N_3668);
and U3710 (N_3710,N_3612,N_3606);
nand U3711 (N_3711,N_3652,N_3662);
xnor U3712 (N_3712,N_3684,N_3651);
nor U3713 (N_3713,N_3611,N_3641);
nand U3714 (N_3714,N_3693,N_3697);
nor U3715 (N_3715,N_3676,N_3630);
nand U3716 (N_3716,N_3604,N_3624);
or U3717 (N_3717,N_3621,N_3608);
nor U3718 (N_3718,N_3681,N_3600);
and U3719 (N_3719,N_3618,N_3622);
nand U3720 (N_3720,N_3626,N_3664);
nand U3721 (N_3721,N_3616,N_3623);
nor U3722 (N_3722,N_3610,N_3613);
and U3723 (N_3723,N_3640,N_3649);
and U3724 (N_3724,N_3692,N_3634);
nor U3725 (N_3725,N_3686,N_3629);
nor U3726 (N_3726,N_3679,N_3643);
xnor U3727 (N_3727,N_3677,N_3670);
nand U3728 (N_3728,N_3603,N_3639);
and U3729 (N_3729,N_3637,N_3698);
and U3730 (N_3730,N_3682,N_3631);
or U3731 (N_3731,N_3633,N_3638);
or U3732 (N_3732,N_3646,N_3671);
nor U3733 (N_3733,N_3601,N_3645);
or U3734 (N_3734,N_3617,N_3687);
nand U3735 (N_3735,N_3632,N_3657);
xor U3736 (N_3736,N_3614,N_3680);
nand U3737 (N_3737,N_3656,N_3694);
nor U3738 (N_3738,N_3648,N_3644);
or U3739 (N_3739,N_3666,N_3605);
nor U3740 (N_3740,N_3689,N_3661);
nor U3741 (N_3741,N_3615,N_3660);
nand U3742 (N_3742,N_3678,N_3672);
nor U3743 (N_3743,N_3636,N_3602);
xor U3744 (N_3744,N_3607,N_3688);
nand U3745 (N_3745,N_3619,N_3655);
or U3746 (N_3746,N_3695,N_3675);
nor U3747 (N_3747,N_3674,N_3647);
xor U3748 (N_3748,N_3691,N_3654);
or U3749 (N_3749,N_3690,N_3663);
and U3750 (N_3750,N_3667,N_3670);
nand U3751 (N_3751,N_3652,N_3619);
nor U3752 (N_3752,N_3685,N_3622);
or U3753 (N_3753,N_3636,N_3692);
or U3754 (N_3754,N_3677,N_3667);
or U3755 (N_3755,N_3622,N_3691);
nand U3756 (N_3756,N_3651,N_3680);
or U3757 (N_3757,N_3623,N_3618);
nor U3758 (N_3758,N_3642,N_3654);
nand U3759 (N_3759,N_3687,N_3607);
and U3760 (N_3760,N_3677,N_3650);
and U3761 (N_3761,N_3672,N_3651);
xnor U3762 (N_3762,N_3693,N_3627);
and U3763 (N_3763,N_3683,N_3634);
nor U3764 (N_3764,N_3634,N_3670);
nand U3765 (N_3765,N_3678,N_3601);
nand U3766 (N_3766,N_3678,N_3674);
and U3767 (N_3767,N_3631,N_3650);
and U3768 (N_3768,N_3695,N_3670);
nand U3769 (N_3769,N_3634,N_3638);
xor U3770 (N_3770,N_3694,N_3647);
xor U3771 (N_3771,N_3690,N_3637);
or U3772 (N_3772,N_3690,N_3656);
or U3773 (N_3773,N_3611,N_3699);
or U3774 (N_3774,N_3634,N_3629);
xnor U3775 (N_3775,N_3689,N_3652);
xnor U3776 (N_3776,N_3641,N_3649);
and U3777 (N_3777,N_3613,N_3664);
and U3778 (N_3778,N_3664,N_3673);
and U3779 (N_3779,N_3630,N_3637);
nand U3780 (N_3780,N_3642,N_3670);
nor U3781 (N_3781,N_3692,N_3632);
or U3782 (N_3782,N_3607,N_3647);
xnor U3783 (N_3783,N_3666,N_3607);
or U3784 (N_3784,N_3645,N_3655);
nor U3785 (N_3785,N_3648,N_3697);
or U3786 (N_3786,N_3677,N_3621);
nand U3787 (N_3787,N_3661,N_3697);
xnor U3788 (N_3788,N_3635,N_3696);
nand U3789 (N_3789,N_3620,N_3618);
xnor U3790 (N_3790,N_3602,N_3619);
and U3791 (N_3791,N_3691,N_3637);
and U3792 (N_3792,N_3601,N_3606);
or U3793 (N_3793,N_3622,N_3629);
nor U3794 (N_3794,N_3604,N_3603);
and U3795 (N_3795,N_3660,N_3610);
and U3796 (N_3796,N_3639,N_3655);
nand U3797 (N_3797,N_3644,N_3627);
nor U3798 (N_3798,N_3682,N_3640);
nand U3799 (N_3799,N_3692,N_3681);
and U3800 (N_3800,N_3738,N_3720);
or U3801 (N_3801,N_3760,N_3787);
nand U3802 (N_3802,N_3757,N_3745);
nor U3803 (N_3803,N_3734,N_3764);
and U3804 (N_3804,N_3726,N_3796);
xor U3805 (N_3805,N_3789,N_3731);
nor U3806 (N_3806,N_3710,N_3759);
nor U3807 (N_3807,N_3761,N_3752);
nand U3808 (N_3808,N_3723,N_3769);
and U3809 (N_3809,N_3724,N_3703);
and U3810 (N_3810,N_3727,N_3777);
nor U3811 (N_3811,N_3729,N_3722);
and U3812 (N_3812,N_3756,N_3762);
or U3813 (N_3813,N_3740,N_3792);
and U3814 (N_3814,N_3750,N_3758);
and U3815 (N_3815,N_3709,N_3728);
nand U3816 (N_3816,N_3798,N_3735);
nand U3817 (N_3817,N_3793,N_3716);
nor U3818 (N_3818,N_3799,N_3784);
nor U3819 (N_3819,N_3737,N_3770);
and U3820 (N_3820,N_3779,N_3744);
and U3821 (N_3821,N_3732,N_3749);
and U3822 (N_3822,N_3781,N_3783);
nor U3823 (N_3823,N_3776,N_3733);
xor U3824 (N_3824,N_3701,N_3771);
and U3825 (N_3825,N_3753,N_3788);
or U3826 (N_3826,N_3713,N_3718);
or U3827 (N_3827,N_3775,N_3700);
and U3828 (N_3828,N_3702,N_3778);
and U3829 (N_3829,N_3767,N_3795);
and U3830 (N_3830,N_3774,N_3707);
nand U3831 (N_3831,N_3785,N_3797);
and U3832 (N_3832,N_3715,N_3721);
or U3833 (N_3833,N_3773,N_3786);
nor U3834 (N_3834,N_3743,N_3790);
nor U3835 (N_3835,N_3711,N_3719);
and U3836 (N_3836,N_3708,N_3747);
or U3837 (N_3837,N_3763,N_3754);
nor U3838 (N_3838,N_3712,N_3766);
nand U3839 (N_3839,N_3751,N_3755);
nor U3840 (N_3840,N_3765,N_3782);
nand U3841 (N_3841,N_3748,N_3714);
nor U3842 (N_3842,N_3742,N_3741);
or U3843 (N_3843,N_3705,N_3794);
nor U3844 (N_3844,N_3772,N_3768);
or U3845 (N_3845,N_3746,N_3725);
nor U3846 (N_3846,N_3704,N_3739);
nor U3847 (N_3847,N_3736,N_3706);
nand U3848 (N_3848,N_3730,N_3780);
or U3849 (N_3849,N_3717,N_3791);
and U3850 (N_3850,N_3736,N_3789);
xnor U3851 (N_3851,N_3796,N_3714);
nand U3852 (N_3852,N_3718,N_3775);
and U3853 (N_3853,N_3747,N_3721);
xor U3854 (N_3854,N_3743,N_3709);
nand U3855 (N_3855,N_3779,N_3762);
and U3856 (N_3856,N_3750,N_3773);
and U3857 (N_3857,N_3712,N_3796);
or U3858 (N_3858,N_3745,N_3709);
nand U3859 (N_3859,N_3797,N_3773);
nor U3860 (N_3860,N_3720,N_3708);
or U3861 (N_3861,N_3761,N_3701);
nand U3862 (N_3862,N_3788,N_3751);
nor U3863 (N_3863,N_3782,N_3778);
xor U3864 (N_3864,N_3715,N_3796);
and U3865 (N_3865,N_3771,N_3717);
xor U3866 (N_3866,N_3759,N_3768);
nor U3867 (N_3867,N_3783,N_3780);
xnor U3868 (N_3868,N_3718,N_3757);
nand U3869 (N_3869,N_3729,N_3785);
nand U3870 (N_3870,N_3751,N_3714);
or U3871 (N_3871,N_3752,N_3730);
and U3872 (N_3872,N_3717,N_3761);
and U3873 (N_3873,N_3781,N_3776);
or U3874 (N_3874,N_3773,N_3718);
nor U3875 (N_3875,N_3731,N_3709);
or U3876 (N_3876,N_3739,N_3767);
nand U3877 (N_3877,N_3719,N_3724);
or U3878 (N_3878,N_3728,N_3706);
or U3879 (N_3879,N_3705,N_3791);
or U3880 (N_3880,N_3765,N_3795);
nor U3881 (N_3881,N_3786,N_3712);
and U3882 (N_3882,N_3700,N_3752);
and U3883 (N_3883,N_3701,N_3784);
nand U3884 (N_3884,N_3761,N_3710);
or U3885 (N_3885,N_3732,N_3754);
xor U3886 (N_3886,N_3777,N_3773);
nor U3887 (N_3887,N_3774,N_3777);
nand U3888 (N_3888,N_3771,N_3733);
xnor U3889 (N_3889,N_3740,N_3720);
xor U3890 (N_3890,N_3703,N_3773);
and U3891 (N_3891,N_3774,N_3794);
nand U3892 (N_3892,N_3721,N_3761);
or U3893 (N_3893,N_3745,N_3724);
or U3894 (N_3894,N_3757,N_3746);
nand U3895 (N_3895,N_3751,N_3766);
xor U3896 (N_3896,N_3760,N_3762);
xor U3897 (N_3897,N_3708,N_3765);
nand U3898 (N_3898,N_3714,N_3798);
nor U3899 (N_3899,N_3771,N_3722);
nand U3900 (N_3900,N_3851,N_3883);
nor U3901 (N_3901,N_3853,N_3821);
or U3902 (N_3902,N_3828,N_3845);
nand U3903 (N_3903,N_3824,N_3865);
and U3904 (N_3904,N_3815,N_3816);
nor U3905 (N_3905,N_3836,N_3849);
or U3906 (N_3906,N_3889,N_3856);
nor U3907 (N_3907,N_3869,N_3826);
or U3908 (N_3908,N_3846,N_3818);
or U3909 (N_3909,N_3823,N_3885);
or U3910 (N_3910,N_3806,N_3878);
and U3911 (N_3911,N_3866,N_3868);
nand U3912 (N_3912,N_3855,N_3841);
nand U3913 (N_3913,N_3873,N_3861);
nand U3914 (N_3914,N_3874,N_3893);
and U3915 (N_3915,N_3842,N_3872);
nor U3916 (N_3916,N_3882,N_3850);
and U3917 (N_3917,N_3870,N_3822);
nor U3918 (N_3918,N_3847,N_3854);
nand U3919 (N_3919,N_3810,N_3860);
or U3920 (N_3920,N_3899,N_3813);
and U3921 (N_3921,N_3890,N_3884);
xor U3922 (N_3922,N_3805,N_3838);
or U3923 (N_3923,N_3829,N_3864);
and U3924 (N_3924,N_3880,N_3814);
or U3925 (N_3925,N_3825,N_3820);
nand U3926 (N_3926,N_3819,N_3831);
nor U3927 (N_3927,N_3858,N_3879);
nor U3928 (N_3928,N_3817,N_3802);
nand U3929 (N_3929,N_3827,N_3895);
and U3930 (N_3930,N_3891,N_3896);
nor U3931 (N_3931,N_3835,N_3833);
or U3932 (N_3932,N_3843,N_3837);
or U3933 (N_3933,N_3871,N_3839);
or U3934 (N_3934,N_3848,N_3830);
and U3935 (N_3935,N_3832,N_3867);
nor U3936 (N_3936,N_3800,N_3862);
and U3937 (N_3937,N_3875,N_3844);
and U3938 (N_3938,N_3894,N_3886);
nor U3939 (N_3939,N_3876,N_3811);
nand U3940 (N_3940,N_3888,N_3808);
nor U3941 (N_3941,N_3834,N_3897);
nand U3942 (N_3942,N_3881,N_3887);
nand U3943 (N_3943,N_3863,N_3877);
and U3944 (N_3944,N_3898,N_3804);
and U3945 (N_3945,N_3807,N_3812);
nor U3946 (N_3946,N_3840,N_3859);
and U3947 (N_3947,N_3852,N_3809);
or U3948 (N_3948,N_3801,N_3803);
nor U3949 (N_3949,N_3892,N_3857);
or U3950 (N_3950,N_3812,N_3882);
and U3951 (N_3951,N_3843,N_3855);
xor U3952 (N_3952,N_3813,N_3889);
nand U3953 (N_3953,N_3868,N_3841);
nand U3954 (N_3954,N_3891,N_3823);
and U3955 (N_3955,N_3864,N_3860);
or U3956 (N_3956,N_3804,N_3810);
nand U3957 (N_3957,N_3845,N_3801);
nor U3958 (N_3958,N_3890,N_3808);
nand U3959 (N_3959,N_3820,N_3863);
nand U3960 (N_3960,N_3819,N_3818);
or U3961 (N_3961,N_3848,N_3877);
xor U3962 (N_3962,N_3811,N_3861);
nand U3963 (N_3963,N_3851,N_3848);
xnor U3964 (N_3964,N_3808,N_3842);
nor U3965 (N_3965,N_3853,N_3862);
nor U3966 (N_3966,N_3862,N_3842);
and U3967 (N_3967,N_3847,N_3862);
and U3968 (N_3968,N_3855,N_3811);
and U3969 (N_3969,N_3847,N_3877);
nor U3970 (N_3970,N_3808,N_3850);
nand U3971 (N_3971,N_3894,N_3878);
nand U3972 (N_3972,N_3838,N_3808);
nand U3973 (N_3973,N_3811,N_3886);
and U3974 (N_3974,N_3857,N_3839);
or U3975 (N_3975,N_3881,N_3893);
or U3976 (N_3976,N_3851,N_3810);
xor U3977 (N_3977,N_3820,N_3899);
nand U3978 (N_3978,N_3812,N_3894);
or U3979 (N_3979,N_3816,N_3860);
or U3980 (N_3980,N_3820,N_3801);
xor U3981 (N_3981,N_3815,N_3814);
or U3982 (N_3982,N_3849,N_3872);
and U3983 (N_3983,N_3829,N_3815);
nand U3984 (N_3984,N_3858,N_3862);
nor U3985 (N_3985,N_3867,N_3869);
or U3986 (N_3986,N_3883,N_3863);
nand U3987 (N_3987,N_3868,N_3895);
nor U3988 (N_3988,N_3809,N_3819);
nor U3989 (N_3989,N_3867,N_3878);
nor U3990 (N_3990,N_3866,N_3843);
nor U3991 (N_3991,N_3833,N_3828);
nor U3992 (N_3992,N_3843,N_3840);
and U3993 (N_3993,N_3815,N_3808);
nand U3994 (N_3994,N_3835,N_3877);
xor U3995 (N_3995,N_3856,N_3877);
and U3996 (N_3996,N_3824,N_3843);
and U3997 (N_3997,N_3834,N_3870);
nor U3998 (N_3998,N_3884,N_3879);
nor U3999 (N_3999,N_3823,N_3835);
or U4000 (N_4000,N_3970,N_3904);
or U4001 (N_4001,N_3960,N_3958);
nand U4002 (N_4002,N_3988,N_3916);
xnor U4003 (N_4003,N_3962,N_3964);
and U4004 (N_4004,N_3972,N_3997);
or U4005 (N_4005,N_3947,N_3941);
or U4006 (N_4006,N_3996,N_3967);
nor U4007 (N_4007,N_3939,N_3991);
and U4008 (N_4008,N_3987,N_3952);
or U4009 (N_4009,N_3909,N_3930);
nor U4010 (N_4010,N_3977,N_3974);
xor U4011 (N_4011,N_3900,N_3995);
nor U4012 (N_4012,N_3968,N_3918);
or U4013 (N_4013,N_3951,N_3901);
nor U4014 (N_4014,N_3902,N_3907);
and U4015 (N_4015,N_3973,N_3926);
xor U4016 (N_4016,N_3966,N_3905);
nand U4017 (N_4017,N_3961,N_3911);
nand U4018 (N_4018,N_3903,N_3913);
and U4019 (N_4019,N_3910,N_3969);
nor U4020 (N_4020,N_3982,N_3917);
nand U4021 (N_4021,N_3983,N_3971);
nand U4022 (N_4022,N_3993,N_3986);
nand U4023 (N_4023,N_3938,N_3906);
and U4024 (N_4024,N_3950,N_3925);
or U4025 (N_4025,N_3985,N_3989);
nand U4026 (N_4026,N_3933,N_3934);
nor U4027 (N_4027,N_3949,N_3979);
nand U4028 (N_4028,N_3990,N_3924);
nor U4029 (N_4029,N_3944,N_3945);
nand U4030 (N_4030,N_3957,N_3942);
or U4031 (N_4031,N_3992,N_3922);
and U4032 (N_4032,N_3959,N_3954);
or U4033 (N_4033,N_3932,N_3928);
or U4034 (N_4034,N_3963,N_3931);
or U4035 (N_4035,N_3935,N_3965);
or U4036 (N_4036,N_3981,N_3937);
nor U4037 (N_4037,N_3999,N_3955);
and U4038 (N_4038,N_3912,N_3921);
nand U4039 (N_4039,N_3998,N_3920);
nand U4040 (N_4040,N_3943,N_3946);
and U4041 (N_4041,N_3914,N_3976);
nand U4042 (N_4042,N_3956,N_3940);
nand U4043 (N_4043,N_3980,N_3919);
and U4044 (N_4044,N_3978,N_3994);
and U4045 (N_4045,N_3929,N_3923);
nand U4046 (N_4046,N_3915,N_3936);
or U4047 (N_4047,N_3984,N_3948);
or U4048 (N_4048,N_3975,N_3908);
nand U4049 (N_4049,N_3953,N_3927);
nor U4050 (N_4050,N_3998,N_3915);
and U4051 (N_4051,N_3917,N_3926);
or U4052 (N_4052,N_3954,N_3910);
nor U4053 (N_4053,N_3908,N_3918);
and U4054 (N_4054,N_3928,N_3926);
nor U4055 (N_4055,N_3916,N_3961);
nand U4056 (N_4056,N_3915,N_3913);
nand U4057 (N_4057,N_3914,N_3911);
and U4058 (N_4058,N_3913,N_3982);
nand U4059 (N_4059,N_3995,N_3989);
or U4060 (N_4060,N_3953,N_3969);
and U4061 (N_4061,N_3931,N_3949);
and U4062 (N_4062,N_3959,N_3947);
and U4063 (N_4063,N_3924,N_3914);
or U4064 (N_4064,N_3908,N_3904);
nand U4065 (N_4065,N_3984,N_3957);
nand U4066 (N_4066,N_3976,N_3977);
nor U4067 (N_4067,N_3936,N_3971);
and U4068 (N_4068,N_3941,N_3987);
nor U4069 (N_4069,N_3950,N_3911);
or U4070 (N_4070,N_3952,N_3968);
or U4071 (N_4071,N_3909,N_3976);
xnor U4072 (N_4072,N_3937,N_3912);
nand U4073 (N_4073,N_3904,N_3935);
or U4074 (N_4074,N_3942,N_3909);
nor U4075 (N_4075,N_3901,N_3997);
or U4076 (N_4076,N_3945,N_3979);
xnor U4077 (N_4077,N_3919,N_3990);
or U4078 (N_4078,N_3921,N_3918);
nand U4079 (N_4079,N_3922,N_3968);
nor U4080 (N_4080,N_3981,N_3952);
nor U4081 (N_4081,N_3982,N_3962);
or U4082 (N_4082,N_3963,N_3905);
nor U4083 (N_4083,N_3925,N_3961);
or U4084 (N_4084,N_3954,N_3991);
or U4085 (N_4085,N_3962,N_3950);
nand U4086 (N_4086,N_3966,N_3996);
and U4087 (N_4087,N_3923,N_3944);
and U4088 (N_4088,N_3934,N_3971);
nor U4089 (N_4089,N_3938,N_3973);
and U4090 (N_4090,N_3927,N_3950);
and U4091 (N_4091,N_3944,N_3991);
or U4092 (N_4092,N_3927,N_3904);
nand U4093 (N_4093,N_3932,N_3917);
xnor U4094 (N_4094,N_3972,N_3994);
nor U4095 (N_4095,N_3983,N_3901);
nor U4096 (N_4096,N_3914,N_3917);
nor U4097 (N_4097,N_3941,N_3986);
nand U4098 (N_4098,N_3900,N_3921);
and U4099 (N_4099,N_3977,N_3999);
or U4100 (N_4100,N_4095,N_4003);
nor U4101 (N_4101,N_4000,N_4050);
and U4102 (N_4102,N_4075,N_4091);
nand U4103 (N_4103,N_4073,N_4042);
or U4104 (N_4104,N_4015,N_4052);
or U4105 (N_4105,N_4069,N_4011);
nand U4106 (N_4106,N_4006,N_4020);
nor U4107 (N_4107,N_4013,N_4096);
or U4108 (N_4108,N_4059,N_4092);
and U4109 (N_4109,N_4061,N_4007);
nor U4110 (N_4110,N_4043,N_4025);
nand U4111 (N_4111,N_4099,N_4037);
nor U4112 (N_4112,N_4082,N_4068);
xnor U4113 (N_4113,N_4019,N_4034);
nor U4114 (N_4114,N_4097,N_4081);
or U4115 (N_4115,N_4077,N_4038);
nand U4116 (N_4116,N_4078,N_4039);
nand U4117 (N_4117,N_4004,N_4065);
nand U4118 (N_4118,N_4067,N_4014);
nor U4119 (N_4119,N_4089,N_4040);
nor U4120 (N_4120,N_4005,N_4098);
or U4121 (N_4121,N_4010,N_4046);
or U4122 (N_4122,N_4047,N_4060);
or U4123 (N_4123,N_4031,N_4035);
nand U4124 (N_4124,N_4063,N_4087);
nand U4125 (N_4125,N_4055,N_4066);
and U4126 (N_4126,N_4008,N_4083);
xor U4127 (N_4127,N_4079,N_4085);
nor U4128 (N_4128,N_4056,N_4002);
and U4129 (N_4129,N_4032,N_4026);
and U4130 (N_4130,N_4053,N_4074);
nand U4131 (N_4131,N_4051,N_4064);
nor U4132 (N_4132,N_4024,N_4045);
or U4133 (N_4133,N_4080,N_4057);
nor U4134 (N_4134,N_4029,N_4027);
nor U4135 (N_4135,N_4023,N_4017);
or U4136 (N_4136,N_4036,N_4054);
and U4137 (N_4137,N_4084,N_4041);
and U4138 (N_4138,N_4072,N_4030);
xor U4139 (N_4139,N_4062,N_4001);
and U4140 (N_4140,N_4070,N_4086);
nor U4141 (N_4141,N_4058,N_4093);
nand U4142 (N_4142,N_4049,N_4094);
or U4143 (N_4143,N_4071,N_4088);
nor U4144 (N_4144,N_4090,N_4018);
or U4145 (N_4145,N_4012,N_4028);
and U4146 (N_4146,N_4016,N_4033);
or U4147 (N_4147,N_4076,N_4044);
or U4148 (N_4148,N_4021,N_4009);
and U4149 (N_4149,N_4048,N_4022);
or U4150 (N_4150,N_4072,N_4016);
nor U4151 (N_4151,N_4085,N_4073);
and U4152 (N_4152,N_4099,N_4040);
or U4153 (N_4153,N_4033,N_4043);
nor U4154 (N_4154,N_4018,N_4017);
nand U4155 (N_4155,N_4006,N_4031);
xnor U4156 (N_4156,N_4000,N_4035);
or U4157 (N_4157,N_4022,N_4066);
nand U4158 (N_4158,N_4081,N_4071);
xnor U4159 (N_4159,N_4098,N_4068);
or U4160 (N_4160,N_4008,N_4023);
nand U4161 (N_4161,N_4082,N_4011);
or U4162 (N_4162,N_4090,N_4084);
nand U4163 (N_4163,N_4033,N_4060);
and U4164 (N_4164,N_4035,N_4071);
nor U4165 (N_4165,N_4009,N_4068);
and U4166 (N_4166,N_4057,N_4046);
or U4167 (N_4167,N_4096,N_4054);
or U4168 (N_4168,N_4047,N_4001);
and U4169 (N_4169,N_4028,N_4083);
nor U4170 (N_4170,N_4048,N_4007);
and U4171 (N_4171,N_4070,N_4054);
and U4172 (N_4172,N_4011,N_4003);
nor U4173 (N_4173,N_4021,N_4000);
nor U4174 (N_4174,N_4098,N_4051);
nor U4175 (N_4175,N_4061,N_4095);
nand U4176 (N_4176,N_4012,N_4080);
nand U4177 (N_4177,N_4083,N_4030);
or U4178 (N_4178,N_4015,N_4059);
nor U4179 (N_4179,N_4021,N_4046);
or U4180 (N_4180,N_4081,N_4078);
or U4181 (N_4181,N_4048,N_4002);
and U4182 (N_4182,N_4056,N_4008);
and U4183 (N_4183,N_4092,N_4075);
nor U4184 (N_4184,N_4067,N_4008);
nor U4185 (N_4185,N_4002,N_4037);
or U4186 (N_4186,N_4002,N_4051);
or U4187 (N_4187,N_4033,N_4014);
or U4188 (N_4188,N_4099,N_4043);
nor U4189 (N_4189,N_4003,N_4064);
nor U4190 (N_4190,N_4058,N_4051);
xnor U4191 (N_4191,N_4049,N_4018);
and U4192 (N_4192,N_4066,N_4051);
or U4193 (N_4193,N_4086,N_4037);
or U4194 (N_4194,N_4005,N_4062);
or U4195 (N_4195,N_4085,N_4016);
xnor U4196 (N_4196,N_4050,N_4056);
or U4197 (N_4197,N_4084,N_4074);
nor U4198 (N_4198,N_4062,N_4003);
nor U4199 (N_4199,N_4022,N_4083);
nor U4200 (N_4200,N_4116,N_4155);
and U4201 (N_4201,N_4184,N_4127);
or U4202 (N_4202,N_4190,N_4168);
and U4203 (N_4203,N_4199,N_4162);
or U4204 (N_4204,N_4181,N_4171);
nand U4205 (N_4205,N_4120,N_4180);
and U4206 (N_4206,N_4132,N_4124);
and U4207 (N_4207,N_4123,N_4117);
xnor U4208 (N_4208,N_4144,N_4154);
nor U4209 (N_4209,N_4156,N_4153);
or U4210 (N_4210,N_4142,N_4119);
nor U4211 (N_4211,N_4126,N_4136);
or U4212 (N_4212,N_4129,N_4186);
nand U4213 (N_4213,N_4170,N_4189);
and U4214 (N_4214,N_4161,N_4130);
and U4215 (N_4215,N_4100,N_4106);
xor U4216 (N_4216,N_4179,N_4118);
nand U4217 (N_4217,N_4112,N_4158);
xnor U4218 (N_4218,N_4128,N_4141);
nand U4219 (N_4219,N_4188,N_4147);
and U4220 (N_4220,N_4148,N_4145);
or U4221 (N_4221,N_4164,N_4177);
nor U4222 (N_4222,N_4185,N_4139);
and U4223 (N_4223,N_4122,N_4163);
nand U4224 (N_4224,N_4134,N_4173);
or U4225 (N_4225,N_4103,N_4101);
and U4226 (N_4226,N_4193,N_4110);
nor U4227 (N_4227,N_4135,N_4146);
nor U4228 (N_4228,N_4104,N_4157);
or U4229 (N_4229,N_4131,N_4196);
nand U4230 (N_4230,N_4111,N_4140);
xor U4231 (N_4231,N_4176,N_4195);
nor U4232 (N_4232,N_4178,N_4143);
nand U4233 (N_4233,N_4125,N_4197);
xor U4234 (N_4234,N_4182,N_4160);
or U4235 (N_4235,N_4183,N_4107);
nand U4236 (N_4236,N_4121,N_4152);
and U4237 (N_4237,N_4174,N_4138);
and U4238 (N_4238,N_4137,N_4167);
xor U4239 (N_4239,N_4192,N_4187);
xor U4240 (N_4240,N_4115,N_4105);
nand U4241 (N_4241,N_4165,N_4149);
nor U4242 (N_4242,N_4102,N_4109);
nor U4243 (N_4243,N_4151,N_4175);
or U4244 (N_4244,N_4194,N_4150);
or U4245 (N_4245,N_4114,N_4133);
and U4246 (N_4246,N_4159,N_4172);
nor U4247 (N_4247,N_4191,N_4108);
and U4248 (N_4248,N_4166,N_4169);
nor U4249 (N_4249,N_4113,N_4198);
or U4250 (N_4250,N_4169,N_4189);
nor U4251 (N_4251,N_4129,N_4174);
nor U4252 (N_4252,N_4165,N_4130);
xor U4253 (N_4253,N_4160,N_4116);
and U4254 (N_4254,N_4109,N_4178);
nor U4255 (N_4255,N_4182,N_4162);
or U4256 (N_4256,N_4127,N_4131);
nor U4257 (N_4257,N_4163,N_4197);
nand U4258 (N_4258,N_4106,N_4184);
and U4259 (N_4259,N_4177,N_4135);
or U4260 (N_4260,N_4160,N_4156);
or U4261 (N_4261,N_4184,N_4194);
nor U4262 (N_4262,N_4182,N_4169);
nor U4263 (N_4263,N_4158,N_4188);
and U4264 (N_4264,N_4125,N_4127);
nor U4265 (N_4265,N_4163,N_4175);
nand U4266 (N_4266,N_4154,N_4100);
and U4267 (N_4267,N_4138,N_4107);
nand U4268 (N_4268,N_4147,N_4172);
nand U4269 (N_4269,N_4178,N_4108);
nor U4270 (N_4270,N_4141,N_4134);
nand U4271 (N_4271,N_4140,N_4187);
or U4272 (N_4272,N_4153,N_4180);
nor U4273 (N_4273,N_4197,N_4141);
or U4274 (N_4274,N_4123,N_4113);
or U4275 (N_4275,N_4150,N_4198);
nor U4276 (N_4276,N_4192,N_4128);
and U4277 (N_4277,N_4172,N_4136);
nand U4278 (N_4278,N_4171,N_4175);
nor U4279 (N_4279,N_4169,N_4175);
nand U4280 (N_4280,N_4126,N_4104);
nand U4281 (N_4281,N_4183,N_4149);
or U4282 (N_4282,N_4103,N_4111);
or U4283 (N_4283,N_4124,N_4135);
nand U4284 (N_4284,N_4121,N_4183);
nand U4285 (N_4285,N_4184,N_4185);
or U4286 (N_4286,N_4114,N_4173);
nand U4287 (N_4287,N_4155,N_4103);
nand U4288 (N_4288,N_4182,N_4163);
or U4289 (N_4289,N_4126,N_4155);
and U4290 (N_4290,N_4114,N_4163);
or U4291 (N_4291,N_4100,N_4111);
or U4292 (N_4292,N_4126,N_4184);
nand U4293 (N_4293,N_4110,N_4120);
xnor U4294 (N_4294,N_4166,N_4103);
xor U4295 (N_4295,N_4150,N_4162);
nor U4296 (N_4296,N_4130,N_4123);
xor U4297 (N_4297,N_4131,N_4181);
nand U4298 (N_4298,N_4151,N_4119);
nand U4299 (N_4299,N_4127,N_4140);
xnor U4300 (N_4300,N_4262,N_4250);
or U4301 (N_4301,N_4239,N_4248);
and U4302 (N_4302,N_4297,N_4260);
or U4303 (N_4303,N_4264,N_4235);
or U4304 (N_4304,N_4233,N_4225);
or U4305 (N_4305,N_4200,N_4237);
nand U4306 (N_4306,N_4280,N_4221);
nand U4307 (N_4307,N_4211,N_4266);
or U4308 (N_4308,N_4257,N_4204);
nor U4309 (N_4309,N_4228,N_4267);
and U4310 (N_4310,N_4271,N_4278);
and U4311 (N_4311,N_4244,N_4254);
xor U4312 (N_4312,N_4238,N_4294);
or U4313 (N_4313,N_4287,N_4212);
and U4314 (N_4314,N_4256,N_4296);
nor U4315 (N_4315,N_4279,N_4202);
and U4316 (N_4316,N_4243,N_4213);
and U4317 (N_4317,N_4298,N_4208);
nand U4318 (N_4318,N_4290,N_4240);
and U4319 (N_4319,N_4283,N_4247);
nand U4320 (N_4320,N_4215,N_4285);
and U4321 (N_4321,N_4273,N_4242);
nand U4322 (N_4322,N_4268,N_4288);
nor U4323 (N_4323,N_4253,N_4209);
nand U4324 (N_4324,N_4207,N_4203);
and U4325 (N_4325,N_4226,N_4276);
nand U4326 (N_4326,N_4214,N_4249);
nand U4327 (N_4327,N_4231,N_4261);
nand U4328 (N_4328,N_4246,N_4265);
or U4329 (N_4329,N_4222,N_4245);
nand U4330 (N_4330,N_4227,N_4216);
nand U4331 (N_4331,N_4223,N_4259);
nor U4332 (N_4332,N_4201,N_4274);
nor U4333 (N_4333,N_4289,N_4299);
and U4334 (N_4334,N_4277,N_4281);
nor U4335 (N_4335,N_4210,N_4269);
xor U4336 (N_4336,N_4206,N_4284);
and U4337 (N_4337,N_4230,N_4293);
nor U4338 (N_4338,N_4205,N_4236);
and U4339 (N_4339,N_4251,N_4282);
nor U4340 (N_4340,N_4258,N_4275);
and U4341 (N_4341,N_4218,N_4291);
or U4342 (N_4342,N_4255,N_4229);
or U4343 (N_4343,N_4224,N_4232);
xnor U4344 (N_4344,N_4295,N_4252);
and U4345 (N_4345,N_4270,N_4217);
or U4346 (N_4346,N_4219,N_4241);
and U4347 (N_4347,N_4292,N_4272);
nand U4348 (N_4348,N_4263,N_4286);
or U4349 (N_4349,N_4234,N_4220);
and U4350 (N_4350,N_4273,N_4275);
and U4351 (N_4351,N_4233,N_4262);
or U4352 (N_4352,N_4266,N_4243);
nor U4353 (N_4353,N_4203,N_4228);
nor U4354 (N_4354,N_4212,N_4242);
or U4355 (N_4355,N_4240,N_4280);
nor U4356 (N_4356,N_4222,N_4253);
or U4357 (N_4357,N_4252,N_4249);
nor U4358 (N_4358,N_4259,N_4296);
or U4359 (N_4359,N_4232,N_4278);
nor U4360 (N_4360,N_4252,N_4230);
nand U4361 (N_4361,N_4271,N_4282);
nor U4362 (N_4362,N_4215,N_4202);
nand U4363 (N_4363,N_4292,N_4204);
and U4364 (N_4364,N_4231,N_4296);
nand U4365 (N_4365,N_4205,N_4269);
or U4366 (N_4366,N_4242,N_4262);
nor U4367 (N_4367,N_4250,N_4226);
nand U4368 (N_4368,N_4220,N_4210);
nor U4369 (N_4369,N_4276,N_4261);
nor U4370 (N_4370,N_4227,N_4289);
nor U4371 (N_4371,N_4205,N_4221);
nor U4372 (N_4372,N_4208,N_4219);
xnor U4373 (N_4373,N_4222,N_4280);
nand U4374 (N_4374,N_4293,N_4251);
nor U4375 (N_4375,N_4200,N_4236);
nor U4376 (N_4376,N_4200,N_4268);
nor U4377 (N_4377,N_4205,N_4287);
or U4378 (N_4378,N_4258,N_4274);
or U4379 (N_4379,N_4293,N_4292);
xor U4380 (N_4380,N_4261,N_4299);
or U4381 (N_4381,N_4267,N_4246);
and U4382 (N_4382,N_4218,N_4262);
or U4383 (N_4383,N_4256,N_4250);
and U4384 (N_4384,N_4203,N_4233);
nor U4385 (N_4385,N_4252,N_4203);
and U4386 (N_4386,N_4269,N_4232);
or U4387 (N_4387,N_4233,N_4230);
and U4388 (N_4388,N_4225,N_4227);
nor U4389 (N_4389,N_4224,N_4239);
nor U4390 (N_4390,N_4229,N_4245);
and U4391 (N_4391,N_4226,N_4225);
or U4392 (N_4392,N_4274,N_4231);
nand U4393 (N_4393,N_4203,N_4223);
xnor U4394 (N_4394,N_4253,N_4269);
xor U4395 (N_4395,N_4208,N_4215);
and U4396 (N_4396,N_4220,N_4291);
nand U4397 (N_4397,N_4278,N_4216);
or U4398 (N_4398,N_4243,N_4219);
and U4399 (N_4399,N_4206,N_4289);
and U4400 (N_4400,N_4307,N_4316);
nor U4401 (N_4401,N_4380,N_4387);
nor U4402 (N_4402,N_4328,N_4326);
or U4403 (N_4403,N_4314,N_4365);
nand U4404 (N_4404,N_4376,N_4395);
nor U4405 (N_4405,N_4330,N_4321);
or U4406 (N_4406,N_4350,N_4397);
nand U4407 (N_4407,N_4324,N_4373);
nor U4408 (N_4408,N_4339,N_4318);
nand U4409 (N_4409,N_4309,N_4305);
xor U4410 (N_4410,N_4356,N_4302);
xor U4411 (N_4411,N_4379,N_4371);
or U4412 (N_4412,N_4312,N_4319);
nor U4413 (N_4413,N_4332,N_4331);
and U4414 (N_4414,N_4337,N_4362);
xor U4415 (N_4415,N_4363,N_4375);
and U4416 (N_4416,N_4349,N_4391);
nand U4417 (N_4417,N_4392,N_4308);
or U4418 (N_4418,N_4357,N_4334);
nor U4419 (N_4419,N_4398,N_4353);
nand U4420 (N_4420,N_4341,N_4385);
nand U4421 (N_4421,N_4369,N_4399);
and U4422 (N_4422,N_4390,N_4370);
nor U4423 (N_4423,N_4364,N_4344);
nor U4424 (N_4424,N_4320,N_4327);
and U4425 (N_4425,N_4381,N_4315);
nor U4426 (N_4426,N_4342,N_4359);
nand U4427 (N_4427,N_4368,N_4393);
nor U4428 (N_4428,N_4306,N_4358);
and U4429 (N_4429,N_4384,N_4313);
or U4430 (N_4430,N_4347,N_4354);
nor U4431 (N_4431,N_4300,N_4396);
xnor U4432 (N_4432,N_4335,N_4345);
or U4433 (N_4433,N_4325,N_4333);
xnor U4434 (N_4434,N_4322,N_4311);
nand U4435 (N_4435,N_4352,N_4372);
nor U4436 (N_4436,N_4377,N_4338);
nand U4437 (N_4437,N_4389,N_4303);
and U4438 (N_4438,N_4323,N_4388);
xnor U4439 (N_4439,N_4348,N_4351);
nor U4440 (N_4440,N_4367,N_4355);
nand U4441 (N_4441,N_4340,N_4378);
nand U4442 (N_4442,N_4343,N_4301);
or U4443 (N_4443,N_4336,N_4382);
nand U4444 (N_4444,N_4329,N_4366);
nor U4445 (N_4445,N_4361,N_4346);
nor U4446 (N_4446,N_4374,N_4304);
nand U4447 (N_4447,N_4383,N_4317);
nand U4448 (N_4448,N_4310,N_4394);
nor U4449 (N_4449,N_4386,N_4360);
or U4450 (N_4450,N_4355,N_4358);
and U4451 (N_4451,N_4336,N_4368);
or U4452 (N_4452,N_4383,N_4324);
or U4453 (N_4453,N_4393,N_4316);
nor U4454 (N_4454,N_4324,N_4312);
xor U4455 (N_4455,N_4358,N_4357);
and U4456 (N_4456,N_4385,N_4334);
nand U4457 (N_4457,N_4306,N_4347);
or U4458 (N_4458,N_4326,N_4381);
or U4459 (N_4459,N_4344,N_4351);
xor U4460 (N_4460,N_4311,N_4391);
and U4461 (N_4461,N_4336,N_4390);
nor U4462 (N_4462,N_4379,N_4311);
nor U4463 (N_4463,N_4397,N_4303);
or U4464 (N_4464,N_4315,N_4300);
nor U4465 (N_4465,N_4385,N_4360);
nand U4466 (N_4466,N_4346,N_4340);
nor U4467 (N_4467,N_4303,N_4326);
xnor U4468 (N_4468,N_4399,N_4339);
nand U4469 (N_4469,N_4336,N_4379);
nand U4470 (N_4470,N_4313,N_4307);
nand U4471 (N_4471,N_4361,N_4333);
or U4472 (N_4472,N_4318,N_4321);
nor U4473 (N_4473,N_4306,N_4384);
nand U4474 (N_4474,N_4306,N_4359);
nand U4475 (N_4475,N_4387,N_4338);
nand U4476 (N_4476,N_4357,N_4309);
nor U4477 (N_4477,N_4308,N_4337);
or U4478 (N_4478,N_4350,N_4371);
nand U4479 (N_4479,N_4386,N_4369);
and U4480 (N_4480,N_4342,N_4331);
nand U4481 (N_4481,N_4383,N_4303);
nor U4482 (N_4482,N_4360,N_4361);
and U4483 (N_4483,N_4365,N_4379);
and U4484 (N_4484,N_4388,N_4376);
nand U4485 (N_4485,N_4359,N_4349);
and U4486 (N_4486,N_4342,N_4384);
nand U4487 (N_4487,N_4370,N_4353);
and U4488 (N_4488,N_4372,N_4394);
nor U4489 (N_4489,N_4388,N_4309);
or U4490 (N_4490,N_4308,N_4354);
nand U4491 (N_4491,N_4394,N_4338);
or U4492 (N_4492,N_4349,N_4332);
and U4493 (N_4493,N_4383,N_4363);
nor U4494 (N_4494,N_4366,N_4312);
xor U4495 (N_4495,N_4314,N_4350);
and U4496 (N_4496,N_4340,N_4319);
and U4497 (N_4497,N_4351,N_4364);
nor U4498 (N_4498,N_4301,N_4361);
nor U4499 (N_4499,N_4395,N_4382);
or U4500 (N_4500,N_4482,N_4423);
nor U4501 (N_4501,N_4420,N_4443);
or U4502 (N_4502,N_4469,N_4434);
and U4503 (N_4503,N_4460,N_4444);
or U4504 (N_4504,N_4494,N_4435);
nor U4505 (N_4505,N_4419,N_4411);
nor U4506 (N_4506,N_4456,N_4436);
nor U4507 (N_4507,N_4474,N_4426);
and U4508 (N_4508,N_4492,N_4413);
and U4509 (N_4509,N_4466,N_4414);
nor U4510 (N_4510,N_4446,N_4430);
nor U4511 (N_4511,N_4491,N_4433);
xor U4512 (N_4512,N_4402,N_4484);
and U4513 (N_4513,N_4406,N_4429);
nor U4514 (N_4514,N_4478,N_4459);
nand U4515 (N_4515,N_4432,N_4452);
nand U4516 (N_4516,N_4496,N_4403);
or U4517 (N_4517,N_4412,N_4417);
nor U4518 (N_4518,N_4464,N_4497);
or U4519 (N_4519,N_4472,N_4455);
or U4520 (N_4520,N_4454,N_4408);
nor U4521 (N_4521,N_4467,N_4441);
nand U4522 (N_4522,N_4415,N_4495);
or U4523 (N_4523,N_4489,N_4439);
and U4524 (N_4524,N_4475,N_4471);
or U4525 (N_4525,N_4404,N_4410);
or U4526 (N_4526,N_4401,N_4445);
and U4527 (N_4527,N_4425,N_4493);
nor U4528 (N_4528,N_4465,N_4463);
xnor U4529 (N_4529,N_4447,N_4450);
nor U4530 (N_4530,N_4473,N_4424);
nand U4531 (N_4531,N_4431,N_4461);
nor U4532 (N_4532,N_4485,N_4437);
nor U4533 (N_4533,N_4486,N_4488);
and U4534 (N_4534,N_4462,N_4453);
xor U4535 (N_4535,N_4418,N_4449);
nand U4536 (N_4536,N_4407,N_4487);
or U4537 (N_4537,N_4483,N_4490);
nand U4538 (N_4538,N_4442,N_4468);
and U4539 (N_4539,N_4499,N_4421);
and U4540 (N_4540,N_4451,N_4409);
xor U4541 (N_4541,N_4479,N_4457);
nand U4542 (N_4542,N_4480,N_4427);
xnor U4543 (N_4543,N_4458,N_4470);
xor U4544 (N_4544,N_4498,N_4438);
and U4545 (N_4545,N_4476,N_4400);
or U4546 (N_4546,N_4405,N_4422);
and U4547 (N_4547,N_4481,N_4477);
nand U4548 (N_4548,N_4440,N_4428);
nand U4549 (N_4549,N_4416,N_4448);
and U4550 (N_4550,N_4483,N_4405);
nor U4551 (N_4551,N_4461,N_4432);
and U4552 (N_4552,N_4456,N_4466);
nor U4553 (N_4553,N_4450,N_4454);
nand U4554 (N_4554,N_4427,N_4453);
and U4555 (N_4555,N_4452,N_4482);
nand U4556 (N_4556,N_4475,N_4451);
nor U4557 (N_4557,N_4449,N_4496);
nor U4558 (N_4558,N_4407,N_4473);
and U4559 (N_4559,N_4400,N_4487);
nor U4560 (N_4560,N_4402,N_4475);
nand U4561 (N_4561,N_4464,N_4460);
or U4562 (N_4562,N_4431,N_4432);
and U4563 (N_4563,N_4411,N_4431);
nor U4564 (N_4564,N_4436,N_4471);
or U4565 (N_4565,N_4463,N_4453);
nor U4566 (N_4566,N_4495,N_4454);
nand U4567 (N_4567,N_4484,N_4423);
and U4568 (N_4568,N_4415,N_4414);
nand U4569 (N_4569,N_4468,N_4406);
nand U4570 (N_4570,N_4448,N_4423);
and U4571 (N_4571,N_4422,N_4441);
or U4572 (N_4572,N_4423,N_4411);
nand U4573 (N_4573,N_4451,N_4408);
nor U4574 (N_4574,N_4428,N_4438);
or U4575 (N_4575,N_4449,N_4409);
nor U4576 (N_4576,N_4431,N_4414);
and U4577 (N_4577,N_4419,N_4461);
and U4578 (N_4578,N_4499,N_4445);
and U4579 (N_4579,N_4435,N_4473);
and U4580 (N_4580,N_4493,N_4478);
nor U4581 (N_4581,N_4448,N_4490);
or U4582 (N_4582,N_4434,N_4443);
nand U4583 (N_4583,N_4471,N_4461);
and U4584 (N_4584,N_4493,N_4443);
or U4585 (N_4585,N_4492,N_4424);
nor U4586 (N_4586,N_4436,N_4483);
nand U4587 (N_4587,N_4416,N_4409);
or U4588 (N_4588,N_4415,N_4457);
or U4589 (N_4589,N_4445,N_4454);
or U4590 (N_4590,N_4473,N_4419);
or U4591 (N_4591,N_4463,N_4483);
and U4592 (N_4592,N_4466,N_4432);
nand U4593 (N_4593,N_4406,N_4428);
nor U4594 (N_4594,N_4426,N_4486);
and U4595 (N_4595,N_4495,N_4440);
or U4596 (N_4596,N_4451,N_4419);
nand U4597 (N_4597,N_4415,N_4431);
nor U4598 (N_4598,N_4459,N_4466);
nor U4599 (N_4599,N_4434,N_4462);
nand U4600 (N_4600,N_4548,N_4598);
and U4601 (N_4601,N_4523,N_4534);
and U4602 (N_4602,N_4599,N_4539);
or U4603 (N_4603,N_4595,N_4527);
nand U4604 (N_4604,N_4545,N_4576);
and U4605 (N_4605,N_4565,N_4572);
nand U4606 (N_4606,N_4588,N_4537);
nand U4607 (N_4607,N_4538,N_4530);
nor U4608 (N_4608,N_4525,N_4524);
or U4609 (N_4609,N_4563,N_4560);
nand U4610 (N_4610,N_4581,N_4506);
nand U4611 (N_4611,N_4569,N_4533);
nand U4612 (N_4612,N_4573,N_4519);
nor U4613 (N_4613,N_4557,N_4567);
nand U4614 (N_4614,N_4587,N_4503);
nor U4615 (N_4615,N_4543,N_4551);
and U4616 (N_4616,N_4584,N_4509);
and U4617 (N_4617,N_4554,N_4580);
xor U4618 (N_4618,N_4561,N_4546);
xor U4619 (N_4619,N_4544,N_4583);
and U4620 (N_4620,N_4514,N_4516);
or U4621 (N_4621,N_4577,N_4555);
or U4622 (N_4622,N_4559,N_4591);
xnor U4623 (N_4623,N_4528,N_4589);
nor U4624 (N_4624,N_4507,N_4585);
nor U4625 (N_4625,N_4542,N_4536);
and U4626 (N_4626,N_4508,N_4579);
nor U4627 (N_4627,N_4556,N_4597);
and U4628 (N_4628,N_4526,N_4570);
nand U4629 (N_4629,N_4571,N_4531);
nand U4630 (N_4630,N_4521,N_4520);
or U4631 (N_4631,N_4593,N_4529);
or U4632 (N_4632,N_4590,N_4541);
or U4633 (N_4633,N_4512,N_4535);
xor U4634 (N_4634,N_4566,N_4574);
and U4635 (N_4635,N_4594,N_4501);
nand U4636 (N_4636,N_4517,N_4552);
nand U4637 (N_4637,N_4547,N_4500);
nand U4638 (N_4638,N_4592,N_4511);
or U4639 (N_4639,N_4515,N_4596);
nor U4640 (N_4640,N_4522,N_4532);
nand U4641 (N_4641,N_4513,N_4558);
xor U4642 (N_4642,N_4582,N_4504);
nand U4643 (N_4643,N_4578,N_4553);
nand U4644 (N_4644,N_4540,N_4510);
nand U4645 (N_4645,N_4550,N_4518);
nor U4646 (N_4646,N_4568,N_4549);
nor U4647 (N_4647,N_4575,N_4564);
or U4648 (N_4648,N_4562,N_4505);
or U4649 (N_4649,N_4502,N_4586);
nand U4650 (N_4650,N_4500,N_4517);
or U4651 (N_4651,N_4586,N_4528);
nand U4652 (N_4652,N_4577,N_4535);
nand U4653 (N_4653,N_4508,N_4531);
or U4654 (N_4654,N_4534,N_4504);
or U4655 (N_4655,N_4530,N_4533);
nor U4656 (N_4656,N_4588,N_4560);
nand U4657 (N_4657,N_4504,N_4551);
or U4658 (N_4658,N_4522,N_4512);
nor U4659 (N_4659,N_4547,N_4566);
nand U4660 (N_4660,N_4530,N_4579);
nand U4661 (N_4661,N_4541,N_4528);
or U4662 (N_4662,N_4598,N_4557);
and U4663 (N_4663,N_4588,N_4567);
or U4664 (N_4664,N_4595,N_4534);
nand U4665 (N_4665,N_4519,N_4542);
and U4666 (N_4666,N_4572,N_4514);
nor U4667 (N_4667,N_4531,N_4592);
or U4668 (N_4668,N_4564,N_4531);
or U4669 (N_4669,N_4560,N_4554);
or U4670 (N_4670,N_4502,N_4513);
xor U4671 (N_4671,N_4506,N_4501);
and U4672 (N_4672,N_4512,N_4581);
or U4673 (N_4673,N_4519,N_4547);
and U4674 (N_4674,N_4577,N_4541);
nor U4675 (N_4675,N_4570,N_4544);
or U4676 (N_4676,N_4567,N_4583);
and U4677 (N_4677,N_4551,N_4506);
or U4678 (N_4678,N_4520,N_4500);
or U4679 (N_4679,N_4504,N_4515);
or U4680 (N_4680,N_4543,N_4579);
nand U4681 (N_4681,N_4502,N_4539);
and U4682 (N_4682,N_4551,N_4570);
xnor U4683 (N_4683,N_4577,N_4582);
nand U4684 (N_4684,N_4573,N_4595);
nand U4685 (N_4685,N_4505,N_4536);
and U4686 (N_4686,N_4537,N_4583);
nand U4687 (N_4687,N_4586,N_4530);
and U4688 (N_4688,N_4572,N_4524);
xor U4689 (N_4689,N_4577,N_4548);
xor U4690 (N_4690,N_4513,N_4501);
nand U4691 (N_4691,N_4524,N_4563);
and U4692 (N_4692,N_4520,N_4560);
nand U4693 (N_4693,N_4507,N_4595);
or U4694 (N_4694,N_4509,N_4533);
nand U4695 (N_4695,N_4506,N_4531);
and U4696 (N_4696,N_4561,N_4579);
and U4697 (N_4697,N_4502,N_4542);
xor U4698 (N_4698,N_4512,N_4504);
xnor U4699 (N_4699,N_4505,N_4540);
nand U4700 (N_4700,N_4614,N_4681);
nand U4701 (N_4701,N_4622,N_4625);
or U4702 (N_4702,N_4654,N_4632);
or U4703 (N_4703,N_4621,N_4666);
nand U4704 (N_4704,N_4601,N_4639);
nor U4705 (N_4705,N_4673,N_4641);
nor U4706 (N_4706,N_4652,N_4698);
nand U4707 (N_4707,N_4602,N_4611);
or U4708 (N_4708,N_4677,N_4695);
or U4709 (N_4709,N_4691,N_4645);
nor U4710 (N_4710,N_4649,N_4675);
nor U4711 (N_4711,N_4640,N_4676);
and U4712 (N_4712,N_4650,N_4637);
nand U4713 (N_4713,N_4628,N_4690);
nand U4714 (N_4714,N_4660,N_4656);
or U4715 (N_4715,N_4616,N_4635);
nor U4716 (N_4716,N_4629,N_4692);
and U4717 (N_4717,N_4647,N_4657);
nor U4718 (N_4718,N_4655,N_4683);
nand U4719 (N_4719,N_4617,N_4604);
nor U4720 (N_4720,N_4659,N_4638);
nor U4721 (N_4721,N_4618,N_4624);
nor U4722 (N_4722,N_4626,N_4615);
or U4723 (N_4723,N_4684,N_4669);
nand U4724 (N_4724,N_4658,N_4651);
nor U4725 (N_4725,N_4643,N_4610);
or U4726 (N_4726,N_4661,N_4633);
nand U4727 (N_4727,N_4646,N_4686);
and U4728 (N_4728,N_4697,N_4603);
and U4729 (N_4729,N_4674,N_4678);
and U4730 (N_4730,N_4620,N_4636);
nor U4731 (N_4731,N_4644,N_4672);
nor U4732 (N_4732,N_4679,N_4662);
xor U4733 (N_4733,N_4642,N_4613);
and U4734 (N_4734,N_4623,N_4653);
or U4735 (N_4735,N_4670,N_4663);
nor U4736 (N_4736,N_4612,N_4667);
or U4737 (N_4737,N_4607,N_4665);
nor U4738 (N_4738,N_4627,N_4689);
or U4739 (N_4739,N_4671,N_4606);
nor U4740 (N_4740,N_4619,N_4699);
nor U4741 (N_4741,N_4668,N_4694);
nand U4742 (N_4742,N_4680,N_4631);
nand U4743 (N_4743,N_4600,N_4648);
or U4744 (N_4744,N_4605,N_4609);
nor U4745 (N_4745,N_4630,N_4634);
or U4746 (N_4746,N_4685,N_4664);
nand U4747 (N_4747,N_4688,N_4682);
nor U4748 (N_4748,N_4687,N_4693);
or U4749 (N_4749,N_4696,N_4608);
nand U4750 (N_4750,N_4643,N_4644);
nor U4751 (N_4751,N_4658,N_4657);
nor U4752 (N_4752,N_4678,N_4665);
nor U4753 (N_4753,N_4687,N_4695);
nor U4754 (N_4754,N_4616,N_4625);
nand U4755 (N_4755,N_4658,N_4690);
nor U4756 (N_4756,N_4671,N_4673);
xor U4757 (N_4757,N_4669,N_4600);
and U4758 (N_4758,N_4655,N_4693);
and U4759 (N_4759,N_4606,N_4643);
nand U4760 (N_4760,N_4638,N_4657);
and U4761 (N_4761,N_4641,N_4633);
and U4762 (N_4762,N_4618,N_4684);
or U4763 (N_4763,N_4661,N_4698);
or U4764 (N_4764,N_4697,N_4676);
or U4765 (N_4765,N_4619,N_4615);
nand U4766 (N_4766,N_4608,N_4605);
and U4767 (N_4767,N_4663,N_4655);
nor U4768 (N_4768,N_4676,N_4678);
nand U4769 (N_4769,N_4630,N_4638);
xnor U4770 (N_4770,N_4663,N_4619);
nand U4771 (N_4771,N_4618,N_4687);
nand U4772 (N_4772,N_4696,N_4675);
nand U4773 (N_4773,N_4621,N_4635);
nand U4774 (N_4774,N_4694,N_4603);
and U4775 (N_4775,N_4686,N_4619);
nand U4776 (N_4776,N_4650,N_4652);
nand U4777 (N_4777,N_4663,N_4669);
nor U4778 (N_4778,N_4653,N_4649);
xor U4779 (N_4779,N_4664,N_4613);
or U4780 (N_4780,N_4619,N_4629);
and U4781 (N_4781,N_4623,N_4627);
nor U4782 (N_4782,N_4647,N_4665);
and U4783 (N_4783,N_4675,N_4671);
nand U4784 (N_4784,N_4605,N_4639);
and U4785 (N_4785,N_4660,N_4685);
and U4786 (N_4786,N_4648,N_4651);
nor U4787 (N_4787,N_4671,N_4622);
and U4788 (N_4788,N_4612,N_4665);
or U4789 (N_4789,N_4619,N_4641);
xnor U4790 (N_4790,N_4694,N_4692);
and U4791 (N_4791,N_4651,N_4601);
nand U4792 (N_4792,N_4671,N_4665);
nor U4793 (N_4793,N_4676,N_4605);
nor U4794 (N_4794,N_4633,N_4693);
nand U4795 (N_4795,N_4615,N_4611);
or U4796 (N_4796,N_4618,N_4615);
nor U4797 (N_4797,N_4641,N_4620);
and U4798 (N_4798,N_4669,N_4643);
nand U4799 (N_4799,N_4602,N_4650);
or U4800 (N_4800,N_4767,N_4783);
or U4801 (N_4801,N_4796,N_4714);
nand U4802 (N_4802,N_4736,N_4779);
nand U4803 (N_4803,N_4733,N_4772);
nand U4804 (N_4804,N_4732,N_4777);
or U4805 (N_4805,N_4780,N_4700);
or U4806 (N_4806,N_4715,N_4747);
and U4807 (N_4807,N_4795,N_4765);
nand U4808 (N_4808,N_4758,N_4737);
nor U4809 (N_4809,N_4768,N_4719);
or U4810 (N_4810,N_4790,N_4748);
nor U4811 (N_4811,N_4757,N_4721);
and U4812 (N_4812,N_4749,N_4708);
or U4813 (N_4813,N_4739,N_4750);
nand U4814 (N_4814,N_4741,N_4752);
and U4815 (N_4815,N_4735,N_4745);
nand U4816 (N_4816,N_4787,N_4717);
xor U4817 (N_4817,N_4794,N_4761);
xor U4818 (N_4818,N_4756,N_4724);
or U4819 (N_4819,N_4774,N_4769);
and U4820 (N_4820,N_4766,N_4778);
nor U4821 (N_4821,N_4771,N_4716);
nor U4822 (N_4822,N_4788,N_4799);
or U4823 (N_4823,N_4728,N_4722);
or U4824 (N_4824,N_4760,N_4707);
xnor U4825 (N_4825,N_4710,N_4781);
nor U4826 (N_4826,N_4743,N_4785);
nand U4827 (N_4827,N_4731,N_4711);
or U4828 (N_4828,N_4759,N_4720);
and U4829 (N_4829,N_4742,N_4763);
and U4830 (N_4830,N_4773,N_4704);
xnor U4831 (N_4831,N_4706,N_4726);
xnor U4832 (N_4832,N_4764,N_4753);
nor U4833 (N_4833,N_4730,N_4770);
and U4834 (N_4834,N_4725,N_4786);
nand U4835 (N_4835,N_4755,N_4709);
or U4836 (N_4836,N_4746,N_4776);
nor U4837 (N_4837,N_4727,N_4734);
and U4838 (N_4838,N_4738,N_4723);
and U4839 (N_4839,N_4791,N_4775);
xor U4840 (N_4840,N_4712,N_4789);
or U4841 (N_4841,N_4713,N_4782);
or U4842 (N_4842,N_4744,N_4762);
xnor U4843 (N_4843,N_4798,N_4792);
and U4844 (N_4844,N_4751,N_4718);
and U4845 (N_4845,N_4754,N_4793);
or U4846 (N_4846,N_4784,N_4740);
and U4847 (N_4847,N_4702,N_4729);
nand U4848 (N_4848,N_4703,N_4701);
or U4849 (N_4849,N_4705,N_4797);
or U4850 (N_4850,N_4735,N_4719);
and U4851 (N_4851,N_4719,N_4764);
and U4852 (N_4852,N_4748,N_4706);
nand U4853 (N_4853,N_4761,N_4732);
or U4854 (N_4854,N_4700,N_4784);
nor U4855 (N_4855,N_4782,N_4720);
or U4856 (N_4856,N_4744,N_4731);
nand U4857 (N_4857,N_4753,N_4706);
nor U4858 (N_4858,N_4711,N_4766);
and U4859 (N_4859,N_4747,N_4788);
and U4860 (N_4860,N_4781,N_4709);
xnor U4861 (N_4861,N_4776,N_4714);
nor U4862 (N_4862,N_4753,N_4711);
nand U4863 (N_4863,N_4746,N_4783);
and U4864 (N_4864,N_4727,N_4768);
nor U4865 (N_4865,N_4779,N_4702);
and U4866 (N_4866,N_4796,N_4705);
nor U4867 (N_4867,N_4700,N_4794);
xnor U4868 (N_4868,N_4778,N_4743);
and U4869 (N_4869,N_4711,N_4758);
or U4870 (N_4870,N_4759,N_4716);
or U4871 (N_4871,N_4761,N_4717);
nand U4872 (N_4872,N_4775,N_4795);
nor U4873 (N_4873,N_4731,N_4740);
or U4874 (N_4874,N_4758,N_4770);
or U4875 (N_4875,N_4717,N_4789);
nor U4876 (N_4876,N_4727,N_4741);
or U4877 (N_4877,N_4786,N_4751);
nand U4878 (N_4878,N_4764,N_4709);
nand U4879 (N_4879,N_4714,N_4708);
or U4880 (N_4880,N_4768,N_4777);
nor U4881 (N_4881,N_4783,N_4740);
or U4882 (N_4882,N_4786,N_4782);
or U4883 (N_4883,N_4790,N_4715);
and U4884 (N_4884,N_4710,N_4749);
xor U4885 (N_4885,N_4760,N_4797);
nand U4886 (N_4886,N_4759,N_4743);
or U4887 (N_4887,N_4749,N_4753);
and U4888 (N_4888,N_4776,N_4755);
or U4889 (N_4889,N_4722,N_4794);
or U4890 (N_4890,N_4745,N_4736);
nand U4891 (N_4891,N_4738,N_4735);
nor U4892 (N_4892,N_4760,N_4757);
or U4893 (N_4893,N_4700,N_4728);
and U4894 (N_4894,N_4748,N_4741);
xor U4895 (N_4895,N_4797,N_4772);
and U4896 (N_4896,N_4742,N_4799);
nand U4897 (N_4897,N_4794,N_4719);
xor U4898 (N_4898,N_4700,N_4733);
or U4899 (N_4899,N_4768,N_4772);
xnor U4900 (N_4900,N_4822,N_4848);
nand U4901 (N_4901,N_4837,N_4867);
and U4902 (N_4902,N_4895,N_4819);
nand U4903 (N_4903,N_4877,N_4879);
nor U4904 (N_4904,N_4857,N_4807);
or U4905 (N_4905,N_4804,N_4833);
and U4906 (N_4906,N_4881,N_4852);
and U4907 (N_4907,N_4893,N_4869);
nor U4908 (N_4908,N_4820,N_4875);
nand U4909 (N_4909,N_4878,N_4871);
nor U4910 (N_4910,N_4821,N_4889);
nor U4911 (N_4911,N_4884,N_4891);
nand U4912 (N_4912,N_4839,N_4854);
nand U4913 (N_4913,N_4800,N_4874);
xnor U4914 (N_4914,N_4817,N_4814);
nand U4915 (N_4915,N_4813,N_4898);
nor U4916 (N_4916,N_4843,N_4835);
nand U4917 (N_4917,N_4894,N_4825);
or U4918 (N_4918,N_4888,N_4860);
and U4919 (N_4919,N_4887,N_4886);
nand U4920 (N_4920,N_4834,N_4865);
or U4921 (N_4921,N_4851,N_4801);
or U4922 (N_4922,N_4832,N_4838);
nand U4923 (N_4923,N_4815,N_4880);
nor U4924 (N_4924,N_4830,N_4872);
nand U4925 (N_4925,N_4890,N_4840);
nor U4926 (N_4926,N_4808,N_4811);
nor U4927 (N_4927,N_4868,N_4803);
nand U4928 (N_4928,N_4850,N_4836);
nor U4929 (N_4929,N_4812,N_4847);
nor U4930 (N_4930,N_4856,N_4897);
nand U4931 (N_4931,N_4816,N_4883);
nor U4932 (N_4932,N_4846,N_4809);
nor U4933 (N_4933,N_4866,N_4802);
or U4934 (N_4934,N_4853,N_4896);
or U4935 (N_4935,N_4859,N_4805);
and U4936 (N_4936,N_4829,N_4845);
or U4937 (N_4937,N_4826,N_4849);
xnor U4938 (N_4938,N_4862,N_4873);
and U4939 (N_4939,N_4824,N_4818);
or U4940 (N_4940,N_4842,N_4823);
and U4941 (N_4941,N_4844,N_4892);
nor U4942 (N_4942,N_4806,N_4831);
xnor U4943 (N_4943,N_4870,N_4864);
or U4944 (N_4944,N_4858,N_4841);
nor U4945 (N_4945,N_4885,N_4863);
nor U4946 (N_4946,N_4827,N_4810);
or U4947 (N_4947,N_4828,N_4855);
xnor U4948 (N_4948,N_4882,N_4861);
and U4949 (N_4949,N_4899,N_4876);
and U4950 (N_4950,N_4812,N_4854);
xor U4951 (N_4951,N_4874,N_4868);
nor U4952 (N_4952,N_4816,N_4851);
and U4953 (N_4953,N_4892,N_4857);
nand U4954 (N_4954,N_4888,N_4845);
and U4955 (N_4955,N_4863,N_4873);
or U4956 (N_4956,N_4883,N_4807);
or U4957 (N_4957,N_4848,N_4814);
nor U4958 (N_4958,N_4827,N_4894);
or U4959 (N_4959,N_4829,N_4833);
and U4960 (N_4960,N_4850,N_4888);
or U4961 (N_4961,N_4846,N_4853);
xor U4962 (N_4962,N_4805,N_4860);
nand U4963 (N_4963,N_4809,N_4894);
and U4964 (N_4964,N_4890,N_4865);
nor U4965 (N_4965,N_4849,N_4890);
nor U4966 (N_4966,N_4881,N_4831);
xnor U4967 (N_4967,N_4840,N_4800);
and U4968 (N_4968,N_4872,N_4828);
or U4969 (N_4969,N_4841,N_4878);
or U4970 (N_4970,N_4801,N_4838);
or U4971 (N_4971,N_4883,N_4896);
or U4972 (N_4972,N_4882,N_4815);
xor U4973 (N_4973,N_4841,N_4821);
nand U4974 (N_4974,N_4840,N_4842);
or U4975 (N_4975,N_4803,N_4875);
or U4976 (N_4976,N_4800,N_4838);
or U4977 (N_4977,N_4805,N_4841);
nand U4978 (N_4978,N_4857,N_4898);
and U4979 (N_4979,N_4817,N_4888);
nand U4980 (N_4980,N_4850,N_4821);
or U4981 (N_4981,N_4824,N_4828);
nor U4982 (N_4982,N_4815,N_4806);
nor U4983 (N_4983,N_4826,N_4859);
xor U4984 (N_4984,N_4834,N_4881);
nand U4985 (N_4985,N_4868,N_4850);
nand U4986 (N_4986,N_4875,N_4879);
or U4987 (N_4987,N_4839,N_4833);
or U4988 (N_4988,N_4837,N_4874);
nor U4989 (N_4989,N_4851,N_4877);
xor U4990 (N_4990,N_4856,N_4862);
or U4991 (N_4991,N_4872,N_4854);
or U4992 (N_4992,N_4812,N_4894);
nand U4993 (N_4993,N_4899,N_4826);
nand U4994 (N_4994,N_4846,N_4880);
nor U4995 (N_4995,N_4891,N_4844);
nor U4996 (N_4996,N_4847,N_4827);
nand U4997 (N_4997,N_4894,N_4836);
nand U4998 (N_4998,N_4887,N_4839);
or U4999 (N_4999,N_4877,N_4866);
and UO_0 (O_0,N_4960,N_4938);
xor UO_1 (O_1,N_4976,N_4905);
nand UO_2 (O_2,N_4988,N_4926);
nor UO_3 (O_3,N_4996,N_4913);
or UO_4 (O_4,N_4921,N_4967);
and UO_5 (O_5,N_4994,N_4971);
nand UO_6 (O_6,N_4922,N_4950);
nor UO_7 (O_7,N_4982,N_4936);
nand UO_8 (O_8,N_4912,N_4991);
nand UO_9 (O_9,N_4984,N_4958);
and UO_10 (O_10,N_4906,N_4903);
xnor UO_11 (O_11,N_4917,N_4948);
or UO_12 (O_12,N_4920,N_4909);
nor UO_13 (O_13,N_4977,N_4992);
nand UO_14 (O_14,N_4980,N_4964);
or UO_15 (O_15,N_4955,N_4978);
nand UO_16 (O_16,N_4981,N_4914);
or UO_17 (O_17,N_4946,N_4933);
nor UO_18 (O_18,N_4911,N_4974);
or UO_19 (O_19,N_4987,N_4932);
nand UO_20 (O_20,N_4986,N_4900);
or UO_21 (O_21,N_4925,N_4910);
nand UO_22 (O_22,N_4953,N_4943);
nor UO_23 (O_23,N_4928,N_4939);
and UO_24 (O_24,N_4944,N_4985);
xnor UO_25 (O_25,N_4947,N_4952);
and UO_26 (O_26,N_4962,N_4957);
nor UO_27 (O_27,N_4918,N_4972);
and UO_28 (O_28,N_4924,N_4940);
nor UO_29 (O_29,N_4966,N_4989);
or UO_30 (O_30,N_4907,N_4915);
nand UO_31 (O_31,N_4908,N_4927);
xnor UO_32 (O_32,N_4951,N_4961);
or UO_33 (O_33,N_4937,N_4902);
or UO_34 (O_34,N_4923,N_4973);
nor UO_35 (O_35,N_4929,N_4945);
or UO_36 (O_36,N_4901,N_4931);
and UO_37 (O_37,N_4995,N_4965);
and UO_38 (O_38,N_4954,N_4979);
nand UO_39 (O_39,N_4963,N_4935);
or UO_40 (O_40,N_4999,N_4975);
and UO_41 (O_41,N_4916,N_4934);
or UO_42 (O_42,N_4969,N_4949);
xor UO_43 (O_43,N_4998,N_4956);
xnor UO_44 (O_44,N_4997,N_4968);
nand UO_45 (O_45,N_4959,N_4990);
nor UO_46 (O_46,N_4930,N_4993);
nor UO_47 (O_47,N_4919,N_4941);
or UO_48 (O_48,N_4942,N_4983);
or UO_49 (O_49,N_4970,N_4904);
nand UO_50 (O_50,N_4950,N_4945);
nand UO_51 (O_51,N_4952,N_4960);
or UO_52 (O_52,N_4995,N_4974);
and UO_53 (O_53,N_4953,N_4926);
xor UO_54 (O_54,N_4974,N_4948);
xnor UO_55 (O_55,N_4974,N_4968);
nand UO_56 (O_56,N_4910,N_4942);
xnor UO_57 (O_57,N_4918,N_4900);
and UO_58 (O_58,N_4987,N_4948);
or UO_59 (O_59,N_4938,N_4997);
nand UO_60 (O_60,N_4967,N_4995);
nor UO_61 (O_61,N_4940,N_4957);
and UO_62 (O_62,N_4944,N_4916);
nand UO_63 (O_63,N_4970,N_4999);
or UO_64 (O_64,N_4943,N_4907);
nor UO_65 (O_65,N_4969,N_4903);
or UO_66 (O_66,N_4913,N_4958);
nand UO_67 (O_67,N_4916,N_4920);
and UO_68 (O_68,N_4969,N_4910);
nor UO_69 (O_69,N_4941,N_4981);
nand UO_70 (O_70,N_4927,N_4947);
nor UO_71 (O_71,N_4939,N_4969);
xor UO_72 (O_72,N_4945,N_4997);
xnor UO_73 (O_73,N_4918,N_4902);
and UO_74 (O_74,N_4928,N_4947);
xor UO_75 (O_75,N_4991,N_4964);
nor UO_76 (O_76,N_4903,N_4993);
xor UO_77 (O_77,N_4913,N_4942);
and UO_78 (O_78,N_4965,N_4989);
xor UO_79 (O_79,N_4966,N_4936);
and UO_80 (O_80,N_4967,N_4982);
nor UO_81 (O_81,N_4997,N_4995);
and UO_82 (O_82,N_4900,N_4993);
nand UO_83 (O_83,N_4936,N_4961);
or UO_84 (O_84,N_4922,N_4910);
nand UO_85 (O_85,N_4961,N_4901);
nand UO_86 (O_86,N_4949,N_4993);
nor UO_87 (O_87,N_4989,N_4954);
nand UO_88 (O_88,N_4924,N_4949);
or UO_89 (O_89,N_4984,N_4975);
nand UO_90 (O_90,N_4907,N_4986);
nor UO_91 (O_91,N_4965,N_4922);
nand UO_92 (O_92,N_4970,N_4939);
nor UO_93 (O_93,N_4962,N_4949);
or UO_94 (O_94,N_4917,N_4971);
xor UO_95 (O_95,N_4998,N_4952);
and UO_96 (O_96,N_4935,N_4958);
nand UO_97 (O_97,N_4958,N_4962);
or UO_98 (O_98,N_4979,N_4996);
and UO_99 (O_99,N_4947,N_4963);
or UO_100 (O_100,N_4944,N_4918);
nor UO_101 (O_101,N_4939,N_4915);
xnor UO_102 (O_102,N_4946,N_4948);
nand UO_103 (O_103,N_4924,N_4906);
or UO_104 (O_104,N_4911,N_4952);
or UO_105 (O_105,N_4988,N_4999);
or UO_106 (O_106,N_4979,N_4959);
nand UO_107 (O_107,N_4933,N_4940);
or UO_108 (O_108,N_4917,N_4939);
xor UO_109 (O_109,N_4941,N_4959);
nand UO_110 (O_110,N_4959,N_4963);
xnor UO_111 (O_111,N_4912,N_4941);
nor UO_112 (O_112,N_4960,N_4962);
nand UO_113 (O_113,N_4905,N_4927);
or UO_114 (O_114,N_4960,N_4964);
or UO_115 (O_115,N_4958,N_4997);
or UO_116 (O_116,N_4919,N_4971);
nor UO_117 (O_117,N_4937,N_4907);
nand UO_118 (O_118,N_4922,N_4932);
or UO_119 (O_119,N_4960,N_4983);
nand UO_120 (O_120,N_4908,N_4975);
or UO_121 (O_121,N_4912,N_4948);
and UO_122 (O_122,N_4914,N_4972);
nor UO_123 (O_123,N_4913,N_4903);
nand UO_124 (O_124,N_4984,N_4942);
nand UO_125 (O_125,N_4983,N_4946);
nor UO_126 (O_126,N_4953,N_4971);
or UO_127 (O_127,N_4927,N_4942);
nor UO_128 (O_128,N_4989,N_4930);
nand UO_129 (O_129,N_4992,N_4991);
nand UO_130 (O_130,N_4916,N_4954);
and UO_131 (O_131,N_4927,N_4972);
nor UO_132 (O_132,N_4981,N_4954);
and UO_133 (O_133,N_4946,N_4936);
or UO_134 (O_134,N_4920,N_4936);
nor UO_135 (O_135,N_4926,N_4958);
nor UO_136 (O_136,N_4908,N_4943);
nand UO_137 (O_137,N_4922,N_4958);
and UO_138 (O_138,N_4936,N_4972);
or UO_139 (O_139,N_4996,N_4980);
nand UO_140 (O_140,N_4961,N_4977);
and UO_141 (O_141,N_4949,N_4937);
and UO_142 (O_142,N_4927,N_4910);
and UO_143 (O_143,N_4926,N_4996);
nor UO_144 (O_144,N_4997,N_4957);
nor UO_145 (O_145,N_4910,N_4957);
or UO_146 (O_146,N_4927,N_4940);
nand UO_147 (O_147,N_4933,N_4921);
or UO_148 (O_148,N_4965,N_4991);
nor UO_149 (O_149,N_4958,N_4945);
and UO_150 (O_150,N_4925,N_4957);
and UO_151 (O_151,N_4936,N_4937);
nand UO_152 (O_152,N_4969,N_4968);
nand UO_153 (O_153,N_4950,N_4971);
and UO_154 (O_154,N_4911,N_4903);
or UO_155 (O_155,N_4966,N_4977);
nand UO_156 (O_156,N_4980,N_4958);
or UO_157 (O_157,N_4933,N_4904);
and UO_158 (O_158,N_4950,N_4941);
or UO_159 (O_159,N_4988,N_4949);
and UO_160 (O_160,N_4952,N_4948);
nand UO_161 (O_161,N_4909,N_4979);
or UO_162 (O_162,N_4945,N_4991);
or UO_163 (O_163,N_4920,N_4928);
nor UO_164 (O_164,N_4991,N_4950);
xor UO_165 (O_165,N_4927,N_4952);
nor UO_166 (O_166,N_4930,N_4938);
and UO_167 (O_167,N_4968,N_4993);
nand UO_168 (O_168,N_4962,N_4945);
or UO_169 (O_169,N_4996,N_4945);
nand UO_170 (O_170,N_4905,N_4975);
nor UO_171 (O_171,N_4910,N_4984);
xor UO_172 (O_172,N_4926,N_4927);
and UO_173 (O_173,N_4921,N_4997);
or UO_174 (O_174,N_4929,N_4980);
or UO_175 (O_175,N_4958,N_4972);
nor UO_176 (O_176,N_4998,N_4915);
nand UO_177 (O_177,N_4903,N_4904);
or UO_178 (O_178,N_4992,N_4939);
or UO_179 (O_179,N_4971,N_4986);
nor UO_180 (O_180,N_4918,N_4937);
and UO_181 (O_181,N_4962,N_4940);
nand UO_182 (O_182,N_4967,N_4946);
or UO_183 (O_183,N_4903,N_4922);
nand UO_184 (O_184,N_4998,N_4962);
or UO_185 (O_185,N_4980,N_4902);
nor UO_186 (O_186,N_4994,N_4945);
nand UO_187 (O_187,N_4968,N_4930);
xnor UO_188 (O_188,N_4955,N_4922);
nor UO_189 (O_189,N_4946,N_4990);
xnor UO_190 (O_190,N_4936,N_4971);
or UO_191 (O_191,N_4975,N_4945);
or UO_192 (O_192,N_4955,N_4961);
nor UO_193 (O_193,N_4935,N_4949);
xor UO_194 (O_194,N_4992,N_4970);
nand UO_195 (O_195,N_4992,N_4995);
nor UO_196 (O_196,N_4961,N_4903);
or UO_197 (O_197,N_4901,N_4988);
nand UO_198 (O_198,N_4938,N_4996);
xor UO_199 (O_199,N_4958,N_4912);
or UO_200 (O_200,N_4919,N_4954);
or UO_201 (O_201,N_4975,N_4916);
or UO_202 (O_202,N_4950,N_4938);
nand UO_203 (O_203,N_4920,N_4980);
nor UO_204 (O_204,N_4990,N_4921);
nand UO_205 (O_205,N_4981,N_4905);
and UO_206 (O_206,N_4985,N_4975);
nor UO_207 (O_207,N_4950,N_4903);
xnor UO_208 (O_208,N_4977,N_4978);
nand UO_209 (O_209,N_4990,N_4999);
and UO_210 (O_210,N_4965,N_4970);
nor UO_211 (O_211,N_4995,N_4932);
nor UO_212 (O_212,N_4929,N_4911);
nor UO_213 (O_213,N_4926,N_4971);
or UO_214 (O_214,N_4945,N_4983);
nand UO_215 (O_215,N_4925,N_4953);
nor UO_216 (O_216,N_4925,N_4937);
nand UO_217 (O_217,N_4917,N_4916);
or UO_218 (O_218,N_4987,N_4934);
xnor UO_219 (O_219,N_4989,N_4903);
nand UO_220 (O_220,N_4925,N_4919);
or UO_221 (O_221,N_4919,N_4924);
or UO_222 (O_222,N_4913,N_4946);
nor UO_223 (O_223,N_4915,N_4950);
nor UO_224 (O_224,N_4913,N_4972);
nand UO_225 (O_225,N_4934,N_4925);
nor UO_226 (O_226,N_4992,N_4976);
nand UO_227 (O_227,N_4949,N_4968);
nor UO_228 (O_228,N_4917,N_4909);
nor UO_229 (O_229,N_4924,N_4954);
nor UO_230 (O_230,N_4983,N_4940);
nand UO_231 (O_231,N_4993,N_4995);
and UO_232 (O_232,N_4940,N_4965);
nor UO_233 (O_233,N_4957,N_4939);
and UO_234 (O_234,N_4918,N_4954);
nand UO_235 (O_235,N_4953,N_4935);
nand UO_236 (O_236,N_4900,N_4906);
or UO_237 (O_237,N_4949,N_4942);
or UO_238 (O_238,N_4954,N_4921);
nand UO_239 (O_239,N_4934,N_4907);
nand UO_240 (O_240,N_4938,N_4904);
nor UO_241 (O_241,N_4909,N_4985);
nor UO_242 (O_242,N_4967,N_4910);
nand UO_243 (O_243,N_4985,N_4955);
xnor UO_244 (O_244,N_4903,N_4971);
and UO_245 (O_245,N_4948,N_4992);
nor UO_246 (O_246,N_4912,N_4924);
nand UO_247 (O_247,N_4936,N_4993);
nor UO_248 (O_248,N_4953,N_4962);
nand UO_249 (O_249,N_4992,N_4965);
nand UO_250 (O_250,N_4932,N_4996);
nor UO_251 (O_251,N_4905,N_4934);
and UO_252 (O_252,N_4941,N_4984);
xnor UO_253 (O_253,N_4929,N_4994);
xor UO_254 (O_254,N_4924,N_4939);
nand UO_255 (O_255,N_4945,N_4931);
and UO_256 (O_256,N_4935,N_4950);
and UO_257 (O_257,N_4964,N_4983);
nor UO_258 (O_258,N_4990,N_4980);
or UO_259 (O_259,N_4905,N_4916);
or UO_260 (O_260,N_4932,N_4912);
xnor UO_261 (O_261,N_4961,N_4974);
and UO_262 (O_262,N_4966,N_4909);
xnor UO_263 (O_263,N_4973,N_4929);
nand UO_264 (O_264,N_4919,N_4903);
and UO_265 (O_265,N_4969,N_4964);
xnor UO_266 (O_266,N_4954,N_4965);
nand UO_267 (O_267,N_4911,N_4918);
xor UO_268 (O_268,N_4976,N_4921);
and UO_269 (O_269,N_4946,N_4929);
or UO_270 (O_270,N_4923,N_4910);
and UO_271 (O_271,N_4977,N_4969);
or UO_272 (O_272,N_4981,N_4901);
nor UO_273 (O_273,N_4939,N_4998);
or UO_274 (O_274,N_4938,N_4953);
xor UO_275 (O_275,N_4909,N_4951);
nand UO_276 (O_276,N_4953,N_4989);
or UO_277 (O_277,N_4965,N_4977);
and UO_278 (O_278,N_4933,N_4955);
or UO_279 (O_279,N_4958,N_4919);
or UO_280 (O_280,N_4977,N_4958);
or UO_281 (O_281,N_4956,N_4910);
nor UO_282 (O_282,N_4912,N_4938);
or UO_283 (O_283,N_4992,N_4987);
nor UO_284 (O_284,N_4964,N_4931);
or UO_285 (O_285,N_4956,N_4970);
nor UO_286 (O_286,N_4937,N_4957);
and UO_287 (O_287,N_4969,N_4978);
nor UO_288 (O_288,N_4951,N_4952);
nor UO_289 (O_289,N_4990,N_4944);
nor UO_290 (O_290,N_4937,N_4922);
nand UO_291 (O_291,N_4925,N_4946);
nand UO_292 (O_292,N_4993,N_4924);
and UO_293 (O_293,N_4989,N_4961);
or UO_294 (O_294,N_4983,N_4943);
xnor UO_295 (O_295,N_4969,N_4959);
and UO_296 (O_296,N_4936,N_4967);
nor UO_297 (O_297,N_4902,N_4915);
or UO_298 (O_298,N_4948,N_4981);
and UO_299 (O_299,N_4956,N_4952);
nor UO_300 (O_300,N_4923,N_4907);
and UO_301 (O_301,N_4906,N_4968);
nand UO_302 (O_302,N_4929,N_4949);
nand UO_303 (O_303,N_4970,N_4917);
nand UO_304 (O_304,N_4962,N_4919);
and UO_305 (O_305,N_4947,N_4929);
nand UO_306 (O_306,N_4905,N_4900);
or UO_307 (O_307,N_4932,N_4961);
xnor UO_308 (O_308,N_4974,N_4940);
and UO_309 (O_309,N_4944,N_4932);
nor UO_310 (O_310,N_4955,N_4963);
or UO_311 (O_311,N_4939,N_4911);
nand UO_312 (O_312,N_4911,N_4931);
nand UO_313 (O_313,N_4969,N_4957);
nand UO_314 (O_314,N_4923,N_4993);
and UO_315 (O_315,N_4975,N_4977);
or UO_316 (O_316,N_4969,N_4911);
and UO_317 (O_317,N_4977,N_4921);
nor UO_318 (O_318,N_4980,N_4928);
nand UO_319 (O_319,N_4997,N_4932);
and UO_320 (O_320,N_4945,N_4995);
xor UO_321 (O_321,N_4908,N_4944);
xor UO_322 (O_322,N_4978,N_4931);
nand UO_323 (O_323,N_4943,N_4942);
or UO_324 (O_324,N_4937,N_4987);
or UO_325 (O_325,N_4938,N_4969);
nand UO_326 (O_326,N_4924,N_4934);
xnor UO_327 (O_327,N_4910,N_4998);
xor UO_328 (O_328,N_4959,N_4904);
or UO_329 (O_329,N_4936,N_4998);
and UO_330 (O_330,N_4945,N_4934);
nor UO_331 (O_331,N_4964,N_4976);
nor UO_332 (O_332,N_4984,N_4943);
and UO_333 (O_333,N_4954,N_4901);
or UO_334 (O_334,N_4999,N_4966);
and UO_335 (O_335,N_4988,N_4934);
or UO_336 (O_336,N_4977,N_4912);
and UO_337 (O_337,N_4957,N_4912);
nand UO_338 (O_338,N_4946,N_4908);
and UO_339 (O_339,N_4961,N_4975);
or UO_340 (O_340,N_4951,N_4997);
nor UO_341 (O_341,N_4955,N_4940);
nand UO_342 (O_342,N_4922,N_4933);
and UO_343 (O_343,N_4998,N_4991);
nor UO_344 (O_344,N_4908,N_4915);
nand UO_345 (O_345,N_4960,N_4922);
or UO_346 (O_346,N_4956,N_4995);
nand UO_347 (O_347,N_4956,N_4957);
nor UO_348 (O_348,N_4991,N_4941);
nand UO_349 (O_349,N_4964,N_4972);
and UO_350 (O_350,N_4953,N_4988);
or UO_351 (O_351,N_4972,N_4902);
nand UO_352 (O_352,N_4940,N_4900);
and UO_353 (O_353,N_4917,N_4925);
nor UO_354 (O_354,N_4919,N_4946);
and UO_355 (O_355,N_4958,N_4934);
nor UO_356 (O_356,N_4904,N_4909);
nor UO_357 (O_357,N_4915,N_4992);
or UO_358 (O_358,N_4979,N_4924);
or UO_359 (O_359,N_4964,N_4933);
nand UO_360 (O_360,N_4957,N_4986);
and UO_361 (O_361,N_4999,N_4936);
and UO_362 (O_362,N_4902,N_4961);
or UO_363 (O_363,N_4949,N_4981);
xor UO_364 (O_364,N_4995,N_4911);
nor UO_365 (O_365,N_4933,N_4935);
nand UO_366 (O_366,N_4914,N_4927);
or UO_367 (O_367,N_4966,N_4946);
nand UO_368 (O_368,N_4902,N_4975);
and UO_369 (O_369,N_4925,N_4924);
or UO_370 (O_370,N_4977,N_4948);
nand UO_371 (O_371,N_4944,N_4929);
nor UO_372 (O_372,N_4983,N_4938);
xor UO_373 (O_373,N_4965,N_4979);
or UO_374 (O_374,N_4959,N_4924);
nand UO_375 (O_375,N_4937,N_4974);
and UO_376 (O_376,N_4927,N_4938);
nand UO_377 (O_377,N_4971,N_4932);
or UO_378 (O_378,N_4911,N_4977);
xor UO_379 (O_379,N_4937,N_4971);
nor UO_380 (O_380,N_4908,N_4934);
nor UO_381 (O_381,N_4921,N_4930);
nand UO_382 (O_382,N_4983,N_4981);
xnor UO_383 (O_383,N_4915,N_4982);
and UO_384 (O_384,N_4916,N_4902);
or UO_385 (O_385,N_4902,N_4985);
nand UO_386 (O_386,N_4949,N_4999);
nand UO_387 (O_387,N_4946,N_4949);
xnor UO_388 (O_388,N_4910,N_4943);
xnor UO_389 (O_389,N_4920,N_4974);
and UO_390 (O_390,N_4905,N_4973);
or UO_391 (O_391,N_4944,N_4975);
nor UO_392 (O_392,N_4915,N_4980);
or UO_393 (O_393,N_4932,N_4954);
nor UO_394 (O_394,N_4919,N_4921);
nor UO_395 (O_395,N_4983,N_4908);
and UO_396 (O_396,N_4986,N_4977);
and UO_397 (O_397,N_4929,N_4908);
nor UO_398 (O_398,N_4975,N_4954);
and UO_399 (O_399,N_4919,N_4936);
nand UO_400 (O_400,N_4916,N_4932);
and UO_401 (O_401,N_4928,N_4993);
nor UO_402 (O_402,N_4997,N_4967);
and UO_403 (O_403,N_4967,N_4904);
and UO_404 (O_404,N_4976,N_4914);
or UO_405 (O_405,N_4941,N_4973);
or UO_406 (O_406,N_4946,N_4904);
nor UO_407 (O_407,N_4993,N_4996);
nand UO_408 (O_408,N_4978,N_4957);
and UO_409 (O_409,N_4951,N_4979);
nor UO_410 (O_410,N_4962,N_4922);
nand UO_411 (O_411,N_4916,N_4906);
nor UO_412 (O_412,N_4973,N_4978);
or UO_413 (O_413,N_4956,N_4961);
nand UO_414 (O_414,N_4906,N_4973);
or UO_415 (O_415,N_4972,N_4965);
nor UO_416 (O_416,N_4927,N_4922);
nand UO_417 (O_417,N_4963,N_4938);
or UO_418 (O_418,N_4932,N_4960);
nand UO_419 (O_419,N_4934,N_4939);
nor UO_420 (O_420,N_4998,N_4931);
and UO_421 (O_421,N_4969,N_4922);
nand UO_422 (O_422,N_4915,N_4964);
and UO_423 (O_423,N_4958,N_4978);
xnor UO_424 (O_424,N_4951,N_4950);
and UO_425 (O_425,N_4952,N_4976);
and UO_426 (O_426,N_4908,N_4998);
xnor UO_427 (O_427,N_4945,N_4942);
and UO_428 (O_428,N_4959,N_4991);
xnor UO_429 (O_429,N_4922,N_4978);
nand UO_430 (O_430,N_4938,N_4943);
nor UO_431 (O_431,N_4931,N_4923);
and UO_432 (O_432,N_4909,N_4910);
or UO_433 (O_433,N_4933,N_4963);
or UO_434 (O_434,N_4954,N_4937);
nor UO_435 (O_435,N_4954,N_4920);
nor UO_436 (O_436,N_4957,N_4934);
nand UO_437 (O_437,N_4960,N_4914);
nand UO_438 (O_438,N_4967,N_4969);
xor UO_439 (O_439,N_4968,N_4957);
nor UO_440 (O_440,N_4902,N_4938);
and UO_441 (O_441,N_4980,N_4953);
xor UO_442 (O_442,N_4982,N_4905);
nor UO_443 (O_443,N_4922,N_4949);
nor UO_444 (O_444,N_4925,N_4943);
nor UO_445 (O_445,N_4933,N_4974);
or UO_446 (O_446,N_4958,N_4928);
nor UO_447 (O_447,N_4947,N_4925);
nor UO_448 (O_448,N_4987,N_4949);
nor UO_449 (O_449,N_4956,N_4982);
nor UO_450 (O_450,N_4956,N_4918);
xor UO_451 (O_451,N_4998,N_4944);
and UO_452 (O_452,N_4909,N_4946);
nand UO_453 (O_453,N_4905,N_4953);
nor UO_454 (O_454,N_4962,N_4975);
nor UO_455 (O_455,N_4948,N_4903);
nor UO_456 (O_456,N_4958,N_4982);
or UO_457 (O_457,N_4912,N_4936);
nor UO_458 (O_458,N_4907,N_4936);
nor UO_459 (O_459,N_4924,N_4986);
nor UO_460 (O_460,N_4976,N_4923);
xnor UO_461 (O_461,N_4935,N_4915);
xnor UO_462 (O_462,N_4951,N_4977);
nor UO_463 (O_463,N_4961,N_4976);
nand UO_464 (O_464,N_4914,N_4983);
nand UO_465 (O_465,N_4972,N_4984);
or UO_466 (O_466,N_4966,N_4945);
nand UO_467 (O_467,N_4919,N_4934);
and UO_468 (O_468,N_4993,N_4952);
nor UO_469 (O_469,N_4901,N_4934);
and UO_470 (O_470,N_4911,N_4915);
or UO_471 (O_471,N_4965,N_4948);
nand UO_472 (O_472,N_4984,N_4938);
xnor UO_473 (O_473,N_4911,N_4971);
and UO_474 (O_474,N_4936,N_4991);
nor UO_475 (O_475,N_4928,N_4951);
and UO_476 (O_476,N_4955,N_4907);
and UO_477 (O_477,N_4946,N_4958);
nor UO_478 (O_478,N_4954,N_4973);
or UO_479 (O_479,N_4989,N_4931);
nor UO_480 (O_480,N_4991,N_4926);
nand UO_481 (O_481,N_4936,N_4968);
nor UO_482 (O_482,N_4990,N_4922);
nand UO_483 (O_483,N_4976,N_4926);
xnor UO_484 (O_484,N_4973,N_4961);
and UO_485 (O_485,N_4918,N_4965);
xor UO_486 (O_486,N_4951,N_4972);
nand UO_487 (O_487,N_4950,N_4999);
nor UO_488 (O_488,N_4994,N_4902);
nor UO_489 (O_489,N_4977,N_4925);
nor UO_490 (O_490,N_4960,N_4994);
nor UO_491 (O_491,N_4923,N_4959);
nor UO_492 (O_492,N_4906,N_4991);
and UO_493 (O_493,N_4994,N_4996);
nor UO_494 (O_494,N_4998,N_4993);
and UO_495 (O_495,N_4949,N_4992);
or UO_496 (O_496,N_4951,N_4942);
or UO_497 (O_497,N_4966,N_4929);
and UO_498 (O_498,N_4999,N_4930);
and UO_499 (O_499,N_4918,N_4909);
or UO_500 (O_500,N_4978,N_4962);
nand UO_501 (O_501,N_4986,N_4909);
xnor UO_502 (O_502,N_4960,N_4981);
nor UO_503 (O_503,N_4923,N_4991);
nand UO_504 (O_504,N_4924,N_4983);
xnor UO_505 (O_505,N_4908,N_4909);
and UO_506 (O_506,N_4955,N_4929);
and UO_507 (O_507,N_4956,N_4942);
and UO_508 (O_508,N_4956,N_4950);
nand UO_509 (O_509,N_4958,N_4988);
or UO_510 (O_510,N_4937,N_4967);
nor UO_511 (O_511,N_4946,N_4905);
or UO_512 (O_512,N_4943,N_4913);
or UO_513 (O_513,N_4995,N_4905);
nand UO_514 (O_514,N_4935,N_4990);
nand UO_515 (O_515,N_4950,N_4926);
nor UO_516 (O_516,N_4984,N_4903);
nor UO_517 (O_517,N_4938,N_4964);
or UO_518 (O_518,N_4997,N_4931);
or UO_519 (O_519,N_4906,N_4974);
nand UO_520 (O_520,N_4990,N_4915);
nor UO_521 (O_521,N_4986,N_4916);
nand UO_522 (O_522,N_4911,N_4975);
nor UO_523 (O_523,N_4904,N_4994);
nand UO_524 (O_524,N_4924,N_4929);
xnor UO_525 (O_525,N_4907,N_4972);
and UO_526 (O_526,N_4910,N_4989);
nand UO_527 (O_527,N_4925,N_4966);
nor UO_528 (O_528,N_4968,N_4941);
or UO_529 (O_529,N_4992,N_4901);
and UO_530 (O_530,N_4973,N_4924);
and UO_531 (O_531,N_4971,N_4914);
or UO_532 (O_532,N_4903,N_4999);
and UO_533 (O_533,N_4916,N_4984);
or UO_534 (O_534,N_4968,N_4960);
xor UO_535 (O_535,N_4973,N_4957);
and UO_536 (O_536,N_4972,N_4956);
nand UO_537 (O_537,N_4910,N_4996);
nand UO_538 (O_538,N_4960,N_4935);
and UO_539 (O_539,N_4918,N_4986);
or UO_540 (O_540,N_4904,N_4960);
or UO_541 (O_541,N_4914,N_4921);
xor UO_542 (O_542,N_4983,N_4906);
nor UO_543 (O_543,N_4984,N_4918);
or UO_544 (O_544,N_4943,N_4971);
xor UO_545 (O_545,N_4926,N_4957);
nor UO_546 (O_546,N_4911,N_4991);
or UO_547 (O_547,N_4915,N_4952);
or UO_548 (O_548,N_4994,N_4932);
or UO_549 (O_549,N_4995,N_4914);
or UO_550 (O_550,N_4997,N_4973);
nand UO_551 (O_551,N_4956,N_4958);
nand UO_552 (O_552,N_4914,N_4905);
and UO_553 (O_553,N_4944,N_4930);
and UO_554 (O_554,N_4915,N_4930);
and UO_555 (O_555,N_4930,N_4980);
xnor UO_556 (O_556,N_4900,N_4957);
or UO_557 (O_557,N_4925,N_4962);
nand UO_558 (O_558,N_4941,N_4994);
nor UO_559 (O_559,N_4914,N_4974);
or UO_560 (O_560,N_4922,N_4946);
nor UO_561 (O_561,N_4999,N_4963);
nor UO_562 (O_562,N_4946,N_4996);
nand UO_563 (O_563,N_4969,N_4992);
or UO_564 (O_564,N_4991,N_4979);
nand UO_565 (O_565,N_4935,N_4936);
and UO_566 (O_566,N_4966,N_4954);
or UO_567 (O_567,N_4950,N_4933);
and UO_568 (O_568,N_4944,N_4951);
or UO_569 (O_569,N_4973,N_4928);
and UO_570 (O_570,N_4906,N_4929);
or UO_571 (O_571,N_4949,N_4961);
xor UO_572 (O_572,N_4939,N_4956);
nor UO_573 (O_573,N_4918,N_4906);
and UO_574 (O_574,N_4902,N_4904);
or UO_575 (O_575,N_4951,N_4934);
nor UO_576 (O_576,N_4916,N_4950);
nor UO_577 (O_577,N_4967,N_4979);
and UO_578 (O_578,N_4993,N_4988);
xnor UO_579 (O_579,N_4942,N_4938);
and UO_580 (O_580,N_4981,N_4920);
nor UO_581 (O_581,N_4971,N_4942);
or UO_582 (O_582,N_4963,N_4936);
nor UO_583 (O_583,N_4904,N_4943);
nor UO_584 (O_584,N_4987,N_4984);
nor UO_585 (O_585,N_4931,N_4977);
nand UO_586 (O_586,N_4963,N_4917);
nor UO_587 (O_587,N_4987,N_4972);
and UO_588 (O_588,N_4998,N_4904);
nand UO_589 (O_589,N_4989,N_4947);
nor UO_590 (O_590,N_4969,N_4912);
xnor UO_591 (O_591,N_4916,N_4941);
nand UO_592 (O_592,N_4986,N_4946);
nand UO_593 (O_593,N_4958,N_4992);
and UO_594 (O_594,N_4981,N_4936);
nand UO_595 (O_595,N_4985,N_4910);
and UO_596 (O_596,N_4908,N_4902);
nand UO_597 (O_597,N_4938,N_4934);
and UO_598 (O_598,N_4948,N_4942);
nor UO_599 (O_599,N_4957,N_4941);
nand UO_600 (O_600,N_4903,N_4966);
nor UO_601 (O_601,N_4958,N_4975);
and UO_602 (O_602,N_4995,N_4958);
nor UO_603 (O_603,N_4901,N_4977);
or UO_604 (O_604,N_4986,N_4915);
nand UO_605 (O_605,N_4982,N_4960);
nand UO_606 (O_606,N_4940,N_4985);
or UO_607 (O_607,N_4984,N_4990);
xor UO_608 (O_608,N_4932,N_4967);
and UO_609 (O_609,N_4935,N_4965);
xnor UO_610 (O_610,N_4970,N_4984);
xnor UO_611 (O_611,N_4964,N_4998);
or UO_612 (O_612,N_4956,N_4947);
and UO_613 (O_613,N_4913,N_4968);
nor UO_614 (O_614,N_4985,N_4926);
xnor UO_615 (O_615,N_4959,N_4948);
or UO_616 (O_616,N_4906,N_4905);
or UO_617 (O_617,N_4996,N_4960);
or UO_618 (O_618,N_4902,N_4906);
xor UO_619 (O_619,N_4978,N_4949);
nand UO_620 (O_620,N_4925,N_4984);
nand UO_621 (O_621,N_4969,N_4970);
and UO_622 (O_622,N_4939,N_4935);
nor UO_623 (O_623,N_4997,N_4985);
nand UO_624 (O_624,N_4961,N_4967);
or UO_625 (O_625,N_4992,N_4931);
and UO_626 (O_626,N_4996,N_4908);
or UO_627 (O_627,N_4960,N_4957);
or UO_628 (O_628,N_4908,N_4970);
nand UO_629 (O_629,N_4959,N_4921);
or UO_630 (O_630,N_4937,N_4985);
nor UO_631 (O_631,N_4934,N_4963);
and UO_632 (O_632,N_4968,N_4924);
xor UO_633 (O_633,N_4906,N_4965);
nand UO_634 (O_634,N_4979,N_4942);
nand UO_635 (O_635,N_4919,N_4923);
nor UO_636 (O_636,N_4958,N_4971);
or UO_637 (O_637,N_4975,N_4990);
nor UO_638 (O_638,N_4981,N_4975);
and UO_639 (O_639,N_4945,N_4918);
and UO_640 (O_640,N_4942,N_4961);
nand UO_641 (O_641,N_4942,N_4935);
or UO_642 (O_642,N_4920,N_4983);
and UO_643 (O_643,N_4982,N_4957);
xor UO_644 (O_644,N_4920,N_4944);
or UO_645 (O_645,N_4999,N_4924);
or UO_646 (O_646,N_4988,N_4902);
xnor UO_647 (O_647,N_4967,N_4968);
nor UO_648 (O_648,N_4918,N_4913);
nand UO_649 (O_649,N_4908,N_4950);
and UO_650 (O_650,N_4960,N_4944);
nor UO_651 (O_651,N_4946,N_4978);
or UO_652 (O_652,N_4906,N_4958);
or UO_653 (O_653,N_4952,N_4932);
and UO_654 (O_654,N_4949,N_4919);
and UO_655 (O_655,N_4949,N_4951);
nand UO_656 (O_656,N_4944,N_4970);
and UO_657 (O_657,N_4937,N_4963);
nand UO_658 (O_658,N_4905,N_4978);
or UO_659 (O_659,N_4957,N_4996);
nand UO_660 (O_660,N_4981,N_4913);
and UO_661 (O_661,N_4907,N_4995);
nor UO_662 (O_662,N_4953,N_4901);
xor UO_663 (O_663,N_4943,N_4912);
and UO_664 (O_664,N_4954,N_4988);
nor UO_665 (O_665,N_4918,N_4989);
or UO_666 (O_666,N_4995,N_4955);
nor UO_667 (O_667,N_4915,N_4979);
xnor UO_668 (O_668,N_4962,N_4990);
or UO_669 (O_669,N_4935,N_4952);
or UO_670 (O_670,N_4992,N_4946);
xor UO_671 (O_671,N_4993,N_4971);
xor UO_672 (O_672,N_4956,N_4980);
or UO_673 (O_673,N_4953,N_4946);
nand UO_674 (O_674,N_4904,N_4947);
or UO_675 (O_675,N_4917,N_4990);
or UO_676 (O_676,N_4973,N_4968);
nor UO_677 (O_677,N_4975,N_4993);
or UO_678 (O_678,N_4963,N_4932);
or UO_679 (O_679,N_4987,N_4941);
nor UO_680 (O_680,N_4988,N_4992);
or UO_681 (O_681,N_4959,N_4971);
or UO_682 (O_682,N_4966,N_4960);
nand UO_683 (O_683,N_4998,N_4926);
nand UO_684 (O_684,N_4977,N_4913);
nand UO_685 (O_685,N_4935,N_4927);
nor UO_686 (O_686,N_4961,N_4916);
nor UO_687 (O_687,N_4927,N_4995);
or UO_688 (O_688,N_4913,N_4973);
nor UO_689 (O_689,N_4951,N_4948);
nor UO_690 (O_690,N_4954,N_4915);
and UO_691 (O_691,N_4995,N_4998);
nand UO_692 (O_692,N_4949,N_4976);
and UO_693 (O_693,N_4952,N_4978);
or UO_694 (O_694,N_4970,N_4933);
xor UO_695 (O_695,N_4951,N_4905);
nor UO_696 (O_696,N_4955,N_4954);
and UO_697 (O_697,N_4984,N_4977);
and UO_698 (O_698,N_4965,N_4942);
or UO_699 (O_699,N_4977,N_4940);
and UO_700 (O_700,N_4906,N_4954);
nand UO_701 (O_701,N_4927,N_4969);
nand UO_702 (O_702,N_4969,N_4942);
and UO_703 (O_703,N_4944,N_4986);
or UO_704 (O_704,N_4910,N_4980);
or UO_705 (O_705,N_4945,N_4941);
xor UO_706 (O_706,N_4922,N_4957);
nor UO_707 (O_707,N_4910,N_4911);
nand UO_708 (O_708,N_4978,N_4915);
and UO_709 (O_709,N_4956,N_4902);
and UO_710 (O_710,N_4916,N_4949);
and UO_711 (O_711,N_4979,N_4970);
nor UO_712 (O_712,N_4900,N_4970);
nand UO_713 (O_713,N_4958,N_4923);
nand UO_714 (O_714,N_4911,N_4950);
or UO_715 (O_715,N_4991,N_4996);
xor UO_716 (O_716,N_4933,N_4944);
or UO_717 (O_717,N_4991,N_4924);
or UO_718 (O_718,N_4953,N_4984);
or UO_719 (O_719,N_4974,N_4938);
nor UO_720 (O_720,N_4933,N_4939);
or UO_721 (O_721,N_4929,N_4913);
nor UO_722 (O_722,N_4942,N_4939);
nand UO_723 (O_723,N_4926,N_4979);
nand UO_724 (O_724,N_4962,N_4948);
and UO_725 (O_725,N_4977,N_4939);
or UO_726 (O_726,N_4956,N_4940);
and UO_727 (O_727,N_4939,N_4961);
or UO_728 (O_728,N_4961,N_4960);
and UO_729 (O_729,N_4914,N_4989);
nand UO_730 (O_730,N_4907,N_4985);
or UO_731 (O_731,N_4988,N_4907);
and UO_732 (O_732,N_4908,N_4937);
and UO_733 (O_733,N_4929,N_4901);
or UO_734 (O_734,N_4907,N_4904);
nor UO_735 (O_735,N_4945,N_4948);
nor UO_736 (O_736,N_4908,N_4952);
nand UO_737 (O_737,N_4923,N_4966);
nor UO_738 (O_738,N_4908,N_4969);
xor UO_739 (O_739,N_4951,N_4927);
nand UO_740 (O_740,N_4997,N_4950);
and UO_741 (O_741,N_4935,N_4984);
and UO_742 (O_742,N_4977,N_4900);
and UO_743 (O_743,N_4993,N_4947);
xor UO_744 (O_744,N_4972,N_4954);
and UO_745 (O_745,N_4943,N_4969);
and UO_746 (O_746,N_4952,N_4986);
xor UO_747 (O_747,N_4902,N_4978);
or UO_748 (O_748,N_4977,N_4950);
and UO_749 (O_749,N_4924,N_4997);
or UO_750 (O_750,N_4952,N_4972);
nor UO_751 (O_751,N_4928,N_4929);
nand UO_752 (O_752,N_4981,N_4923);
nand UO_753 (O_753,N_4986,N_4913);
or UO_754 (O_754,N_4946,N_4974);
and UO_755 (O_755,N_4996,N_4905);
nor UO_756 (O_756,N_4937,N_4965);
nand UO_757 (O_757,N_4905,N_4904);
and UO_758 (O_758,N_4978,N_4907);
or UO_759 (O_759,N_4978,N_4966);
nor UO_760 (O_760,N_4980,N_4947);
nor UO_761 (O_761,N_4927,N_4911);
or UO_762 (O_762,N_4918,N_4935);
xnor UO_763 (O_763,N_4914,N_4982);
nor UO_764 (O_764,N_4920,N_4925);
or UO_765 (O_765,N_4982,N_4920);
or UO_766 (O_766,N_4982,N_4944);
or UO_767 (O_767,N_4917,N_4966);
or UO_768 (O_768,N_4939,N_4908);
or UO_769 (O_769,N_4973,N_4995);
nor UO_770 (O_770,N_4984,N_4960);
nand UO_771 (O_771,N_4935,N_4947);
nand UO_772 (O_772,N_4998,N_4986);
xnor UO_773 (O_773,N_4947,N_4996);
nand UO_774 (O_774,N_4907,N_4910);
or UO_775 (O_775,N_4901,N_4917);
nand UO_776 (O_776,N_4912,N_4935);
nand UO_777 (O_777,N_4934,N_4910);
nand UO_778 (O_778,N_4939,N_4904);
and UO_779 (O_779,N_4906,N_4901);
and UO_780 (O_780,N_4981,N_4927);
or UO_781 (O_781,N_4975,N_4918);
and UO_782 (O_782,N_4978,N_4916);
nor UO_783 (O_783,N_4984,N_4956);
nor UO_784 (O_784,N_4980,N_4998);
nor UO_785 (O_785,N_4905,N_4991);
nand UO_786 (O_786,N_4944,N_4947);
or UO_787 (O_787,N_4989,N_4991);
nand UO_788 (O_788,N_4911,N_4957);
xor UO_789 (O_789,N_4978,N_4933);
and UO_790 (O_790,N_4971,N_4913);
and UO_791 (O_791,N_4994,N_4911);
xnor UO_792 (O_792,N_4960,N_4943);
nand UO_793 (O_793,N_4994,N_4927);
nand UO_794 (O_794,N_4963,N_4910);
nand UO_795 (O_795,N_4955,N_4997);
or UO_796 (O_796,N_4960,N_4930);
nor UO_797 (O_797,N_4970,N_4946);
nor UO_798 (O_798,N_4976,N_4939);
nand UO_799 (O_799,N_4923,N_4936);
nand UO_800 (O_800,N_4985,N_4978);
xnor UO_801 (O_801,N_4900,N_4979);
or UO_802 (O_802,N_4935,N_4905);
nor UO_803 (O_803,N_4955,N_4959);
nand UO_804 (O_804,N_4949,N_4982);
nand UO_805 (O_805,N_4952,N_4966);
and UO_806 (O_806,N_4949,N_4997);
or UO_807 (O_807,N_4938,N_4911);
or UO_808 (O_808,N_4904,N_4979);
nand UO_809 (O_809,N_4947,N_4969);
nand UO_810 (O_810,N_4902,N_4935);
nand UO_811 (O_811,N_4997,N_4943);
nand UO_812 (O_812,N_4920,N_4965);
or UO_813 (O_813,N_4975,N_4939);
and UO_814 (O_814,N_4971,N_4970);
or UO_815 (O_815,N_4955,N_4932);
or UO_816 (O_816,N_4900,N_4949);
nor UO_817 (O_817,N_4964,N_4949);
or UO_818 (O_818,N_4911,N_4956);
nor UO_819 (O_819,N_4987,N_4938);
and UO_820 (O_820,N_4933,N_4924);
or UO_821 (O_821,N_4944,N_4966);
nand UO_822 (O_822,N_4929,N_4912);
and UO_823 (O_823,N_4942,N_4977);
or UO_824 (O_824,N_4990,N_4988);
nand UO_825 (O_825,N_4900,N_4910);
and UO_826 (O_826,N_4949,N_4945);
or UO_827 (O_827,N_4906,N_4922);
nor UO_828 (O_828,N_4978,N_4901);
nor UO_829 (O_829,N_4970,N_4927);
and UO_830 (O_830,N_4958,N_4943);
nor UO_831 (O_831,N_4997,N_4902);
nand UO_832 (O_832,N_4978,N_4990);
nand UO_833 (O_833,N_4977,N_4990);
and UO_834 (O_834,N_4932,N_4948);
xor UO_835 (O_835,N_4920,N_4919);
nand UO_836 (O_836,N_4956,N_4999);
or UO_837 (O_837,N_4958,N_4983);
nor UO_838 (O_838,N_4940,N_4996);
or UO_839 (O_839,N_4938,N_4990);
nand UO_840 (O_840,N_4957,N_4943);
nor UO_841 (O_841,N_4936,N_4988);
nand UO_842 (O_842,N_4996,N_4935);
nor UO_843 (O_843,N_4967,N_4972);
nor UO_844 (O_844,N_4989,N_4913);
and UO_845 (O_845,N_4943,N_4991);
nor UO_846 (O_846,N_4915,N_4941);
nand UO_847 (O_847,N_4929,N_4988);
nand UO_848 (O_848,N_4945,N_4963);
nor UO_849 (O_849,N_4910,N_4901);
nand UO_850 (O_850,N_4959,N_4999);
or UO_851 (O_851,N_4958,N_4915);
or UO_852 (O_852,N_4910,N_4953);
and UO_853 (O_853,N_4926,N_4954);
and UO_854 (O_854,N_4988,N_4981);
or UO_855 (O_855,N_4911,N_4951);
or UO_856 (O_856,N_4966,N_4918);
or UO_857 (O_857,N_4904,N_4965);
nand UO_858 (O_858,N_4976,N_4986);
nand UO_859 (O_859,N_4956,N_4955);
nor UO_860 (O_860,N_4962,N_4983);
and UO_861 (O_861,N_4956,N_4991);
or UO_862 (O_862,N_4993,N_4932);
nand UO_863 (O_863,N_4924,N_4905);
nor UO_864 (O_864,N_4984,N_4913);
nand UO_865 (O_865,N_4907,N_4900);
or UO_866 (O_866,N_4999,N_4991);
and UO_867 (O_867,N_4950,N_4936);
nand UO_868 (O_868,N_4943,N_4924);
nor UO_869 (O_869,N_4973,N_4980);
nand UO_870 (O_870,N_4938,N_4944);
nand UO_871 (O_871,N_4922,N_4983);
nand UO_872 (O_872,N_4990,N_4954);
or UO_873 (O_873,N_4917,N_4951);
nor UO_874 (O_874,N_4970,N_4975);
xor UO_875 (O_875,N_4921,N_4911);
nor UO_876 (O_876,N_4984,N_4929);
and UO_877 (O_877,N_4998,N_4933);
nor UO_878 (O_878,N_4972,N_4933);
nand UO_879 (O_879,N_4967,N_4934);
nor UO_880 (O_880,N_4957,N_4974);
nor UO_881 (O_881,N_4937,N_4966);
nor UO_882 (O_882,N_4966,N_4988);
and UO_883 (O_883,N_4926,N_4989);
nor UO_884 (O_884,N_4972,N_4940);
nand UO_885 (O_885,N_4976,N_4970);
nor UO_886 (O_886,N_4981,N_4964);
nor UO_887 (O_887,N_4917,N_4935);
and UO_888 (O_888,N_4985,N_4951);
nor UO_889 (O_889,N_4930,N_4965);
or UO_890 (O_890,N_4923,N_4927);
xor UO_891 (O_891,N_4981,N_4944);
or UO_892 (O_892,N_4963,N_4927);
and UO_893 (O_893,N_4976,N_4959);
nand UO_894 (O_894,N_4949,N_4914);
nand UO_895 (O_895,N_4929,N_4962);
nor UO_896 (O_896,N_4967,N_4987);
or UO_897 (O_897,N_4966,N_4932);
nand UO_898 (O_898,N_4908,N_4987);
or UO_899 (O_899,N_4979,N_4969);
nand UO_900 (O_900,N_4907,N_4926);
and UO_901 (O_901,N_4981,N_4916);
nand UO_902 (O_902,N_4904,N_4976);
xor UO_903 (O_903,N_4925,N_4955);
xnor UO_904 (O_904,N_4985,N_4994);
xnor UO_905 (O_905,N_4951,N_4967);
nor UO_906 (O_906,N_4941,N_4921);
and UO_907 (O_907,N_4997,N_4926);
and UO_908 (O_908,N_4948,N_4908);
nor UO_909 (O_909,N_4920,N_4914);
or UO_910 (O_910,N_4960,N_4999);
nor UO_911 (O_911,N_4946,N_4994);
or UO_912 (O_912,N_4999,N_4910);
nor UO_913 (O_913,N_4963,N_4918);
nand UO_914 (O_914,N_4985,N_4949);
nor UO_915 (O_915,N_4968,N_4971);
or UO_916 (O_916,N_4946,N_4900);
or UO_917 (O_917,N_4917,N_4902);
or UO_918 (O_918,N_4976,N_4912);
or UO_919 (O_919,N_4958,N_4949);
nand UO_920 (O_920,N_4970,N_4909);
or UO_921 (O_921,N_4928,N_4917);
and UO_922 (O_922,N_4926,N_4912);
and UO_923 (O_923,N_4963,N_4930);
nand UO_924 (O_924,N_4934,N_4953);
xor UO_925 (O_925,N_4992,N_4952);
xnor UO_926 (O_926,N_4925,N_4972);
nor UO_927 (O_927,N_4920,N_4930);
nor UO_928 (O_928,N_4976,N_4965);
nand UO_929 (O_929,N_4959,N_4930);
xor UO_930 (O_930,N_4959,N_4915);
nor UO_931 (O_931,N_4979,N_4995);
nand UO_932 (O_932,N_4907,N_4917);
or UO_933 (O_933,N_4998,N_4953);
xnor UO_934 (O_934,N_4946,N_4998);
and UO_935 (O_935,N_4912,N_4971);
nand UO_936 (O_936,N_4916,N_4924);
or UO_937 (O_937,N_4935,N_4948);
nor UO_938 (O_938,N_4900,N_4928);
and UO_939 (O_939,N_4980,N_4974);
or UO_940 (O_940,N_4988,N_4974);
or UO_941 (O_941,N_4972,N_4930);
nand UO_942 (O_942,N_4983,N_4995);
nor UO_943 (O_943,N_4960,N_4970);
nor UO_944 (O_944,N_4965,N_4996);
nor UO_945 (O_945,N_4965,N_4944);
nand UO_946 (O_946,N_4905,N_4950);
and UO_947 (O_947,N_4920,N_4987);
nand UO_948 (O_948,N_4908,N_4986);
and UO_949 (O_949,N_4953,N_4939);
nand UO_950 (O_950,N_4954,N_4925);
nor UO_951 (O_951,N_4946,N_4915);
nor UO_952 (O_952,N_4919,N_4928);
and UO_953 (O_953,N_4920,N_4907);
nor UO_954 (O_954,N_4902,N_4992);
and UO_955 (O_955,N_4924,N_4918);
and UO_956 (O_956,N_4975,N_4960);
xor UO_957 (O_957,N_4963,N_4901);
or UO_958 (O_958,N_4906,N_4999);
nor UO_959 (O_959,N_4958,N_4961);
xor UO_960 (O_960,N_4951,N_4971);
and UO_961 (O_961,N_4947,N_4938);
nor UO_962 (O_962,N_4938,N_4907);
and UO_963 (O_963,N_4992,N_4945);
and UO_964 (O_964,N_4940,N_4951);
or UO_965 (O_965,N_4960,N_4919);
nor UO_966 (O_966,N_4933,N_4986);
nand UO_967 (O_967,N_4935,N_4971);
nand UO_968 (O_968,N_4992,N_4998);
nor UO_969 (O_969,N_4939,N_4936);
and UO_970 (O_970,N_4926,N_4914);
xnor UO_971 (O_971,N_4933,N_4936);
nand UO_972 (O_972,N_4981,N_4987);
xor UO_973 (O_973,N_4915,N_4940);
nand UO_974 (O_974,N_4914,N_4961);
and UO_975 (O_975,N_4999,N_4902);
xor UO_976 (O_976,N_4951,N_4975);
and UO_977 (O_977,N_4927,N_4906);
nor UO_978 (O_978,N_4949,N_4956);
or UO_979 (O_979,N_4988,N_4952);
nor UO_980 (O_980,N_4982,N_4964);
nor UO_981 (O_981,N_4977,N_4932);
nand UO_982 (O_982,N_4967,N_4944);
or UO_983 (O_983,N_4990,N_4918);
nor UO_984 (O_984,N_4946,N_4977);
nor UO_985 (O_985,N_4905,N_4992);
nand UO_986 (O_986,N_4942,N_4966);
nand UO_987 (O_987,N_4993,N_4972);
nand UO_988 (O_988,N_4921,N_4995);
xnor UO_989 (O_989,N_4958,N_4987);
nor UO_990 (O_990,N_4912,N_4939);
and UO_991 (O_991,N_4939,N_4983);
xor UO_992 (O_992,N_4968,N_4914);
nand UO_993 (O_993,N_4985,N_4935);
and UO_994 (O_994,N_4995,N_4936);
or UO_995 (O_995,N_4912,N_4921);
nand UO_996 (O_996,N_4980,N_4993);
nand UO_997 (O_997,N_4963,N_4943);
xnor UO_998 (O_998,N_4961,N_4971);
nand UO_999 (O_999,N_4952,N_4902);
endmodule