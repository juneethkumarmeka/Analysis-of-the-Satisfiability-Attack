module basic_1000_10000_1500_5_levels_1xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_804,In_393);
nor U1 (N_1,In_775,In_958);
nor U2 (N_2,In_491,In_989);
or U3 (N_3,In_311,In_808);
nor U4 (N_4,In_157,In_684);
nand U5 (N_5,In_801,In_730);
and U6 (N_6,In_881,In_639);
and U7 (N_7,In_670,In_585);
or U8 (N_8,In_446,In_758);
nor U9 (N_9,In_27,In_54);
or U10 (N_10,In_498,In_256);
nand U11 (N_11,In_332,In_742);
nand U12 (N_12,In_611,In_705);
and U13 (N_13,In_188,In_479);
or U14 (N_14,In_923,In_221);
nand U15 (N_15,In_316,In_325);
nor U16 (N_16,In_367,In_592);
nor U17 (N_17,In_568,In_744);
or U18 (N_18,In_652,In_64);
nand U19 (N_19,In_388,In_732);
nand U20 (N_20,In_233,In_244);
nor U21 (N_21,In_867,In_455);
nor U22 (N_22,In_628,In_603);
or U23 (N_23,In_712,In_999);
or U24 (N_24,In_165,In_594);
nand U25 (N_25,In_1,In_132);
nand U26 (N_26,In_547,In_212);
nor U27 (N_27,In_394,In_154);
nor U28 (N_28,In_841,In_770);
or U29 (N_29,In_751,In_747);
nor U30 (N_30,In_726,In_395);
nand U31 (N_31,In_102,In_475);
or U32 (N_32,In_86,In_908);
nand U33 (N_33,In_492,In_284);
nand U34 (N_34,In_624,In_831);
or U35 (N_35,In_225,In_308);
or U36 (N_36,In_363,In_882);
or U37 (N_37,In_607,In_650);
and U38 (N_38,In_623,In_408);
nor U39 (N_39,In_482,In_901);
nand U40 (N_40,In_272,In_60);
nor U41 (N_41,In_172,In_985);
or U42 (N_42,In_876,In_135);
or U43 (N_43,In_532,In_505);
or U44 (N_44,In_277,In_569);
or U45 (N_45,In_640,In_508);
nor U46 (N_46,In_609,In_231);
and U47 (N_47,In_126,In_754);
and U48 (N_48,In_762,In_506);
nor U49 (N_49,In_761,In_340);
nor U50 (N_50,In_701,In_648);
and U51 (N_51,In_200,In_784);
nor U52 (N_52,In_629,In_227);
nor U53 (N_53,In_436,In_655);
nor U54 (N_54,In_45,In_702);
nor U55 (N_55,In_734,In_144);
and U56 (N_56,In_44,In_28);
nand U57 (N_57,In_974,In_261);
nor U58 (N_58,In_121,In_134);
nor U59 (N_59,In_169,In_971);
or U60 (N_60,In_427,In_865);
nor U61 (N_61,In_793,In_571);
nand U62 (N_62,In_829,In_21);
and U63 (N_63,In_599,In_187);
or U64 (N_64,In_107,In_907);
and U65 (N_65,In_666,In_916);
nor U66 (N_66,In_385,In_360);
and U67 (N_67,In_746,In_168);
or U68 (N_68,In_315,In_950);
nand U69 (N_69,In_370,In_428);
and U70 (N_70,In_145,In_292);
and U71 (N_71,In_774,In_53);
nor U72 (N_72,In_893,In_996);
nand U73 (N_73,In_429,In_151);
nor U74 (N_74,In_912,In_539);
or U75 (N_75,In_303,In_296);
and U76 (N_76,In_987,In_649);
nor U77 (N_77,In_782,In_727);
nand U78 (N_78,In_725,In_405);
or U79 (N_79,In_119,In_517);
and U80 (N_80,In_35,In_103);
nand U81 (N_81,In_619,In_304);
nor U82 (N_82,In_219,In_80);
nand U83 (N_83,In_323,In_201);
nand U84 (N_84,In_495,In_170);
or U85 (N_85,In_889,In_764);
and U86 (N_86,In_438,In_65);
nand U87 (N_87,In_935,In_92);
nor U88 (N_88,In_471,In_536);
nor U89 (N_89,In_91,In_0);
or U90 (N_90,In_739,In_736);
nand U91 (N_91,In_554,In_377);
nor U92 (N_92,In_910,In_812);
nand U93 (N_93,In_616,In_690);
nor U94 (N_94,In_478,In_735);
nor U95 (N_95,In_982,In_937);
nor U96 (N_96,In_869,In_731);
and U97 (N_97,In_693,In_887);
nand U98 (N_98,In_980,In_620);
xor U99 (N_99,In_976,In_826);
nor U100 (N_100,In_673,In_513);
nor U101 (N_101,In_936,In_326);
nand U102 (N_102,In_286,In_274);
or U103 (N_103,In_417,In_259);
nand U104 (N_104,In_207,In_424);
and U105 (N_105,In_464,In_660);
nor U106 (N_106,In_983,In_663);
nand U107 (N_107,In_444,In_493);
nand U108 (N_108,In_290,In_546);
or U109 (N_109,In_249,In_115);
nor U110 (N_110,In_988,In_596);
nand U111 (N_111,In_755,In_205);
and U112 (N_112,In_575,In_266);
and U113 (N_113,In_15,In_827);
nor U114 (N_114,In_338,In_952);
or U115 (N_115,In_819,In_969);
nor U116 (N_116,In_551,In_716);
nor U117 (N_117,In_542,In_919);
nor U118 (N_118,In_462,In_209);
nand U119 (N_119,In_34,In_838);
and U120 (N_120,In_267,In_737);
and U121 (N_121,In_839,In_713);
nor U122 (N_122,In_572,In_563);
nand U123 (N_123,In_485,In_503);
and U124 (N_124,In_669,In_959);
nand U125 (N_125,In_548,In_589);
nor U126 (N_126,In_242,In_617);
and U127 (N_127,In_501,In_389);
or U128 (N_128,In_431,In_36);
or U129 (N_129,In_788,In_940);
or U130 (N_130,In_89,In_677);
and U131 (N_131,In_473,In_280);
and U132 (N_132,In_559,In_371);
or U133 (N_133,In_946,In_23);
nor U134 (N_134,In_264,In_351);
and U135 (N_135,In_738,In_341);
nor U136 (N_136,In_911,In_415);
nor U137 (N_137,In_73,In_275);
or U138 (N_138,In_419,In_239);
nor U139 (N_139,In_885,In_81);
nand U140 (N_140,In_997,In_871);
or U141 (N_141,In_88,In_857);
or U142 (N_142,In_844,In_566);
nand U143 (N_143,In_357,In_855);
or U144 (N_144,In_216,In_842);
and U145 (N_145,In_720,In_349);
or U146 (N_146,In_260,In_872);
or U147 (N_147,In_703,In_777);
nand U148 (N_148,In_153,In_120);
nor U149 (N_149,In_7,In_49);
or U150 (N_150,In_306,In_704);
or U151 (N_151,In_248,In_918);
and U152 (N_152,In_376,In_156);
nor U153 (N_153,In_711,In_378);
or U154 (N_154,In_874,In_480);
nand U155 (N_155,In_101,In_97);
or U156 (N_156,In_171,In_30);
nor U157 (N_157,In_366,In_769);
nor U158 (N_158,In_553,In_133);
nand U159 (N_159,In_850,In_832);
nor U160 (N_160,In_710,In_317);
xnor U161 (N_161,In_84,In_469);
nor U162 (N_162,In_615,In_198);
or U163 (N_163,In_387,In_598);
nor U164 (N_164,In_155,In_964);
nor U165 (N_165,In_752,In_500);
or U166 (N_166,In_320,In_468);
nor U167 (N_167,In_128,In_421);
nand U168 (N_168,In_287,In_318);
nand U169 (N_169,In_886,In_676);
or U170 (N_170,In_509,In_197);
nor U171 (N_171,In_805,In_833);
or U172 (N_172,In_443,In_434);
and U173 (N_173,In_61,In_582);
or U174 (N_174,In_772,In_557);
or U175 (N_175,In_890,In_140);
and U176 (N_176,In_333,In_526);
or U177 (N_177,In_581,In_496);
nor U178 (N_178,In_6,In_519);
and U179 (N_179,In_131,In_82);
nor U180 (N_180,In_866,In_226);
nand U181 (N_181,In_815,In_18);
or U182 (N_182,In_399,In_797);
nor U183 (N_183,In_373,In_270);
xor U184 (N_184,In_564,In_977);
xnor U185 (N_185,In_743,In_196);
or U186 (N_186,In_917,In_892);
and U187 (N_187,In_531,In_671);
nand U188 (N_188,In_268,In_386);
nor U189 (N_189,In_58,In_760);
and U190 (N_190,In_477,In_873);
and U191 (N_191,In_689,In_520);
and U192 (N_192,In_347,In_597);
or U193 (N_193,In_423,In_236);
or U194 (N_194,In_262,In_861);
or U195 (N_195,In_939,In_411);
nor U196 (N_196,In_860,In_214);
and U197 (N_197,In_973,In_185);
or U198 (N_198,In_282,In_125);
nor U199 (N_199,In_359,In_828);
nor U200 (N_200,In_608,In_740);
nor U201 (N_201,In_159,In_765);
nand U202 (N_202,In_729,In_147);
and U203 (N_203,In_285,In_184);
and U204 (N_204,In_382,In_281);
and U205 (N_205,In_13,In_954);
and U206 (N_206,In_612,In_409);
or U207 (N_207,In_926,In_646);
and U208 (N_208,In_442,In_8);
and U209 (N_209,In_297,In_83);
and U210 (N_210,In_179,In_110);
or U211 (N_211,In_858,In_55);
nand U212 (N_212,In_915,In_342);
or U213 (N_213,In_695,In_149);
nand U214 (N_214,In_237,In_990);
or U215 (N_215,In_961,In_803);
or U216 (N_216,In_903,In_957);
or U217 (N_217,In_447,In_524);
or U218 (N_218,In_194,In_979);
and U219 (N_219,In_20,In_692);
or U220 (N_220,In_204,In_358);
and U221 (N_221,In_899,In_220);
and U222 (N_222,In_218,In_694);
nand U223 (N_223,In_263,In_851);
and U224 (N_224,In_700,In_426);
nand U225 (N_225,In_484,In_780);
nor U226 (N_226,In_552,In_404);
and U227 (N_227,In_158,In_331);
and U228 (N_228,In_502,In_927);
or U229 (N_229,In_641,In_779);
and U230 (N_230,In_681,In_246);
or U231 (N_231,In_883,In_654);
nand U232 (N_232,In_470,In_944);
or U233 (N_233,In_163,In_813);
nor U234 (N_234,In_820,In_512);
nand U235 (N_235,In_191,In_733);
and U236 (N_236,In_778,In_71);
or U237 (N_237,In_391,In_25);
nand U238 (N_238,In_435,In_223);
or U239 (N_239,In_230,In_11);
nand U240 (N_240,In_560,In_487);
nor U241 (N_241,In_814,In_79);
and U242 (N_242,In_661,In_369);
nand U243 (N_243,In_806,In_425);
nand U244 (N_244,In_488,In_621);
or U245 (N_245,In_322,In_837);
or U246 (N_246,In_610,In_454);
or U247 (N_247,In_875,In_458);
nor U248 (N_248,In_356,In_241);
and U249 (N_249,In_580,In_213);
nand U250 (N_250,In_398,In_16);
nor U251 (N_251,In_537,In_474);
and U252 (N_252,In_76,In_934);
nor U253 (N_253,In_578,In_909);
nand U254 (N_254,In_544,In_402);
nor U255 (N_255,In_776,In_709);
nor U256 (N_256,In_794,In_476);
or U257 (N_257,In_38,In_452);
or U258 (N_258,In_515,In_117);
and U259 (N_259,In_483,In_416);
nor U260 (N_260,In_161,In_657);
nand U261 (N_261,In_407,In_978);
nand U262 (N_262,In_309,In_966);
and U263 (N_263,In_384,In_283);
nand U264 (N_264,In_183,In_632);
nand U265 (N_265,In_664,In_111);
or U266 (N_266,In_577,In_998);
nand U267 (N_267,In_522,In_527);
or U268 (N_268,In_991,In_699);
nand U269 (N_269,In_529,In_863);
nand U270 (N_270,In_822,In_634);
and U271 (N_271,In_148,In_37);
and U272 (N_272,In_307,In_400);
or U273 (N_273,In_606,In_523);
nor U274 (N_274,In_708,In_69);
nand U275 (N_275,In_334,In_714);
nand U276 (N_276,In_439,In_583);
nand U277 (N_277,In_51,In_698);
and U278 (N_278,In_186,In_335);
nand U279 (N_279,In_904,In_301);
and U280 (N_280,In_561,In_706);
nor U281 (N_281,In_138,In_771);
nand U282 (N_282,In_339,In_795);
nor U283 (N_283,In_674,In_630);
nor U284 (N_284,In_593,In_511);
nand U285 (N_285,In_251,In_984);
and U286 (N_286,In_662,In_445);
and U287 (N_287,In_12,In_178);
nor U288 (N_288,In_289,In_951);
nand U289 (N_289,In_933,In_925);
nor U290 (N_290,In_365,In_176);
nand U291 (N_291,In_809,In_109);
nand U292 (N_292,In_106,In_59);
nand U293 (N_293,In_122,In_127);
or U294 (N_294,In_210,In_897);
nor U295 (N_295,In_570,In_799);
and U296 (N_296,In_636,In_792);
and U297 (N_297,In_942,In_245);
nand U298 (N_298,In_217,In_556);
and U299 (N_299,In_528,In_968);
or U300 (N_300,In_77,In_175);
nor U301 (N_301,In_767,In_362);
nand U302 (N_302,In_879,In_541);
nand U303 (N_303,In_459,In_401);
and U304 (N_304,In_229,In_234);
and U305 (N_305,In_328,In_651);
nor U306 (N_306,In_880,In_24);
nand U307 (N_307,In_228,In_626);
or U308 (N_308,In_255,In_816);
and U309 (N_309,In_412,In_123);
and U310 (N_310,In_913,In_642);
xor U311 (N_311,In_896,In_291);
nand U312 (N_312,In_852,In_46);
nand U313 (N_313,In_540,In_108);
or U314 (N_314,In_825,In_414);
and U315 (N_315,In_258,In_273);
and U316 (N_316,In_167,In_222);
nand U317 (N_317,In_22,In_675);
nand U318 (N_318,In_584,In_202);
nor U319 (N_319,In_848,In_811);
nand U320 (N_320,In_3,In_271);
and U321 (N_321,In_905,In_243);
nor U322 (N_322,In_807,In_862);
or U323 (N_323,In_203,In_265);
nand U324 (N_324,In_457,In_497);
or U325 (N_325,In_643,In_50);
nand U326 (N_326,In_836,In_87);
and U327 (N_327,In_240,In_90);
and U328 (N_328,In_891,In_160);
and U329 (N_329,In_208,In_948);
nand U330 (N_330,In_392,In_679);
nand U331 (N_331,In_330,In_588);
and U332 (N_332,In_486,In_379);
and U333 (N_333,In_31,In_722);
nand U334 (N_334,In_63,In_975);
and U335 (N_335,In_830,In_723);
or U336 (N_336,In_164,In_374);
nand U337 (N_337,In_372,In_42);
nor U338 (N_338,In_574,In_321);
nor U339 (N_339,In_96,In_380);
nor U340 (N_340,In_19,In_849);
nand U341 (N_341,In_136,In_656);
and U342 (N_342,In_845,In_105);
nor U343 (N_343,In_549,In_510);
nor U344 (N_344,In_895,In_545);
nand U345 (N_345,In_902,In_678);
nand U346 (N_346,In_56,In_930);
and U347 (N_347,In_461,In_965);
or U348 (N_348,In_295,In_637);
or U349 (N_349,In_749,In_667);
or U350 (N_350,In_152,In_305);
and U351 (N_351,In_898,In_450);
nand U352 (N_352,In_361,In_573);
nand U353 (N_353,In_352,In_253);
or U354 (N_354,In_141,In_192);
nand U355 (N_355,In_41,In_162);
nor U356 (N_356,In_565,In_453);
and U357 (N_357,In_48,In_177);
nor U358 (N_358,In_972,In_579);
and U359 (N_359,In_252,In_166);
nand U360 (N_360,In_100,In_943);
and U361 (N_361,In_397,In_319);
nor U362 (N_362,In_688,In_768);
or U363 (N_363,In_601,In_718);
or U364 (N_364,In_2,In_215);
nand U365 (N_365,In_78,In_659);
xor U366 (N_366,In_62,In_312);
and U367 (N_367,In_460,In_142);
or U368 (N_368,In_113,In_324);
or U369 (N_369,In_888,In_489);
and U370 (N_370,In_894,In_864);
nand U371 (N_371,In_550,In_810);
and U372 (N_372,In_293,In_514);
or U373 (N_373,In_691,In_420);
nand U374 (N_374,In_586,In_254);
nand U375 (N_375,In_250,In_85);
nand U376 (N_376,In_66,In_441);
or U377 (N_377,In_817,In_668);
or U378 (N_378,In_576,In_99);
nor U379 (N_379,In_75,In_143);
and U380 (N_380,In_992,In_354);
nor U381 (N_381,In_390,In_472);
nor U382 (N_382,In_276,In_150);
nor U383 (N_383,In_114,In_381);
or U384 (N_384,In_685,In_786);
or U385 (N_385,In_70,In_783);
and U386 (N_386,In_644,In_790);
nor U387 (N_387,In_481,In_967);
and U388 (N_388,In_840,In_32);
or U389 (N_389,In_884,In_555);
or U390 (N_390,In_190,In_67);
xnor U391 (N_391,In_921,In_658);
and U392 (N_392,In_530,In_375);
nor U393 (N_393,In_211,In_986);
or U394 (N_394,In_494,In_635);
or U395 (N_395,In_298,In_970);
and U396 (N_396,In_336,In_52);
and U397 (N_397,In_95,In_17);
or U398 (N_398,In_602,In_345);
and U399 (N_399,In_614,In_538);
nor U400 (N_400,In_789,In_900);
or U401 (N_401,In_707,In_174);
nand U402 (N_402,In_173,In_525);
nor U403 (N_403,In_928,In_947);
or U404 (N_404,In_129,In_856);
nand U405 (N_405,In_766,In_355);
or U406 (N_406,In_40,In_956);
nand U407 (N_407,In_344,In_504);
or U408 (N_408,In_451,In_633);
nor U409 (N_409,In_313,In_748);
nor U410 (N_410,In_631,In_995);
nor U411 (N_411,In_802,In_39);
or U412 (N_412,In_232,In_449);
nor U413 (N_413,In_697,In_963);
and U414 (N_414,In_72,In_665);
and U415 (N_415,In_724,In_257);
and U416 (N_416,In_567,In_906);
or U417 (N_417,In_364,In_763);
or U418 (N_418,In_962,In_499);
nor U419 (N_419,In_432,In_279);
and U420 (N_420,In_410,In_47);
nor U421 (N_421,In_924,In_139);
nand U422 (N_422,In_638,In_941);
and U423 (N_423,In_302,In_757);
or U424 (N_424,In_853,In_953);
nor U425 (N_425,In_604,In_195);
nand U426 (N_426,In_796,In_433);
or U427 (N_427,In_74,In_300);
nor U428 (N_428,In_847,In_413);
nand U429 (N_429,In_193,In_235);
or U430 (N_430,In_773,In_846);
and U431 (N_431,In_299,In_741);
or U432 (N_432,In_353,In_112);
nand U433 (N_433,In_337,In_756);
or U434 (N_434,In_294,In_94);
nor U435 (N_435,In_465,In_627);
nor U436 (N_436,In_696,In_800);
and U437 (N_437,In_721,In_868);
nand U438 (N_438,In_247,In_914);
nand U439 (N_439,In_683,In_93);
and U440 (N_440,In_877,In_118);
nand U441 (N_441,In_329,In_745);
nand U442 (N_442,In_422,In_396);
nor U443 (N_443,In_124,In_653);
and U444 (N_444,In_348,In_945);
and U445 (N_445,In_682,In_920);
or U446 (N_446,In_467,In_613);
or U447 (N_447,In_278,In_587);
nand U448 (N_448,In_955,In_931);
and U449 (N_449,In_605,In_821);
nand U450 (N_450,In_180,In_33);
or U451 (N_451,In_728,In_558);
nand U452 (N_452,In_43,In_835);
nand U453 (N_453,In_463,In_9);
and U454 (N_454,In_647,In_680);
or U455 (N_455,In_750,In_818);
nand U456 (N_456,In_622,In_181);
or U457 (N_457,In_137,In_14);
or U458 (N_458,In_368,In_98);
nand U459 (N_459,In_625,In_687);
and U460 (N_460,In_116,In_715);
nor U461 (N_461,In_785,In_238);
nand U462 (N_462,In_929,In_878);
or U463 (N_463,In_686,In_533);
nor U464 (N_464,In_843,In_600);
nor U465 (N_465,In_516,In_932);
or U466 (N_466,In_5,In_834);
or U467 (N_467,In_645,In_466);
nand U468 (N_468,In_448,In_791);
nand U469 (N_469,In_4,In_595);
xnor U470 (N_470,In_29,In_490);
nor U471 (N_471,In_759,In_993);
xnor U472 (N_472,In_406,In_57);
nor U473 (N_473,In_981,In_753);
nand U474 (N_474,In_403,In_269);
nand U475 (N_475,In_343,In_994);
xnor U476 (N_476,In_224,In_591);
or U477 (N_477,In_672,In_189);
nand U478 (N_478,In_787,In_922);
and U479 (N_479,In_383,In_562);
nand U480 (N_480,In_518,In_521);
nand U481 (N_481,In_781,In_418);
and U482 (N_482,In_346,In_870);
and U483 (N_483,In_440,In_590);
or U484 (N_484,In_146,In_938);
nor U485 (N_485,In_350,In_798);
nor U486 (N_486,In_104,In_437);
nor U487 (N_487,In_288,In_68);
and U488 (N_488,In_859,In_182);
and U489 (N_489,In_854,In_206);
and U490 (N_490,In_10,In_824);
nand U491 (N_491,In_314,In_949);
or U492 (N_492,In_618,In_543);
nor U493 (N_493,In_960,In_26);
or U494 (N_494,In_130,In_717);
nand U495 (N_495,In_535,In_507);
or U496 (N_496,In_310,In_823);
or U497 (N_497,In_719,In_327);
or U498 (N_498,In_199,In_430);
or U499 (N_499,In_456,In_534);
nor U500 (N_500,In_164,In_773);
nor U501 (N_501,In_97,In_714);
and U502 (N_502,In_75,In_81);
nand U503 (N_503,In_538,In_466);
nor U504 (N_504,In_746,In_987);
and U505 (N_505,In_107,In_654);
and U506 (N_506,In_715,In_44);
nor U507 (N_507,In_718,In_211);
nand U508 (N_508,In_322,In_291);
and U509 (N_509,In_695,In_942);
and U510 (N_510,In_724,In_909);
nand U511 (N_511,In_633,In_853);
nor U512 (N_512,In_904,In_974);
and U513 (N_513,In_119,In_543);
and U514 (N_514,In_841,In_953);
nor U515 (N_515,In_839,In_539);
or U516 (N_516,In_993,In_999);
nand U517 (N_517,In_418,In_216);
nand U518 (N_518,In_166,In_632);
nor U519 (N_519,In_730,In_814);
and U520 (N_520,In_495,In_457);
nand U521 (N_521,In_22,In_350);
or U522 (N_522,In_342,In_984);
or U523 (N_523,In_428,In_512);
nor U524 (N_524,In_911,In_651);
nor U525 (N_525,In_481,In_302);
and U526 (N_526,In_160,In_808);
or U527 (N_527,In_986,In_814);
nand U528 (N_528,In_675,In_919);
nor U529 (N_529,In_885,In_159);
nand U530 (N_530,In_673,In_808);
nor U531 (N_531,In_575,In_43);
nand U532 (N_532,In_347,In_901);
and U533 (N_533,In_431,In_96);
nor U534 (N_534,In_356,In_295);
nand U535 (N_535,In_948,In_955);
or U536 (N_536,In_649,In_886);
and U537 (N_537,In_148,In_14);
nand U538 (N_538,In_527,In_476);
nor U539 (N_539,In_636,In_336);
or U540 (N_540,In_468,In_697);
nor U541 (N_541,In_939,In_654);
nor U542 (N_542,In_271,In_320);
nand U543 (N_543,In_40,In_916);
nand U544 (N_544,In_650,In_266);
or U545 (N_545,In_624,In_961);
and U546 (N_546,In_868,In_607);
or U547 (N_547,In_807,In_885);
nor U548 (N_548,In_885,In_476);
and U549 (N_549,In_316,In_788);
or U550 (N_550,In_565,In_332);
nand U551 (N_551,In_865,In_657);
xnor U552 (N_552,In_870,In_679);
and U553 (N_553,In_991,In_202);
and U554 (N_554,In_238,In_426);
and U555 (N_555,In_366,In_916);
nor U556 (N_556,In_453,In_907);
nand U557 (N_557,In_324,In_512);
and U558 (N_558,In_819,In_74);
and U559 (N_559,In_143,In_276);
nor U560 (N_560,In_118,In_529);
nor U561 (N_561,In_956,In_155);
or U562 (N_562,In_439,In_946);
and U563 (N_563,In_951,In_689);
nand U564 (N_564,In_276,In_666);
nand U565 (N_565,In_512,In_754);
or U566 (N_566,In_507,In_786);
xor U567 (N_567,In_556,In_352);
nand U568 (N_568,In_697,In_333);
nand U569 (N_569,In_674,In_110);
nand U570 (N_570,In_953,In_607);
and U571 (N_571,In_436,In_525);
nand U572 (N_572,In_308,In_274);
or U573 (N_573,In_254,In_769);
nor U574 (N_574,In_120,In_52);
nand U575 (N_575,In_618,In_161);
nand U576 (N_576,In_69,In_665);
and U577 (N_577,In_66,In_282);
and U578 (N_578,In_330,In_406);
nor U579 (N_579,In_627,In_51);
nand U580 (N_580,In_479,In_723);
nand U581 (N_581,In_277,In_982);
or U582 (N_582,In_370,In_455);
and U583 (N_583,In_222,In_907);
or U584 (N_584,In_102,In_264);
and U585 (N_585,In_955,In_499);
nor U586 (N_586,In_274,In_925);
and U587 (N_587,In_283,In_240);
or U588 (N_588,In_793,In_12);
nor U589 (N_589,In_530,In_579);
nor U590 (N_590,In_346,In_831);
nor U591 (N_591,In_740,In_864);
or U592 (N_592,In_43,In_998);
nand U593 (N_593,In_399,In_515);
nor U594 (N_594,In_905,In_674);
nor U595 (N_595,In_939,In_862);
nor U596 (N_596,In_560,In_417);
nor U597 (N_597,In_327,In_226);
nor U598 (N_598,In_709,In_290);
nor U599 (N_599,In_675,In_409);
nor U600 (N_600,In_204,In_562);
nor U601 (N_601,In_936,In_286);
nand U602 (N_602,In_266,In_101);
nand U603 (N_603,In_818,In_106);
and U604 (N_604,In_814,In_941);
or U605 (N_605,In_14,In_86);
or U606 (N_606,In_194,In_882);
and U607 (N_607,In_867,In_881);
nand U608 (N_608,In_210,In_313);
and U609 (N_609,In_708,In_89);
nand U610 (N_610,In_652,In_644);
and U611 (N_611,In_464,In_363);
and U612 (N_612,In_6,In_142);
nor U613 (N_613,In_503,In_614);
nand U614 (N_614,In_768,In_839);
or U615 (N_615,In_439,In_62);
and U616 (N_616,In_929,In_329);
nand U617 (N_617,In_989,In_223);
and U618 (N_618,In_99,In_954);
nand U619 (N_619,In_225,In_473);
and U620 (N_620,In_17,In_329);
nand U621 (N_621,In_840,In_885);
nand U622 (N_622,In_909,In_26);
nand U623 (N_623,In_357,In_305);
and U624 (N_624,In_684,In_10);
xnor U625 (N_625,In_891,In_831);
or U626 (N_626,In_161,In_92);
xnor U627 (N_627,In_731,In_907);
nor U628 (N_628,In_867,In_813);
nor U629 (N_629,In_334,In_367);
nor U630 (N_630,In_419,In_889);
and U631 (N_631,In_684,In_132);
nor U632 (N_632,In_692,In_92);
xor U633 (N_633,In_970,In_255);
nor U634 (N_634,In_180,In_939);
and U635 (N_635,In_887,In_453);
nor U636 (N_636,In_176,In_36);
and U637 (N_637,In_437,In_192);
nor U638 (N_638,In_942,In_986);
or U639 (N_639,In_72,In_115);
nor U640 (N_640,In_749,In_719);
nand U641 (N_641,In_479,In_573);
nor U642 (N_642,In_387,In_201);
nand U643 (N_643,In_851,In_29);
and U644 (N_644,In_563,In_378);
nand U645 (N_645,In_387,In_934);
nand U646 (N_646,In_692,In_294);
nor U647 (N_647,In_634,In_202);
nand U648 (N_648,In_569,In_688);
nand U649 (N_649,In_220,In_560);
nand U650 (N_650,In_268,In_853);
nor U651 (N_651,In_146,In_974);
nand U652 (N_652,In_333,In_906);
nor U653 (N_653,In_868,In_990);
nand U654 (N_654,In_604,In_491);
nor U655 (N_655,In_660,In_629);
and U656 (N_656,In_857,In_747);
nand U657 (N_657,In_569,In_28);
or U658 (N_658,In_99,In_40);
and U659 (N_659,In_212,In_775);
nor U660 (N_660,In_872,In_828);
and U661 (N_661,In_853,In_531);
nor U662 (N_662,In_331,In_49);
and U663 (N_663,In_6,In_951);
or U664 (N_664,In_776,In_397);
nand U665 (N_665,In_13,In_921);
nand U666 (N_666,In_127,In_24);
nand U667 (N_667,In_82,In_287);
or U668 (N_668,In_673,In_420);
nor U669 (N_669,In_989,In_58);
nor U670 (N_670,In_178,In_716);
nor U671 (N_671,In_208,In_268);
or U672 (N_672,In_548,In_663);
nor U673 (N_673,In_920,In_814);
nor U674 (N_674,In_882,In_931);
nor U675 (N_675,In_509,In_805);
nand U676 (N_676,In_264,In_558);
and U677 (N_677,In_531,In_196);
and U678 (N_678,In_337,In_454);
nor U679 (N_679,In_410,In_576);
or U680 (N_680,In_714,In_818);
or U681 (N_681,In_690,In_498);
or U682 (N_682,In_313,In_610);
nor U683 (N_683,In_657,In_600);
nor U684 (N_684,In_87,In_777);
or U685 (N_685,In_869,In_629);
and U686 (N_686,In_942,In_128);
nand U687 (N_687,In_200,In_261);
and U688 (N_688,In_715,In_271);
nor U689 (N_689,In_917,In_885);
and U690 (N_690,In_402,In_415);
and U691 (N_691,In_984,In_270);
nand U692 (N_692,In_785,In_999);
nand U693 (N_693,In_142,In_35);
and U694 (N_694,In_85,In_781);
nand U695 (N_695,In_760,In_804);
and U696 (N_696,In_84,In_570);
nor U697 (N_697,In_62,In_636);
xnor U698 (N_698,In_786,In_132);
or U699 (N_699,In_579,In_951);
or U700 (N_700,In_151,In_744);
and U701 (N_701,In_217,In_11);
and U702 (N_702,In_563,In_333);
or U703 (N_703,In_187,In_968);
nor U704 (N_704,In_305,In_546);
or U705 (N_705,In_562,In_419);
and U706 (N_706,In_497,In_227);
or U707 (N_707,In_9,In_967);
nand U708 (N_708,In_897,In_735);
nor U709 (N_709,In_38,In_955);
xnor U710 (N_710,In_810,In_872);
nand U711 (N_711,In_579,In_195);
nor U712 (N_712,In_212,In_443);
nand U713 (N_713,In_581,In_91);
nand U714 (N_714,In_217,In_133);
or U715 (N_715,In_532,In_543);
and U716 (N_716,In_128,In_928);
nand U717 (N_717,In_280,In_606);
nor U718 (N_718,In_255,In_953);
nor U719 (N_719,In_542,In_475);
nor U720 (N_720,In_182,In_578);
and U721 (N_721,In_768,In_400);
nand U722 (N_722,In_671,In_703);
or U723 (N_723,In_929,In_218);
and U724 (N_724,In_277,In_858);
or U725 (N_725,In_882,In_820);
or U726 (N_726,In_493,In_317);
or U727 (N_727,In_859,In_714);
nor U728 (N_728,In_641,In_659);
and U729 (N_729,In_164,In_743);
and U730 (N_730,In_661,In_561);
nor U731 (N_731,In_124,In_816);
nand U732 (N_732,In_485,In_671);
or U733 (N_733,In_291,In_765);
and U734 (N_734,In_181,In_257);
or U735 (N_735,In_497,In_567);
or U736 (N_736,In_279,In_756);
and U737 (N_737,In_436,In_929);
and U738 (N_738,In_488,In_252);
or U739 (N_739,In_224,In_29);
and U740 (N_740,In_706,In_916);
or U741 (N_741,In_710,In_356);
or U742 (N_742,In_928,In_977);
and U743 (N_743,In_909,In_650);
nor U744 (N_744,In_961,In_394);
nor U745 (N_745,In_589,In_141);
nor U746 (N_746,In_511,In_952);
nor U747 (N_747,In_981,In_130);
nand U748 (N_748,In_556,In_969);
and U749 (N_749,In_39,In_860);
and U750 (N_750,In_516,In_371);
or U751 (N_751,In_244,In_92);
or U752 (N_752,In_236,In_253);
and U753 (N_753,In_532,In_707);
xor U754 (N_754,In_475,In_223);
and U755 (N_755,In_470,In_899);
nor U756 (N_756,In_87,In_941);
nand U757 (N_757,In_918,In_956);
nand U758 (N_758,In_747,In_566);
nor U759 (N_759,In_713,In_142);
nand U760 (N_760,In_959,In_511);
or U761 (N_761,In_530,In_125);
and U762 (N_762,In_263,In_306);
nor U763 (N_763,In_615,In_16);
or U764 (N_764,In_340,In_933);
nor U765 (N_765,In_85,In_816);
nor U766 (N_766,In_983,In_875);
and U767 (N_767,In_458,In_564);
xor U768 (N_768,In_377,In_495);
nand U769 (N_769,In_996,In_256);
or U770 (N_770,In_131,In_652);
or U771 (N_771,In_609,In_755);
and U772 (N_772,In_913,In_667);
or U773 (N_773,In_176,In_871);
nor U774 (N_774,In_971,In_302);
nand U775 (N_775,In_742,In_682);
nand U776 (N_776,In_666,In_958);
nor U777 (N_777,In_810,In_633);
nor U778 (N_778,In_730,In_34);
nor U779 (N_779,In_734,In_504);
nand U780 (N_780,In_975,In_394);
nor U781 (N_781,In_675,In_86);
or U782 (N_782,In_404,In_941);
or U783 (N_783,In_42,In_57);
nand U784 (N_784,In_192,In_542);
nor U785 (N_785,In_66,In_330);
nor U786 (N_786,In_758,In_361);
nor U787 (N_787,In_86,In_511);
nor U788 (N_788,In_459,In_764);
nor U789 (N_789,In_554,In_373);
or U790 (N_790,In_269,In_263);
nor U791 (N_791,In_206,In_756);
nor U792 (N_792,In_2,In_164);
nand U793 (N_793,In_32,In_509);
and U794 (N_794,In_766,In_548);
and U795 (N_795,In_546,In_2);
nand U796 (N_796,In_482,In_375);
nand U797 (N_797,In_381,In_294);
nor U798 (N_798,In_587,In_18);
or U799 (N_799,In_119,In_846);
or U800 (N_800,In_530,In_613);
nor U801 (N_801,In_887,In_612);
or U802 (N_802,In_492,In_464);
and U803 (N_803,In_854,In_398);
nand U804 (N_804,In_218,In_530);
or U805 (N_805,In_373,In_338);
nand U806 (N_806,In_336,In_859);
nor U807 (N_807,In_58,In_643);
and U808 (N_808,In_639,In_719);
and U809 (N_809,In_988,In_90);
nand U810 (N_810,In_931,In_297);
or U811 (N_811,In_863,In_930);
and U812 (N_812,In_980,In_985);
nor U813 (N_813,In_238,In_887);
and U814 (N_814,In_785,In_46);
nand U815 (N_815,In_32,In_714);
or U816 (N_816,In_239,In_109);
and U817 (N_817,In_452,In_796);
nand U818 (N_818,In_433,In_594);
or U819 (N_819,In_874,In_758);
nand U820 (N_820,In_99,In_39);
and U821 (N_821,In_240,In_670);
or U822 (N_822,In_484,In_687);
or U823 (N_823,In_765,In_566);
or U824 (N_824,In_536,In_613);
and U825 (N_825,In_901,In_169);
nand U826 (N_826,In_685,In_429);
or U827 (N_827,In_2,In_993);
nor U828 (N_828,In_710,In_8);
nor U829 (N_829,In_790,In_245);
and U830 (N_830,In_387,In_26);
and U831 (N_831,In_320,In_418);
nand U832 (N_832,In_512,In_232);
and U833 (N_833,In_543,In_265);
nor U834 (N_834,In_882,In_791);
or U835 (N_835,In_428,In_409);
or U836 (N_836,In_317,In_700);
or U837 (N_837,In_251,In_823);
and U838 (N_838,In_361,In_982);
nand U839 (N_839,In_71,In_425);
nand U840 (N_840,In_625,In_632);
or U841 (N_841,In_413,In_614);
and U842 (N_842,In_879,In_305);
nand U843 (N_843,In_884,In_439);
and U844 (N_844,In_530,In_818);
or U845 (N_845,In_849,In_694);
or U846 (N_846,In_460,In_235);
and U847 (N_847,In_723,In_333);
nor U848 (N_848,In_214,In_322);
or U849 (N_849,In_628,In_609);
or U850 (N_850,In_886,In_859);
nor U851 (N_851,In_449,In_143);
nor U852 (N_852,In_618,In_781);
or U853 (N_853,In_162,In_396);
nand U854 (N_854,In_505,In_60);
and U855 (N_855,In_218,In_907);
nor U856 (N_856,In_956,In_204);
nand U857 (N_857,In_869,In_172);
or U858 (N_858,In_951,In_147);
nor U859 (N_859,In_203,In_372);
and U860 (N_860,In_746,In_792);
nand U861 (N_861,In_833,In_510);
nand U862 (N_862,In_50,In_429);
or U863 (N_863,In_887,In_753);
or U864 (N_864,In_959,In_210);
xnor U865 (N_865,In_366,In_747);
or U866 (N_866,In_457,In_565);
or U867 (N_867,In_103,In_826);
nand U868 (N_868,In_697,In_238);
nor U869 (N_869,In_142,In_364);
nand U870 (N_870,In_800,In_542);
and U871 (N_871,In_318,In_429);
nand U872 (N_872,In_478,In_957);
and U873 (N_873,In_961,In_354);
nand U874 (N_874,In_444,In_411);
nor U875 (N_875,In_318,In_649);
and U876 (N_876,In_173,In_110);
and U877 (N_877,In_932,In_372);
or U878 (N_878,In_263,In_475);
nand U879 (N_879,In_121,In_290);
and U880 (N_880,In_598,In_115);
and U881 (N_881,In_363,In_247);
or U882 (N_882,In_701,In_273);
nor U883 (N_883,In_764,In_796);
or U884 (N_884,In_953,In_173);
nor U885 (N_885,In_65,In_627);
or U886 (N_886,In_741,In_585);
or U887 (N_887,In_129,In_268);
nand U888 (N_888,In_53,In_790);
nor U889 (N_889,In_741,In_818);
and U890 (N_890,In_636,In_404);
nor U891 (N_891,In_979,In_357);
and U892 (N_892,In_766,In_710);
xor U893 (N_893,In_896,In_798);
and U894 (N_894,In_673,In_391);
or U895 (N_895,In_288,In_722);
nor U896 (N_896,In_675,In_269);
nand U897 (N_897,In_993,In_989);
nor U898 (N_898,In_665,In_697);
and U899 (N_899,In_977,In_247);
nand U900 (N_900,In_550,In_150);
nand U901 (N_901,In_178,In_240);
nor U902 (N_902,In_63,In_641);
and U903 (N_903,In_743,In_616);
nand U904 (N_904,In_562,In_158);
or U905 (N_905,In_978,In_690);
nand U906 (N_906,In_179,In_578);
or U907 (N_907,In_555,In_181);
nand U908 (N_908,In_995,In_404);
nand U909 (N_909,In_397,In_342);
or U910 (N_910,In_262,In_856);
or U911 (N_911,In_598,In_640);
nor U912 (N_912,In_51,In_942);
or U913 (N_913,In_264,In_965);
nand U914 (N_914,In_934,In_339);
and U915 (N_915,In_985,In_988);
nand U916 (N_916,In_832,In_190);
or U917 (N_917,In_13,In_885);
nor U918 (N_918,In_893,In_610);
nor U919 (N_919,In_642,In_15);
or U920 (N_920,In_539,In_950);
or U921 (N_921,In_876,In_914);
nor U922 (N_922,In_374,In_860);
and U923 (N_923,In_959,In_625);
and U924 (N_924,In_952,In_208);
or U925 (N_925,In_443,In_220);
or U926 (N_926,In_993,In_855);
nand U927 (N_927,In_310,In_943);
or U928 (N_928,In_254,In_629);
and U929 (N_929,In_522,In_24);
or U930 (N_930,In_635,In_236);
and U931 (N_931,In_5,In_522);
nand U932 (N_932,In_884,In_787);
and U933 (N_933,In_968,In_125);
or U934 (N_934,In_143,In_924);
nor U935 (N_935,In_796,In_431);
and U936 (N_936,In_254,In_293);
nor U937 (N_937,In_288,In_426);
and U938 (N_938,In_78,In_913);
nand U939 (N_939,In_396,In_113);
and U940 (N_940,In_620,In_774);
or U941 (N_941,In_510,In_982);
nor U942 (N_942,In_543,In_794);
nor U943 (N_943,In_42,In_19);
nand U944 (N_944,In_414,In_79);
nor U945 (N_945,In_667,In_22);
nor U946 (N_946,In_536,In_974);
nor U947 (N_947,In_297,In_154);
or U948 (N_948,In_719,In_118);
and U949 (N_949,In_875,In_661);
nor U950 (N_950,In_622,In_145);
nand U951 (N_951,In_837,In_736);
and U952 (N_952,In_737,In_677);
nand U953 (N_953,In_376,In_886);
nor U954 (N_954,In_39,In_156);
and U955 (N_955,In_228,In_243);
nand U956 (N_956,In_787,In_571);
nand U957 (N_957,In_731,In_622);
nor U958 (N_958,In_570,In_685);
and U959 (N_959,In_590,In_732);
nand U960 (N_960,In_193,In_678);
and U961 (N_961,In_371,In_266);
or U962 (N_962,In_767,In_542);
nor U963 (N_963,In_306,In_560);
and U964 (N_964,In_527,In_514);
nand U965 (N_965,In_864,In_190);
and U966 (N_966,In_833,In_826);
nor U967 (N_967,In_157,In_241);
nor U968 (N_968,In_800,In_678);
nand U969 (N_969,In_827,In_198);
nor U970 (N_970,In_220,In_26);
or U971 (N_971,In_234,In_412);
or U972 (N_972,In_41,In_406);
or U973 (N_973,In_86,In_216);
or U974 (N_974,In_905,In_57);
nand U975 (N_975,In_931,In_944);
or U976 (N_976,In_421,In_548);
and U977 (N_977,In_17,In_302);
nand U978 (N_978,In_268,In_270);
or U979 (N_979,In_676,In_285);
nor U980 (N_980,In_880,In_914);
nand U981 (N_981,In_731,In_818);
nand U982 (N_982,In_183,In_382);
nor U983 (N_983,In_829,In_797);
nor U984 (N_984,In_858,In_77);
nand U985 (N_985,In_740,In_762);
nand U986 (N_986,In_225,In_962);
and U987 (N_987,In_934,In_578);
nor U988 (N_988,In_673,In_427);
or U989 (N_989,In_546,In_594);
nor U990 (N_990,In_823,In_252);
and U991 (N_991,In_737,In_689);
nor U992 (N_992,In_936,In_156);
and U993 (N_993,In_728,In_770);
nor U994 (N_994,In_94,In_368);
and U995 (N_995,In_878,In_302);
and U996 (N_996,In_382,In_105);
nor U997 (N_997,In_460,In_90);
and U998 (N_998,In_221,In_49);
nand U999 (N_999,In_752,In_518);
or U1000 (N_1000,In_218,In_544);
nand U1001 (N_1001,In_477,In_461);
nand U1002 (N_1002,In_940,In_976);
or U1003 (N_1003,In_339,In_790);
or U1004 (N_1004,In_743,In_34);
nor U1005 (N_1005,In_938,In_612);
nand U1006 (N_1006,In_570,In_466);
nand U1007 (N_1007,In_812,In_615);
nor U1008 (N_1008,In_247,In_820);
nand U1009 (N_1009,In_453,In_567);
nor U1010 (N_1010,In_302,In_104);
nor U1011 (N_1011,In_745,In_727);
nand U1012 (N_1012,In_112,In_282);
nor U1013 (N_1013,In_510,In_48);
nor U1014 (N_1014,In_282,In_290);
or U1015 (N_1015,In_452,In_457);
and U1016 (N_1016,In_409,In_819);
or U1017 (N_1017,In_541,In_105);
and U1018 (N_1018,In_892,In_369);
nand U1019 (N_1019,In_42,In_609);
or U1020 (N_1020,In_992,In_763);
nand U1021 (N_1021,In_754,In_579);
or U1022 (N_1022,In_967,In_994);
nor U1023 (N_1023,In_18,In_764);
nor U1024 (N_1024,In_179,In_64);
or U1025 (N_1025,In_972,In_715);
nand U1026 (N_1026,In_298,In_788);
or U1027 (N_1027,In_579,In_34);
nand U1028 (N_1028,In_675,In_199);
and U1029 (N_1029,In_113,In_591);
nor U1030 (N_1030,In_661,In_220);
and U1031 (N_1031,In_145,In_662);
or U1032 (N_1032,In_214,In_384);
or U1033 (N_1033,In_489,In_175);
nor U1034 (N_1034,In_750,In_49);
and U1035 (N_1035,In_215,In_274);
and U1036 (N_1036,In_309,In_814);
and U1037 (N_1037,In_331,In_119);
nand U1038 (N_1038,In_713,In_261);
nor U1039 (N_1039,In_684,In_160);
or U1040 (N_1040,In_58,In_173);
nand U1041 (N_1041,In_415,In_414);
and U1042 (N_1042,In_878,In_423);
nor U1043 (N_1043,In_59,In_513);
and U1044 (N_1044,In_271,In_120);
and U1045 (N_1045,In_873,In_173);
or U1046 (N_1046,In_182,In_305);
or U1047 (N_1047,In_456,In_289);
or U1048 (N_1048,In_295,In_780);
or U1049 (N_1049,In_673,In_428);
nor U1050 (N_1050,In_831,In_414);
nor U1051 (N_1051,In_849,In_43);
nor U1052 (N_1052,In_428,In_362);
nor U1053 (N_1053,In_623,In_562);
nor U1054 (N_1054,In_797,In_531);
nor U1055 (N_1055,In_403,In_980);
nand U1056 (N_1056,In_706,In_94);
nand U1057 (N_1057,In_632,In_211);
or U1058 (N_1058,In_629,In_117);
or U1059 (N_1059,In_566,In_448);
nor U1060 (N_1060,In_657,In_831);
nor U1061 (N_1061,In_277,In_699);
nor U1062 (N_1062,In_863,In_199);
nor U1063 (N_1063,In_718,In_902);
and U1064 (N_1064,In_560,In_983);
nand U1065 (N_1065,In_18,In_126);
and U1066 (N_1066,In_193,In_412);
nor U1067 (N_1067,In_480,In_803);
nor U1068 (N_1068,In_809,In_498);
and U1069 (N_1069,In_650,In_926);
or U1070 (N_1070,In_570,In_211);
and U1071 (N_1071,In_303,In_275);
and U1072 (N_1072,In_95,In_907);
and U1073 (N_1073,In_555,In_810);
nor U1074 (N_1074,In_713,In_937);
and U1075 (N_1075,In_688,In_433);
or U1076 (N_1076,In_374,In_270);
nand U1077 (N_1077,In_770,In_947);
nand U1078 (N_1078,In_837,In_291);
nand U1079 (N_1079,In_122,In_96);
nor U1080 (N_1080,In_478,In_744);
nand U1081 (N_1081,In_673,In_456);
nand U1082 (N_1082,In_331,In_352);
nand U1083 (N_1083,In_681,In_186);
or U1084 (N_1084,In_757,In_637);
nand U1085 (N_1085,In_391,In_528);
or U1086 (N_1086,In_991,In_345);
or U1087 (N_1087,In_341,In_402);
and U1088 (N_1088,In_293,In_553);
or U1089 (N_1089,In_793,In_125);
nand U1090 (N_1090,In_782,In_843);
and U1091 (N_1091,In_548,In_62);
and U1092 (N_1092,In_854,In_249);
nand U1093 (N_1093,In_467,In_657);
nand U1094 (N_1094,In_214,In_373);
nor U1095 (N_1095,In_581,In_592);
nor U1096 (N_1096,In_36,In_803);
nor U1097 (N_1097,In_630,In_871);
and U1098 (N_1098,In_428,In_894);
nor U1099 (N_1099,In_61,In_855);
and U1100 (N_1100,In_987,In_442);
nor U1101 (N_1101,In_762,In_245);
nand U1102 (N_1102,In_888,In_212);
and U1103 (N_1103,In_48,In_731);
nor U1104 (N_1104,In_564,In_463);
or U1105 (N_1105,In_962,In_847);
nand U1106 (N_1106,In_620,In_400);
nand U1107 (N_1107,In_273,In_339);
and U1108 (N_1108,In_569,In_686);
or U1109 (N_1109,In_645,In_298);
nor U1110 (N_1110,In_297,In_590);
nand U1111 (N_1111,In_48,In_863);
and U1112 (N_1112,In_342,In_232);
or U1113 (N_1113,In_790,In_328);
or U1114 (N_1114,In_611,In_850);
and U1115 (N_1115,In_997,In_283);
or U1116 (N_1116,In_785,In_259);
and U1117 (N_1117,In_832,In_322);
nand U1118 (N_1118,In_517,In_456);
nor U1119 (N_1119,In_75,In_520);
and U1120 (N_1120,In_111,In_632);
nor U1121 (N_1121,In_636,In_638);
nor U1122 (N_1122,In_679,In_497);
and U1123 (N_1123,In_514,In_405);
or U1124 (N_1124,In_317,In_300);
and U1125 (N_1125,In_673,In_166);
or U1126 (N_1126,In_101,In_390);
and U1127 (N_1127,In_362,In_338);
nand U1128 (N_1128,In_543,In_700);
or U1129 (N_1129,In_227,In_212);
nor U1130 (N_1130,In_228,In_70);
nand U1131 (N_1131,In_583,In_661);
nor U1132 (N_1132,In_878,In_56);
nand U1133 (N_1133,In_989,In_440);
and U1134 (N_1134,In_797,In_123);
nand U1135 (N_1135,In_102,In_175);
or U1136 (N_1136,In_85,In_994);
nor U1137 (N_1137,In_105,In_538);
nand U1138 (N_1138,In_505,In_697);
or U1139 (N_1139,In_699,In_889);
and U1140 (N_1140,In_655,In_235);
or U1141 (N_1141,In_24,In_101);
or U1142 (N_1142,In_151,In_341);
or U1143 (N_1143,In_293,In_45);
nor U1144 (N_1144,In_159,In_890);
and U1145 (N_1145,In_231,In_361);
nand U1146 (N_1146,In_692,In_986);
xnor U1147 (N_1147,In_763,In_471);
nand U1148 (N_1148,In_936,In_25);
nor U1149 (N_1149,In_862,In_269);
or U1150 (N_1150,In_201,In_463);
nand U1151 (N_1151,In_465,In_433);
nand U1152 (N_1152,In_125,In_927);
nand U1153 (N_1153,In_946,In_283);
or U1154 (N_1154,In_47,In_824);
xnor U1155 (N_1155,In_980,In_859);
nor U1156 (N_1156,In_408,In_36);
nor U1157 (N_1157,In_960,In_915);
or U1158 (N_1158,In_57,In_675);
and U1159 (N_1159,In_346,In_569);
nand U1160 (N_1160,In_642,In_400);
and U1161 (N_1161,In_723,In_239);
nor U1162 (N_1162,In_549,In_123);
and U1163 (N_1163,In_455,In_294);
or U1164 (N_1164,In_881,In_684);
or U1165 (N_1165,In_476,In_976);
nand U1166 (N_1166,In_365,In_193);
and U1167 (N_1167,In_319,In_48);
nor U1168 (N_1168,In_384,In_579);
nor U1169 (N_1169,In_622,In_163);
or U1170 (N_1170,In_136,In_936);
nor U1171 (N_1171,In_556,In_673);
or U1172 (N_1172,In_361,In_83);
nand U1173 (N_1173,In_758,In_897);
or U1174 (N_1174,In_259,In_664);
nor U1175 (N_1175,In_48,In_375);
or U1176 (N_1176,In_556,In_851);
nand U1177 (N_1177,In_490,In_475);
xor U1178 (N_1178,In_27,In_924);
nor U1179 (N_1179,In_679,In_53);
nor U1180 (N_1180,In_981,In_514);
nor U1181 (N_1181,In_960,In_71);
nand U1182 (N_1182,In_44,In_40);
nand U1183 (N_1183,In_789,In_836);
and U1184 (N_1184,In_337,In_659);
or U1185 (N_1185,In_560,In_837);
or U1186 (N_1186,In_630,In_213);
and U1187 (N_1187,In_102,In_991);
nor U1188 (N_1188,In_119,In_855);
and U1189 (N_1189,In_100,In_394);
and U1190 (N_1190,In_147,In_652);
nor U1191 (N_1191,In_726,In_936);
and U1192 (N_1192,In_752,In_299);
and U1193 (N_1193,In_489,In_564);
or U1194 (N_1194,In_455,In_80);
and U1195 (N_1195,In_973,In_556);
nand U1196 (N_1196,In_668,In_747);
nor U1197 (N_1197,In_70,In_248);
nand U1198 (N_1198,In_263,In_332);
or U1199 (N_1199,In_119,In_521);
nand U1200 (N_1200,In_675,In_85);
and U1201 (N_1201,In_141,In_204);
and U1202 (N_1202,In_813,In_653);
nand U1203 (N_1203,In_881,In_381);
and U1204 (N_1204,In_389,In_27);
nor U1205 (N_1205,In_890,In_617);
or U1206 (N_1206,In_936,In_202);
and U1207 (N_1207,In_755,In_462);
and U1208 (N_1208,In_31,In_138);
nand U1209 (N_1209,In_530,In_854);
nor U1210 (N_1210,In_595,In_563);
or U1211 (N_1211,In_812,In_166);
or U1212 (N_1212,In_193,In_145);
and U1213 (N_1213,In_409,In_876);
nor U1214 (N_1214,In_40,In_724);
and U1215 (N_1215,In_729,In_739);
nand U1216 (N_1216,In_125,In_995);
nor U1217 (N_1217,In_205,In_750);
nor U1218 (N_1218,In_31,In_146);
and U1219 (N_1219,In_387,In_150);
or U1220 (N_1220,In_452,In_102);
nor U1221 (N_1221,In_613,In_497);
and U1222 (N_1222,In_551,In_553);
nor U1223 (N_1223,In_832,In_206);
and U1224 (N_1224,In_193,In_612);
nor U1225 (N_1225,In_620,In_635);
and U1226 (N_1226,In_724,In_225);
nor U1227 (N_1227,In_400,In_623);
and U1228 (N_1228,In_127,In_383);
nor U1229 (N_1229,In_289,In_622);
or U1230 (N_1230,In_970,In_799);
or U1231 (N_1231,In_32,In_684);
nor U1232 (N_1232,In_214,In_561);
nand U1233 (N_1233,In_693,In_607);
and U1234 (N_1234,In_978,In_394);
and U1235 (N_1235,In_738,In_615);
nor U1236 (N_1236,In_287,In_647);
or U1237 (N_1237,In_108,In_697);
or U1238 (N_1238,In_639,In_702);
nor U1239 (N_1239,In_751,In_538);
and U1240 (N_1240,In_937,In_809);
and U1241 (N_1241,In_629,In_250);
nand U1242 (N_1242,In_228,In_298);
nand U1243 (N_1243,In_262,In_320);
and U1244 (N_1244,In_614,In_945);
and U1245 (N_1245,In_429,In_24);
or U1246 (N_1246,In_494,In_318);
and U1247 (N_1247,In_148,In_416);
nand U1248 (N_1248,In_275,In_133);
nand U1249 (N_1249,In_250,In_102);
nor U1250 (N_1250,In_703,In_195);
or U1251 (N_1251,In_885,In_645);
or U1252 (N_1252,In_750,In_640);
or U1253 (N_1253,In_553,In_963);
or U1254 (N_1254,In_97,In_382);
nor U1255 (N_1255,In_308,In_74);
and U1256 (N_1256,In_850,In_241);
nand U1257 (N_1257,In_801,In_268);
nor U1258 (N_1258,In_378,In_771);
or U1259 (N_1259,In_531,In_837);
and U1260 (N_1260,In_38,In_291);
or U1261 (N_1261,In_418,In_403);
nor U1262 (N_1262,In_464,In_192);
and U1263 (N_1263,In_996,In_864);
and U1264 (N_1264,In_641,In_862);
nand U1265 (N_1265,In_698,In_170);
and U1266 (N_1266,In_535,In_134);
nand U1267 (N_1267,In_108,In_838);
or U1268 (N_1268,In_753,In_655);
and U1269 (N_1269,In_470,In_178);
and U1270 (N_1270,In_252,In_985);
or U1271 (N_1271,In_955,In_682);
and U1272 (N_1272,In_502,In_443);
nor U1273 (N_1273,In_635,In_323);
and U1274 (N_1274,In_577,In_623);
nor U1275 (N_1275,In_838,In_835);
or U1276 (N_1276,In_452,In_824);
and U1277 (N_1277,In_368,In_138);
and U1278 (N_1278,In_816,In_424);
and U1279 (N_1279,In_395,In_204);
nor U1280 (N_1280,In_287,In_123);
nand U1281 (N_1281,In_831,In_780);
or U1282 (N_1282,In_814,In_644);
nand U1283 (N_1283,In_604,In_44);
nand U1284 (N_1284,In_370,In_833);
and U1285 (N_1285,In_447,In_42);
or U1286 (N_1286,In_949,In_514);
nor U1287 (N_1287,In_235,In_116);
nand U1288 (N_1288,In_442,In_448);
or U1289 (N_1289,In_210,In_430);
or U1290 (N_1290,In_235,In_674);
and U1291 (N_1291,In_127,In_930);
and U1292 (N_1292,In_765,In_211);
or U1293 (N_1293,In_877,In_556);
nand U1294 (N_1294,In_610,In_729);
and U1295 (N_1295,In_167,In_372);
and U1296 (N_1296,In_951,In_628);
nand U1297 (N_1297,In_218,In_921);
nand U1298 (N_1298,In_383,In_591);
nor U1299 (N_1299,In_260,In_876);
nor U1300 (N_1300,In_997,In_594);
or U1301 (N_1301,In_681,In_687);
and U1302 (N_1302,In_126,In_535);
nor U1303 (N_1303,In_9,In_902);
and U1304 (N_1304,In_610,In_143);
and U1305 (N_1305,In_421,In_646);
nor U1306 (N_1306,In_238,In_745);
or U1307 (N_1307,In_674,In_63);
or U1308 (N_1308,In_709,In_256);
or U1309 (N_1309,In_585,In_2);
and U1310 (N_1310,In_214,In_221);
and U1311 (N_1311,In_974,In_611);
nand U1312 (N_1312,In_994,In_925);
and U1313 (N_1313,In_993,In_460);
nand U1314 (N_1314,In_706,In_345);
nand U1315 (N_1315,In_926,In_511);
nand U1316 (N_1316,In_418,In_996);
nand U1317 (N_1317,In_783,In_418);
or U1318 (N_1318,In_842,In_596);
nor U1319 (N_1319,In_967,In_460);
and U1320 (N_1320,In_603,In_75);
or U1321 (N_1321,In_301,In_156);
and U1322 (N_1322,In_425,In_185);
or U1323 (N_1323,In_903,In_102);
and U1324 (N_1324,In_900,In_600);
nor U1325 (N_1325,In_267,In_524);
xor U1326 (N_1326,In_583,In_463);
and U1327 (N_1327,In_219,In_310);
nand U1328 (N_1328,In_598,In_889);
nand U1329 (N_1329,In_589,In_697);
and U1330 (N_1330,In_290,In_657);
xnor U1331 (N_1331,In_302,In_584);
or U1332 (N_1332,In_228,In_553);
or U1333 (N_1333,In_627,In_310);
xnor U1334 (N_1334,In_397,In_437);
and U1335 (N_1335,In_708,In_710);
nor U1336 (N_1336,In_552,In_575);
or U1337 (N_1337,In_294,In_109);
nor U1338 (N_1338,In_164,In_241);
nor U1339 (N_1339,In_554,In_78);
nand U1340 (N_1340,In_796,In_266);
and U1341 (N_1341,In_504,In_590);
and U1342 (N_1342,In_357,In_89);
or U1343 (N_1343,In_624,In_657);
nor U1344 (N_1344,In_535,In_85);
nand U1345 (N_1345,In_218,In_141);
nand U1346 (N_1346,In_876,In_938);
or U1347 (N_1347,In_854,In_642);
and U1348 (N_1348,In_754,In_958);
nor U1349 (N_1349,In_779,In_464);
or U1350 (N_1350,In_724,In_231);
nand U1351 (N_1351,In_726,In_365);
or U1352 (N_1352,In_435,In_553);
nor U1353 (N_1353,In_858,In_366);
nor U1354 (N_1354,In_753,In_947);
nor U1355 (N_1355,In_104,In_808);
or U1356 (N_1356,In_241,In_183);
nor U1357 (N_1357,In_545,In_450);
and U1358 (N_1358,In_827,In_230);
nor U1359 (N_1359,In_48,In_266);
and U1360 (N_1360,In_122,In_581);
nor U1361 (N_1361,In_834,In_955);
and U1362 (N_1362,In_154,In_741);
nor U1363 (N_1363,In_87,In_935);
nand U1364 (N_1364,In_448,In_428);
nor U1365 (N_1365,In_426,In_372);
or U1366 (N_1366,In_39,In_600);
nand U1367 (N_1367,In_591,In_630);
nor U1368 (N_1368,In_441,In_684);
nand U1369 (N_1369,In_809,In_43);
and U1370 (N_1370,In_469,In_867);
or U1371 (N_1371,In_61,In_472);
nand U1372 (N_1372,In_701,In_469);
and U1373 (N_1373,In_779,In_286);
or U1374 (N_1374,In_919,In_698);
or U1375 (N_1375,In_176,In_30);
and U1376 (N_1376,In_301,In_777);
nand U1377 (N_1377,In_858,In_933);
nor U1378 (N_1378,In_664,In_333);
nand U1379 (N_1379,In_244,In_234);
nor U1380 (N_1380,In_512,In_734);
or U1381 (N_1381,In_731,In_134);
nor U1382 (N_1382,In_977,In_785);
or U1383 (N_1383,In_860,In_864);
nand U1384 (N_1384,In_162,In_816);
or U1385 (N_1385,In_247,In_448);
nor U1386 (N_1386,In_230,In_252);
nand U1387 (N_1387,In_325,In_408);
or U1388 (N_1388,In_528,In_998);
nand U1389 (N_1389,In_160,In_721);
or U1390 (N_1390,In_631,In_396);
nand U1391 (N_1391,In_649,In_306);
nand U1392 (N_1392,In_655,In_485);
nand U1393 (N_1393,In_261,In_663);
nand U1394 (N_1394,In_204,In_353);
or U1395 (N_1395,In_633,In_579);
and U1396 (N_1396,In_120,In_838);
or U1397 (N_1397,In_538,In_393);
and U1398 (N_1398,In_324,In_980);
and U1399 (N_1399,In_25,In_789);
nand U1400 (N_1400,In_584,In_795);
nor U1401 (N_1401,In_375,In_407);
and U1402 (N_1402,In_556,In_604);
nand U1403 (N_1403,In_818,In_805);
and U1404 (N_1404,In_953,In_889);
nand U1405 (N_1405,In_734,In_45);
and U1406 (N_1406,In_189,In_699);
and U1407 (N_1407,In_135,In_789);
nor U1408 (N_1408,In_551,In_800);
nor U1409 (N_1409,In_465,In_116);
nand U1410 (N_1410,In_973,In_529);
or U1411 (N_1411,In_92,In_726);
or U1412 (N_1412,In_56,In_501);
nor U1413 (N_1413,In_820,In_989);
and U1414 (N_1414,In_51,In_304);
and U1415 (N_1415,In_544,In_464);
nor U1416 (N_1416,In_986,In_741);
nand U1417 (N_1417,In_884,In_642);
and U1418 (N_1418,In_550,In_246);
and U1419 (N_1419,In_323,In_188);
nand U1420 (N_1420,In_858,In_388);
or U1421 (N_1421,In_164,In_610);
or U1422 (N_1422,In_232,In_369);
nand U1423 (N_1423,In_820,In_855);
and U1424 (N_1424,In_432,In_635);
nor U1425 (N_1425,In_525,In_121);
and U1426 (N_1426,In_722,In_468);
and U1427 (N_1427,In_313,In_304);
nand U1428 (N_1428,In_274,In_749);
nand U1429 (N_1429,In_573,In_939);
and U1430 (N_1430,In_330,In_440);
or U1431 (N_1431,In_58,In_870);
and U1432 (N_1432,In_384,In_6);
nor U1433 (N_1433,In_651,In_360);
nand U1434 (N_1434,In_511,In_426);
or U1435 (N_1435,In_81,In_880);
and U1436 (N_1436,In_494,In_934);
and U1437 (N_1437,In_593,In_719);
and U1438 (N_1438,In_701,In_981);
nor U1439 (N_1439,In_135,In_305);
or U1440 (N_1440,In_505,In_341);
and U1441 (N_1441,In_925,In_420);
and U1442 (N_1442,In_159,In_237);
or U1443 (N_1443,In_568,In_734);
or U1444 (N_1444,In_271,In_761);
nor U1445 (N_1445,In_879,In_459);
or U1446 (N_1446,In_95,In_661);
nor U1447 (N_1447,In_798,In_587);
and U1448 (N_1448,In_605,In_501);
nand U1449 (N_1449,In_628,In_383);
and U1450 (N_1450,In_152,In_649);
and U1451 (N_1451,In_778,In_272);
or U1452 (N_1452,In_283,In_963);
nor U1453 (N_1453,In_423,In_727);
nand U1454 (N_1454,In_212,In_271);
nand U1455 (N_1455,In_191,In_886);
nor U1456 (N_1456,In_624,In_325);
or U1457 (N_1457,In_644,In_698);
and U1458 (N_1458,In_182,In_838);
nand U1459 (N_1459,In_941,In_644);
and U1460 (N_1460,In_635,In_291);
nand U1461 (N_1461,In_804,In_426);
nand U1462 (N_1462,In_394,In_143);
nand U1463 (N_1463,In_442,In_367);
nand U1464 (N_1464,In_408,In_134);
nand U1465 (N_1465,In_780,In_657);
nand U1466 (N_1466,In_358,In_534);
and U1467 (N_1467,In_516,In_65);
or U1468 (N_1468,In_527,In_354);
nand U1469 (N_1469,In_578,In_694);
nand U1470 (N_1470,In_450,In_65);
nand U1471 (N_1471,In_924,In_135);
nand U1472 (N_1472,In_439,In_84);
nand U1473 (N_1473,In_224,In_228);
and U1474 (N_1474,In_926,In_421);
nand U1475 (N_1475,In_825,In_794);
nor U1476 (N_1476,In_981,In_955);
nor U1477 (N_1477,In_684,In_9);
and U1478 (N_1478,In_536,In_763);
and U1479 (N_1479,In_555,In_574);
nand U1480 (N_1480,In_573,In_596);
nor U1481 (N_1481,In_326,In_917);
or U1482 (N_1482,In_465,In_295);
or U1483 (N_1483,In_867,In_18);
nand U1484 (N_1484,In_78,In_491);
or U1485 (N_1485,In_245,In_959);
nor U1486 (N_1486,In_463,In_536);
nor U1487 (N_1487,In_302,In_710);
and U1488 (N_1488,In_731,In_231);
or U1489 (N_1489,In_609,In_590);
and U1490 (N_1490,In_769,In_944);
nand U1491 (N_1491,In_512,In_909);
nand U1492 (N_1492,In_907,In_735);
nor U1493 (N_1493,In_66,In_531);
or U1494 (N_1494,In_51,In_531);
and U1495 (N_1495,In_515,In_908);
nor U1496 (N_1496,In_279,In_862);
xor U1497 (N_1497,In_638,In_780);
and U1498 (N_1498,In_472,In_657);
nor U1499 (N_1499,In_570,In_677);
nand U1500 (N_1500,In_240,In_63);
nand U1501 (N_1501,In_688,In_201);
nand U1502 (N_1502,In_309,In_968);
or U1503 (N_1503,In_970,In_29);
nor U1504 (N_1504,In_101,In_963);
nand U1505 (N_1505,In_110,In_843);
and U1506 (N_1506,In_485,In_733);
and U1507 (N_1507,In_57,In_978);
or U1508 (N_1508,In_600,In_367);
and U1509 (N_1509,In_338,In_724);
or U1510 (N_1510,In_376,In_517);
nor U1511 (N_1511,In_158,In_387);
nand U1512 (N_1512,In_741,In_844);
or U1513 (N_1513,In_601,In_864);
nor U1514 (N_1514,In_732,In_683);
nor U1515 (N_1515,In_444,In_543);
nand U1516 (N_1516,In_989,In_27);
and U1517 (N_1517,In_983,In_549);
nor U1518 (N_1518,In_683,In_746);
or U1519 (N_1519,In_75,In_606);
nand U1520 (N_1520,In_327,In_59);
nand U1521 (N_1521,In_178,In_428);
or U1522 (N_1522,In_625,In_711);
nor U1523 (N_1523,In_982,In_774);
or U1524 (N_1524,In_925,In_196);
or U1525 (N_1525,In_703,In_499);
nor U1526 (N_1526,In_89,In_398);
nand U1527 (N_1527,In_738,In_511);
nor U1528 (N_1528,In_30,In_498);
nand U1529 (N_1529,In_759,In_401);
and U1530 (N_1530,In_496,In_933);
nor U1531 (N_1531,In_39,In_574);
nand U1532 (N_1532,In_252,In_425);
nor U1533 (N_1533,In_571,In_422);
nand U1534 (N_1534,In_105,In_665);
and U1535 (N_1535,In_210,In_839);
nand U1536 (N_1536,In_368,In_200);
nand U1537 (N_1537,In_904,In_600);
and U1538 (N_1538,In_987,In_828);
or U1539 (N_1539,In_952,In_68);
nand U1540 (N_1540,In_579,In_706);
and U1541 (N_1541,In_892,In_780);
and U1542 (N_1542,In_419,In_25);
nand U1543 (N_1543,In_61,In_557);
nor U1544 (N_1544,In_979,In_502);
and U1545 (N_1545,In_290,In_190);
and U1546 (N_1546,In_197,In_458);
nor U1547 (N_1547,In_623,In_597);
or U1548 (N_1548,In_31,In_409);
or U1549 (N_1549,In_224,In_410);
or U1550 (N_1550,In_751,In_869);
nand U1551 (N_1551,In_772,In_232);
nor U1552 (N_1552,In_120,In_642);
and U1553 (N_1553,In_234,In_506);
and U1554 (N_1554,In_227,In_245);
and U1555 (N_1555,In_411,In_209);
or U1556 (N_1556,In_80,In_557);
or U1557 (N_1557,In_766,In_852);
and U1558 (N_1558,In_648,In_758);
and U1559 (N_1559,In_389,In_33);
and U1560 (N_1560,In_120,In_134);
and U1561 (N_1561,In_500,In_516);
and U1562 (N_1562,In_92,In_266);
and U1563 (N_1563,In_955,In_932);
nor U1564 (N_1564,In_968,In_427);
and U1565 (N_1565,In_790,In_340);
nand U1566 (N_1566,In_251,In_80);
and U1567 (N_1567,In_992,In_391);
and U1568 (N_1568,In_681,In_577);
or U1569 (N_1569,In_367,In_965);
and U1570 (N_1570,In_590,In_124);
nor U1571 (N_1571,In_813,In_123);
and U1572 (N_1572,In_864,In_382);
or U1573 (N_1573,In_300,In_723);
nor U1574 (N_1574,In_142,In_668);
nor U1575 (N_1575,In_590,In_415);
nor U1576 (N_1576,In_780,In_208);
nand U1577 (N_1577,In_502,In_754);
or U1578 (N_1578,In_628,In_424);
or U1579 (N_1579,In_857,In_872);
and U1580 (N_1580,In_462,In_725);
nor U1581 (N_1581,In_910,In_239);
and U1582 (N_1582,In_637,In_244);
and U1583 (N_1583,In_63,In_387);
nand U1584 (N_1584,In_743,In_638);
and U1585 (N_1585,In_905,In_284);
or U1586 (N_1586,In_166,In_577);
and U1587 (N_1587,In_754,In_937);
nor U1588 (N_1588,In_967,In_573);
nor U1589 (N_1589,In_308,In_240);
and U1590 (N_1590,In_950,In_623);
nand U1591 (N_1591,In_926,In_590);
and U1592 (N_1592,In_121,In_542);
nor U1593 (N_1593,In_30,In_105);
nor U1594 (N_1594,In_467,In_669);
nor U1595 (N_1595,In_694,In_185);
or U1596 (N_1596,In_714,In_717);
nand U1597 (N_1597,In_567,In_731);
nor U1598 (N_1598,In_563,In_506);
or U1599 (N_1599,In_481,In_722);
nand U1600 (N_1600,In_317,In_665);
or U1601 (N_1601,In_379,In_686);
nand U1602 (N_1602,In_223,In_554);
nor U1603 (N_1603,In_842,In_812);
nor U1604 (N_1604,In_255,In_848);
and U1605 (N_1605,In_569,In_783);
nor U1606 (N_1606,In_155,In_318);
or U1607 (N_1607,In_161,In_154);
nor U1608 (N_1608,In_633,In_647);
nor U1609 (N_1609,In_535,In_795);
or U1610 (N_1610,In_335,In_226);
nor U1611 (N_1611,In_698,In_419);
nor U1612 (N_1612,In_259,In_119);
or U1613 (N_1613,In_633,In_990);
nor U1614 (N_1614,In_850,In_336);
nand U1615 (N_1615,In_418,In_621);
and U1616 (N_1616,In_71,In_525);
and U1617 (N_1617,In_408,In_820);
nor U1618 (N_1618,In_332,In_517);
nand U1619 (N_1619,In_809,In_323);
nor U1620 (N_1620,In_802,In_783);
nor U1621 (N_1621,In_641,In_14);
and U1622 (N_1622,In_848,In_329);
nor U1623 (N_1623,In_779,In_237);
or U1624 (N_1624,In_720,In_566);
nand U1625 (N_1625,In_786,In_232);
and U1626 (N_1626,In_873,In_958);
nor U1627 (N_1627,In_449,In_568);
or U1628 (N_1628,In_189,In_181);
or U1629 (N_1629,In_874,In_975);
nor U1630 (N_1630,In_413,In_514);
nor U1631 (N_1631,In_496,In_587);
or U1632 (N_1632,In_26,In_144);
nand U1633 (N_1633,In_996,In_528);
nand U1634 (N_1634,In_817,In_421);
nand U1635 (N_1635,In_979,In_207);
nand U1636 (N_1636,In_505,In_135);
nand U1637 (N_1637,In_28,In_634);
nor U1638 (N_1638,In_192,In_388);
nand U1639 (N_1639,In_602,In_436);
and U1640 (N_1640,In_265,In_770);
nor U1641 (N_1641,In_827,In_624);
and U1642 (N_1642,In_684,In_197);
nor U1643 (N_1643,In_208,In_677);
nand U1644 (N_1644,In_276,In_690);
nor U1645 (N_1645,In_812,In_473);
and U1646 (N_1646,In_616,In_928);
and U1647 (N_1647,In_678,In_375);
and U1648 (N_1648,In_531,In_915);
nand U1649 (N_1649,In_501,In_486);
and U1650 (N_1650,In_797,In_686);
nand U1651 (N_1651,In_279,In_514);
or U1652 (N_1652,In_527,In_734);
nand U1653 (N_1653,In_738,In_861);
and U1654 (N_1654,In_477,In_331);
or U1655 (N_1655,In_195,In_315);
and U1656 (N_1656,In_346,In_650);
nor U1657 (N_1657,In_314,In_313);
nand U1658 (N_1658,In_841,In_798);
and U1659 (N_1659,In_772,In_273);
or U1660 (N_1660,In_945,In_377);
nand U1661 (N_1661,In_398,In_383);
and U1662 (N_1662,In_894,In_506);
nor U1663 (N_1663,In_229,In_447);
nor U1664 (N_1664,In_9,In_931);
or U1665 (N_1665,In_902,In_750);
and U1666 (N_1666,In_789,In_751);
or U1667 (N_1667,In_474,In_348);
and U1668 (N_1668,In_742,In_777);
nand U1669 (N_1669,In_609,In_504);
nor U1670 (N_1670,In_116,In_576);
and U1671 (N_1671,In_955,In_924);
nor U1672 (N_1672,In_991,In_365);
nand U1673 (N_1673,In_379,In_64);
or U1674 (N_1674,In_732,In_823);
nand U1675 (N_1675,In_621,In_317);
or U1676 (N_1676,In_362,In_956);
and U1677 (N_1677,In_108,In_405);
nand U1678 (N_1678,In_585,In_217);
or U1679 (N_1679,In_255,In_605);
or U1680 (N_1680,In_366,In_288);
and U1681 (N_1681,In_181,In_626);
or U1682 (N_1682,In_704,In_117);
nor U1683 (N_1683,In_828,In_199);
nor U1684 (N_1684,In_72,In_570);
and U1685 (N_1685,In_170,In_562);
or U1686 (N_1686,In_829,In_662);
nor U1687 (N_1687,In_827,In_863);
nor U1688 (N_1688,In_708,In_673);
nand U1689 (N_1689,In_695,In_271);
nand U1690 (N_1690,In_938,In_216);
and U1691 (N_1691,In_182,In_467);
and U1692 (N_1692,In_626,In_970);
nand U1693 (N_1693,In_726,In_657);
nor U1694 (N_1694,In_646,In_850);
nor U1695 (N_1695,In_822,In_566);
and U1696 (N_1696,In_601,In_774);
nor U1697 (N_1697,In_619,In_346);
and U1698 (N_1698,In_412,In_561);
nor U1699 (N_1699,In_650,In_114);
nand U1700 (N_1700,In_680,In_768);
or U1701 (N_1701,In_952,In_976);
and U1702 (N_1702,In_876,In_17);
xor U1703 (N_1703,In_346,In_417);
nor U1704 (N_1704,In_950,In_501);
nand U1705 (N_1705,In_87,In_783);
nand U1706 (N_1706,In_52,In_257);
nand U1707 (N_1707,In_729,In_495);
nor U1708 (N_1708,In_990,In_926);
and U1709 (N_1709,In_768,In_256);
nor U1710 (N_1710,In_257,In_879);
nand U1711 (N_1711,In_464,In_235);
nor U1712 (N_1712,In_807,In_869);
nand U1713 (N_1713,In_569,In_888);
nand U1714 (N_1714,In_454,In_353);
nor U1715 (N_1715,In_644,In_522);
or U1716 (N_1716,In_578,In_810);
and U1717 (N_1717,In_28,In_82);
nand U1718 (N_1718,In_480,In_768);
and U1719 (N_1719,In_842,In_913);
nor U1720 (N_1720,In_590,In_605);
or U1721 (N_1721,In_492,In_312);
and U1722 (N_1722,In_88,In_787);
nand U1723 (N_1723,In_569,In_374);
nor U1724 (N_1724,In_745,In_443);
or U1725 (N_1725,In_190,In_792);
and U1726 (N_1726,In_704,In_607);
nor U1727 (N_1727,In_204,In_743);
or U1728 (N_1728,In_841,In_97);
or U1729 (N_1729,In_104,In_316);
nand U1730 (N_1730,In_57,In_489);
and U1731 (N_1731,In_563,In_838);
and U1732 (N_1732,In_662,In_424);
and U1733 (N_1733,In_828,In_482);
nand U1734 (N_1734,In_972,In_967);
nor U1735 (N_1735,In_972,In_334);
nor U1736 (N_1736,In_527,In_337);
nor U1737 (N_1737,In_905,In_393);
nand U1738 (N_1738,In_994,In_978);
and U1739 (N_1739,In_671,In_627);
or U1740 (N_1740,In_248,In_672);
nand U1741 (N_1741,In_113,In_458);
or U1742 (N_1742,In_680,In_557);
or U1743 (N_1743,In_781,In_38);
or U1744 (N_1744,In_541,In_503);
and U1745 (N_1745,In_85,In_727);
nand U1746 (N_1746,In_233,In_931);
or U1747 (N_1747,In_358,In_914);
nor U1748 (N_1748,In_515,In_512);
nor U1749 (N_1749,In_690,In_322);
and U1750 (N_1750,In_992,In_775);
nand U1751 (N_1751,In_99,In_150);
and U1752 (N_1752,In_706,In_721);
or U1753 (N_1753,In_443,In_208);
nand U1754 (N_1754,In_772,In_210);
nand U1755 (N_1755,In_973,In_138);
nand U1756 (N_1756,In_167,In_522);
nor U1757 (N_1757,In_595,In_816);
nor U1758 (N_1758,In_125,In_941);
nor U1759 (N_1759,In_114,In_521);
and U1760 (N_1760,In_229,In_296);
nand U1761 (N_1761,In_100,In_560);
or U1762 (N_1762,In_378,In_63);
nand U1763 (N_1763,In_410,In_453);
nor U1764 (N_1764,In_111,In_354);
xnor U1765 (N_1765,In_42,In_956);
nand U1766 (N_1766,In_799,In_216);
nor U1767 (N_1767,In_696,In_336);
nor U1768 (N_1768,In_554,In_587);
nor U1769 (N_1769,In_310,In_94);
or U1770 (N_1770,In_902,In_356);
nand U1771 (N_1771,In_17,In_977);
and U1772 (N_1772,In_449,In_494);
nand U1773 (N_1773,In_359,In_283);
nand U1774 (N_1774,In_455,In_383);
nor U1775 (N_1775,In_446,In_491);
nand U1776 (N_1776,In_381,In_520);
or U1777 (N_1777,In_919,In_958);
or U1778 (N_1778,In_999,In_572);
nor U1779 (N_1779,In_387,In_68);
and U1780 (N_1780,In_217,In_928);
nand U1781 (N_1781,In_304,In_5);
nand U1782 (N_1782,In_635,In_271);
or U1783 (N_1783,In_675,In_703);
and U1784 (N_1784,In_393,In_848);
nor U1785 (N_1785,In_300,In_154);
or U1786 (N_1786,In_458,In_784);
nor U1787 (N_1787,In_935,In_214);
or U1788 (N_1788,In_458,In_264);
nor U1789 (N_1789,In_750,In_383);
nor U1790 (N_1790,In_133,In_635);
nor U1791 (N_1791,In_555,In_100);
nor U1792 (N_1792,In_277,In_857);
and U1793 (N_1793,In_644,In_527);
and U1794 (N_1794,In_224,In_833);
and U1795 (N_1795,In_48,In_281);
and U1796 (N_1796,In_334,In_143);
or U1797 (N_1797,In_685,In_715);
nor U1798 (N_1798,In_403,In_30);
and U1799 (N_1799,In_505,In_645);
nor U1800 (N_1800,In_830,In_7);
nor U1801 (N_1801,In_85,In_730);
nor U1802 (N_1802,In_760,In_830);
nand U1803 (N_1803,In_227,In_554);
or U1804 (N_1804,In_386,In_873);
and U1805 (N_1805,In_369,In_324);
nor U1806 (N_1806,In_603,In_446);
and U1807 (N_1807,In_408,In_282);
nor U1808 (N_1808,In_691,In_579);
or U1809 (N_1809,In_832,In_791);
or U1810 (N_1810,In_219,In_513);
nand U1811 (N_1811,In_38,In_782);
or U1812 (N_1812,In_302,In_9);
nand U1813 (N_1813,In_906,In_822);
nand U1814 (N_1814,In_978,In_69);
nor U1815 (N_1815,In_685,In_2);
nand U1816 (N_1816,In_709,In_5);
or U1817 (N_1817,In_94,In_19);
nand U1818 (N_1818,In_480,In_29);
nand U1819 (N_1819,In_725,In_445);
nand U1820 (N_1820,In_925,In_282);
or U1821 (N_1821,In_532,In_302);
nand U1822 (N_1822,In_601,In_482);
nor U1823 (N_1823,In_63,In_93);
nor U1824 (N_1824,In_459,In_954);
nor U1825 (N_1825,In_412,In_866);
or U1826 (N_1826,In_78,In_878);
nor U1827 (N_1827,In_676,In_1);
nor U1828 (N_1828,In_884,In_975);
nor U1829 (N_1829,In_860,In_145);
or U1830 (N_1830,In_12,In_742);
and U1831 (N_1831,In_728,In_539);
or U1832 (N_1832,In_870,In_336);
nand U1833 (N_1833,In_636,In_292);
or U1834 (N_1834,In_952,In_688);
and U1835 (N_1835,In_501,In_767);
and U1836 (N_1836,In_717,In_819);
and U1837 (N_1837,In_671,In_176);
and U1838 (N_1838,In_922,In_386);
nor U1839 (N_1839,In_680,In_137);
or U1840 (N_1840,In_622,In_603);
nor U1841 (N_1841,In_88,In_946);
nor U1842 (N_1842,In_657,In_884);
and U1843 (N_1843,In_569,In_194);
and U1844 (N_1844,In_585,In_651);
nand U1845 (N_1845,In_883,In_214);
nor U1846 (N_1846,In_19,In_319);
and U1847 (N_1847,In_976,In_311);
or U1848 (N_1848,In_170,In_999);
or U1849 (N_1849,In_529,In_120);
nor U1850 (N_1850,In_757,In_313);
nand U1851 (N_1851,In_972,In_554);
nor U1852 (N_1852,In_799,In_453);
and U1853 (N_1853,In_721,In_321);
nor U1854 (N_1854,In_299,In_13);
and U1855 (N_1855,In_641,In_612);
and U1856 (N_1856,In_251,In_224);
nor U1857 (N_1857,In_161,In_882);
nand U1858 (N_1858,In_429,In_542);
or U1859 (N_1859,In_158,In_243);
nand U1860 (N_1860,In_427,In_99);
nand U1861 (N_1861,In_757,In_877);
and U1862 (N_1862,In_902,In_310);
nor U1863 (N_1863,In_643,In_932);
nor U1864 (N_1864,In_560,In_683);
or U1865 (N_1865,In_194,In_925);
nor U1866 (N_1866,In_479,In_20);
nor U1867 (N_1867,In_264,In_823);
nand U1868 (N_1868,In_581,In_299);
nand U1869 (N_1869,In_528,In_785);
and U1870 (N_1870,In_782,In_879);
xor U1871 (N_1871,In_703,In_709);
nor U1872 (N_1872,In_343,In_751);
nor U1873 (N_1873,In_857,In_98);
and U1874 (N_1874,In_804,In_964);
and U1875 (N_1875,In_43,In_674);
nand U1876 (N_1876,In_571,In_29);
and U1877 (N_1877,In_239,In_493);
nor U1878 (N_1878,In_622,In_664);
or U1879 (N_1879,In_460,In_387);
nor U1880 (N_1880,In_645,In_124);
nor U1881 (N_1881,In_465,In_306);
nor U1882 (N_1882,In_882,In_570);
nor U1883 (N_1883,In_893,In_476);
or U1884 (N_1884,In_373,In_44);
nor U1885 (N_1885,In_209,In_410);
nor U1886 (N_1886,In_396,In_653);
nor U1887 (N_1887,In_171,In_663);
nand U1888 (N_1888,In_444,In_701);
or U1889 (N_1889,In_596,In_993);
nand U1890 (N_1890,In_401,In_559);
and U1891 (N_1891,In_929,In_771);
nand U1892 (N_1892,In_98,In_442);
or U1893 (N_1893,In_772,In_50);
or U1894 (N_1894,In_749,In_688);
and U1895 (N_1895,In_32,In_199);
nor U1896 (N_1896,In_191,In_286);
or U1897 (N_1897,In_253,In_771);
nand U1898 (N_1898,In_916,In_672);
and U1899 (N_1899,In_444,In_889);
and U1900 (N_1900,In_556,In_663);
and U1901 (N_1901,In_678,In_179);
and U1902 (N_1902,In_372,In_724);
nand U1903 (N_1903,In_803,In_908);
xnor U1904 (N_1904,In_898,In_817);
nor U1905 (N_1905,In_906,In_807);
nor U1906 (N_1906,In_353,In_381);
nor U1907 (N_1907,In_100,In_183);
and U1908 (N_1908,In_690,In_679);
and U1909 (N_1909,In_910,In_612);
nor U1910 (N_1910,In_456,In_463);
and U1911 (N_1911,In_327,In_565);
xor U1912 (N_1912,In_679,In_627);
or U1913 (N_1913,In_795,In_111);
or U1914 (N_1914,In_152,In_513);
or U1915 (N_1915,In_107,In_19);
nor U1916 (N_1916,In_333,In_440);
and U1917 (N_1917,In_82,In_139);
xnor U1918 (N_1918,In_155,In_305);
nand U1919 (N_1919,In_798,In_125);
or U1920 (N_1920,In_267,In_615);
nand U1921 (N_1921,In_679,In_195);
nor U1922 (N_1922,In_804,In_510);
nor U1923 (N_1923,In_245,In_793);
and U1924 (N_1924,In_859,In_461);
and U1925 (N_1925,In_754,In_542);
nor U1926 (N_1926,In_292,In_665);
nand U1927 (N_1927,In_760,In_427);
nor U1928 (N_1928,In_702,In_903);
or U1929 (N_1929,In_692,In_94);
nor U1930 (N_1930,In_878,In_424);
nor U1931 (N_1931,In_730,In_347);
nand U1932 (N_1932,In_97,In_451);
nand U1933 (N_1933,In_393,In_868);
and U1934 (N_1934,In_254,In_528);
or U1935 (N_1935,In_940,In_420);
or U1936 (N_1936,In_242,In_588);
and U1937 (N_1937,In_908,In_958);
nand U1938 (N_1938,In_549,In_445);
nor U1939 (N_1939,In_466,In_45);
and U1940 (N_1940,In_749,In_634);
nand U1941 (N_1941,In_893,In_478);
nand U1942 (N_1942,In_335,In_182);
nor U1943 (N_1943,In_898,In_225);
nor U1944 (N_1944,In_89,In_714);
or U1945 (N_1945,In_825,In_214);
and U1946 (N_1946,In_151,In_557);
and U1947 (N_1947,In_938,In_843);
and U1948 (N_1948,In_999,In_849);
and U1949 (N_1949,In_191,In_173);
nor U1950 (N_1950,In_236,In_411);
xor U1951 (N_1951,In_66,In_589);
nor U1952 (N_1952,In_683,In_611);
or U1953 (N_1953,In_704,In_382);
nand U1954 (N_1954,In_115,In_35);
and U1955 (N_1955,In_573,In_222);
nand U1956 (N_1956,In_646,In_316);
or U1957 (N_1957,In_768,In_163);
nor U1958 (N_1958,In_160,In_887);
and U1959 (N_1959,In_737,In_408);
nand U1960 (N_1960,In_954,In_66);
nand U1961 (N_1961,In_709,In_25);
nand U1962 (N_1962,In_948,In_432);
nor U1963 (N_1963,In_705,In_744);
and U1964 (N_1964,In_868,In_1);
and U1965 (N_1965,In_719,In_987);
and U1966 (N_1966,In_528,In_35);
or U1967 (N_1967,In_896,In_221);
nor U1968 (N_1968,In_235,In_84);
nor U1969 (N_1969,In_426,In_412);
nand U1970 (N_1970,In_876,In_533);
and U1971 (N_1971,In_461,In_100);
or U1972 (N_1972,In_587,In_754);
or U1973 (N_1973,In_768,In_531);
nand U1974 (N_1974,In_574,In_883);
nor U1975 (N_1975,In_158,In_539);
or U1976 (N_1976,In_704,In_77);
or U1977 (N_1977,In_514,In_580);
or U1978 (N_1978,In_401,In_570);
and U1979 (N_1979,In_378,In_609);
nor U1980 (N_1980,In_932,In_515);
nor U1981 (N_1981,In_83,In_920);
or U1982 (N_1982,In_597,In_475);
nor U1983 (N_1983,In_463,In_338);
and U1984 (N_1984,In_140,In_122);
or U1985 (N_1985,In_788,In_283);
and U1986 (N_1986,In_16,In_665);
nor U1987 (N_1987,In_343,In_676);
or U1988 (N_1988,In_152,In_682);
and U1989 (N_1989,In_632,In_884);
or U1990 (N_1990,In_82,In_878);
nor U1991 (N_1991,In_110,In_71);
nand U1992 (N_1992,In_771,In_986);
nor U1993 (N_1993,In_58,In_234);
and U1994 (N_1994,In_719,In_262);
and U1995 (N_1995,In_851,In_602);
xnor U1996 (N_1996,In_878,In_804);
nand U1997 (N_1997,In_461,In_699);
or U1998 (N_1998,In_497,In_297);
nand U1999 (N_1999,In_987,In_806);
and U2000 (N_2000,N_1442,N_1709);
and U2001 (N_2001,N_1331,N_1135);
nand U2002 (N_2002,N_1077,N_464);
and U2003 (N_2003,N_923,N_1248);
and U2004 (N_2004,N_1382,N_1172);
or U2005 (N_2005,N_1512,N_782);
and U2006 (N_2006,N_1116,N_1040);
and U2007 (N_2007,N_264,N_569);
nor U2008 (N_2008,N_1106,N_1974);
nand U2009 (N_2009,N_114,N_600);
nor U2010 (N_2010,N_1858,N_292);
and U2011 (N_2011,N_1544,N_1255);
and U2012 (N_2012,N_127,N_1239);
and U2013 (N_2013,N_1816,N_1180);
nand U2014 (N_2014,N_1198,N_1062);
or U2015 (N_2015,N_479,N_1189);
and U2016 (N_2016,N_1938,N_481);
and U2017 (N_2017,N_1251,N_528);
and U2018 (N_2018,N_70,N_1081);
or U2019 (N_2019,N_410,N_1961);
and U2020 (N_2020,N_494,N_972);
nor U2021 (N_2021,N_1837,N_1827);
nand U2022 (N_2022,N_1394,N_201);
nor U2023 (N_2023,N_1607,N_1450);
or U2024 (N_2024,N_194,N_910);
and U2025 (N_2025,N_1810,N_1963);
or U2026 (N_2026,N_221,N_1949);
and U2027 (N_2027,N_297,N_1353);
nor U2028 (N_2028,N_1803,N_701);
nand U2029 (N_2029,N_1675,N_1917);
nor U2030 (N_2030,N_1128,N_1290);
or U2031 (N_2031,N_873,N_296);
nor U2032 (N_2032,N_807,N_1867);
nand U2033 (N_2033,N_273,N_882);
or U2034 (N_2034,N_710,N_780);
nand U2035 (N_2035,N_1279,N_324);
and U2036 (N_2036,N_1628,N_1638);
and U2037 (N_2037,N_497,N_151);
nor U2038 (N_2038,N_939,N_54);
nand U2039 (N_2039,N_203,N_1604);
and U2040 (N_2040,N_861,N_1433);
and U2041 (N_2041,N_963,N_593);
or U2042 (N_2042,N_738,N_805);
nand U2043 (N_2043,N_1818,N_1013);
nor U2044 (N_2044,N_330,N_1984);
xnor U2045 (N_2045,N_427,N_1975);
and U2046 (N_2046,N_523,N_1894);
nand U2047 (N_2047,N_1393,N_1035);
nand U2048 (N_2048,N_684,N_914);
and U2049 (N_2049,N_1031,N_912);
and U2050 (N_2050,N_709,N_862);
and U2051 (N_2051,N_1103,N_654);
nand U2052 (N_2052,N_35,N_1112);
and U2053 (N_2053,N_418,N_1388);
nor U2054 (N_2054,N_705,N_144);
and U2055 (N_2055,N_694,N_502);
nor U2056 (N_2056,N_988,N_1807);
or U2057 (N_2057,N_510,N_104);
or U2058 (N_2058,N_1943,N_1806);
or U2059 (N_2059,N_1569,N_350);
nand U2060 (N_2060,N_656,N_1434);
and U2061 (N_2061,N_1828,N_552);
nor U2062 (N_2062,N_214,N_1699);
and U2063 (N_2063,N_1733,N_567);
and U2064 (N_2064,N_348,N_171);
and U2065 (N_2065,N_1888,N_142);
nand U2066 (N_2066,N_145,N_1033);
or U2067 (N_2067,N_1101,N_1320);
nand U2068 (N_2068,N_1207,N_1413);
or U2069 (N_2069,N_1371,N_840);
or U2070 (N_2070,N_165,N_1579);
nand U2071 (N_2071,N_1585,N_565);
or U2072 (N_2072,N_764,N_1562);
nor U2073 (N_2073,N_985,N_1832);
nand U2074 (N_2074,N_1223,N_680);
and U2075 (N_2075,N_88,N_484);
nor U2076 (N_2076,N_859,N_1968);
nand U2077 (N_2077,N_1366,N_676);
nand U2078 (N_2078,N_1740,N_280);
xor U2079 (N_2079,N_531,N_997);
and U2080 (N_2080,N_1946,N_1854);
or U2081 (N_2081,N_474,N_1362);
and U2082 (N_2082,N_1278,N_785);
and U2083 (N_2083,N_1155,N_1613);
nand U2084 (N_2084,N_773,N_1276);
or U2085 (N_2085,N_1439,N_812);
and U2086 (N_2086,N_1504,N_1752);
and U2087 (N_2087,N_846,N_1408);
nor U2088 (N_2088,N_1289,N_1497);
and U2089 (N_2089,N_760,N_1325);
or U2090 (N_2090,N_1250,N_1783);
nor U2091 (N_2091,N_548,N_551);
or U2092 (N_2092,N_1852,N_642);
or U2093 (N_2093,N_1519,N_63);
and U2094 (N_2094,N_855,N_217);
nand U2095 (N_2095,N_1953,N_436);
and U2096 (N_2096,N_361,N_1932);
and U2097 (N_2097,N_1549,N_1652);
nor U2098 (N_2098,N_1058,N_626);
and U2099 (N_2099,N_1731,N_700);
or U2100 (N_2100,N_1057,N_1417);
or U2101 (N_2101,N_1340,N_1923);
and U2102 (N_2102,N_1677,N_331);
nand U2103 (N_2103,N_20,N_1778);
nand U2104 (N_2104,N_1650,N_1422);
nor U2105 (N_2105,N_1517,N_1684);
and U2106 (N_2106,N_1065,N_1564);
nor U2107 (N_2107,N_1884,N_1187);
or U2108 (N_2108,N_1751,N_1967);
nand U2109 (N_2109,N_532,N_1225);
and U2110 (N_2110,N_699,N_970);
nand U2111 (N_2111,N_645,N_1700);
and U2112 (N_2112,N_1485,N_1337);
nand U2113 (N_2113,N_390,N_668);
nand U2114 (N_2114,N_962,N_1855);
and U2115 (N_2115,N_1219,N_893);
xor U2116 (N_2116,N_170,N_1964);
nand U2117 (N_2117,N_45,N_400);
nor U2118 (N_2118,N_869,N_1666);
or U2119 (N_2119,N_1808,N_1727);
nor U2120 (N_2120,N_908,N_482);
or U2121 (N_2121,N_1174,N_1516);
nand U2122 (N_2122,N_850,N_17);
nor U2123 (N_2123,N_1679,N_1142);
and U2124 (N_2124,N_453,N_944);
and U2125 (N_2125,N_1299,N_1499);
nor U2126 (N_2126,N_34,N_877);
nand U2127 (N_2127,N_1070,N_1994);
or U2128 (N_2128,N_1351,N_1835);
or U2129 (N_2129,N_200,N_284);
nand U2130 (N_2130,N_1614,N_679);
and U2131 (N_2131,N_1910,N_1794);
nor U2132 (N_2132,N_1238,N_996);
or U2133 (N_2133,N_1271,N_779);
nand U2134 (N_2134,N_1472,N_362);
or U2135 (N_2135,N_105,N_247);
or U2136 (N_2136,N_1399,N_745);
nor U2137 (N_2137,N_409,N_211);
or U2138 (N_2138,N_1181,N_1334);
or U2139 (N_2139,N_351,N_352);
and U2140 (N_2140,N_298,N_713);
and U2141 (N_2141,N_1507,N_1635);
and U2142 (N_2142,N_1527,N_1498);
xnor U2143 (N_2143,N_951,N_43);
or U2144 (N_2144,N_176,N_309);
and U2145 (N_2145,N_977,N_1011);
or U2146 (N_2146,N_627,N_279);
and U2147 (N_2147,N_1988,N_108);
and U2148 (N_2148,N_225,N_1830);
and U2149 (N_2149,N_1339,N_466);
nand U2150 (N_2150,N_1034,N_371);
nor U2151 (N_2151,N_1622,N_1547);
and U2152 (N_2152,N_1895,N_377);
nor U2153 (N_2153,N_72,N_156);
nand U2154 (N_2154,N_432,N_1158);
nor U2155 (N_2155,N_29,N_1697);
and U2156 (N_2156,N_174,N_771);
and U2157 (N_2157,N_911,N_1078);
or U2158 (N_2158,N_1269,N_78);
nand U2159 (N_2159,N_1678,N_570);
nand U2160 (N_2160,N_438,N_1490);
nor U2161 (N_2161,N_1649,N_1283);
nand U2162 (N_2162,N_1372,N_1762);
or U2163 (N_2163,N_1117,N_1669);
and U2164 (N_2164,N_1049,N_276);
or U2165 (N_2165,N_1188,N_1476);
nand U2166 (N_2166,N_1360,N_451);
nand U2167 (N_2167,N_653,N_533);
or U2168 (N_2168,N_1014,N_802);
and U2169 (N_2169,N_1051,N_1822);
nand U2170 (N_2170,N_832,N_1235);
or U2171 (N_2171,N_596,N_1277);
xnor U2172 (N_2172,N_1061,N_1589);
nand U2173 (N_2173,N_1068,N_966);
and U2174 (N_2174,N_845,N_353);
or U2175 (N_2175,N_1798,N_1716);
nor U2176 (N_2176,N_793,N_1495);
nor U2177 (N_2177,N_719,N_1267);
or U2178 (N_2178,N_887,N_1839);
nand U2179 (N_2179,N_1621,N_393);
nand U2180 (N_2180,N_55,N_1880);
nor U2181 (N_2181,N_714,N_277);
nand U2182 (N_2182,N_1991,N_1411);
nor U2183 (N_2183,N_928,N_506);
and U2184 (N_2184,N_1484,N_711);
or U2185 (N_2185,N_1183,N_1119);
and U2186 (N_2186,N_1004,N_218);
nor U2187 (N_2187,N_1471,N_159);
nand U2188 (N_2188,N_1902,N_148);
nand U2189 (N_2189,N_1573,N_942);
nand U2190 (N_2190,N_1330,N_818);
and U2191 (N_2191,N_237,N_73);
nor U2192 (N_2192,N_1319,N_830);
nand U2193 (N_2193,N_918,N_1620);
or U2194 (N_2194,N_266,N_15);
and U2195 (N_2195,N_447,N_109);
nand U2196 (N_2196,N_1899,N_103);
or U2197 (N_2197,N_251,N_204);
and U2198 (N_2198,N_1987,N_139);
nand U2199 (N_2199,N_872,N_1924);
nor U2200 (N_2200,N_1287,N_106);
or U2201 (N_2201,N_538,N_121);
nor U2202 (N_2202,N_1210,N_1378);
or U2203 (N_2203,N_1651,N_1390);
nor U2204 (N_2204,N_1170,N_575);
or U2205 (N_2205,N_4,N_450);
and U2206 (N_2206,N_1344,N_1936);
nor U2207 (N_2207,N_1097,N_1066);
and U2208 (N_2208,N_930,N_367);
nor U2209 (N_2209,N_913,N_1550);
nand U2210 (N_2210,N_856,N_530);
or U2211 (N_2211,N_265,N_857);
and U2212 (N_2212,N_511,N_534);
and U2213 (N_2213,N_1275,N_245);
nand U2214 (N_2214,N_235,N_1797);
and U2215 (N_2215,N_490,N_295);
and U2216 (N_2216,N_617,N_876);
or U2217 (N_2217,N_1745,N_226);
or U2218 (N_2218,N_1653,N_1313);
nor U2219 (N_2219,N_308,N_1851);
nand U2220 (N_2220,N_820,N_1515);
nand U2221 (N_2221,N_1788,N_469);
nor U2222 (N_2222,N_1195,N_1947);
nor U2223 (N_2223,N_1201,N_1298);
or U2224 (N_2224,N_1680,N_412);
nand U2225 (N_2225,N_1771,N_195);
and U2226 (N_2226,N_925,N_734);
or U2227 (N_2227,N_1359,N_1217);
and U2228 (N_2228,N_1608,N_1701);
nor U2229 (N_2229,N_249,N_1506);
nand U2230 (N_2230,N_448,N_852);
nor U2231 (N_2231,N_1431,N_491);
or U2232 (N_2232,N_116,N_622);
or U2233 (N_2233,N_1599,N_1995);
nand U2234 (N_2234,N_1916,N_314);
and U2235 (N_2235,N_1615,N_118);
or U2236 (N_2236,N_1829,N_1776);
nand U2237 (N_2237,N_422,N_563);
or U2238 (N_2238,N_141,N_936);
or U2239 (N_2239,N_1721,N_1148);
and U2240 (N_2240,N_580,N_0);
and U2241 (N_2241,N_1875,N_1941);
nor U2242 (N_2242,N_99,N_463);
and U2243 (N_2243,N_1163,N_496);
or U2244 (N_2244,N_13,N_46);
nand U2245 (N_2245,N_1132,N_1426);
and U2246 (N_2246,N_662,N_87);
xnor U2247 (N_2247,N_166,N_1878);
or U2248 (N_2248,N_863,N_1202);
nor U2249 (N_2249,N_1427,N_744);
nand U2250 (N_2250,N_1996,N_489);
and U2251 (N_2251,N_3,N_136);
and U2252 (N_2252,N_1374,N_1000);
nand U2253 (N_2253,N_205,N_442);
and U2254 (N_2254,N_1083,N_1118);
and U2255 (N_2255,N_1882,N_1139);
nor U2256 (N_2256,N_1841,N_1557);
nand U2257 (N_2257,N_1111,N_1877);
or U2258 (N_2258,N_1715,N_1896);
nor U2259 (N_2259,N_1785,N_1959);
or U2260 (N_2260,N_1594,N_1780);
nand U2261 (N_2261,N_1322,N_761);
nand U2262 (N_2262,N_210,N_815);
nand U2263 (N_2263,N_839,N_1800);
and U2264 (N_2264,N_8,N_774);
or U2265 (N_2265,N_597,N_664);
and U2266 (N_2266,N_1206,N_843);
or U2267 (N_2267,N_206,N_844);
and U2268 (N_2268,N_1312,N_186);
and U2269 (N_2269,N_378,N_998);
nor U2270 (N_2270,N_1392,N_290);
and U2271 (N_2271,N_824,N_1746);
nand U2272 (N_2272,N_1747,N_767);
nor U2273 (N_2273,N_509,N_437);
and U2274 (N_2274,N_1933,N_1587);
nand U2275 (N_2275,N_1496,N_1503);
nand U2276 (N_2276,N_1843,N_598);
and U2277 (N_2277,N_1718,N_544);
nand U2278 (N_2278,N_665,N_1449);
and U2279 (N_2279,N_1345,N_310);
or U2280 (N_2280,N_1976,N_59);
nor U2281 (N_2281,N_1094,N_742);
and U2282 (N_2282,N_1805,N_1026);
nor U2283 (N_2283,N_1140,N_620);
and U2284 (N_2284,N_1518,N_1897);
nand U2285 (N_2285,N_178,N_746);
nor U2286 (N_2286,N_1326,N_1826);
nor U2287 (N_2287,N_443,N_1335);
and U2288 (N_2288,N_1510,N_588);
and U2289 (N_2289,N_1212,N_380);
and U2290 (N_2290,N_1368,N_585);
and U2291 (N_2291,N_1153,N_1689);
nor U2292 (N_2292,N_1059,N_161);
and U2293 (N_2293,N_1912,N_633);
nand U2294 (N_2294,N_1908,N_130);
nand U2295 (N_2295,N_1999,N_1811);
nand U2296 (N_2296,N_1759,N_888);
or U2297 (N_2297,N_1577,N_94);
nor U2298 (N_2298,N_135,N_456);
nand U2299 (N_2299,N_1421,N_1921);
and U2300 (N_2300,N_1205,N_715);
nor U2301 (N_2301,N_404,N_1071);
or U2302 (N_2302,N_1537,N_1245);
and U2303 (N_2303,N_1475,N_690);
nand U2304 (N_2304,N_49,N_1981);
nor U2305 (N_2305,N_119,N_301);
or U2306 (N_2306,N_1461,N_1447);
nor U2307 (N_2307,N_1539,N_553);
or U2308 (N_2308,N_1892,N_65);
nor U2309 (N_2309,N_560,N_1571);
and U2310 (N_2310,N_623,N_6);
nor U2311 (N_2311,N_1177,N_982);
xor U2312 (N_2312,N_838,N_1010);
nor U2313 (N_2313,N_1859,N_1487);
nor U2314 (N_2314,N_638,N_955);
nand U2315 (N_2315,N_1384,N_1674);
nor U2316 (N_2316,N_909,N_1869);
and U2317 (N_2317,N_1470,N_1024);
nand U2318 (N_2318,N_1664,N_747);
and U2319 (N_2319,N_1355,N_1179);
nand U2320 (N_2320,N_1559,N_1823);
nor U2321 (N_2321,N_1074,N_1324);
and U2322 (N_2322,N_1758,N_117);
and U2323 (N_2323,N_224,N_1333);
xnor U2324 (N_2324,N_1847,N_834);
and U2325 (N_2325,N_306,N_1619);
nor U2326 (N_2326,N_399,N_707);
and U2327 (N_2327,N_1753,N_646);
and U2328 (N_2328,N_1021,N_1416);
nand U2329 (N_2329,N_776,N_234);
nor U2330 (N_2330,N_1088,N_967);
xnor U2331 (N_2331,N_101,N_1568);
nor U2332 (N_2332,N_935,N_722);
or U2333 (N_2333,N_907,N_986);
nand U2334 (N_2334,N_1911,N_125);
or U2335 (N_2335,N_637,N_529);
and U2336 (N_2336,N_1790,N_1872);
nand U2337 (N_2337,N_1369,N_37);
nand U2338 (N_2338,N_1171,N_1317);
nand U2339 (N_2339,N_299,N_193);
and U2340 (N_2340,N_402,N_1246);
or U2341 (N_2341,N_1046,N_1134);
and U2342 (N_2342,N_2,N_107);
nand U2343 (N_2343,N_1428,N_883);
nor U2344 (N_2344,N_1970,N_431);
nor U2345 (N_2345,N_659,N_56);
nand U2346 (N_2346,N_480,N_196);
or U2347 (N_2347,N_591,N_1723);
or U2348 (N_2348,N_487,N_697);
nand U2349 (N_2349,N_870,N_708);
or U2350 (N_2350,N_1636,N_1098);
nand U2351 (N_2351,N_1376,N_1280);
nand U2352 (N_2352,N_572,N_991);
nor U2353 (N_2353,N_1136,N_613);
nand U2354 (N_2354,N_1572,N_546);
and U2355 (N_2355,N_554,N_571);
nor U2356 (N_2356,N_1842,N_387);
and U2357 (N_2357,N_1072,N_667);
nand U2358 (N_2358,N_149,N_1231);
and U2359 (N_2359,N_1809,N_1091);
nand U2360 (N_2360,N_547,N_688);
nor U2361 (N_2361,N_1184,N_1030);
and U2362 (N_2362,N_5,N_836);
nor U2363 (N_2363,N_1131,N_516);
nand U2364 (N_2364,N_163,N_1402);
nor U2365 (N_2365,N_550,N_1696);
nand U2366 (N_2366,N_905,N_407);
or U2367 (N_2367,N_961,N_1993);
xor U2368 (N_2368,N_758,N_169);
nand U2369 (N_2369,N_1474,N_1348);
nor U2370 (N_2370,N_1467,N_1926);
nor U2371 (N_2371,N_270,N_1303);
or U2372 (N_2372,N_147,N_64);
or U2373 (N_2373,N_369,N_1272);
or U2374 (N_2374,N_1092,N_1063);
nor U2375 (N_2375,N_1942,N_1533);
nand U2376 (N_2376,N_449,N_250);
and U2377 (N_2377,N_85,N_1254);
or U2378 (N_2378,N_246,N_175);
nor U2379 (N_2379,N_655,N_599);
and U2380 (N_2380,N_1919,N_96);
and U2381 (N_2381,N_1554,N_1200);
or U2382 (N_2382,N_417,N_634);
nand U2383 (N_2383,N_1270,N_32);
and U2384 (N_2384,N_240,N_590);
nor U2385 (N_2385,N_712,N_987);
and U2386 (N_2386,N_415,N_1769);
or U2387 (N_2387,N_1266,N_1138);
and U2388 (N_2388,N_720,N_1149);
or U2389 (N_2389,N_1575,N_629);
or U2390 (N_2390,N_1463,N_248);
and U2391 (N_2391,N_1354,N_207);
or U2392 (N_2392,N_1958,N_275);
or U2393 (N_2393,N_304,N_1401);
or U2394 (N_2394,N_359,N_1927);
and U2395 (N_2395,N_1609,N_440);
and U2396 (N_2396,N_1242,N_446);
and U2397 (N_2397,N_1720,N_1704);
nand U2398 (N_2398,N_770,N_691);
and U2399 (N_2399,N_1658,N_80);
nor U2400 (N_2400,N_355,N_1125);
and U2401 (N_2401,N_1403,N_537);
nand U2402 (N_2402,N_258,N_1089);
or U2403 (N_2403,N_558,N_215);
nand U2404 (N_2404,N_202,N_26);
and U2405 (N_2405,N_79,N_1584);
and U2406 (N_2406,N_1915,N_917);
nor U2407 (N_2407,N_527,N_1479);
and U2408 (N_2408,N_1015,N_1361);
or U2409 (N_2409,N_1123,N_1222);
nor U2410 (N_2410,N_1883,N_1944);
and U2411 (N_2411,N_1777,N_1813);
nand U2412 (N_2412,N_357,N_1860);
and U2413 (N_2413,N_1918,N_1237);
nand U2414 (N_2414,N_227,N_229);
nor U2415 (N_2415,N_381,N_1310);
or U2416 (N_2416,N_1914,N_1044);
nand U2417 (N_2417,N_1432,N_1095);
nor U2418 (N_2418,N_871,N_894);
nand U2419 (N_2419,N_503,N_1849);
and U2420 (N_2420,N_1193,N_1338);
or U2421 (N_2421,N_926,N_1726);
or U2422 (N_2422,N_1151,N_1157);
nor U2423 (N_2423,N_549,N_334);
nor U2424 (N_2424,N_1781,N_505);
nor U2425 (N_2425,N_1526,N_733);
or U2426 (N_2426,N_233,N_583);
nand U2427 (N_2427,N_1692,N_254);
or U2428 (N_2428,N_256,N_189);
nor U2429 (N_2429,N_1052,N_837);
nor U2430 (N_2430,N_1380,N_1815);
nor U2431 (N_2431,N_1349,N_1948);
nand U2432 (N_2432,N_1284,N_1352);
or U2433 (N_2433,N_687,N_467);
nand U2434 (N_2434,N_1901,N_616);
and U2435 (N_2435,N_1363,N_1913);
nand U2436 (N_2436,N_1309,N_740);
or U2437 (N_2437,N_1711,N_1850);
nand U2438 (N_2438,N_1076,N_1191);
nor U2439 (N_2439,N_1130,N_1006);
or U2440 (N_2440,N_97,N_1165);
and U2441 (N_2441,N_157,N_1846);
and U2442 (N_2442,N_133,N_1682);
nand U2443 (N_2443,N_1929,N_423);
or U2444 (N_2444,N_154,N_472);
and U2445 (N_2445,N_398,N_851);
and U2446 (N_2446,N_1249,N_609);
nand U2447 (N_2447,N_1121,N_841);
and U2448 (N_2448,N_1623,N_822);
nand U2449 (N_2449,N_1318,N_1705);
and U2450 (N_2450,N_230,N_1928);
or U2451 (N_2451,N_1258,N_1304);
nand U2452 (N_2452,N_929,N_848);
and U2453 (N_2453,N_92,N_539);
or U2454 (N_2454,N_1655,N_606);
and U2455 (N_2455,N_1950,N_1323);
nand U2456 (N_2456,N_631,N_1952);
and U2457 (N_2457,N_1764,N_397);
nand U2458 (N_2458,N_1446,N_396);
or U2459 (N_2459,N_1531,N_1002);
and U2460 (N_2460,N_829,N_1488);
nand U2461 (N_2461,N_500,N_1306);
or U2462 (N_2462,N_754,N_1377);
nand U2463 (N_2463,N_460,N_1538);
nand U2464 (N_2464,N_1291,N_51);
nand U2465 (N_2465,N_1164,N_833);
nand U2466 (N_2466,N_1032,N_792);
and U2467 (N_2467,N_342,N_74);
nor U2468 (N_2468,N_242,N_1316);
or U2469 (N_2469,N_1395,N_328);
or U2470 (N_2470,N_168,N_1028);
nand U2471 (N_2471,N_683,N_1586);
nor U2472 (N_2472,N_405,N_1185);
or U2473 (N_2473,N_7,N_641);
and U2474 (N_2474,N_1668,N_896);
nor U2475 (N_2475,N_1418,N_769);
nor U2476 (N_2476,N_1937,N_408);
nand U2477 (N_2477,N_1690,N_316);
or U2478 (N_2478,N_1553,N_1603);
nor U2479 (N_2479,N_1373,N_1717);
and U2480 (N_2480,N_766,N_21);
and U2481 (N_2481,N_678,N_777);
or U2482 (N_2482,N_1243,N_568);
and U2483 (N_2483,N_394,N_1760);
and U2484 (N_2484,N_180,N_373);
nand U2485 (N_2485,N_974,N_134);
and U2486 (N_2486,N_756,N_957);
or U2487 (N_2487,N_1529,N_1514);
nand U2488 (N_2488,N_1473,N_1260);
or U2489 (N_2489,N_1702,N_18);
nand U2490 (N_2490,N_753,N_724);
or U2491 (N_2491,N_1775,N_809);
and U2492 (N_2492,N_799,N_625);
nand U2493 (N_2493,N_1945,N_302);
nor U2494 (N_2494,N_1631,N_1425);
and U2495 (N_2495,N_1989,N_1025);
or U2496 (N_2496,N_473,N_260);
or U2497 (N_2497,N_263,N_1169);
nand U2498 (N_2498,N_1451,N_152);
or U2499 (N_2499,N_1956,N_1090);
nor U2500 (N_2500,N_90,N_383);
nand U2501 (N_2501,N_765,N_1966);
nand U2502 (N_2502,N_735,N_1863);
or U2503 (N_2503,N_1367,N_971);
nand U2504 (N_2504,N_1898,N_915);
nand U2505 (N_2505,N_1660,N_340);
nand U2506 (N_2506,N_1465,N_884);
and U2507 (N_2507,N_1645,N_471);
nor U2508 (N_2508,N_198,N_1285);
or U2509 (N_2509,N_60,N_1152);
nor U2510 (N_2510,N_1167,N_749);
or U2511 (N_2511,N_727,N_1814);
nand U2512 (N_2512,N_1096,N_1890);
nand U2513 (N_2513,N_1166,N_999);
nor U2514 (N_2514,N_732,N_689);
nand U2515 (N_2515,N_864,N_470);
or U2516 (N_2516,N_1998,N_375);
and U2517 (N_2517,N_1227,N_847);
and U2518 (N_2518,N_1412,N_1199);
nand U2519 (N_2519,N_1983,N_1505);
nor U2520 (N_2520,N_475,N_1694);
and U2521 (N_2521,N_736,N_1556);
and U2522 (N_2522,N_1834,N_311);
nand U2523 (N_2523,N_608,N_752);
nand U2524 (N_2524,N_1922,N_1224);
nor U2525 (N_2525,N_934,N_1560);
nand U2526 (N_2526,N_1532,N_695);
or U2527 (N_2527,N_236,N_126);
and U2528 (N_2528,N_1687,N_445);
or U2529 (N_2529,N_1329,N_1821);
nor U2530 (N_2530,N_269,N_858);
nor U2531 (N_2531,N_1824,N_1646);
and U2532 (N_2532,N_685,N_1561);
and U2533 (N_2533,N_1468,N_160);
or U2534 (N_2534,N_1307,N_1295);
nor U2535 (N_2535,N_1060,N_522);
and U2536 (N_2536,N_1146,N_696);
or U2537 (N_2537,N_89,N_179);
or U2538 (N_2538,N_562,N_1410);
nor U2539 (N_2539,N_1124,N_1602);
and U2540 (N_2540,N_938,N_521);
and U2541 (N_2541,N_525,N_555);
and U2542 (N_2542,N_1161,N_19);
nor U2543 (N_2543,N_115,N_958);
and U2544 (N_2544,N_384,N_557);
and U2545 (N_2545,N_1729,N_1612);
or U2546 (N_2546,N_755,N_177);
nor U2547 (N_2547,N_388,N_1292);
nand U2548 (N_2548,N_1749,N_1773);
and U2549 (N_2549,N_1486,N_584);
or U2550 (N_2550,N_1494,N_1197);
nor U2551 (N_2551,N_1887,N_1424);
and U2552 (N_2552,N_759,N_932);
and U2553 (N_2553,N_183,N_1302);
or U2554 (N_2554,N_878,N_1951);
nand U2555 (N_2555,N_979,N_1383);
nand U2556 (N_2556,N_940,N_77);
nand U2557 (N_2557,N_1574,N_1301);
or U2558 (N_2558,N_48,N_27);
nand U2559 (N_2559,N_541,N_797);
nor U2560 (N_2560,N_559,N_1228);
nand U2561 (N_2561,N_1196,N_831);
or U2562 (N_2562,N_167,N_804);
or U2563 (N_2563,N_1480,N_1005);
nand U2564 (N_2564,N_1583,N_675);
and U2565 (N_2565,N_389,N_75);
nor U2566 (N_2566,N_1750,N_698);
or U2567 (N_2567,N_1105,N_1840);
nor U2568 (N_2568,N_1102,N_564);
nand U2569 (N_2569,N_671,N_1268);
and U2570 (N_2570,N_919,N_478);
and U2571 (N_2571,N_382,N_1904);
nand U2572 (N_2572,N_1257,N_1300);
nand U2573 (N_2573,N_1216,N_1535);
nor U2574 (N_2574,N_138,N_1685);
nor U2575 (N_2575,N_1168,N_798);
and U2576 (N_2576,N_842,N_155);
or U2577 (N_2577,N_916,N_716);
nor U2578 (N_2578,N_775,N_1232);
or U2579 (N_2579,N_976,N_341);
nor U2580 (N_2580,N_1695,N_1017);
nor U2581 (N_2581,N_561,N_1763);
nor U2582 (N_2582,N_1159,N_370);
nor U2583 (N_2583,N_83,N_86);
nor U2584 (N_2584,N_731,N_31);
nand U2585 (N_2585,N_636,N_1430);
nand U2586 (N_2586,N_1833,N_651);
nor U2587 (N_2587,N_321,N_499);
nor U2588 (N_2588,N_100,N_223);
nor U2589 (N_2589,N_57,N_262);
nand U2590 (N_2590,N_1606,N_1703);
nor U2591 (N_2591,N_674,N_945);
nor U2592 (N_2592,N_1099,N_704);
nand U2593 (N_2593,N_1812,N_50);
nor U2594 (N_2594,N_823,N_455);
or U2595 (N_2595,N_1252,N_730);
nand U2596 (N_2596,N_498,N_640);
nand U2597 (N_2597,N_162,N_128);
and U2598 (N_2598,N_1862,N_781);
and U2599 (N_2599,N_1903,N_372);
nor U2600 (N_2600,N_890,N_123);
nand U2601 (N_2601,N_140,N_1047);
nand U2602 (N_2602,N_1647,N_868);
nor U2603 (N_2603,N_946,N_1525);
nor U2604 (N_2604,N_1969,N_1761);
or U2605 (N_2605,N_212,N_826);
nand U2606 (N_2606,N_150,N_1802);
or U2607 (N_2607,N_1209,N_1540);
nand U2608 (N_2608,N_430,N_421);
and U2609 (N_2609,N_1971,N_1502);
or U2610 (N_2610,N_1454,N_615);
or U2611 (N_2611,N_1286,N_191);
and U2612 (N_2612,N_1972,N_403);
nand U2613 (N_2613,N_1893,N_866);
or U2614 (N_2614,N_1419,N_1436);
nand U2615 (N_2615,N_990,N_1524);
and U2616 (N_2616,N_1263,N_1667);
and U2617 (N_2617,N_604,N_1445);
and U2618 (N_2618,N_1229,N_1194);
or U2619 (N_2619,N_542,N_337);
nor U2620 (N_2620,N_1457,N_197);
nor U2621 (N_2621,N_1548,N_1511);
or U2622 (N_2622,N_1160,N_1713);
nand U2623 (N_2623,N_725,N_433);
nand U2624 (N_2624,N_1043,N_1768);
nand U2625 (N_2625,N_1234,N_347);
nand U2626 (N_2626,N_892,N_1455);
nor U2627 (N_2627,N_1069,N_42);
nor U2628 (N_2628,N_1203,N_810);
nand U2629 (N_2629,N_978,N_1154);
nor U2630 (N_2630,N_146,N_723);
nand U2631 (N_2631,N_1444,N_1874);
nor U2632 (N_2632,N_1437,N_1293);
nor U2633 (N_2633,N_1641,N_587);
or U2634 (N_2634,N_803,N_1848);
nand U2635 (N_2635,N_898,N_743);
nor U2636 (N_2636,N_1520,N_1233);
and U2637 (N_2637,N_922,N_791);
nand U2638 (N_2638,N_1240,N_1336);
or U2639 (N_2639,N_786,N_426);
nand U2640 (N_2640,N_989,N_401);
or U2641 (N_2641,N_392,N_835);
or U2642 (N_2642,N_307,N_458);
nand U2643 (N_2643,N_454,N_1960);
or U2644 (N_2644,N_1350,N_1523);
nor U2645 (N_2645,N_1779,N_58);
nand U2646 (N_2646,N_1477,N_1670);
and U2647 (N_2647,N_1459,N_995);
and U2648 (N_2648,N_853,N_1870);
nor U2649 (N_2649,N_1605,N_1642);
or U2650 (N_2650,N_1466,N_241);
nor U2651 (N_2651,N_1029,N_483);
nor U2652 (N_2652,N_1007,N_1321);
and U2653 (N_2653,N_1672,N_1909);
nor U2654 (N_2654,N_827,N_1086);
or U2655 (N_2655,N_949,N_875);
nand U2656 (N_2656,N_783,N_1930);
or U2657 (N_2657,N_1691,N_435);
or U2658 (N_2658,N_1037,N_1055);
or U2659 (N_2659,N_1085,N_574);
or U2660 (N_2660,N_333,N_1469);
nor U2661 (N_2661,N_1920,N_952);
and U2662 (N_2662,N_1400,N_1997);
nand U2663 (N_2663,N_452,N_1534);
nor U2664 (N_2664,N_158,N_1087);
nand U2665 (N_2665,N_461,N_1150);
nor U2666 (N_2666,N_1110,N_44);
or U2667 (N_2667,N_1581,N_881);
or U2668 (N_2668,N_1178,N_1555);
or U2669 (N_2669,N_411,N_28);
nand U2670 (N_2670,N_1838,N_1627);
and U2671 (N_2671,N_293,N_1084);
nand U2672 (N_2672,N_578,N_906);
nor U2673 (N_2673,N_789,N_1656);
nor U2674 (N_2674,N_573,N_338);
nand U2675 (N_2675,N_524,N_232);
and U2676 (N_2676,N_1708,N_886);
nand U2677 (N_2677,N_1483,N_25);
or U2678 (N_2678,N_501,N_1772);
and U2679 (N_2679,N_885,N_504);
and U2680 (N_2680,N_122,N_305);
and U2681 (N_2681,N_1415,N_1563);
or U2682 (N_2682,N_1643,N_1873);
or U2683 (N_2683,N_648,N_428);
and U2684 (N_2684,N_579,N_1597);
nand U2685 (N_2685,N_1804,N_1662);
and U2686 (N_2686,N_414,N_239);
nand U2687 (N_2687,N_1173,N_343);
or U2688 (N_2688,N_1443,N_84);
and U2689 (N_2689,N_540,N_520);
nor U2690 (N_2690,N_874,N_1601);
and U2691 (N_2691,N_1681,N_1879);
nand U2692 (N_2692,N_602,N_751);
or U2693 (N_2693,N_209,N_1104);
or U2694 (N_2694,N_1965,N_1985);
nand U2695 (N_2695,N_768,N_1625);
or U2696 (N_2696,N_1792,N_953);
nor U2697 (N_2697,N_1143,N_1332);
nand U2698 (N_2698,N_1748,N_1346);
and U2699 (N_2699,N_1856,N_1365);
nand U2700 (N_2700,N_317,N_1441);
nand U2701 (N_2701,N_112,N_1513);
and U2702 (N_2702,N_1221,N_950);
nand U2703 (N_2703,N_1639,N_983);
or U2704 (N_2704,N_319,N_897);
xor U2705 (N_2705,N_322,N_181);
or U2706 (N_2706,N_252,N_52);
nand U2707 (N_2707,N_1939,N_790);
nand U2708 (N_2708,N_728,N_1676);
or U2709 (N_2709,N_1082,N_1825);
or U2710 (N_2710,N_1012,N_30);
nand U2711 (N_2711,N_69,N_335);
or U2712 (N_2712,N_1844,N_339);
nand U2713 (N_2713,N_536,N_652);
and U2714 (N_2714,N_1464,N_1986);
or U2715 (N_2715,N_649,N_1688);
and U2716 (N_2716,N_1698,N_1114);
nor U2717 (N_2717,N_682,N_1767);
or U2718 (N_2718,N_1016,N_53);
nor U2719 (N_2719,N_1385,N_1962);
or U2720 (N_2720,N_23,N_772);
nand U2721 (N_2721,N_22,N_1595);
or U2722 (N_2722,N_1598,N_346);
and U2723 (N_2723,N_336,N_1784);
or U2724 (N_2724,N_1429,N_1108);
nand U2725 (N_2725,N_184,N_1448);
nand U2726 (N_2726,N_1236,N_964);
nor U2727 (N_2727,N_1610,N_315);
and U2728 (N_2728,N_784,N_1934);
nor U2729 (N_2729,N_1632,N_903);
or U2730 (N_2730,N_981,N_1774);
nor U2731 (N_2731,N_289,N_1509);
and U2732 (N_2732,N_1045,N_1876);
nor U2733 (N_2733,N_1868,N_1175);
or U2734 (N_2734,N_1905,N_968);
nor U2735 (N_2735,N_924,N_39);
nand U2736 (N_2736,N_1719,N_129);
nor U2737 (N_2737,N_1398,N_391);
or U2738 (N_2738,N_190,N_365);
and U2739 (N_2739,N_624,N_291);
nand U2740 (N_2740,N_993,N_814);
nor U2741 (N_2741,N_1754,N_1054);
or U2742 (N_2742,N_891,N_1391);
and U2743 (N_2743,N_960,N_795);
and U2744 (N_2744,N_1831,N_444);
nor U2745 (N_2745,N_632,N_406);
or U2746 (N_2746,N_1050,N_1648);
and U2747 (N_2747,N_621,N_1462);
nor U2748 (N_2748,N_644,N_1686);
and U2749 (N_2749,N_379,N_93);
nand U2750 (N_2750,N_1654,N_1405);
nor U2751 (N_2751,N_1737,N_95);
and U2752 (N_2752,N_1253,N_595);
nor U2753 (N_2753,N_323,N_1294);
and U2754 (N_2754,N_1001,N_737);
nand U2755 (N_2755,N_931,N_1633);
nand U2756 (N_2756,N_1420,N_543);
nor U2757 (N_2757,N_937,N_1940);
nand U2758 (N_2758,N_376,N_1009);
nand U2759 (N_2759,N_618,N_111);
nor U2760 (N_2760,N_1528,N_1836);
nand U2761 (N_2761,N_1141,N_1992);
nor U2762 (N_2762,N_921,N_1973);
and U2763 (N_2763,N_1552,N_1640);
or U2764 (N_2764,N_965,N_137);
xor U2765 (N_2765,N_1397,N_1795);
and U2766 (N_2766,N_1671,N_61);
and U2767 (N_2767,N_1693,N_948);
and U2768 (N_2768,N_1891,N_1342);
and U2769 (N_2769,N_345,N_681);
and U2770 (N_2770,N_828,N_1409);
nor U2771 (N_2771,N_326,N_821);
or U2772 (N_2772,N_650,N_927);
and U2773 (N_2773,N_750,N_1256);
nand U2774 (N_2774,N_1712,N_1770);
or U2775 (N_2775,N_1262,N_1226);
and U2776 (N_2776,N_1282,N_825);
or U2777 (N_2777,N_1980,N_879);
and U2778 (N_2778,N_630,N_199);
and U2779 (N_2779,N_1008,N_1744);
nand U2780 (N_2780,N_904,N_880);
or U2781 (N_2781,N_325,N_1389);
nand U2782 (N_2782,N_1954,N_692);
nor U2783 (N_2783,N_1220,N_672);
nand U2784 (N_2784,N_1038,N_172);
nor U2785 (N_2785,N_1305,N_261);
nand U2786 (N_2786,N_76,N_1724);
and U2787 (N_2787,N_364,N_1327);
nor U2788 (N_2788,N_300,N_788);
nor U2789 (N_2789,N_1617,N_288);
nor U2790 (N_2790,N_320,N_1990);
or U2791 (N_2791,N_1736,N_581);
nand U2792 (N_2792,N_1730,N_1739);
and U2793 (N_2793,N_969,N_956);
nor U2794 (N_2794,N_259,N_1358);
nor U2795 (N_2795,N_901,N_366);
nand U2796 (N_2796,N_192,N_657);
and U2797 (N_2797,N_1931,N_1742);
nand U2798 (N_2798,N_1728,N_1864);
or U2799 (N_2799,N_356,N_854);
or U2800 (N_2800,N_1789,N_1264);
or U2801 (N_2801,N_281,N_1162);
and U2802 (N_2802,N_895,N_268);
and U2803 (N_2803,N_71,N_1982);
and U2804 (N_2804,N_40,N_661);
or U2805 (N_2805,N_943,N_718);
nand U2806 (N_2806,N_68,N_1710);
nand U2807 (N_2807,N_1755,N_286);
nor U2808 (N_2808,N_702,N_1596);
or U2809 (N_2809,N_1543,N_1213);
nand U2810 (N_2810,N_1787,N_282);
or U2811 (N_2811,N_1080,N_1567);
nor U2812 (N_2812,N_12,N_1530);
nand U2813 (N_2813,N_1056,N_1857);
and U2814 (N_2814,N_1881,N_669);
nor U2815 (N_2815,N_1659,N_354);
and U2816 (N_2816,N_368,N_1799);
or U2817 (N_2817,N_1900,N_1551);
nor U2818 (N_2818,N_1208,N_1156);
nor U2819 (N_2819,N_1616,N_434);
or U2820 (N_2820,N_285,N_813);
and U2821 (N_2821,N_614,N_1315);
or U2822 (N_2822,N_1381,N_220);
nand U2823 (N_2823,N_468,N_1861);
nand U2824 (N_2824,N_643,N_1493);
nand U2825 (N_2825,N_219,N_1375);
nand U2826 (N_2826,N_1296,N_1735);
and U2827 (N_2827,N_187,N_318);
nand U2828 (N_2828,N_1536,N_592);
or U2829 (N_2829,N_1663,N_902);
nand U2830 (N_2830,N_477,N_741);
nor U2831 (N_2831,N_1265,N_1683);
nor U2832 (N_2832,N_493,N_14);
or U2833 (N_2833,N_611,N_1423);
and U2834 (N_2834,N_994,N_1732);
nand U2835 (N_2835,N_806,N_586);
or U2836 (N_2836,N_1611,N_327);
nand U2837 (N_2837,N_899,N_1297);
and U2838 (N_2838,N_603,N_1801);
nor U2839 (N_2839,N_514,N_1145);
nor U2840 (N_2840,N_693,N_1576);
nor U2841 (N_2841,N_1853,N_267);
nor U2842 (N_2842,N_1817,N_1396);
and U2843 (N_2843,N_796,N_941);
and U2844 (N_2844,N_794,N_1845);
nand U2845 (N_2845,N_1501,N_1665);
or U2846 (N_2846,N_973,N_577);
xor U2847 (N_2847,N_594,N_954);
nand U2848 (N_2848,N_663,N_1176);
nand U2849 (N_2849,N_385,N_1478);
or U2850 (N_2850,N_120,N_1741);
and U2851 (N_2851,N_476,N_82);
or U2852 (N_2852,N_1558,N_1624);
xor U2853 (N_2853,N_706,N_1182);
nor U2854 (N_2854,N_441,N_244);
or U2855 (N_2855,N_228,N_1003);
and U2856 (N_2856,N_1955,N_124);
or U2857 (N_2857,N_1886,N_748);
and U2858 (N_2858,N_1288,N_1356);
nand U2859 (N_2859,N_257,N_1935);
xor U2860 (N_2860,N_1387,N_1618);
and U2861 (N_2861,N_1341,N_216);
or U2862 (N_2862,N_143,N_1657);
and U2863 (N_2863,N_1482,N_1364);
and U2864 (N_2864,N_1,N_947);
nand U2865 (N_2865,N_589,N_1067);
nor U2866 (N_2866,N_91,N_1311);
nand U2867 (N_2867,N_1041,N_131);
or U2868 (N_2868,N_1796,N_243);
nor U2869 (N_2869,N_1786,N_36);
or U2870 (N_2870,N_457,N_253);
nor U2871 (N_2871,N_1244,N_920);
and U2872 (N_2872,N_518,N_612);
nor U2873 (N_2873,N_566,N_272);
nand U2874 (N_2874,N_666,N_424);
or U2875 (N_2875,N_1093,N_658);
nor U2876 (N_2876,N_762,N_1522);
nand U2877 (N_2877,N_647,N_1706);
and U2878 (N_2878,N_303,N_980);
or U2879 (N_2879,N_1192,N_1190);
or U2880 (N_2880,N_1541,N_67);
or U2881 (N_2881,N_819,N_959);
and U2882 (N_2882,N_416,N_1259);
or U2883 (N_2883,N_1453,N_16);
nor U2884 (N_2884,N_164,N_1889);
nor U2885 (N_2885,N_486,N_11);
nor U2886 (N_2886,N_1765,N_1215);
nand U2887 (N_2887,N_1906,N_1521);
nand U2888 (N_2888,N_1137,N_717);
and U2889 (N_2889,N_1492,N_1075);
nand U2890 (N_2890,N_1211,N_1120);
and U2891 (N_2891,N_867,N_1820);
or U2892 (N_2892,N_1404,N_1907);
and U2893 (N_2893,N_1100,N_1722);
nand U2894 (N_2894,N_778,N_1230);
nor U2895 (N_2895,N_24,N_173);
nand U2896 (N_2896,N_1819,N_1115);
or U2897 (N_2897,N_1629,N_1042);
nor U2898 (N_2898,N_507,N_349);
nor U2899 (N_2899,N_1129,N_1566);
nor U2900 (N_2900,N_726,N_607);
and U2901 (N_2901,N_673,N_1570);
nand U2902 (N_2902,N_1456,N_703);
and U2903 (N_2903,N_208,N_374);
or U2904 (N_2904,N_628,N_1379);
or U2905 (N_2905,N_1791,N_1406);
and U2906 (N_2906,N_386,N_1756);
nand U2907 (N_2907,N_1546,N_294);
or U2908 (N_2908,N_808,N_1064);
or U2909 (N_2909,N_1489,N_81);
nand U2910 (N_2910,N_1023,N_677);
or U2911 (N_2911,N_1273,N_1626);
nand U2912 (N_2912,N_439,N_1578);
nor U2913 (N_2913,N_1637,N_395);
nand U2914 (N_2914,N_459,N_865);
or U2915 (N_2915,N_1328,N_1630);
and U2916 (N_2916,N_992,N_344);
and U2917 (N_2917,N_933,N_1126);
or U2918 (N_2918,N_787,N_1147);
and U2919 (N_2919,N_1978,N_801);
or U2920 (N_2920,N_1545,N_508);
and U2921 (N_2921,N_488,N_1027);
nor U2922 (N_2922,N_420,N_984);
or U2923 (N_2923,N_1343,N_800);
or U2924 (N_2924,N_419,N_271);
xor U2925 (N_2925,N_1386,N_278);
or U2926 (N_2926,N_238,N_287);
nand U2927 (N_2927,N_182,N_556);
nor U2928 (N_2928,N_1588,N_526);
nand U2929 (N_2929,N_757,N_1592);
nor U2930 (N_2930,N_413,N_255);
nor U2931 (N_2931,N_102,N_900);
and U2932 (N_2932,N_1673,N_1580);
or U2933 (N_2933,N_38,N_1500);
and U2934 (N_2934,N_113,N_763);
nor U2935 (N_2935,N_849,N_462);
nand U2936 (N_2936,N_1079,N_1491);
and U2937 (N_2937,N_62,N_1885);
or U2938 (N_2938,N_660,N_1582);
and U2939 (N_2939,N_1634,N_1247);
nor U2940 (N_2940,N_1073,N_816);
and U2941 (N_2941,N_429,N_1314);
nor U2942 (N_2942,N_1782,N_601);
or U2943 (N_2943,N_1766,N_47);
and U2944 (N_2944,N_1957,N_1707);
and U2945 (N_2945,N_975,N_670);
and U2946 (N_2946,N_492,N_1308);
and U2947 (N_2947,N_312,N_363);
nor U2948 (N_2948,N_222,N_535);
nor U2949 (N_2949,N_1107,N_1186);
nor U2950 (N_2950,N_1113,N_1347);
or U2951 (N_2951,N_10,N_1925);
nor U2952 (N_2952,N_635,N_739);
or U2953 (N_2953,N_1357,N_889);
and U2954 (N_2954,N_1743,N_610);
and U2955 (N_2955,N_1036,N_1218);
and U2956 (N_2956,N_515,N_1407);
and U2957 (N_2957,N_1370,N_1738);
or U2958 (N_2958,N_1435,N_1542);
nand U2959 (N_2959,N_41,N_1865);
or U2960 (N_2960,N_110,N_132);
nand U2961 (N_2961,N_1274,N_1438);
and U2962 (N_2962,N_1214,N_1053);
nand U2963 (N_2963,N_1109,N_1661);
or U2964 (N_2964,N_639,N_686);
or U2965 (N_2965,N_729,N_1979);
nor U2966 (N_2966,N_519,N_1565);
nor U2967 (N_2967,N_1871,N_1020);
nand U2968 (N_2968,N_1725,N_1144);
nor U2969 (N_2969,N_517,N_1022);
or U2970 (N_2970,N_582,N_545);
nor U2971 (N_2971,N_98,N_1460);
or U2972 (N_2972,N_465,N_1481);
nand U2973 (N_2973,N_495,N_9);
or U2974 (N_2974,N_1133,N_360);
and U2975 (N_2975,N_1414,N_605);
and U2976 (N_2976,N_513,N_1508);
and U2977 (N_2977,N_1793,N_66);
nand U2978 (N_2978,N_1757,N_283);
or U2979 (N_2979,N_619,N_1204);
and U2980 (N_2980,N_1048,N_1122);
or U2981 (N_2981,N_1600,N_1440);
and U2982 (N_2982,N_1977,N_188);
nand U2983 (N_2983,N_817,N_329);
or U2984 (N_2984,N_1452,N_1591);
nand U2985 (N_2985,N_1593,N_213);
and U2986 (N_2986,N_1241,N_332);
nand U2987 (N_2987,N_811,N_1261);
or U2988 (N_2988,N_153,N_860);
nor U2989 (N_2989,N_33,N_231);
or U2990 (N_2990,N_721,N_1018);
nand U2991 (N_2991,N_425,N_1019);
and U2992 (N_2992,N_313,N_1866);
xor U2993 (N_2993,N_1127,N_358);
and U2994 (N_2994,N_576,N_1039);
nor U2995 (N_2995,N_1458,N_1714);
or U2996 (N_2996,N_274,N_1734);
nand U2997 (N_2997,N_1590,N_485);
and U2998 (N_2998,N_185,N_1644);
nand U2999 (N_2999,N_1281,N_512);
and U3000 (N_3000,N_214,N_543);
nand U3001 (N_3001,N_1453,N_965);
nor U3002 (N_3002,N_1030,N_1919);
nand U3003 (N_3003,N_1127,N_1573);
nor U3004 (N_3004,N_1616,N_684);
and U3005 (N_3005,N_621,N_1783);
and U3006 (N_3006,N_1504,N_1869);
or U3007 (N_3007,N_212,N_1793);
or U3008 (N_3008,N_769,N_608);
nor U3009 (N_3009,N_884,N_1906);
or U3010 (N_3010,N_1733,N_1955);
nand U3011 (N_3011,N_1488,N_825);
nor U3012 (N_3012,N_344,N_177);
and U3013 (N_3013,N_1568,N_1230);
or U3014 (N_3014,N_1984,N_773);
and U3015 (N_3015,N_1106,N_1623);
nor U3016 (N_3016,N_126,N_1387);
nor U3017 (N_3017,N_176,N_872);
nor U3018 (N_3018,N_412,N_491);
and U3019 (N_3019,N_486,N_530);
nand U3020 (N_3020,N_1027,N_661);
and U3021 (N_3021,N_841,N_1141);
and U3022 (N_3022,N_35,N_1788);
or U3023 (N_3023,N_1666,N_1040);
and U3024 (N_3024,N_1683,N_526);
nor U3025 (N_3025,N_1578,N_1711);
nand U3026 (N_3026,N_220,N_1926);
and U3027 (N_3027,N_1102,N_1617);
or U3028 (N_3028,N_1368,N_434);
or U3029 (N_3029,N_928,N_826);
nor U3030 (N_3030,N_407,N_794);
nor U3031 (N_3031,N_931,N_1814);
nor U3032 (N_3032,N_1702,N_1204);
and U3033 (N_3033,N_1931,N_1721);
and U3034 (N_3034,N_352,N_1204);
nand U3035 (N_3035,N_696,N_460);
xor U3036 (N_3036,N_1315,N_1933);
nor U3037 (N_3037,N_399,N_1944);
nand U3038 (N_3038,N_1371,N_1213);
and U3039 (N_3039,N_672,N_1590);
or U3040 (N_3040,N_1501,N_1446);
or U3041 (N_3041,N_612,N_485);
and U3042 (N_3042,N_1956,N_1238);
nand U3043 (N_3043,N_543,N_235);
and U3044 (N_3044,N_1498,N_1932);
nor U3045 (N_3045,N_393,N_470);
or U3046 (N_3046,N_997,N_387);
nand U3047 (N_3047,N_997,N_1574);
nand U3048 (N_3048,N_677,N_749);
nor U3049 (N_3049,N_599,N_1813);
or U3050 (N_3050,N_391,N_1544);
and U3051 (N_3051,N_610,N_1351);
or U3052 (N_3052,N_1843,N_688);
nand U3053 (N_3053,N_1787,N_1923);
nor U3054 (N_3054,N_1961,N_1125);
nor U3055 (N_3055,N_821,N_1452);
nor U3056 (N_3056,N_384,N_868);
or U3057 (N_3057,N_1087,N_660);
nor U3058 (N_3058,N_1773,N_710);
or U3059 (N_3059,N_38,N_671);
or U3060 (N_3060,N_1450,N_1297);
xnor U3061 (N_3061,N_401,N_1592);
and U3062 (N_3062,N_1226,N_364);
nand U3063 (N_3063,N_640,N_1545);
nor U3064 (N_3064,N_1056,N_1893);
nand U3065 (N_3065,N_511,N_1153);
nor U3066 (N_3066,N_608,N_352);
and U3067 (N_3067,N_1427,N_547);
nand U3068 (N_3068,N_376,N_223);
or U3069 (N_3069,N_1319,N_38);
nand U3070 (N_3070,N_700,N_190);
or U3071 (N_3071,N_766,N_1715);
nor U3072 (N_3072,N_779,N_1984);
nor U3073 (N_3073,N_1444,N_274);
nand U3074 (N_3074,N_260,N_1380);
nor U3075 (N_3075,N_367,N_676);
nor U3076 (N_3076,N_1616,N_1715);
xor U3077 (N_3077,N_1370,N_1775);
and U3078 (N_3078,N_1023,N_107);
nor U3079 (N_3079,N_500,N_608);
nor U3080 (N_3080,N_324,N_991);
nor U3081 (N_3081,N_292,N_327);
nand U3082 (N_3082,N_1608,N_739);
nand U3083 (N_3083,N_770,N_1006);
or U3084 (N_3084,N_294,N_147);
or U3085 (N_3085,N_53,N_1872);
or U3086 (N_3086,N_1945,N_549);
nor U3087 (N_3087,N_426,N_1980);
nand U3088 (N_3088,N_815,N_649);
and U3089 (N_3089,N_41,N_1657);
and U3090 (N_3090,N_1236,N_733);
nor U3091 (N_3091,N_532,N_1093);
nand U3092 (N_3092,N_1164,N_1292);
and U3093 (N_3093,N_1301,N_877);
or U3094 (N_3094,N_1345,N_1061);
or U3095 (N_3095,N_653,N_1067);
or U3096 (N_3096,N_796,N_1311);
nand U3097 (N_3097,N_177,N_86);
nand U3098 (N_3098,N_1306,N_1753);
nor U3099 (N_3099,N_812,N_1231);
nand U3100 (N_3100,N_1265,N_126);
or U3101 (N_3101,N_990,N_1698);
and U3102 (N_3102,N_479,N_832);
and U3103 (N_3103,N_1166,N_1488);
and U3104 (N_3104,N_1678,N_924);
and U3105 (N_3105,N_1439,N_424);
nand U3106 (N_3106,N_472,N_1969);
or U3107 (N_3107,N_981,N_557);
xor U3108 (N_3108,N_203,N_1415);
or U3109 (N_3109,N_1889,N_725);
nor U3110 (N_3110,N_841,N_790);
nand U3111 (N_3111,N_1966,N_1496);
nor U3112 (N_3112,N_1181,N_971);
xnor U3113 (N_3113,N_1089,N_1516);
nor U3114 (N_3114,N_1466,N_65);
or U3115 (N_3115,N_327,N_348);
and U3116 (N_3116,N_668,N_1718);
nor U3117 (N_3117,N_297,N_1905);
nor U3118 (N_3118,N_464,N_468);
nor U3119 (N_3119,N_1611,N_1690);
or U3120 (N_3120,N_658,N_1066);
nand U3121 (N_3121,N_952,N_259);
nand U3122 (N_3122,N_1841,N_14);
or U3123 (N_3123,N_1103,N_177);
and U3124 (N_3124,N_1126,N_1021);
nand U3125 (N_3125,N_1900,N_259);
nand U3126 (N_3126,N_10,N_71);
or U3127 (N_3127,N_1324,N_1100);
and U3128 (N_3128,N_1049,N_1544);
or U3129 (N_3129,N_1728,N_1677);
nor U3130 (N_3130,N_1012,N_875);
or U3131 (N_3131,N_56,N_1878);
nand U3132 (N_3132,N_1711,N_1073);
and U3133 (N_3133,N_1792,N_750);
xor U3134 (N_3134,N_1510,N_1598);
nand U3135 (N_3135,N_1503,N_1284);
nor U3136 (N_3136,N_1129,N_1629);
nand U3137 (N_3137,N_387,N_1723);
and U3138 (N_3138,N_440,N_180);
nand U3139 (N_3139,N_564,N_1632);
and U3140 (N_3140,N_213,N_1360);
nand U3141 (N_3141,N_285,N_413);
nor U3142 (N_3142,N_1872,N_328);
or U3143 (N_3143,N_943,N_860);
nand U3144 (N_3144,N_521,N_1177);
nor U3145 (N_3145,N_1574,N_490);
and U3146 (N_3146,N_1550,N_1895);
nand U3147 (N_3147,N_132,N_497);
and U3148 (N_3148,N_290,N_894);
and U3149 (N_3149,N_1028,N_1831);
nor U3150 (N_3150,N_467,N_1289);
nor U3151 (N_3151,N_734,N_1949);
or U3152 (N_3152,N_181,N_736);
nand U3153 (N_3153,N_10,N_1728);
or U3154 (N_3154,N_1079,N_1066);
and U3155 (N_3155,N_635,N_1233);
or U3156 (N_3156,N_1158,N_1750);
nand U3157 (N_3157,N_204,N_1169);
and U3158 (N_3158,N_649,N_88);
or U3159 (N_3159,N_1846,N_1779);
nor U3160 (N_3160,N_482,N_1669);
nor U3161 (N_3161,N_26,N_153);
nand U3162 (N_3162,N_1792,N_1406);
and U3163 (N_3163,N_689,N_1967);
nand U3164 (N_3164,N_314,N_497);
nand U3165 (N_3165,N_1599,N_474);
or U3166 (N_3166,N_434,N_233);
nand U3167 (N_3167,N_1059,N_1274);
nand U3168 (N_3168,N_474,N_1029);
nand U3169 (N_3169,N_1896,N_336);
nand U3170 (N_3170,N_285,N_441);
or U3171 (N_3171,N_1689,N_842);
or U3172 (N_3172,N_1893,N_898);
nand U3173 (N_3173,N_1737,N_1065);
or U3174 (N_3174,N_1071,N_1625);
and U3175 (N_3175,N_616,N_726);
nand U3176 (N_3176,N_672,N_1027);
nor U3177 (N_3177,N_1941,N_1931);
nor U3178 (N_3178,N_1658,N_242);
nor U3179 (N_3179,N_91,N_1238);
nor U3180 (N_3180,N_462,N_904);
or U3181 (N_3181,N_1330,N_972);
nor U3182 (N_3182,N_183,N_1168);
nand U3183 (N_3183,N_1877,N_1063);
nor U3184 (N_3184,N_1587,N_866);
or U3185 (N_3185,N_73,N_287);
or U3186 (N_3186,N_1056,N_360);
nor U3187 (N_3187,N_706,N_1786);
nor U3188 (N_3188,N_868,N_1587);
nand U3189 (N_3189,N_295,N_346);
and U3190 (N_3190,N_1132,N_511);
or U3191 (N_3191,N_1648,N_1623);
nor U3192 (N_3192,N_1346,N_661);
or U3193 (N_3193,N_1356,N_1752);
or U3194 (N_3194,N_1764,N_1476);
nand U3195 (N_3195,N_209,N_384);
and U3196 (N_3196,N_1336,N_1420);
or U3197 (N_3197,N_883,N_1232);
or U3198 (N_3198,N_324,N_370);
or U3199 (N_3199,N_1205,N_253);
and U3200 (N_3200,N_862,N_1310);
nor U3201 (N_3201,N_1453,N_1760);
nand U3202 (N_3202,N_76,N_852);
or U3203 (N_3203,N_68,N_1617);
nand U3204 (N_3204,N_1834,N_333);
or U3205 (N_3205,N_363,N_1693);
and U3206 (N_3206,N_511,N_729);
and U3207 (N_3207,N_1177,N_920);
nor U3208 (N_3208,N_334,N_1170);
nand U3209 (N_3209,N_932,N_1160);
nand U3210 (N_3210,N_1515,N_953);
nand U3211 (N_3211,N_768,N_751);
nor U3212 (N_3212,N_28,N_1904);
nand U3213 (N_3213,N_1893,N_315);
nand U3214 (N_3214,N_1486,N_1545);
nor U3215 (N_3215,N_1174,N_883);
nor U3216 (N_3216,N_926,N_169);
or U3217 (N_3217,N_1467,N_1894);
nand U3218 (N_3218,N_701,N_962);
and U3219 (N_3219,N_420,N_861);
nand U3220 (N_3220,N_1206,N_1931);
and U3221 (N_3221,N_1242,N_113);
nand U3222 (N_3222,N_474,N_1260);
xor U3223 (N_3223,N_1762,N_1748);
nand U3224 (N_3224,N_1076,N_682);
or U3225 (N_3225,N_744,N_477);
or U3226 (N_3226,N_798,N_105);
nor U3227 (N_3227,N_164,N_1131);
nand U3228 (N_3228,N_458,N_1181);
nor U3229 (N_3229,N_490,N_619);
nand U3230 (N_3230,N_1479,N_758);
or U3231 (N_3231,N_1346,N_1917);
nand U3232 (N_3232,N_741,N_869);
nor U3233 (N_3233,N_102,N_258);
or U3234 (N_3234,N_1224,N_865);
nor U3235 (N_3235,N_15,N_1154);
and U3236 (N_3236,N_1870,N_93);
nand U3237 (N_3237,N_1382,N_1036);
or U3238 (N_3238,N_166,N_453);
nand U3239 (N_3239,N_765,N_812);
nor U3240 (N_3240,N_415,N_128);
and U3241 (N_3241,N_103,N_1407);
nor U3242 (N_3242,N_1423,N_1113);
and U3243 (N_3243,N_972,N_1515);
or U3244 (N_3244,N_1267,N_776);
nor U3245 (N_3245,N_1467,N_622);
or U3246 (N_3246,N_1757,N_573);
or U3247 (N_3247,N_457,N_1984);
xnor U3248 (N_3248,N_1151,N_593);
and U3249 (N_3249,N_6,N_1131);
nor U3250 (N_3250,N_1100,N_1038);
and U3251 (N_3251,N_318,N_206);
and U3252 (N_3252,N_1503,N_784);
nand U3253 (N_3253,N_470,N_1209);
or U3254 (N_3254,N_825,N_370);
nor U3255 (N_3255,N_175,N_1107);
and U3256 (N_3256,N_926,N_361);
nand U3257 (N_3257,N_1198,N_864);
or U3258 (N_3258,N_1045,N_248);
and U3259 (N_3259,N_1840,N_1531);
nand U3260 (N_3260,N_1655,N_1148);
xnor U3261 (N_3261,N_1421,N_1819);
or U3262 (N_3262,N_1124,N_1854);
nor U3263 (N_3263,N_608,N_1989);
nand U3264 (N_3264,N_1030,N_638);
nand U3265 (N_3265,N_697,N_1881);
or U3266 (N_3266,N_698,N_743);
and U3267 (N_3267,N_53,N_102);
and U3268 (N_3268,N_562,N_799);
and U3269 (N_3269,N_65,N_142);
or U3270 (N_3270,N_1630,N_1680);
and U3271 (N_3271,N_280,N_814);
or U3272 (N_3272,N_590,N_1806);
nor U3273 (N_3273,N_1409,N_816);
nand U3274 (N_3274,N_1873,N_1715);
nor U3275 (N_3275,N_697,N_731);
nor U3276 (N_3276,N_476,N_449);
and U3277 (N_3277,N_1452,N_745);
nand U3278 (N_3278,N_1879,N_898);
or U3279 (N_3279,N_83,N_240);
and U3280 (N_3280,N_39,N_281);
or U3281 (N_3281,N_626,N_1594);
nor U3282 (N_3282,N_1842,N_1113);
nor U3283 (N_3283,N_1929,N_884);
nand U3284 (N_3284,N_567,N_755);
or U3285 (N_3285,N_1435,N_1883);
or U3286 (N_3286,N_90,N_794);
and U3287 (N_3287,N_554,N_535);
nand U3288 (N_3288,N_381,N_373);
and U3289 (N_3289,N_1693,N_1347);
nand U3290 (N_3290,N_615,N_1893);
nand U3291 (N_3291,N_404,N_1269);
and U3292 (N_3292,N_1275,N_782);
and U3293 (N_3293,N_1867,N_888);
or U3294 (N_3294,N_146,N_1774);
nand U3295 (N_3295,N_167,N_588);
nand U3296 (N_3296,N_31,N_1944);
and U3297 (N_3297,N_301,N_202);
nor U3298 (N_3298,N_1879,N_1283);
nor U3299 (N_3299,N_955,N_1194);
nand U3300 (N_3300,N_576,N_1157);
and U3301 (N_3301,N_1223,N_1301);
or U3302 (N_3302,N_190,N_1120);
or U3303 (N_3303,N_658,N_803);
nor U3304 (N_3304,N_227,N_767);
nand U3305 (N_3305,N_685,N_1169);
nor U3306 (N_3306,N_1870,N_905);
nor U3307 (N_3307,N_893,N_1032);
xnor U3308 (N_3308,N_328,N_546);
and U3309 (N_3309,N_1075,N_417);
nor U3310 (N_3310,N_18,N_818);
nand U3311 (N_3311,N_466,N_710);
nand U3312 (N_3312,N_472,N_422);
nand U3313 (N_3313,N_608,N_1832);
nand U3314 (N_3314,N_1397,N_433);
nor U3315 (N_3315,N_621,N_863);
nor U3316 (N_3316,N_1529,N_1550);
xnor U3317 (N_3317,N_67,N_379);
or U3318 (N_3318,N_635,N_188);
or U3319 (N_3319,N_1111,N_1795);
or U3320 (N_3320,N_744,N_534);
and U3321 (N_3321,N_1053,N_1025);
nor U3322 (N_3322,N_787,N_1612);
nor U3323 (N_3323,N_74,N_1848);
or U3324 (N_3324,N_828,N_746);
nor U3325 (N_3325,N_293,N_1953);
nand U3326 (N_3326,N_1719,N_60);
nand U3327 (N_3327,N_1702,N_1769);
nand U3328 (N_3328,N_1589,N_329);
nand U3329 (N_3329,N_1572,N_1907);
nor U3330 (N_3330,N_1969,N_1852);
or U3331 (N_3331,N_902,N_1537);
or U3332 (N_3332,N_1858,N_568);
nand U3333 (N_3333,N_888,N_304);
and U3334 (N_3334,N_1210,N_1368);
nand U3335 (N_3335,N_686,N_399);
and U3336 (N_3336,N_1727,N_1247);
or U3337 (N_3337,N_1508,N_1494);
nor U3338 (N_3338,N_713,N_28);
xnor U3339 (N_3339,N_1967,N_287);
nand U3340 (N_3340,N_838,N_1257);
nor U3341 (N_3341,N_712,N_1169);
and U3342 (N_3342,N_785,N_1356);
xor U3343 (N_3343,N_445,N_770);
or U3344 (N_3344,N_968,N_655);
nor U3345 (N_3345,N_842,N_368);
and U3346 (N_3346,N_1945,N_411);
nand U3347 (N_3347,N_1987,N_969);
or U3348 (N_3348,N_567,N_1679);
nand U3349 (N_3349,N_1337,N_1003);
nor U3350 (N_3350,N_1792,N_1621);
nand U3351 (N_3351,N_768,N_451);
or U3352 (N_3352,N_1559,N_149);
or U3353 (N_3353,N_167,N_932);
or U3354 (N_3354,N_1314,N_1862);
nor U3355 (N_3355,N_1866,N_261);
nor U3356 (N_3356,N_511,N_1938);
nor U3357 (N_3357,N_1125,N_314);
nand U3358 (N_3358,N_1975,N_497);
nand U3359 (N_3359,N_1997,N_1787);
and U3360 (N_3360,N_1140,N_1603);
or U3361 (N_3361,N_1217,N_1017);
nor U3362 (N_3362,N_865,N_265);
nor U3363 (N_3363,N_116,N_1214);
and U3364 (N_3364,N_1789,N_417);
and U3365 (N_3365,N_1897,N_1048);
or U3366 (N_3366,N_41,N_203);
nor U3367 (N_3367,N_1054,N_1707);
nor U3368 (N_3368,N_909,N_1535);
nor U3369 (N_3369,N_705,N_1025);
nor U3370 (N_3370,N_1878,N_1116);
and U3371 (N_3371,N_860,N_1680);
nand U3372 (N_3372,N_1538,N_1856);
nor U3373 (N_3373,N_1966,N_1337);
or U3374 (N_3374,N_1413,N_1855);
and U3375 (N_3375,N_588,N_48);
nand U3376 (N_3376,N_1258,N_173);
and U3377 (N_3377,N_95,N_173);
nor U3378 (N_3378,N_501,N_1621);
and U3379 (N_3379,N_684,N_1401);
and U3380 (N_3380,N_1654,N_1423);
nor U3381 (N_3381,N_562,N_530);
or U3382 (N_3382,N_95,N_138);
or U3383 (N_3383,N_1042,N_448);
and U3384 (N_3384,N_147,N_783);
nand U3385 (N_3385,N_961,N_151);
nand U3386 (N_3386,N_1959,N_512);
or U3387 (N_3387,N_1164,N_1758);
nor U3388 (N_3388,N_689,N_1671);
nor U3389 (N_3389,N_1930,N_1883);
and U3390 (N_3390,N_1741,N_163);
nor U3391 (N_3391,N_1937,N_893);
and U3392 (N_3392,N_1176,N_1088);
or U3393 (N_3393,N_1542,N_1035);
and U3394 (N_3394,N_162,N_571);
nand U3395 (N_3395,N_1583,N_1178);
nor U3396 (N_3396,N_344,N_963);
and U3397 (N_3397,N_1175,N_1975);
nand U3398 (N_3398,N_523,N_822);
and U3399 (N_3399,N_998,N_679);
and U3400 (N_3400,N_778,N_1956);
nand U3401 (N_3401,N_1106,N_1026);
and U3402 (N_3402,N_259,N_1091);
nand U3403 (N_3403,N_1943,N_750);
nor U3404 (N_3404,N_1641,N_1090);
nand U3405 (N_3405,N_1847,N_1631);
nand U3406 (N_3406,N_891,N_233);
nand U3407 (N_3407,N_1419,N_529);
nor U3408 (N_3408,N_159,N_1513);
nand U3409 (N_3409,N_680,N_1930);
nand U3410 (N_3410,N_462,N_1524);
or U3411 (N_3411,N_241,N_1781);
or U3412 (N_3412,N_1631,N_65);
nand U3413 (N_3413,N_1932,N_1115);
nor U3414 (N_3414,N_1918,N_1083);
and U3415 (N_3415,N_1092,N_1603);
and U3416 (N_3416,N_1279,N_236);
nand U3417 (N_3417,N_325,N_108);
and U3418 (N_3418,N_1632,N_745);
and U3419 (N_3419,N_1499,N_144);
nor U3420 (N_3420,N_130,N_609);
nor U3421 (N_3421,N_681,N_1399);
nor U3422 (N_3422,N_1398,N_1058);
and U3423 (N_3423,N_612,N_812);
nand U3424 (N_3424,N_1845,N_541);
nor U3425 (N_3425,N_1508,N_45);
or U3426 (N_3426,N_1711,N_538);
nand U3427 (N_3427,N_115,N_866);
nand U3428 (N_3428,N_310,N_167);
nor U3429 (N_3429,N_234,N_1555);
and U3430 (N_3430,N_1419,N_849);
nor U3431 (N_3431,N_244,N_1148);
or U3432 (N_3432,N_235,N_452);
nand U3433 (N_3433,N_948,N_1568);
nor U3434 (N_3434,N_1468,N_1600);
or U3435 (N_3435,N_257,N_1506);
nor U3436 (N_3436,N_1408,N_1969);
or U3437 (N_3437,N_1185,N_150);
or U3438 (N_3438,N_339,N_17);
and U3439 (N_3439,N_1788,N_292);
or U3440 (N_3440,N_1545,N_641);
nor U3441 (N_3441,N_262,N_1615);
nand U3442 (N_3442,N_808,N_1836);
or U3443 (N_3443,N_1726,N_365);
and U3444 (N_3444,N_621,N_1784);
nor U3445 (N_3445,N_1353,N_661);
and U3446 (N_3446,N_1471,N_1549);
or U3447 (N_3447,N_1282,N_1212);
or U3448 (N_3448,N_1070,N_1662);
or U3449 (N_3449,N_254,N_844);
or U3450 (N_3450,N_424,N_743);
and U3451 (N_3451,N_1981,N_281);
nor U3452 (N_3452,N_1710,N_1644);
nand U3453 (N_3453,N_35,N_165);
and U3454 (N_3454,N_963,N_1624);
nand U3455 (N_3455,N_860,N_1026);
or U3456 (N_3456,N_1681,N_828);
and U3457 (N_3457,N_626,N_300);
nand U3458 (N_3458,N_903,N_1225);
and U3459 (N_3459,N_1668,N_1660);
nor U3460 (N_3460,N_1195,N_1306);
or U3461 (N_3461,N_1004,N_1220);
nor U3462 (N_3462,N_100,N_266);
and U3463 (N_3463,N_70,N_939);
nand U3464 (N_3464,N_733,N_1122);
nand U3465 (N_3465,N_1421,N_438);
nor U3466 (N_3466,N_1531,N_390);
nand U3467 (N_3467,N_1897,N_81);
or U3468 (N_3468,N_876,N_1171);
and U3469 (N_3469,N_277,N_1281);
nor U3470 (N_3470,N_1406,N_1806);
or U3471 (N_3471,N_219,N_1541);
nor U3472 (N_3472,N_1932,N_1601);
xnor U3473 (N_3473,N_119,N_1784);
nand U3474 (N_3474,N_1601,N_1524);
and U3475 (N_3475,N_1333,N_1282);
nor U3476 (N_3476,N_341,N_1469);
nand U3477 (N_3477,N_917,N_580);
and U3478 (N_3478,N_247,N_100);
nor U3479 (N_3479,N_319,N_97);
or U3480 (N_3480,N_447,N_748);
nand U3481 (N_3481,N_315,N_449);
nor U3482 (N_3482,N_1615,N_1746);
nor U3483 (N_3483,N_526,N_1250);
or U3484 (N_3484,N_1606,N_1457);
nor U3485 (N_3485,N_1714,N_571);
and U3486 (N_3486,N_1282,N_1992);
or U3487 (N_3487,N_705,N_943);
nor U3488 (N_3488,N_583,N_532);
nor U3489 (N_3489,N_326,N_1201);
or U3490 (N_3490,N_464,N_542);
nand U3491 (N_3491,N_836,N_1064);
or U3492 (N_3492,N_645,N_1251);
or U3493 (N_3493,N_1019,N_434);
nor U3494 (N_3494,N_1822,N_711);
or U3495 (N_3495,N_924,N_1439);
and U3496 (N_3496,N_1661,N_128);
or U3497 (N_3497,N_532,N_1767);
and U3498 (N_3498,N_622,N_1099);
nor U3499 (N_3499,N_396,N_1398);
nor U3500 (N_3500,N_604,N_997);
nand U3501 (N_3501,N_1536,N_19);
and U3502 (N_3502,N_860,N_266);
nand U3503 (N_3503,N_712,N_1508);
nor U3504 (N_3504,N_427,N_421);
nand U3505 (N_3505,N_769,N_380);
nor U3506 (N_3506,N_1525,N_1547);
nand U3507 (N_3507,N_1925,N_1493);
nor U3508 (N_3508,N_127,N_182);
nor U3509 (N_3509,N_366,N_506);
or U3510 (N_3510,N_1939,N_117);
or U3511 (N_3511,N_78,N_691);
nand U3512 (N_3512,N_1246,N_867);
nor U3513 (N_3513,N_743,N_1464);
nor U3514 (N_3514,N_1173,N_1652);
or U3515 (N_3515,N_851,N_179);
and U3516 (N_3516,N_922,N_1073);
and U3517 (N_3517,N_1172,N_941);
nand U3518 (N_3518,N_1749,N_868);
nor U3519 (N_3519,N_542,N_783);
or U3520 (N_3520,N_715,N_447);
and U3521 (N_3521,N_1761,N_1135);
and U3522 (N_3522,N_375,N_785);
nand U3523 (N_3523,N_411,N_1431);
nand U3524 (N_3524,N_1786,N_1082);
and U3525 (N_3525,N_1714,N_1733);
or U3526 (N_3526,N_1902,N_1118);
or U3527 (N_3527,N_98,N_475);
or U3528 (N_3528,N_602,N_285);
nand U3529 (N_3529,N_882,N_181);
or U3530 (N_3530,N_1670,N_1671);
nand U3531 (N_3531,N_1926,N_569);
nor U3532 (N_3532,N_1592,N_1743);
nand U3533 (N_3533,N_1772,N_327);
nor U3534 (N_3534,N_1758,N_1248);
or U3535 (N_3535,N_918,N_1890);
nor U3536 (N_3536,N_643,N_1896);
or U3537 (N_3537,N_1228,N_1464);
and U3538 (N_3538,N_1045,N_1595);
or U3539 (N_3539,N_802,N_398);
and U3540 (N_3540,N_1352,N_1974);
and U3541 (N_3541,N_1926,N_831);
nand U3542 (N_3542,N_1964,N_1214);
and U3543 (N_3543,N_441,N_343);
nand U3544 (N_3544,N_474,N_1911);
and U3545 (N_3545,N_47,N_1321);
and U3546 (N_3546,N_632,N_48);
or U3547 (N_3547,N_1099,N_1694);
or U3548 (N_3548,N_895,N_1114);
nor U3549 (N_3549,N_1309,N_657);
nand U3550 (N_3550,N_636,N_1934);
or U3551 (N_3551,N_431,N_480);
or U3552 (N_3552,N_642,N_1189);
or U3553 (N_3553,N_1974,N_1937);
or U3554 (N_3554,N_78,N_369);
or U3555 (N_3555,N_865,N_1757);
nand U3556 (N_3556,N_1192,N_401);
or U3557 (N_3557,N_1716,N_1137);
and U3558 (N_3558,N_1810,N_283);
and U3559 (N_3559,N_925,N_1001);
and U3560 (N_3560,N_769,N_1266);
and U3561 (N_3561,N_1870,N_633);
nor U3562 (N_3562,N_1974,N_1863);
and U3563 (N_3563,N_225,N_415);
or U3564 (N_3564,N_771,N_1716);
and U3565 (N_3565,N_326,N_239);
nor U3566 (N_3566,N_1198,N_367);
nor U3567 (N_3567,N_229,N_1370);
nor U3568 (N_3568,N_1388,N_1350);
nand U3569 (N_3569,N_1583,N_412);
or U3570 (N_3570,N_607,N_266);
or U3571 (N_3571,N_1899,N_688);
or U3572 (N_3572,N_1750,N_465);
nand U3573 (N_3573,N_515,N_1742);
nand U3574 (N_3574,N_1377,N_867);
or U3575 (N_3575,N_1350,N_595);
nor U3576 (N_3576,N_1657,N_1140);
or U3577 (N_3577,N_1475,N_1055);
and U3578 (N_3578,N_1989,N_287);
or U3579 (N_3579,N_1477,N_1855);
and U3580 (N_3580,N_1167,N_836);
nand U3581 (N_3581,N_1161,N_1052);
nand U3582 (N_3582,N_1657,N_563);
nand U3583 (N_3583,N_17,N_570);
or U3584 (N_3584,N_901,N_549);
nor U3585 (N_3585,N_1271,N_826);
nand U3586 (N_3586,N_1713,N_32);
nor U3587 (N_3587,N_1365,N_1486);
nor U3588 (N_3588,N_197,N_1817);
nand U3589 (N_3589,N_1155,N_282);
nor U3590 (N_3590,N_525,N_747);
nor U3591 (N_3591,N_1589,N_1201);
nand U3592 (N_3592,N_1803,N_830);
nor U3593 (N_3593,N_307,N_998);
or U3594 (N_3594,N_1368,N_169);
nand U3595 (N_3595,N_1801,N_1444);
and U3596 (N_3596,N_629,N_1412);
nand U3597 (N_3597,N_167,N_1324);
or U3598 (N_3598,N_30,N_1562);
and U3599 (N_3599,N_691,N_87);
nand U3600 (N_3600,N_980,N_1672);
nand U3601 (N_3601,N_311,N_1538);
nor U3602 (N_3602,N_1636,N_1370);
and U3603 (N_3603,N_1475,N_371);
nand U3604 (N_3604,N_259,N_1565);
nand U3605 (N_3605,N_1112,N_1373);
or U3606 (N_3606,N_609,N_8);
nor U3607 (N_3607,N_1019,N_378);
nor U3608 (N_3608,N_436,N_980);
and U3609 (N_3609,N_1106,N_1136);
nor U3610 (N_3610,N_873,N_1303);
nor U3611 (N_3611,N_725,N_1891);
or U3612 (N_3612,N_1517,N_719);
or U3613 (N_3613,N_1886,N_551);
xnor U3614 (N_3614,N_122,N_1219);
or U3615 (N_3615,N_1546,N_53);
or U3616 (N_3616,N_1673,N_758);
and U3617 (N_3617,N_856,N_1173);
nand U3618 (N_3618,N_1678,N_747);
nor U3619 (N_3619,N_631,N_7);
and U3620 (N_3620,N_1407,N_1469);
nand U3621 (N_3621,N_722,N_1955);
nand U3622 (N_3622,N_1252,N_1349);
and U3623 (N_3623,N_62,N_254);
or U3624 (N_3624,N_590,N_766);
or U3625 (N_3625,N_1109,N_1866);
nand U3626 (N_3626,N_927,N_1735);
nand U3627 (N_3627,N_416,N_533);
nand U3628 (N_3628,N_1515,N_238);
nand U3629 (N_3629,N_1766,N_1300);
nand U3630 (N_3630,N_782,N_1079);
nor U3631 (N_3631,N_1006,N_268);
and U3632 (N_3632,N_609,N_1767);
or U3633 (N_3633,N_1687,N_1902);
nor U3634 (N_3634,N_1494,N_1129);
nand U3635 (N_3635,N_878,N_1707);
or U3636 (N_3636,N_880,N_1415);
nand U3637 (N_3637,N_624,N_1620);
nand U3638 (N_3638,N_1387,N_925);
nor U3639 (N_3639,N_759,N_1269);
nor U3640 (N_3640,N_549,N_265);
and U3641 (N_3641,N_171,N_1611);
nor U3642 (N_3642,N_315,N_387);
and U3643 (N_3643,N_544,N_1943);
and U3644 (N_3644,N_72,N_600);
and U3645 (N_3645,N_415,N_10);
nor U3646 (N_3646,N_838,N_1752);
nand U3647 (N_3647,N_1090,N_956);
or U3648 (N_3648,N_1005,N_812);
nand U3649 (N_3649,N_1899,N_371);
and U3650 (N_3650,N_672,N_327);
or U3651 (N_3651,N_1438,N_501);
nand U3652 (N_3652,N_1730,N_927);
nor U3653 (N_3653,N_72,N_253);
and U3654 (N_3654,N_510,N_902);
and U3655 (N_3655,N_297,N_129);
or U3656 (N_3656,N_791,N_737);
or U3657 (N_3657,N_1080,N_713);
nand U3658 (N_3658,N_1457,N_569);
or U3659 (N_3659,N_1472,N_1253);
nand U3660 (N_3660,N_509,N_1571);
and U3661 (N_3661,N_130,N_238);
nor U3662 (N_3662,N_816,N_1744);
nand U3663 (N_3663,N_1269,N_1293);
or U3664 (N_3664,N_678,N_1977);
nor U3665 (N_3665,N_801,N_142);
nor U3666 (N_3666,N_425,N_1670);
and U3667 (N_3667,N_1380,N_1088);
or U3668 (N_3668,N_968,N_1711);
nor U3669 (N_3669,N_398,N_1586);
nand U3670 (N_3670,N_879,N_845);
nand U3671 (N_3671,N_1367,N_1236);
and U3672 (N_3672,N_1062,N_1626);
or U3673 (N_3673,N_450,N_1280);
nor U3674 (N_3674,N_788,N_237);
or U3675 (N_3675,N_1104,N_1369);
nor U3676 (N_3676,N_1338,N_1831);
nor U3677 (N_3677,N_1573,N_940);
nand U3678 (N_3678,N_761,N_1689);
and U3679 (N_3679,N_1997,N_509);
nor U3680 (N_3680,N_1364,N_715);
or U3681 (N_3681,N_1661,N_829);
nor U3682 (N_3682,N_1326,N_1586);
or U3683 (N_3683,N_1019,N_999);
nor U3684 (N_3684,N_793,N_709);
nand U3685 (N_3685,N_1875,N_101);
nand U3686 (N_3686,N_1518,N_1064);
nand U3687 (N_3687,N_542,N_1002);
or U3688 (N_3688,N_1904,N_297);
and U3689 (N_3689,N_1801,N_846);
or U3690 (N_3690,N_988,N_1391);
nor U3691 (N_3691,N_1387,N_967);
nor U3692 (N_3692,N_337,N_1966);
xor U3693 (N_3693,N_1927,N_205);
nand U3694 (N_3694,N_1062,N_1225);
and U3695 (N_3695,N_1452,N_885);
nand U3696 (N_3696,N_52,N_1666);
nor U3697 (N_3697,N_1633,N_1948);
and U3698 (N_3698,N_1418,N_469);
or U3699 (N_3699,N_1166,N_1863);
or U3700 (N_3700,N_1126,N_1336);
or U3701 (N_3701,N_1462,N_754);
nor U3702 (N_3702,N_1405,N_1101);
and U3703 (N_3703,N_440,N_245);
nand U3704 (N_3704,N_1735,N_1812);
and U3705 (N_3705,N_1365,N_484);
nand U3706 (N_3706,N_1433,N_814);
and U3707 (N_3707,N_546,N_829);
nand U3708 (N_3708,N_280,N_144);
nor U3709 (N_3709,N_1120,N_217);
nand U3710 (N_3710,N_336,N_765);
and U3711 (N_3711,N_561,N_983);
or U3712 (N_3712,N_124,N_1179);
and U3713 (N_3713,N_384,N_736);
nor U3714 (N_3714,N_1634,N_1087);
nor U3715 (N_3715,N_903,N_1232);
nand U3716 (N_3716,N_1465,N_1886);
nor U3717 (N_3717,N_1238,N_1147);
nor U3718 (N_3718,N_1044,N_1812);
or U3719 (N_3719,N_838,N_854);
and U3720 (N_3720,N_498,N_1136);
nor U3721 (N_3721,N_1207,N_892);
xor U3722 (N_3722,N_355,N_810);
nor U3723 (N_3723,N_1585,N_1375);
nor U3724 (N_3724,N_1338,N_7);
or U3725 (N_3725,N_372,N_254);
or U3726 (N_3726,N_631,N_1696);
nor U3727 (N_3727,N_1639,N_1445);
or U3728 (N_3728,N_1620,N_1203);
and U3729 (N_3729,N_1448,N_1972);
nand U3730 (N_3730,N_1556,N_353);
nor U3731 (N_3731,N_754,N_1403);
or U3732 (N_3732,N_286,N_803);
nor U3733 (N_3733,N_276,N_389);
nor U3734 (N_3734,N_1110,N_1204);
nand U3735 (N_3735,N_410,N_31);
nand U3736 (N_3736,N_1404,N_1898);
nand U3737 (N_3737,N_1248,N_897);
nand U3738 (N_3738,N_789,N_999);
or U3739 (N_3739,N_1688,N_1025);
or U3740 (N_3740,N_53,N_784);
nand U3741 (N_3741,N_1154,N_801);
and U3742 (N_3742,N_409,N_1383);
and U3743 (N_3743,N_1732,N_1775);
and U3744 (N_3744,N_487,N_322);
and U3745 (N_3745,N_1330,N_1772);
or U3746 (N_3746,N_138,N_1153);
nand U3747 (N_3747,N_259,N_1222);
or U3748 (N_3748,N_1957,N_141);
nor U3749 (N_3749,N_320,N_860);
or U3750 (N_3750,N_1687,N_1875);
and U3751 (N_3751,N_655,N_1164);
nor U3752 (N_3752,N_1160,N_705);
nand U3753 (N_3753,N_1006,N_796);
nor U3754 (N_3754,N_1896,N_1569);
nand U3755 (N_3755,N_192,N_741);
nor U3756 (N_3756,N_641,N_119);
or U3757 (N_3757,N_38,N_748);
nand U3758 (N_3758,N_1352,N_1677);
nor U3759 (N_3759,N_990,N_363);
and U3760 (N_3760,N_1307,N_1713);
nor U3761 (N_3761,N_1203,N_733);
nor U3762 (N_3762,N_1271,N_1448);
nand U3763 (N_3763,N_180,N_1036);
nor U3764 (N_3764,N_1759,N_1541);
nor U3765 (N_3765,N_1536,N_696);
or U3766 (N_3766,N_1817,N_99);
nor U3767 (N_3767,N_281,N_1271);
and U3768 (N_3768,N_880,N_362);
and U3769 (N_3769,N_1357,N_1469);
nand U3770 (N_3770,N_495,N_1860);
or U3771 (N_3771,N_1902,N_674);
xnor U3772 (N_3772,N_810,N_495);
and U3773 (N_3773,N_1146,N_482);
nor U3774 (N_3774,N_196,N_1001);
nor U3775 (N_3775,N_508,N_1692);
and U3776 (N_3776,N_1373,N_1979);
nand U3777 (N_3777,N_897,N_1257);
and U3778 (N_3778,N_525,N_1109);
nand U3779 (N_3779,N_1420,N_607);
nor U3780 (N_3780,N_1062,N_721);
or U3781 (N_3781,N_405,N_241);
nor U3782 (N_3782,N_459,N_1715);
or U3783 (N_3783,N_1459,N_209);
nor U3784 (N_3784,N_52,N_80);
nor U3785 (N_3785,N_1239,N_708);
nor U3786 (N_3786,N_1788,N_1547);
or U3787 (N_3787,N_922,N_1417);
and U3788 (N_3788,N_179,N_1273);
nand U3789 (N_3789,N_1905,N_1683);
nand U3790 (N_3790,N_1608,N_117);
and U3791 (N_3791,N_917,N_1138);
nor U3792 (N_3792,N_1131,N_751);
and U3793 (N_3793,N_1178,N_1908);
nand U3794 (N_3794,N_194,N_1193);
nand U3795 (N_3795,N_171,N_850);
and U3796 (N_3796,N_1576,N_584);
nor U3797 (N_3797,N_1700,N_1926);
or U3798 (N_3798,N_1040,N_1817);
nor U3799 (N_3799,N_1274,N_812);
or U3800 (N_3800,N_1504,N_1855);
nand U3801 (N_3801,N_1895,N_437);
and U3802 (N_3802,N_1315,N_1603);
nor U3803 (N_3803,N_223,N_1264);
nor U3804 (N_3804,N_1442,N_1242);
and U3805 (N_3805,N_348,N_1022);
or U3806 (N_3806,N_1709,N_1814);
nand U3807 (N_3807,N_1331,N_217);
nor U3808 (N_3808,N_681,N_536);
nand U3809 (N_3809,N_1803,N_185);
and U3810 (N_3810,N_881,N_49);
and U3811 (N_3811,N_1657,N_788);
nand U3812 (N_3812,N_1735,N_1184);
or U3813 (N_3813,N_396,N_591);
nor U3814 (N_3814,N_31,N_1947);
nor U3815 (N_3815,N_1855,N_509);
nor U3816 (N_3816,N_1239,N_440);
and U3817 (N_3817,N_885,N_55);
or U3818 (N_3818,N_1037,N_241);
nor U3819 (N_3819,N_1472,N_20);
nor U3820 (N_3820,N_366,N_567);
nor U3821 (N_3821,N_60,N_1417);
nand U3822 (N_3822,N_1474,N_397);
nor U3823 (N_3823,N_1170,N_1618);
or U3824 (N_3824,N_658,N_297);
nor U3825 (N_3825,N_503,N_1442);
nor U3826 (N_3826,N_1610,N_1871);
or U3827 (N_3827,N_1708,N_540);
and U3828 (N_3828,N_1127,N_368);
or U3829 (N_3829,N_227,N_1647);
or U3830 (N_3830,N_1621,N_252);
xor U3831 (N_3831,N_332,N_850);
nor U3832 (N_3832,N_918,N_519);
nand U3833 (N_3833,N_815,N_1531);
and U3834 (N_3834,N_879,N_1706);
nand U3835 (N_3835,N_435,N_427);
and U3836 (N_3836,N_1306,N_182);
nand U3837 (N_3837,N_222,N_1176);
nor U3838 (N_3838,N_1717,N_1847);
nor U3839 (N_3839,N_1591,N_1095);
xnor U3840 (N_3840,N_1068,N_1959);
and U3841 (N_3841,N_1258,N_1460);
nor U3842 (N_3842,N_1279,N_1985);
nand U3843 (N_3843,N_722,N_690);
and U3844 (N_3844,N_200,N_982);
or U3845 (N_3845,N_822,N_274);
nor U3846 (N_3846,N_1958,N_1105);
or U3847 (N_3847,N_614,N_1212);
nor U3848 (N_3848,N_637,N_1695);
and U3849 (N_3849,N_224,N_1583);
nor U3850 (N_3850,N_1609,N_1297);
nand U3851 (N_3851,N_1972,N_890);
and U3852 (N_3852,N_176,N_1311);
and U3853 (N_3853,N_540,N_1852);
nor U3854 (N_3854,N_1289,N_950);
or U3855 (N_3855,N_1450,N_1868);
and U3856 (N_3856,N_1822,N_881);
nor U3857 (N_3857,N_726,N_1890);
and U3858 (N_3858,N_1911,N_580);
and U3859 (N_3859,N_1269,N_863);
or U3860 (N_3860,N_420,N_968);
and U3861 (N_3861,N_806,N_1891);
nand U3862 (N_3862,N_950,N_200);
and U3863 (N_3863,N_1944,N_264);
or U3864 (N_3864,N_1264,N_1703);
and U3865 (N_3865,N_923,N_978);
nor U3866 (N_3866,N_1543,N_1873);
nand U3867 (N_3867,N_1399,N_583);
nand U3868 (N_3868,N_1514,N_448);
nand U3869 (N_3869,N_1160,N_1657);
nor U3870 (N_3870,N_1223,N_703);
nor U3871 (N_3871,N_925,N_168);
nor U3872 (N_3872,N_657,N_646);
nand U3873 (N_3873,N_1905,N_633);
or U3874 (N_3874,N_317,N_1666);
nor U3875 (N_3875,N_51,N_167);
nand U3876 (N_3876,N_1182,N_460);
nand U3877 (N_3877,N_239,N_331);
nor U3878 (N_3878,N_1590,N_1166);
nand U3879 (N_3879,N_1152,N_732);
nor U3880 (N_3880,N_923,N_1986);
xnor U3881 (N_3881,N_1456,N_230);
nand U3882 (N_3882,N_1316,N_945);
nor U3883 (N_3883,N_8,N_1893);
nand U3884 (N_3884,N_1869,N_1604);
xnor U3885 (N_3885,N_656,N_370);
nor U3886 (N_3886,N_1857,N_802);
and U3887 (N_3887,N_1640,N_705);
nor U3888 (N_3888,N_1897,N_1132);
nor U3889 (N_3889,N_776,N_405);
nand U3890 (N_3890,N_516,N_614);
nor U3891 (N_3891,N_447,N_1909);
and U3892 (N_3892,N_248,N_1678);
nor U3893 (N_3893,N_1471,N_1597);
and U3894 (N_3894,N_1036,N_535);
nand U3895 (N_3895,N_217,N_561);
nor U3896 (N_3896,N_1542,N_1782);
nor U3897 (N_3897,N_1566,N_768);
or U3898 (N_3898,N_192,N_1980);
and U3899 (N_3899,N_1566,N_1136);
nand U3900 (N_3900,N_1114,N_1949);
or U3901 (N_3901,N_912,N_602);
nand U3902 (N_3902,N_1602,N_290);
or U3903 (N_3903,N_187,N_1700);
nand U3904 (N_3904,N_85,N_1723);
nor U3905 (N_3905,N_1914,N_1564);
and U3906 (N_3906,N_584,N_948);
nor U3907 (N_3907,N_340,N_1071);
nor U3908 (N_3908,N_1431,N_654);
and U3909 (N_3909,N_1280,N_766);
nor U3910 (N_3910,N_250,N_544);
or U3911 (N_3911,N_1002,N_750);
and U3912 (N_3912,N_936,N_923);
nand U3913 (N_3913,N_112,N_1424);
nor U3914 (N_3914,N_1531,N_806);
xnor U3915 (N_3915,N_1509,N_935);
and U3916 (N_3916,N_945,N_720);
nand U3917 (N_3917,N_211,N_1712);
or U3918 (N_3918,N_1911,N_1976);
nand U3919 (N_3919,N_1136,N_494);
or U3920 (N_3920,N_1027,N_675);
nor U3921 (N_3921,N_696,N_1717);
and U3922 (N_3922,N_865,N_1754);
nand U3923 (N_3923,N_1242,N_1434);
or U3924 (N_3924,N_364,N_635);
nand U3925 (N_3925,N_1603,N_1998);
or U3926 (N_3926,N_1434,N_1464);
or U3927 (N_3927,N_1067,N_723);
or U3928 (N_3928,N_1596,N_821);
nor U3929 (N_3929,N_1955,N_594);
nand U3930 (N_3930,N_788,N_422);
and U3931 (N_3931,N_1276,N_1125);
nor U3932 (N_3932,N_596,N_1334);
and U3933 (N_3933,N_992,N_50);
or U3934 (N_3934,N_1749,N_697);
and U3935 (N_3935,N_1834,N_1511);
nor U3936 (N_3936,N_219,N_447);
or U3937 (N_3937,N_1186,N_27);
nor U3938 (N_3938,N_897,N_1994);
or U3939 (N_3939,N_639,N_34);
and U3940 (N_3940,N_1322,N_1040);
or U3941 (N_3941,N_816,N_571);
nor U3942 (N_3942,N_518,N_866);
or U3943 (N_3943,N_837,N_500);
and U3944 (N_3944,N_985,N_1255);
nor U3945 (N_3945,N_822,N_1434);
nor U3946 (N_3946,N_522,N_808);
or U3947 (N_3947,N_788,N_1507);
nand U3948 (N_3948,N_1320,N_1584);
nand U3949 (N_3949,N_1391,N_498);
nand U3950 (N_3950,N_1492,N_1336);
nand U3951 (N_3951,N_1961,N_592);
nand U3952 (N_3952,N_1743,N_1075);
xor U3953 (N_3953,N_1544,N_408);
or U3954 (N_3954,N_1089,N_1452);
xnor U3955 (N_3955,N_723,N_240);
nor U3956 (N_3956,N_1626,N_1928);
or U3957 (N_3957,N_1908,N_131);
nor U3958 (N_3958,N_588,N_1313);
nand U3959 (N_3959,N_125,N_1934);
nand U3960 (N_3960,N_1835,N_1384);
nand U3961 (N_3961,N_1500,N_214);
or U3962 (N_3962,N_756,N_1622);
or U3963 (N_3963,N_326,N_1112);
and U3964 (N_3964,N_1463,N_301);
nor U3965 (N_3965,N_1232,N_1559);
or U3966 (N_3966,N_1205,N_161);
nand U3967 (N_3967,N_940,N_352);
and U3968 (N_3968,N_562,N_1146);
or U3969 (N_3969,N_730,N_1739);
or U3970 (N_3970,N_1121,N_1852);
and U3971 (N_3971,N_1634,N_804);
nand U3972 (N_3972,N_911,N_1439);
and U3973 (N_3973,N_1842,N_1612);
or U3974 (N_3974,N_1888,N_1068);
nand U3975 (N_3975,N_1483,N_1780);
nand U3976 (N_3976,N_1440,N_327);
xnor U3977 (N_3977,N_260,N_1294);
or U3978 (N_3978,N_501,N_1912);
nor U3979 (N_3979,N_769,N_837);
nor U3980 (N_3980,N_669,N_1134);
nand U3981 (N_3981,N_309,N_1434);
nand U3982 (N_3982,N_857,N_961);
and U3983 (N_3983,N_997,N_198);
nand U3984 (N_3984,N_740,N_1676);
nor U3985 (N_3985,N_1295,N_1827);
and U3986 (N_3986,N_179,N_549);
nand U3987 (N_3987,N_1400,N_1602);
nand U3988 (N_3988,N_667,N_390);
and U3989 (N_3989,N_1670,N_1263);
or U3990 (N_3990,N_1466,N_1878);
or U3991 (N_3991,N_1921,N_982);
nor U3992 (N_3992,N_1095,N_209);
nor U3993 (N_3993,N_1439,N_1329);
or U3994 (N_3994,N_269,N_1376);
nand U3995 (N_3995,N_1772,N_940);
or U3996 (N_3996,N_474,N_1328);
nor U3997 (N_3997,N_1708,N_1148);
nand U3998 (N_3998,N_364,N_1573);
or U3999 (N_3999,N_304,N_236);
nor U4000 (N_4000,N_2097,N_2943);
nor U4001 (N_4001,N_3452,N_2286);
and U4002 (N_4002,N_2839,N_3979);
or U4003 (N_4003,N_2612,N_3212);
or U4004 (N_4004,N_3889,N_3069);
or U4005 (N_4005,N_3735,N_2776);
nand U4006 (N_4006,N_2379,N_2605);
and U4007 (N_4007,N_3969,N_3325);
nor U4008 (N_4008,N_2210,N_3068);
and U4009 (N_4009,N_2534,N_2955);
nor U4010 (N_4010,N_3010,N_3363);
nor U4011 (N_4011,N_3284,N_3082);
nor U4012 (N_4012,N_2141,N_2034);
and U4013 (N_4013,N_2278,N_3860);
nor U4014 (N_4014,N_3977,N_2136);
nand U4015 (N_4015,N_3169,N_3794);
nor U4016 (N_4016,N_2145,N_2731);
nor U4017 (N_4017,N_3438,N_3317);
or U4018 (N_4018,N_3527,N_3358);
nor U4019 (N_4019,N_3526,N_2398);
or U4020 (N_4020,N_2639,N_3428);
and U4021 (N_4021,N_2434,N_2303);
or U4022 (N_4022,N_2483,N_3901);
nor U4023 (N_4023,N_2827,N_2894);
nor U4024 (N_4024,N_2608,N_2510);
or U4025 (N_4025,N_3194,N_3795);
and U4026 (N_4026,N_3639,N_2227);
nand U4027 (N_4027,N_3046,N_2637);
or U4028 (N_4028,N_3830,N_3383);
nand U4029 (N_4029,N_2522,N_3876);
nand U4030 (N_4030,N_2897,N_3832);
nor U4031 (N_4031,N_2266,N_3401);
or U4032 (N_4032,N_2563,N_3618);
and U4033 (N_4033,N_2866,N_2087);
or U4034 (N_4034,N_2855,N_3851);
and U4035 (N_4035,N_2797,N_3582);
or U4036 (N_4036,N_2710,N_3017);
nor U4037 (N_4037,N_2626,N_2718);
nor U4038 (N_4038,N_2935,N_2372);
nand U4039 (N_4039,N_3297,N_3481);
nor U4040 (N_4040,N_2105,N_2255);
nor U4041 (N_4041,N_3610,N_2983);
and U4042 (N_4042,N_2975,N_3588);
and U4043 (N_4043,N_2016,N_2144);
nand U4044 (N_4044,N_3395,N_3932);
nand U4045 (N_4045,N_2519,N_2734);
or U4046 (N_4046,N_2913,N_2359);
and U4047 (N_4047,N_2625,N_3165);
nor U4048 (N_4048,N_2369,N_2505);
and U4049 (N_4049,N_2442,N_3965);
nor U4050 (N_4050,N_2553,N_2331);
and U4051 (N_4051,N_3692,N_3565);
or U4052 (N_4052,N_2100,N_3559);
or U4053 (N_4053,N_2853,N_2095);
nor U4054 (N_4054,N_2856,N_2854);
nand U4055 (N_4055,N_3249,N_3463);
nor U4056 (N_4056,N_2769,N_3804);
and U4057 (N_4057,N_3403,N_2516);
and U4058 (N_4058,N_3024,N_2116);
nand U4059 (N_4059,N_3602,N_3035);
nor U4060 (N_4060,N_2479,N_3285);
or U4061 (N_4061,N_2989,N_2251);
and U4062 (N_4062,N_2150,N_2705);
nand U4063 (N_4063,N_2480,N_3528);
nor U4064 (N_4064,N_2934,N_2536);
and U4065 (N_4065,N_3311,N_3086);
xnor U4066 (N_4066,N_2777,N_2887);
nor U4067 (N_4067,N_2566,N_3942);
or U4068 (N_4068,N_2584,N_2167);
and U4069 (N_4069,N_2194,N_2630);
nor U4070 (N_4070,N_2977,N_3567);
or U4071 (N_4071,N_3562,N_2944);
or U4072 (N_4072,N_3608,N_3073);
nor U4073 (N_4073,N_3952,N_3020);
nor U4074 (N_4074,N_2492,N_2383);
nand U4075 (N_4075,N_2312,N_3984);
and U4076 (N_4076,N_2545,N_2321);
nor U4077 (N_4077,N_3672,N_2790);
and U4078 (N_4078,N_3259,N_3546);
or U4079 (N_4079,N_3126,N_2015);
nor U4080 (N_4080,N_3990,N_3516);
nor U4081 (N_4081,N_3025,N_3778);
nor U4082 (N_4082,N_2692,N_3552);
or U4083 (N_4083,N_3278,N_3710);
and U4084 (N_4084,N_2476,N_2815);
and U4085 (N_4085,N_3571,N_3508);
nand U4086 (N_4086,N_2942,N_3486);
nor U4087 (N_4087,N_3127,N_3006);
nor U4088 (N_4088,N_2698,N_3023);
nand U4089 (N_4089,N_3504,N_3107);
nand U4090 (N_4090,N_2757,N_2783);
and U4091 (N_4091,N_2949,N_3584);
or U4092 (N_4092,N_2773,N_3738);
nor U4093 (N_4093,N_2373,N_2513);
or U4094 (N_4094,N_2403,N_2669);
and U4095 (N_4095,N_2080,N_3364);
and U4096 (N_4096,N_3682,N_3339);
nor U4097 (N_4097,N_2471,N_2067);
or U4098 (N_4098,N_2952,N_2524);
or U4099 (N_4099,N_3004,N_3427);
or U4100 (N_4100,N_3730,N_2759);
and U4101 (N_4101,N_3976,N_2556);
nor U4102 (N_4102,N_3789,N_2904);
nand U4103 (N_4103,N_2154,N_2305);
nand U4104 (N_4104,N_2209,N_2488);
nand U4105 (N_4105,N_3464,N_2157);
nor U4106 (N_4106,N_2835,N_2579);
nor U4107 (N_4107,N_2207,N_3859);
and U4108 (N_4108,N_3695,N_3919);
or U4109 (N_4109,N_2039,N_2966);
nand U4110 (N_4110,N_2928,N_2939);
or U4111 (N_4111,N_2256,N_2829);
and U4112 (N_4112,N_2262,N_3717);
and U4113 (N_4113,N_3589,N_2561);
nand U4114 (N_4114,N_3656,N_3091);
and U4115 (N_4115,N_3606,N_2618);
or U4116 (N_4116,N_2348,N_2414);
and U4117 (N_4117,N_2073,N_2253);
nor U4118 (N_4118,N_2875,N_3745);
nand U4119 (N_4119,N_2281,N_3170);
nand U4120 (N_4120,N_2493,N_2697);
nand U4121 (N_4121,N_2911,N_3372);
and U4122 (N_4122,N_2104,N_3579);
or U4123 (N_4123,N_3908,N_3479);
or U4124 (N_4124,N_2115,N_3030);
nand U4125 (N_4125,N_3515,N_2551);
and U4126 (N_4126,N_3113,N_3449);
or U4127 (N_4127,N_3764,N_2784);
nand U4128 (N_4128,N_3232,N_3742);
and U4129 (N_4129,N_2018,N_3114);
and U4130 (N_4130,N_3135,N_3043);
nor U4131 (N_4131,N_3946,N_2463);
and U4132 (N_4132,N_3629,N_3718);
nand U4133 (N_4133,N_3061,N_3992);
and U4134 (N_4134,N_2717,N_2086);
and U4135 (N_4135,N_3276,N_2751);
nor U4136 (N_4136,N_3609,N_2441);
or U4137 (N_4137,N_2003,N_2313);
or U4138 (N_4138,N_3262,N_2109);
nand U4139 (N_4139,N_3802,N_3161);
nor U4140 (N_4140,N_3723,N_3757);
nand U4141 (N_4141,N_3586,N_2345);
nand U4142 (N_4142,N_3986,N_2602);
nor U4143 (N_4143,N_2182,N_2096);
and U4144 (N_4144,N_2661,N_2946);
and U4145 (N_4145,N_3911,N_3595);
nor U4146 (N_4146,N_3484,N_2867);
or U4147 (N_4147,N_2238,N_3172);
or U4148 (N_4148,N_2953,N_3236);
nand U4149 (N_4149,N_3825,N_2469);
and U4150 (N_4150,N_3497,N_3774);
and U4151 (N_4151,N_2766,N_3845);
or U4152 (N_4152,N_3168,N_3597);
and U4153 (N_4153,N_2660,N_3386);
and U4154 (N_4154,N_3580,N_2526);
and U4155 (N_4155,N_2040,N_2288);
nor U4156 (N_4156,N_3347,N_2284);
and U4157 (N_4157,N_3775,N_2054);
nand U4158 (N_4158,N_3222,N_3868);
and U4159 (N_4159,N_3177,N_2409);
nor U4160 (N_4160,N_3028,N_2482);
and U4161 (N_4161,N_3088,N_3381);
or U4162 (N_4162,N_3397,N_3419);
nand U4163 (N_4163,N_2060,N_2754);
nand U4164 (N_4164,N_3097,N_2367);
or U4165 (N_4165,N_2357,N_2009);
nand U4166 (N_4166,N_2870,N_2410);
nand U4167 (N_4167,N_2258,N_2417);
nor U4168 (N_4168,N_3233,N_2174);
nand U4169 (N_4169,N_2301,N_2613);
nor U4170 (N_4170,N_3677,N_2007);
nand U4171 (N_4171,N_2057,N_3539);
and U4172 (N_4172,N_3944,N_2749);
nor U4173 (N_4173,N_2923,N_2098);
or U4174 (N_4174,N_2549,N_2416);
and U4175 (N_4175,N_3807,N_2239);
nand U4176 (N_4176,N_3400,N_3142);
nand U4177 (N_4177,N_2791,N_2930);
nand U4178 (N_4178,N_3517,N_3708);
nand U4179 (N_4179,N_2232,N_2577);
or U4180 (N_4180,N_3153,N_3784);
and U4181 (N_4181,N_3534,N_3290);
and U4182 (N_4182,N_3267,N_3931);
nor U4183 (N_4183,N_3008,N_2940);
or U4184 (N_4184,N_2223,N_3596);
nand U4185 (N_4185,N_3664,N_2272);
nand U4186 (N_4186,N_2686,N_3129);
and U4187 (N_4187,N_2092,N_3522);
or U4188 (N_4188,N_2428,N_2846);
or U4189 (N_4189,N_2511,N_2828);
and U4190 (N_4190,N_2302,N_3027);
and U4191 (N_4191,N_2364,N_3836);
and U4192 (N_4192,N_3987,N_3365);
and U4193 (N_4193,N_3195,N_3281);
nor U4194 (N_4194,N_2544,N_2518);
nand U4195 (N_4195,N_3145,N_2451);
nand U4196 (N_4196,N_2538,N_2882);
or U4197 (N_4197,N_3870,N_2076);
and U4198 (N_4198,N_3144,N_2599);
and U4199 (N_4199,N_2653,N_3346);
nor U4200 (N_4200,N_3079,N_3343);
nand U4201 (N_4201,N_2622,N_3150);
nand U4202 (N_4202,N_2937,N_2183);
nand U4203 (N_4203,N_3092,N_2520);
and U4204 (N_4204,N_3143,N_2557);
and U4205 (N_4205,N_2716,N_3301);
nand U4206 (N_4206,N_2999,N_3242);
or U4207 (N_4207,N_2090,N_3408);
nand U4208 (N_4208,N_2822,N_2899);
nor U4209 (N_4209,N_2184,N_2103);
and U4210 (N_4210,N_2346,N_3714);
or U4211 (N_4211,N_2322,N_3304);
or U4212 (N_4212,N_3506,N_3551);
nand U4213 (N_4213,N_2800,N_3728);
or U4214 (N_4214,N_3881,N_3048);
nor U4215 (N_4215,N_2648,N_2261);
or U4216 (N_4216,N_2725,N_3287);
or U4217 (N_4217,N_3469,N_2964);
and U4218 (N_4218,N_3635,N_2876);
and U4219 (N_4219,N_3754,N_2069);
and U4220 (N_4220,N_3805,N_3821);
nor U4221 (N_4221,N_3455,N_2594);
and U4222 (N_4222,N_2267,N_2588);
nor U4223 (N_4223,N_3186,N_2699);
or U4224 (N_4224,N_3159,N_3075);
nor U4225 (N_4225,N_2743,N_3003);
nand U4226 (N_4226,N_3070,N_3737);
nand U4227 (N_4227,N_2327,N_3548);
and U4228 (N_4228,N_3149,N_2657);
or U4229 (N_4229,N_2289,N_2555);
or U4230 (N_4230,N_2126,N_2874);
or U4231 (N_4231,N_3255,N_3724);
nand U4232 (N_4232,N_2037,N_2580);
or U4233 (N_4233,N_3943,N_2540);
xnor U4234 (N_4234,N_2914,N_3308);
nor U4235 (N_4235,N_3840,N_3575);
and U4236 (N_4236,N_2593,N_2093);
and U4237 (N_4237,N_3101,N_2504);
nand U4238 (N_4238,N_3827,N_2912);
and U4239 (N_4239,N_3537,N_2195);
and U4240 (N_4240,N_3362,N_3653);
and U4241 (N_4241,N_3513,N_2459);
nor U4242 (N_4242,N_3445,N_3012);
and U4243 (N_4243,N_2980,N_3797);
or U4244 (N_4244,N_3252,N_2454);
nor U4245 (N_4245,N_3507,N_2547);
and U4246 (N_4246,N_2742,N_3733);
nor U4247 (N_4247,N_2125,N_2212);
nand U4248 (N_4248,N_3855,N_3566);
nor U4249 (N_4249,N_2811,N_3077);
nor U4250 (N_4250,N_2401,N_2623);
nand U4251 (N_4251,N_3060,N_2640);
or U4252 (N_4252,N_2431,N_2606);
and U4253 (N_4253,N_2241,N_2748);
and U4254 (N_4254,N_2390,N_2248);
and U4255 (N_4255,N_2527,N_3390);
nand U4256 (N_4256,N_2885,N_3247);
or U4257 (N_4257,N_2224,N_2172);
and U4258 (N_4258,N_3426,N_2666);
nand U4259 (N_4259,N_3510,N_3810);
nor U4260 (N_4260,N_2269,N_2539);
or U4261 (N_4261,N_3839,N_2252);
nand U4262 (N_4262,N_2211,N_2685);
and U4263 (N_4263,N_2512,N_2064);
and U4264 (N_4264,N_2767,N_2896);
or U4265 (N_4265,N_2466,N_2772);
and U4266 (N_4266,N_2906,N_2208);
nand U4267 (N_4267,N_2575,N_2435);
nor U4268 (N_4268,N_3394,N_3666);
or U4269 (N_4269,N_2392,N_3348);
and U4270 (N_4270,N_2189,N_3747);
nand U4271 (N_4271,N_3019,N_2316);
nand U4272 (N_4272,N_2014,N_3554);
nand U4273 (N_4273,N_2521,N_3156);
nor U4274 (N_4274,N_3047,N_3116);
or U4275 (N_4275,N_3109,N_2049);
nor U4276 (N_4276,N_3644,N_3366);
and U4277 (N_4277,N_3229,N_2166);
and U4278 (N_4278,N_3310,N_3322);
or U4279 (N_4279,N_2865,N_3475);
nand U4280 (N_4280,N_3632,N_3736);
nand U4281 (N_4281,N_3995,N_2532);
and U4282 (N_4282,N_2795,N_3154);
and U4283 (N_4283,N_2981,N_2857);
or U4284 (N_4284,N_2333,N_3342);
nor U4285 (N_4285,N_3897,N_2655);
nand U4286 (N_4286,N_2399,N_2374);
nand U4287 (N_4287,N_2407,N_3947);
and U4288 (N_4288,N_3907,N_3514);
nor U4289 (N_4289,N_3961,N_3040);
or U4290 (N_4290,N_2834,N_3975);
or U4291 (N_4291,N_2196,N_2782);
or U4292 (N_4292,N_2436,N_3558);
or U4293 (N_4293,N_2432,N_2475);
and U4294 (N_4294,N_2050,N_2794);
and U4295 (N_4295,N_2738,N_3788);
and U4296 (N_4296,N_3219,N_3543);
nand U4297 (N_4297,N_2775,N_3146);
nor U4298 (N_4298,N_3227,N_3835);
or U4299 (N_4299,N_2733,N_2378);
or U4300 (N_4300,N_2338,N_3076);
or U4301 (N_4301,N_3329,N_2259);
nor U4302 (N_4302,N_2677,N_2156);
nand U4303 (N_4303,N_2153,N_2437);
and U4304 (N_4304,N_2192,N_2525);
or U4305 (N_4305,N_3124,N_2936);
and U4306 (N_4306,N_2112,N_2106);
and U4307 (N_4307,N_2271,N_3895);
or U4308 (N_4308,N_3903,N_3785);
nand U4309 (N_4309,N_3972,N_2631);
or U4310 (N_4310,N_2761,N_3703);
or U4311 (N_4311,N_3509,N_2927);
and U4312 (N_4312,N_2567,N_3341);
and U4313 (N_4313,N_3777,N_2349);
nor U4314 (N_4314,N_2426,N_3521);
nor U4315 (N_4315,N_3257,N_2375);
and U4316 (N_4316,N_2721,N_2978);
nand U4317 (N_4317,N_2832,N_3388);
nor U4318 (N_4318,N_2696,N_2358);
and U4319 (N_4319,N_2231,N_3123);
and U4320 (N_4320,N_2394,N_2276);
nand U4321 (N_4321,N_3791,N_3598);
nor U4322 (N_4322,N_2307,N_3251);
nand U4323 (N_4323,N_3237,N_3239);
and U4324 (N_4324,N_2711,N_3748);
or U4325 (N_4325,N_2879,N_3253);
or U4326 (N_4326,N_2135,N_2214);
and U4327 (N_4327,N_2177,N_2023);
or U4328 (N_4328,N_2113,N_3857);
nand U4329 (N_4329,N_2508,N_2658);
and U4330 (N_4330,N_2117,N_3679);
or U4331 (N_4331,N_2051,N_3300);
and U4332 (N_4332,N_2031,N_2771);
and U4333 (N_4333,N_2796,N_3496);
nor U4334 (N_4334,N_2781,N_2991);
nor U4335 (N_4335,N_3781,N_3241);
or U4336 (N_4336,N_3918,N_2993);
nand U4337 (N_4337,N_2148,N_3104);
or U4338 (N_4338,N_3448,N_3711);
and U4339 (N_4339,N_2821,N_2035);
and U4340 (N_4340,N_3410,N_3822);
nor U4341 (N_4341,N_2164,N_3636);
or U4342 (N_4342,N_2306,N_2809);
or U4343 (N_4343,N_3258,N_3938);
nor U4344 (N_4344,N_3535,N_3456);
nor U4345 (N_4345,N_2205,N_2165);
and U4346 (N_4346,N_3122,N_3207);
nand U4347 (N_4347,N_3896,N_2816);
or U4348 (N_4348,N_3225,N_3953);
nand U4349 (N_4349,N_3190,N_3056);
and U4350 (N_4350,N_2843,N_2503);
or U4351 (N_4351,N_3704,N_3963);
nor U4352 (N_4352,N_3356,N_2714);
nor U4353 (N_4353,N_3051,N_3874);
nand U4354 (N_4354,N_3327,N_3293);
nand U4355 (N_4355,N_3796,N_2474);
nor U4356 (N_4356,N_3478,N_3299);
nand U4357 (N_4357,N_2689,N_3181);
and U4358 (N_4358,N_3640,N_2558);
and U4359 (N_4359,N_3015,N_3274);
nor U4360 (N_4360,N_3768,N_2737);
and U4361 (N_4361,N_3173,N_2443);
or U4362 (N_4362,N_2900,N_2541);
nand U4363 (N_4363,N_2181,N_3487);
nand U4364 (N_4364,N_2491,N_3180);
nor U4365 (N_4365,N_3049,N_3062);
and U4366 (N_4366,N_2802,N_3275);
nand U4367 (N_4367,N_2114,N_2941);
and U4368 (N_4368,N_2121,N_3420);
nor U4369 (N_4369,N_3996,N_3915);
and U4370 (N_4370,N_2600,N_3937);
or U4371 (N_4371,N_2022,N_3661);
and U4372 (N_4372,N_3729,N_2514);
nor U4373 (N_4373,N_2188,N_2901);
or U4374 (N_4374,N_2812,N_2841);
nand U4375 (N_4375,N_2011,N_3380);
or U4376 (N_4376,N_3862,N_2645);
or U4377 (N_4377,N_2158,N_3220);
and U4378 (N_4378,N_3888,N_3941);
nor U4379 (N_4379,N_2310,N_2614);
or U4380 (N_4380,N_3950,N_3871);
nor U4381 (N_4381,N_2235,N_3741);
nor U4382 (N_4382,N_3503,N_2485);
xor U4383 (N_4383,N_2481,N_2386);
or U4384 (N_4384,N_3430,N_3044);
or U4385 (N_4385,N_2895,N_2120);
nor U4386 (N_4386,N_3688,N_3878);
nand U4387 (N_4387,N_2667,N_2452);
nor U4388 (N_4388,N_2762,N_2176);
or U4389 (N_4389,N_2308,N_2130);
and U4390 (N_4390,N_2074,N_3282);
or U4391 (N_4391,N_3964,N_2543);
or U4392 (N_4392,N_3384,N_2633);
nor U4393 (N_4393,N_2945,N_2724);
or U4394 (N_4394,N_3819,N_3319);
nor U4395 (N_4395,N_2651,N_2969);
or U4396 (N_4396,N_2339,N_2601);
nor U4397 (N_4397,N_2799,N_2293);
nor U4398 (N_4398,N_3887,N_3226);
nand U4399 (N_4399,N_2573,N_3645);
nor U4400 (N_4400,N_2460,N_3432);
or U4401 (N_4401,N_3725,N_2328);
nor U4402 (N_4402,N_3041,N_2755);
or U4403 (N_4403,N_2610,N_3106);
nand U4404 (N_4404,N_3910,N_2420);
or U4405 (N_4405,N_2218,N_3934);
nand U4406 (N_4406,N_3641,N_2082);
nor U4407 (N_4407,N_2429,N_2706);
nand U4408 (N_4408,N_2068,N_3817);
nor U4409 (N_4409,N_2823,N_3560);
or U4410 (N_4410,N_3812,N_3250);
or U4411 (N_4411,N_2909,N_2179);
nor U4412 (N_4412,N_3296,N_3416);
nand U4413 (N_4413,N_3681,N_2758);
or U4414 (N_4414,N_3800,N_3529);
nor U4415 (N_4415,N_3201,N_3425);
and U4416 (N_4416,N_2851,N_2006);
nand U4417 (N_4417,N_3011,N_2529);
nor U4418 (N_4418,N_2788,N_3734);
and U4419 (N_4419,N_3368,N_2350);
nand U4420 (N_4420,N_3096,N_2884);
nand U4421 (N_4421,N_2523,N_2384);
nand U4422 (N_4422,N_3002,N_3962);
nand U4423 (N_4423,N_2243,N_3863);
nor U4424 (N_4424,N_3370,N_3739);
nand U4425 (N_4425,N_2285,N_3891);
nand U4426 (N_4426,N_3525,N_2604);
nand U4427 (N_4427,N_3532,N_3906);
nor U4428 (N_4428,N_2101,N_3099);
or U4429 (N_4429,N_3133,N_2917);
nand U4430 (N_4430,N_3080,N_2583);
or U4431 (N_4431,N_2304,N_2956);
or U4432 (N_4432,N_2961,N_2680);
nor U4433 (N_4433,N_3763,N_2032);
and U4434 (N_4434,N_2603,N_2779);
nand U4435 (N_4435,N_2260,N_2656);
or U4436 (N_4436,N_2628,N_2395);
or U4437 (N_4437,N_2217,N_3790);
nand U4438 (N_4438,N_2270,N_2642);
nand U4439 (N_4439,N_2780,N_3877);
or U4440 (N_4440,N_3451,N_3094);
or U4441 (N_4441,N_3928,N_3131);
or U4442 (N_4442,N_2702,N_2905);
nand U4443 (N_4443,N_3228,N_2311);
and U4444 (N_4444,N_2550,N_2299);
nor U4445 (N_4445,N_2746,N_3273);
or U4446 (N_4446,N_2219,N_3850);
nor U4447 (N_4447,N_2155,N_3326);
nand U4448 (N_4448,N_2146,N_3671);
nand U4449 (N_4449,N_3604,N_3336);
or U4450 (N_4450,N_3031,N_3470);
nand U4451 (N_4451,N_3187,N_3780);
and U4452 (N_4452,N_3178,N_2110);
and U4453 (N_4453,N_3890,N_2672);
or U4454 (N_4454,N_2915,N_3647);
or U4455 (N_4455,N_2048,N_2447);
nor U4456 (N_4456,N_3377,N_3089);
nand U4457 (N_4457,N_3176,N_3309);
nand U4458 (N_4458,N_3256,N_3511);
or U4459 (N_4459,N_3519,N_2967);
and U4460 (N_4460,N_3691,N_3667);
nand U4461 (N_4461,N_3930,N_3939);
nor U4462 (N_4462,N_2903,N_2959);
nor U4463 (N_4463,N_3268,N_2764);
nand U4464 (N_4464,N_3956,N_2996);
and U4465 (N_4465,N_2674,N_2620);
nor U4466 (N_4466,N_2134,N_3715);
and U4467 (N_4467,N_2152,N_3686);
nor U4468 (N_4468,N_3271,N_2741);
or U4469 (N_4469,N_3553,N_3151);
nand U4470 (N_4470,N_3899,N_2650);
nor U4471 (N_4471,N_3501,N_2000);
and U4472 (N_4472,N_2890,N_3196);
nand U4473 (N_4473,N_3743,N_2198);
and U4474 (N_4474,N_2458,N_2619);
nand U4475 (N_4475,N_3429,N_2237);
nand U4476 (N_4476,N_3373,N_2203);
or U4477 (N_4477,N_3406,N_3826);
nand U4478 (N_4478,N_2888,N_2472);
nand U4479 (N_4479,N_2542,N_3959);
nor U4480 (N_4480,N_3261,N_2891);
nand U4481 (N_4481,N_3141,N_2922);
nor U4482 (N_4482,N_2047,N_2139);
or U4483 (N_4483,N_3994,N_3098);
nand U4484 (N_4484,N_3536,N_2222);
and U4485 (N_4485,N_2634,N_3422);
or U4486 (N_4486,N_3767,N_2963);
nor U4487 (N_4487,N_2213,N_2353);
nor U4488 (N_4488,N_3759,N_3318);
nor U4489 (N_4489,N_2277,N_2785);
nand U4490 (N_4490,N_2043,N_3678);
or U4491 (N_4491,N_3643,N_3633);
nand U4492 (N_4492,N_3164,N_2400);
or U4493 (N_4493,N_3337,N_3731);
or U4494 (N_4494,N_3920,N_3622);
or U4495 (N_4495,N_3152,N_3245);
xor U4496 (N_4496,N_3960,N_2046);
or U4497 (N_4497,N_3018,N_3493);
nand U4498 (N_4498,N_3974,N_3833);
or U4499 (N_4499,N_3696,N_3034);
nand U4500 (N_4500,N_2202,N_3084);
nand U4501 (N_4501,N_2319,N_2484);
nand U4502 (N_4502,N_2065,N_2282);
or U4503 (N_4503,N_2701,N_3295);
and U4504 (N_4504,N_3058,N_2257);
and U4505 (N_4505,N_2703,N_2127);
nor U4506 (N_4506,N_2030,N_3846);
nand U4507 (N_4507,N_2137,N_3087);
and U4508 (N_4508,N_3443,N_2753);
or U4509 (N_4509,N_3824,N_3055);
and U4510 (N_4510,N_3576,N_3147);
and U4511 (N_4511,N_3541,N_2986);
nor U4512 (N_4512,N_3700,N_3533);
nor U4513 (N_4513,N_2582,N_2659);
and U4514 (N_4514,N_3856,N_3036);
nand U4515 (N_4515,N_3721,N_2792);
and U4516 (N_4516,N_3680,N_3663);
nor U4517 (N_4517,N_2236,N_3892);
nor U4518 (N_4518,N_3162,N_2820);
and U4519 (N_4519,N_3866,N_2789);
and U4520 (N_4520,N_3673,N_2671);
and U4521 (N_4521,N_3078,N_2836);
or U4522 (N_4522,N_2948,N_3627);
nor U4523 (N_4523,N_2842,N_2433);
or U4524 (N_4524,N_3264,N_2111);
nand U4525 (N_4525,N_2535,N_3900);
nand U4526 (N_4526,N_2726,N_3770);
nor U4527 (N_4527,N_2586,N_3185);
and U4528 (N_4528,N_2161,N_3205);
or U4529 (N_4529,N_2123,N_3894);
or U4530 (N_4530,N_3454,N_3561);
nand U4531 (N_4531,N_2574,N_2768);
nor U4532 (N_4532,N_2838,N_3307);
or U4533 (N_4533,N_2760,N_2185);
nor U4534 (N_4534,N_2024,N_2814);
nor U4535 (N_4535,N_2868,N_3477);
or U4536 (N_4536,N_2552,N_3110);
and U4537 (N_4537,N_3375,N_3413);
nand U4538 (N_4538,N_3848,N_3354);
nor U4539 (N_4539,N_3948,N_3631);
nor U4540 (N_4540,N_3459,N_3235);
and U4541 (N_4541,N_2062,N_3393);
and U4542 (N_4542,N_2347,N_3806);
and U4543 (N_4543,N_2793,N_2872);
nor U4544 (N_4544,N_3726,N_2490);
nand U4545 (N_4545,N_2770,N_3001);
and U4546 (N_4546,N_3230,N_2254);
nand U4547 (N_4547,N_2860,N_3709);
nand U4548 (N_4548,N_2193,N_2691);
or U4549 (N_4549,N_2094,N_2931);
nand U4550 (N_4550,N_3732,N_3240);
nand U4551 (N_4551,N_2440,N_3634);
nand U4552 (N_4552,N_2831,N_2589);
nand U4553 (N_4553,N_3139,N_3340);
and U4554 (N_4554,N_3512,N_3217);
nor U4555 (N_4555,N_3547,N_3657);
nor U4556 (N_4556,N_3376,N_3988);
nand U4557 (N_4557,N_2226,N_3292);
xor U4558 (N_4558,N_2361,N_3861);
nand U4559 (N_4559,N_3136,N_2422);
nor U4560 (N_4560,N_2974,N_3216);
nand U4561 (N_4561,N_3587,N_3902);
nor U4562 (N_4562,N_3072,N_2204);
nand U4563 (N_4563,N_3214,N_3756);
nand U4564 (N_4564,N_2273,N_2715);
or U4565 (N_4565,N_3621,N_2225);
nand U4566 (N_4566,N_2881,N_3065);
and U4567 (N_4567,N_2690,N_2938);
or U4568 (N_4568,N_2274,N_3753);
nor U4569 (N_4569,N_2119,N_3210);
or U4570 (N_4570,N_2537,N_2376);
or U4571 (N_4571,N_2590,N_3494);
or U4572 (N_4572,N_3021,N_2979);
nor U4573 (N_4573,N_3603,N_3776);
and U4574 (N_4574,N_3014,N_3660);
nor U4575 (N_4575,N_2929,N_3490);
nor U4576 (N_4576,N_3200,N_3349);
nor U4577 (N_4577,N_3614,N_2334);
and U4578 (N_4578,N_2804,N_3052);
nand U4579 (N_4579,N_3699,N_3531);
nor U4580 (N_4580,N_2958,N_3005);
and U4581 (N_4581,N_3916,N_3769);
and U4582 (N_4582,N_3361,N_3707);
or U4583 (N_4583,N_3244,N_2438);
nor U4584 (N_4584,N_3545,N_2886);
and U4585 (N_4585,N_3137,N_2533);
nor U4586 (N_4586,N_2180,N_2995);
nor U4587 (N_4587,N_2215,N_2708);
and U4588 (N_4588,N_3303,N_2187);
nor U4589 (N_4589,N_2300,N_3765);
nor U4590 (N_4590,N_2078,N_2041);
or U4591 (N_4591,N_2246,N_3352);
nand U4592 (N_4592,N_3211,N_3458);
nor U4593 (N_4593,N_2406,N_2002);
or U4594 (N_4594,N_3179,N_2233);
nor U4595 (N_4595,N_3409,N_2221);
nor U4596 (N_4596,N_3782,N_3059);
nor U4597 (N_4597,N_3404,N_2220);
and U4598 (N_4598,N_3243,N_3460);
nor U4599 (N_4599,N_3993,N_2240);
and U4600 (N_4600,N_3933,N_2283);
nand U4601 (N_4601,N_3439,N_2295);
and U4602 (N_4602,N_2486,N_2752);
or U4603 (N_4603,N_3331,N_3359);
nand U4604 (N_4604,N_3157,N_3809);
nor U4605 (N_4605,N_3392,N_2982);
and U4606 (N_4606,N_3298,N_2200);
or U4607 (N_4607,N_2419,N_3755);
or U4608 (N_4608,N_2990,N_2858);
and U4609 (N_4609,N_2391,N_3029);
and U4610 (N_4610,N_2728,N_2170);
and U4611 (N_4611,N_2918,N_3045);
xnor U4612 (N_4612,N_3160,N_3476);
nor U4613 (N_4613,N_3951,N_3389);
and U4614 (N_4614,N_2739,N_3945);
and U4615 (N_4615,N_3617,N_2173);
and U4616 (N_4616,N_2693,N_3694);
nor U4617 (N_4617,N_3263,N_3578);
nor U4618 (N_4618,N_2336,N_2635);
and U4619 (N_4619,N_2494,N_3831);
nand U4620 (N_4620,N_2160,N_3206);
nor U4621 (N_4621,N_3549,N_2803);
or U4622 (N_4622,N_2013,N_3816);
or U4623 (N_4623,N_2947,N_3837);
nor U4624 (N_4624,N_2102,N_2572);
nor U4625 (N_4625,N_2997,N_3716);
and U4626 (N_4626,N_3405,N_3446);
nand U4627 (N_4627,N_2960,N_3407);
nand U4628 (N_4628,N_3885,N_2385);
and U4629 (N_4629,N_3619,N_3971);
and U4630 (N_4630,N_3814,N_3033);
nand U4631 (N_4631,N_2169,N_2778);
or U4632 (N_4632,N_2430,N_3314);
nand U4633 (N_4633,N_3813,N_2597);
or U4634 (N_4634,N_3936,N_3713);
or U4635 (N_4635,N_2824,N_2370);
nor U4636 (N_4636,N_2765,N_2644);
and U4637 (N_4637,N_2864,N_3202);
or U4638 (N_4638,N_2649,N_3022);
nor U4639 (N_4639,N_3642,N_3668);
nand U4640 (N_4640,N_3648,N_2501);
nand U4641 (N_4641,N_3385,N_2850);
and U4642 (N_4642,N_2627,N_3898);
nor U4643 (N_4643,N_2340,N_2320);
or U4644 (N_4644,N_2515,N_2467);
nor U4645 (N_4645,N_2723,N_2206);
nor U4646 (N_4646,N_2323,N_3057);
nand U4647 (N_4647,N_2817,N_2228);
nand U4648 (N_4648,N_2564,N_2609);
nor U4649 (N_4649,N_2084,N_2898);
and U4650 (N_4650,N_3213,N_2678);
or U4651 (N_4651,N_2560,N_2191);
nand U4652 (N_4652,N_2089,N_3880);
and U4653 (N_4653,N_3053,N_3183);
or U4654 (N_4654,N_3599,N_3630);
nand U4655 (N_4655,N_3758,N_2162);
or U4656 (N_4656,N_2813,N_2061);
and U4657 (N_4657,N_2869,N_3654);
and U4658 (N_4658,N_2694,N_2457);
nand U4659 (N_4659,N_2495,N_2825);
nor U4660 (N_4660,N_3612,N_2056);
nand U4661 (N_4661,N_2017,N_2968);
or U4662 (N_4662,N_2412,N_3698);
nor U4663 (N_4663,N_3203,N_3434);
or U4664 (N_4664,N_2423,N_3367);
nor U4665 (N_4665,N_3556,N_3499);
or U4666 (N_4666,N_3313,N_3949);
or U4667 (N_4667,N_3265,N_3415);
and U4668 (N_4668,N_2448,N_2801);
nand U4669 (N_4669,N_3081,N_3254);
nor U4670 (N_4670,N_3909,N_3590);
or U4671 (N_4671,N_2352,N_2337);
xnor U4672 (N_4672,N_2163,N_2315);
and U4673 (N_4673,N_3382,N_2925);
or U4674 (N_4674,N_2029,N_3125);
and U4675 (N_4675,N_2216,N_3570);
nand U4676 (N_4676,N_3676,N_2388);
and U4677 (N_4677,N_2679,N_2908);
nor U4678 (N_4678,N_2279,N_3488);
nor U4679 (N_4679,N_2987,N_3231);
or U4680 (N_4680,N_3652,N_3128);
and U4681 (N_4681,N_2444,N_3280);
or U4682 (N_4682,N_3266,N_2411);
and U4683 (N_4683,N_2250,N_3134);
and U4684 (N_4684,N_3842,N_2197);
and U4685 (N_4685,N_3815,N_3269);
or U4686 (N_4686,N_2028,N_3038);
nand U4687 (N_4687,N_3520,N_2636);
nand U4688 (N_4688,N_2830,N_2341);
and U4689 (N_4689,N_2565,N_2292);
nor U4690 (N_4690,N_2971,N_2124);
nand U4691 (N_4691,N_2291,N_3433);
and U4692 (N_4692,N_3037,N_3009);
and U4693 (N_4693,N_3685,N_3760);
nand U4694 (N_4694,N_2424,N_3492);
or U4695 (N_4695,N_3093,N_3074);
and U4696 (N_4696,N_2883,N_3193);
and U4697 (N_4697,N_2988,N_3138);
and U4698 (N_4698,N_2175,N_3007);
nand U4699 (N_4699,N_3912,N_3424);
nor U4700 (N_4700,N_3498,N_3378);
or U4701 (N_4701,N_2787,N_2902);
nand U4702 (N_4702,N_2456,N_3396);
and U4703 (N_4703,N_2498,N_3117);
and U4704 (N_4704,N_3786,N_3130);
nor U4705 (N_4705,N_3369,N_2445);
or U4706 (N_4706,N_2496,N_2178);
nor U4707 (N_4707,N_2298,N_2688);
nor U4708 (N_4708,N_3398,N_2735);
and U4709 (N_4709,N_3435,N_3719);
nor U4710 (N_4710,N_2362,N_3722);
or U4711 (N_4711,N_3431,N_2617);
or U4712 (N_4712,N_3893,N_3771);
nor U4713 (N_4713,N_3155,N_2242);
nand U4714 (N_4714,N_2893,N_2833);
and U4715 (N_4715,N_3917,N_2402);
and U4716 (N_4716,N_3924,N_3148);
and U4717 (N_4717,N_3638,N_2368);
and U4718 (N_4718,N_2329,N_2487);
nand U4719 (N_4719,N_3783,N_3332);
or U4720 (N_4720,N_3120,N_2360);
nand U4721 (N_4721,N_3873,N_3544);
or U4722 (N_4722,N_3312,N_2932);
nand U4723 (N_4723,N_3338,N_2118);
nand U4724 (N_4724,N_3849,N_3192);
nand U4725 (N_4725,N_2585,N_3683);
nand U4726 (N_4726,N_2632,N_2763);
and U4727 (N_4727,N_2712,N_3904);
nor U4728 (N_4728,N_3869,N_3277);
nor U4729 (N_4729,N_3935,N_2500);
or U4730 (N_4730,N_3985,N_3973);
or U4731 (N_4731,N_3823,N_3925);
and U4732 (N_4732,N_2965,N_3740);
nor U4733 (N_4733,N_2849,N_3752);
nand U4734 (N_4734,N_3118,N_3316);
or U4735 (N_4735,N_3286,N_2280);
or U4736 (N_4736,N_2138,N_2470);
and U4737 (N_4737,N_2365,N_3453);
nor U4738 (N_4738,N_2425,N_3000);
or U4739 (N_4739,N_3171,N_2477);
and U4740 (N_4740,N_3357,N_2607);
or U4741 (N_4741,N_2393,N_2151);
nand U4742 (N_4742,N_2027,N_2707);
nor U4743 (N_4743,N_2806,N_3474);
nand U4744 (N_4744,N_3335,N_3997);
nor U4745 (N_4745,N_3412,N_3108);
nand U4746 (N_4746,N_3538,N_3613);
nand U4747 (N_4747,N_2862,N_3411);
and U4748 (N_4748,N_2081,N_2265);
and U4749 (N_4749,N_3843,N_2380);
or U4750 (N_4750,N_2736,N_3746);
or U4751 (N_4751,N_3967,N_3355);
nor U4752 (N_4752,N_3980,N_3467);
or U4753 (N_4753,N_3854,N_3697);
nor U4754 (N_4754,N_3289,N_2665);
nand U4755 (N_4755,N_3524,N_2042);
or U4756 (N_4756,N_2294,N_2976);
nand U4757 (N_4757,N_3970,N_3270);
and U4758 (N_4758,N_3626,N_3982);
nand U4759 (N_4759,N_2020,N_3215);
nor U4760 (N_4760,N_3163,N_3158);
and U4761 (N_4761,N_2070,N_3828);
nor U4762 (N_4762,N_2462,N_2818);
and U4763 (N_4763,N_2578,N_3847);
nand U4764 (N_4764,N_3350,N_2871);
and U4765 (N_4765,N_2026,N_3121);
and U4766 (N_4766,N_2363,N_2465);
and U4767 (N_4767,N_2229,N_3199);
and U4768 (N_4768,N_2848,N_2296);
and U4769 (N_4769,N_3540,N_3198);
or U4770 (N_4770,N_2892,N_2140);
nand U4771 (N_4771,N_3462,N_3705);
or U4772 (N_4772,N_2861,N_2554);
and U4773 (N_4773,N_3593,N_2171);
nor U4774 (N_4774,N_3224,N_3921);
and U4775 (N_4775,N_3450,N_3675);
or U4776 (N_4776,N_2919,N_3095);
or U4777 (N_4777,N_3218,N_2149);
or U4778 (N_4778,N_3583,N_2774);
and U4779 (N_4779,N_2837,N_2747);
and U4780 (N_4780,N_3867,N_3808);
nand U4781 (N_4781,N_2950,N_3864);
nand U4782 (N_4782,N_2729,N_2343);
xor U4783 (N_4783,N_2287,N_2506);
or U4784 (N_4784,N_3379,N_3208);
nor U4785 (N_4785,N_2559,N_3371);
nand U4786 (N_4786,N_2389,N_3766);
and U4787 (N_4787,N_2719,N_3750);
nand U4788 (N_4788,N_2910,N_2335);
and U4789 (N_4789,N_2985,N_3345);
and U4790 (N_4790,N_2970,N_3574);
and U4791 (N_4791,N_2684,N_3662);
nor U4792 (N_4792,N_3374,N_3323);
nor U4793 (N_4793,N_2852,N_2954);
or U4794 (N_4794,N_3983,N_3841);
and U4795 (N_4795,N_2001,N_2351);
nand U4796 (N_4796,N_3421,N_3792);
or U4797 (N_4797,N_3927,N_3607);
and U4798 (N_4798,N_2099,N_2446);
or U4799 (N_4799,N_2108,N_2654);
and U4800 (N_4800,N_2889,N_3221);
or U4801 (N_4801,N_2621,N_3601);
nand U4802 (N_4802,N_2053,N_3701);
nor U4803 (N_4803,N_2663,N_2290);
or U4804 (N_4804,N_2951,N_2807);
nand U4805 (N_4805,N_3702,N_3328);
nor U4806 (N_4806,N_3550,N_3013);
nand U4807 (N_4807,N_3090,N_2992);
xor U4808 (N_4808,N_2190,N_3204);
or U4809 (N_4809,N_2921,N_3564);
nand U4810 (N_4810,N_2808,N_3572);
nor U4811 (N_4811,N_2647,N_3085);
and U4812 (N_4812,N_3940,N_3140);
nand U4813 (N_4813,N_2756,N_2330);
nand U4814 (N_4814,N_2012,N_2038);
nor U4815 (N_4815,N_2973,N_2933);
or U4816 (N_4816,N_2528,N_2847);
or U4817 (N_4817,N_2531,N_2810);
nor U4818 (N_4818,N_3853,N_3600);
and U4819 (N_4819,N_2058,N_2008);
and U4820 (N_4820,N_2924,N_2615);
xor U4821 (N_4821,N_3188,N_3905);
nand U4822 (N_4822,N_3865,N_2010);
and U4823 (N_4823,N_3344,N_3050);
or U4824 (N_4824,N_2071,N_3112);
and U4825 (N_4825,N_2464,N_2413);
nor U4826 (N_4826,N_2722,N_2878);
nand U4827 (N_4827,N_2088,N_2616);
nand U4828 (N_4828,N_2840,N_2131);
and U4829 (N_4829,N_2247,N_3913);
or U4830 (N_4830,N_3690,N_2122);
nand U4831 (N_4831,N_3167,N_3981);
or U4832 (N_4832,N_3751,N_2880);
and U4833 (N_4833,N_2382,N_2342);
nor U4834 (N_4834,N_2507,N_2730);
nor U4835 (N_4835,N_2355,N_2859);
or U4836 (N_4836,N_2681,N_2354);
and U4837 (N_4837,N_3999,N_3387);
or U4838 (N_4838,N_3886,N_3465);
or U4839 (N_4839,N_2907,N_3563);
and U4840 (N_4840,N_2427,N_3957);
nor U4841 (N_4841,N_2421,N_2662);
or U4842 (N_4842,N_3568,N_3238);
nor U4843 (N_4843,N_3829,N_3628);
or U4844 (N_4844,N_3105,N_3761);
and U4845 (N_4845,N_2845,N_3466);
and U4846 (N_4846,N_3442,N_3294);
and U4847 (N_4847,N_3067,N_3879);
nor U4848 (N_4848,N_2638,N_2332);
and U4849 (N_4849,N_3779,N_2576);
nand U4850 (N_4850,N_2548,N_3649);
or U4851 (N_4851,N_2325,N_3883);
and U4852 (N_4852,N_2019,N_2004);
and U4853 (N_4853,N_2075,N_3444);
or U4854 (N_4854,N_2264,N_2168);
nor U4855 (N_4855,N_3111,N_3820);
nor U4856 (N_4856,N_3624,N_2920);
or U4857 (N_4857,N_3414,N_2497);
nor U4858 (N_4858,N_2581,N_2668);
nand U4859 (N_4859,N_2377,N_2641);
and U4860 (N_4860,N_3417,N_3557);
and U4861 (N_4861,N_3399,N_2077);
and U4862 (N_4862,N_2439,N_2596);
or U4863 (N_4863,N_3441,N_2275);
and U4864 (N_4864,N_2396,N_3042);
and U4865 (N_4865,N_3016,N_3542);
and U4866 (N_4866,N_2309,N_3625);
nor U4867 (N_4867,N_2128,N_2450);
or U4868 (N_4868,N_3926,N_2568);
or U4869 (N_4869,N_2682,N_2449);
or U4870 (N_4870,N_2044,N_2063);
and U4871 (N_4871,N_3391,N_2356);
or U4872 (N_4872,N_2798,N_2624);
and U4873 (N_4873,N_2072,N_3620);
or U4874 (N_4874,N_2727,N_3689);
and U4875 (N_4875,N_3914,N_2687);
nor U4876 (N_4876,N_2052,N_3569);
and U4877 (N_4877,N_3523,N_3480);
and U4878 (N_4878,N_2461,N_2066);
or U4879 (N_4879,N_2079,N_2036);
or U4880 (N_4880,N_3616,N_3063);
and U4881 (N_4881,N_2750,N_2598);
nor U4882 (N_4882,N_2670,N_2546);
nand U4883 (N_4883,N_3834,N_3103);
nor U4884 (N_4884,N_3083,N_3321);
or U4885 (N_4885,N_3720,N_3646);
nand U4886 (N_4886,N_3793,N_2957);
or U4887 (N_4887,N_2468,N_2478);
nor U4888 (N_4888,N_2132,N_2744);
or U4889 (N_4889,N_3054,N_3762);
and U4890 (N_4890,N_3530,N_3637);
and U4891 (N_4891,N_3306,N_3119);
nand U4892 (N_4892,N_2502,N_2571);
and U4893 (N_4893,N_2740,N_3315);
nand U4894 (N_4894,N_3305,N_3991);
nand U4895 (N_4895,N_2234,N_2314);
or U4896 (N_4896,N_3605,N_2720);
nor U4897 (N_4897,N_2673,N_3811);
and U4898 (N_4898,N_3518,N_3334);
and U4899 (N_4899,N_3182,N_3650);
nand U4900 (N_4900,N_2418,N_2873);
and U4901 (N_4901,N_2404,N_2268);
or U4902 (N_4902,N_3727,N_2562);
or U4903 (N_4903,N_3594,N_3989);
nand U4904 (N_4904,N_3884,N_3858);
nor U4905 (N_4905,N_3502,N_3283);
or U4906 (N_4906,N_3447,N_3223);
and U4907 (N_4907,N_2025,N_3872);
nor U4908 (N_4908,N_2297,N_3958);
nor U4909 (N_4909,N_3320,N_2186);
and U4910 (N_4910,N_3184,N_3330);
or U4911 (N_4911,N_3260,N_3922);
and U4912 (N_4912,N_2201,N_2366);
nand U4913 (N_4913,N_2709,N_3674);
or U4914 (N_4914,N_2489,N_3818);
and U4915 (N_4915,N_2805,N_2317);
or U4916 (N_4916,N_3032,N_2591);
and U4917 (N_4917,N_2408,N_2405);
nand U4918 (N_4918,N_3471,N_3978);
or U4919 (N_4919,N_2326,N_3333);
and U4920 (N_4920,N_2676,N_3468);
nand U4921 (N_4921,N_2675,N_3573);
and U4922 (N_4922,N_3066,N_3787);
nand U4923 (N_4923,N_2005,N_2387);
nand U4924 (N_4924,N_3482,N_3585);
nor U4925 (N_4925,N_3457,N_2877);
or U4926 (N_4926,N_3658,N_3803);
nor U4927 (N_4927,N_2611,N_3651);
or U4928 (N_4928,N_2263,N_3246);
and U4929 (N_4929,N_2998,N_3670);
nand U4930 (N_4930,N_2926,N_3248);
and U4931 (N_4931,N_3852,N_2324);
or U4932 (N_4932,N_3875,N_3272);
nand U4933 (N_4933,N_3712,N_2509);
nor U4934 (N_4934,N_3324,N_3485);
nor U4935 (N_4935,N_2646,N_3744);
and U4936 (N_4936,N_2994,N_3234);
nor U4937 (N_4937,N_2819,N_2199);
and U4938 (N_4938,N_3591,N_3611);
and U4939 (N_4939,N_2085,N_3882);
and U4940 (N_4940,N_3505,N_2683);
or U4941 (N_4941,N_2142,N_2133);
and U4942 (N_4942,N_3659,N_3577);
and U4943 (N_4943,N_3798,N_2732);
and U4944 (N_4944,N_2147,N_3026);
nor U4945 (N_4945,N_3115,N_3749);
or U4946 (N_4946,N_3669,N_3191);
nand U4947 (N_4947,N_3132,N_3423);
nand U4948 (N_4948,N_3353,N_2570);
and U4949 (N_4949,N_2664,N_3174);
nand U4950 (N_4950,N_3039,N_2045);
xnor U4951 (N_4951,N_3472,N_2652);
nand U4952 (N_4952,N_3655,N_2713);
nand U4953 (N_4953,N_3175,N_2473);
or U4954 (N_4954,N_3440,N_2569);
nor U4955 (N_4955,N_2397,N_3064);
nor U4956 (N_4956,N_3473,N_2244);
nand U4957 (N_4957,N_2704,N_2344);
and U4958 (N_4958,N_3801,N_3555);
and U4959 (N_4959,N_2786,N_3166);
nand U4960 (N_4960,N_2453,N_3291);
and U4961 (N_4961,N_3592,N_2962);
and U4962 (N_4962,N_3665,N_2826);
nand U4963 (N_4963,N_3360,N_3500);
nand U4964 (N_4964,N_3288,N_3436);
and U4965 (N_4965,N_2381,N_3495);
xor U4966 (N_4966,N_2643,N_2984);
nand U4967 (N_4967,N_2595,N_2629);
nor U4968 (N_4968,N_3772,N_3844);
or U4969 (N_4969,N_2517,N_3954);
nand U4970 (N_4970,N_2249,N_2107);
or U4971 (N_4971,N_3693,N_3437);
and U4972 (N_4972,N_3351,N_3838);
nand U4973 (N_4973,N_2129,N_3706);
nor U4974 (N_4974,N_2745,N_3799);
or U4975 (N_4975,N_3102,N_2159);
nand U4976 (N_4976,N_2371,N_2592);
nor U4977 (N_4977,N_3955,N_3968);
and U4978 (N_4978,N_3197,N_2530);
nand U4979 (N_4979,N_2972,N_3209);
or U4980 (N_4980,N_2021,N_3491);
or U4981 (N_4981,N_3402,N_3923);
or U4982 (N_4982,N_2844,N_3279);
or U4983 (N_4983,N_3998,N_3489);
nor U4984 (N_4984,N_2059,N_2230);
and U4985 (N_4985,N_3687,N_3483);
and U4986 (N_4986,N_2415,N_3966);
and U4987 (N_4987,N_2863,N_2245);
nand U4988 (N_4988,N_2916,N_3461);
nor U4989 (N_4989,N_3071,N_3302);
nand U4990 (N_4990,N_2695,N_2033);
nor U4991 (N_4991,N_3929,N_3581);
nor U4992 (N_4992,N_3418,N_2455);
or U4993 (N_4993,N_3615,N_2055);
nor U4994 (N_4994,N_3189,N_2143);
nand U4995 (N_4995,N_2083,N_3623);
and U4996 (N_4996,N_2587,N_3100);
and U4997 (N_4997,N_2700,N_2318);
xor U4998 (N_4998,N_2091,N_2499);
nand U4999 (N_4999,N_3773,N_3684);
or U5000 (N_5000,N_3215,N_3898);
nor U5001 (N_5001,N_3227,N_3186);
or U5002 (N_5002,N_3859,N_3175);
nand U5003 (N_5003,N_2258,N_2605);
nand U5004 (N_5004,N_2224,N_3836);
or U5005 (N_5005,N_2292,N_2522);
or U5006 (N_5006,N_2228,N_3647);
or U5007 (N_5007,N_3201,N_3239);
nand U5008 (N_5008,N_3222,N_3444);
or U5009 (N_5009,N_2552,N_2077);
and U5010 (N_5010,N_2717,N_3505);
and U5011 (N_5011,N_3692,N_3770);
nand U5012 (N_5012,N_2847,N_3066);
and U5013 (N_5013,N_3050,N_2807);
and U5014 (N_5014,N_2793,N_2573);
and U5015 (N_5015,N_3605,N_2849);
nand U5016 (N_5016,N_3020,N_2497);
nor U5017 (N_5017,N_2587,N_3909);
and U5018 (N_5018,N_3071,N_3688);
nor U5019 (N_5019,N_2115,N_2631);
and U5020 (N_5020,N_2672,N_3873);
nand U5021 (N_5021,N_3144,N_2222);
nor U5022 (N_5022,N_2997,N_2662);
nor U5023 (N_5023,N_2664,N_2445);
or U5024 (N_5024,N_3534,N_2594);
and U5025 (N_5025,N_3953,N_3831);
xor U5026 (N_5026,N_3258,N_3115);
nand U5027 (N_5027,N_2868,N_3045);
xor U5028 (N_5028,N_3134,N_2457);
nand U5029 (N_5029,N_2147,N_2749);
or U5030 (N_5030,N_3560,N_3373);
or U5031 (N_5031,N_3652,N_3296);
nor U5032 (N_5032,N_2125,N_3228);
nor U5033 (N_5033,N_2518,N_3646);
nand U5034 (N_5034,N_2150,N_3083);
and U5035 (N_5035,N_3789,N_3971);
and U5036 (N_5036,N_3678,N_3638);
and U5037 (N_5037,N_2244,N_2409);
and U5038 (N_5038,N_3569,N_2388);
and U5039 (N_5039,N_3033,N_2232);
and U5040 (N_5040,N_3308,N_2907);
nor U5041 (N_5041,N_3356,N_3433);
nor U5042 (N_5042,N_3290,N_2754);
nand U5043 (N_5043,N_3780,N_3310);
nand U5044 (N_5044,N_3575,N_3088);
nand U5045 (N_5045,N_3906,N_3864);
nand U5046 (N_5046,N_2802,N_2814);
and U5047 (N_5047,N_3007,N_3868);
nand U5048 (N_5048,N_2976,N_2949);
or U5049 (N_5049,N_2051,N_2344);
nand U5050 (N_5050,N_3741,N_2224);
nand U5051 (N_5051,N_2560,N_2249);
nand U5052 (N_5052,N_3894,N_3973);
nand U5053 (N_5053,N_3816,N_2591);
nor U5054 (N_5054,N_3925,N_3351);
or U5055 (N_5055,N_3440,N_2842);
and U5056 (N_5056,N_2395,N_3213);
nor U5057 (N_5057,N_2212,N_2585);
nand U5058 (N_5058,N_3880,N_3097);
nor U5059 (N_5059,N_3143,N_2036);
and U5060 (N_5060,N_3395,N_3058);
nand U5061 (N_5061,N_3452,N_3716);
nor U5062 (N_5062,N_3259,N_3756);
nor U5063 (N_5063,N_3012,N_3679);
nand U5064 (N_5064,N_2503,N_2732);
or U5065 (N_5065,N_3964,N_2427);
xor U5066 (N_5066,N_2854,N_2985);
nand U5067 (N_5067,N_2736,N_2143);
nand U5068 (N_5068,N_3400,N_3959);
nand U5069 (N_5069,N_3762,N_3392);
nand U5070 (N_5070,N_3872,N_3925);
nand U5071 (N_5071,N_2498,N_2497);
nor U5072 (N_5072,N_3591,N_3068);
and U5073 (N_5073,N_2317,N_3445);
or U5074 (N_5074,N_2258,N_3470);
nor U5075 (N_5075,N_2162,N_2663);
nand U5076 (N_5076,N_2035,N_3439);
nor U5077 (N_5077,N_3726,N_3453);
nor U5078 (N_5078,N_3092,N_2056);
nand U5079 (N_5079,N_3358,N_2572);
or U5080 (N_5080,N_2584,N_3589);
or U5081 (N_5081,N_2287,N_2152);
nor U5082 (N_5082,N_2259,N_2709);
nor U5083 (N_5083,N_2236,N_2499);
nand U5084 (N_5084,N_3542,N_3245);
or U5085 (N_5085,N_3470,N_2032);
and U5086 (N_5086,N_3974,N_3995);
and U5087 (N_5087,N_3280,N_2529);
or U5088 (N_5088,N_2769,N_3346);
and U5089 (N_5089,N_2983,N_2130);
or U5090 (N_5090,N_3503,N_3387);
nor U5091 (N_5091,N_2102,N_2537);
nand U5092 (N_5092,N_2229,N_2196);
nor U5093 (N_5093,N_2310,N_2153);
nand U5094 (N_5094,N_3048,N_2824);
nand U5095 (N_5095,N_3809,N_3554);
and U5096 (N_5096,N_3248,N_2695);
nand U5097 (N_5097,N_2010,N_3545);
nor U5098 (N_5098,N_3588,N_3634);
and U5099 (N_5099,N_3300,N_3236);
nand U5100 (N_5100,N_2831,N_2836);
nand U5101 (N_5101,N_2998,N_2807);
and U5102 (N_5102,N_3393,N_3347);
nor U5103 (N_5103,N_3899,N_2600);
nand U5104 (N_5104,N_2661,N_2245);
nand U5105 (N_5105,N_3465,N_3176);
nor U5106 (N_5106,N_2459,N_2233);
nand U5107 (N_5107,N_2552,N_3111);
or U5108 (N_5108,N_3068,N_2708);
and U5109 (N_5109,N_2308,N_2781);
and U5110 (N_5110,N_3458,N_3962);
nand U5111 (N_5111,N_3482,N_2247);
nor U5112 (N_5112,N_3590,N_3623);
nor U5113 (N_5113,N_2329,N_3242);
and U5114 (N_5114,N_3430,N_2223);
nor U5115 (N_5115,N_3411,N_2776);
xnor U5116 (N_5116,N_2965,N_2160);
xor U5117 (N_5117,N_3716,N_2312);
nand U5118 (N_5118,N_3095,N_3167);
and U5119 (N_5119,N_3404,N_3833);
xnor U5120 (N_5120,N_3766,N_3378);
nor U5121 (N_5121,N_3491,N_2467);
nand U5122 (N_5122,N_2030,N_3015);
nor U5123 (N_5123,N_3744,N_3004);
or U5124 (N_5124,N_3453,N_2514);
nor U5125 (N_5125,N_3362,N_2982);
nand U5126 (N_5126,N_3682,N_3454);
nand U5127 (N_5127,N_2648,N_2191);
and U5128 (N_5128,N_2796,N_3308);
nand U5129 (N_5129,N_2837,N_3922);
and U5130 (N_5130,N_3655,N_2161);
and U5131 (N_5131,N_3106,N_3949);
nand U5132 (N_5132,N_2884,N_3992);
and U5133 (N_5133,N_3743,N_3279);
nor U5134 (N_5134,N_2509,N_2686);
and U5135 (N_5135,N_2795,N_3210);
nand U5136 (N_5136,N_3074,N_3398);
and U5137 (N_5137,N_2166,N_2501);
and U5138 (N_5138,N_3103,N_2877);
or U5139 (N_5139,N_3627,N_2734);
or U5140 (N_5140,N_2580,N_3478);
and U5141 (N_5141,N_3725,N_2372);
nor U5142 (N_5142,N_2100,N_3237);
or U5143 (N_5143,N_2419,N_2208);
nor U5144 (N_5144,N_3398,N_3582);
nand U5145 (N_5145,N_3493,N_3960);
or U5146 (N_5146,N_2942,N_3526);
and U5147 (N_5147,N_3619,N_3948);
or U5148 (N_5148,N_2437,N_3554);
nand U5149 (N_5149,N_3312,N_2608);
nand U5150 (N_5150,N_2844,N_3549);
or U5151 (N_5151,N_2336,N_3726);
or U5152 (N_5152,N_2730,N_2101);
nand U5153 (N_5153,N_3653,N_2534);
nor U5154 (N_5154,N_2922,N_3222);
and U5155 (N_5155,N_2069,N_3602);
or U5156 (N_5156,N_2503,N_2950);
nor U5157 (N_5157,N_3473,N_2792);
and U5158 (N_5158,N_3935,N_2873);
nand U5159 (N_5159,N_3791,N_2060);
or U5160 (N_5160,N_2977,N_3350);
or U5161 (N_5161,N_2459,N_2375);
nor U5162 (N_5162,N_3873,N_2394);
and U5163 (N_5163,N_3809,N_3699);
and U5164 (N_5164,N_2950,N_3499);
nand U5165 (N_5165,N_2115,N_2875);
and U5166 (N_5166,N_3608,N_2830);
nand U5167 (N_5167,N_3403,N_3958);
and U5168 (N_5168,N_2189,N_2544);
nand U5169 (N_5169,N_3361,N_3873);
nand U5170 (N_5170,N_2014,N_3573);
nor U5171 (N_5171,N_3626,N_3262);
and U5172 (N_5172,N_2112,N_3386);
nand U5173 (N_5173,N_3857,N_2224);
nand U5174 (N_5174,N_2927,N_3195);
nor U5175 (N_5175,N_3423,N_2304);
or U5176 (N_5176,N_2483,N_3536);
nand U5177 (N_5177,N_3525,N_2018);
nor U5178 (N_5178,N_2179,N_2604);
nor U5179 (N_5179,N_3454,N_2944);
nand U5180 (N_5180,N_3139,N_2190);
and U5181 (N_5181,N_3060,N_2846);
or U5182 (N_5182,N_2923,N_3564);
or U5183 (N_5183,N_2692,N_3742);
and U5184 (N_5184,N_2426,N_2899);
and U5185 (N_5185,N_3423,N_3367);
nand U5186 (N_5186,N_2512,N_3257);
nor U5187 (N_5187,N_2260,N_3061);
nand U5188 (N_5188,N_2434,N_3568);
and U5189 (N_5189,N_3306,N_3944);
or U5190 (N_5190,N_3760,N_3134);
and U5191 (N_5191,N_3186,N_2844);
and U5192 (N_5192,N_3002,N_2817);
nand U5193 (N_5193,N_3357,N_3894);
and U5194 (N_5194,N_2243,N_2459);
nand U5195 (N_5195,N_2199,N_3249);
or U5196 (N_5196,N_3951,N_2104);
or U5197 (N_5197,N_2847,N_3824);
or U5198 (N_5198,N_3296,N_3697);
and U5199 (N_5199,N_2471,N_3075);
nor U5200 (N_5200,N_2140,N_2324);
or U5201 (N_5201,N_3986,N_3469);
nor U5202 (N_5202,N_3163,N_3997);
and U5203 (N_5203,N_3158,N_3736);
or U5204 (N_5204,N_2170,N_2035);
or U5205 (N_5205,N_3405,N_3323);
or U5206 (N_5206,N_2183,N_2495);
nor U5207 (N_5207,N_2006,N_3022);
nand U5208 (N_5208,N_2879,N_3487);
or U5209 (N_5209,N_2041,N_3294);
nor U5210 (N_5210,N_3713,N_3125);
and U5211 (N_5211,N_2168,N_2014);
and U5212 (N_5212,N_2393,N_3257);
or U5213 (N_5213,N_2480,N_2263);
nor U5214 (N_5214,N_2581,N_3035);
or U5215 (N_5215,N_3823,N_2192);
or U5216 (N_5216,N_3606,N_3718);
and U5217 (N_5217,N_2870,N_3305);
nand U5218 (N_5218,N_3733,N_2251);
nand U5219 (N_5219,N_3191,N_2632);
nor U5220 (N_5220,N_2856,N_2982);
and U5221 (N_5221,N_3117,N_3191);
nor U5222 (N_5222,N_3360,N_2544);
nand U5223 (N_5223,N_3297,N_3533);
and U5224 (N_5224,N_3583,N_2168);
and U5225 (N_5225,N_3831,N_3847);
and U5226 (N_5226,N_3494,N_2843);
nor U5227 (N_5227,N_3700,N_3602);
nor U5228 (N_5228,N_2297,N_3382);
nor U5229 (N_5229,N_2468,N_2497);
and U5230 (N_5230,N_3848,N_2608);
or U5231 (N_5231,N_2711,N_2615);
and U5232 (N_5232,N_2026,N_2906);
nor U5233 (N_5233,N_3049,N_2069);
nand U5234 (N_5234,N_3607,N_2269);
nand U5235 (N_5235,N_3075,N_3770);
nor U5236 (N_5236,N_2994,N_2098);
and U5237 (N_5237,N_2058,N_2083);
nor U5238 (N_5238,N_3455,N_3558);
or U5239 (N_5239,N_2653,N_3961);
nand U5240 (N_5240,N_2907,N_3977);
or U5241 (N_5241,N_2640,N_2419);
nor U5242 (N_5242,N_2246,N_3679);
nand U5243 (N_5243,N_3856,N_3542);
nor U5244 (N_5244,N_2071,N_2447);
nor U5245 (N_5245,N_2722,N_3361);
xor U5246 (N_5246,N_2872,N_2897);
nor U5247 (N_5247,N_2105,N_2828);
nand U5248 (N_5248,N_3901,N_3738);
and U5249 (N_5249,N_3054,N_2663);
or U5250 (N_5250,N_3568,N_3539);
nand U5251 (N_5251,N_2549,N_2445);
or U5252 (N_5252,N_3313,N_3907);
and U5253 (N_5253,N_3342,N_3228);
nor U5254 (N_5254,N_3051,N_3940);
and U5255 (N_5255,N_2437,N_3347);
and U5256 (N_5256,N_2639,N_2552);
nand U5257 (N_5257,N_3821,N_2186);
or U5258 (N_5258,N_2211,N_3150);
nor U5259 (N_5259,N_3645,N_3160);
nor U5260 (N_5260,N_3185,N_2145);
and U5261 (N_5261,N_2731,N_3454);
nor U5262 (N_5262,N_3748,N_2626);
or U5263 (N_5263,N_2355,N_2729);
or U5264 (N_5264,N_2847,N_3275);
or U5265 (N_5265,N_3105,N_3923);
nand U5266 (N_5266,N_2960,N_3799);
or U5267 (N_5267,N_2246,N_2783);
and U5268 (N_5268,N_3521,N_3646);
or U5269 (N_5269,N_3971,N_2929);
or U5270 (N_5270,N_3549,N_3217);
and U5271 (N_5271,N_2988,N_3566);
nand U5272 (N_5272,N_3905,N_2944);
nand U5273 (N_5273,N_3682,N_2687);
nor U5274 (N_5274,N_3805,N_3738);
and U5275 (N_5275,N_2295,N_3514);
or U5276 (N_5276,N_2606,N_3735);
nand U5277 (N_5277,N_3978,N_3145);
and U5278 (N_5278,N_3417,N_2791);
or U5279 (N_5279,N_3329,N_3198);
nand U5280 (N_5280,N_3290,N_3794);
nand U5281 (N_5281,N_2506,N_3876);
nand U5282 (N_5282,N_2950,N_2223);
nor U5283 (N_5283,N_2418,N_3864);
or U5284 (N_5284,N_3066,N_2117);
or U5285 (N_5285,N_2829,N_3501);
and U5286 (N_5286,N_3084,N_2267);
and U5287 (N_5287,N_2891,N_3332);
nor U5288 (N_5288,N_3769,N_2670);
and U5289 (N_5289,N_2734,N_3293);
nand U5290 (N_5290,N_3728,N_2071);
and U5291 (N_5291,N_3604,N_3572);
and U5292 (N_5292,N_2859,N_2380);
nand U5293 (N_5293,N_2672,N_3439);
nand U5294 (N_5294,N_3741,N_3264);
nand U5295 (N_5295,N_3040,N_3475);
nor U5296 (N_5296,N_2347,N_2150);
nand U5297 (N_5297,N_2498,N_3063);
or U5298 (N_5298,N_2925,N_3010);
or U5299 (N_5299,N_2230,N_3282);
nand U5300 (N_5300,N_2983,N_2646);
or U5301 (N_5301,N_3835,N_2263);
nand U5302 (N_5302,N_3060,N_2775);
and U5303 (N_5303,N_2447,N_3787);
or U5304 (N_5304,N_3043,N_3728);
nand U5305 (N_5305,N_3069,N_3758);
nor U5306 (N_5306,N_3517,N_2358);
and U5307 (N_5307,N_3002,N_2123);
nand U5308 (N_5308,N_2500,N_2518);
or U5309 (N_5309,N_3386,N_3092);
and U5310 (N_5310,N_3541,N_2804);
or U5311 (N_5311,N_3464,N_3380);
and U5312 (N_5312,N_2612,N_2432);
and U5313 (N_5313,N_2044,N_2685);
nor U5314 (N_5314,N_3078,N_3303);
nor U5315 (N_5315,N_3569,N_3538);
or U5316 (N_5316,N_3357,N_2287);
or U5317 (N_5317,N_3781,N_3338);
nand U5318 (N_5318,N_3727,N_2544);
nor U5319 (N_5319,N_2537,N_2031);
or U5320 (N_5320,N_2504,N_3335);
and U5321 (N_5321,N_3211,N_3742);
or U5322 (N_5322,N_2311,N_3887);
nand U5323 (N_5323,N_2191,N_3242);
nor U5324 (N_5324,N_3485,N_3661);
nor U5325 (N_5325,N_3308,N_3693);
and U5326 (N_5326,N_3110,N_3898);
and U5327 (N_5327,N_2429,N_2599);
and U5328 (N_5328,N_3499,N_3684);
xor U5329 (N_5329,N_3272,N_2488);
or U5330 (N_5330,N_3859,N_2704);
or U5331 (N_5331,N_2577,N_3798);
nor U5332 (N_5332,N_3818,N_3566);
and U5333 (N_5333,N_2590,N_2735);
or U5334 (N_5334,N_3195,N_2719);
nand U5335 (N_5335,N_2371,N_3024);
or U5336 (N_5336,N_2000,N_3771);
or U5337 (N_5337,N_3468,N_3644);
nor U5338 (N_5338,N_2278,N_3903);
or U5339 (N_5339,N_3494,N_2278);
and U5340 (N_5340,N_3820,N_2586);
nand U5341 (N_5341,N_3410,N_2554);
nand U5342 (N_5342,N_3258,N_3176);
and U5343 (N_5343,N_2907,N_3348);
or U5344 (N_5344,N_2944,N_3828);
nor U5345 (N_5345,N_3272,N_2842);
and U5346 (N_5346,N_2864,N_3279);
nor U5347 (N_5347,N_3620,N_2935);
and U5348 (N_5348,N_3859,N_2225);
nand U5349 (N_5349,N_2938,N_2030);
or U5350 (N_5350,N_2013,N_3595);
and U5351 (N_5351,N_3295,N_2153);
nand U5352 (N_5352,N_3755,N_2035);
or U5353 (N_5353,N_3699,N_3927);
or U5354 (N_5354,N_3212,N_2945);
or U5355 (N_5355,N_3745,N_2503);
nand U5356 (N_5356,N_3149,N_3386);
nor U5357 (N_5357,N_2113,N_2801);
nand U5358 (N_5358,N_2226,N_2937);
and U5359 (N_5359,N_2261,N_3810);
nand U5360 (N_5360,N_3633,N_3851);
nor U5361 (N_5361,N_2381,N_3249);
and U5362 (N_5362,N_2035,N_2091);
or U5363 (N_5363,N_2170,N_3887);
xnor U5364 (N_5364,N_2741,N_2389);
nand U5365 (N_5365,N_2944,N_3124);
and U5366 (N_5366,N_3633,N_3296);
or U5367 (N_5367,N_3117,N_2465);
and U5368 (N_5368,N_2655,N_2396);
nand U5369 (N_5369,N_2156,N_3972);
or U5370 (N_5370,N_2278,N_2074);
nand U5371 (N_5371,N_3272,N_3048);
and U5372 (N_5372,N_2369,N_3750);
or U5373 (N_5373,N_2365,N_3764);
and U5374 (N_5374,N_3201,N_3780);
or U5375 (N_5375,N_3232,N_3823);
or U5376 (N_5376,N_2847,N_2188);
or U5377 (N_5377,N_3903,N_3440);
or U5378 (N_5378,N_3803,N_3883);
nand U5379 (N_5379,N_2662,N_2666);
or U5380 (N_5380,N_2441,N_3906);
nor U5381 (N_5381,N_2889,N_2412);
and U5382 (N_5382,N_2554,N_2976);
nand U5383 (N_5383,N_3564,N_2203);
or U5384 (N_5384,N_2591,N_3595);
or U5385 (N_5385,N_2533,N_2255);
or U5386 (N_5386,N_3147,N_2942);
nand U5387 (N_5387,N_3157,N_2190);
or U5388 (N_5388,N_2567,N_2163);
and U5389 (N_5389,N_2263,N_2036);
or U5390 (N_5390,N_2554,N_3960);
or U5391 (N_5391,N_2310,N_2911);
or U5392 (N_5392,N_3898,N_3453);
nand U5393 (N_5393,N_2139,N_3858);
and U5394 (N_5394,N_3120,N_3580);
nor U5395 (N_5395,N_3028,N_3293);
or U5396 (N_5396,N_3045,N_3543);
nand U5397 (N_5397,N_2390,N_2497);
nand U5398 (N_5398,N_2792,N_3922);
and U5399 (N_5399,N_3046,N_3494);
nand U5400 (N_5400,N_2817,N_3620);
and U5401 (N_5401,N_3666,N_3552);
nand U5402 (N_5402,N_2542,N_2825);
and U5403 (N_5403,N_2563,N_2452);
nor U5404 (N_5404,N_2598,N_3950);
nor U5405 (N_5405,N_3247,N_3504);
or U5406 (N_5406,N_3317,N_2017);
nand U5407 (N_5407,N_3925,N_3099);
or U5408 (N_5408,N_3370,N_3488);
or U5409 (N_5409,N_3640,N_3758);
nor U5410 (N_5410,N_2157,N_2520);
or U5411 (N_5411,N_2198,N_2487);
and U5412 (N_5412,N_3944,N_3429);
nor U5413 (N_5413,N_2986,N_2265);
nand U5414 (N_5414,N_3066,N_2714);
nand U5415 (N_5415,N_2454,N_2990);
nand U5416 (N_5416,N_3061,N_3190);
or U5417 (N_5417,N_2800,N_2699);
nand U5418 (N_5418,N_2163,N_3225);
or U5419 (N_5419,N_3473,N_2208);
nor U5420 (N_5420,N_3781,N_3970);
or U5421 (N_5421,N_3531,N_2147);
nand U5422 (N_5422,N_3401,N_3971);
nor U5423 (N_5423,N_3721,N_3746);
nand U5424 (N_5424,N_2674,N_2159);
nand U5425 (N_5425,N_2519,N_2885);
and U5426 (N_5426,N_3242,N_2648);
or U5427 (N_5427,N_2991,N_3263);
or U5428 (N_5428,N_3264,N_2600);
or U5429 (N_5429,N_2934,N_2329);
nand U5430 (N_5430,N_2101,N_2432);
nand U5431 (N_5431,N_2816,N_2622);
and U5432 (N_5432,N_3181,N_3043);
and U5433 (N_5433,N_3167,N_3166);
or U5434 (N_5434,N_3340,N_2720);
xnor U5435 (N_5435,N_3333,N_3458);
and U5436 (N_5436,N_3858,N_3350);
nor U5437 (N_5437,N_3987,N_2351);
nor U5438 (N_5438,N_2694,N_3355);
and U5439 (N_5439,N_2567,N_2561);
nor U5440 (N_5440,N_2553,N_2432);
nor U5441 (N_5441,N_3376,N_3675);
nand U5442 (N_5442,N_2351,N_2933);
xor U5443 (N_5443,N_3125,N_2440);
nand U5444 (N_5444,N_2929,N_2051);
nand U5445 (N_5445,N_3261,N_2823);
or U5446 (N_5446,N_3796,N_2079);
nor U5447 (N_5447,N_3636,N_2605);
nor U5448 (N_5448,N_2158,N_2491);
and U5449 (N_5449,N_3199,N_3668);
and U5450 (N_5450,N_2445,N_2601);
or U5451 (N_5451,N_2500,N_2383);
and U5452 (N_5452,N_2827,N_2272);
and U5453 (N_5453,N_3436,N_3507);
or U5454 (N_5454,N_2939,N_3723);
nor U5455 (N_5455,N_2860,N_2004);
or U5456 (N_5456,N_2909,N_2193);
nor U5457 (N_5457,N_2120,N_3660);
and U5458 (N_5458,N_2938,N_3921);
and U5459 (N_5459,N_2593,N_2129);
and U5460 (N_5460,N_2087,N_3536);
nor U5461 (N_5461,N_2627,N_3686);
and U5462 (N_5462,N_2671,N_3340);
nor U5463 (N_5463,N_2831,N_3049);
and U5464 (N_5464,N_3717,N_2752);
nor U5465 (N_5465,N_2997,N_3138);
and U5466 (N_5466,N_3257,N_3644);
nand U5467 (N_5467,N_2580,N_2415);
nand U5468 (N_5468,N_2753,N_2245);
nor U5469 (N_5469,N_2553,N_2563);
or U5470 (N_5470,N_2590,N_2281);
nand U5471 (N_5471,N_2889,N_2956);
and U5472 (N_5472,N_2972,N_2001);
nor U5473 (N_5473,N_2517,N_2010);
and U5474 (N_5474,N_2094,N_2493);
nand U5475 (N_5475,N_3326,N_2472);
nand U5476 (N_5476,N_2734,N_3443);
or U5477 (N_5477,N_3333,N_3524);
nand U5478 (N_5478,N_2421,N_2143);
or U5479 (N_5479,N_3203,N_2604);
and U5480 (N_5480,N_2409,N_2068);
nor U5481 (N_5481,N_3670,N_2837);
nand U5482 (N_5482,N_2290,N_3684);
and U5483 (N_5483,N_2118,N_3516);
nor U5484 (N_5484,N_3000,N_3760);
and U5485 (N_5485,N_2917,N_2542);
and U5486 (N_5486,N_2182,N_2290);
nor U5487 (N_5487,N_2881,N_3875);
nor U5488 (N_5488,N_2611,N_2711);
or U5489 (N_5489,N_2457,N_3810);
or U5490 (N_5490,N_2512,N_2998);
and U5491 (N_5491,N_2849,N_2015);
and U5492 (N_5492,N_3453,N_2907);
nor U5493 (N_5493,N_3501,N_2606);
or U5494 (N_5494,N_2743,N_2254);
nor U5495 (N_5495,N_2570,N_3449);
or U5496 (N_5496,N_2564,N_3166);
nor U5497 (N_5497,N_3315,N_2147);
nor U5498 (N_5498,N_2919,N_2383);
or U5499 (N_5499,N_3741,N_2807);
or U5500 (N_5500,N_2578,N_3824);
nand U5501 (N_5501,N_3830,N_3169);
nor U5502 (N_5502,N_2826,N_2424);
nand U5503 (N_5503,N_3738,N_2659);
nand U5504 (N_5504,N_2678,N_3890);
nand U5505 (N_5505,N_3813,N_3928);
or U5506 (N_5506,N_2079,N_3359);
nor U5507 (N_5507,N_2475,N_2229);
nand U5508 (N_5508,N_3629,N_3082);
and U5509 (N_5509,N_3800,N_2259);
and U5510 (N_5510,N_2150,N_2099);
nor U5511 (N_5511,N_2377,N_3241);
nand U5512 (N_5512,N_2990,N_3235);
and U5513 (N_5513,N_3477,N_3771);
nor U5514 (N_5514,N_2394,N_2210);
and U5515 (N_5515,N_3238,N_3936);
nand U5516 (N_5516,N_2711,N_3692);
nand U5517 (N_5517,N_3969,N_2488);
nand U5518 (N_5518,N_3811,N_2677);
nor U5519 (N_5519,N_3252,N_2127);
nor U5520 (N_5520,N_2546,N_3030);
nand U5521 (N_5521,N_2235,N_2863);
and U5522 (N_5522,N_2670,N_3592);
nand U5523 (N_5523,N_3890,N_2226);
and U5524 (N_5524,N_2120,N_2712);
or U5525 (N_5525,N_3649,N_3779);
or U5526 (N_5526,N_3222,N_3088);
nor U5527 (N_5527,N_2302,N_2817);
or U5528 (N_5528,N_3618,N_3034);
or U5529 (N_5529,N_3719,N_2927);
nand U5530 (N_5530,N_2137,N_3652);
and U5531 (N_5531,N_3328,N_2644);
or U5532 (N_5532,N_3365,N_2087);
and U5533 (N_5533,N_2864,N_2980);
or U5534 (N_5534,N_3288,N_3153);
nor U5535 (N_5535,N_2874,N_2047);
nand U5536 (N_5536,N_3300,N_3119);
nor U5537 (N_5537,N_2505,N_3919);
and U5538 (N_5538,N_3783,N_2513);
nand U5539 (N_5539,N_3608,N_3244);
and U5540 (N_5540,N_3931,N_2282);
or U5541 (N_5541,N_2087,N_2119);
and U5542 (N_5542,N_2379,N_2874);
or U5543 (N_5543,N_2333,N_3415);
and U5544 (N_5544,N_2101,N_2813);
and U5545 (N_5545,N_2529,N_2072);
nand U5546 (N_5546,N_2119,N_2454);
and U5547 (N_5547,N_3910,N_2921);
and U5548 (N_5548,N_3010,N_3039);
nand U5549 (N_5549,N_2545,N_2410);
nor U5550 (N_5550,N_3985,N_2132);
or U5551 (N_5551,N_3676,N_2772);
and U5552 (N_5552,N_3876,N_3721);
or U5553 (N_5553,N_2341,N_3627);
nand U5554 (N_5554,N_2002,N_3557);
nor U5555 (N_5555,N_2074,N_2086);
nor U5556 (N_5556,N_3763,N_2522);
nand U5557 (N_5557,N_3893,N_3889);
nor U5558 (N_5558,N_3814,N_3344);
and U5559 (N_5559,N_2378,N_3147);
and U5560 (N_5560,N_3285,N_2607);
or U5561 (N_5561,N_2427,N_3918);
or U5562 (N_5562,N_3188,N_2160);
and U5563 (N_5563,N_2140,N_2110);
nor U5564 (N_5564,N_3111,N_2447);
xor U5565 (N_5565,N_3663,N_3328);
nand U5566 (N_5566,N_2105,N_2529);
nor U5567 (N_5567,N_2506,N_2316);
nand U5568 (N_5568,N_2295,N_3580);
nor U5569 (N_5569,N_3296,N_2413);
and U5570 (N_5570,N_2815,N_2166);
and U5571 (N_5571,N_2383,N_2774);
nand U5572 (N_5572,N_2938,N_3537);
nor U5573 (N_5573,N_2269,N_2628);
nor U5574 (N_5574,N_3279,N_3395);
nand U5575 (N_5575,N_3915,N_3113);
or U5576 (N_5576,N_2110,N_3873);
nor U5577 (N_5577,N_3611,N_3294);
or U5578 (N_5578,N_2941,N_3120);
and U5579 (N_5579,N_3191,N_3850);
nor U5580 (N_5580,N_3839,N_2198);
nand U5581 (N_5581,N_3205,N_2250);
nand U5582 (N_5582,N_3115,N_2022);
nand U5583 (N_5583,N_3525,N_3739);
nor U5584 (N_5584,N_2319,N_2878);
and U5585 (N_5585,N_2142,N_2831);
nand U5586 (N_5586,N_3244,N_2963);
nand U5587 (N_5587,N_3284,N_3171);
and U5588 (N_5588,N_3925,N_2929);
nand U5589 (N_5589,N_3508,N_3250);
nand U5590 (N_5590,N_2598,N_2801);
and U5591 (N_5591,N_2429,N_3819);
nor U5592 (N_5592,N_2733,N_2282);
and U5593 (N_5593,N_2141,N_3995);
and U5594 (N_5594,N_3062,N_2979);
or U5595 (N_5595,N_2280,N_2979);
nand U5596 (N_5596,N_3797,N_2290);
nor U5597 (N_5597,N_2549,N_2319);
or U5598 (N_5598,N_2167,N_2772);
and U5599 (N_5599,N_3189,N_3076);
or U5600 (N_5600,N_3407,N_2206);
or U5601 (N_5601,N_3132,N_3399);
and U5602 (N_5602,N_2620,N_3339);
nor U5603 (N_5603,N_2985,N_3929);
and U5604 (N_5604,N_3009,N_3688);
nand U5605 (N_5605,N_3111,N_2496);
and U5606 (N_5606,N_3981,N_2250);
and U5607 (N_5607,N_3662,N_2622);
or U5608 (N_5608,N_2050,N_3791);
xor U5609 (N_5609,N_2658,N_3689);
and U5610 (N_5610,N_2462,N_3792);
xnor U5611 (N_5611,N_3028,N_3074);
and U5612 (N_5612,N_2358,N_2107);
nor U5613 (N_5613,N_2717,N_3834);
and U5614 (N_5614,N_3106,N_2585);
nand U5615 (N_5615,N_2593,N_3725);
nor U5616 (N_5616,N_3971,N_2967);
or U5617 (N_5617,N_3532,N_3124);
or U5618 (N_5618,N_2530,N_3638);
or U5619 (N_5619,N_2529,N_3048);
or U5620 (N_5620,N_2495,N_3419);
and U5621 (N_5621,N_2640,N_3587);
and U5622 (N_5622,N_3027,N_2319);
nor U5623 (N_5623,N_2650,N_2642);
nand U5624 (N_5624,N_2911,N_2820);
or U5625 (N_5625,N_2339,N_2505);
and U5626 (N_5626,N_3372,N_2527);
nand U5627 (N_5627,N_3640,N_3587);
and U5628 (N_5628,N_2576,N_3513);
xor U5629 (N_5629,N_3160,N_2780);
or U5630 (N_5630,N_2943,N_3306);
nor U5631 (N_5631,N_3026,N_2240);
nor U5632 (N_5632,N_3604,N_2611);
nand U5633 (N_5633,N_2499,N_3433);
or U5634 (N_5634,N_3681,N_3787);
or U5635 (N_5635,N_3689,N_2378);
or U5636 (N_5636,N_2666,N_3453);
or U5637 (N_5637,N_2091,N_2298);
nor U5638 (N_5638,N_3930,N_3398);
nor U5639 (N_5639,N_3657,N_3079);
or U5640 (N_5640,N_3036,N_2891);
or U5641 (N_5641,N_3598,N_2180);
and U5642 (N_5642,N_3288,N_2130);
and U5643 (N_5643,N_2444,N_2981);
or U5644 (N_5644,N_2182,N_3065);
xor U5645 (N_5645,N_3871,N_2847);
or U5646 (N_5646,N_2695,N_2085);
or U5647 (N_5647,N_3934,N_2162);
nand U5648 (N_5648,N_3422,N_3079);
or U5649 (N_5649,N_3393,N_3715);
nor U5650 (N_5650,N_2104,N_2211);
nand U5651 (N_5651,N_3657,N_2617);
nor U5652 (N_5652,N_2548,N_2468);
and U5653 (N_5653,N_2133,N_2136);
or U5654 (N_5654,N_2006,N_2020);
and U5655 (N_5655,N_2293,N_3612);
nand U5656 (N_5656,N_2379,N_2153);
and U5657 (N_5657,N_2559,N_2274);
nor U5658 (N_5658,N_3816,N_2344);
nor U5659 (N_5659,N_2604,N_2287);
nor U5660 (N_5660,N_3730,N_2697);
and U5661 (N_5661,N_3458,N_3280);
or U5662 (N_5662,N_3495,N_3509);
and U5663 (N_5663,N_3191,N_2416);
or U5664 (N_5664,N_3451,N_2985);
nor U5665 (N_5665,N_3931,N_3504);
or U5666 (N_5666,N_2552,N_3557);
nor U5667 (N_5667,N_2386,N_2644);
or U5668 (N_5668,N_2793,N_2379);
nor U5669 (N_5669,N_3636,N_2956);
nor U5670 (N_5670,N_2412,N_2762);
or U5671 (N_5671,N_3513,N_3591);
and U5672 (N_5672,N_3626,N_2764);
or U5673 (N_5673,N_2436,N_3792);
nand U5674 (N_5674,N_3076,N_3632);
nor U5675 (N_5675,N_3513,N_3320);
and U5676 (N_5676,N_2578,N_3699);
or U5677 (N_5677,N_3779,N_3360);
nor U5678 (N_5678,N_2304,N_3402);
or U5679 (N_5679,N_2839,N_3212);
nand U5680 (N_5680,N_2242,N_3156);
nor U5681 (N_5681,N_3657,N_2504);
and U5682 (N_5682,N_3851,N_2616);
and U5683 (N_5683,N_3256,N_3569);
and U5684 (N_5684,N_3161,N_3652);
nand U5685 (N_5685,N_2138,N_3981);
nor U5686 (N_5686,N_3168,N_3233);
nor U5687 (N_5687,N_3498,N_2633);
xor U5688 (N_5688,N_3526,N_3365);
nand U5689 (N_5689,N_3597,N_3051);
nor U5690 (N_5690,N_3413,N_3348);
or U5691 (N_5691,N_2199,N_2945);
nor U5692 (N_5692,N_3952,N_2460);
nor U5693 (N_5693,N_3886,N_2609);
or U5694 (N_5694,N_2552,N_2369);
or U5695 (N_5695,N_2961,N_3394);
nand U5696 (N_5696,N_3570,N_3009);
or U5697 (N_5697,N_3737,N_2926);
nand U5698 (N_5698,N_3004,N_3606);
and U5699 (N_5699,N_2653,N_3181);
and U5700 (N_5700,N_3824,N_3474);
or U5701 (N_5701,N_3733,N_2018);
xor U5702 (N_5702,N_2072,N_3933);
or U5703 (N_5703,N_2599,N_3073);
and U5704 (N_5704,N_3250,N_3477);
or U5705 (N_5705,N_2309,N_2978);
xor U5706 (N_5706,N_2618,N_3966);
nand U5707 (N_5707,N_3877,N_2176);
and U5708 (N_5708,N_3577,N_3512);
nor U5709 (N_5709,N_3912,N_2917);
nor U5710 (N_5710,N_2866,N_2794);
or U5711 (N_5711,N_2277,N_3467);
nand U5712 (N_5712,N_3925,N_3203);
nor U5713 (N_5713,N_2849,N_3582);
and U5714 (N_5714,N_3789,N_2748);
nand U5715 (N_5715,N_2470,N_3659);
nand U5716 (N_5716,N_3641,N_3343);
nand U5717 (N_5717,N_2589,N_2699);
or U5718 (N_5718,N_3159,N_2411);
nor U5719 (N_5719,N_2078,N_3755);
or U5720 (N_5720,N_3129,N_2634);
nand U5721 (N_5721,N_3600,N_2599);
nor U5722 (N_5722,N_2865,N_3838);
or U5723 (N_5723,N_2105,N_2709);
nand U5724 (N_5724,N_2584,N_3199);
or U5725 (N_5725,N_3733,N_3722);
nand U5726 (N_5726,N_3610,N_3735);
or U5727 (N_5727,N_3001,N_3571);
and U5728 (N_5728,N_3879,N_3191);
nor U5729 (N_5729,N_2619,N_2745);
or U5730 (N_5730,N_2694,N_3751);
or U5731 (N_5731,N_3305,N_2248);
and U5732 (N_5732,N_3832,N_3661);
or U5733 (N_5733,N_2577,N_2554);
and U5734 (N_5734,N_3405,N_3752);
nand U5735 (N_5735,N_2046,N_3730);
or U5736 (N_5736,N_3824,N_3243);
nand U5737 (N_5737,N_3038,N_2824);
nand U5738 (N_5738,N_2513,N_3126);
and U5739 (N_5739,N_2734,N_3155);
or U5740 (N_5740,N_3555,N_2685);
nand U5741 (N_5741,N_2848,N_3027);
or U5742 (N_5742,N_3173,N_2362);
or U5743 (N_5743,N_2101,N_3487);
nand U5744 (N_5744,N_3821,N_2273);
nor U5745 (N_5745,N_2264,N_3450);
nand U5746 (N_5746,N_3551,N_2228);
and U5747 (N_5747,N_3227,N_2121);
nand U5748 (N_5748,N_2597,N_2765);
or U5749 (N_5749,N_3552,N_3419);
or U5750 (N_5750,N_2197,N_2427);
nor U5751 (N_5751,N_3088,N_2007);
nand U5752 (N_5752,N_3358,N_2320);
nand U5753 (N_5753,N_3073,N_2749);
or U5754 (N_5754,N_3706,N_3481);
nand U5755 (N_5755,N_3925,N_2321);
nor U5756 (N_5756,N_2698,N_2346);
or U5757 (N_5757,N_2358,N_2905);
or U5758 (N_5758,N_2121,N_2979);
or U5759 (N_5759,N_2707,N_2408);
nand U5760 (N_5760,N_3204,N_3386);
or U5761 (N_5761,N_2102,N_2715);
nor U5762 (N_5762,N_2051,N_3018);
and U5763 (N_5763,N_3421,N_3985);
or U5764 (N_5764,N_2182,N_2731);
nor U5765 (N_5765,N_2872,N_3366);
nor U5766 (N_5766,N_3457,N_2918);
and U5767 (N_5767,N_3922,N_3740);
and U5768 (N_5768,N_2805,N_2378);
nor U5769 (N_5769,N_2962,N_2183);
nor U5770 (N_5770,N_2252,N_3484);
and U5771 (N_5771,N_2966,N_3377);
and U5772 (N_5772,N_2171,N_2652);
or U5773 (N_5773,N_3339,N_3220);
and U5774 (N_5774,N_2815,N_2165);
or U5775 (N_5775,N_2029,N_3052);
or U5776 (N_5776,N_2987,N_3770);
nand U5777 (N_5777,N_2726,N_2785);
or U5778 (N_5778,N_3963,N_2298);
or U5779 (N_5779,N_2705,N_2357);
nor U5780 (N_5780,N_3623,N_3749);
nand U5781 (N_5781,N_3448,N_2601);
or U5782 (N_5782,N_2271,N_2559);
and U5783 (N_5783,N_3053,N_2136);
nor U5784 (N_5784,N_2666,N_3560);
nor U5785 (N_5785,N_3426,N_3690);
or U5786 (N_5786,N_2268,N_3507);
nor U5787 (N_5787,N_2076,N_2775);
or U5788 (N_5788,N_2628,N_2405);
nor U5789 (N_5789,N_2599,N_2028);
nand U5790 (N_5790,N_2079,N_3515);
or U5791 (N_5791,N_2848,N_2733);
nand U5792 (N_5792,N_2762,N_3469);
nand U5793 (N_5793,N_3632,N_2742);
and U5794 (N_5794,N_3808,N_2645);
and U5795 (N_5795,N_2503,N_2839);
and U5796 (N_5796,N_2285,N_2152);
nand U5797 (N_5797,N_2496,N_2014);
or U5798 (N_5798,N_3309,N_3562);
and U5799 (N_5799,N_3042,N_3337);
nor U5800 (N_5800,N_2265,N_3974);
or U5801 (N_5801,N_2405,N_2097);
nor U5802 (N_5802,N_3228,N_3133);
or U5803 (N_5803,N_3384,N_3682);
nor U5804 (N_5804,N_2909,N_3500);
or U5805 (N_5805,N_3687,N_2146);
nor U5806 (N_5806,N_2352,N_2753);
nor U5807 (N_5807,N_3467,N_3862);
and U5808 (N_5808,N_2594,N_3668);
nor U5809 (N_5809,N_3373,N_2853);
or U5810 (N_5810,N_2248,N_2727);
nand U5811 (N_5811,N_2753,N_3067);
and U5812 (N_5812,N_2477,N_3638);
or U5813 (N_5813,N_3260,N_2436);
nor U5814 (N_5814,N_3835,N_2532);
nand U5815 (N_5815,N_3778,N_3763);
nor U5816 (N_5816,N_3824,N_2981);
nor U5817 (N_5817,N_3434,N_3842);
nand U5818 (N_5818,N_2058,N_2957);
xnor U5819 (N_5819,N_2709,N_2995);
nand U5820 (N_5820,N_3469,N_2009);
nand U5821 (N_5821,N_2878,N_2720);
and U5822 (N_5822,N_3601,N_3185);
and U5823 (N_5823,N_2653,N_2261);
or U5824 (N_5824,N_3325,N_3863);
and U5825 (N_5825,N_2929,N_2817);
or U5826 (N_5826,N_2104,N_2222);
nor U5827 (N_5827,N_2781,N_2337);
nor U5828 (N_5828,N_2513,N_3562);
nand U5829 (N_5829,N_3821,N_2594);
nand U5830 (N_5830,N_3405,N_2078);
nand U5831 (N_5831,N_3099,N_2505);
nor U5832 (N_5832,N_2813,N_3627);
nor U5833 (N_5833,N_2691,N_2747);
and U5834 (N_5834,N_3734,N_3025);
nand U5835 (N_5835,N_3030,N_3618);
nor U5836 (N_5836,N_2380,N_3778);
and U5837 (N_5837,N_3238,N_2787);
nor U5838 (N_5838,N_2672,N_3337);
nor U5839 (N_5839,N_3069,N_2589);
nand U5840 (N_5840,N_3393,N_3985);
nand U5841 (N_5841,N_2439,N_2777);
nor U5842 (N_5842,N_2361,N_3821);
and U5843 (N_5843,N_2533,N_3882);
nor U5844 (N_5844,N_3906,N_3090);
or U5845 (N_5845,N_3586,N_2455);
and U5846 (N_5846,N_2920,N_3799);
nor U5847 (N_5847,N_3251,N_3562);
nor U5848 (N_5848,N_3111,N_2810);
nor U5849 (N_5849,N_2980,N_2923);
nor U5850 (N_5850,N_2208,N_3039);
and U5851 (N_5851,N_2138,N_2044);
nor U5852 (N_5852,N_2264,N_2384);
nand U5853 (N_5853,N_3796,N_2741);
or U5854 (N_5854,N_3501,N_3850);
and U5855 (N_5855,N_2502,N_2204);
and U5856 (N_5856,N_2969,N_3117);
and U5857 (N_5857,N_3527,N_2692);
xnor U5858 (N_5858,N_3298,N_2682);
nor U5859 (N_5859,N_3645,N_3699);
nand U5860 (N_5860,N_3312,N_3809);
or U5861 (N_5861,N_3976,N_3136);
and U5862 (N_5862,N_3424,N_3968);
and U5863 (N_5863,N_2954,N_2973);
or U5864 (N_5864,N_2807,N_3556);
nor U5865 (N_5865,N_2308,N_3138);
and U5866 (N_5866,N_3564,N_3721);
or U5867 (N_5867,N_3304,N_2766);
nand U5868 (N_5868,N_2906,N_3332);
nor U5869 (N_5869,N_3749,N_3022);
nand U5870 (N_5870,N_3532,N_2541);
nand U5871 (N_5871,N_3792,N_3741);
and U5872 (N_5872,N_3930,N_3410);
or U5873 (N_5873,N_3058,N_3786);
nand U5874 (N_5874,N_3649,N_3566);
nor U5875 (N_5875,N_3426,N_3643);
and U5876 (N_5876,N_2206,N_3965);
nor U5877 (N_5877,N_2461,N_2700);
and U5878 (N_5878,N_2671,N_2393);
nand U5879 (N_5879,N_3741,N_3965);
or U5880 (N_5880,N_2022,N_2646);
or U5881 (N_5881,N_2807,N_3848);
or U5882 (N_5882,N_3580,N_2253);
nor U5883 (N_5883,N_2822,N_2142);
or U5884 (N_5884,N_2947,N_2167);
and U5885 (N_5885,N_2007,N_2244);
and U5886 (N_5886,N_3370,N_3758);
nor U5887 (N_5887,N_3400,N_2448);
and U5888 (N_5888,N_3729,N_3659);
or U5889 (N_5889,N_2962,N_2890);
and U5890 (N_5890,N_3224,N_2334);
or U5891 (N_5891,N_3969,N_3230);
and U5892 (N_5892,N_3054,N_3009);
nor U5893 (N_5893,N_2394,N_2693);
nor U5894 (N_5894,N_2074,N_2505);
and U5895 (N_5895,N_3033,N_2089);
nand U5896 (N_5896,N_3237,N_2211);
nor U5897 (N_5897,N_3262,N_2673);
nor U5898 (N_5898,N_3873,N_3307);
or U5899 (N_5899,N_2318,N_2725);
or U5900 (N_5900,N_2314,N_3241);
and U5901 (N_5901,N_2560,N_3270);
and U5902 (N_5902,N_3721,N_2951);
or U5903 (N_5903,N_3558,N_2608);
nand U5904 (N_5904,N_2320,N_2566);
and U5905 (N_5905,N_2311,N_3762);
and U5906 (N_5906,N_2889,N_3292);
nand U5907 (N_5907,N_2363,N_3881);
or U5908 (N_5908,N_2631,N_3252);
nor U5909 (N_5909,N_3429,N_3877);
or U5910 (N_5910,N_3603,N_2293);
and U5911 (N_5911,N_2595,N_2077);
nand U5912 (N_5912,N_2175,N_2537);
nor U5913 (N_5913,N_2093,N_2831);
nand U5914 (N_5914,N_3909,N_2501);
nor U5915 (N_5915,N_2224,N_2953);
nand U5916 (N_5916,N_2215,N_3836);
nand U5917 (N_5917,N_3393,N_2687);
nand U5918 (N_5918,N_3086,N_3901);
nor U5919 (N_5919,N_2949,N_3763);
and U5920 (N_5920,N_2437,N_2983);
or U5921 (N_5921,N_3149,N_3553);
nand U5922 (N_5922,N_3426,N_2616);
nand U5923 (N_5923,N_3764,N_3685);
and U5924 (N_5924,N_3882,N_2891);
nand U5925 (N_5925,N_3475,N_2744);
nor U5926 (N_5926,N_3954,N_2671);
nand U5927 (N_5927,N_2498,N_2660);
nor U5928 (N_5928,N_2413,N_2102);
and U5929 (N_5929,N_2943,N_3229);
nand U5930 (N_5930,N_3034,N_3436);
or U5931 (N_5931,N_3838,N_3821);
or U5932 (N_5932,N_2490,N_3531);
and U5933 (N_5933,N_2416,N_3119);
and U5934 (N_5934,N_2170,N_3611);
or U5935 (N_5935,N_2162,N_3066);
and U5936 (N_5936,N_2978,N_2751);
nor U5937 (N_5937,N_2247,N_2725);
and U5938 (N_5938,N_3098,N_2764);
or U5939 (N_5939,N_2767,N_2908);
nor U5940 (N_5940,N_2649,N_3010);
and U5941 (N_5941,N_2502,N_3511);
and U5942 (N_5942,N_3518,N_2548);
nor U5943 (N_5943,N_2565,N_2219);
and U5944 (N_5944,N_3022,N_2255);
and U5945 (N_5945,N_3312,N_3471);
or U5946 (N_5946,N_3857,N_3741);
or U5947 (N_5947,N_3429,N_3662);
or U5948 (N_5948,N_2145,N_2465);
nor U5949 (N_5949,N_2586,N_3200);
and U5950 (N_5950,N_2657,N_2021);
nand U5951 (N_5951,N_3506,N_3842);
or U5952 (N_5952,N_3928,N_3620);
nand U5953 (N_5953,N_2934,N_3054);
nand U5954 (N_5954,N_2132,N_2584);
and U5955 (N_5955,N_3661,N_3525);
nand U5956 (N_5956,N_2635,N_2674);
or U5957 (N_5957,N_2416,N_3781);
xor U5958 (N_5958,N_2974,N_3121);
or U5959 (N_5959,N_2110,N_2717);
nand U5960 (N_5960,N_3876,N_2975);
nor U5961 (N_5961,N_3261,N_2560);
nor U5962 (N_5962,N_3500,N_2357);
nor U5963 (N_5963,N_3821,N_3379);
nor U5964 (N_5964,N_3737,N_3100);
nand U5965 (N_5965,N_2929,N_2486);
nor U5966 (N_5966,N_2751,N_3539);
or U5967 (N_5967,N_3539,N_2256);
or U5968 (N_5968,N_3518,N_2389);
or U5969 (N_5969,N_2394,N_2515);
and U5970 (N_5970,N_3255,N_2940);
nor U5971 (N_5971,N_2577,N_2125);
or U5972 (N_5972,N_2345,N_2513);
and U5973 (N_5973,N_3820,N_2162);
and U5974 (N_5974,N_3603,N_3044);
nor U5975 (N_5975,N_3649,N_2763);
nand U5976 (N_5976,N_3583,N_2051);
nand U5977 (N_5977,N_3234,N_3555);
or U5978 (N_5978,N_3900,N_2787);
and U5979 (N_5979,N_3404,N_2021);
nor U5980 (N_5980,N_2774,N_3689);
or U5981 (N_5981,N_3346,N_2254);
nand U5982 (N_5982,N_3400,N_2860);
nor U5983 (N_5983,N_2471,N_2339);
and U5984 (N_5984,N_3403,N_3141);
or U5985 (N_5985,N_2002,N_3051);
nand U5986 (N_5986,N_3209,N_2570);
and U5987 (N_5987,N_2925,N_2011);
nand U5988 (N_5988,N_3161,N_3020);
and U5989 (N_5989,N_2746,N_3024);
nand U5990 (N_5990,N_2902,N_2994);
nor U5991 (N_5991,N_3270,N_2170);
nand U5992 (N_5992,N_3981,N_3680);
or U5993 (N_5993,N_3531,N_3546);
nor U5994 (N_5994,N_3300,N_2329);
xor U5995 (N_5995,N_3507,N_2463);
and U5996 (N_5996,N_3145,N_2203);
and U5997 (N_5997,N_2002,N_3693);
nand U5998 (N_5998,N_2369,N_3232);
nand U5999 (N_5999,N_2125,N_2962);
nor U6000 (N_6000,N_5233,N_5547);
or U6001 (N_6001,N_4762,N_5357);
and U6002 (N_6002,N_5155,N_5039);
and U6003 (N_6003,N_5344,N_5782);
or U6004 (N_6004,N_4819,N_5127);
or U6005 (N_6005,N_4879,N_5413);
nor U6006 (N_6006,N_4282,N_5460);
nor U6007 (N_6007,N_4798,N_4694);
nor U6008 (N_6008,N_5142,N_5154);
and U6009 (N_6009,N_4579,N_4485);
and U6010 (N_6010,N_5196,N_5482);
nand U6011 (N_6011,N_4179,N_5559);
nand U6012 (N_6012,N_5485,N_5377);
or U6013 (N_6013,N_4688,N_5809);
or U6014 (N_6014,N_4086,N_4549);
or U6015 (N_6015,N_4994,N_4202);
and U6016 (N_6016,N_5964,N_5544);
nor U6017 (N_6017,N_4333,N_4831);
nand U6018 (N_6018,N_5991,N_4397);
nand U6019 (N_6019,N_5268,N_5309);
nand U6020 (N_6020,N_5030,N_4175);
nand U6021 (N_6021,N_5402,N_5669);
nor U6022 (N_6022,N_5063,N_4371);
nor U6023 (N_6023,N_5525,N_4207);
nor U6024 (N_6024,N_5845,N_4035);
nor U6025 (N_6025,N_4536,N_4808);
nor U6026 (N_6026,N_4319,N_4356);
nor U6027 (N_6027,N_5683,N_5311);
nor U6028 (N_6028,N_5748,N_5803);
and U6029 (N_6029,N_4653,N_4911);
nand U6030 (N_6030,N_4242,N_4028);
nand U6031 (N_6031,N_4865,N_4968);
or U6032 (N_6032,N_5033,N_4575);
and U6033 (N_6033,N_5812,N_4592);
nand U6034 (N_6034,N_5625,N_4064);
nand U6035 (N_6035,N_5407,N_5631);
nand U6036 (N_6036,N_4238,N_4609);
or U6037 (N_6037,N_4452,N_4613);
or U6038 (N_6038,N_4499,N_5215);
or U6039 (N_6039,N_4862,N_4644);
or U6040 (N_6040,N_4039,N_5581);
or U6041 (N_6041,N_5056,N_4321);
or U6042 (N_6042,N_5840,N_4413);
nand U6043 (N_6043,N_5347,N_5982);
xor U6044 (N_6044,N_5259,N_5785);
nor U6045 (N_6045,N_4334,N_4110);
and U6046 (N_6046,N_4813,N_4699);
or U6047 (N_6047,N_5073,N_4636);
and U6048 (N_6048,N_5510,N_5505);
or U6049 (N_6049,N_5206,N_4287);
or U6050 (N_6050,N_5834,N_4511);
nor U6051 (N_6051,N_5754,N_5476);
or U6052 (N_6052,N_4446,N_4915);
nor U6053 (N_6053,N_5511,N_4978);
and U6054 (N_6054,N_4317,N_4444);
or U6055 (N_6055,N_5284,N_4366);
nor U6056 (N_6056,N_4670,N_4427);
nor U6057 (N_6057,N_4059,N_4336);
nor U6058 (N_6058,N_4948,N_4729);
nand U6059 (N_6059,N_5151,N_4061);
nor U6060 (N_6060,N_5839,N_5288);
or U6061 (N_6061,N_5883,N_4363);
nand U6062 (N_6062,N_4735,N_5540);
nor U6063 (N_6063,N_5700,N_5159);
and U6064 (N_6064,N_5121,N_5753);
xor U6065 (N_6065,N_5863,N_5003);
and U6066 (N_6066,N_4558,N_4628);
and U6067 (N_6067,N_5324,N_5022);
and U6068 (N_6068,N_4290,N_5950);
and U6069 (N_6069,N_5795,N_4426);
nand U6070 (N_6070,N_4781,N_5008);
or U6071 (N_6071,N_4203,N_4137);
nand U6072 (N_6072,N_4351,N_5287);
nand U6073 (N_6073,N_4461,N_5556);
or U6074 (N_6074,N_4856,N_4313);
nand U6075 (N_6075,N_4494,N_5943);
and U6076 (N_6076,N_5780,N_5589);
or U6077 (N_6077,N_4042,N_4600);
or U6078 (N_6078,N_5112,N_5874);
nand U6079 (N_6079,N_4706,N_5423);
nand U6080 (N_6080,N_5549,N_4765);
and U6081 (N_6081,N_4764,N_4986);
and U6082 (N_6082,N_4314,N_4920);
nor U6083 (N_6083,N_5374,N_5786);
nor U6084 (N_6084,N_5571,N_5273);
and U6085 (N_6085,N_4622,N_5679);
or U6086 (N_6086,N_4298,N_5521);
or U6087 (N_6087,N_4142,N_5147);
and U6088 (N_6088,N_5739,N_4153);
nand U6089 (N_6089,N_5368,N_5997);
or U6090 (N_6090,N_5531,N_4068);
or U6091 (N_6091,N_4014,N_5441);
or U6092 (N_6092,N_4106,N_5418);
and U6093 (N_6093,N_4795,N_5322);
nand U6094 (N_6094,N_5980,N_5861);
or U6095 (N_6095,N_5468,N_5904);
or U6096 (N_6096,N_5977,N_4256);
or U6097 (N_6097,N_5255,N_4807);
nand U6098 (N_6098,N_4604,N_4825);
and U6099 (N_6099,N_5775,N_5299);
or U6100 (N_6100,N_4777,N_4253);
and U6101 (N_6101,N_4851,N_5504);
and U6102 (N_6102,N_4265,N_5434);
xnor U6103 (N_6103,N_5937,N_5075);
or U6104 (N_6104,N_5929,N_4353);
and U6105 (N_6105,N_4890,N_4416);
nand U6106 (N_6106,N_4800,N_5973);
nand U6107 (N_6107,N_5432,N_4013);
or U6108 (N_6108,N_4180,N_5626);
nand U6109 (N_6109,N_5506,N_4517);
nand U6110 (N_6110,N_4547,N_5523);
or U6111 (N_6111,N_5331,N_5602);
nand U6112 (N_6112,N_5466,N_5794);
nand U6113 (N_6113,N_4633,N_5960);
and U6114 (N_6114,N_5806,N_5566);
and U6115 (N_6115,N_4476,N_4933);
and U6116 (N_6116,N_4286,N_4006);
nand U6117 (N_6117,N_5193,N_5723);
nand U6118 (N_6118,N_5718,N_5009);
nand U6119 (N_6119,N_5366,N_5736);
nand U6120 (N_6120,N_5333,N_5171);
nor U6121 (N_6121,N_5616,N_4681);
and U6122 (N_6122,N_4501,N_4742);
nor U6123 (N_6123,N_4508,N_5918);
nand U6124 (N_6124,N_4462,N_4026);
nand U6125 (N_6125,N_5232,N_4768);
and U6126 (N_6126,N_4418,N_5978);
nand U6127 (N_6127,N_5647,N_4659);
and U6128 (N_6128,N_4873,N_4896);
nor U6129 (N_6129,N_5724,N_5654);
or U6130 (N_6130,N_4977,N_4231);
and U6131 (N_6131,N_5406,N_4975);
nand U6132 (N_6132,N_4724,N_4770);
nor U6133 (N_6133,N_5188,N_5939);
nor U6134 (N_6134,N_4998,N_5446);
and U6135 (N_6135,N_5887,N_4894);
nor U6136 (N_6136,N_4664,N_5303);
nand U6137 (N_6137,N_5719,N_5797);
and U6138 (N_6138,N_5867,N_4859);
and U6139 (N_6139,N_5080,N_4956);
or U6140 (N_6140,N_5774,N_4582);
nand U6141 (N_6141,N_4845,N_4936);
and U6142 (N_6142,N_4853,N_4897);
nand U6143 (N_6143,N_5308,N_4081);
nor U6144 (N_6144,N_5732,N_5089);
nor U6145 (N_6145,N_4697,N_4837);
nand U6146 (N_6146,N_5928,N_4638);
nor U6147 (N_6147,N_5006,N_5953);
nor U6148 (N_6148,N_5038,N_5164);
xnor U6149 (N_6149,N_5551,N_5034);
nor U6150 (N_6150,N_4751,N_4545);
nor U6151 (N_6151,N_4331,N_5078);
nand U6152 (N_6152,N_5760,N_4274);
and U6153 (N_6153,N_5065,N_5479);
nor U6154 (N_6154,N_4297,N_5126);
or U6155 (N_6155,N_4273,N_4468);
or U6156 (N_6156,N_5143,N_5518);
and U6157 (N_6157,N_4021,N_5516);
nor U6158 (N_6158,N_4570,N_5120);
and U6159 (N_6159,N_5156,N_4224);
and U6160 (N_6160,N_5049,N_4131);
nor U6161 (N_6161,N_4560,N_4390);
nand U6162 (N_6162,N_4323,N_5614);
and U6163 (N_6163,N_5856,N_4748);
and U6164 (N_6164,N_5796,N_5742);
nor U6165 (N_6165,N_5452,N_5296);
or U6166 (N_6166,N_5409,N_4782);
xor U6167 (N_6167,N_4525,N_4861);
and U6168 (N_6168,N_4692,N_4693);
nand U6169 (N_6169,N_4191,N_5852);
xnor U6170 (N_6170,N_5059,N_4164);
nand U6171 (N_6171,N_5777,N_5588);
and U6172 (N_6172,N_4250,N_5734);
or U6173 (N_6173,N_5111,N_5575);
or U6174 (N_6174,N_5227,N_5220);
or U6175 (N_6175,N_5335,N_5998);
and U6176 (N_6176,N_4054,N_4677);
and U6177 (N_6177,N_5241,N_4025);
nor U6178 (N_6178,N_4210,N_5972);
nand U6179 (N_6179,N_4712,N_5312);
or U6180 (N_6180,N_5594,N_4587);
nand U6181 (N_6181,N_5642,N_5655);
or U6182 (N_6182,N_5539,N_4208);
or U6183 (N_6183,N_4548,N_5425);
nand U6184 (N_6184,N_5316,N_4899);
nor U6185 (N_6185,N_5408,N_4221);
nand U6186 (N_6186,N_5162,N_4473);
or U6187 (N_6187,N_4071,N_4490);
nor U6188 (N_6188,N_4996,N_4802);
or U6189 (N_6189,N_5167,N_5586);
nand U6190 (N_6190,N_5947,N_4037);
nand U6191 (N_6191,N_5955,N_5032);
and U6192 (N_6192,N_5823,N_4130);
nor U6193 (N_6193,N_5590,N_5661);
and U6194 (N_6194,N_4611,N_4305);
and U6195 (N_6195,N_5744,N_5873);
or U6196 (N_6196,N_5985,N_4119);
or U6197 (N_6197,N_4518,N_5779);
and U6198 (N_6198,N_4612,N_5414);
and U6199 (N_6199,N_4198,N_5858);
and U6200 (N_6200,N_4451,N_4731);
and U6201 (N_6201,N_5798,N_5680);
nand U6202 (N_6202,N_5005,N_4687);
xnor U6203 (N_6203,N_5150,N_4541);
nand U6204 (N_6204,N_4176,N_4821);
nor U6205 (N_6205,N_4085,N_4151);
nor U6206 (N_6206,N_4120,N_5440);
nand U6207 (N_6207,N_5692,N_4850);
nand U6208 (N_6208,N_4438,N_5389);
nand U6209 (N_6209,N_4673,N_4597);
or U6210 (N_6210,N_5189,N_5971);
nand U6211 (N_6211,N_5424,N_4236);
and U6212 (N_6212,N_5119,N_5144);
nand U6213 (N_6213,N_4520,N_4095);
nand U6214 (N_6214,N_5848,N_4874);
and U6215 (N_6215,N_4190,N_4369);
or U6216 (N_6216,N_5292,N_4642);
and U6217 (N_6217,N_5745,N_5791);
nand U6218 (N_6218,N_5604,N_5580);
and U6219 (N_6219,N_4489,N_5496);
and U6220 (N_6220,N_4146,N_5054);
and U6221 (N_6221,N_4552,N_4041);
or U6222 (N_6222,N_5532,N_5743);
or U6223 (N_6223,N_5562,N_4109);
nor U6224 (N_6224,N_4602,N_5857);
nor U6225 (N_6225,N_4820,N_5050);
or U6226 (N_6226,N_4531,N_5271);
nand U6227 (N_6227,N_4684,N_5223);
nand U6228 (N_6228,N_5727,N_5746);
nor U6229 (N_6229,N_5272,N_4185);
nor U6230 (N_6230,N_5134,N_5105);
or U6231 (N_6231,N_4421,N_5174);
nand U6232 (N_6232,N_4240,N_4206);
nand U6233 (N_6233,N_5543,N_4078);
nor U6234 (N_6234,N_5702,N_5367);
or U6235 (N_6235,N_4778,N_4395);
xor U6236 (N_6236,N_4268,N_5417);
and U6237 (N_6237,N_4754,N_5689);
nand U6238 (N_6238,N_5841,N_4847);
nand U6239 (N_6239,N_5278,N_5252);
or U6240 (N_6240,N_4056,N_5747);
and U6241 (N_6241,N_4783,N_5137);
nor U6242 (N_6242,N_4004,N_5662);
nand U6243 (N_6243,N_4848,N_5709);
nor U6244 (N_6244,N_4671,N_5045);
nand U6245 (N_6245,N_5457,N_4789);
nor U6246 (N_6246,N_5190,N_5900);
nor U6247 (N_6247,N_5920,N_5690);
or U6248 (N_6248,N_4099,N_4625);
nand U6249 (N_6249,N_4507,N_5618);
and U6250 (N_6250,N_5988,N_4551);
nor U6251 (N_6251,N_5691,N_5014);
or U6252 (N_6252,N_5450,N_5866);
nor U6253 (N_6253,N_5847,N_4347);
nand U6254 (N_6254,N_5390,N_5088);
and U6255 (N_6255,N_5563,N_4741);
nand U6256 (N_6256,N_5429,N_5258);
or U6257 (N_6257,N_5433,N_4219);
nand U6258 (N_6258,N_4855,N_4954);
and U6259 (N_6259,N_4784,N_5875);
and U6260 (N_6260,N_5491,N_5936);
or U6261 (N_6261,N_4901,N_5375);
nor U6262 (N_6262,N_5577,N_4247);
nor U6263 (N_6263,N_4965,N_5788);
nor U6264 (N_6264,N_5400,N_5350);
nor U6265 (N_6265,N_5097,N_5674);
nand U6266 (N_6266,N_4048,N_4230);
and U6267 (N_6267,N_4415,N_4150);
and U6268 (N_6268,N_5676,N_5619);
nand U6269 (N_6269,N_5109,N_4569);
nand U6270 (N_6270,N_4912,N_5229);
or U6271 (N_6271,N_5909,N_4118);
and U6272 (N_6272,N_5698,N_5401);
nand U6273 (N_6273,N_5200,N_5093);
and U6274 (N_6274,N_4701,N_5031);
nand U6275 (N_6275,N_4393,N_4944);
nor U6276 (N_6276,N_5023,N_4133);
nand U6277 (N_6277,N_5094,N_4196);
or U6278 (N_6278,N_4074,N_4985);
or U6279 (N_6279,N_5289,N_5285);
and U6280 (N_6280,N_4477,N_4704);
xnor U6281 (N_6281,N_4621,N_5872);
nor U6282 (N_6282,N_5565,N_4630);
nand U6283 (N_6283,N_4683,N_4033);
or U6284 (N_6284,N_4480,N_5851);
or U6285 (N_6285,N_5339,N_5697);
or U6286 (N_6286,N_5512,N_5952);
or U6287 (N_6287,N_4112,N_4339);
nand U6288 (N_6288,N_5475,N_5761);
nor U6289 (N_6289,N_4727,N_5069);
nor U6290 (N_6290,N_4358,N_5981);
or U6291 (N_6291,N_4771,N_5079);
or U6292 (N_6292,N_4018,N_4824);
nand U6293 (N_6293,N_5751,N_4195);
or U6294 (N_6294,N_4102,N_4918);
or U6295 (N_6295,N_4939,N_5705);
or U6296 (N_6296,N_5870,N_4445);
nand U6297 (N_6297,N_5681,N_4893);
nor U6298 (N_6298,N_5963,N_5437);
nor U6299 (N_6299,N_4870,N_5314);
and U6300 (N_6300,N_5325,N_4010);
and U6301 (N_6301,N_5684,N_5945);
nand U6302 (N_6302,N_5204,N_5520);
nand U6303 (N_6303,N_5387,N_5941);
nor U6304 (N_6304,N_5462,N_4315);
and U6305 (N_6305,N_4093,N_4182);
nand U6306 (N_6306,N_5508,N_5652);
nor U6307 (N_6307,N_4001,N_4809);
nor U6308 (N_6308,N_5092,N_5608);
nand U6309 (N_6309,N_4844,N_5996);
nor U6310 (N_6310,N_5102,N_5301);
or U6311 (N_6311,N_4411,N_5778);
nand U6312 (N_6312,N_4482,N_4329);
or U6313 (N_6313,N_5793,N_4378);
nand U6314 (N_6314,N_5694,N_5878);
nor U6315 (N_6315,N_5965,N_5313);
nor U6316 (N_6316,N_4752,N_5716);
nor U6317 (N_6317,N_4005,N_5923);
nand U6318 (N_6318,N_4318,N_5246);
nand U6319 (N_6319,N_4410,N_5587);
nor U6320 (N_6320,N_4303,N_4690);
nor U6321 (N_6321,N_4386,N_4891);
nand U6322 (N_6322,N_4733,N_4121);
nor U6323 (N_6323,N_5430,N_5884);
and U6324 (N_6324,N_5323,N_5671);
nor U6325 (N_6325,N_5624,N_5098);
and U6326 (N_6326,N_5037,N_5472);
nand U6327 (N_6327,N_4407,N_4738);
nor U6328 (N_6328,N_4846,N_4737);
nor U6329 (N_6329,N_4326,N_4740);
or U6330 (N_6330,N_4361,N_5805);
and U6331 (N_6331,N_5320,N_5051);
nand U6332 (N_6332,N_5893,N_4436);
nor U6333 (N_6333,N_5113,N_4437);
nor U6334 (N_6334,N_5758,N_5058);
or U6335 (N_6335,N_4324,N_5264);
or U6336 (N_6336,N_5293,N_4646);
or U6337 (N_6337,N_4254,N_4383);
or U6338 (N_6338,N_5769,N_4201);
or U6339 (N_6339,N_4239,N_5582);
xnor U6340 (N_6340,N_5628,N_4029);
nand U6341 (N_6341,N_5244,N_4345);
and U6342 (N_6342,N_5849,N_4730);
nand U6343 (N_6343,N_4047,N_5426);
nand U6344 (N_6344,N_5012,N_4365);
xnor U6345 (N_6345,N_4199,N_5627);
xnor U6346 (N_6346,N_4745,N_4101);
nand U6347 (N_6347,N_5818,N_4755);
and U6348 (N_6348,N_4760,N_5186);
nor U6349 (N_6349,N_4550,N_5890);
nor U6350 (N_6350,N_5819,N_4011);
nand U6351 (N_6351,N_4759,N_5047);
nand U6352 (N_6352,N_5275,N_4951);
or U6353 (N_6353,N_5052,N_4949);
xor U6354 (N_6354,N_4953,N_4065);
and U6355 (N_6355,N_5235,N_4617);
or U6356 (N_6356,N_5254,N_4116);
or U6357 (N_6357,N_5804,N_4373);
nand U6358 (N_6358,N_4937,N_4909);
and U6359 (N_6359,N_4398,N_4513);
nand U6360 (N_6360,N_4155,N_4934);
nand U6361 (N_6361,N_5021,N_4999);
or U6362 (N_6362,N_4493,N_5552);
nor U6363 (N_6363,N_4982,N_4259);
nand U6364 (N_6364,N_4127,N_4301);
nand U6365 (N_6365,N_5341,N_5269);
and U6366 (N_6366,N_4539,N_5926);
nor U6367 (N_6367,N_5281,N_5621);
and U6368 (N_6368,N_4655,N_5938);
nor U6369 (N_6369,N_4000,N_4063);
nor U6370 (N_6370,N_4554,N_5474);
nand U6371 (N_6371,N_4723,N_5854);
or U6372 (N_6372,N_5198,N_4362);
nor U6373 (N_6373,N_4157,N_5974);
or U6374 (N_6374,N_5166,N_4581);
or U6375 (N_6375,N_4177,N_5949);
nor U6376 (N_6376,N_5172,N_5713);
or U6377 (N_6377,N_5454,N_5427);
nor U6378 (N_6378,N_4970,N_5610);
and U6379 (N_6379,N_4328,N_5074);
and U6380 (N_6380,N_5226,N_4172);
nor U6381 (N_6381,N_5000,N_4610);
nor U6382 (N_6382,N_4432,N_4635);
nor U6383 (N_6383,N_5001,N_5675);
or U6384 (N_6384,N_4359,N_4555);
or U6385 (N_6385,N_4060,N_4838);
xor U6386 (N_6386,N_4641,N_4495);
and U6387 (N_6387,N_5930,N_4139);
nand U6388 (N_6388,N_5787,N_4586);
nand U6389 (N_6389,N_5535,N_5572);
nor U6390 (N_6390,N_5411,N_4192);
or U6391 (N_6391,N_4674,N_5799);
nor U6392 (N_6392,N_4425,N_4769);
and U6393 (N_6393,N_5574,N_5213);
or U6394 (N_6394,N_4211,N_5456);
or U6395 (N_6395,N_4491,N_5099);
nand U6396 (N_6396,N_4077,N_4966);
nor U6397 (N_6397,N_4335,N_5752);
or U6398 (N_6398,N_4459,N_4750);
and U6399 (N_6399,N_5044,N_5912);
or U6400 (N_6400,N_4352,N_5541);
or U6401 (N_6401,N_5885,N_5025);
and U6402 (N_6402,N_4827,N_5927);
or U6403 (N_6403,N_5976,N_5706);
or U6404 (N_6404,N_4027,N_4559);
and U6405 (N_6405,N_4627,N_5983);
and U6406 (N_6406,N_4036,N_5392);
or U6407 (N_6407,N_5792,N_5548);
nor U6408 (N_6408,N_4705,N_5125);
or U6409 (N_6409,N_4388,N_4618);
nor U6410 (N_6410,N_5160,N_4235);
nand U6411 (N_6411,N_5286,N_4104);
nor U6412 (N_6412,N_5763,N_4498);
nor U6413 (N_6413,N_4124,N_5494);
nand U6414 (N_6414,N_5640,N_4082);
or U6415 (N_6415,N_4910,N_4527);
nor U6416 (N_6416,N_5495,N_5877);
and U6417 (N_6417,N_5721,N_5591);
nand U6418 (N_6418,N_4608,N_4500);
or U6419 (N_6419,N_4565,N_4528);
or U6420 (N_6420,N_5236,N_4563);
or U6421 (N_6421,N_4780,N_5707);
xor U6422 (N_6422,N_4756,N_5247);
nor U6423 (N_6423,N_5886,N_5342);
and U6424 (N_6424,N_5340,N_5536);
or U6425 (N_6425,N_4216,N_4979);
or U6426 (N_6426,N_5567,N_4404);
and U6427 (N_6427,N_4981,N_4184);
and U6428 (N_6428,N_4823,N_4003);
nor U6429 (N_6429,N_5360,N_5564);
nand U6430 (N_6430,N_5224,N_5915);
nor U6431 (N_6431,N_5598,N_5528);
nand U6432 (N_6432,N_5183,N_4594);
nand U6433 (N_6433,N_5428,N_4512);
and U6434 (N_6434,N_5067,N_5944);
nand U6435 (N_6435,N_4799,N_4143);
nor U6436 (N_6436,N_5898,N_5569);
nor U6437 (N_6437,N_4430,N_4775);
or U6438 (N_6438,N_5613,N_5061);
nand U6439 (N_6439,N_5391,N_4295);
or U6440 (N_6440,N_5612,N_5659);
nor U6441 (N_6441,N_4149,N_4387);
xnor U6442 (N_6442,N_4908,N_5527);
and U6443 (N_6443,N_5816,N_5968);
and U6444 (N_6444,N_4719,N_4249);
nor U6445 (N_6445,N_5913,N_5029);
and U6446 (N_6446,N_5202,N_4412);
or U6447 (N_6447,N_4168,N_4533);
nor U6448 (N_6448,N_4080,N_5507);
and U6449 (N_6449,N_5648,N_5328);
nand U6450 (N_6450,N_4652,N_4803);
and U6451 (N_6451,N_4812,N_4877);
or U6452 (N_6452,N_5643,N_5601);
nand U6453 (N_6453,N_4504,N_4117);
and U6454 (N_6454,N_4995,N_4228);
and U6455 (N_6455,N_4876,N_4632);
or U6456 (N_6456,N_4805,N_5420);
or U6457 (N_6457,N_5573,N_5583);
or U6458 (N_6458,N_4007,N_5265);
and U6459 (N_6459,N_5864,N_5597);
nand U6460 (N_6460,N_4811,N_4220);
nand U6461 (N_6461,N_4766,N_5629);
xnor U6462 (N_6462,N_4330,N_4884);
nand U6463 (N_6463,N_5305,N_5415);
and U6464 (N_6464,N_5405,N_5934);
nor U6465 (N_6465,N_4816,N_5889);
nand U6466 (N_6466,N_4030,N_5260);
and U6467 (N_6467,N_4299,N_4349);
nor U6468 (N_6468,N_5735,N_4840);
and U6469 (N_6469,N_4648,N_4929);
nor U6470 (N_6470,N_4523,N_5942);
or U6471 (N_6471,N_4836,N_4163);
and U6472 (N_6472,N_5245,N_4159);
nand U6473 (N_6473,N_5488,N_4218);
and U6474 (N_6474,N_4538,N_5464);
and U6475 (N_6475,N_4343,N_4797);
or U6476 (N_6476,N_4928,N_4757);
or U6477 (N_6477,N_4261,N_4215);
nand U6478 (N_6478,N_4532,N_5931);
nand U6479 (N_6479,N_5678,N_4450);
xnor U6480 (N_6480,N_5040,N_4974);
and U6481 (N_6481,N_5519,N_5458);
nor U6482 (N_6482,N_5141,N_4785);
or U6483 (N_6483,N_4881,N_5703);
or U6484 (N_6484,N_5493,N_5999);
nand U6485 (N_6485,N_5209,N_5179);
nor U6486 (N_6486,N_4573,N_5550);
nor U6487 (N_6487,N_5827,N_4478);
or U6488 (N_6488,N_5948,N_5055);
nand U6489 (N_6489,N_5500,N_5249);
xnor U6490 (N_6490,N_4232,N_4747);
nand U6491 (N_6491,N_4125,N_5738);
and U6492 (N_6492,N_4726,N_4283);
and U6493 (N_6493,N_4574,N_4584);
or U6494 (N_6494,N_5710,N_5962);
or U6495 (N_6495,N_5214,N_5242);
or U6496 (N_6496,N_4103,N_5140);
and U6497 (N_6497,N_5892,N_5385);
or U6498 (N_6498,N_4391,N_4817);
or U6499 (N_6499,N_4833,N_5146);
nor U6500 (N_6500,N_5534,N_4225);
nor U6501 (N_6501,N_5345,N_5492);
nor U6502 (N_6502,N_4464,N_5899);
or U6503 (N_6503,N_4370,N_5810);
or U6504 (N_6504,N_5257,N_4524);
and U6505 (N_6505,N_4243,N_5149);
nor U6506 (N_6506,N_4340,N_5180);
nor U6507 (N_6507,N_4868,N_5095);
nand U6508 (N_6508,N_4883,N_4709);
nand U6509 (N_6509,N_4834,N_4668);
or U6510 (N_6510,N_4346,N_4736);
and U6511 (N_6511,N_4591,N_5276);
nand U6512 (N_6512,N_5473,N_4886);
nor U6513 (N_6513,N_5741,N_5077);
or U6514 (N_6514,N_5380,N_5068);
nand U6515 (N_6515,N_4631,N_5533);
and U6516 (N_6516,N_5832,N_4138);
nor U6517 (N_6517,N_5961,N_4009);
nor U6518 (N_6518,N_5986,N_4680);
or U6519 (N_6519,N_4431,N_4698);
nand U6520 (N_6520,N_4293,N_4420);
or U6521 (N_6521,N_5959,N_4790);
or U6522 (N_6522,N_5036,N_5356);
and U6523 (N_6523,N_5321,N_5595);
and U6524 (N_6524,N_4960,N_4156);
nor U6525 (N_6525,N_5994,N_5178);
and U6526 (N_6526,N_4914,N_4720);
xnor U6527 (N_6527,N_4058,N_5995);
nor U6528 (N_6528,N_4307,N_4440);
nand U6529 (N_6529,N_5731,N_5445);
nor U6530 (N_6530,N_5637,N_5808);
and U6531 (N_6531,N_4713,N_4200);
and U6532 (N_6532,N_5131,N_5070);
nor U6533 (N_6533,N_4113,N_5225);
and U6534 (N_6534,N_4663,N_5636);
nor U6535 (N_6535,N_5181,N_4522);
and U6536 (N_6536,N_4017,N_5489);
xor U6537 (N_6537,N_5091,N_5064);
and U6538 (N_6538,N_4822,N_5813);
or U6539 (N_6539,N_4734,N_5665);
and U6540 (N_6540,N_5764,N_5924);
nand U6541 (N_6541,N_5940,N_4166);
and U6542 (N_6542,N_4381,N_4758);
nand U6543 (N_6543,N_5471,N_4983);
nand U6544 (N_6544,N_5205,N_4173);
nor U6545 (N_6545,N_4097,N_5910);
or U6546 (N_6546,N_5267,N_4672);
or U6547 (N_6547,N_4959,N_5300);
nand U6548 (N_6548,N_5192,N_5772);
or U6549 (N_6549,N_4572,N_5100);
and U6550 (N_6550,N_4379,N_4553);
nor U6551 (N_6551,N_5053,N_5755);
or U6552 (N_6552,N_4987,N_4019);
nand U6553 (N_6553,N_5908,N_5704);
and U6554 (N_6554,N_4576,N_4044);
nand U6555 (N_6555,N_4643,N_4094);
nand U6556 (N_6556,N_5989,N_5243);
nor U6557 (N_6557,N_4792,N_5175);
nand U6558 (N_6558,N_5568,N_5733);
and U6559 (N_6559,N_4835,N_4588);
nor U6560 (N_6560,N_5830,N_4843);
or U6561 (N_6561,N_4640,N_4488);
nor U6562 (N_6562,N_4794,N_4129);
and U6563 (N_6563,N_4900,N_4542);
or U6564 (N_6564,N_4327,N_4392);
or U6565 (N_6565,N_5295,N_5853);
or U6566 (N_6566,N_4197,N_4496);
nand U6567 (N_6567,N_4031,N_5599);
nor U6568 (N_6568,N_5115,N_4922);
nor U6569 (N_6569,N_5990,N_4463);
nand U6570 (N_6570,N_4372,N_4629);
nand U6571 (N_6571,N_4275,N_5634);
or U6572 (N_6572,N_4364,N_4024);
nor U6573 (N_6573,N_4312,N_5641);
nand U6574 (N_6574,N_5355,N_4791);
nor U6575 (N_6575,N_4417,N_5714);
or U6576 (N_6576,N_5838,N_4401);
or U6577 (N_6577,N_5210,N_4375);
nand U6578 (N_6578,N_4540,N_5199);
nor U6579 (N_6579,N_4389,N_5712);
and U6580 (N_6580,N_5279,N_5783);
nand U6581 (N_6581,N_5352,N_5579);
or U6582 (N_6582,N_5979,N_5645);
nor U6583 (N_6583,N_5262,N_5646);
xnor U6584 (N_6584,N_4374,N_4530);
nor U6585 (N_6585,N_5644,N_5184);
nand U6586 (N_6586,N_5110,N_5682);
nor U6587 (N_6587,N_5951,N_4067);
and U6588 (N_6588,N_4442,N_5018);
or U6589 (N_6589,N_4107,N_5194);
or U6590 (N_6590,N_4585,N_5101);
or U6591 (N_6591,N_4645,N_5957);
and U6592 (N_6592,N_4849,N_4241);
nand U6593 (N_6593,N_5876,N_4384);
nand U6594 (N_6594,N_5169,N_4237);
or U6595 (N_6595,N_5394,N_5455);
nand U6596 (N_6596,N_4973,N_5197);
or U6597 (N_6597,N_4767,N_4952);
nor U6598 (N_6598,N_5836,N_4456);
nor U6599 (N_6599,N_5526,N_5517);
nand U6600 (N_6600,N_5860,N_5750);
nand U6601 (N_6601,N_4471,N_5467);
and U6602 (N_6602,N_4062,N_5701);
nand U6603 (N_6603,N_4718,N_5365);
nand U6604 (N_6604,N_5992,N_5277);
nand U6605 (N_6605,N_5332,N_5399);
nor U6606 (N_6606,N_4863,N_4815);
nor U6607 (N_6607,N_5326,N_4360);
nor U6608 (N_6608,N_4961,N_5503);
or U6609 (N_6609,N_4487,N_5336);
xnor U6610 (N_6610,N_4832,N_4852);
or U6611 (N_6611,N_5081,N_5954);
or U6612 (N_6612,N_5919,N_5606);
and U6613 (N_6613,N_4470,N_4875);
nand U6614 (N_6614,N_5762,N_5578);
and U6615 (N_6615,N_5057,N_4145);
nor U6616 (N_6616,N_4474,N_5208);
nand U6617 (N_6617,N_4739,N_4926);
or U6618 (N_6618,N_4806,N_5801);
or U6619 (N_6619,N_4135,N_4676);
or U6620 (N_6620,N_5555,N_5351);
and U6621 (N_6621,N_5017,N_5237);
and U6622 (N_6622,N_4971,N_4828);
or U6623 (N_6623,N_5603,N_4930);
nor U6624 (N_6624,N_4076,N_5358);
nor U6625 (N_6625,N_5894,N_4714);
nand U6626 (N_6626,N_4957,N_4046);
and U6627 (N_6627,N_4543,N_4990);
or U6628 (N_6628,N_4399,N_5596);
or U6629 (N_6629,N_4213,N_4568);
or U6630 (N_6630,N_4492,N_5248);
nand U6631 (N_6631,N_5509,N_5846);
or U6632 (N_6632,N_4309,N_4126);
and U6633 (N_6633,N_4226,N_4651);
nand U6634 (N_6634,N_5315,N_5686);
or U6635 (N_6635,N_5715,N_4079);
or U6636 (N_6636,N_5693,N_5219);
or U6637 (N_6637,N_5699,N_4872);
nor U6638 (N_6638,N_5607,N_4906);
nand U6639 (N_6639,N_4658,N_4049);
and U6640 (N_6640,N_4776,N_5781);
nand U6641 (N_6641,N_4284,N_5135);
and U6642 (N_6642,N_4419,N_5263);
xnor U6643 (N_6643,N_5490,N_5130);
nand U6644 (N_6644,N_5916,N_5771);
or U6645 (N_6645,N_5048,N_5379);
nand U6646 (N_6646,N_4935,N_4596);
nor U6647 (N_6647,N_5843,N_4428);
nor U6648 (N_6648,N_5035,N_4396);
or U6649 (N_6649,N_5459,N_4447);
nor U6650 (N_6650,N_5107,N_4154);
nand U6651 (N_6651,N_4089,N_5497);
or U6652 (N_6652,N_4593,N_5905);
and U6653 (N_6653,N_5768,N_4087);
nor U6654 (N_6654,N_5274,N_4557);
nor U6655 (N_6655,N_4084,N_4967);
nor U6656 (N_6656,N_4889,N_4885);
nand U6657 (N_6657,N_4408,N_5203);
nand U6658 (N_6658,N_4400,N_4932);
nor U6659 (N_6659,N_4786,N_5486);
or U6660 (N_6660,N_5895,N_4607);
or U6661 (N_6661,N_4316,N_5880);
or U6662 (N_6662,N_4073,N_4269);
or U6663 (N_6663,N_5234,N_5449);
or U6664 (N_6664,N_4368,N_4669);
nand U6665 (N_6665,N_5163,N_5118);
nor U6666 (N_6666,N_5502,N_5967);
nor U6667 (N_6667,N_5145,N_5891);
or U6668 (N_6668,N_4302,N_4728);
nor U6669 (N_6669,N_5862,N_5842);
or U6670 (N_6670,N_4616,N_5371);
and U6671 (N_6671,N_4660,N_5825);
or U6672 (N_6672,N_4519,N_5042);
and U6673 (N_6673,N_5086,N_5668);
nor U6674 (N_6674,N_4291,N_4262);
or U6675 (N_6675,N_4940,N_5765);
nor U6676 (N_6676,N_4251,N_4429);
nand U6677 (N_6677,N_5663,N_5465);
or U6678 (N_6678,N_5396,N_4144);
nor U6679 (N_6679,N_4289,N_5439);
and U6680 (N_6680,N_4433,N_4980);
and U6681 (N_6681,N_5478,N_5253);
nand U6682 (N_6682,N_5283,N_4818);
and U6683 (N_6683,N_5221,N_5651);
nand U6684 (N_6684,N_4564,N_4969);
nor U6685 (N_6685,N_4964,N_5170);
or U6686 (N_6686,N_5729,N_5650);
nor U6687 (N_6687,N_5932,N_4382);
nor U6688 (N_6688,N_5238,N_4189);
and U6689 (N_6689,N_5844,N_4483);
nor U6690 (N_6690,N_4285,N_5438);
nor U6691 (N_6691,N_4725,N_5222);
nor U6692 (N_6692,N_4248,N_5513);
nor U6693 (N_6693,N_5633,N_4458);
or U6694 (N_6694,N_4266,N_5403);
or U6695 (N_6695,N_5327,N_4942);
and U6696 (N_6696,N_5436,N_4072);
nand U6697 (N_6697,N_5330,N_4787);
or U6698 (N_6698,N_4749,N_4304);
nor U6699 (N_6699,N_5231,N_5658);
xnor U6700 (N_6700,N_4123,N_4296);
and U6701 (N_6701,N_5956,N_4946);
or U6702 (N_6702,N_5561,N_4308);
and U6703 (N_6703,N_4376,N_4722);
or U6704 (N_6704,N_4869,N_5191);
and U6705 (N_6705,N_4354,N_5882);
and U6706 (N_6706,N_4469,N_4475);
nand U6707 (N_6707,N_4280,N_5007);
nor U6708 (N_6708,N_4717,N_4546);
xnor U6709 (N_6709,N_4535,N_5463);
or U6710 (N_6710,N_5653,N_4516);
or U6711 (N_6711,N_4577,N_5136);
or U6712 (N_6712,N_4279,N_4105);
or U6713 (N_6713,N_5696,N_4702);
nor U6714 (N_6714,N_4796,N_5013);
nand U6715 (N_6715,N_4793,N_4448);
or U6716 (N_6716,N_4115,N_4092);
nor U6717 (N_6717,N_5630,N_4887);
and U6718 (N_6718,N_5290,N_4578);
or U6719 (N_6719,N_5868,N_5087);
and U6720 (N_6720,N_5906,N_5010);
xnor U6721 (N_6721,N_4252,N_4204);
nand U6722 (N_6722,N_4271,N_4763);
nor U6723 (N_6723,N_4913,N_4255);
and U6724 (N_6724,N_5002,N_4453);
and U6725 (N_6725,N_5807,N_4066);
or U6726 (N_6726,N_4923,N_4583);
and U6727 (N_6727,N_5896,N_5338);
and U6728 (N_6728,N_4310,N_4955);
nor U6729 (N_6729,N_4695,N_4650);
nand U6730 (N_6730,N_5104,N_5987);
and U6731 (N_6731,N_4357,N_5122);
nand U6732 (N_6732,N_4294,N_5302);
nor U6733 (N_6733,N_4788,N_4023);
nand U6734 (N_6734,N_4605,N_5656);
nand U6735 (N_6735,N_4866,N_5822);
or U6736 (N_6736,N_5935,N_5664);
or U6737 (N_6737,N_5529,N_5802);
nand U6738 (N_6738,N_5800,N_4521);
and U6739 (N_6739,N_4320,N_5685);
and U6740 (N_6740,N_4128,N_4991);
or U6741 (N_6741,N_5514,N_5469);
and U6742 (N_6742,N_4245,N_4505);
nand U6743 (N_6743,N_4941,N_4132);
or U6744 (N_6744,N_5673,N_5261);
nand U6745 (N_6745,N_4526,N_5381);
and U6746 (N_6746,N_5487,N_4486);
nand U6747 (N_6747,N_4311,N_4841);
nor U6748 (N_6748,N_4070,N_5638);
nor U6749 (N_6749,N_5975,N_4022);
nand U6750 (N_6750,N_4544,N_5297);
nor U6751 (N_6751,N_4882,N_5384);
nor U6752 (N_6752,N_4229,N_5461);
or U6753 (N_6753,N_4598,N_5828);
nor U6754 (N_6754,N_4779,N_4744);
or U6755 (N_6755,N_5431,N_4715);
and U6756 (N_6756,N_5337,N_5334);
or U6757 (N_6757,N_5132,N_5576);
and U6758 (N_6758,N_5670,N_5416);
nor U6759 (N_6759,N_5970,N_4761);
or U6760 (N_6760,N_5280,N_4810);
nand U6761 (N_6761,N_5593,N_4619);
and U6762 (N_6762,N_4222,N_5383);
and U6763 (N_6763,N_5307,N_5826);
or U6764 (N_6764,N_4732,N_5821);
and U6765 (N_6765,N_5158,N_4716);
or U6766 (N_6766,N_5397,N_5138);
or U6767 (N_6767,N_4506,N_4403);
nor U6768 (N_6768,N_4606,N_5216);
xnor U6769 (N_6769,N_4924,N_5066);
or U6770 (N_6770,N_4441,N_4051);
nor U6771 (N_6771,N_5240,N_4406);
nor U6772 (N_6772,N_5364,N_4774);
nor U6773 (N_6773,N_4615,N_5027);
nor U6774 (N_6774,N_4595,N_4842);
or U6775 (N_6775,N_5766,N_4394);
or U6776 (N_6776,N_5770,N_4140);
nand U6777 (N_6777,N_4703,N_4580);
nor U6778 (N_6778,N_5740,N_4455);
and U6779 (N_6779,N_5480,N_4534);
or U6780 (N_6780,N_5865,N_4147);
nand U6781 (N_6781,N_4829,N_4993);
nor U6782 (N_6782,N_4160,N_5108);
and U6783 (N_6783,N_5609,N_4514);
nand U6784 (N_6784,N_5922,N_5695);
and U6785 (N_6785,N_4342,N_5393);
and U6786 (N_6786,N_5855,N_4355);
nor U6787 (N_6787,N_4152,N_5817);
nand U6788 (N_6788,N_5725,N_5869);
nand U6789 (N_6789,N_5717,N_5096);
nor U6790 (N_6790,N_4134,N_5076);
or U6791 (N_6791,N_4258,N_5453);
nor U6792 (N_6792,N_5421,N_5349);
or U6793 (N_6793,N_4055,N_4566);
or U6794 (N_6794,N_5914,N_5966);
and U6795 (N_6795,N_4032,N_4903);
or U6796 (N_6796,N_4624,N_4167);
and U6797 (N_6797,N_5304,N_4148);
nor U6798 (N_6798,N_4707,N_4466);
nand U6799 (N_6799,N_4332,N_5318);
nor U6800 (N_6800,N_4626,N_4826);
and U6801 (N_6801,N_4992,N_4214);
or U6802 (N_6802,N_4227,N_4424);
nor U6803 (N_6803,N_4989,N_4804);
nor U6804 (N_6804,N_4053,N_5370);
nand U6805 (N_6805,N_4743,N_5306);
nor U6806 (N_6806,N_5168,N_4963);
xnor U6807 (N_6807,N_5124,N_5498);
or U6808 (N_6808,N_4246,N_5726);
and U6809 (N_6809,N_4878,N_5019);
or U6810 (N_6810,N_4423,N_5660);
nand U6811 (N_6811,N_5362,N_4943);
or U6812 (N_6812,N_5711,N_5114);
nor U6813 (N_6813,N_4350,N_5903);
and U6814 (N_6814,N_4814,N_4409);
nor U6815 (N_6815,N_5133,N_4300);
or U6816 (N_6816,N_5632,N_5026);
nand U6817 (N_6817,N_5835,N_4634);
nor U6818 (N_6818,N_4008,N_5270);
nand U6819 (N_6819,N_4435,N_5443);
nand U6820 (N_6820,N_5850,N_5969);
and U6821 (N_6821,N_4801,N_5173);
nor U6822 (N_6822,N_4919,N_5558);
or U6823 (N_6823,N_4927,N_4682);
nor U6824 (N_6824,N_4503,N_5251);
nor U6825 (N_6825,N_5218,N_5784);
or U6826 (N_6826,N_5071,N_5925);
nor U6827 (N_6827,N_4997,N_5165);
or U6828 (N_6828,N_5759,N_5195);
and U6829 (N_6829,N_4637,N_5211);
and U6830 (N_6830,N_4857,N_5570);
and U6831 (N_6831,N_4223,N_5106);
or U6832 (N_6832,N_5622,N_4002);
or U6833 (N_6833,N_4871,N_4916);
or U6834 (N_6834,N_5062,N_4015);
nand U6835 (N_6835,N_4260,N_5917);
nand U6836 (N_6836,N_5617,N_5444);
or U6837 (N_6837,N_5911,N_5666);
nand U6838 (N_6838,N_4141,N_4170);
or U6839 (N_6839,N_5090,N_4457);
nor U6840 (N_6840,N_5282,N_5363);
nand U6841 (N_6841,N_5388,N_4270);
xor U6842 (N_6842,N_5442,N_4034);
nand U6843 (N_6843,N_4947,N_5833);
or U6844 (N_6844,N_4467,N_4988);
nor U6845 (N_6845,N_4665,N_5560);
or U6846 (N_6846,N_5720,N_4341);
or U6847 (N_6847,N_5139,N_5790);
and U6848 (N_6848,N_5020,N_5623);
nor U6849 (N_6849,N_4348,N_4292);
or U6850 (N_6850,N_4620,N_4898);
nand U6851 (N_6851,N_5343,N_4169);
or U6852 (N_6852,N_4069,N_4052);
nor U6853 (N_6853,N_5933,N_4122);
and U6854 (N_6854,N_5515,N_5085);
or U6855 (N_6855,N_4460,N_5250);
or U6856 (N_6856,N_4325,N_4892);
and U6857 (N_6857,N_4306,N_5161);
nand U6858 (N_6858,N_5946,N_4562);
and U6859 (N_6859,N_5522,N_5103);
and U6860 (N_6860,N_5410,N_5028);
or U6861 (N_6861,N_4561,N_4661);
nor U6862 (N_6862,N_5756,N_5201);
or U6863 (N_6863,N_5611,N_5592);
and U6864 (N_6864,N_4601,N_5829);
xor U6865 (N_6865,N_4205,N_5524);
nand U6866 (N_6866,N_4686,N_4016);
nor U6867 (N_6867,N_4194,N_4590);
and U6868 (N_6868,N_5538,N_5470);
nand U6869 (N_6869,N_4267,N_4098);
nor U6870 (N_6870,N_4667,N_5435);
and U6871 (N_6871,N_5688,N_5984);
xnor U6872 (N_6872,N_5228,N_4614);
nand U6873 (N_6873,N_5310,N_5814);
nor U6874 (N_6874,N_5217,N_4839);
nor U6875 (N_6875,N_5398,N_4111);
nor U6876 (N_6876,N_5116,N_4057);
and U6877 (N_6877,N_5767,N_5294);
or U6878 (N_6878,N_5620,N_4281);
and U6879 (N_6879,N_5298,N_5605);
nor U6880 (N_6880,N_5128,N_5354);
nand U6881 (N_6881,N_5557,N_4272);
nor U6882 (N_6882,N_5011,N_5378);
nand U6883 (N_6883,N_4657,N_5353);
or U6884 (N_6884,N_4711,N_4976);
nand U6885 (N_6885,N_4083,N_5542);
nor U6886 (N_6886,N_4649,N_4114);
nand U6887 (N_6887,N_5831,N_5448);
nand U6888 (N_6888,N_5901,N_4234);
nor U6889 (N_6889,N_4277,N_4905);
and U6890 (N_6890,N_4867,N_4043);
or U6891 (N_6891,N_5395,N_4193);
or U6892 (N_6892,N_4472,N_5346);
or U6893 (N_6893,N_5649,N_4958);
xnor U6894 (N_6894,N_4188,N_5546);
or U6895 (N_6895,N_5043,N_5483);
nor U6896 (N_6896,N_4984,N_4385);
or U6897 (N_6897,N_5657,N_4537);
nand U6898 (N_6898,N_5773,N_4603);
nand U6899 (N_6899,N_4858,N_5993);
and U6900 (N_6900,N_5820,N_4556);
nor U6901 (N_6901,N_4217,N_4656);
or U6902 (N_6902,N_4050,N_5553);
nor U6903 (N_6903,N_4931,N_5239);
or U6904 (N_6904,N_5386,N_4515);
or U6905 (N_6905,N_4088,N_5266);
nor U6906 (N_6906,N_4405,N_5041);
nand U6907 (N_6907,N_5888,N_5708);
nor U6908 (N_6908,N_5015,N_5737);
or U6909 (N_6909,N_4449,N_4938);
nor U6910 (N_6910,N_4479,N_5148);
nand U6911 (N_6911,N_4186,N_5902);
or U6912 (N_6912,N_5348,N_5256);
nor U6913 (N_6913,N_5451,N_5958);
and U6914 (N_6914,N_5060,N_4443);
nor U6915 (N_6915,N_5382,N_4454);
and U6916 (N_6916,N_4162,N_5728);
nand U6917 (N_6917,N_5373,N_4666);
and U6918 (N_6918,N_4721,N_5359);
nand U6919 (N_6919,N_4161,N_5585);
nor U6920 (N_6920,N_5317,N_4647);
or U6921 (N_6921,N_5639,N_5530);
or U6922 (N_6922,N_4244,N_5811);
nand U6923 (N_6923,N_5481,N_4481);
and U6924 (N_6924,N_5687,N_4696);
nor U6925 (N_6925,N_5376,N_4708);
nor U6926 (N_6926,N_5789,N_5072);
or U6927 (N_6927,N_4100,N_4917);
or U6928 (N_6928,N_4171,N_4108);
and U6929 (N_6929,N_5123,N_4571);
xor U6930 (N_6930,N_5369,N_5477);
or U6931 (N_6931,N_4322,N_4888);
and U6932 (N_6932,N_5672,N_5859);
or U6933 (N_6933,N_5881,N_5722);
nand U6934 (N_6934,N_4174,N_4689);
or U6935 (N_6935,N_5083,N_5084);
nor U6936 (N_6936,N_4045,N_5879);
or U6937 (N_6937,N_5422,N_4165);
nor U6938 (N_6938,N_5361,N_4367);
nand U6939 (N_6939,N_4921,N_4830);
nand U6940 (N_6940,N_5185,N_5554);
nand U6941 (N_6941,N_4263,N_4950);
and U6942 (N_6942,N_5584,N_5447);
nor U6943 (N_6943,N_5329,N_5921);
or U6944 (N_6944,N_4907,N_5176);
or U6945 (N_6945,N_4639,N_4038);
and U6946 (N_6946,N_5615,N_5152);
or U6947 (N_6947,N_4181,N_4414);
or U6948 (N_6948,N_4178,N_4710);
nor U6949 (N_6949,N_4484,N_4589);
nor U6950 (N_6950,N_4678,N_5545);
or U6951 (N_6951,N_4183,N_5319);
nor U6952 (N_6952,N_5871,N_4040);
or U6953 (N_6953,N_4773,N_5730);
nor U6954 (N_6954,N_4623,N_4700);
nor U6955 (N_6955,N_5537,N_4567);
nand U6956 (N_6956,N_4187,N_5182);
nand U6957 (N_6957,N_5667,N_5635);
nor U6958 (N_6958,N_4902,N_5177);
nor U6959 (N_6959,N_4380,N_4925);
or U6960 (N_6960,N_5749,N_4497);
nor U6961 (N_6961,N_5499,N_4422);
xnor U6962 (N_6962,N_4233,N_4096);
and U6963 (N_6963,N_5484,N_5907);
or U6964 (N_6964,N_5412,N_4090);
and U6965 (N_6965,N_4502,N_4278);
and U6966 (N_6966,N_5207,N_5824);
and U6967 (N_6967,N_4509,N_4864);
or U6968 (N_6968,N_4904,N_5212);
and U6969 (N_6969,N_4158,N_4860);
nor U6970 (N_6970,N_4020,N_4276);
nor U6971 (N_6971,N_4337,N_4945);
nand U6972 (N_6972,N_5757,N_5837);
nor U6973 (N_6973,N_4880,N_5187);
nand U6974 (N_6974,N_4753,N_5776);
nand U6975 (N_6975,N_4685,N_5157);
and U6976 (N_6976,N_5046,N_4529);
nand U6977 (N_6977,N_4599,N_4510);
or U6978 (N_6978,N_4264,N_5677);
or U6979 (N_6979,N_4344,N_5291);
nand U6980 (N_6980,N_4654,N_4465);
or U6981 (N_6981,N_5419,N_5372);
nor U6982 (N_6982,N_4675,N_4338);
nand U6983 (N_6983,N_5153,N_4212);
nor U6984 (N_6984,N_4075,N_4091);
and U6985 (N_6985,N_4962,N_4662);
or U6986 (N_6986,N_5004,N_4691);
or U6987 (N_6987,N_4972,N_5230);
or U6988 (N_6988,N_5129,N_4288);
and U6989 (N_6989,N_4209,N_5117);
and U6990 (N_6990,N_5600,N_4402);
nand U6991 (N_6991,N_4895,N_5024);
or U6992 (N_6992,N_4746,N_4679);
or U6993 (N_6993,N_4012,N_4377);
nor U6994 (N_6994,N_5897,N_5404);
nor U6995 (N_6995,N_4854,N_5082);
and U6996 (N_6996,N_4772,N_5501);
nor U6997 (N_6997,N_4257,N_4136);
nor U6998 (N_6998,N_4439,N_5815);
and U6999 (N_6999,N_4434,N_5016);
and U7000 (N_7000,N_5557,N_4615);
nor U7001 (N_7001,N_4896,N_4550);
nor U7002 (N_7002,N_5802,N_4046);
or U7003 (N_7003,N_5668,N_5867);
and U7004 (N_7004,N_5827,N_5626);
and U7005 (N_7005,N_4022,N_4584);
or U7006 (N_7006,N_5539,N_4876);
and U7007 (N_7007,N_4539,N_5380);
nand U7008 (N_7008,N_5348,N_4023);
and U7009 (N_7009,N_5533,N_4717);
or U7010 (N_7010,N_4089,N_5947);
nor U7011 (N_7011,N_4021,N_4742);
nor U7012 (N_7012,N_4242,N_5258);
nor U7013 (N_7013,N_4085,N_4079);
and U7014 (N_7014,N_4118,N_5298);
nand U7015 (N_7015,N_4086,N_5010);
or U7016 (N_7016,N_5516,N_5586);
and U7017 (N_7017,N_4299,N_4997);
or U7018 (N_7018,N_4377,N_4696);
nand U7019 (N_7019,N_4115,N_4943);
and U7020 (N_7020,N_5996,N_4000);
and U7021 (N_7021,N_5010,N_4376);
or U7022 (N_7022,N_4891,N_4578);
and U7023 (N_7023,N_5071,N_4571);
nand U7024 (N_7024,N_5330,N_5693);
nand U7025 (N_7025,N_4250,N_5816);
and U7026 (N_7026,N_5076,N_5726);
nor U7027 (N_7027,N_5709,N_5011);
and U7028 (N_7028,N_4079,N_4819);
nand U7029 (N_7029,N_4011,N_5987);
or U7030 (N_7030,N_5122,N_5058);
or U7031 (N_7031,N_4306,N_5227);
and U7032 (N_7032,N_4269,N_5354);
or U7033 (N_7033,N_4522,N_4695);
and U7034 (N_7034,N_4763,N_5397);
and U7035 (N_7035,N_5411,N_4697);
or U7036 (N_7036,N_5362,N_4411);
or U7037 (N_7037,N_4521,N_5203);
or U7038 (N_7038,N_4507,N_5778);
nor U7039 (N_7039,N_4746,N_5261);
nor U7040 (N_7040,N_5094,N_5380);
nor U7041 (N_7041,N_5190,N_4650);
or U7042 (N_7042,N_4576,N_4530);
or U7043 (N_7043,N_5384,N_4438);
or U7044 (N_7044,N_4706,N_5871);
and U7045 (N_7045,N_4703,N_4047);
nor U7046 (N_7046,N_4045,N_4639);
and U7047 (N_7047,N_5493,N_4784);
or U7048 (N_7048,N_5185,N_5634);
and U7049 (N_7049,N_4488,N_5502);
and U7050 (N_7050,N_5151,N_5437);
and U7051 (N_7051,N_4600,N_4449);
or U7052 (N_7052,N_5313,N_5897);
or U7053 (N_7053,N_4343,N_4644);
and U7054 (N_7054,N_5531,N_5446);
nor U7055 (N_7055,N_4709,N_5399);
and U7056 (N_7056,N_5713,N_4095);
nand U7057 (N_7057,N_4227,N_4201);
or U7058 (N_7058,N_4345,N_5585);
or U7059 (N_7059,N_5142,N_4435);
or U7060 (N_7060,N_5075,N_4125);
nor U7061 (N_7061,N_4308,N_4739);
nand U7062 (N_7062,N_5592,N_5072);
or U7063 (N_7063,N_4032,N_5202);
and U7064 (N_7064,N_5211,N_5315);
or U7065 (N_7065,N_4192,N_5701);
and U7066 (N_7066,N_5540,N_5938);
and U7067 (N_7067,N_5709,N_5082);
and U7068 (N_7068,N_5418,N_5054);
or U7069 (N_7069,N_5434,N_4502);
and U7070 (N_7070,N_4800,N_4839);
nor U7071 (N_7071,N_5137,N_4241);
nor U7072 (N_7072,N_5165,N_4745);
and U7073 (N_7073,N_5167,N_5982);
and U7074 (N_7074,N_4748,N_4011);
nor U7075 (N_7075,N_5206,N_5466);
or U7076 (N_7076,N_4592,N_5986);
nand U7077 (N_7077,N_4449,N_5632);
or U7078 (N_7078,N_4507,N_4038);
or U7079 (N_7079,N_4375,N_5906);
nor U7080 (N_7080,N_4169,N_4124);
and U7081 (N_7081,N_4017,N_5410);
and U7082 (N_7082,N_4991,N_5304);
nor U7083 (N_7083,N_5651,N_4697);
nor U7084 (N_7084,N_4473,N_5821);
or U7085 (N_7085,N_5691,N_5939);
and U7086 (N_7086,N_5944,N_4366);
nor U7087 (N_7087,N_5257,N_5734);
nor U7088 (N_7088,N_4932,N_5875);
and U7089 (N_7089,N_5472,N_5467);
xor U7090 (N_7090,N_4802,N_5592);
nor U7091 (N_7091,N_5588,N_5146);
nor U7092 (N_7092,N_5900,N_5235);
nand U7093 (N_7093,N_5515,N_4708);
or U7094 (N_7094,N_4872,N_5232);
and U7095 (N_7095,N_5425,N_4510);
nor U7096 (N_7096,N_5134,N_4786);
nor U7097 (N_7097,N_4869,N_5192);
and U7098 (N_7098,N_4850,N_5770);
or U7099 (N_7099,N_5752,N_5646);
or U7100 (N_7100,N_5642,N_4468);
nand U7101 (N_7101,N_4727,N_4502);
and U7102 (N_7102,N_4715,N_4584);
and U7103 (N_7103,N_5866,N_5733);
nand U7104 (N_7104,N_4441,N_5469);
nor U7105 (N_7105,N_5664,N_4971);
nand U7106 (N_7106,N_4174,N_4794);
and U7107 (N_7107,N_5745,N_4339);
and U7108 (N_7108,N_5366,N_5471);
nor U7109 (N_7109,N_4764,N_4586);
nor U7110 (N_7110,N_5388,N_4117);
nand U7111 (N_7111,N_5837,N_4597);
and U7112 (N_7112,N_5204,N_4295);
and U7113 (N_7113,N_5076,N_4496);
or U7114 (N_7114,N_4868,N_4629);
nor U7115 (N_7115,N_5552,N_4410);
nor U7116 (N_7116,N_5657,N_5779);
nand U7117 (N_7117,N_4692,N_5766);
and U7118 (N_7118,N_4455,N_5491);
and U7119 (N_7119,N_4377,N_5705);
and U7120 (N_7120,N_4196,N_4534);
or U7121 (N_7121,N_4862,N_5802);
nor U7122 (N_7122,N_5849,N_4933);
nor U7123 (N_7123,N_5344,N_4901);
nand U7124 (N_7124,N_4781,N_5256);
and U7125 (N_7125,N_5704,N_5998);
nand U7126 (N_7126,N_5246,N_4767);
and U7127 (N_7127,N_5097,N_4545);
and U7128 (N_7128,N_5155,N_4831);
nand U7129 (N_7129,N_4036,N_5753);
nor U7130 (N_7130,N_4027,N_4030);
nand U7131 (N_7131,N_4257,N_4768);
nor U7132 (N_7132,N_4438,N_4936);
and U7133 (N_7133,N_5712,N_4204);
nand U7134 (N_7134,N_5386,N_5030);
nor U7135 (N_7135,N_4120,N_5268);
and U7136 (N_7136,N_5226,N_4406);
nand U7137 (N_7137,N_4722,N_4958);
and U7138 (N_7138,N_4057,N_5284);
and U7139 (N_7139,N_5718,N_4876);
nand U7140 (N_7140,N_4015,N_5976);
and U7141 (N_7141,N_4244,N_5060);
nand U7142 (N_7142,N_4721,N_4588);
or U7143 (N_7143,N_5413,N_5124);
nand U7144 (N_7144,N_5018,N_5406);
or U7145 (N_7145,N_4568,N_5452);
nor U7146 (N_7146,N_5365,N_5010);
nand U7147 (N_7147,N_4560,N_5509);
and U7148 (N_7148,N_5632,N_5187);
or U7149 (N_7149,N_4460,N_5605);
and U7150 (N_7150,N_4796,N_4488);
nand U7151 (N_7151,N_5165,N_4583);
or U7152 (N_7152,N_4924,N_5231);
nand U7153 (N_7153,N_4643,N_4130);
nor U7154 (N_7154,N_4940,N_4760);
and U7155 (N_7155,N_4575,N_5218);
or U7156 (N_7156,N_5032,N_5718);
nor U7157 (N_7157,N_5559,N_5446);
and U7158 (N_7158,N_5519,N_4133);
nand U7159 (N_7159,N_4306,N_4948);
and U7160 (N_7160,N_5302,N_5088);
nor U7161 (N_7161,N_5256,N_5776);
nand U7162 (N_7162,N_5365,N_5853);
and U7163 (N_7163,N_5673,N_4747);
and U7164 (N_7164,N_4879,N_5755);
or U7165 (N_7165,N_5723,N_4258);
or U7166 (N_7166,N_4561,N_4743);
and U7167 (N_7167,N_5475,N_4738);
or U7168 (N_7168,N_4415,N_4323);
or U7169 (N_7169,N_5661,N_5680);
or U7170 (N_7170,N_4589,N_5878);
nand U7171 (N_7171,N_4739,N_5160);
nor U7172 (N_7172,N_5582,N_5478);
nand U7173 (N_7173,N_4409,N_4800);
nor U7174 (N_7174,N_4062,N_4102);
or U7175 (N_7175,N_5879,N_4682);
nor U7176 (N_7176,N_5327,N_5836);
or U7177 (N_7177,N_5801,N_4011);
nand U7178 (N_7178,N_5996,N_5698);
nand U7179 (N_7179,N_5958,N_5048);
or U7180 (N_7180,N_4207,N_4565);
or U7181 (N_7181,N_4425,N_4946);
nand U7182 (N_7182,N_4561,N_5998);
or U7183 (N_7183,N_5892,N_4006);
nor U7184 (N_7184,N_5109,N_4938);
or U7185 (N_7185,N_4095,N_5926);
and U7186 (N_7186,N_5319,N_4341);
xor U7187 (N_7187,N_5348,N_5557);
and U7188 (N_7188,N_4220,N_4877);
nor U7189 (N_7189,N_5549,N_5095);
nand U7190 (N_7190,N_5680,N_4171);
or U7191 (N_7191,N_5484,N_5805);
and U7192 (N_7192,N_4170,N_5347);
nor U7193 (N_7193,N_4208,N_4795);
nor U7194 (N_7194,N_4288,N_5408);
and U7195 (N_7195,N_5664,N_4853);
or U7196 (N_7196,N_5308,N_4582);
nand U7197 (N_7197,N_5372,N_4926);
or U7198 (N_7198,N_4938,N_4051);
or U7199 (N_7199,N_4825,N_5917);
nand U7200 (N_7200,N_4057,N_5990);
and U7201 (N_7201,N_4847,N_4488);
or U7202 (N_7202,N_5040,N_4013);
nand U7203 (N_7203,N_4307,N_5586);
and U7204 (N_7204,N_4609,N_5746);
nand U7205 (N_7205,N_5991,N_5074);
and U7206 (N_7206,N_4463,N_4455);
or U7207 (N_7207,N_4122,N_4243);
nand U7208 (N_7208,N_5266,N_4833);
and U7209 (N_7209,N_5532,N_5492);
nor U7210 (N_7210,N_5611,N_5416);
nand U7211 (N_7211,N_5216,N_5880);
or U7212 (N_7212,N_4371,N_4392);
nor U7213 (N_7213,N_5655,N_4854);
and U7214 (N_7214,N_4437,N_5921);
or U7215 (N_7215,N_5333,N_5922);
nor U7216 (N_7216,N_4913,N_5138);
nand U7217 (N_7217,N_5866,N_4094);
xor U7218 (N_7218,N_5113,N_5723);
and U7219 (N_7219,N_4878,N_5547);
and U7220 (N_7220,N_5304,N_4444);
and U7221 (N_7221,N_4570,N_5835);
and U7222 (N_7222,N_4040,N_5703);
nor U7223 (N_7223,N_4328,N_5882);
nor U7224 (N_7224,N_5193,N_4994);
and U7225 (N_7225,N_4614,N_4151);
and U7226 (N_7226,N_5749,N_4532);
and U7227 (N_7227,N_4011,N_5993);
and U7228 (N_7228,N_5785,N_4726);
nor U7229 (N_7229,N_4435,N_5927);
and U7230 (N_7230,N_4890,N_5604);
nand U7231 (N_7231,N_5951,N_5701);
nand U7232 (N_7232,N_4510,N_5439);
nor U7233 (N_7233,N_5240,N_5310);
or U7234 (N_7234,N_5340,N_5378);
and U7235 (N_7235,N_5371,N_5423);
nor U7236 (N_7236,N_5796,N_5979);
xor U7237 (N_7237,N_4374,N_4358);
nor U7238 (N_7238,N_4675,N_4633);
nand U7239 (N_7239,N_4513,N_4496);
nor U7240 (N_7240,N_5335,N_5320);
nand U7241 (N_7241,N_5871,N_5476);
or U7242 (N_7242,N_5099,N_5575);
nand U7243 (N_7243,N_4379,N_4213);
and U7244 (N_7244,N_5319,N_5804);
nand U7245 (N_7245,N_4489,N_4496);
nand U7246 (N_7246,N_5735,N_5829);
or U7247 (N_7247,N_4762,N_5418);
nand U7248 (N_7248,N_5171,N_5262);
or U7249 (N_7249,N_4270,N_4991);
or U7250 (N_7250,N_5616,N_4187);
and U7251 (N_7251,N_4959,N_4456);
nor U7252 (N_7252,N_5104,N_4292);
or U7253 (N_7253,N_4994,N_4297);
or U7254 (N_7254,N_5569,N_5896);
nand U7255 (N_7255,N_5228,N_4748);
and U7256 (N_7256,N_4839,N_5507);
and U7257 (N_7257,N_5112,N_5815);
and U7258 (N_7258,N_4066,N_5206);
nand U7259 (N_7259,N_4250,N_4482);
and U7260 (N_7260,N_4243,N_4990);
or U7261 (N_7261,N_5443,N_4376);
and U7262 (N_7262,N_5433,N_5923);
nor U7263 (N_7263,N_4820,N_5816);
nor U7264 (N_7264,N_4181,N_5722);
nor U7265 (N_7265,N_5218,N_4665);
and U7266 (N_7266,N_5181,N_5726);
xnor U7267 (N_7267,N_4137,N_5502);
nor U7268 (N_7268,N_4650,N_4341);
xnor U7269 (N_7269,N_5499,N_4825);
and U7270 (N_7270,N_5456,N_4495);
nor U7271 (N_7271,N_5752,N_4500);
nor U7272 (N_7272,N_5759,N_4021);
nand U7273 (N_7273,N_5947,N_4958);
nand U7274 (N_7274,N_4220,N_4825);
nand U7275 (N_7275,N_5447,N_4658);
and U7276 (N_7276,N_4194,N_5808);
or U7277 (N_7277,N_5747,N_5877);
or U7278 (N_7278,N_5343,N_5480);
and U7279 (N_7279,N_5762,N_5120);
or U7280 (N_7280,N_5713,N_5219);
nand U7281 (N_7281,N_5753,N_4045);
nor U7282 (N_7282,N_5092,N_5201);
or U7283 (N_7283,N_5047,N_4685);
nand U7284 (N_7284,N_5743,N_4069);
nand U7285 (N_7285,N_4116,N_5745);
and U7286 (N_7286,N_5774,N_5240);
and U7287 (N_7287,N_5977,N_5813);
nand U7288 (N_7288,N_4860,N_4363);
or U7289 (N_7289,N_5600,N_5404);
and U7290 (N_7290,N_5573,N_4730);
or U7291 (N_7291,N_5049,N_4427);
nand U7292 (N_7292,N_5757,N_5564);
nor U7293 (N_7293,N_5991,N_4851);
nand U7294 (N_7294,N_4094,N_5060);
and U7295 (N_7295,N_5829,N_5772);
or U7296 (N_7296,N_4139,N_4256);
nor U7297 (N_7297,N_5281,N_5241);
xnor U7298 (N_7298,N_4754,N_4144);
and U7299 (N_7299,N_4489,N_5194);
or U7300 (N_7300,N_5234,N_4090);
nand U7301 (N_7301,N_5085,N_5065);
and U7302 (N_7302,N_4204,N_4474);
nand U7303 (N_7303,N_4107,N_5095);
nand U7304 (N_7304,N_4701,N_5145);
nor U7305 (N_7305,N_4097,N_4725);
and U7306 (N_7306,N_5511,N_5671);
and U7307 (N_7307,N_4969,N_5460);
nor U7308 (N_7308,N_4691,N_5206);
or U7309 (N_7309,N_4016,N_5274);
nand U7310 (N_7310,N_4426,N_4441);
and U7311 (N_7311,N_5796,N_4536);
and U7312 (N_7312,N_5794,N_4693);
or U7313 (N_7313,N_5261,N_5427);
nor U7314 (N_7314,N_5323,N_5106);
nor U7315 (N_7315,N_4967,N_4590);
nand U7316 (N_7316,N_4570,N_5480);
nand U7317 (N_7317,N_4893,N_4512);
or U7318 (N_7318,N_4809,N_5543);
and U7319 (N_7319,N_5362,N_5310);
or U7320 (N_7320,N_4351,N_5367);
and U7321 (N_7321,N_5437,N_4171);
or U7322 (N_7322,N_5169,N_5566);
and U7323 (N_7323,N_5007,N_4103);
nor U7324 (N_7324,N_5839,N_4369);
or U7325 (N_7325,N_5920,N_4730);
and U7326 (N_7326,N_5958,N_4882);
nand U7327 (N_7327,N_4314,N_4421);
or U7328 (N_7328,N_5068,N_4183);
nor U7329 (N_7329,N_4815,N_5414);
nor U7330 (N_7330,N_5996,N_5492);
nand U7331 (N_7331,N_5183,N_5875);
and U7332 (N_7332,N_4768,N_4870);
nand U7333 (N_7333,N_5313,N_4281);
and U7334 (N_7334,N_5038,N_5172);
or U7335 (N_7335,N_4411,N_4550);
and U7336 (N_7336,N_4432,N_5407);
nor U7337 (N_7337,N_5478,N_4359);
or U7338 (N_7338,N_4862,N_5856);
nor U7339 (N_7339,N_4446,N_4206);
or U7340 (N_7340,N_5382,N_4824);
nand U7341 (N_7341,N_4994,N_5492);
and U7342 (N_7342,N_5978,N_5170);
and U7343 (N_7343,N_5223,N_5136);
nor U7344 (N_7344,N_4220,N_4987);
or U7345 (N_7345,N_4524,N_5453);
nor U7346 (N_7346,N_4604,N_4688);
and U7347 (N_7347,N_5207,N_5924);
nand U7348 (N_7348,N_4776,N_5975);
and U7349 (N_7349,N_4765,N_4847);
and U7350 (N_7350,N_5023,N_5888);
or U7351 (N_7351,N_5885,N_4632);
and U7352 (N_7352,N_4846,N_5491);
nand U7353 (N_7353,N_4145,N_4557);
nor U7354 (N_7354,N_5781,N_4902);
and U7355 (N_7355,N_4111,N_4439);
or U7356 (N_7356,N_5075,N_4110);
and U7357 (N_7357,N_5471,N_5019);
nand U7358 (N_7358,N_4685,N_4241);
nor U7359 (N_7359,N_5520,N_4345);
or U7360 (N_7360,N_4557,N_5071);
or U7361 (N_7361,N_5639,N_4038);
or U7362 (N_7362,N_5363,N_4550);
nor U7363 (N_7363,N_5163,N_4924);
or U7364 (N_7364,N_5528,N_4319);
and U7365 (N_7365,N_5357,N_4424);
nand U7366 (N_7366,N_4057,N_5902);
or U7367 (N_7367,N_4765,N_5920);
or U7368 (N_7368,N_5234,N_4817);
or U7369 (N_7369,N_5207,N_4456);
and U7370 (N_7370,N_4571,N_5832);
nor U7371 (N_7371,N_5830,N_4642);
or U7372 (N_7372,N_5531,N_5889);
nor U7373 (N_7373,N_5409,N_5333);
or U7374 (N_7374,N_5936,N_5154);
nand U7375 (N_7375,N_5860,N_4912);
or U7376 (N_7376,N_5820,N_5376);
nor U7377 (N_7377,N_5985,N_5257);
nor U7378 (N_7378,N_5818,N_4523);
nand U7379 (N_7379,N_4302,N_5135);
and U7380 (N_7380,N_4815,N_5010);
nor U7381 (N_7381,N_5943,N_5314);
and U7382 (N_7382,N_5647,N_5397);
or U7383 (N_7383,N_5659,N_4861);
nand U7384 (N_7384,N_5592,N_4348);
and U7385 (N_7385,N_5976,N_5557);
nand U7386 (N_7386,N_5908,N_5011);
nand U7387 (N_7387,N_5662,N_4374);
nor U7388 (N_7388,N_5119,N_4417);
or U7389 (N_7389,N_5768,N_5975);
nand U7390 (N_7390,N_4319,N_5606);
and U7391 (N_7391,N_5359,N_4406);
nor U7392 (N_7392,N_4157,N_4923);
and U7393 (N_7393,N_5920,N_4791);
nor U7394 (N_7394,N_4071,N_4006);
nor U7395 (N_7395,N_5573,N_4298);
nand U7396 (N_7396,N_5329,N_5805);
and U7397 (N_7397,N_4269,N_5959);
nand U7398 (N_7398,N_4651,N_4847);
nor U7399 (N_7399,N_5026,N_4189);
nor U7400 (N_7400,N_5462,N_5934);
nand U7401 (N_7401,N_5231,N_4857);
nor U7402 (N_7402,N_5931,N_4039);
or U7403 (N_7403,N_4389,N_4845);
and U7404 (N_7404,N_5734,N_5206);
or U7405 (N_7405,N_4741,N_5725);
or U7406 (N_7406,N_5691,N_4193);
and U7407 (N_7407,N_5368,N_5397);
nand U7408 (N_7408,N_4911,N_5033);
or U7409 (N_7409,N_5380,N_5990);
and U7410 (N_7410,N_5594,N_4020);
and U7411 (N_7411,N_5208,N_5116);
and U7412 (N_7412,N_4051,N_4439);
and U7413 (N_7413,N_4331,N_4814);
nand U7414 (N_7414,N_5920,N_5112);
nor U7415 (N_7415,N_4297,N_4602);
nand U7416 (N_7416,N_5559,N_4055);
and U7417 (N_7417,N_4034,N_5479);
or U7418 (N_7418,N_5600,N_4557);
or U7419 (N_7419,N_4744,N_5233);
and U7420 (N_7420,N_5896,N_5501);
or U7421 (N_7421,N_5562,N_4077);
nand U7422 (N_7422,N_4185,N_4392);
or U7423 (N_7423,N_5901,N_5259);
or U7424 (N_7424,N_5760,N_4176);
or U7425 (N_7425,N_5631,N_5218);
nor U7426 (N_7426,N_5339,N_4946);
and U7427 (N_7427,N_5064,N_5422);
xnor U7428 (N_7428,N_5395,N_5924);
nor U7429 (N_7429,N_5085,N_5916);
and U7430 (N_7430,N_5174,N_5023);
nor U7431 (N_7431,N_4389,N_5433);
and U7432 (N_7432,N_4717,N_4109);
nand U7433 (N_7433,N_4164,N_5911);
nor U7434 (N_7434,N_4921,N_4089);
nand U7435 (N_7435,N_4756,N_4136);
and U7436 (N_7436,N_4610,N_5746);
nor U7437 (N_7437,N_5173,N_4384);
nor U7438 (N_7438,N_4969,N_4416);
or U7439 (N_7439,N_5961,N_4089);
or U7440 (N_7440,N_5512,N_4370);
or U7441 (N_7441,N_4392,N_5640);
or U7442 (N_7442,N_5366,N_5491);
nor U7443 (N_7443,N_4835,N_4148);
nand U7444 (N_7444,N_4775,N_5110);
nor U7445 (N_7445,N_4747,N_5830);
nand U7446 (N_7446,N_4663,N_4698);
or U7447 (N_7447,N_4150,N_5756);
and U7448 (N_7448,N_4383,N_4621);
and U7449 (N_7449,N_5583,N_4523);
or U7450 (N_7450,N_5682,N_5809);
nand U7451 (N_7451,N_5316,N_5412);
nor U7452 (N_7452,N_5954,N_5019);
or U7453 (N_7453,N_4456,N_4255);
or U7454 (N_7454,N_4513,N_5269);
nor U7455 (N_7455,N_5724,N_4626);
and U7456 (N_7456,N_5932,N_4425);
or U7457 (N_7457,N_5012,N_4187);
nand U7458 (N_7458,N_4682,N_5968);
nor U7459 (N_7459,N_5119,N_4591);
nor U7460 (N_7460,N_4292,N_5455);
nand U7461 (N_7461,N_5834,N_4210);
or U7462 (N_7462,N_5049,N_4491);
nand U7463 (N_7463,N_4473,N_5565);
nor U7464 (N_7464,N_5111,N_5591);
or U7465 (N_7465,N_4346,N_5500);
nand U7466 (N_7466,N_5539,N_4483);
nand U7467 (N_7467,N_4050,N_4781);
nand U7468 (N_7468,N_5807,N_4997);
or U7469 (N_7469,N_4107,N_5688);
nor U7470 (N_7470,N_5508,N_4919);
and U7471 (N_7471,N_4197,N_5395);
and U7472 (N_7472,N_4655,N_5068);
nor U7473 (N_7473,N_5986,N_5753);
nor U7474 (N_7474,N_4411,N_5767);
nor U7475 (N_7475,N_4662,N_4417);
nor U7476 (N_7476,N_4935,N_5366);
or U7477 (N_7477,N_4216,N_4036);
or U7478 (N_7478,N_5269,N_5990);
or U7479 (N_7479,N_5812,N_4455);
nand U7480 (N_7480,N_5888,N_5151);
nand U7481 (N_7481,N_4955,N_4493);
and U7482 (N_7482,N_5437,N_5609);
or U7483 (N_7483,N_5631,N_4573);
and U7484 (N_7484,N_4067,N_4127);
or U7485 (N_7485,N_4084,N_5037);
and U7486 (N_7486,N_5177,N_5276);
and U7487 (N_7487,N_4589,N_5004);
nor U7488 (N_7488,N_5776,N_5164);
and U7489 (N_7489,N_5356,N_4355);
xnor U7490 (N_7490,N_5976,N_4755);
or U7491 (N_7491,N_5947,N_5503);
and U7492 (N_7492,N_5439,N_4795);
and U7493 (N_7493,N_4281,N_5807);
nand U7494 (N_7494,N_4856,N_4098);
and U7495 (N_7495,N_4909,N_5240);
and U7496 (N_7496,N_4512,N_4364);
or U7497 (N_7497,N_5599,N_4063);
nand U7498 (N_7498,N_4818,N_5405);
nand U7499 (N_7499,N_5938,N_5606);
or U7500 (N_7500,N_5270,N_5778);
nand U7501 (N_7501,N_5158,N_4905);
nor U7502 (N_7502,N_5840,N_4036);
and U7503 (N_7503,N_4715,N_4469);
and U7504 (N_7504,N_5422,N_5822);
nor U7505 (N_7505,N_4404,N_5023);
and U7506 (N_7506,N_4299,N_4264);
nor U7507 (N_7507,N_5893,N_5469);
or U7508 (N_7508,N_4282,N_4945);
nand U7509 (N_7509,N_4301,N_5308);
nor U7510 (N_7510,N_5991,N_4245);
nand U7511 (N_7511,N_4685,N_5116);
or U7512 (N_7512,N_5521,N_4765);
or U7513 (N_7513,N_5479,N_5143);
and U7514 (N_7514,N_5406,N_4663);
nor U7515 (N_7515,N_4575,N_5895);
nand U7516 (N_7516,N_4075,N_5407);
nand U7517 (N_7517,N_5019,N_5079);
or U7518 (N_7518,N_4110,N_5857);
nand U7519 (N_7519,N_4633,N_4394);
nor U7520 (N_7520,N_5429,N_5404);
nor U7521 (N_7521,N_5606,N_5972);
nor U7522 (N_7522,N_4383,N_4120);
nor U7523 (N_7523,N_4018,N_4313);
nand U7524 (N_7524,N_4963,N_4875);
nor U7525 (N_7525,N_5928,N_4399);
and U7526 (N_7526,N_4528,N_4370);
and U7527 (N_7527,N_4388,N_4419);
or U7528 (N_7528,N_5838,N_4066);
or U7529 (N_7529,N_5196,N_5647);
and U7530 (N_7530,N_4968,N_4900);
nand U7531 (N_7531,N_5013,N_4091);
and U7532 (N_7532,N_5682,N_4826);
nor U7533 (N_7533,N_5212,N_5965);
nor U7534 (N_7534,N_5261,N_4771);
nor U7535 (N_7535,N_4566,N_5852);
and U7536 (N_7536,N_5159,N_4111);
or U7537 (N_7537,N_4663,N_5073);
nand U7538 (N_7538,N_4176,N_4363);
nand U7539 (N_7539,N_4382,N_5220);
nand U7540 (N_7540,N_4862,N_4908);
and U7541 (N_7541,N_4726,N_5641);
or U7542 (N_7542,N_5841,N_4999);
or U7543 (N_7543,N_4297,N_4244);
and U7544 (N_7544,N_5648,N_5940);
and U7545 (N_7545,N_5122,N_5313);
or U7546 (N_7546,N_4153,N_5862);
or U7547 (N_7547,N_4188,N_5512);
nand U7548 (N_7548,N_5114,N_5236);
and U7549 (N_7549,N_4564,N_4548);
or U7550 (N_7550,N_5924,N_4766);
nand U7551 (N_7551,N_5594,N_5830);
nor U7552 (N_7552,N_4790,N_5730);
or U7553 (N_7553,N_4858,N_5242);
and U7554 (N_7554,N_4405,N_5530);
and U7555 (N_7555,N_4478,N_5146);
nand U7556 (N_7556,N_5766,N_4922);
nand U7557 (N_7557,N_4934,N_4690);
and U7558 (N_7558,N_5070,N_4912);
nor U7559 (N_7559,N_5498,N_4825);
nor U7560 (N_7560,N_5470,N_5831);
or U7561 (N_7561,N_5265,N_4414);
nor U7562 (N_7562,N_4779,N_4118);
nor U7563 (N_7563,N_4346,N_4186);
nand U7564 (N_7564,N_4730,N_4251);
or U7565 (N_7565,N_5704,N_4163);
nand U7566 (N_7566,N_5965,N_4555);
or U7567 (N_7567,N_4916,N_5471);
nor U7568 (N_7568,N_4219,N_5662);
nor U7569 (N_7569,N_5132,N_4470);
or U7570 (N_7570,N_5362,N_5224);
nand U7571 (N_7571,N_4271,N_4627);
nor U7572 (N_7572,N_5703,N_5444);
or U7573 (N_7573,N_4088,N_5679);
or U7574 (N_7574,N_5514,N_5389);
nor U7575 (N_7575,N_5851,N_5216);
or U7576 (N_7576,N_5855,N_4687);
nand U7577 (N_7577,N_4200,N_4625);
and U7578 (N_7578,N_4657,N_5336);
and U7579 (N_7579,N_5980,N_4911);
nor U7580 (N_7580,N_5564,N_4479);
nand U7581 (N_7581,N_5912,N_4856);
or U7582 (N_7582,N_4308,N_5226);
nor U7583 (N_7583,N_5262,N_4226);
and U7584 (N_7584,N_5111,N_5230);
or U7585 (N_7585,N_5497,N_4002);
and U7586 (N_7586,N_4570,N_5092);
or U7587 (N_7587,N_5814,N_5366);
nor U7588 (N_7588,N_5593,N_4554);
nor U7589 (N_7589,N_4718,N_4234);
nand U7590 (N_7590,N_5638,N_4686);
nand U7591 (N_7591,N_4496,N_4646);
and U7592 (N_7592,N_5790,N_5989);
and U7593 (N_7593,N_4024,N_5674);
or U7594 (N_7594,N_4182,N_4595);
nor U7595 (N_7595,N_4294,N_5456);
or U7596 (N_7596,N_4252,N_5705);
nand U7597 (N_7597,N_4006,N_4646);
or U7598 (N_7598,N_5833,N_5242);
and U7599 (N_7599,N_4115,N_5180);
or U7600 (N_7600,N_5470,N_5344);
nor U7601 (N_7601,N_5190,N_4733);
or U7602 (N_7602,N_4877,N_4960);
and U7603 (N_7603,N_5804,N_4103);
or U7604 (N_7604,N_5696,N_4303);
and U7605 (N_7605,N_5921,N_5060);
or U7606 (N_7606,N_5228,N_5162);
and U7607 (N_7607,N_5128,N_5472);
nor U7608 (N_7608,N_4265,N_4530);
nor U7609 (N_7609,N_4889,N_4427);
nand U7610 (N_7610,N_5926,N_4325);
nor U7611 (N_7611,N_4894,N_5805);
nor U7612 (N_7612,N_5833,N_5979);
and U7613 (N_7613,N_4414,N_4430);
nor U7614 (N_7614,N_5406,N_5026);
and U7615 (N_7615,N_5408,N_5120);
and U7616 (N_7616,N_4981,N_4701);
and U7617 (N_7617,N_5713,N_4469);
and U7618 (N_7618,N_4409,N_4053);
nor U7619 (N_7619,N_5951,N_4488);
and U7620 (N_7620,N_5705,N_5285);
or U7621 (N_7621,N_5030,N_4858);
nor U7622 (N_7622,N_4858,N_4438);
nand U7623 (N_7623,N_4395,N_4453);
or U7624 (N_7624,N_5130,N_5109);
nor U7625 (N_7625,N_5653,N_4383);
nand U7626 (N_7626,N_5700,N_4158);
or U7627 (N_7627,N_4515,N_4933);
nor U7628 (N_7628,N_5950,N_4706);
or U7629 (N_7629,N_4493,N_4011);
nand U7630 (N_7630,N_4455,N_5332);
nand U7631 (N_7631,N_5208,N_5316);
nand U7632 (N_7632,N_5555,N_4368);
and U7633 (N_7633,N_4086,N_4043);
and U7634 (N_7634,N_4350,N_4062);
and U7635 (N_7635,N_4402,N_5124);
nor U7636 (N_7636,N_5029,N_4629);
or U7637 (N_7637,N_4436,N_4463);
or U7638 (N_7638,N_5445,N_5996);
nand U7639 (N_7639,N_5287,N_5166);
nor U7640 (N_7640,N_5838,N_5719);
or U7641 (N_7641,N_5644,N_5276);
nand U7642 (N_7642,N_5824,N_5795);
nor U7643 (N_7643,N_4203,N_5764);
and U7644 (N_7644,N_4074,N_5361);
nand U7645 (N_7645,N_4666,N_4821);
nand U7646 (N_7646,N_5680,N_5078);
and U7647 (N_7647,N_5781,N_5068);
nor U7648 (N_7648,N_5461,N_5589);
and U7649 (N_7649,N_5322,N_4187);
nand U7650 (N_7650,N_4792,N_5975);
nand U7651 (N_7651,N_5660,N_5167);
and U7652 (N_7652,N_5937,N_5735);
or U7653 (N_7653,N_4417,N_4115);
nand U7654 (N_7654,N_5544,N_4175);
nor U7655 (N_7655,N_4361,N_4184);
nor U7656 (N_7656,N_5284,N_4907);
or U7657 (N_7657,N_4129,N_5373);
nor U7658 (N_7658,N_5013,N_5481);
or U7659 (N_7659,N_4107,N_5793);
nand U7660 (N_7660,N_5362,N_4777);
or U7661 (N_7661,N_5121,N_4369);
and U7662 (N_7662,N_5698,N_5507);
or U7663 (N_7663,N_5156,N_5160);
or U7664 (N_7664,N_5507,N_4922);
and U7665 (N_7665,N_4614,N_4009);
nor U7666 (N_7666,N_4985,N_5763);
and U7667 (N_7667,N_5594,N_4823);
or U7668 (N_7668,N_5652,N_5698);
and U7669 (N_7669,N_4153,N_5788);
or U7670 (N_7670,N_4450,N_4480);
or U7671 (N_7671,N_5841,N_5765);
or U7672 (N_7672,N_5226,N_5825);
nand U7673 (N_7673,N_5553,N_5059);
nand U7674 (N_7674,N_4852,N_5891);
or U7675 (N_7675,N_5493,N_4295);
and U7676 (N_7676,N_4571,N_5428);
or U7677 (N_7677,N_5362,N_5814);
nor U7678 (N_7678,N_5596,N_5665);
nand U7679 (N_7679,N_4674,N_5924);
nand U7680 (N_7680,N_4466,N_5786);
and U7681 (N_7681,N_5238,N_5727);
or U7682 (N_7682,N_5880,N_4515);
nand U7683 (N_7683,N_4043,N_5896);
nor U7684 (N_7684,N_4228,N_5024);
nor U7685 (N_7685,N_5292,N_5012);
nand U7686 (N_7686,N_4971,N_5077);
and U7687 (N_7687,N_4531,N_5665);
and U7688 (N_7688,N_5397,N_4032);
nor U7689 (N_7689,N_4207,N_5387);
nor U7690 (N_7690,N_4653,N_5615);
and U7691 (N_7691,N_4971,N_5789);
and U7692 (N_7692,N_5446,N_5297);
nor U7693 (N_7693,N_5959,N_5310);
nand U7694 (N_7694,N_5374,N_4123);
or U7695 (N_7695,N_5963,N_4041);
or U7696 (N_7696,N_4903,N_5579);
or U7697 (N_7697,N_4680,N_4030);
nor U7698 (N_7698,N_5104,N_5903);
nand U7699 (N_7699,N_5755,N_5270);
or U7700 (N_7700,N_4766,N_4146);
or U7701 (N_7701,N_4711,N_5960);
or U7702 (N_7702,N_4208,N_5516);
nand U7703 (N_7703,N_4104,N_4902);
nor U7704 (N_7704,N_5717,N_5468);
nand U7705 (N_7705,N_5142,N_4484);
nor U7706 (N_7706,N_5723,N_4960);
nor U7707 (N_7707,N_4313,N_4588);
or U7708 (N_7708,N_4818,N_5859);
nand U7709 (N_7709,N_5039,N_4767);
nand U7710 (N_7710,N_4825,N_4312);
and U7711 (N_7711,N_5840,N_5563);
or U7712 (N_7712,N_5748,N_4057);
nand U7713 (N_7713,N_4294,N_4615);
nor U7714 (N_7714,N_4568,N_5623);
and U7715 (N_7715,N_5444,N_4903);
and U7716 (N_7716,N_5200,N_5932);
nor U7717 (N_7717,N_4072,N_5373);
and U7718 (N_7718,N_5153,N_4297);
and U7719 (N_7719,N_4162,N_4147);
nand U7720 (N_7720,N_4818,N_4135);
nor U7721 (N_7721,N_5545,N_5755);
and U7722 (N_7722,N_4639,N_5377);
or U7723 (N_7723,N_5560,N_5349);
nor U7724 (N_7724,N_5863,N_5574);
nor U7725 (N_7725,N_5406,N_4777);
nand U7726 (N_7726,N_4555,N_4170);
nor U7727 (N_7727,N_4448,N_4648);
or U7728 (N_7728,N_4067,N_4988);
or U7729 (N_7729,N_4228,N_5742);
and U7730 (N_7730,N_4356,N_4902);
or U7731 (N_7731,N_5246,N_4926);
and U7732 (N_7732,N_4351,N_4438);
nand U7733 (N_7733,N_4377,N_4591);
nor U7734 (N_7734,N_4398,N_5367);
or U7735 (N_7735,N_4722,N_4155);
nand U7736 (N_7736,N_5711,N_5166);
or U7737 (N_7737,N_5987,N_4601);
or U7738 (N_7738,N_4243,N_4147);
or U7739 (N_7739,N_5359,N_4300);
or U7740 (N_7740,N_4448,N_4858);
and U7741 (N_7741,N_4928,N_5421);
and U7742 (N_7742,N_4726,N_5101);
nor U7743 (N_7743,N_4092,N_5737);
nand U7744 (N_7744,N_5423,N_4108);
nor U7745 (N_7745,N_4570,N_4539);
or U7746 (N_7746,N_4123,N_4461);
nand U7747 (N_7747,N_4725,N_5764);
nor U7748 (N_7748,N_4604,N_4754);
or U7749 (N_7749,N_4787,N_4782);
or U7750 (N_7750,N_4468,N_4492);
and U7751 (N_7751,N_5349,N_5851);
nand U7752 (N_7752,N_5326,N_4170);
and U7753 (N_7753,N_4753,N_5925);
nand U7754 (N_7754,N_5871,N_4170);
nand U7755 (N_7755,N_4413,N_5328);
and U7756 (N_7756,N_5477,N_5539);
and U7757 (N_7757,N_5744,N_5327);
or U7758 (N_7758,N_5745,N_4695);
or U7759 (N_7759,N_4897,N_5567);
nor U7760 (N_7760,N_4888,N_5153);
or U7761 (N_7761,N_4789,N_5858);
nand U7762 (N_7762,N_4465,N_4755);
or U7763 (N_7763,N_4767,N_5404);
nand U7764 (N_7764,N_4699,N_5717);
or U7765 (N_7765,N_4627,N_5206);
nor U7766 (N_7766,N_5205,N_4363);
nor U7767 (N_7767,N_5564,N_4227);
and U7768 (N_7768,N_4273,N_5577);
or U7769 (N_7769,N_5410,N_4739);
nand U7770 (N_7770,N_4352,N_5000);
and U7771 (N_7771,N_4819,N_5966);
nand U7772 (N_7772,N_4060,N_5189);
nor U7773 (N_7773,N_4984,N_5428);
nand U7774 (N_7774,N_4368,N_5207);
nand U7775 (N_7775,N_5432,N_5197);
and U7776 (N_7776,N_4814,N_4400);
nor U7777 (N_7777,N_4474,N_5485);
nand U7778 (N_7778,N_5224,N_5866);
nand U7779 (N_7779,N_4897,N_5789);
and U7780 (N_7780,N_4978,N_4769);
nand U7781 (N_7781,N_4614,N_4909);
nor U7782 (N_7782,N_5138,N_4305);
nor U7783 (N_7783,N_5916,N_4542);
or U7784 (N_7784,N_4971,N_4537);
nor U7785 (N_7785,N_5582,N_5702);
nand U7786 (N_7786,N_4559,N_4823);
nor U7787 (N_7787,N_4498,N_5208);
nand U7788 (N_7788,N_5820,N_5065);
nand U7789 (N_7789,N_4499,N_5714);
nor U7790 (N_7790,N_4835,N_4490);
nand U7791 (N_7791,N_4976,N_4062);
nor U7792 (N_7792,N_4891,N_5373);
and U7793 (N_7793,N_5142,N_5659);
and U7794 (N_7794,N_5020,N_5769);
and U7795 (N_7795,N_4005,N_4982);
and U7796 (N_7796,N_4813,N_4406);
and U7797 (N_7797,N_5204,N_5855);
nand U7798 (N_7798,N_4301,N_4864);
or U7799 (N_7799,N_5761,N_5675);
or U7800 (N_7800,N_4127,N_4612);
or U7801 (N_7801,N_5214,N_4139);
nor U7802 (N_7802,N_4815,N_4998);
or U7803 (N_7803,N_5899,N_4250);
and U7804 (N_7804,N_5133,N_5995);
nand U7805 (N_7805,N_5622,N_4840);
or U7806 (N_7806,N_4864,N_4428);
nand U7807 (N_7807,N_4075,N_4848);
and U7808 (N_7808,N_5664,N_5731);
and U7809 (N_7809,N_5672,N_5819);
and U7810 (N_7810,N_5451,N_5733);
nor U7811 (N_7811,N_5428,N_5645);
nand U7812 (N_7812,N_5204,N_5530);
or U7813 (N_7813,N_4317,N_4926);
and U7814 (N_7814,N_4322,N_4947);
xnor U7815 (N_7815,N_5540,N_4739);
and U7816 (N_7816,N_4138,N_4113);
and U7817 (N_7817,N_5939,N_5007);
nand U7818 (N_7818,N_5084,N_5889);
or U7819 (N_7819,N_4012,N_4756);
or U7820 (N_7820,N_4383,N_5350);
xnor U7821 (N_7821,N_5819,N_5953);
nor U7822 (N_7822,N_4244,N_5407);
nor U7823 (N_7823,N_4215,N_5884);
or U7824 (N_7824,N_5278,N_4632);
nor U7825 (N_7825,N_5700,N_4160);
nand U7826 (N_7826,N_4961,N_5632);
xor U7827 (N_7827,N_5971,N_5701);
nand U7828 (N_7828,N_5828,N_5451);
nand U7829 (N_7829,N_4314,N_5728);
or U7830 (N_7830,N_5752,N_4107);
or U7831 (N_7831,N_4208,N_5507);
nand U7832 (N_7832,N_4404,N_5170);
and U7833 (N_7833,N_4017,N_4885);
nand U7834 (N_7834,N_5620,N_5084);
xnor U7835 (N_7835,N_5384,N_5610);
or U7836 (N_7836,N_5695,N_4424);
or U7837 (N_7837,N_4808,N_5263);
or U7838 (N_7838,N_5831,N_4797);
or U7839 (N_7839,N_5031,N_5353);
nand U7840 (N_7840,N_5139,N_5213);
nand U7841 (N_7841,N_4810,N_5352);
nand U7842 (N_7842,N_4133,N_5963);
nor U7843 (N_7843,N_5933,N_5173);
nor U7844 (N_7844,N_5262,N_5280);
and U7845 (N_7845,N_4096,N_4261);
nand U7846 (N_7846,N_4262,N_4000);
and U7847 (N_7847,N_4524,N_4892);
nand U7848 (N_7848,N_5970,N_4784);
nand U7849 (N_7849,N_4603,N_5744);
nor U7850 (N_7850,N_4221,N_4413);
nor U7851 (N_7851,N_5691,N_4952);
and U7852 (N_7852,N_4502,N_5413);
nor U7853 (N_7853,N_4591,N_5036);
nor U7854 (N_7854,N_4610,N_5160);
nand U7855 (N_7855,N_4259,N_4990);
nor U7856 (N_7856,N_5676,N_5622);
and U7857 (N_7857,N_4853,N_4217);
nand U7858 (N_7858,N_4225,N_5352);
nand U7859 (N_7859,N_5720,N_4743);
or U7860 (N_7860,N_4110,N_5682);
nor U7861 (N_7861,N_4984,N_4059);
and U7862 (N_7862,N_4392,N_5781);
nand U7863 (N_7863,N_5931,N_4785);
xnor U7864 (N_7864,N_4211,N_4331);
and U7865 (N_7865,N_4848,N_4712);
and U7866 (N_7866,N_5016,N_5535);
nand U7867 (N_7867,N_4823,N_4487);
nor U7868 (N_7868,N_5291,N_4379);
nand U7869 (N_7869,N_5027,N_5699);
nor U7870 (N_7870,N_4930,N_4255);
or U7871 (N_7871,N_5261,N_5787);
and U7872 (N_7872,N_5603,N_5897);
nor U7873 (N_7873,N_5969,N_4588);
and U7874 (N_7874,N_4426,N_4332);
nor U7875 (N_7875,N_5227,N_5781);
and U7876 (N_7876,N_4948,N_4473);
nand U7877 (N_7877,N_4984,N_4045);
nor U7878 (N_7878,N_4336,N_4654);
nand U7879 (N_7879,N_5673,N_4787);
nor U7880 (N_7880,N_5725,N_4328);
and U7881 (N_7881,N_4193,N_4240);
nand U7882 (N_7882,N_5193,N_5252);
or U7883 (N_7883,N_5653,N_5481);
nand U7884 (N_7884,N_5145,N_5616);
nand U7885 (N_7885,N_4204,N_5635);
nor U7886 (N_7886,N_4748,N_4956);
and U7887 (N_7887,N_5392,N_5518);
and U7888 (N_7888,N_5113,N_4028);
or U7889 (N_7889,N_5045,N_4426);
or U7890 (N_7890,N_5251,N_4736);
nand U7891 (N_7891,N_4243,N_5292);
and U7892 (N_7892,N_5042,N_5216);
or U7893 (N_7893,N_5978,N_4598);
or U7894 (N_7894,N_5264,N_4611);
nor U7895 (N_7895,N_5979,N_5625);
and U7896 (N_7896,N_5967,N_4221);
xnor U7897 (N_7897,N_4209,N_4727);
and U7898 (N_7898,N_4740,N_4060);
and U7899 (N_7899,N_5135,N_4741);
nor U7900 (N_7900,N_5525,N_5395);
nand U7901 (N_7901,N_4832,N_5581);
or U7902 (N_7902,N_4026,N_5546);
or U7903 (N_7903,N_5465,N_4555);
and U7904 (N_7904,N_5700,N_4056);
nand U7905 (N_7905,N_5279,N_5804);
nand U7906 (N_7906,N_5465,N_5787);
and U7907 (N_7907,N_4860,N_4452);
nand U7908 (N_7908,N_4413,N_5730);
nand U7909 (N_7909,N_5086,N_5183);
and U7910 (N_7910,N_5806,N_5479);
nand U7911 (N_7911,N_5537,N_4157);
nand U7912 (N_7912,N_5803,N_5250);
or U7913 (N_7913,N_4168,N_4649);
or U7914 (N_7914,N_4316,N_4236);
nand U7915 (N_7915,N_5748,N_4522);
and U7916 (N_7916,N_4343,N_5524);
and U7917 (N_7917,N_4658,N_4997);
xor U7918 (N_7918,N_5175,N_5362);
and U7919 (N_7919,N_4007,N_4594);
nand U7920 (N_7920,N_4414,N_5869);
or U7921 (N_7921,N_4325,N_5622);
or U7922 (N_7922,N_5458,N_4026);
or U7923 (N_7923,N_4481,N_4804);
nand U7924 (N_7924,N_5122,N_4366);
nor U7925 (N_7925,N_4047,N_5485);
nor U7926 (N_7926,N_4464,N_5557);
and U7927 (N_7927,N_5236,N_5989);
or U7928 (N_7928,N_5134,N_5436);
nor U7929 (N_7929,N_5138,N_4216);
nor U7930 (N_7930,N_5141,N_5114);
and U7931 (N_7931,N_5187,N_5281);
nor U7932 (N_7932,N_5735,N_5064);
nand U7933 (N_7933,N_4861,N_5532);
nor U7934 (N_7934,N_5171,N_4852);
nand U7935 (N_7935,N_5224,N_4878);
xnor U7936 (N_7936,N_4724,N_4026);
nor U7937 (N_7937,N_4805,N_5347);
nor U7938 (N_7938,N_5161,N_5079);
or U7939 (N_7939,N_5158,N_4500);
and U7940 (N_7940,N_5396,N_4931);
nor U7941 (N_7941,N_4530,N_5742);
and U7942 (N_7942,N_4005,N_4705);
nand U7943 (N_7943,N_5649,N_5900);
nor U7944 (N_7944,N_4850,N_5756);
nand U7945 (N_7945,N_4195,N_5018);
nor U7946 (N_7946,N_5683,N_5602);
or U7947 (N_7947,N_4352,N_4156);
or U7948 (N_7948,N_4306,N_4664);
nand U7949 (N_7949,N_5418,N_5739);
nor U7950 (N_7950,N_4863,N_5877);
or U7951 (N_7951,N_4033,N_5268);
nand U7952 (N_7952,N_5299,N_5695);
or U7953 (N_7953,N_4318,N_4717);
nor U7954 (N_7954,N_5440,N_5778);
nand U7955 (N_7955,N_4584,N_5193);
or U7956 (N_7956,N_5245,N_5987);
nand U7957 (N_7957,N_4478,N_4607);
and U7958 (N_7958,N_5470,N_4819);
and U7959 (N_7959,N_5546,N_4514);
nand U7960 (N_7960,N_5656,N_4256);
or U7961 (N_7961,N_5982,N_4736);
nand U7962 (N_7962,N_4056,N_4775);
nor U7963 (N_7963,N_4437,N_4310);
nor U7964 (N_7964,N_4471,N_5011);
nor U7965 (N_7965,N_5822,N_4670);
nand U7966 (N_7966,N_4901,N_5673);
nand U7967 (N_7967,N_5965,N_4757);
nor U7968 (N_7968,N_5595,N_5143);
nand U7969 (N_7969,N_5019,N_4961);
or U7970 (N_7970,N_5301,N_5615);
or U7971 (N_7971,N_4747,N_5813);
nor U7972 (N_7972,N_5759,N_5616);
and U7973 (N_7973,N_4994,N_4616);
nand U7974 (N_7974,N_5370,N_5967);
nor U7975 (N_7975,N_4300,N_5281);
or U7976 (N_7976,N_4472,N_4756);
and U7977 (N_7977,N_5376,N_5383);
and U7978 (N_7978,N_5356,N_5487);
nor U7979 (N_7979,N_5497,N_5962);
and U7980 (N_7980,N_4055,N_4777);
nand U7981 (N_7981,N_4275,N_4814);
nand U7982 (N_7982,N_5621,N_4214);
nand U7983 (N_7983,N_5942,N_5894);
nor U7984 (N_7984,N_4731,N_5974);
nor U7985 (N_7985,N_4599,N_5385);
xor U7986 (N_7986,N_5879,N_4259);
nand U7987 (N_7987,N_4717,N_5254);
or U7988 (N_7988,N_5469,N_5479);
and U7989 (N_7989,N_4104,N_5041);
nand U7990 (N_7990,N_4094,N_5755);
or U7991 (N_7991,N_4665,N_5474);
or U7992 (N_7992,N_5664,N_5022);
and U7993 (N_7993,N_4075,N_5671);
nand U7994 (N_7994,N_4456,N_5488);
nor U7995 (N_7995,N_5530,N_5420);
nor U7996 (N_7996,N_5531,N_5702);
nand U7997 (N_7997,N_4296,N_5540);
nand U7998 (N_7998,N_5671,N_5992);
and U7999 (N_7999,N_4838,N_4752);
or U8000 (N_8000,N_6795,N_7186);
nand U8001 (N_8001,N_6265,N_7851);
nor U8002 (N_8002,N_6197,N_7165);
and U8003 (N_8003,N_7459,N_6561);
and U8004 (N_8004,N_6010,N_6823);
and U8005 (N_8005,N_7502,N_7416);
or U8006 (N_8006,N_7290,N_7021);
nand U8007 (N_8007,N_6152,N_7286);
and U8008 (N_8008,N_6635,N_7526);
nand U8009 (N_8009,N_7027,N_7926);
or U8010 (N_8010,N_6456,N_7220);
and U8011 (N_8011,N_6579,N_6689);
nor U8012 (N_8012,N_6644,N_6298);
nand U8013 (N_8013,N_7256,N_7732);
xor U8014 (N_8014,N_7744,N_7966);
or U8015 (N_8015,N_6072,N_6826);
nor U8016 (N_8016,N_6380,N_7728);
or U8017 (N_8017,N_7706,N_6590);
and U8018 (N_8018,N_6700,N_7367);
nor U8019 (N_8019,N_6078,N_6271);
nand U8020 (N_8020,N_7661,N_7497);
or U8021 (N_8021,N_7109,N_7203);
nor U8022 (N_8022,N_6522,N_6601);
nand U8023 (N_8023,N_7140,N_7542);
xor U8024 (N_8024,N_6482,N_6731);
and U8025 (N_8025,N_6486,N_7360);
nand U8026 (N_8026,N_7099,N_7339);
and U8027 (N_8027,N_6870,N_6841);
nand U8028 (N_8028,N_7805,N_6300);
or U8029 (N_8029,N_7535,N_7260);
nand U8030 (N_8030,N_7052,N_7415);
nand U8031 (N_8031,N_6762,N_7869);
nor U8032 (N_8032,N_7493,N_7714);
nor U8033 (N_8033,N_6773,N_7187);
nand U8034 (N_8034,N_6118,N_7531);
and U8035 (N_8035,N_7619,N_6819);
nor U8036 (N_8036,N_6704,N_6965);
and U8037 (N_8037,N_7891,N_7268);
nand U8038 (N_8038,N_7469,N_6939);
and U8039 (N_8039,N_7825,N_7972);
nand U8040 (N_8040,N_6085,N_7738);
or U8041 (N_8041,N_6835,N_7467);
or U8042 (N_8042,N_6181,N_7918);
nor U8043 (N_8043,N_6126,N_6595);
or U8044 (N_8044,N_7568,N_7720);
or U8045 (N_8045,N_6972,N_7337);
nor U8046 (N_8046,N_6370,N_6260);
nand U8047 (N_8047,N_6283,N_7422);
or U8048 (N_8048,N_7802,N_7973);
xor U8049 (N_8049,N_7201,N_7277);
nor U8050 (N_8050,N_7997,N_7250);
or U8051 (N_8051,N_7060,N_6004);
nor U8052 (N_8052,N_6887,N_6089);
or U8053 (N_8053,N_7451,N_7346);
and U8054 (N_8054,N_6099,N_7480);
nor U8055 (N_8055,N_6792,N_7310);
nand U8056 (N_8056,N_7832,N_6041);
nor U8057 (N_8057,N_6481,N_7300);
nor U8058 (N_8058,N_6431,N_7734);
and U8059 (N_8059,N_6882,N_6788);
nor U8060 (N_8060,N_6301,N_6050);
or U8061 (N_8061,N_6065,N_6473);
nand U8062 (N_8062,N_6307,N_7879);
and U8063 (N_8063,N_7331,N_7767);
or U8064 (N_8064,N_7089,N_7287);
nor U8065 (N_8065,N_7715,N_7653);
and U8066 (N_8066,N_6386,N_6613);
or U8067 (N_8067,N_6190,N_6504);
or U8068 (N_8068,N_7597,N_6142);
nand U8069 (N_8069,N_6937,N_7830);
nand U8070 (N_8070,N_7281,N_7991);
nor U8071 (N_8071,N_7944,N_6999);
xor U8072 (N_8072,N_7115,N_6318);
nor U8073 (N_8073,N_7192,N_7026);
and U8074 (N_8074,N_6991,N_7387);
nor U8075 (N_8075,N_7611,N_6311);
nand U8076 (N_8076,N_7334,N_7325);
nand U8077 (N_8077,N_7782,N_7092);
or U8078 (N_8078,N_6694,N_7838);
nand U8079 (N_8079,N_7769,N_6061);
nor U8080 (N_8080,N_7839,N_6114);
nand U8081 (N_8081,N_7697,N_7080);
or U8082 (N_8082,N_7309,N_6852);
nand U8083 (N_8083,N_6828,N_6611);
nand U8084 (N_8084,N_7071,N_6912);
xor U8085 (N_8085,N_6450,N_7410);
nand U8086 (N_8086,N_6638,N_7279);
nand U8087 (N_8087,N_6840,N_7970);
nor U8088 (N_8088,N_7584,N_6183);
nor U8089 (N_8089,N_6376,N_6323);
nor U8090 (N_8090,N_6393,N_7401);
or U8091 (N_8091,N_7053,N_6657);
nand U8092 (N_8092,N_6096,N_6603);
nor U8093 (N_8093,N_7793,N_6645);
xor U8094 (N_8094,N_6862,N_6199);
nand U8095 (N_8095,N_7960,N_7341);
and U8096 (N_8096,N_7432,N_7875);
and U8097 (N_8097,N_7116,N_7986);
nand U8098 (N_8098,N_6620,N_7847);
nor U8099 (N_8099,N_7441,N_6916);
or U8100 (N_8100,N_7788,N_7554);
nor U8101 (N_8101,N_7274,N_6173);
nor U8102 (N_8102,N_7583,N_6392);
nor U8103 (N_8103,N_6411,N_6746);
or U8104 (N_8104,N_6684,N_6772);
nand U8105 (N_8105,N_7481,N_6924);
nor U8106 (N_8106,N_6629,N_6902);
nand U8107 (N_8107,N_6453,N_6637);
nor U8108 (N_8108,N_7942,N_6572);
and U8109 (N_8109,N_6817,N_6593);
nand U8110 (N_8110,N_7166,N_7100);
nand U8111 (N_8111,N_6354,N_6060);
or U8112 (N_8112,N_7063,N_7385);
and U8113 (N_8113,N_6594,N_7984);
or U8114 (N_8114,N_6653,N_7555);
or U8115 (N_8115,N_7082,N_6258);
nand U8116 (N_8116,N_6727,N_7212);
and U8117 (N_8117,N_7707,N_6996);
nor U8118 (N_8118,N_6812,N_7664);
and U8119 (N_8119,N_6586,N_6209);
nor U8120 (N_8120,N_7029,N_6867);
or U8121 (N_8121,N_7428,N_7392);
or U8122 (N_8122,N_6102,N_7488);
nor U8123 (N_8123,N_7292,N_7076);
and U8124 (N_8124,N_6668,N_6455);
and U8125 (N_8125,N_6331,N_6496);
or U8126 (N_8126,N_6945,N_6702);
or U8127 (N_8127,N_6294,N_6641);
and U8128 (N_8128,N_6110,N_6843);
or U8129 (N_8129,N_6967,N_6277);
nand U8130 (N_8130,N_7755,N_7215);
nand U8131 (N_8131,N_7307,N_7864);
and U8132 (N_8132,N_6753,N_6926);
nor U8133 (N_8133,N_7579,N_6013);
or U8134 (N_8134,N_6970,N_6137);
nand U8135 (N_8135,N_7421,N_7022);
or U8136 (N_8136,N_6591,N_7735);
nand U8137 (N_8137,N_7238,N_6674);
nor U8138 (N_8138,N_7686,N_6597);
or U8139 (N_8139,N_7153,N_6315);
or U8140 (N_8140,N_6745,N_7983);
or U8141 (N_8141,N_7491,N_7721);
or U8142 (N_8142,N_7400,N_7204);
nor U8143 (N_8143,N_7362,N_6950);
nand U8144 (N_8144,N_7097,N_6712);
nor U8145 (N_8145,N_7407,N_6176);
or U8146 (N_8146,N_7070,N_7709);
nand U8147 (N_8147,N_6871,N_7976);
nand U8148 (N_8148,N_7935,N_7898);
nand U8149 (N_8149,N_6309,N_7678);
nor U8150 (N_8150,N_6328,N_7396);
xnor U8151 (N_8151,N_7477,N_6037);
nor U8152 (N_8152,N_7899,N_7179);
nand U8153 (N_8153,N_6441,N_7807);
nor U8154 (N_8154,N_6313,N_6723);
nand U8155 (N_8155,N_6241,N_6989);
xnor U8156 (N_8156,N_7137,N_7573);
and U8157 (N_8157,N_6440,N_7448);
and U8158 (N_8158,N_6346,N_7431);
and U8159 (N_8159,N_7595,N_6350);
nand U8160 (N_8160,N_6454,N_7656);
nand U8161 (N_8161,N_6351,N_6851);
or U8162 (N_8162,N_7110,N_6555);
or U8163 (N_8163,N_6514,N_6632);
nand U8164 (N_8164,N_7787,N_7083);
or U8165 (N_8165,N_7023,N_7327);
and U8166 (N_8166,N_7336,N_7282);
nand U8167 (N_8167,N_6774,N_6742);
and U8168 (N_8168,N_7181,N_6216);
or U8169 (N_8169,N_7642,N_6364);
and U8170 (N_8170,N_7740,N_6825);
nand U8171 (N_8171,N_6776,N_6739);
nor U8172 (N_8172,N_7081,N_6266);
nor U8173 (N_8173,N_6129,N_6439);
nor U8174 (N_8174,N_7106,N_7230);
nor U8175 (N_8175,N_6535,N_6711);
or U8176 (N_8176,N_6659,N_6278);
nand U8177 (N_8177,N_7501,N_6680);
and U8178 (N_8178,N_6108,N_7848);
nand U8179 (N_8179,N_7602,N_6730);
nor U8180 (N_8180,N_7378,N_6302);
and U8181 (N_8181,N_6856,N_6803);
or U8182 (N_8182,N_6539,N_6565);
nand U8183 (N_8183,N_7885,N_6786);
and U8184 (N_8184,N_7638,N_7121);
or U8185 (N_8185,N_6771,N_7996);
and U8186 (N_8186,N_6269,N_7958);
or U8187 (N_8187,N_6047,N_6575);
nor U8188 (N_8188,N_6284,N_7645);
or U8189 (N_8189,N_6896,N_7919);
and U8190 (N_8190,N_6703,N_6459);
nand U8191 (N_8191,N_6663,N_6449);
nor U8192 (N_8192,N_6566,N_6042);
and U8193 (N_8193,N_7739,N_6526);
or U8194 (N_8194,N_6073,N_6097);
or U8195 (N_8195,N_7833,N_7527);
or U8196 (N_8196,N_7357,N_6818);
nand U8197 (N_8197,N_7677,N_7746);
nand U8198 (N_8198,N_6732,N_7954);
nor U8199 (N_8199,N_7024,N_7999);
xor U8200 (N_8200,N_6317,N_7061);
or U8201 (N_8201,N_7945,N_6192);
nor U8202 (N_8202,N_6813,N_7532);
and U8203 (N_8203,N_6884,N_7790);
and U8204 (N_8204,N_7852,N_7130);
and U8205 (N_8205,N_6985,N_7688);
nand U8206 (N_8206,N_7067,N_7540);
nand U8207 (N_8207,N_7444,N_7601);
nand U8208 (N_8208,N_6292,N_7759);
and U8209 (N_8209,N_6669,N_6503);
and U8210 (N_8210,N_6760,N_6027);
xor U8211 (N_8211,N_7786,N_7373);
and U8212 (N_8212,N_6787,N_6132);
nor U8213 (N_8213,N_7837,N_7921);
nor U8214 (N_8214,N_7162,N_6305);
or U8215 (N_8215,N_6428,N_7939);
or U8216 (N_8216,N_6296,N_7988);
and U8217 (N_8217,N_7580,N_6343);
and U8218 (N_8218,N_6978,N_6515);
nand U8219 (N_8219,N_6264,N_7030);
or U8220 (N_8220,N_6255,N_6903);
nand U8221 (N_8221,N_7364,N_6665);
nor U8222 (N_8222,N_7870,N_6658);
and U8223 (N_8223,N_7409,N_7056);
nor U8224 (N_8224,N_7783,N_6600);
or U8225 (N_8225,N_7271,N_7667);
and U8226 (N_8226,N_7980,N_6465);
or U8227 (N_8227,N_6675,N_6009);
nand U8228 (N_8228,N_7452,N_6366);
or U8229 (N_8229,N_7668,N_6942);
nand U8230 (N_8230,N_7154,N_6589);
or U8231 (N_8231,N_6673,N_7150);
or U8232 (N_8232,N_6766,N_6827);
and U8233 (N_8233,N_7625,N_6157);
xnor U8234 (N_8234,N_6627,N_6966);
nor U8235 (N_8235,N_6372,N_7332);
and U8236 (N_8236,N_7761,N_6604);
and U8237 (N_8237,N_7299,N_7840);
nor U8238 (N_8238,N_7445,N_6218);
and U8239 (N_8239,N_7095,N_6164);
nor U8240 (N_8240,N_6034,N_6430);
nand U8241 (N_8241,N_6713,N_7992);
nor U8242 (N_8242,N_7222,N_6532);
nand U8243 (N_8243,N_7589,N_7388);
nor U8244 (N_8244,N_7375,N_7824);
xor U8245 (N_8245,N_6560,N_7188);
or U8246 (N_8246,N_7486,N_7032);
and U8247 (N_8247,N_7485,N_7841);
and U8248 (N_8248,N_7529,N_6246);
or U8249 (N_8249,N_7365,N_7125);
nand U8250 (N_8250,N_6934,N_6876);
and U8251 (N_8251,N_7672,N_6375);
and U8252 (N_8252,N_6281,N_7647);
and U8253 (N_8253,N_6239,N_7685);
or U8254 (N_8254,N_7120,N_6425);
nand U8255 (N_8255,N_7247,N_7995);
nand U8256 (N_8256,N_6094,N_7436);
and U8257 (N_8257,N_6518,N_6634);
nand U8258 (N_8258,N_6121,N_7046);
nor U8259 (N_8259,N_7406,N_6576);
nor U8260 (N_8260,N_6419,N_7363);
and U8261 (N_8261,N_7005,N_6633);
or U8262 (N_8262,N_6549,N_6784);
nor U8263 (N_8263,N_6193,N_6074);
nand U8264 (N_8264,N_6697,N_6385);
nor U8265 (N_8265,N_6329,N_7940);
nand U8266 (N_8266,N_6930,N_6794);
nand U8267 (N_8267,N_6754,N_7135);
nor U8268 (N_8268,N_6617,N_7171);
or U8269 (N_8269,N_6039,N_6326);
nor U8270 (N_8270,N_7141,N_6626);
or U8271 (N_8271,N_6799,N_6736);
and U8272 (N_8272,N_6347,N_7967);
nor U8273 (N_8273,N_7794,N_6420);
and U8274 (N_8274,N_6605,N_6223);
and U8275 (N_8275,N_7408,N_6769);
nand U8276 (N_8276,N_7896,N_7016);
nor U8277 (N_8277,N_6915,N_6112);
and U8278 (N_8278,N_6960,N_7598);
or U8279 (N_8279,N_7207,N_6435);
or U8280 (N_8280,N_6136,N_7311);
nor U8281 (N_8281,N_6306,N_6184);
nor U8282 (N_8282,N_6342,N_7610);
nor U8283 (N_8283,N_7713,N_6396);
or U8284 (N_8284,N_6369,N_7284);
and U8285 (N_8285,N_6820,N_7159);
or U8286 (N_8286,N_7644,N_6761);
or U8287 (N_8287,N_7433,N_6768);
nand U8288 (N_8288,N_6213,N_7742);
nand U8289 (N_8289,N_7893,N_7169);
nand U8290 (N_8290,N_7572,N_7934);
nor U8291 (N_8291,N_6524,N_7102);
nor U8292 (N_8292,N_6415,N_6242);
nor U8293 (N_8293,N_6451,N_7887);
nor U8294 (N_8294,N_6172,N_6563);
nor U8295 (N_8295,N_6686,N_6071);
nor U8296 (N_8296,N_7434,N_6869);
nand U8297 (N_8297,N_7087,N_7276);
nand U8298 (N_8298,N_6954,N_7062);
nand U8299 (N_8299,N_6195,N_7425);
nor U8300 (N_8300,N_7231,N_7041);
and U8301 (N_8301,N_6161,N_7058);
nand U8302 (N_8302,N_7132,N_7103);
nor U8303 (N_8303,N_6452,N_7161);
and U8304 (N_8304,N_7640,N_7711);
or U8305 (N_8305,N_6297,N_7539);
or U8306 (N_8306,N_6839,N_7265);
and U8307 (N_8307,N_6837,N_7324);
and U8308 (N_8308,N_6012,N_7189);
or U8309 (N_8309,N_7679,N_7209);
or U8310 (N_8310,N_7578,N_6188);
nor U8311 (N_8311,N_7000,N_7004);
nor U8312 (N_8312,N_7612,N_7698);
nand U8313 (N_8313,N_6763,N_6357);
or U8314 (N_8314,N_7468,N_7733);
or U8315 (N_8315,N_7516,N_7163);
and U8316 (N_8316,N_7774,N_7391);
or U8317 (N_8317,N_6226,N_7338);
or U8318 (N_8318,N_7438,N_6378);
nand U8319 (N_8319,N_6618,N_7350);
nand U8320 (N_8320,N_7571,N_7237);
nand U8321 (N_8321,N_7909,N_6339);
or U8322 (N_8322,N_6494,N_6807);
nor U8323 (N_8323,N_6938,N_7957);
and U8324 (N_8324,N_7756,N_7423);
or U8325 (N_8325,N_7297,N_7641);
or U8326 (N_8326,N_6053,N_6580);
or U8327 (N_8327,N_7775,N_7315);
and U8328 (N_8328,N_6358,N_7766);
nor U8329 (N_8329,N_6981,N_7419);
or U8330 (N_8330,N_6725,N_7561);
nand U8331 (N_8331,N_7553,N_7009);
nor U8332 (N_8332,N_7143,N_6356);
and U8333 (N_8333,N_7006,N_7902);
and U8334 (N_8334,N_6406,N_6588);
and U8335 (N_8335,N_6033,N_7628);
nor U8336 (N_8336,N_7812,N_6201);
nand U8337 (N_8337,N_6254,N_7904);
and U8338 (N_8338,N_6379,N_6891);
or U8339 (N_8339,N_7430,N_6511);
nand U8340 (N_8340,N_7442,N_7569);
and U8341 (N_8341,N_7587,N_6516);
or U8342 (N_8342,N_6308,N_6348);
or U8343 (N_8343,N_6335,N_6052);
nand U8344 (N_8344,N_7886,N_7737);
nand U8345 (N_8345,N_7040,N_6476);
or U8346 (N_8346,N_7541,N_7007);
and U8347 (N_8347,N_7917,N_7908);
nand U8348 (N_8348,N_6952,N_6830);
xor U8349 (N_8349,N_6457,N_6365);
and U8350 (N_8350,N_7465,N_7458);
nor U8351 (N_8351,N_6546,N_6858);
or U8352 (N_8352,N_7753,N_6997);
nor U8353 (N_8353,N_6214,N_6554);
or U8354 (N_8354,N_6969,N_7461);
nand U8355 (N_8355,N_7895,N_6525);
nand U8356 (N_8356,N_6800,N_6401);
or U8357 (N_8357,N_7399,N_7915);
and U8358 (N_8358,N_6474,N_6655);
and U8359 (N_8359,N_7494,N_7213);
nor U8360 (N_8360,N_6253,N_7949);
and U8361 (N_8361,N_7931,N_6014);
nor U8362 (N_8362,N_6186,N_7152);
nor U8363 (N_8363,N_6983,N_6749);
nor U8364 (N_8364,N_7077,N_7476);
nand U8365 (N_8365,N_6433,N_7088);
nand U8366 (N_8366,N_7924,N_6314);
nor U8367 (N_8367,N_6528,N_7621);
or U8368 (N_8368,N_7705,N_6087);
and U8369 (N_8369,N_7402,N_6026);
and U8370 (N_8370,N_7033,N_7242);
or U8371 (N_8371,N_6815,N_7090);
and U8372 (N_8372,N_7994,N_6035);
and U8373 (N_8373,N_7462,N_6607);
nor U8374 (N_8374,N_7558,N_7129);
xor U8375 (N_8375,N_6345,N_7693);
nor U8376 (N_8376,N_6685,N_6683);
nand U8377 (N_8377,N_7792,N_7550);
nand U8378 (N_8378,N_7182,N_7151);
nand U8379 (N_8379,N_7971,N_6544);
or U8380 (N_8380,N_6295,N_7085);
and U8381 (N_8381,N_7439,N_6489);
nor U8382 (N_8382,N_7352,N_6402);
nor U8383 (N_8383,N_6276,N_7499);
and U8384 (N_8384,N_7803,N_6616);
or U8385 (N_8385,N_7795,N_6988);
nor U8386 (N_8386,N_7293,N_7845);
or U8387 (N_8387,N_6921,N_6881);
nor U8388 (N_8388,N_6404,N_7884);
and U8389 (N_8389,N_7221,N_6834);
and U8390 (N_8390,N_7910,N_7313);
and U8391 (N_8391,N_7874,N_6533);
nand U8392 (N_8392,N_7564,N_7586);
and U8393 (N_8393,N_6340,N_6225);
nor U8394 (N_8394,N_6583,N_6520);
nand U8395 (N_8395,N_7823,N_6462);
nand U8396 (N_8396,N_6286,N_6116);
nor U8397 (N_8397,N_6986,N_7801);
and U8398 (N_8398,N_7294,N_6510);
nand U8399 (N_8399,N_6529,N_7142);
and U8400 (N_8400,N_6168,N_6066);
and U8401 (N_8401,N_7609,N_7927);
and U8402 (N_8402,N_7235,N_6540);
and U8403 (N_8403,N_6568,N_7225);
and U8404 (N_8404,N_6319,N_7475);
nor U8405 (N_8405,N_7968,N_7723);
nand U8406 (N_8406,N_6144,N_6070);
nand U8407 (N_8407,N_7528,N_6202);
nor U8408 (N_8408,N_6198,N_6105);
or U8409 (N_8409,N_6490,N_7637);
and U8410 (N_8410,N_6421,N_6383);
or U8411 (N_8411,N_6387,N_7280);
nor U8412 (N_8412,N_7546,N_7665);
or U8413 (N_8413,N_7930,N_6793);
or U8414 (N_8414,N_6067,N_6946);
nand U8415 (N_8415,N_7544,N_7112);
nor U8416 (N_8416,N_7456,N_7218);
nor U8417 (N_8417,N_6512,N_7606);
and U8418 (N_8418,N_7119,N_6885);
nor U8419 (N_8419,N_6699,N_7473);
nand U8420 (N_8420,N_6362,N_7897);
and U8421 (N_8421,N_6941,N_6992);
and U8422 (N_8422,N_7929,N_6467);
nor U8423 (N_8423,N_6864,N_6117);
or U8424 (N_8424,N_6215,N_6692);
nand U8425 (N_8425,N_6990,N_7349);
nand U8426 (N_8426,N_6007,N_7505);
nand U8427 (N_8427,N_6846,N_6910);
or U8428 (N_8428,N_6248,N_7916);
xnor U8429 (N_8429,N_6656,N_6899);
nor U8430 (N_8430,N_7747,N_7694);
or U8431 (N_8431,N_6150,N_6288);
nand U8432 (N_8432,N_7328,N_7599);
nand U8433 (N_8433,N_6581,N_6898);
or U8434 (N_8434,N_6531,N_7173);
or U8435 (N_8435,N_7214,N_6208);
nor U8436 (N_8436,N_6232,N_7857);
and U8437 (N_8437,N_6537,N_7435);
and U8438 (N_8438,N_6003,N_6040);
and U8439 (N_8439,N_7947,N_7050);
nor U8440 (N_8440,N_7860,N_6897);
nand U8441 (N_8441,N_7028,N_6321);
or U8442 (N_8442,N_7245,N_7748);
nand U8443 (N_8443,N_7227,N_6821);
and U8444 (N_8444,N_7199,N_6382);
xnor U8445 (N_8445,N_6123,N_6437);
or U8446 (N_8446,N_7008,N_6274);
or U8447 (N_8447,N_7622,N_6923);
or U8448 (N_8448,N_6879,N_7556);
and U8449 (N_8449,N_7871,N_7390);
and U8450 (N_8450,N_6664,N_7138);
nor U8451 (N_8451,N_6417,N_6088);
or U8452 (N_8452,N_6621,N_7513);
xnor U8453 (N_8453,N_6714,N_6245);
and U8454 (N_8454,N_6968,N_6180);
or U8455 (N_8455,N_7420,N_7107);
nor U8456 (N_8456,N_6801,N_6316);
nand U8457 (N_8457,N_6980,N_6780);
or U8458 (N_8458,N_7719,N_6081);
or U8459 (N_8459,N_6671,N_7702);
nor U8460 (N_8460,N_7591,N_7646);
and U8461 (N_8461,N_7155,N_6883);
nand U8462 (N_8462,N_7384,N_7472);
nand U8463 (N_8463,N_7716,N_7371);
or U8464 (N_8464,N_7736,N_6287);
and U8465 (N_8465,N_7254,N_6374);
nor U8466 (N_8466,N_6464,N_7136);
or U8467 (N_8467,N_6844,N_7892);
and U8468 (N_8468,N_6904,N_6691);
nor U8469 (N_8469,N_7521,N_7859);
and U8470 (N_8470,N_6949,N_6219);
or U8471 (N_8471,N_6811,N_7312);
and U8472 (N_8472,N_7515,N_6359);
and U8473 (N_8473,N_7514,N_6470);
or U8474 (N_8474,N_7074,N_6107);
and U8475 (N_8475,N_7275,N_6259);
nor U8476 (N_8476,N_6715,N_7370);
and U8477 (N_8477,N_6163,N_6677);
nor U8478 (N_8478,N_6006,N_7623);
or U8479 (N_8479,N_7533,N_6207);
nor U8480 (N_8480,N_6483,N_6976);
or U8481 (N_8481,N_6928,N_7139);
and U8482 (N_8482,N_7117,N_7266);
nor U8483 (N_8483,N_7043,N_6538);
nor U8484 (N_8484,N_6023,N_7068);
and U8485 (N_8485,N_7278,N_7504);
nand U8486 (N_8486,N_6847,N_7650);
and U8487 (N_8487,N_6082,N_7849);
nor U8488 (N_8488,N_7447,N_6083);
or U8489 (N_8489,N_6032,N_6974);
or U8490 (N_8490,N_6391,N_6252);
nand U8491 (N_8491,N_7069,N_7019);
nor U8492 (N_8492,N_6019,N_6251);
and U8493 (N_8493,N_7306,N_7633);
and U8494 (N_8494,N_7634,N_6360);
or U8495 (N_8495,N_7345,N_6979);
and U8496 (N_8496,N_7635,N_7750);
and U8497 (N_8497,N_6493,N_7843);
nand U8498 (N_8498,N_6418,N_6001);
and U8499 (N_8499,N_7455,N_7938);
nor U8500 (N_8500,N_7333,N_6571);
nor U8501 (N_8501,N_7956,N_6808);
nor U8502 (N_8502,N_6759,N_7636);
and U8503 (N_8503,N_6709,N_7791);
nor U8504 (N_8504,N_7093,N_7366);
and U8505 (N_8505,N_6488,N_6130);
or U8506 (N_8506,N_6853,N_7835);
and U8507 (N_8507,N_6741,N_7096);
nor U8508 (N_8508,N_6000,N_6502);
nand U8509 (N_8509,N_6495,N_7039);
nor U8510 (N_8510,N_6466,N_7890);
nand U8511 (N_8511,N_6695,N_7557);
nand U8512 (N_8512,N_6028,N_6458);
and U8513 (N_8513,N_6361,N_7604);
and U8514 (N_8514,N_6303,N_7552);
nor U8515 (N_8515,N_7822,N_6636);
and U8516 (N_8516,N_7881,N_7379);
and U8517 (N_8517,N_7820,N_6854);
and U8518 (N_8518,N_7975,N_6506);
or U8519 (N_8519,N_6212,N_7819);
nor U8520 (N_8520,N_7358,N_7581);
nand U8521 (N_8521,N_7343,N_7876);
or U8522 (N_8522,N_6534,N_7726);
nor U8523 (N_8523,N_6649,N_7174);
nor U8524 (N_8524,N_6064,N_7217);
or U8525 (N_8525,N_6958,N_6519);
or U8526 (N_8526,N_7412,N_7122);
nand U8527 (N_8527,N_6757,N_6256);
or U8528 (N_8528,N_6115,N_6210);
nor U8529 (N_8529,N_7252,N_7014);
nor U8530 (N_8530,N_7652,N_6892);
nand U8531 (N_8531,N_7608,N_7335);
or U8532 (N_8532,N_6153,N_6735);
nand U8533 (N_8533,N_6389,N_7348);
nor U8534 (N_8534,N_6666,N_7785);
or U8535 (N_8535,N_6109,N_7317);
and U8536 (N_8536,N_6204,N_6625);
nand U8537 (N_8537,N_7285,N_7249);
or U8538 (N_8538,N_7522,N_7614);
or U8539 (N_8539,N_6722,N_7549);
and U8540 (N_8540,N_7405,N_7180);
nand U8541 (N_8541,N_7907,N_7648);
nand U8542 (N_8542,N_7322,N_7190);
or U8543 (N_8543,N_7751,N_7079);
or U8544 (N_8544,N_6833,N_6149);
nand U8545 (N_8545,N_7510,N_6973);
and U8546 (N_8546,N_7104,N_6189);
nor U8547 (N_8547,N_7543,N_6147);
and U8548 (N_8548,N_6243,N_6491);
nand U8549 (N_8549,N_6220,N_7066);
or U8550 (N_8550,N_7781,N_7565);
nand U8551 (N_8551,N_6816,N_7816);
and U8552 (N_8552,N_7758,N_6146);
nand U8553 (N_8553,N_6499,N_6721);
nor U8554 (N_8554,N_7655,N_6015);
nor U8555 (N_8555,N_6922,N_6475);
or U8556 (N_8556,N_6077,N_7865);
and U8557 (N_8557,N_7002,N_7684);
and U8558 (N_8558,N_6492,N_7156);
nor U8559 (N_8559,N_6178,N_7763);
nor U8560 (N_8560,N_7963,N_6536);
or U8561 (N_8561,N_6872,N_6138);
or U8562 (N_8562,N_6337,N_6679);
nand U8563 (N_8563,N_7003,N_6599);
nor U8564 (N_8564,N_6250,N_6249);
and U8565 (N_8565,N_6913,N_7817);
nor U8566 (N_8566,N_7205,N_6446);
and U8567 (N_8567,N_6063,N_7613);
nand U8568 (N_8568,N_6282,N_7660);
or U8569 (N_8569,N_7243,N_7932);
nor U8570 (N_8570,N_6895,N_7398);
or U8571 (N_8571,N_6688,N_6874);
xnor U8572 (N_8572,N_6963,N_6257);
nor U8573 (N_8573,N_7498,N_6235);
nor U8574 (N_8574,N_7424,N_7867);
or U8575 (N_8575,N_6547,N_6918);
nand U8576 (N_8576,N_7340,N_7773);
nor U8577 (N_8577,N_7134,N_6765);
and U8578 (N_8578,N_7905,N_7471);
and U8579 (N_8579,N_6310,N_6447);
and U8580 (N_8580,N_6409,N_6086);
nand U8581 (N_8581,N_6609,N_6681);
and U8582 (N_8582,N_7200,N_7687);
nand U8583 (N_8583,N_7234,N_6654);
and U8584 (N_8584,N_6338,N_6472);
and U8585 (N_8585,N_7224,N_7086);
nor U8586 (N_8586,N_6200,N_7084);
or U8587 (N_8587,N_6877,N_7001);
nor U8588 (N_8588,N_7226,N_7457);
and U8589 (N_8589,N_7042,N_6553);
nor U8590 (N_8590,N_7862,N_6615);
or U8591 (N_8591,N_7811,N_7196);
nand U8592 (N_8592,N_7038,N_6622);
and U8593 (N_8593,N_6234,N_7146);
and U8594 (N_8594,N_6640,N_6237);
nand U8595 (N_8595,N_7075,N_7809);
or U8596 (N_8596,N_6975,N_7208);
and U8597 (N_8597,N_6038,N_6124);
or U8598 (N_8598,N_7314,N_6530);
and U8599 (N_8599,N_7673,N_6848);
nor U8600 (N_8600,N_6919,N_6054);
or U8601 (N_8601,N_6280,N_7351);
xnor U8602 (N_8602,N_7320,N_6487);
nand U8603 (N_8603,N_7482,N_6845);
and U8604 (N_8604,N_6423,N_7206);
or U8605 (N_8605,N_6341,N_6353);
nor U8606 (N_8606,N_7523,N_7631);
nor U8607 (N_8607,N_6577,N_7760);
nor U8608 (N_8608,N_7354,N_7717);
nand U8609 (N_8609,N_6785,N_7177);
nand U8610 (N_8610,N_6002,N_6720);
nand U8611 (N_8611,N_6717,N_7228);
or U8612 (N_8612,N_7657,N_6729);
and U8613 (N_8613,N_6894,N_7045);
nor U8614 (N_8614,N_7072,N_6805);
and U8615 (N_8615,N_6371,N_6399);
nor U8616 (N_8616,N_7211,N_7308);
or U8617 (N_8617,N_6587,N_7426);
and U8618 (N_8618,N_7128,N_6501);
nand U8619 (N_8619,N_7202,N_6127);
or U8620 (N_8620,N_6719,N_7073);
nand U8621 (N_8621,N_7288,N_6145);
nand U8622 (N_8622,N_6111,N_7962);
and U8623 (N_8623,N_7810,N_7977);
or U8624 (N_8624,N_7013,N_6394);
nand U8625 (N_8625,N_7987,N_6905);
and U8626 (N_8626,N_7518,N_6931);
nor U8627 (N_8627,N_6333,N_7624);
nor U8628 (N_8628,N_7630,N_6718);
and U8629 (N_8629,N_6174,N_6194);
nor U8630 (N_8630,N_6750,N_7178);
or U8631 (N_8631,N_7846,N_7440);
and U8632 (N_8632,N_6646,N_7126);
nand U8633 (N_8633,N_6789,N_6390);
or U8634 (N_8634,N_6324,N_7157);
or U8635 (N_8635,N_7844,N_7536);
and U8636 (N_8636,N_6782,N_6030);
nand U8637 (N_8637,N_6293,N_7158);
nand U8638 (N_8638,N_6233,N_6602);
nand U8639 (N_8639,N_7663,N_6485);
nor U8640 (N_8640,N_6171,N_7961);
nor U8641 (N_8641,N_7464,N_6222);
nor U8642 (N_8642,N_7700,N_7853);
nor U8643 (N_8643,N_6550,N_6866);
nor U8644 (N_8644,N_7779,N_6170);
nor U8645 (N_8645,N_7952,N_6971);
nor U8646 (N_8646,N_7295,N_7743);
or U8647 (N_8647,N_6527,N_6564);
nor U8648 (N_8648,N_6878,N_7632);
nor U8649 (N_8649,N_6940,N_7605);
or U8650 (N_8650,N_7114,N_7361);
or U8651 (N_8651,N_7559,N_6412);
or U8652 (N_8652,N_6809,N_6046);
nor U8653 (N_8653,N_7659,N_6156);
nor U8654 (N_8654,N_6935,N_7374);
or U8655 (N_8655,N_7669,N_6961);
nand U8656 (N_8656,N_7683,N_6024);
nor U8657 (N_8657,N_7629,N_6095);
nor U8658 (N_8658,N_7517,N_7031);
nor U8659 (N_8659,N_6998,N_7863);
and U8660 (N_8660,N_6770,N_6838);
or U8661 (N_8661,N_7981,N_7925);
nand U8662 (N_8662,N_6327,N_7725);
nand U8663 (N_8663,N_7463,N_6631);
and U8664 (N_8664,N_6098,N_6020);
nor U8665 (N_8665,N_6076,N_6651);
and U8666 (N_8666,N_7731,N_6247);
and U8667 (N_8667,N_6948,N_6850);
nor U8668 (N_8668,N_7044,N_7699);
or U8669 (N_8669,N_7048,N_7262);
and U8670 (N_8670,N_6570,N_6687);
or U8671 (N_8671,N_6018,N_7283);
nor U8672 (N_8672,N_7316,N_7449);
nor U8673 (N_8673,N_7718,N_7382);
and U8674 (N_8674,N_6263,N_6890);
or U8675 (N_8675,N_7427,N_6804);
nand U8676 (N_8676,N_6062,N_7035);
nand U8677 (N_8677,N_7959,N_7393);
nor U8678 (N_8678,N_6517,N_7834);
xnor U8679 (N_8679,N_6336,N_7185);
nand U8680 (N_8680,N_7417,N_7359);
nand U8681 (N_8681,N_6943,N_7244);
or U8682 (N_8682,N_7800,N_6322);
nand U8683 (N_8683,N_7496,N_6624);
nor U8684 (N_8684,N_7562,N_7567);
nand U8685 (N_8685,N_7403,N_6332);
nand U8686 (N_8686,N_6959,N_6914);
and U8687 (N_8687,N_7305,N_6751);
nor U8688 (N_8688,N_6925,N_7797);
or U8689 (N_8689,N_6125,N_6203);
and U8690 (N_8690,N_6977,N_6798);
and U8691 (N_8691,N_7563,N_7025);
nor U8692 (N_8692,N_6951,N_7730);
nor U8693 (N_8693,N_7856,N_7508);
and U8694 (N_8694,N_6806,N_7912);
and U8695 (N_8695,N_6873,N_7184);
nand U8696 (N_8696,N_7566,N_6831);
or U8697 (N_8697,N_6160,N_7034);
or U8698 (N_8698,N_6708,N_6448);
nor U8699 (N_8699,N_6747,N_7500);
nor U8700 (N_8700,N_6855,N_6230);
nand U8701 (N_8701,N_7487,N_6384);
and U8702 (N_8702,N_7627,N_7489);
nand U8703 (N_8703,N_7330,N_6471);
or U8704 (N_8704,N_7708,N_7933);
and U8705 (N_8705,N_6436,N_7955);
or U8706 (N_8706,N_6148,N_7261);
or U8707 (N_8707,N_6573,N_6987);
or U8708 (N_8708,N_6407,N_7826);
and U8709 (N_8709,N_7701,N_6755);
xnor U8710 (N_8710,N_6021,N_7167);
nand U8711 (N_8711,N_7454,N_6557);
nor U8712 (N_8712,N_6434,N_6344);
and U8713 (N_8713,N_7289,N_6408);
nand U8714 (N_8714,N_7724,N_7397);
nor U8715 (N_8715,N_6484,N_6155);
and U8716 (N_8716,N_6106,N_7534);
or U8717 (N_8717,N_7347,N_6400);
nor U8718 (N_8718,N_6927,N_6128);
and U8719 (N_8719,N_6767,N_6444);
nand U8720 (N_8720,N_7054,N_7133);
nand U8721 (N_8721,N_6758,N_7344);
and U8722 (N_8722,N_7877,N_7978);
nand U8723 (N_8723,N_6008,N_6429);
or U8724 (N_8724,N_7749,N_6701);
and U8725 (N_8725,N_6426,N_6802);
and U8726 (N_8726,N_7617,N_6104);
or U8727 (N_8727,N_7789,N_7111);
nand U8728 (N_8728,N_6497,N_7524);
or U8729 (N_8729,N_7466,N_6598);
nor U8730 (N_8730,N_7239,N_6143);
nor U8731 (N_8731,N_6724,N_6084);
nor U8732 (N_8732,N_6995,N_6079);
and U8733 (N_8733,N_6058,N_7548);
nand U8734 (N_8734,N_7411,N_7160);
or U8735 (N_8735,N_7273,N_7443);
nor U8736 (N_8736,N_7078,N_6388);
and U8737 (N_8737,N_6438,N_6779);
or U8738 (N_8738,N_7253,N_6690);
nand U8739 (N_8739,N_6710,N_6505);
nor U8740 (N_8740,N_6051,N_6608);
nor U8741 (N_8741,N_7883,N_7091);
nor U8742 (N_8742,N_6224,N_6381);
nand U8743 (N_8743,N_6628,N_7113);
nand U8744 (N_8744,N_7982,N_6352);
or U8745 (N_8745,N_6545,N_7979);
nand U8746 (N_8746,N_7483,N_7511);
and U8747 (N_8747,N_6863,N_7386);
nor U8748 (N_8748,N_6796,N_7241);
or U8749 (N_8749,N_6822,N_6238);
or U8750 (N_8750,N_6612,N_6036);
nand U8751 (N_8751,N_6460,N_7223);
nand U8752 (N_8752,N_6480,N_7670);
or U8753 (N_8753,N_7772,N_7251);
or U8754 (N_8754,N_7804,N_7872);
and U8755 (N_8755,N_7729,N_7263);
nor U8756 (N_8756,N_6728,N_6596);
or U8757 (N_8757,N_6477,N_7413);
or U8758 (N_8758,N_7389,N_6217);
and U8759 (N_8759,N_7017,N_7574);
nand U8760 (N_8760,N_6578,N_6562);
or U8761 (N_8761,N_7594,N_6080);
xnor U8762 (N_8762,N_7355,N_7191);
or U8763 (N_8763,N_6752,N_6069);
or U8764 (N_8764,N_7974,N_6211);
or U8765 (N_8765,N_7850,N_7784);
and U8766 (N_8766,N_6911,N_7148);
or U8767 (N_8767,N_7615,N_6888);
or U8768 (N_8768,N_6101,N_7353);
nor U8769 (N_8769,N_7593,N_6029);
nor U8770 (N_8770,N_7828,N_7882);
and U8771 (N_8771,N_7990,N_7302);
nor U8772 (N_8772,N_7814,N_7356);
or U8773 (N_8773,N_7799,N_6177);
nor U8774 (N_8774,N_6908,N_7183);
and U8775 (N_8775,N_7936,N_6698);
nor U8776 (N_8776,N_7240,N_6231);
or U8777 (N_8777,N_7696,N_7768);
nand U8778 (N_8778,N_6982,N_6610);
nor U8779 (N_8779,N_7551,N_6165);
nand U8780 (N_8780,N_6781,N_7258);
nand U8781 (N_8781,N_7394,N_7592);
nor U8782 (N_8782,N_6574,N_6733);
and U8783 (N_8783,N_7953,N_6678);
nand U8784 (N_8784,N_7639,N_7671);
nand U8785 (N_8785,N_7855,N_6648);
and U8786 (N_8786,N_6582,N_6442);
and U8787 (N_8787,N_7020,N_6373);
and U8788 (N_8788,N_7131,N_7323);
and U8789 (N_8789,N_7303,N_6289);
nor U8790 (N_8790,N_6865,N_7603);
nand U8791 (N_8791,N_6569,N_6929);
and U8792 (N_8792,N_6140,N_6463);
nand U8793 (N_8793,N_7922,N_6944);
nand U8794 (N_8794,N_7296,N_7168);
and U8795 (N_8795,N_6558,N_7291);
or U8796 (N_8796,N_6187,N_7827);
and U8797 (N_8797,N_6122,N_7059);
and U8798 (N_8798,N_7395,N_6778);
and U8799 (N_8799,N_7806,N_6661);
nand U8800 (N_8800,N_6410,N_7478);
and U8801 (N_8801,N_7525,N_7170);
nor U8802 (N_8802,N_7888,N_7329);
nor U8803 (N_8803,N_7727,N_7951);
or U8804 (N_8804,N_6134,N_6956);
and U8805 (N_8805,N_6413,N_6092);
nor U8806 (N_8806,N_6416,N_7576);
and U8807 (N_8807,N_6670,N_6662);
and U8808 (N_8808,N_6642,N_6268);
and U8809 (N_8809,N_6403,N_6705);
nor U8810 (N_8810,N_6920,N_7689);
or U8811 (N_8811,N_6777,N_6859);
or U8812 (N_8812,N_6131,N_7369);
nor U8813 (N_8813,N_6240,N_7304);
or U8814 (N_8814,N_7446,N_7255);
nand U8815 (N_8815,N_7470,N_7969);
nand U8816 (N_8816,N_6933,N_7770);
xnor U8817 (N_8817,N_6045,N_6016);
or U8818 (N_8818,N_7246,N_7829);
nand U8819 (N_8819,N_6167,N_6880);
or U8820 (N_8820,N_7607,N_7643);
nor U8821 (N_8821,N_7948,N_6221);
nand U8822 (N_8822,N_6893,N_7771);
nand U8823 (N_8823,N_7989,N_7965);
or U8824 (N_8824,N_6405,N_6151);
or U8825 (N_8825,N_6368,N_6162);
nor U8826 (N_8826,N_7741,N_6445);
nor U8827 (N_8827,N_7570,N_7490);
or U8828 (N_8828,N_7752,N_6120);
nor U8829 (N_8829,N_7538,N_6623);
or U8830 (N_8830,N_6643,N_7232);
or U8831 (N_8831,N_6542,N_7764);
and U8832 (N_8832,N_6179,N_7216);
or U8833 (N_8833,N_7512,N_7065);
nand U8834 (N_8834,N_6541,N_6395);
or U8835 (N_8835,N_7108,N_7680);
or U8836 (N_8836,N_6875,N_7318);
and U8837 (N_8837,N_6469,N_6367);
nand U8838 (N_8838,N_6461,N_7172);
nand U8839 (N_8839,N_6706,N_6182);
and U8840 (N_8840,N_6135,N_6206);
nor U8841 (N_8841,N_6025,N_6056);
nand U8842 (N_8842,N_6824,N_7298);
or U8843 (N_8843,N_6559,N_6279);
nor U8844 (N_8844,N_6744,N_7906);
nand U8845 (N_8845,N_6427,N_7590);
and U8846 (N_8846,N_7690,N_6290);
and U8847 (N_8847,N_7654,N_7036);
or U8848 (N_8848,N_7012,N_7149);
nand U8849 (N_8849,N_7236,N_7015);
or U8850 (N_8850,N_7450,N_6205);
nor U8851 (N_8851,N_7858,N_6398);
and U8852 (N_8852,N_7124,N_7878);
nor U8853 (N_8853,N_7901,N_7651);
xor U8854 (N_8854,N_6667,N_7175);
and U8855 (N_8855,N_6228,N_6191);
nor U8856 (N_8856,N_7620,N_7695);
nor U8857 (N_8857,N_6955,N_6842);
or U8858 (N_8858,N_7519,N_7560);
nand U8859 (N_8859,N_6113,N_7722);
and U8860 (N_8860,N_7194,N_7821);
nor U8861 (N_8861,N_7176,N_7198);
or U8862 (N_8862,N_6270,N_7808);
or U8863 (N_8863,N_6175,N_6424);
or U8864 (N_8864,N_7460,N_7537);
and U8865 (N_8865,N_6909,N_7105);
nand U8866 (N_8866,N_6272,N_6861);
or U8867 (N_8867,N_6227,N_7368);
or U8868 (N_8868,N_6614,N_6068);
nand U8869 (N_8869,N_7064,N_7195);
nand U8870 (N_8870,N_6091,N_6639);
nor U8871 (N_8871,N_7272,N_7666);
nand U8872 (N_8872,N_7229,N_7585);
nor U8873 (N_8873,N_6330,N_7745);
nor U8874 (N_8874,N_6285,N_6797);
nand U8875 (N_8875,N_7658,N_6261);
or U8876 (N_8876,N_6422,N_7815);
nand U8877 (N_8877,N_7941,N_6548);
and U8878 (N_8878,N_7780,N_7626);
nand U8879 (N_8879,N_7437,N_7676);
nand U8880 (N_8880,N_7575,N_6836);
nand U8881 (N_8881,N_6196,N_7492);
nor U8882 (N_8882,N_6141,N_6543);
and U8883 (N_8883,N_6707,N_6244);
nand U8884 (N_8884,N_6584,N_7507);
nand U8885 (N_8885,N_7055,N_7011);
nor U8886 (N_8886,N_7010,N_7484);
nor U8887 (N_8887,N_7582,N_6468);
nand U8888 (N_8888,N_7616,N_6185);
or U8889 (N_8889,N_6139,N_6267);
nand U8890 (N_8890,N_6443,N_7453);
and U8891 (N_8891,N_7928,N_6849);
and U8892 (N_8892,N_7319,N_7429);
nor U8893 (N_8893,N_6682,N_7649);
and U8894 (N_8894,N_7520,N_7873);
or U8895 (N_8895,N_7681,N_6049);
and U8896 (N_8896,N_7703,N_6748);
and U8897 (N_8897,N_7778,N_6159);
nor U8898 (N_8898,N_6957,N_7530);
nand U8899 (N_8899,N_7547,N_7911);
or U8900 (N_8900,N_6810,N_6273);
or U8901 (N_8901,N_7342,N_7964);
nor U8902 (N_8902,N_7691,N_6650);
nand U8903 (N_8903,N_7164,N_7037);
nor U8904 (N_8904,N_7662,N_6291);
and U8905 (N_8905,N_7414,N_6057);
or U8906 (N_8906,N_6055,N_7937);
and U8907 (N_8907,N_7950,N_6962);
or U8908 (N_8908,N_7831,N_7710);
or U8909 (N_8909,N_6783,N_7923);
nor U8910 (N_8910,N_7854,N_6498);
nand U8911 (N_8911,N_7600,N_6889);
nor U8912 (N_8912,N_7762,N_7596);
or U8913 (N_8913,N_6262,N_6275);
or U8914 (N_8914,N_7682,N_6630);
and U8915 (N_8915,N_7577,N_7145);
or U8916 (N_8916,N_7998,N_7372);
and U8917 (N_8917,N_6059,N_6936);
or U8918 (N_8918,N_7094,N_6964);
nand U8919 (N_8919,N_7267,N_7270);
nand U8920 (N_8920,N_7588,N_7868);
nor U8921 (N_8921,N_6044,N_7675);
or U8922 (N_8922,N_6672,N_6693);
or U8923 (N_8923,N_6508,N_7506);
nand U8924 (N_8924,N_7985,N_7889);
and U8925 (N_8925,N_6900,N_6432);
nand U8926 (N_8926,N_6479,N_7383);
or U8927 (N_8927,N_6647,N_6133);
nand U8928 (N_8928,N_7842,N_7049);
or U8929 (N_8929,N_7377,N_6043);
nor U8930 (N_8930,N_6552,N_6901);
or U8931 (N_8931,N_7712,N_7993);
and U8932 (N_8932,N_7248,N_7210);
nor U8933 (N_8933,N_7796,N_6775);
nor U8934 (N_8934,N_6523,N_7813);
and U8935 (N_8935,N_6790,N_7101);
or U8936 (N_8936,N_6737,N_7193);
or U8937 (N_8937,N_6377,N_6397);
or U8938 (N_8938,N_6860,N_7381);
nor U8939 (N_8939,N_7123,N_7127);
nor U8940 (N_8940,N_6756,N_6093);
or U8941 (N_8941,N_6660,N_7257);
nand U8942 (N_8942,N_7900,N_7798);
nand U8943 (N_8943,N_6906,N_6363);
nor U8944 (N_8944,N_6676,N_7946);
and U8945 (N_8945,N_6740,N_7776);
nor U8946 (N_8946,N_6169,N_6154);
or U8947 (N_8947,N_6993,N_6606);
or U8948 (N_8948,N_7259,N_7147);
or U8949 (N_8949,N_6814,N_6166);
and U8950 (N_8950,N_6334,N_6738);
or U8951 (N_8951,N_6917,N_6349);
nand U8952 (N_8952,N_6652,N_7376);
nand U8953 (N_8953,N_6947,N_6100);
nand U8954 (N_8954,N_6791,N_6031);
and U8955 (N_8955,N_6696,N_7943);
and U8956 (N_8956,N_6886,N_7913);
nor U8957 (N_8957,N_6017,N_7866);
nor U8958 (N_8958,N_7509,N_7144);
nor U8959 (N_8959,N_7495,N_7861);
nor U8960 (N_8960,N_6932,N_6567);
nor U8961 (N_8961,N_7321,N_7047);
and U8962 (N_8962,N_7018,N_7757);
and U8963 (N_8963,N_7674,N_6478);
nor U8964 (N_8964,N_7326,N_7765);
nor U8965 (N_8965,N_6414,N_6005);
nor U8966 (N_8966,N_6857,N_6984);
or U8967 (N_8967,N_6592,N_6507);
or U8968 (N_8968,N_7380,N_6619);
nand U8969 (N_8969,N_6103,N_7836);
and U8970 (N_8970,N_7051,N_7057);
or U8971 (N_8971,N_7474,N_7704);
nand U8972 (N_8972,N_7098,N_6119);
nand U8973 (N_8973,N_7479,N_7418);
or U8974 (N_8974,N_7197,N_7219);
or U8975 (N_8975,N_6829,N_6236);
or U8976 (N_8976,N_7404,N_6716);
or U8977 (N_8977,N_7894,N_6320);
and U8978 (N_8978,N_6764,N_7503);
and U8979 (N_8979,N_6726,N_6312);
nand U8980 (N_8980,N_6994,N_7914);
or U8981 (N_8981,N_6325,N_6734);
and U8982 (N_8982,N_6551,N_7903);
nor U8983 (N_8983,N_6304,N_6509);
nor U8984 (N_8984,N_6355,N_6090);
and U8985 (N_8985,N_6832,N_6022);
and U8986 (N_8986,N_7692,N_7818);
nor U8987 (N_8987,N_6513,N_6158);
or U8988 (N_8988,N_7301,N_6075);
nor U8989 (N_8989,N_6585,N_6229);
and U8990 (N_8990,N_6556,N_7920);
nor U8991 (N_8991,N_7777,N_6011);
or U8992 (N_8992,N_6868,N_7880);
and U8993 (N_8993,N_6907,N_7754);
and U8994 (N_8994,N_6500,N_6048);
and U8995 (N_8995,N_6299,N_7264);
or U8996 (N_8996,N_7269,N_7233);
nand U8997 (N_8997,N_7545,N_7118);
nor U8998 (N_8998,N_6521,N_7618);
and U8999 (N_8999,N_6953,N_6743);
or U9000 (N_9000,N_7505,N_7062);
or U9001 (N_9001,N_6268,N_6511);
and U9002 (N_9002,N_6280,N_6392);
xor U9003 (N_9003,N_6507,N_6148);
or U9004 (N_9004,N_7741,N_6012);
nor U9005 (N_9005,N_7210,N_7045);
nor U9006 (N_9006,N_7449,N_7905);
and U9007 (N_9007,N_6989,N_7461);
nand U9008 (N_9008,N_6434,N_6269);
nand U9009 (N_9009,N_6571,N_6264);
nor U9010 (N_9010,N_6152,N_6608);
and U9011 (N_9011,N_6718,N_6386);
nor U9012 (N_9012,N_6017,N_7625);
nor U9013 (N_9013,N_7555,N_6460);
or U9014 (N_9014,N_6763,N_7238);
or U9015 (N_9015,N_7794,N_7972);
or U9016 (N_9016,N_7711,N_6003);
or U9017 (N_9017,N_6008,N_6423);
nand U9018 (N_9018,N_6804,N_6815);
and U9019 (N_9019,N_7385,N_6009);
nor U9020 (N_9020,N_7835,N_6347);
nand U9021 (N_9021,N_6815,N_6393);
nand U9022 (N_9022,N_7159,N_6854);
and U9023 (N_9023,N_6306,N_6265);
nor U9024 (N_9024,N_6615,N_6674);
nor U9025 (N_9025,N_6156,N_6452);
nand U9026 (N_9026,N_6078,N_7261);
nand U9027 (N_9027,N_6545,N_6587);
nand U9028 (N_9028,N_7844,N_6502);
nand U9029 (N_9029,N_6273,N_7728);
or U9030 (N_9030,N_6691,N_7211);
or U9031 (N_9031,N_6028,N_7350);
nor U9032 (N_9032,N_6225,N_6457);
nand U9033 (N_9033,N_7273,N_6707);
nor U9034 (N_9034,N_7161,N_7821);
or U9035 (N_9035,N_6530,N_6138);
or U9036 (N_9036,N_6649,N_7027);
nor U9037 (N_9037,N_7592,N_7120);
nor U9038 (N_9038,N_6931,N_7621);
or U9039 (N_9039,N_7285,N_6037);
nand U9040 (N_9040,N_6837,N_7842);
or U9041 (N_9041,N_7359,N_6314);
and U9042 (N_9042,N_6528,N_6110);
or U9043 (N_9043,N_7795,N_7366);
nand U9044 (N_9044,N_6540,N_6139);
or U9045 (N_9045,N_6583,N_6059);
nand U9046 (N_9046,N_7133,N_7353);
nand U9047 (N_9047,N_7378,N_6354);
and U9048 (N_9048,N_7623,N_6010);
or U9049 (N_9049,N_6498,N_7375);
or U9050 (N_9050,N_7952,N_7528);
nor U9051 (N_9051,N_7165,N_7838);
nor U9052 (N_9052,N_7447,N_6818);
nand U9053 (N_9053,N_7683,N_7660);
nor U9054 (N_9054,N_7351,N_6644);
or U9055 (N_9055,N_7286,N_6253);
and U9056 (N_9056,N_6476,N_7742);
nor U9057 (N_9057,N_6500,N_6228);
and U9058 (N_9058,N_7622,N_6717);
and U9059 (N_9059,N_6663,N_6399);
nand U9060 (N_9060,N_7152,N_7576);
nand U9061 (N_9061,N_6642,N_6572);
nor U9062 (N_9062,N_7046,N_6840);
or U9063 (N_9063,N_7886,N_6874);
nand U9064 (N_9064,N_7587,N_7954);
nand U9065 (N_9065,N_7066,N_7738);
nor U9066 (N_9066,N_7576,N_7930);
nor U9067 (N_9067,N_7678,N_7309);
or U9068 (N_9068,N_6823,N_7477);
nor U9069 (N_9069,N_6679,N_6563);
and U9070 (N_9070,N_7145,N_6031);
nor U9071 (N_9071,N_7028,N_7128);
and U9072 (N_9072,N_7980,N_7697);
nor U9073 (N_9073,N_6558,N_6551);
or U9074 (N_9074,N_6766,N_6969);
and U9075 (N_9075,N_7108,N_7916);
nand U9076 (N_9076,N_7823,N_7730);
nor U9077 (N_9077,N_6481,N_7329);
or U9078 (N_9078,N_6351,N_6638);
nor U9079 (N_9079,N_7093,N_7162);
nand U9080 (N_9080,N_7278,N_6013);
nand U9081 (N_9081,N_6095,N_7973);
nor U9082 (N_9082,N_6792,N_6485);
nand U9083 (N_9083,N_7400,N_6477);
nor U9084 (N_9084,N_7295,N_6853);
and U9085 (N_9085,N_6625,N_6598);
or U9086 (N_9086,N_7174,N_6393);
or U9087 (N_9087,N_6672,N_6778);
and U9088 (N_9088,N_7466,N_7318);
xor U9089 (N_9089,N_6925,N_6911);
or U9090 (N_9090,N_7295,N_6393);
nor U9091 (N_9091,N_7217,N_6845);
and U9092 (N_9092,N_7977,N_7344);
nor U9093 (N_9093,N_7157,N_7563);
and U9094 (N_9094,N_6081,N_7793);
and U9095 (N_9095,N_6244,N_6902);
nor U9096 (N_9096,N_6338,N_7806);
nand U9097 (N_9097,N_6138,N_6280);
and U9098 (N_9098,N_7783,N_7709);
nand U9099 (N_9099,N_6787,N_6665);
or U9100 (N_9100,N_6066,N_7735);
or U9101 (N_9101,N_6553,N_6398);
or U9102 (N_9102,N_6443,N_7526);
or U9103 (N_9103,N_6932,N_7190);
nand U9104 (N_9104,N_6614,N_6399);
or U9105 (N_9105,N_6992,N_6721);
and U9106 (N_9106,N_6285,N_7337);
and U9107 (N_9107,N_7087,N_6592);
nand U9108 (N_9108,N_6838,N_7849);
or U9109 (N_9109,N_7535,N_7647);
nand U9110 (N_9110,N_7412,N_7503);
and U9111 (N_9111,N_7217,N_7674);
and U9112 (N_9112,N_6890,N_6873);
or U9113 (N_9113,N_7155,N_7234);
nand U9114 (N_9114,N_7158,N_6064);
nor U9115 (N_9115,N_7413,N_7922);
nor U9116 (N_9116,N_6799,N_6615);
and U9117 (N_9117,N_6024,N_6226);
or U9118 (N_9118,N_6693,N_6204);
or U9119 (N_9119,N_6601,N_7800);
nor U9120 (N_9120,N_6019,N_6046);
and U9121 (N_9121,N_7890,N_6661);
or U9122 (N_9122,N_6645,N_7978);
and U9123 (N_9123,N_6503,N_7361);
and U9124 (N_9124,N_6202,N_7068);
nand U9125 (N_9125,N_6183,N_7560);
and U9126 (N_9126,N_7565,N_7727);
and U9127 (N_9127,N_6379,N_7377);
and U9128 (N_9128,N_6711,N_7258);
nor U9129 (N_9129,N_6681,N_7565);
or U9130 (N_9130,N_6854,N_7181);
nor U9131 (N_9131,N_7000,N_6926);
nor U9132 (N_9132,N_7978,N_6153);
nor U9133 (N_9133,N_6702,N_7358);
and U9134 (N_9134,N_6975,N_7294);
nor U9135 (N_9135,N_6018,N_7876);
nand U9136 (N_9136,N_7168,N_6254);
nor U9137 (N_9137,N_7764,N_7424);
and U9138 (N_9138,N_7974,N_7970);
and U9139 (N_9139,N_7057,N_7917);
nand U9140 (N_9140,N_7167,N_7827);
nand U9141 (N_9141,N_6719,N_7701);
and U9142 (N_9142,N_6087,N_7393);
nand U9143 (N_9143,N_7418,N_6285);
nor U9144 (N_9144,N_6064,N_6213);
or U9145 (N_9145,N_7202,N_7174);
or U9146 (N_9146,N_6092,N_7441);
or U9147 (N_9147,N_7042,N_6831);
and U9148 (N_9148,N_6790,N_6736);
or U9149 (N_9149,N_7097,N_6591);
and U9150 (N_9150,N_6594,N_6485);
nand U9151 (N_9151,N_7421,N_7476);
and U9152 (N_9152,N_7542,N_7425);
nor U9153 (N_9153,N_7429,N_7946);
nand U9154 (N_9154,N_6490,N_6818);
and U9155 (N_9155,N_6556,N_6659);
nor U9156 (N_9156,N_7780,N_6019);
nor U9157 (N_9157,N_7971,N_6840);
nor U9158 (N_9158,N_6969,N_7208);
nor U9159 (N_9159,N_7914,N_7694);
nor U9160 (N_9160,N_7668,N_6102);
and U9161 (N_9161,N_6107,N_6298);
nor U9162 (N_9162,N_6930,N_6419);
and U9163 (N_9163,N_7784,N_6123);
nand U9164 (N_9164,N_7744,N_7281);
nand U9165 (N_9165,N_6379,N_7894);
nor U9166 (N_9166,N_7894,N_7756);
and U9167 (N_9167,N_6351,N_6034);
nor U9168 (N_9168,N_6217,N_7607);
nor U9169 (N_9169,N_7653,N_7427);
nor U9170 (N_9170,N_6478,N_7277);
nor U9171 (N_9171,N_6142,N_6344);
nand U9172 (N_9172,N_7703,N_6939);
nor U9173 (N_9173,N_6871,N_7179);
or U9174 (N_9174,N_7502,N_7157);
nand U9175 (N_9175,N_6182,N_7880);
and U9176 (N_9176,N_6780,N_6059);
or U9177 (N_9177,N_6136,N_6804);
nor U9178 (N_9178,N_6914,N_7601);
nor U9179 (N_9179,N_6581,N_7395);
and U9180 (N_9180,N_6897,N_7263);
or U9181 (N_9181,N_6596,N_7836);
nand U9182 (N_9182,N_7073,N_7452);
nand U9183 (N_9183,N_6107,N_7724);
nand U9184 (N_9184,N_7074,N_7592);
and U9185 (N_9185,N_6038,N_7043);
and U9186 (N_9186,N_6109,N_6824);
nand U9187 (N_9187,N_7242,N_6194);
and U9188 (N_9188,N_7838,N_7151);
and U9189 (N_9189,N_6002,N_6108);
or U9190 (N_9190,N_7114,N_7185);
nand U9191 (N_9191,N_6154,N_7870);
and U9192 (N_9192,N_7996,N_7103);
or U9193 (N_9193,N_6513,N_6172);
or U9194 (N_9194,N_6611,N_6187);
and U9195 (N_9195,N_6957,N_7487);
or U9196 (N_9196,N_6844,N_6289);
or U9197 (N_9197,N_7657,N_7339);
and U9198 (N_9198,N_6125,N_6785);
nand U9199 (N_9199,N_6676,N_7377);
nor U9200 (N_9200,N_7561,N_6853);
and U9201 (N_9201,N_6769,N_7566);
or U9202 (N_9202,N_7474,N_6668);
nor U9203 (N_9203,N_7054,N_7872);
or U9204 (N_9204,N_6510,N_6491);
and U9205 (N_9205,N_6309,N_6371);
and U9206 (N_9206,N_7509,N_6671);
or U9207 (N_9207,N_6710,N_7834);
nand U9208 (N_9208,N_7089,N_6094);
nor U9209 (N_9209,N_6260,N_6738);
and U9210 (N_9210,N_7733,N_6983);
nand U9211 (N_9211,N_7417,N_6635);
and U9212 (N_9212,N_7720,N_6858);
nand U9213 (N_9213,N_7626,N_7862);
nand U9214 (N_9214,N_7769,N_6087);
nand U9215 (N_9215,N_6039,N_6526);
or U9216 (N_9216,N_6343,N_6619);
nand U9217 (N_9217,N_7856,N_6880);
nand U9218 (N_9218,N_7485,N_7483);
nor U9219 (N_9219,N_7942,N_6364);
nand U9220 (N_9220,N_7007,N_7699);
nor U9221 (N_9221,N_7384,N_6700);
and U9222 (N_9222,N_6091,N_6521);
nand U9223 (N_9223,N_6644,N_6280);
or U9224 (N_9224,N_7192,N_7222);
nor U9225 (N_9225,N_7496,N_7484);
and U9226 (N_9226,N_7151,N_7225);
nand U9227 (N_9227,N_6785,N_6291);
nand U9228 (N_9228,N_7946,N_7498);
nor U9229 (N_9229,N_6155,N_7739);
and U9230 (N_9230,N_6548,N_7999);
nor U9231 (N_9231,N_7899,N_6511);
or U9232 (N_9232,N_7083,N_6177);
nor U9233 (N_9233,N_7944,N_7866);
nand U9234 (N_9234,N_7792,N_7500);
nor U9235 (N_9235,N_7830,N_6427);
nor U9236 (N_9236,N_6563,N_7077);
nand U9237 (N_9237,N_6551,N_6651);
nand U9238 (N_9238,N_6345,N_7457);
nor U9239 (N_9239,N_6832,N_7262);
nand U9240 (N_9240,N_6561,N_7152);
and U9241 (N_9241,N_7058,N_6924);
or U9242 (N_9242,N_6677,N_6324);
or U9243 (N_9243,N_7232,N_6242);
nor U9244 (N_9244,N_6131,N_7824);
and U9245 (N_9245,N_7323,N_7479);
or U9246 (N_9246,N_7738,N_6466);
and U9247 (N_9247,N_6894,N_7331);
nand U9248 (N_9248,N_6564,N_7849);
nand U9249 (N_9249,N_7248,N_7199);
or U9250 (N_9250,N_7897,N_6533);
nor U9251 (N_9251,N_7107,N_6562);
or U9252 (N_9252,N_6723,N_6868);
nand U9253 (N_9253,N_7149,N_7673);
or U9254 (N_9254,N_7014,N_6050);
nand U9255 (N_9255,N_7716,N_7352);
nand U9256 (N_9256,N_6742,N_6295);
or U9257 (N_9257,N_7487,N_6141);
or U9258 (N_9258,N_7333,N_6344);
or U9259 (N_9259,N_7373,N_7400);
or U9260 (N_9260,N_7526,N_7749);
nor U9261 (N_9261,N_6359,N_7603);
nand U9262 (N_9262,N_7490,N_7740);
and U9263 (N_9263,N_7682,N_6118);
and U9264 (N_9264,N_6698,N_7821);
nor U9265 (N_9265,N_6219,N_7767);
nand U9266 (N_9266,N_7762,N_7048);
and U9267 (N_9267,N_6757,N_6048);
nand U9268 (N_9268,N_6351,N_7372);
nor U9269 (N_9269,N_6408,N_7159);
and U9270 (N_9270,N_6449,N_6349);
or U9271 (N_9271,N_6566,N_7558);
nor U9272 (N_9272,N_6763,N_7422);
and U9273 (N_9273,N_6550,N_6771);
nand U9274 (N_9274,N_7967,N_6937);
nor U9275 (N_9275,N_6222,N_6976);
nor U9276 (N_9276,N_7994,N_7661);
and U9277 (N_9277,N_7916,N_7764);
nor U9278 (N_9278,N_7901,N_7356);
or U9279 (N_9279,N_6135,N_6154);
nor U9280 (N_9280,N_7163,N_7887);
nor U9281 (N_9281,N_6703,N_6617);
nor U9282 (N_9282,N_7662,N_7185);
nor U9283 (N_9283,N_7415,N_7147);
or U9284 (N_9284,N_7475,N_6263);
or U9285 (N_9285,N_6354,N_7039);
and U9286 (N_9286,N_6198,N_6358);
and U9287 (N_9287,N_7252,N_6729);
nand U9288 (N_9288,N_7187,N_6984);
or U9289 (N_9289,N_6293,N_7528);
and U9290 (N_9290,N_6442,N_7564);
and U9291 (N_9291,N_7879,N_7658);
and U9292 (N_9292,N_6468,N_6742);
nand U9293 (N_9293,N_7554,N_7032);
nand U9294 (N_9294,N_6086,N_7548);
nor U9295 (N_9295,N_7653,N_7419);
and U9296 (N_9296,N_7345,N_6865);
and U9297 (N_9297,N_7348,N_7493);
and U9298 (N_9298,N_6165,N_7797);
and U9299 (N_9299,N_7627,N_7368);
nor U9300 (N_9300,N_6813,N_7289);
nand U9301 (N_9301,N_6263,N_7142);
or U9302 (N_9302,N_6787,N_6356);
nor U9303 (N_9303,N_7937,N_6743);
or U9304 (N_9304,N_6128,N_7801);
nand U9305 (N_9305,N_6444,N_6433);
and U9306 (N_9306,N_6704,N_6530);
nor U9307 (N_9307,N_6171,N_7953);
nor U9308 (N_9308,N_7783,N_7331);
nand U9309 (N_9309,N_7697,N_6041);
nor U9310 (N_9310,N_6181,N_6936);
nand U9311 (N_9311,N_6834,N_6289);
or U9312 (N_9312,N_6362,N_6582);
and U9313 (N_9313,N_6475,N_7253);
and U9314 (N_9314,N_7199,N_6219);
nor U9315 (N_9315,N_7082,N_7930);
and U9316 (N_9316,N_6127,N_6251);
and U9317 (N_9317,N_7953,N_7603);
and U9318 (N_9318,N_7463,N_7748);
or U9319 (N_9319,N_6791,N_7708);
nor U9320 (N_9320,N_7897,N_7481);
and U9321 (N_9321,N_6564,N_6352);
nor U9322 (N_9322,N_7714,N_7716);
nor U9323 (N_9323,N_7420,N_6708);
and U9324 (N_9324,N_7502,N_7003);
nor U9325 (N_9325,N_7814,N_6495);
and U9326 (N_9326,N_6241,N_7846);
nand U9327 (N_9327,N_7125,N_7560);
nand U9328 (N_9328,N_7325,N_7030);
nor U9329 (N_9329,N_6962,N_7230);
nor U9330 (N_9330,N_7883,N_6228);
or U9331 (N_9331,N_6293,N_6289);
or U9332 (N_9332,N_6609,N_7023);
nand U9333 (N_9333,N_7767,N_7838);
and U9334 (N_9334,N_7497,N_7528);
nor U9335 (N_9335,N_6479,N_7753);
nor U9336 (N_9336,N_6685,N_7718);
and U9337 (N_9337,N_7151,N_6541);
or U9338 (N_9338,N_6758,N_6799);
and U9339 (N_9339,N_6150,N_6589);
nand U9340 (N_9340,N_6567,N_6890);
or U9341 (N_9341,N_6490,N_6640);
and U9342 (N_9342,N_6872,N_7728);
and U9343 (N_9343,N_6641,N_6601);
nor U9344 (N_9344,N_6439,N_7605);
nand U9345 (N_9345,N_6379,N_7991);
or U9346 (N_9346,N_7596,N_6654);
or U9347 (N_9347,N_7184,N_7240);
nand U9348 (N_9348,N_6649,N_7494);
nor U9349 (N_9349,N_7685,N_6126);
nand U9350 (N_9350,N_7100,N_7458);
and U9351 (N_9351,N_6926,N_6510);
nor U9352 (N_9352,N_7006,N_6820);
and U9353 (N_9353,N_7434,N_7841);
or U9354 (N_9354,N_7058,N_7756);
or U9355 (N_9355,N_6730,N_6606);
nor U9356 (N_9356,N_6517,N_7664);
nor U9357 (N_9357,N_7365,N_6797);
nor U9358 (N_9358,N_6293,N_7902);
nand U9359 (N_9359,N_7477,N_6239);
nand U9360 (N_9360,N_6815,N_7040);
or U9361 (N_9361,N_6103,N_7599);
and U9362 (N_9362,N_7121,N_6253);
or U9363 (N_9363,N_7764,N_7392);
and U9364 (N_9364,N_7437,N_6997);
nor U9365 (N_9365,N_7816,N_7023);
and U9366 (N_9366,N_6351,N_7612);
nand U9367 (N_9367,N_7144,N_6184);
nand U9368 (N_9368,N_7468,N_7687);
or U9369 (N_9369,N_7707,N_6574);
nand U9370 (N_9370,N_7366,N_6160);
nand U9371 (N_9371,N_6071,N_6643);
or U9372 (N_9372,N_7357,N_7692);
nand U9373 (N_9373,N_7119,N_6952);
and U9374 (N_9374,N_7694,N_6074);
nor U9375 (N_9375,N_7257,N_7072);
nand U9376 (N_9376,N_6716,N_6686);
or U9377 (N_9377,N_7632,N_7704);
nand U9378 (N_9378,N_6059,N_6600);
nand U9379 (N_9379,N_6965,N_6446);
nand U9380 (N_9380,N_6746,N_6006);
or U9381 (N_9381,N_7301,N_7643);
and U9382 (N_9382,N_7072,N_7956);
nand U9383 (N_9383,N_6761,N_6580);
and U9384 (N_9384,N_6655,N_6823);
nor U9385 (N_9385,N_6223,N_6330);
nor U9386 (N_9386,N_6334,N_6992);
nor U9387 (N_9387,N_6950,N_6877);
nor U9388 (N_9388,N_6664,N_7669);
nor U9389 (N_9389,N_7567,N_6276);
or U9390 (N_9390,N_7880,N_6071);
nor U9391 (N_9391,N_6472,N_6712);
and U9392 (N_9392,N_6369,N_6328);
or U9393 (N_9393,N_6447,N_6630);
and U9394 (N_9394,N_7889,N_6037);
xnor U9395 (N_9395,N_6390,N_6775);
nand U9396 (N_9396,N_7214,N_6363);
and U9397 (N_9397,N_6181,N_7843);
nor U9398 (N_9398,N_7498,N_6570);
nor U9399 (N_9399,N_6442,N_6727);
nand U9400 (N_9400,N_6222,N_6661);
nor U9401 (N_9401,N_7894,N_6120);
or U9402 (N_9402,N_6841,N_7249);
or U9403 (N_9403,N_7903,N_6501);
and U9404 (N_9404,N_7371,N_7709);
and U9405 (N_9405,N_6309,N_6173);
nor U9406 (N_9406,N_6153,N_6078);
nor U9407 (N_9407,N_7917,N_7116);
and U9408 (N_9408,N_7463,N_7839);
nand U9409 (N_9409,N_7390,N_7018);
nor U9410 (N_9410,N_6810,N_6084);
nand U9411 (N_9411,N_7763,N_6601);
or U9412 (N_9412,N_6305,N_7556);
or U9413 (N_9413,N_7099,N_7997);
or U9414 (N_9414,N_7959,N_6605);
or U9415 (N_9415,N_6792,N_7521);
and U9416 (N_9416,N_6327,N_7350);
and U9417 (N_9417,N_7346,N_6380);
nor U9418 (N_9418,N_7586,N_6219);
and U9419 (N_9419,N_6983,N_6360);
nor U9420 (N_9420,N_6802,N_7330);
nor U9421 (N_9421,N_7006,N_6993);
or U9422 (N_9422,N_7557,N_7333);
and U9423 (N_9423,N_7796,N_6919);
nand U9424 (N_9424,N_7338,N_7440);
xnor U9425 (N_9425,N_7915,N_6153);
and U9426 (N_9426,N_7958,N_7225);
or U9427 (N_9427,N_7870,N_6465);
or U9428 (N_9428,N_6597,N_6692);
nor U9429 (N_9429,N_6228,N_6361);
nor U9430 (N_9430,N_7691,N_6223);
nor U9431 (N_9431,N_7114,N_6007);
and U9432 (N_9432,N_6636,N_7081);
and U9433 (N_9433,N_7519,N_6824);
and U9434 (N_9434,N_7942,N_6141);
nor U9435 (N_9435,N_6687,N_6301);
nor U9436 (N_9436,N_6052,N_7793);
xor U9437 (N_9437,N_7817,N_6459);
and U9438 (N_9438,N_6262,N_6729);
xnor U9439 (N_9439,N_6203,N_7711);
or U9440 (N_9440,N_7562,N_7612);
nand U9441 (N_9441,N_7794,N_6860);
or U9442 (N_9442,N_6944,N_6869);
or U9443 (N_9443,N_6922,N_6342);
and U9444 (N_9444,N_6618,N_6811);
nor U9445 (N_9445,N_6841,N_7986);
and U9446 (N_9446,N_7215,N_7062);
and U9447 (N_9447,N_6673,N_7058);
nand U9448 (N_9448,N_7289,N_7015);
nor U9449 (N_9449,N_7691,N_6774);
or U9450 (N_9450,N_7014,N_6234);
nor U9451 (N_9451,N_6243,N_6549);
nor U9452 (N_9452,N_7670,N_6359);
or U9453 (N_9453,N_6174,N_6575);
or U9454 (N_9454,N_7404,N_6451);
and U9455 (N_9455,N_6735,N_6309);
nand U9456 (N_9456,N_6567,N_7726);
or U9457 (N_9457,N_6481,N_7572);
nor U9458 (N_9458,N_6273,N_7839);
nor U9459 (N_9459,N_7833,N_7818);
nand U9460 (N_9460,N_7175,N_7236);
or U9461 (N_9461,N_6225,N_7495);
nand U9462 (N_9462,N_6331,N_6637);
nand U9463 (N_9463,N_7736,N_7975);
or U9464 (N_9464,N_7928,N_6557);
and U9465 (N_9465,N_7608,N_6773);
or U9466 (N_9466,N_6826,N_6093);
and U9467 (N_9467,N_7850,N_7945);
nor U9468 (N_9468,N_6038,N_6421);
or U9469 (N_9469,N_7299,N_6384);
or U9470 (N_9470,N_6965,N_6857);
and U9471 (N_9471,N_7121,N_7323);
nor U9472 (N_9472,N_7894,N_7196);
nor U9473 (N_9473,N_7007,N_6570);
and U9474 (N_9474,N_7759,N_6285);
nor U9475 (N_9475,N_6745,N_7222);
and U9476 (N_9476,N_6256,N_7718);
nand U9477 (N_9477,N_6286,N_7981);
and U9478 (N_9478,N_7704,N_7785);
or U9479 (N_9479,N_7230,N_7728);
or U9480 (N_9480,N_7742,N_6902);
nand U9481 (N_9481,N_6972,N_6433);
nand U9482 (N_9482,N_7176,N_7994);
nand U9483 (N_9483,N_6670,N_6691);
and U9484 (N_9484,N_6833,N_6343);
nand U9485 (N_9485,N_6349,N_6423);
or U9486 (N_9486,N_6738,N_6458);
and U9487 (N_9487,N_7334,N_7004);
nor U9488 (N_9488,N_7398,N_7835);
or U9489 (N_9489,N_7482,N_6567);
or U9490 (N_9490,N_6900,N_7382);
nand U9491 (N_9491,N_6453,N_6278);
or U9492 (N_9492,N_7824,N_6213);
and U9493 (N_9493,N_7902,N_6617);
nand U9494 (N_9494,N_6853,N_7524);
or U9495 (N_9495,N_6626,N_6854);
and U9496 (N_9496,N_7940,N_7632);
nand U9497 (N_9497,N_6450,N_6872);
and U9498 (N_9498,N_7582,N_6979);
nor U9499 (N_9499,N_7340,N_7007);
and U9500 (N_9500,N_6932,N_6806);
and U9501 (N_9501,N_6733,N_6312);
or U9502 (N_9502,N_6818,N_6798);
or U9503 (N_9503,N_6506,N_7102);
or U9504 (N_9504,N_6159,N_6956);
or U9505 (N_9505,N_7740,N_6901);
and U9506 (N_9506,N_6434,N_6035);
and U9507 (N_9507,N_7642,N_6344);
nor U9508 (N_9508,N_6476,N_6473);
and U9509 (N_9509,N_6717,N_6102);
nand U9510 (N_9510,N_6025,N_6751);
or U9511 (N_9511,N_7243,N_7359);
nand U9512 (N_9512,N_7245,N_7526);
nor U9513 (N_9513,N_7314,N_7370);
nand U9514 (N_9514,N_7579,N_6562);
or U9515 (N_9515,N_7776,N_7102);
nand U9516 (N_9516,N_6472,N_7738);
or U9517 (N_9517,N_7907,N_6027);
nand U9518 (N_9518,N_6009,N_6108);
nor U9519 (N_9519,N_6378,N_6711);
or U9520 (N_9520,N_6343,N_6465);
or U9521 (N_9521,N_7864,N_6433);
and U9522 (N_9522,N_6906,N_6978);
nand U9523 (N_9523,N_7019,N_7567);
nor U9524 (N_9524,N_7349,N_6111);
nand U9525 (N_9525,N_7412,N_6285);
and U9526 (N_9526,N_6411,N_6168);
or U9527 (N_9527,N_6325,N_6011);
nor U9528 (N_9528,N_7962,N_7511);
nand U9529 (N_9529,N_6492,N_7253);
nand U9530 (N_9530,N_6877,N_7846);
nor U9531 (N_9531,N_6933,N_7822);
and U9532 (N_9532,N_7647,N_6641);
and U9533 (N_9533,N_7762,N_7106);
nor U9534 (N_9534,N_7231,N_7558);
nand U9535 (N_9535,N_6490,N_7828);
nor U9536 (N_9536,N_7626,N_6071);
or U9537 (N_9537,N_7530,N_7164);
or U9538 (N_9538,N_6523,N_7502);
and U9539 (N_9539,N_6345,N_6566);
and U9540 (N_9540,N_6048,N_7416);
and U9541 (N_9541,N_6149,N_7568);
nor U9542 (N_9542,N_7242,N_7723);
nor U9543 (N_9543,N_6603,N_7080);
and U9544 (N_9544,N_6798,N_7457);
nor U9545 (N_9545,N_6489,N_6086);
or U9546 (N_9546,N_7135,N_6064);
nand U9547 (N_9547,N_7953,N_6457);
or U9548 (N_9548,N_6537,N_7623);
and U9549 (N_9549,N_7750,N_6815);
and U9550 (N_9550,N_6348,N_7752);
and U9551 (N_9551,N_7162,N_7062);
or U9552 (N_9552,N_6090,N_7300);
nor U9553 (N_9553,N_7391,N_7488);
or U9554 (N_9554,N_7226,N_7711);
nand U9555 (N_9555,N_6930,N_7182);
nand U9556 (N_9556,N_7754,N_6681);
nor U9557 (N_9557,N_7202,N_6406);
and U9558 (N_9558,N_6899,N_7367);
nand U9559 (N_9559,N_6615,N_6414);
and U9560 (N_9560,N_7844,N_7469);
nand U9561 (N_9561,N_7078,N_7892);
nor U9562 (N_9562,N_6164,N_6383);
nand U9563 (N_9563,N_7311,N_7504);
and U9564 (N_9564,N_7722,N_6067);
nor U9565 (N_9565,N_7558,N_6984);
nand U9566 (N_9566,N_7255,N_7609);
or U9567 (N_9567,N_7301,N_6370);
or U9568 (N_9568,N_7183,N_6730);
nand U9569 (N_9569,N_6942,N_6780);
and U9570 (N_9570,N_7744,N_6969);
and U9571 (N_9571,N_7581,N_7974);
and U9572 (N_9572,N_6671,N_7319);
nor U9573 (N_9573,N_7328,N_7539);
nor U9574 (N_9574,N_6941,N_6041);
or U9575 (N_9575,N_6224,N_7881);
or U9576 (N_9576,N_7765,N_6625);
nor U9577 (N_9577,N_6720,N_6582);
or U9578 (N_9578,N_6736,N_6547);
or U9579 (N_9579,N_7089,N_6639);
or U9580 (N_9580,N_6110,N_7200);
nand U9581 (N_9581,N_7416,N_6792);
or U9582 (N_9582,N_7938,N_7727);
nand U9583 (N_9583,N_6764,N_6051);
or U9584 (N_9584,N_7861,N_7352);
and U9585 (N_9585,N_6979,N_7929);
or U9586 (N_9586,N_6659,N_7410);
nand U9587 (N_9587,N_7664,N_7550);
or U9588 (N_9588,N_6444,N_7471);
or U9589 (N_9589,N_7144,N_6187);
nor U9590 (N_9590,N_7021,N_7598);
or U9591 (N_9591,N_7345,N_7534);
and U9592 (N_9592,N_6195,N_7533);
or U9593 (N_9593,N_7075,N_7764);
and U9594 (N_9594,N_7954,N_6584);
or U9595 (N_9595,N_6580,N_7658);
nor U9596 (N_9596,N_6755,N_7842);
nand U9597 (N_9597,N_7435,N_6723);
and U9598 (N_9598,N_6370,N_6028);
or U9599 (N_9599,N_7352,N_7794);
and U9600 (N_9600,N_6825,N_7662);
or U9601 (N_9601,N_7222,N_6822);
and U9602 (N_9602,N_6798,N_6363);
nand U9603 (N_9603,N_6268,N_7944);
and U9604 (N_9604,N_7946,N_7455);
nor U9605 (N_9605,N_6089,N_7782);
or U9606 (N_9606,N_7637,N_6166);
nor U9607 (N_9607,N_6738,N_6820);
nand U9608 (N_9608,N_6584,N_7514);
or U9609 (N_9609,N_6271,N_7680);
nor U9610 (N_9610,N_7362,N_6431);
nor U9611 (N_9611,N_7189,N_7186);
nand U9612 (N_9612,N_6277,N_7353);
nand U9613 (N_9613,N_7641,N_7070);
nand U9614 (N_9614,N_7413,N_6291);
and U9615 (N_9615,N_7105,N_6334);
nand U9616 (N_9616,N_6075,N_7224);
nor U9617 (N_9617,N_7815,N_7136);
nor U9618 (N_9618,N_7012,N_6496);
nor U9619 (N_9619,N_7869,N_7996);
xnor U9620 (N_9620,N_6939,N_7441);
and U9621 (N_9621,N_7654,N_6024);
and U9622 (N_9622,N_6118,N_7382);
and U9623 (N_9623,N_6771,N_6577);
or U9624 (N_9624,N_7948,N_7365);
and U9625 (N_9625,N_7600,N_7662);
or U9626 (N_9626,N_7910,N_6127);
or U9627 (N_9627,N_7295,N_6189);
nand U9628 (N_9628,N_7172,N_7331);
or U9629 (N_9629,N_7474,N_6907);
nor U9630 (N_9630,N_7685,N_7793);
nand U9631 (N_9631,N_7800,N_6830);
nand U9632 (N_9632,N_6710,N_7167);
and U9633 (N_9633,N_6741,N_6560);
nor U9634 (N_9634,N_7876,N_7310);
and U9635 (N_9635,N_6164,N_7211);
or U9636 (N_9636,N_6994,N_6963);
and U9637 (N_9637,N_6098,N_7514);
and U9638 (N_9638,N_6736,N_6522);
or U9639 (N_9639,N_6630,N_6195);
and U9640 (N_9640,N_6611,N_7783);
xnor U9641 (N_9641,N_7456,N_6852);
and U9642 (N_9642,N_7608,N_7238);
nor U9643 (N_9643,N_7591,N_6611);
and U9644 (N_9644,N_6457,N_7147);
and U9645 (N_9645,N_7427,N_6098);
nor U9646 (N_9646,N_6376,N_7827);
or U9647 (N_9647,N_7582,N_7626);
or U9648 (N_9648,N_7603,N_6779);
nor U9649 (N_9649,N_6199,N_7608);
or U9650 (N_9650,N_7343,N_6967);
nor U9651 (N_9651,N_7009,N_6883);
nor U9652 (N_9652,N_7282,N_6562);
nand U9653 (N_9653,N_7608,N_6070);
and U9654 (N_9654,N_6745,N_7872);
and U9655 (N_9655,N_6032,N_7137);
or U9656 (N_9656,N_7943,N_6256);
nor U9657 (N_9657,N_7499,N_7370);
or U9658 (N_9658,N_7646,N_6390);
and U9659 (N_9659,N_7184,N_7818);
nand U9660 (N_9660,N_7140,N_6801);
nand U9661 (N_9661,N_6952,N_6381);
nor U9662 (N_9662,N_6948,N_6273);
nand U9663 (N_9663,N_7154,N_6919);
nand U9664 (N_9664,N_7838,N_7947);
nor U9665 (N_9665,N_6138,N_7780);
and U9666 (N_9666,N_7871,N_7795);
nor U9667 (N_9667,N_7648,N_7747);
or U9668 (N_9668,N_7957,N_7903);
nor U9669 (N_9669,N_7231,N_7050);
nand U9670 (N_9670,N_7016,N_6834);
nand U9671 (N_9671,N_6638,N_6589);
nand U9672 (N_9672,N_7836,N_6032);
and U9673 (N_9673,N_6751,N_6183);
nand U9674 (N_9674,N_6276,N_6191);
and U9675 (N_9675,N_6566,N_7211);
nor U9676 (N_9676,N_7173,N_6779);
nor U9677 (N_9677,N_6122,N_7892);
or U9678 (N_9678,N_7691,N_7761);
nor U9679 (N_9679,N_7559,N_6924);
or U9680 (N_9680,N_7100,N_7704);
and U9681 (N_9681,N_7848,N_7872);
or U9682 (N_9682,N_7797,N_6532);
or U9683 (N_9683,N_6779,N_6962);
or U9684 (N_9684,N_7959,N_7053);
or U9685 (N_9685,N_7897,N_7891);
nor U9686 (N_9686,N_6188,N_6132);
nor U9687 (N_9687,N_6980,N_7908);
nor U9688 (N_9688,N_6349,N_6785);
nor U9689 (N_9689,N_6980,N_6862);
nor U9690 (N_9690,N_6520,N_7071);
nand U9691 (N_9691,N_6224,N_7974);
nand U9692 (N_9692,N_7419,N_6537);
nand U9693 (N_9693,N_7263,N_7773);
nand U9694 (N_9694,N_6516,N_6505);
nand U9695 (N_9695,N_6534,N_6559);
or U9696 (N_9696,N_7761,N_6789);
nand U9697 (N_9697,N_6750,N_6400);
nor U9698 (N_9698,N_6779,N_6478);
nand U9699 (N_9699,N_7331,N_6839);
or U9700 (N_9700,N_7679,N_6156);
nand U9701 (N_9701,N_6576,N_7195);
nand U9702 (N_9702,N_7745,N_7089);
or U9703 (N_9703,N_6246,N_6024);
and U9704 (N_9704,N_7283,N_6593);
nor U9705 (N_9705,N_6166,N_6899);
and U9706 (N_9706,N_6740,N_6262);
nand U9707 (N_9707,N_7681,N_7011);
nand U9708 (N_9708,N_7373,N_7104);
and U9709 (N_9709,N_6608,N_7826);
nand U9710 (N_9710,N_7338,N_7457);
nand U9711 (N_9711,N_6119,N_7892);
or U9712 (N_9712,N_7149,N_6209);
or U9713 (N_9713,N_6968,N_6612);
nor U9714 (N_9714,N_6140,N_7973);
nand U9715 (N_9715,N_7745,N_6589);
nor U9716 (N_9716,N_7448,N_7843);
or U9717 (N_9717,N_7414,N_6695);
or U9718 (N_9718,N_6251,N_6079);
nor U9719 (N_9719,N_6826,N_6095);
or U9720 (N_9720,N_6392,N_7549);
or U9721 (N_9721,N_7314,N_6063);
or U9722 (N_9722,N_6722,N_7089);
nand U9723 (N_9723,N_6144,N_6148);
nand U9724 (N_9724,N_6557,N_6479);
or U9725 (N_9725,N_7733,N_7742);
and U9726 (N_9726,N_7750,N_7273);
nor U9727 (N_9727,N_7653,N_7889);
nor U9728 (N_9728,N_7553,N_6287);
and U9729 (N_9729,N_6678,N_6639);
nor U9730 (N_9730,N_6421,N_6786);
nand U9731 (N_9731,N_6980,N_6913);
and U9732 (N_9732,N_6713,N_7387);
nand U9733 (N_9733,N_7804,N_6974);
nor U9734 (N_9734,N_6688,N_6880);
nor U9735 (N_9735,N_6594,N_7893);
nor U9736 (N_9736,N_6156,N_7625);
or U9737 (N_9737,N_6514,N_7777);
or U9738 (N_9738,N_7987,N_7114);
nand U9739 (N_9739,N_7218,N_6439);
nor U9740 (N_9740,N_7754,N_6809);
nand U9741 (N_9741,N_6362,N_6891);
nor U9742 (N_9742,N_7868,N_7073);
or U9743 (N_9743,N_6885,N_6312);
nand U9744 (N_9744,N_7833,N_6048);
nor U9745 (N_9745,N_6530,N_6355);
nand U9746 (N_9746,N_7301,N_6556);
and U9747 (N_9747,N_7205,N_7410);
nand U9748 (N_9748,N_6230,N_6391);
or U9749 (N_9749,N_6404,N_7593);
and U9750 (N_9750,N_7058,N_6433);
nand U9751 (N_9751,N_7998,N_6680);
nor U9752 (N_9752,N_6673,N_7165);
nand U9753 (N_9753,N_6199,N_7671);
nor U9754 (N_9754,N_6708,N_6477);
nor U9755 (N_9755,N_7155,N_7227);
nand U9756 (N_9756,N_7727,N_7818);
and U9757 (N_9757,N_7038,N_7397);
nor U9758 (N_9758,N_7800,N_7400);
nand U9759 (N_9759,N_7473,N_6730);
nand U9760 (N_9760,N_6007,N_6078);
and U9761 (N_9761,N_6226,N_7434);
or U9762 (N_9762,N_6840,N_7955);
and U9763 (N_9763,N_6628,N_7689);
and U9764 (N_9764,N_7006,N_6595);
nand U9765 (N_9765,N_6338,N_7820);
nand U9766 (N_9766,N_7357,N_7151);
nand U9767 (N_9767,N_7055,N_6532);
and U9768 (N_9768,N_6466,N_6674);
nand U9769 (N_9769,N_6541,N_6301);
nor U9770 (N_9770,N_7384,N_7074);
nor U9771 (N_9771,N_6049,N_7027);
or U9772 (N_9772,N_6827,N_6817);
nor U9773 (N_9773,N_7587,N_7076);
or U9774 (N_9774,N_6045,N_7831);
or U9775 (N_9775,N_6672,N_6665);
or U9776 (N_9776,N_6312,N_6414);
and U9777 (N_9777,N_7879,N_6000);
nand U9778 (N_9778,N_7849,N_7809);
nor U9779 (N_9779,N_7468,N_7412);
and U9780 (N_9780,N_6984,N_6409);
and U9781 (N_9781,N_7824,N_6540);
nor U9782 (N_9782,N_6215,N_7395);
nand U9783 (N_9783,N_7206,N_7145);
or U9784 (N_9784,N_7917,N_7774);
nor U9785 (N_9785,N_6656,N_6389);
nand U9786 (N_9786,N_7532,N_6475);
or U9787 (N_9787,N_7454,N_7088);
nor U9788 (N_9788,N_6346,N_7290);
or U9789 (N_9789,N_7215,N_6844);
or U9790 (N_9790,N_7261,N_6849);
nor U9791 (N_9791,N_7839,N_6626);
nand U9792 (N_9792,N_6521,N_6084);
and U9793 (N_9793,N_7525,N_7719);
nor U9794 (N_9794,N_7611,N_7729);
or U9795 (N_9795,N_6473,N_7971);
nand U9796 (N_9796,N_7227,N_7240);
or U9797 (N_9797,N_6011,N_7739);
and U9798 (N_9798,N_7551,N_6448);
nand U9799 (N_9799,N_7129,N_7719);
nand U9800 (N_9800,N_6866,N_7221);
or U9801 (N_9801,N_6360,N_7815);
or U9802 (N_9802,N_7020,N_6261);
or U9803 (N_9803,N_6604,N_7582);
or U9804 (N_9804,N_7390,N_6663);
and U9805 (N_9805,N_6038,N_7420);
nand U9806 (N_9806,N_6455,N_7562);
nor U9807 (N_9807,N_6334,N_6893);
nor U9808 (N_9808,N_6435,N_7585);
and U9809 (N_9809,N_7175,N_6600);
or U9810 (N_9810,N_6968,N_7318);
and U9811 (N_9811,N_6877,N_7928);
nor U9812 (N_9812,N_7677,N_6709);
nor U9813 (N_9813,N_6591,N_7847);
nand U9814 (N_9814,N_6702,N_7244);
xnor U9815 (N_9815,N_6380,N_6241);
nor U9816 (N_9816,N_6478,N_7622);
or U9817 (N_9817,N_6704,N_7602);
or U9818 (N_9818,N_6436,N_6959);
or U9819 (N_9819,N_6826,N_6240);
or U9820 (N_9820,N_7019,N_6133);
nand U9821 (N_9821,N_7794,N_6076);
and U9822 (N_9822,N_6474,N_6468);
and U9823 (N_9823,N_6098,N_7937);
nor U9824 (N_9824,N_6371,N_6546);
and U9825 (N_9825,N_7620,N_6074);
nand U9826 (N_9826,N_6155,N_7633);
and U9827 (N_9827,N_6658,N_6270);
nand U9828 (N_9828,N_6989,N_6284);
nand U9829 (N_9829,N_7814,N_6220);
or U9830 (N_9830,N_7701,N_6369);
and U9831 (N_9831,N_7976,N_7433);
nand U9832 (N_9832,N_7339,N_6955);
nor U9833 (N_9833,N_7376,N_6041);
nor U9834 (N_9834,N_7980,N_7146);
or U9835 (N_9835,N_7033,N_7155);
nor U9836 (N_9836,N_7490,N_7449);
nor U9837 (N_9837,N_7180,N_7284);
nor U9838 (N_9838,N_6896,N_7033);
nand U9839 (N_9839,N_7059,N_7269);
or U9840 (N_9840,N_6409,N_7268);
nor U9841 (N_9841,N_6923,N_6455);
and U9842 (N_9842,N_7421,N_6154);
nand U9843 (N_9843,N_7770,N_6894);
or U9844 (N_9844,N_7800,N_7093);
or U9845 (N_9845,N_7661,N_6238);
xor U9846 (N_9846,N_7053,N_6928);
and U9847 (N_9847,N_7636,N_7994);
nand U9848 (N_9848,N_6005,N_7472);
nor U9849 (N_9849,N_6717,N_7504);
nor U9850 (N_9850,N_6153,N_6421);
nor U9851 (N_9851,N_6239,N_7145);
or U9852 (N_9852,N_7610,N_6246);
nor U9853 (N_9853,N_7927,N_6671);
nor U9854 (N_9854,N_6604,N_7279);
and U9855 (N_9855,N_7264,N_6564);
nor U9856 (N_9856,N_6878,N_6288);
nor U9857 (N_9857,N_6891,N_7616);
nor U9858 (N_9858,N_7604,N_7640);
and U9859 (N_9859,N_6738,N_6733);
nand U9860 (N_9860,N_7286,N_7118);
and U9861 (N_9861,N_6668,N_6971);
nor U9862 (N_9862,N_7858,N_7526);
nand U9863 (N_9863,N_7182,N_6855);
nand U9864 (N_9864,N_7381,N_6724);
nand U9865 (N_9865,N_7001,N_7156);
nor U9866 (N_9866,N_6861,N_7956);
and U9867 (N_9867,N_6587,N_7223);
nand U9868 (N_9868,N_7982,N_6565);
or U9869 (N_9869,N_6042,N_7725);
or U9870 (N_9870,N_7167,N_6316);
nand U9871 (N_9871,N_7725,N_6139);
and U9872 (N_9872,N_6235,N_7665);
or U9873 (N_9873,N_7271,N_7337);
nand U9874 (N_9874,N_6112,N_7836);
nand U9875 (N_9875,N_6327,N_6856);
and U9876 (N_9876,N_6326,N_7075);
and U9877 (N_9877,N_7424,N_6846);
and U9878 (N_9878,N_6403,N_7974);
or U9879 (N_9879,N_7510,N_7941);
or U9880 (N_9880,N_6901,N_6935);
or U9881 (N_9881,N_6890,N_7947);
nor U9882 (N_9882,N_6015,N_7912);
or U9883 (N_9883,N_6093,N_6327);
nand U9884 (N_9884,N_6419,N_7466);
or U9885 (N_9885,N_7135,N_6444);
nor U9886 (N_9886,N_6542,N_6908);
and U9887 (N_9887,N_7232,N_7003);
or U9888 (N_9888,N_7230,N_7944);
or U9889 (N_9889,N_7213,N_6446);
nor U9890 (N_9890,N_7198,N_7130);
or U9891 (N_9891,N_7318,N_6794);
or U9892 (N_9892,N_6122,N_7173);
or U9893 (N_9893,N_7701,N_7690);
and U9894 (N_9894,N_6992,N_6858);
and U9895 (N_9895,N_6727,N_6166);
nor U9896 (N_9896,N_6378,N_6234);
or U9897 (N_9897,N_6453,N_7565);
and U9898 (N_9898,N_7850,N_6279);
and U9899 (N_9899,N_6191,N_6516);
nor U9900 (N_9900,N_7765,N_7322);
nand U9901 (N_9901,N_6081,N_7096);
nand U9902 (N_9902,N_7242,N_7706);
and U9903 (N_9903,N_6213,N_7933);
nand U9904 (N_9904,N_6131,N_7996);
nand U9905 (N_9905,N_7448,N_6743);
or U9906 (N_9906,N_7266,N_6153);
nand U9907 (N_9907,N_7767,N_6846);
and U9908 (N_9908,N_7980,N_6603);
and U9909 (N_9909,N_6793,N_6065);
nor U9910 (N_9910,N_7558,N_6462);
and U9911 (N_9911,N_7811,N_7917);
or U9912 (N_9912,N_7303,N_7445);
or U9913 (N_9913,N_6594,N_6623);
nand U9914 (N_9914,N_6206,N_6130);
and U9915 (N_9915,N_7953,N_6468);
and U9916 (N_9916,N_6602,N_7106);
or U9917 (N_9917,N_6583,N_6952);
or U9918 (N_9918,N_7710,N_7480);
or U9919 (N_9919,N_6143,N_7203);
nand U9920 (N_9920,N_6340,N_6933);
nand U9921 (N_9921,N_7397,N_6186);
nor U9922 (N_9922,N_6130,N_6767);
and U9923 (N_9923,N_7301,N_7587);
or U9924 (N_9924,N_6417,N_7191);
and U9925 (N_9925,N_7230,N_6503);
and U9926 (N_9926,N_7768,N_6591);
and U9927 (N_9927,N_6315,N_7228);
and U9928 (N_9928,N_6773,N_6396);
nand U9929 (N_9929,N_7119,N_7635);
and U9930 (N_9930,N_6887,N_7429);
nor U9931 (N_9931,N_6962,N_7891);
nor U9932 (N_9932,N_6756,N_6352);
and U9933 (N_9933,N_7805,N_6087);
xor U9934 (N_9934,N_6680,N_6352);
and U9935 (N_9935,N_6608,N_6403);
or U9936 (N_9936,N_6115,N_6147);
nand U9937 (N_9937,N_7387,N_7380);
and U9938 (N_9938,N_7813,N_6791);
nand U9939 (N_9939,N_6194,N_7703);
or U9940 (N_9940,N_7356,N_7963);
nand U9941 (N_9941,N_6983,N_6892);
or U9942 (N_9942,N_7541,N_7299);
nand U9943 (N_9943,N_6490,N_7279);
nor U9944 (N_9944,N_6701,N_7462);
and U9945 (N_9945,N_7391,N_7634);
or U9946 (N_9946,N_7095,N_7003);
nor U9947 (N_9947,N_6440,N_6377);
and U9948 (N_9948,N_7954,N_7962);
and U9949 (N_9949,N_6205,N_7305);
and U9950 (N_9950,N_6980,N_6598);
nand U9951 (N_9951,N_7731,N_7232);
or U9952 (N_9952,N_6740,N_7287);
nor U9953 (N_9953,N_7485,N_7609);
and U9954 (N_9954,N_6159,N_6632);
and U9955 (N_9955,N_7016,N_6516);
nand U9956 (N_9956,N_6137,N_7112);
or U9957 (N_9957,N_7343,N_7799);
nor U9958 (N_9958,N_7070,N_7335);
and U9959 (N_9959,N_6549,N_6736);
and U9960 (N_9960,N_7367,N_7959);
or U9961 (N_9961,N_6372,N_7557);
and U9962 (N_9962,N_7202,N_6277);
and U9963 (N_9963,N_6740,N_6858);
and U9964 (N_9964,N_6086,N_7305);
and U9965 (N_9965,N_6217,N_6097);
and U9966 (N_9966,N_6811,N_7266);
or U9967 (N_9967,N_6561,N_7046);
and U9968 (N_9968,N_6245,N_7384);
and U9969 (N_9969,N_6668,N_7464);
or U9970 (N_9970,N_6060,N_6216);
and U9971 (N_9971,N_6693,N_7936);
and U9972 (N_9972,N_6375,N_6744);
and U9973 (N_9973,N_6659,N_6315);
nand U9974 (N_9974,N_7944,N_6576);
and U9975 (N_9975,N_7524,N_6343);
nor U9976 (N_9976,N_7967,N_6373);
or U9977 (N_9977,N_6038,N_7135);
nand U9978 (N_9978,N_7846,N_6829);
nand U9979 (N_9979,N_6022,N_6681);
or U9980 (N_9980,N_6439,N_6713);
nand U9981 (N_9981,N_7416,N_6201);
or U9982 (N_9982,N_6145,N_7817);
or U9983 (N_9983,N_6205,N_6670);
and U9984 (N_9984,N_6040,N_7707);
and U9985 (N_9985,N_7682,N_6929);
nand U9986 (N_9986,N_6256,N_6155);
and U9987 (N_9987,N_7432,N_7764);
nand U9988 (N_9988,N_7480,N_6785);
nand U9989 (N_9989,N_7968,N_6696);
nand U9990 (N_9990,N_7130,N_6366);
nand U9991 (N_9991,N_7882,N_6182);
nand U9992 (N_9992,N_7904,N_7349);
nor U9993 (N_9993,N_6063,N_7735);
nor U9994 (N_9994,N_7846,N_6936);
or U9995 (N_9995,N_6031,N_6096);
or U9996 (N_9996,N_6050,N_7509);
nand U9997 (N_9997,N_7767,N_7957);
nand U9998 (N_9998,N_7864,N_6281);
and U9999 (N_9999,N_7755,N_7974);
nand UO_0 (O_0,N_9363,N_8849);
and UO_1 (O_1,N_9354,N_9880);
or UO_2 (O_2,N_9488,N_8780);
nand UO_3 (O_3,N_8594,N_9955);
nand UO_4 (O_4,N_8407,N_8256);
nor UO_5 (O_5,N_8518,N_9306);
or UO_6 (O_6,N_8272,N_8588);
nor UO_7 (O_7,N_9201,N_8776);
and UO_8 (O_8,N_9774,N_9501);
and UO_9 (O_9,N_8522,N_8812);
nand UO_10 (O_10,N_9924,N_8612);
nand UO_11 (O_11,N_8335,N_9146);
or UO_12 (O_12,N_9797,N_9013);
nor UO_13 (O_13,N_9632,N_8135);
and UO_14 (O_14,N_8813,N_8241);
and UO_15 (O_15,N_9034,N_9159);
nor UO_16 (O_16,N_8056,N_9929);
nor UO_17 (O_17,N_9733,N_8419);
or UO_18 (O_18,N_9224,N_9826);
nand UO_19 (O_19,N_9556,N_8327);
or UO_20 (O_20,N_9567,N_8159);
nor UO_21 (O_21,N_9435,N_9782);
nor UO_22 (O_22,N_9220,N_9778);
or UO_23 (O_23,N_9407,N_8942);
and UO_24 (O_24,N_9158,N_9859);
or UO_25 (O_25,N_8834,N_8699);
or UO_26 (O_26,N_9063,N_8300);
and UO_27 (O_27,N_9537,N_9545);
and UO_28 (O_28,N_8158,N_8284);
and UO_29 (O_29,N_8265,N_8662);
and UO_30 (O_30,N_9166,N_9033);
nand UO_31 (O_31,N_8477,N_8986);
nand UO_32 (O_32,N_9142,N_8050);
or UO_33 (O_33,N_9236,N_9311);
and UO_34 (O_34,N_9706,N_8784);
or UO_35 (O_35,N_8826,N_9934);
and UO_36 (O_36,N_8862,N_9234);
and UO_37 (O_37,N_9599,N_9834);
nor UO_38 (O_38,N_9522,N_9066);
nand UO_39 (O_39,N_9564,N_9662);
nor UO_40 (O_40,N_9459,N_9770);
nor UO_41 (O_41,N_9839,N_8153);
and UO_42 (O_42,N_8424,N_9412);
or UO_43 (O_43,N_9669,N_9956);
or UO_44 (O_44,N_8463,N_9173);
nand UO_45 (O_45,N_8114,N_9205);
or UO_46 (O_46,N_9796,N_9865);
xnor UO_47 (O_47,N_9560,N_9195);
nor UO_48 (O_48,N_8680,N_8336);
and UO_49 (O_49,N_9993,N_9252);
and UO_50 (O_50,N_9894,N_8352);
and UO_51 (O_51,N_9029,N_8916);
and UO_52 (O_52,N_9485,N_9366);
or UO_53 (O_53,N_8537,N_8372);
nand UO_54 (O_54,N_8868,N_8166);
nand UO_55 (O_55,N_9727,N_9190);
and UO_56 (O_56,N_9020,N_9153);
and UO_57 (O_57,N_9926,N_9010);
nand UO_58 (O_58,N_9845,N_8276);
and UO_59 (O_59,N_8016,N_9584);
nor UO_60 (O_60,N_9886,N_9810);
nand UO_61 (O_61,N_8347,N_8240);
nand UO_62 (O_62,N_9285,N_8572);
nand UO_63 (O_63,N_9474,N_9805);
and UO_64 (O_64,N_9215,N_8179);
or UO_65 (O_65,N_8669,N_8764);
nor UO_66 (O_66,N_8449,N_9572);
nand UO_67 (O_67,N_8033,N_8546);
or UO_68 (O_68,N_8438,N_8028);
nand UO_69 (O_69,N_8478,N_9822);
nor UO_70 (O_70,N_9512,N_9719);
or UO_71 (O_71,N_9581,N_8896);
nand UO_72 (O_72,N_9301,N_9809);
and UO_73 (O_73,N_9611,N_8009);
nand UO_74 (O_74,N_9574,N_9896);
nor UO_75 (O_75,N_9766,N_8182);
and UO_76 (O_76,N_9469,N_8941);
or UO_77 (O_77,N_9867,N_9253);
nand UO_78 (O_78,N_8138,N_9247);
nor UO_79 (O_79,N_8509,N_9053);
xor UO_80 (O_80,N_8185,N_8589);
nor UO_81 (O_81,N_8386,N_9788);
and UO_82 (O_82,N_8340,N_8674);
or UO_83 (O_83,N_8548,N_9911);
or UO_84 (O_84,N_9019,N_8991);
nand UO_85 (O_85,N_9089,N_9273);
nor UO_86 (O_86,N_8931,N_8006);
nand UO_87 (O_87,N_9418,N_8750);
nand UO_88 (O_88,N_9267,N_8183);
and UO_89 (O_89,N_9704,N_9232);
xnor UO_90 (O_90,N_8793,N_9198);
nor UO_91 (O_91,N_8308,N_8306);
and UO_92 (O_92,N_9295,N_8876);
nor UO_93 (O_93,N_9968,N_8057);
nand UO_94 (O_94,N_8687,N_8609);
or UO_95 (O_95,N_9106,N_9051);
nand UO_96 (O_96,N_8365,N_8923);
or UO_97 (O_97,N_9180,N_8553);
or UO_98 (O_98,N_8133,N_8520);
nand UO_99 (O_99,N_8037,N_8606);
nor UO_100 (O_100,N_8137,N_9851);
nand UO_101 (O_101,N_9745,N_9933);
nand UO_102 (O_102,N_8889,N_9124);
nand UO_103 (O_103,N_8301,N_8429);
nor UO_104 (O_104,N_8038,N_9920);
nor UO_105 (O_105,N_9773,N_9039);
or UO_106 (O_106,N_9950,N_9561);
nor UO_107 (O_107,N_8355,N_9907);
nand UO_108 (O_108,N_8026,N_9134);
nand UO_109 (O_109,N_8995,N_8186);
or UO_110 (O_110,N_8011,N_8852);
nand UO_111 (O_111,N_8229,N_8385);
nor UO_112 (O_112,N_8632,N_9111);
nand UO_113 (O_113,N_9084,N_8154);
and UO_114 (O_114,N_9888,N_9948);
nand UO_115 (O_115,N_9589,N_9401);
and UO_116 (O_116,N_8358,N_8543);
nor UO_117 (O_117,N_8302,N_9470);
nand UO_118 (O_118,N_8789,N_8967);
and UO_119 (O_119,N_8078,N_9712);
nand UO_120 (O_120,N_8234,N_8310);
nand UO_121 (O_121,N_8072,N_9375);
or UO_122 (O_122,N_8112,N_8743);
and UO_123 (O_123,N_9223,N_8255);
or UO_124 (O_124,N_8107,N_8953);
xnor UO_125 (O_125,N_8309,N_8101);
and UO_126 (O_126,N_8118,N_8314);
nor UO_127 (O_127,N_8432,N_9447);
nor UO_128 (O_128,N_8875,N_9622);
nor UO_129 (O_129,N_9991,N_9693);
nand UO_130 (O_130,N_9972,N_8911);
nor UO_131 (O_131,N_9879,N_9518);
and UO_132 (O_132,N_8701,N_9453);
nand UO_133 (O_133,N_8927,N_8773);
nand UO_134 (O_134,N_9131,N_8210);
or UO_135 (O_135,N_9898,N_8748);
nor UO_136 (O_136,N_9428,N_9919);
and UO_137 (O_137,N_8587,N_8192);
or UO_138 (O_138,N_9332,N_8295);
nand UO_139 (O_139,N_9061,N_8469);
nand UO_140 (O_140,N_8581,N_9214);
or UO_141 (O_141,N_9484,N_8913);
or UO_142 (O_142,N_9597,N_9024);
and UO_143 (O_143,N_9498,N_8547);
nand UO_144 (O_144,N_9906,N_8541);
or UO_145 (O_145,N_9709,N_9272);
and UO_146 (O_146,N_8966,N_8874);
or UO_147 (O_147,N_8517,N_8257);
or UO_148 (O_148,N_9482,N_9682);
nand UO_149 (O_149,N_8400,N_8245);
and UO_150 (O_150,N_8956,N_8232);
nor UO_151 (O_151,N_9877,N_9566);
or UO_152 (O_152,N_8569,N_8296);
nand UO_153 (O_153,N_8254,N_9094);
nand UO_154 (O_154,N_9698,N_9192);
and UO_155 (O_155,N_8924,N_8729);
and UO_156 (O_156,N_8962,N_9749);
or UO_157 (O_157,N_9722,N_8381);
nand UO_158 (O_158,N_8062,N_8387);
nor UO_159 (O_159,N_9360,N_9160);
nand UO_160 (O_160,N_8024,N_9486);
or UO_161 (O_161,N_8582,N_8426);
or UO_162 (O_162,N_9526,N_8249);
nand UO_163 (O_163,N_8790,N_9603);
or UO_164 (O_164,N_9230,N_9813);
nor UO_165 (O_165,N_9771,N_8728);
nor UO_166 (O_166,N_8502,N_8655);
nand UO_167 (O_167,N_9128,N_9940);
or UO_168 (O_168,N_8274,N_8762);
and UO_169 (O_169,N_8197,N_9202);
nand UO_170 (O_170,N_8918,N_8753);
nor UO_171 (O_171,N_8077,N_8361);
nor UO_172 (O_172,N_8298,N_8975);
nor UO_173 (O_173,N_9154,N_8435);
nand UO_174 (O_174,N_9515,N_8823);
nand UO_175 (O_175,N_8236,N_8129);
and UO_176 (O_176,N_8146,N_8124);
nand UO_177 (O_177,N_9041,N_9901);
and UO_178 (O_178,N_9994,N_9710);
nor UO_179 (O_179,N_9186,N_9049);
nand UO_180 (O_180,N_9246,N_8626);
and UO_181 (O_181,N_8635,N_8903);
or UO_182 (O_182,N_8693,N_8817);
nor UO_183 (O_183,N_9695,N_8299);
nor UO_184 (O_184,N_9777,N_9502);
nor UO_185 (O_185,N_8628,N_8872);
or UO_186 (O_186,N_8007,N_8499);
or UO_187 (O_187,N_8204,N_8659);
nor UO_188 (O_188,N_8223,N_9481);
nand UO_189 (O_189,N_8476,N_8108);
nand UO_190 (O_190,N_8858,N_9511);
nor UO_191 (O_191,N_8712,N_8744);
xor UO_192 (O_192,N_9099,N_8644);
nor UO_193 (O_193,N_8253,N_9553);
or UO_194 (O_194,N_9421,N_8677);
nand UO_195 (O_195,N_8866,N_9605);
or UO_196 (O_196,N_8187,N_9768);
or UO_197 (O_197,N_9213,N_8267);
nor UO_198 (O_198,N_8897,N_8494);
nand UO_199 (O_199,N_9643,N_8778);
and UO_200 (O_200,N_9118,N_9419);
nor UO_201 (O_201,N_9003,N_8000);
and UO_202 (O_202,N_8763,N_8919);
nor UO_203 (O_203,N_9821,N_9137);
or UO_204 (O_204,N_8195,N_8189);
and UO_205 (O_205,N_8610,N_9320);
and UO_206 (O_206,N_8554,N_9221);
and UO_207 (O_207,N_9838,N_8354);
nand UO_208 (O_208,N_8831,N_8880);
nand UO_209 (O_209,N_9734,N_8676);
and UO_210 (O_210,N_8036,N_9536);
nand UO_211 (O_211,N_9895,N_9984);
or UO_212 (O_212,N_9073,N_8155);
or UO_213 (O_213,N_9516,N_8578);
nand UO_214 (O_214,N_9754,N_9046);
nor UO_215 (O_215,N_9310,N_8117);
nand UO_216 (O_216,N_9943,N_9374);
or UO_217 (O_217,N_8341,N_8263);
nand UO_218 (O_218,N_8969,N_9659);
nor UO_219 (O_219,N_9740,N_8539);
nand UO_220 (O_220,N_9070,N_8516);
nor UO_221 (O_221,N_8273,N_8691);
and UO_222 (O_222,N_9623,N_8248);
nand UO_223 (O_223,N_9136,N_8280);
or UO_224 (O_224,N_9244,N_8590);
and UO_225 (O_225,N_9119,N_8870);
nand UO_226 (O_226,N_9963,N_8226);
and UO_227 (O_227,N_8796,N_9074);
nor UO_228 (O_228,N_8115,N_9226);
nand UO_229 (O_229,N_8964,N_8735);
or UO_230 (O_230,N_8461,N_8225);
and UO_231 (O_231,N_8201,N_9638);
or UO_232 (O_232,N_9296,N_9784);
or UO_233 (O_233,N_8389,N_8902);
nand UO_234 (O_234,N_9831,N_8425);
nor UO_235 (O_235,N_9613,N_8867);
or UO_236 (O_236,N_9853,N_9305);
nor UO_237 (O_237,N_9197,N_8468);
nand UO_238 (O_238,N_8067,N_8622);
or UO_239 (O_239,N_8066,N_9842);
and UO_240 (O_240,N_8109,N_9278);
or UO_241 (O_241,N_9811,N_9716);
nor UO_242 (O_242,N_8297,N_9833);
nor UO_243 (O_243,N_9723,N_8807);
nand UO_244 (O_244,N_8528,N_8087);
or UO_245 (O_245,N_8379,N_8549);
and UO_246 (O_246,N_8261,N_9109);
and UO_247 (O_247,N_8312,N_9140);
or UO_248 (O_248,N_9508,N_9673);
and UO_249 (O_249,N_9489,N_9125);
nand UO_250 (O_250,N_9958,N_9799);
or UO_251 (O_251,N_9054,N_8544);
nand UO_252 (O_252,N_8636,N_8286);
or UO_253 (O_253,N_9103,N_9027);
nor UO_254 (O_254,N_9528,N_9250);
or UO_255 (O_255,N_8392,N_8180);
nand UO_256 (O_256,N_8250,N_8997);
nor UO_257 (O_257,N_9827,N_8181);
nand UO_258 (O_258,N_8947,N_8761);
and UO_259 (O_259,N_9730,N_8627);
nor UO_260 (O_260,N_9806,N_8716);
and UO_261 (O_261,N_8799,N_8151);
nor UO_262 (O_262,N_8134,N_9113);
nand UO_263 (O_263,N_9022,N_8832);
or UO_264 (O_264,N_9304,N_9960);
nor UO_265 (O_265,N_8471,N_9059);
or UO_266 (O_266,N_8084,N_8085);
and UO_267 (O_267,N_8642,N_9076);
or UO_268 (O_268,N_8216,N_8104);
or UO_269 (O_269,N_8491,N_9598);
or UO_270 (O_270,N_9973,N_8739);
nand UO_271 (O_271,N_9513,N_9222);
or UO_272 (O_272,N_8570,N_8656);
or UO_273 (O_273,N_8816,N_9530);
or UO_274 (O_274,N_9961,N_8961);
nand UO_275 (O_275,N_9259,N_9446);
or UO_276 (O_276,N_9665,N_9860);
or UO_277 (O_277,N_8019,N_9868);
or UO_278 (O_278,N_8160,N_8139);
nand UO_279 (O_279,N_9442,N_8908);
nand UO_280 (O_280,N_9590,N_8618);
and UO_281 (O_281,N_9656,N_8861);
nor UO_282 (O_282,N_9472,N_9229);
nor UO_283 (O_283,N_8527,N_8555);
nor UO_284 (O_284,N_8080,N_9286);
and UO_285 (O_285,N_9619,N_9276);
and UO_286 (O_286,N_8156,N_9008);
nor UO_287 (O_287,N_9448,N_9458);
nor UO_288 (O_288,N_8357,N_9930);
or UO_289 (O_289,N_9437,N_9275);
nor UO_290 (O_290,N_8305,N_9760);
nor UO_291 (O_291,N_9429,N_8498);
or UO_292 (O_292,N_9303,N_9517);
or UO_293 (O_293,N_9580,N_8999);
nand UO_294 (O_294,N_8076,N_8212);
or UO_295 (O_295,N_8682,N_9378);
or UO_296 (O_296,N_9630,N_8611);
nor UO_297 (O_297,N_8696,N_8633);
nand UO_298 (O_298,N_9725,N_9357);
nor UO_299 (O_299,N_9163,N_8152);
or UO_300 (O_300,N_9152,N_9162);
and UO_301 (O_301,N_9044,N_8821);
nand UO_302 (O_302,N_9443,N_8456);
or UO_303 (O_303,N_9322,N_9400);
nor UO_304 (O_304,N_9728,N_8992);
nand UO_305 (O_305,N_8690,N_9342);
xor UO_306 (O_306,N_8206,N_8012);
nor UO_307 (O_307,N_8172,N_8113);
nand UO_308 (O_308,N_8128,N_9832);
or UO_309 (O_309,N_9829,N_9424);
nand UO_310 (O_310,N_8891,N_9413);
or UO_311 (O_311,N_9300,N_9193);
nor UO_312 (O_312,N_9718,N_9887);
or UO_313 (O_313,N_8219,N_9942);
and UO_314 (O_314,N_8487,N_9185);
nor UO_315 (O_315,N_9713,N_9552);
or UO_316 (O_316,N_8607,N_8714);
nor UO_317 (O_317,N_9776,N_8447);
or UO_318 (O_318,N_8619,N_9212);
and UO_319 (O_319,N_9686,N_8470);
nand UO_320 (O_320,N_8830,N_8132);
nor UO_321 (O_321,N_9431,N_9941);
and UO_322 (O_322,N_8629,N_9565);
nand UO_323 (O_323,N_9157,N_8538);
or UO_324 (O_324,N_8493,N_9441);
or UO_325 (O_325,N_8342,N_9820);
nor UO_326 (O_326,N_9248,N_8373);
nor UO_327 (O_327,N_9945,N_9529);
and UO_328 (O_328,N_8140,N_8247);
nor UO_329 (O_329,N_9846,N_9289);
nor UO_330 (O_330,N_8339,N_8162);
nand UO_331 (O_331,N_8787,N_8721);
nor UO_332 (O_332,N_8333,N_8779);
nand UO_333 (O_333,N_8021,N_8806);
or UO_334 (O_334,N_8856,N_8285);
nand UO_335 (O_335,N_9753,N_8514);
or UO_336 (O_336,N_8311,N_9618);
or UO_337 (O_337,N_9258,N_8414);
and UO_338 (O_338,N_9977,N_8706);
or UO_339 (O_339,N_9633,N_9913);
nand UO_340 (O_340,N_8370,N_9280);
nor UO_341 (O_341,N_8631,N_9959);
or UO_342 (O_342,N_9260,N_8736);
nor UO_343 (O_343,N_8412,N_9194);
and UO_344 (O_344,N_9661,N_8458);
nor UO_345 (O_345,N_9081,N_9592);
or UO_346 (O_346,N_8005,N_9916);
nand UO_347 (O_347,N_9112,N_8397);
nand UO_348 (O_348,N_9921,N_8829);
nand UO_349 (O_349,N_9571,N_9225);
nor UO_350 (O_350,N_9711,N_9792);
and UO_351 (O_351,N_9889,N_8568);
nor UO_352 (O_352,N_9483,N_8959);
and UO_353 (O_353,N_8865,N_8266);
and UO_354 (O_354,N_8725,N_8142);
or UO_355 (O_355,N_8409,N_9679);
or UO_356 (O_356,N_8824,N_9938);
or UO_357 (O_357,N_8243,N_9602);
and UO_358 (O_358,N_9087,N_8413);
nand UO_359 (O_359,N_9683,N_9825);
nor UO_360 (O_360,N_9292,N_9245);
nand UO_361 (O_361,N_9601,N_8754);
nand UO_362 (O_362,N_8625,N_8068);
nor UO_363 (O_363,N_9903,N_8808);
nor UO_364 (O_364,N_8641,N_8454);
nor UO_365 (O_365,N_8390,N_8334);
or UO_366 (O_366,N_8233,N_9747);
nor UO_367 (O_367,N_9761,N_9624);
nand UO_368 (O_368,N_9082,N_9384);
or UO_369 (O_369,N_9816,N_9461);
nor UO_370 (O_370,N_9161,N_8848);
and UO_371 (O_371,N_8937,N_9692);
xnor UO_372 (O_372,N_8987,N_8887);
nand UO_373 (O_373,N_9557,N_8377);
nand UO_374 (O_374,N_8921,N_8580);
or UO_375 (O_375,N_8681,N_8765);
nor UO_376 (O_376,N_9023,N_9983);
nand UO_377 (O_377,N_9875,N_9884);
and UO_378 (O_378,N_9001,N_8427);
or UO_379 (O_379,N_9257,N_8174);
nand UO_380 (O_380,N_9040,N_8860);
nor UO_381 (O_381,N_8820,N_8320);
and UO_382 (O_382,N_9700,N_9650);
and UO_383 (O_383,N_8394,N_9585);
nand UO_384 (O_384,N_9535,N_9882);
nand UO_385 (O_385,N_9341,N_8455);
and UO_386 (O_386,N_9372,N_9336);
or UO_387 (O_387,N_9642,N_8375);
or UO_388 (O_388,N_8939,N_9697);
and UO_389 (O_389,N_9107,N_9385);
or UO_390 (O_390,N_8781,N_9358);
nand UO_391 (O_391,N_9607,N_9703);
and UO_392 (O_392,N_9018,N_8605);
nor UO_393 (O_393,N_9586,N_8045);
and UO_394 (O_394,N_9348,N_8178);
nand UO_395 (O_395,N_8446,N_8071);
nor UO_396 (O_396,N_8363,N_9670);
or UO_397 (O_397,N_8202,N_8620);
nand UO_398 (O_398,N_8873,N_8825);
and UO_399 (O_399,N_8805,N_8023);
nand UO_400 (O_400,N_9450,N_9048);
nor UO_401 (O_401,N_8899,N_9892);
nor UO_402 (O_402,N_8958,N_8733);
nor UO_403 (O_403,N_8742,N_8402);
or UO_404 (O_404,N_8445,N_9379);
nand UO_405 (O_405,N_9735,N_9951);
and UO_406 (O_406,N_8657,N_9786);
or UO_407 (O_407,N_9655,N_9864);
nor UO_408 (O_408,N_9325,N_9017);
or UO_409 (O_409,N_8100,N_9386);
and UO_410 (O_410,N_9433,N_8575);
and UO_411 (O_411,N_8048,N_8671);
nor UO_412 (O_412,N_8367,N_9038);
and UO_413 (O_413,N_8399,N_9012);
xnor UO_414 (O_414,N_9815,N_8214);
nand UO_415 (O_415,N_9299,N_8475);
or UO_416 (O_416,N_8176,N_8405);
and UO_417 (O_417,N_9854,N_9425);
and UO_418 (O_418,N_8073,N_9396);
or UO_419 (O_419,N_8551,N_8283);
nor UO_420 (O_420,N_9037,N_8416);
or UO_421 (O_421,N_8359,N_9351);
or UO_422 (O_422,N_9615,N_8864);
nor UO_423 (O_423,N_8705,N_9402);
nor UO_424 (O_424,N_9803,N_8331);
nor UO_425 (O_425,N_9759,N_8244);
or UO_426 (O_426,N_9802,N_8535);
nand UO_427 (O_427,N_9151,N_8859);
or UO_428 (O_428,N_8842,N_9079);
or UO_429 (O_429,N_9177,N_8708);
or UO_430 (O_430,N_8685,N_9026);
or UO_431 (O_431,N_9724,N_8384);
or UO_432 (O_432,N_9849,N_8508);
xnor UO_433 (O_433,N_8246,N_9239);
nor UO_434 (O_434,N_9664,N_8759);
nand UO_435 (O_435,N_8043,N_9191);
nor UO_436 (O_436,N_8511,N_8663);
or UO_437 (O_437,N_9269,N_9494);
xnor UO_438 (O_438,N_8558,N_8900);
or UO_439 (O_439,N_9416,N_8252);
nand UO_440 (O_440,N_9476,N_8022);
or UO_441 (O_441,N_9736,N_9687);
or UO_442 (O_442,N_9741,N_9016);
and UO_443 (O_443,N_8871,N_8515);
and UO_444 (O_444,N_8788,N_9947);
and UO_445 (O_445,N_9523,N_9254);
and UO_446 (O_446,N_8205,N_9264);
nor UO_447 (O_447,N_9126,N_8700);
or UO_448 (O_448,N_8586,N_8772);
and UO_449 (O_449,N_9847,N_8540);
and UO_450 (O_450,N_9218,N_9293);
or UO_451 (O_451,N_8815,N_9312);
nand UO_452 (O_452,N_9268,N_8083);
or UO_453 (O_453,N_8944,N_8980);
nor UO_454 (O_454,N_8457,N_8188);
nor UO_455 (O_455,N_9966,N_9355);
nand UO_456 (O_456,N_8495,N_8271);
nor UO_457 (O_457,N_9319,N_9387);
and UO_458 (O_458,N_8561,N_8979);
nand UO_459 (O_459,N_8208,N_8421);
nor UO_460 (O_460,N_9690,N_8228);
nand UO_461 (O_461,N_9653,N_8269);
and UO_462 (O_462,N_9540,N_8161);
or UO_463 (O_463,N_9787,N_8089);
nor UO_464 (O_464,N_9600,N_9509);
nor UO_465 (O_465,N_9078,N_9701);
or UO_466 (O_466,N_9065,N_8519);
nand UO_467 (O_467,N_8369,N_9620);
xor UO_468 (O_468,N_9328,N_9043);
nor UO_469 (O_469,N_9183,N_9702);
or UO_470 (O_470,N_9284,N_8415);
and UO_471 (O_471,N_8175,N_8719);
nor UO_472 (O_472,N_8675,N_9231);
and UO_473 (O_473,N_9965,N_8168);
nor UO_474 (O_474,N_9594,N_9685);
nand UO_475 (O_475,N_8091,N_8207);
nand UO_476 (O_476,N_8492,N_9009);
or UO_477 (O_477,N_9333,N_9243);
nor UO_478 (O_478,N_9912,N_9971);
or UO_479 (O_479,N_9869,N_9365);
or UO_480 (O_480,N_8120,N_9148);
nand UO_481 (O_481,N_9576,N_9808);
nor UO_482 (O_482,N_8660,N_8801);
nor UO_483 (O_483,N_8965,N_9477);
and UO_484 (O_484,N_8653,N_8709);
or UO_485 (O_485,N_8337,N_9343);
or UO_486 (O_486,N_8098,N_9500);
nor UO_487 (O_487,N_8075,N_9233);
nor UO_488 (O_488,N_9651,N_9345);
or UO_489 (O_489,N_8661,N_9302);
nand UO_490 (O_490,N_9793,N_9069);
nor UO_491 (O_491,N_9781,N_9436);
and UO_492 (O_492,N_9840,N_9691);
nand UO_493 (O_493,N_9967,N_8533);
nand UO_494 (O_494,N_8760,N_8722);
nor UO_495 (O_495,N_8069,N_8093);
nor UO_496 (O_496,N_9287,N_8224);
nor UO_497 (O_497,N_8326,N_8512);
or UO_498 (O_498,N_9902,N_9393);
and UO_499 (O_499,N_9473,N_8623);
nor UO_500 (O_500,N_8526,N_9823);
or UO_501 (O_501,N_9149,N_8797);
or UO_502 (O_502,N_9612,N_9743);
or UO_503 (O_503,N_9775,N_8988);
nor UO_504 (O_504,N_9055,N_9169);
and UO_505 (O_505,N_8974,N_8404);
or UO_506 (O_506,N_8095,N_9885);
nor UO_507 (O_507,N_9294,N_8782);
nand UO_508 (O_508,N_9228,N_8666);
and UO_509 (O_509,N_9588,N_8665);
and UO_510 (O_510,N_9392,N_8396);
and UO_511 (O_511,N_9750,N_8819);
nor UO_512 (O_512,N_9634,N_9497);
xor UO_513 (O_513,N_8550,N_8251);
or UO_514 (O_514,N_8268,N_8530);
or UO_515 (O_515,N_8751,N_8791);
nor UO_516 (O_516,N_9795,N_8562);
nor UO_517 (O_517,N_9262,N_9621);
nand UO_518 (O_518,N_9417,N_8645);
nand UO_519 (O_519,N_9852,N_8008);
nor UO_520 (O_520,N_8563,N_8658);
and UO_521 (O_521,N_8448,N_9184);
or UO_522 (O_522,N_9558,N_9818);
nand UO_523 (O_523,N_8640,N_9841);
nand UO_524 (O_524,N_9203,N_8319);
and UO_525 (O_525,N_8374,N_8191);
nor UO_526 (O_526,N_8488,N_9689);
or UO_527 (O_527,N_8131,N_9814);
or UO_528 (O_528,N_8040,N_9654);
or UO_529 (O_529,N_8809,N_8324);
nor UO_530 (O_530,N_9871,N_9110);
or UO_531 (O_531,N_9524,N_8603);
nor UO_532 (O_532,N_9648,N_8949);
nor UO_533 (O_533,N_9726,N_8330);
nor UO_534 (O_534,N_8884,N_9227);
or UO_535 (O_535,N_9617,N_9321);
nand UO_536 (O_536,N_9627,N_9979);
and UO_537 (O_537,N_9200,N_8262);
nor UO_538 (O_538,N_9139,N_9096);
nand UO_539 (O_539,N_8850,N_8452);
nor UO_540 (O_540,N_8945,N_8698);
nor UO_541 (O_541,N_9986,N_8732);
nor UO_542 (O_542,N_8275,N_8501);
nand UO_543 (O_543,N_8929,N_9757);
nor UO_544 (O_544,N_8288,N_8745);
nand UO_545 (O_545,N_9779,N_8099);
nand UO_546 (O_546,N_9699,N_8479);
nor UO_547 (O_547,N_8686,N_9120);
nand UO_548 (O_548,N_8014,N_9188);
and UO_549 (O_549,N_9872,N_9804);
and UO_550 (O_550,N_9178,N_9990);
nor UO_551 (O_551,N_9835,N_9505);
or UO_552 (O_552,N_8651,N_8922);
or UO_553 (O_553,N_9209,N_8450);
nand UO_554 (O_554,N_9032,N_9207);
nand UO_555 (O_555,N_8740,N_9405);
and UO_556 (O_556,N_8652,N_9145);
and UO_557 (O_557,N_9998,N_8837);
nor UO_558 (O_558,N_9098,N_9547);
nand UO_559 (O_559,N_9144,N_9807);
nor UO_560 (O_560,N_9863,N_9861);
or UO_561 (O_561,N_9937,N_9527);
nand UO_562 (O_562,N_9791,N_8046);
nand UO_563 (O_563,N_9954,N_8993);
or UO_564 (O_564,N_8981,N_9646);
and UO_565 (O_565,N_9671,N_8473);
nor UO_566 (O_566,N_8704,N_9931);
or UO_567 (O_567,N_9471,N_8345);
nor UO_568 (O_568,N_8847,N_9391);
and UO_569 (O_569,N_8777,N_9095);
nand UO_570 (O_570,N_8125,N_9812);
nor UO_571 (O_571,N_8441,N_8844);
or UO_572 (O_572,N_8697,N_9168);
and UO_573 (O_573,N_8798,N_8976);
nor UO_574 (O_574,N_8481,N_8378);
and UO_575 (O_575,N_9408,N_9438);
or UO_576 (O_576,N_9492,N_9684);
nor UO_577 (O_577,N_8054,N_9729);
and UO_578 (O_578,N_8094,N_8503);
nor UO_579 (O_579,N_8074,N_9932);
nor UO_580 (O_580,N_9147,N_8954);
or UO_581 (O_581,N_9062,N_9746);
nand UO_582 (O_582,N_9367,N_8741);
nor UO_583 (O_583,N_8235,N_8116);
or UO_584 (O_584,N_9506,N_9307);
and UO_585 (O_585,N_9427,N_8453);
nand UO_586 (O_586,N_9397,N_9326);
nand UO_587 (O_587,N_8804,N_9411);
nor UO_588 (O_588,N_9196,N_8123);
nor UO_589 (O_589,N_8523,N_9339);
nand UO_590 (O_590,N_9800,N_9964);
nand UO_591 (O_591,N_8785,N_8096);
nand UO_592 (O_592,N_8909,N_8795);
and UO_593 (O_593,N_8483,N_9676);
or UO_594 (O_594,N_8936,N_8525);
and UO_595 (O_595,N_8757,N_9315);
or UO_596 (O_596,N_8869,N_9072);
and UO_597 (O_597,N_9538,N_9491);
nand UO_598 (O_598,N_9204,N_8422);
or UO_599 (O_599,N_8018,N_8049);
or UO_600 (O_600,N_8940,N_9675);
nor UO_601 (O_601,N_9071,N_8393);
nand UO_602 (O_602,N_8755,N_9171);
nor UO_603 (O_603,N_9962,N_8282);
nor UO_604 (O_604,N_9064,N_8451);
nor UO_605 (O_605,N_8227,N_8338);
nor UO_606 (O_606,N_8726,N_8507);
nand UO_607 (O_607,N_9910,N_9116);
nand UO_608 (O_608,N_8010,N_9609);
nor UO_609 (O_609,N_9790,N_9696);
nand UO_610 (O_610,N_9460,N_8892);
nor UO_611 (O_611,N_8482,N_8560);
nor UO_612 (O_612,N_8792,N_9608);
and UO_613 (O_613,N_9463,N_8027);
or UO_614 (O_614,N_9208,N_9789);
or UO_615 (O_615,N_8730,N_9249);
nor UO_616 (O_616,N_9668,N_9383);
nand UO_617 (O_617,N_8213,N_8443);
nand UO_618 (O_618,N_9390,N_9242);
or UO_619 (O_619,N_8906,N_8177);
or UO_620 (O_620,N_8474,N_8410);
nor UO_621 (O_621,N_8839,N_8835);
and UO_622 (O_622,N_9011,N_9007);
nand UO_623 (O_623,N_9394,N_8065);
or UO_624 (O_624,N_8362,N_8614);
xnor UO_625 (O_625,N_8770,N_9369);
and UO_626 (O_626,N_9568,N_8307);
nand UO_627 (O_627,N_9042,N_9974);
nor UO_628 (O_628,N_8715,N_8649);
or UO_629 (O_629,N_9644,N_9677);
nand UO_630 (O_630,N_8294,N_9751);
nand UO_631 (O_631,N_9021,N_8231);
nor UO_632 (O_632,N_9133,N_8032);
nand UO_633 (O_633,N_8654,N_9904);
or UO_634 (O_634,N_8703,N_8034);
or UO_635 (O_635,N_9143,N_9263);
nor UO_636 (O_636,N_8688,N_9318);
nor UO_637 (O_637,N_9923,N_8592);
nand UO_638 (O_638,N_8200,N_9122);
nand UO_639 (O_639,N_9058,N_9891);
nor UO_640 (O_640,N_8332,N_8170);
nand UO_641 (O_641,N_8105,N_8052);
and UO_642 (O_642,N_9414,N_8127);
nand UO_643 (O_643,N_9025,N_8524);
nand UO_644 (O_644,N_8148,N_8364);
or UO_645 (O_645,N_8439,N_8926);
or UO_646 (O_646,N_8149,N_9175);
nor UO_647 (O_647,N_9334,N_8583);
and UO_648 (O_648,N_8190,N_8624);
nand UO_649 (O_649,N_8020,N_9794);
nand UO_650 (O_650,N_9674,N_8692);
or UO_651 (O_651,N_9067,N_8667);
or UO_652 (O_652,N_8122,N_9189);
or UO_653 (O_653,N_8600,N_8843);
nand UO_654 (O_654,N_9652,N_9454);
nor UO_655 (O_655,N_9444,N_9909);
nor UO_656 (O_656,N_8238,N_9308);
or UO_657 (O_657,N_9206,N_8559);
nand UO_658 (O_658,N_8221,N_8291);
nand UO_659 (O_659,N_9739,N_8376);
and UO_660 (O_660,N_8346,N_8395);
xor UO_661 (O_661,N_8702,N_8531);
nand UO_662 (O_662,N_9216,N_9997);
or UO_663 (O_663,N_8890,N_8599);
and UO_664 (O_664,N_8584,N_8984);
or UO_665 (O_665,N_8029,N_8811);
nand UO_666 (O_666,N_8086,N_8313);
nand UO_667 (O_667,N_9667,N_9758);
nand UO_668 (O_668,N_8838,N_9174);
nand UO_669 (O_669,N_9637,N_8604);
nor UO_670 (O_670,N_8593,N_9976);
xor UO_671 (O_671,N_8934,N_9434);
or UO_672 (O_672,N_8002,N_9970);
or UO_673 (O_673,N_9298,N_9551);
or UO_674 (O_674,N_8462,N_9261);
nor UO_675 (O_675,N_8914,N_9337);
nor UO_676 (O_676,N_9935,N_8879);
nor UO_677 (O_677,N_9004,N_9499);
or UO_678 (O_678,N_8430,N_8978);
or UO_679 (O_679,N_9830,N_8731);
and UO_680 (O_680,N_8943,N_9217);
or UO_681 (O_681,N_8106,N_9091);
nand UO_682 (O_682,N_9503,N_9187);
nand UO_683 (O_683,N_9115,N_8001);
or UO_684 (O_684,N_8646,N_9456);
and UO_685 (O_685,N_8215,N_8329);
nand UO_686 (O_686,N_9093,N_8775);
and UO_687 (O_687,N_8747,N_9015);
and UO_688 (O_688,N_9819,N_8143);
nand UO_689 (O_689,N_8564,N_8111);
nor UO_690 (O_690,N_9987,N_9475);
and UO_691 (O_691,N_9415,N_8950);
nand UO_692 (O_692,N_9346,N_9000);
nor UO_693 (O_693,N_8466,N_8678);
and UO_694 (O_694,N_8948,N_8989);
and UO_695 (O_695,N_9409,N_9404);
nand UO_696 (O_696,N_8707,N_8391);
nor UO_697 (O_697,N_9645,N_9595);
nor UO_698 (O_698,N_9256,N_8800);
and UO_699 (O_699,N_9088,N_9335);
or UO_700 (O_700,N_8794,N_9647);
and UO_701 (O_701,N_9395,N_9949);
nor UO_702 (O_702,N_8472,N_8968);
or UO_703 (O_703,N_8343,N_8290);
or UO_704 (O_704,N_8510,N_9593);
nor UO_705 (O_705,N_8672,N_8436);
and UO_706 (O_706,N_9610,N_8467);
or UO_707 (O_707,N_9550,N_9451);
or UO_708 (O_708,N_8841,N_8574);
or UO_709 (O_709,N_9999,N_8786);
and UO_710 (O_710,N_9406,N_9297);
nor UO_711 (O_711,N_9090,N_8289);
or UO_712 (O_712,N_9767,N_9495);
nand UO_713 (O_713,N_8292,N_9897);
nand UO_714 (O_714,N_9543,N_8220);
xor UO_715 (O_715,N_8556,N_9635);
and UO_716 (O_716,N_9544,N_9182);
or UO_717 (O_717,N_9563,N_9085);
nor UO_718 (O_718,N_8110,N_9525);
and UO_719 (O_719,N_8576,N_9549);
or UO_720 (O_720,N_8169,N_9579);
and UO_721 (O_721,N_9780,N_8695);
and UO_722 (O_722,N_9837,N_9944);
nor UO_723 (O_723,N_8571,N_9744);
xnor UO_724 (O_724,N_9291,N_9533);
and UO_725 (O_725,N_8917,N_8840);
and UO_726 (O_726,N_9376,N_9327);
nand UO_727 (O_727,N_9762,N_9344);
nor UO_728 (O_728,N_9672,N_9927);
nand UO_729 (O_729,N_8673,N_8711);
nor UO_730 (O_730,N_8895,N_9641);
nor UO_731 (O_731,N_8193,N_9569);
and UO_732 (O_732,N_9554,N_8985);
and UO_733 (O_733,N_9824,N_8070);
nor UO_734 (O_734,N_9519,N_8534);
and UO_735 (O_735,N_9714,N_9150);
nand UO_736 (O_736,N_9573,N_8259);
nand UO_737 (O_737,N_8318,N_8602);
and UO_738 (O_738,N_9083,N_9423);
nand UO_739 (O_739,N_9577,N_8601);
or UO_740 (O_740,N_8723,N_8496);
or UO_741 (O_741,N_8147,N_9510);
or UO_742 (O_742,N_9100,N_9359);
or UO_743 (O_743,N_9108,N_9953);
nand UO_744 (O_744,N_9165,N_8303);
and UO_745 (O_745,N_9873,N_8088);
nor UO_746 (O_746,N_8293,N_8042);
nor UO_747 (O_747,N_8063,N_8552);
and UO_748 (O_748,N_9769,N_8766);
nor UO_749 (O_749,N_9317,N_8854);
or UO_750 (O_750,N_8203,N_9870);
and UO_751 (O_751,N_8529,N_8047);
nand UO_752 (O_752,N_8670,N_8165);
nand UO_753 (O_753,N_9720,N_9199);
and UO_754 (O_754,N_9487,N_9465);
xor UO_755 (O_755,N_8738,N_8542);
nor UO_756 (O_756,N_8017,N_9399);
xor UO_757 (O_757,N_8081,N_9878);
nor UO_758 (O_758,N_9117,N_9606);
nor UO_759 (O_759,N_9445,N_9316);
or UO_760 (O_760,N_9649,N_8260);
nor UO_761 (O_761,N_9541,N_8323);
nand UO_762 (O_762,N_8103,N_8428);
nand UO_763 (O_763,N_9271,N_9715);
and UO_764 (O_764,N_8912,N_8863);
nor UO_765 (O_765,N_8064,N_8910);
nand UO_766 (O_766,N_9490,N_9559);
nor UO_767 (O_767,N_8970,N_8039);
or UO_768 (O_768,N_9862,N_9975);
nand UO_769 (O_769,N_9596,N_8828);
and UO_770 (O_770,N_9052,N_8881);
nand UO_771 (O_771,N_8411,N_9420);
nor UO_772 (O_772,N_9857,N_9981);
and UO_773 (O_773,N_8015,N_8694);
or UO_774 (O_774,N_8783,N_9548);
or UO_775 (O_775,N_9449,N_9164);
nand UO_776 (O_776,N_9179,N_8668);
nand UO_777 (O_777,N_9353,N_9002);
and UO_778 (O_778,N_9874,N_9364);
nor UO_779 (O_779,N_9238,N_8713);
nand UO_780 (O_780,N_8925,N_8768);
or UO_781 (O_781,N_8893,N_8497);
or UO_782 (O_782,N_8746,N_8643);
nand UO_783 (O_783,N_9855,N_8938);
xor UO_784 (O_784,N_9075,N_9288);
and UO_785 (O_785,N_8486,N_9658);
nand UO_786 (O_786,N_9265,N_8060);
and UO_787 (O_787,N_9466,N_8465);
or UO_788 (O_788,N_9050,N_8403);
or UO_789 (O_789,N_9266,N_9057);
nor UO_790 (O_790,N_8935,N_8097);
and UO_791 (O_791,N_8960,N_9985);
and UO_792 (O_792,N_9045,N_8505);
or UO_793 (O_793,N_8774,N_9917);
and UO_794 (O_794,N_8637,N_8683);
and UO_795 (O_795,N_8933,N_8464);
or UO_796 (O_796,N_9373,N_8930);
and UO_797 (O_797,N_9097,N_8350);
and UO_798 (O_798,N_8079,N_9123);
and UO_799 (O_799,N_9721,N_8270);
nor UO_800 (O_800,N_9370,N_9480);
or UO_801 (O_801,N_8973,N_8737);
nand UO_802 (O_802,N_9468,N_8664);
or UO_803 (O_803,N_8905,N_8258);
nand UO_804 (O_804,N_8406,N_8536);
or UO_805 (O_805,N_9132,N_9240);
nor UO_806 (O_806,N_8130,N_8833);
or UO_807 (O_807,N_8222,N_9531);
or UO_808 (O_808,N_8030,N_8164);
nor UO_809 (O_809,N_8366,N_9707);
nand UO_810 (O_810,N_8490,N_8932);
and UO_811 (O_811,N_8353,N_8418);
or UO_812 (O_812,N_8752,N_8126);
or UO_813 (O_813,N_9989,N_9534);
and UO_814 (O_814,N_8990,N_9866);
and UO_815 (O_815,N_9764,N_9455);
nor UO_816 (O_816,N_8638,N_8322);
nand UO_817 (O_817,N_9114,N_9507);
nand UO_818 (O_818,N_8579,N_9381);
or UO_819 (O_819,N_8596,N_9347);
and UO_820 (O_820,N_9587,N_9277);
nand UO_821 (O_821,N_9432,N_8237);
nor UO_822 (O_822,N_8004,N_9352);
nor UO_823 (O_823,N_8356,N_8615);
nor UO_824 (O_824,N_9241,N_8157);
xnor UO_825 (O_825,N_9582,N_8898);
or UO_826 (O_826,N_9282,N_9056);
or UO_827 (O_827,N_8351,N_8035);
nand UO_828 (O_828,N_9219,N_9127);
nor UO_829 (O_829,N_8920,N_8198);
and UO_830 (O_830,N_8836,N_8344);
or UO_831 (O_831,N_8217,N_9102);
or UO_832 (O_832,N_9900,N_8591);
or UO_833 (O_833,N_8184,N_9848);
and UO_834 (O_834,N_9639,N_9398);
and UO_835 (O_835,N_9464,N_8720);
nor UO_836 (O_836,N_8317,N_8194);
or UO_837 (O_837,N_8894,N_9636);
and UO_838 (O_838,N_8171,N_9361);
nand UO_839 (O_839,N_9748,N_9324);
nor UO_840 (O_840,N_9439,N_8504);
nor UO_841 (O_841,N_9104,N_8287);
and UO_842 (O_842,N_9130,N_8882);
nand UO_843 (O_843,N_9957,N_8857);
or UO_844 (O_844,N_9614,N_9135);
nand UO_845 (O_845,N_9349,N_9388);
and UO_846 (O_846,N_8598,N_9426);
and UO_847 (O_847,N_8613,N_9678);
or UO_848 (O_848,N_8545,N_8437);
nand UO_849 (O_849,N_9922,N_9350);
nand UO_850 (O_850,N_9330,N_9462);
or UO_851 (O_851,N_8577,N_8810);
nor UO_852 (O_852,N_8061,N_8423);
nor UO_853 (O_853,N_8460,N_9338);
nand UO_854 (O_854,N_8484,N_9542);
or UO_855 (O_855,N_8971,N_8886);
or UO_856 (O_856,N_8383,N_8368);
nor UO_857 (O_857,N_9532,N_8444);
and UO_858 (O_858,N_8822,N_8121);
nor UO_859 (O_859,N_8431,N_8982);
nor UO_860 (O_860,N_8717,N_9939);
and UO_861 (O_861,N_8281,N_8557);
nand UO_862 (O_862,N_9604,N_8994);
nand UO_863 (O_863,N_9251,N_8888);
or UO_864 (O_864,N_9493,N_9660);
and UO_865 (O_865,N_9331,N_8532);
and UO_866 (O_866,N_8382,N_9752);
and UO_867 (O_867,N_9129,N_9323);
or UO_868 (O_868,N_9626,N_8209);
nand UO_869 (O_869,N_8506,N_8316);
nand UO_870 (O_870,N_8885,N_9080);
and UO_871 (O_871,N_9893,N_8141);
nor UO_872 (O_872,N_8597,N_9628);
nand UO_873 (O_873,N_9996,N_9801);
nand UO_874 (O_874,N_9514,N_8734);
or UO_875 (O_875,N_8845,N_9520);
and UO_876 (O_876,N_8710,N_8901);
and UO_877 (O_877,N_9828,N_9283);
nor UO_878 (O_878,N_8092,N_8951);
nor UO_879 (O_879,N_9755,N_9410);
or UO_880 (O_880,N_8102,N_8566);
nor UO_881 (O_881,N_8749,N_9181);
and UO_882 (O_882,N_8398,N_9340);
nand UO_883 (O_883,N_9680,N_8348);
or UO_884 (O_884,N_8758,N_9742);
or UO_885 (O_885,N_8044,N_9995);
nor UO_886 (O_886,N_8082,N_8818);
nor UO_887 (O_887,N_9035,N_9031);
and UO_888 (O_888,N_9060,N_9172);
xor UO_889 (O_889,N_8401,N_8878);
and UO_890 (O_890,N_9170,N_8996);
nor UO_891 (O_891,N_8621,N_8883);
nand UO_892 (O_892,N_8434,N_9274);
or UO_893 (O_893,N_9737,N_8442);
and UO_894 (O_894,N_8196,N_9657);
or UO_895 (O_895,N_8264,N_9356);
and UO_896 (O_896,N_8724,N_8058);
nand UO_897 (O_897,N_9629,N_8616);
nor UO_898 (O_898,N_9969,N_8877);
or UO_899 (O_899,N_8349,N_8163);
and UO_900 (O_900,N_9496,N_9856);
xnor UO_901 (O_901,N_9844,N_8485);
or UO_902 (O_902,N_9783,N_8013);
nor UO_903 (O_903,N_9329,N_8380);
or UO_904 (O_904,N_8031,N_8173);
nand UO_905 (O_905,N_9138,N_9270);
or UO_906 (O_906,N_9798,N_8648);
nand UO_907 (O_907,N_8814,N_9235);
nand UO_908 (O_908,N_8321,N_9156);
and UO_909 (O_909,N_9858,N_8041);
or UO_910 (O_910,N_8420,N_9899);
or UO_911 (O_911,N_9467,N_9918);
or UO_912 (O_912,N_9210,N_9167);
nand UO_913 (O_913,N_9141,N_9309);
nor UO_914 (O_914,N_9105,N_9570);
or UO_915 (O_915,N_8647,N_9881);
or UO_916 (O_916,N_8802,N_9279);
nand UO_917 (O_917,N_9028,N_9430);
nor UO_918 (O_918,N_9237,N_8167);
nor UO_919 (O_919,N_8500,N_8277);
nor UO_920 (O_920,N_9915,N_8963);
nor UO_921 (O_921,N_9086,N_8846);
or UO_922 (O_922,N_8278,N_8567);
nor UO_923 (O_923,N_8279,N_9980);
or UO_924 (O_924,N_8242,N_9583);
nand UO_925 (O_925,N_8459,N_8803);
nand UO_926 (O_926,N_9928,N_8928);
nor UO_927 (O_927,N_9914,N_9850);
nand UO_928 (O_928,N_8059,N_8417);
or UO_929 (O_929,N_9936,N_8145);
and UO_930 (O_930,N_9555,N_8328);
nand UO_931 (O_931,N_9666,N_9708);
nor UO_932 (O_932,N_9663,N_8679);
and UO_933 (O_933,N_9422,N_9368);
or UO_934 (O_934,N_9717,N_9988);
or UO_935 (O_935,N_9281,N_8983);
nor UO_936 (O_936,N_9625,N_9521);
or UO_937 (O_937,N_8767,N_9836);
nor UO_938 (O_938,N_8433,N_9925);
or UO_939 (O_939,N_8239,N_8634);
nor UO_940 (O_940,N_9562,N_8360);
and UO_941 (O_941,N_8521,N_8769);
or UO_942 (O_942,N_9785,N_8977);
nor UO_943 (O_943,N_9578,N_9705);
nor UO_944 (O_944,N_9732,N_9403);
nor UO_945 (O_945,N_8003,N_8053);
or UO_946 (O_946,N_9314,N_9992);
and UO_947 (O_947,N_9006,N_9591);
and UO_948 (O_948,N_9843,N_9014);
or UO_949 (O_949,N_9068,N_8851);
and UO_950 (O_950,N_9092,N_8315);
and UO_951 (O_951,N_8025,N_8998);
or UO_952 (O_952,N_9756,N_8218);
nor UO_953 (O_953,N_9640,N_9313);
or UO_954 (O_954,N_9155,N_9616);
nand UO_955 (O_955,N_8055,N_8440);
nand UO_956 (O_956,N_8907,N_9478);
nor UO_957 (O_957,N_9731,N_8972);
and UO_958 (O_958,N_8585,N_8573);
and UO_959 (O_959,N_8150,N_9908);
nand UO_960 (O_960,N_8727,N_8051);
nor UO_961 (O_961,N_8771,N_8608);
nor UO_962 (O_962,N_9978,N_8617);
nand UO_963 (O_963,N_8513,N_9763);
nor UO_964 (O_964,N_9362,N_8957);
nand UO_965 (O_965,N_8595,N_9077);
nor UO_966 (O_966,N_9952,N_8144);
nor UO_967 (O_967,N_9005,N_9905);
nor UO_968 (O_968,N_9030,N_8489);
nand UO_969 (O_969,N_8211,N_9255);
or UO_970 (O_970,N_8199,N_8136);
nand UO_971 (O_971,N_9946,N_9101);
nand UO_972 (O_972,N_9176,N_8565);
or UO_973 (O_973,N_9631,N_9575);
nand UO_974 (O_974,N_8915,N_8388);
nor UO_975 (O_975,N_9539,N_8855);
or UO_976 (O_976,N_9817,N_9982);
and UO_977 (O_977,N_9121,N_8630);
or UO_978 (O_978,N_9371,N_9883);
and UO_979 (O_979,N_8119,N_8325);
and UO_980 (O_980,N_9738,N_8756);
and UO_981 (O_981,N_9546,N_8371);
or UO_982 (O_982,N_8639,N_9457);
nand UO_983 (O_983,N_8684,N_9890);
and UO_984 (O_984,N_9772,N_9440);
and UO_985 (O_985,N_8650,N_9377);
and UO_986 (O_986,N_9452,N_8689);
nor UO_987 (O_987,N_8230,N_9047);
nor UO_988 (O_988,N_8304,N_8904);
nand UO_989 (O_989,N_9211,N_9036);
or UO_990 (O_990,N_9380,N_8718);
and UO_991 (O_991,N_9382,N_9479);
and UO_992 (O_992,N_9681,N_9694);
nand UO_993 (O_993,N_8090,N_8480);
nand UO_994 (O_994,N_9290,N_8853);
nand UO_995 (O_995,N_9688,N_9504);
or UO_996 (O_996,N_8408,N_9765);
and UO_997 (O_997,N_9389,N_8827);
nand UO_998 (O_998,N_9876,N_8955);
or UO_999 (O_999,N_8952,N_8946);
nand UO_1000 (O_1000,N_9022,N_9649);
or UO_1001 (O_1001,N_8522,N_8957);
nor UO_1002 (O_1002,N_9517,N_8559);
or UO_1003 (O_1003,N_8101,N_9722);
or UO_1004 (O_1004,N_8172,N_9463);
and UO_1005 (O_1005,N_8215,N_9652);
nor UO_1006 (O_1006,N_8876,N_8646);
nor UO_1007 (O_1007,N_9480,N_9586);
or UO_1008 (O_1008,N_8028,N_9206);
or UO_1009 (O_1009,N_8366,N_8549);
nand UO_1010 (O_1010,N_8477,N_9779);
or UO_1011 (O_1011,N_8436,N_8112);
nand UO_1012 (O_1012,N_9345,N_8743);
nor UO_1013 (O_1013,N_9170,N_9004);
or UO_1014 (O_1014,N_9904,N_8564);
nor UO_1015 (O_1015,N_8209,N_8824);
nand UO_1016 (O_1016,N_9017,N_9456);
nand UO_1017 (O_1017,N_9395,N_8529);
and UO_1018 (O_1018,N_9527,N_8754);
nand UO_1019 (O_1019,N_9019,N_9143);
or UO_1020 (O_1020,N_9251,N_8013);
nand UO_1021 (O_1021,N_9975,N_8124);
nand UO_1022 (O_1022,N_8824,N_8771);
and UO_1023 (O_1023,N_8259,N_8898);
or UO_1024 (O_1024,N_9807,N_9112);
and UO_1025 (O_1025,N_9298,N_8338);
and UO_1026 (O_1026,N_8637,N_9486);
nand UO_1027 (O_1027,N_8316,N_8676);
and UO_1028 (O_1028,N_9740,N_9750);
and UO_1029 (O_1029,N_8613,N_8234);
nor UO_1030 (O_1030,N_8727,N_9618);
nand UO_1031 (O_1031,N_8599,N_9467);
and UO_1032 (O_1032,N_8455,N_9024);
and UO_1033 (O_1033,N_9438,N_8377);
or UO_1034 (O_1034,N_9752,N_9695);
or UO_1035 (O_1035,N_9416,N_8752);
nor UO_1036 (O_1036,N_9942,N_9106);
nand UO_1037 (O_1037,N_9365,N_9537);
nand UO_1038 (O_1038,N_9620,N_9968);
nand UO_1039 (O_1039,N_9795,N_9061);
and UO_1040 (O_1040,N_9137,N_9078);
nor UO_1041 (O_1041,N_8485,N_8976);
or UO_1042 (O_1042,N_9524,N_8255);
nor UO_1043 (O_1043,N_8396,N_9657);
nand UO_1044 (O_1044,N_8559,N_8271);
or UO_1045 (O_1045,N_8230,N_8769);
nor UO_1046 (O_1046,N_9369,N_8315);
nor UO_1047 (O_1047,N_9637,N_8492);
or UO_1048 (O_1048,N_9513,N_8235);
or UO_1049 (O_1049,N_9985,N_9993);
nand UO_1050 (O_1050,N_8672,N_9067);
nand UO_1051 (O_1051,N_8954,N_9961);
and UO_1052 (O_1052,N_8600,N_9300);
nor UO_1053 (O_1053,N_9213,N_9166);
nor UO_1054 (O_1054,N_8137,N_8341);
or UO_1055 (O_1055,N_8231,N_9248);
nor UO_1056 (O_1056,N_8171,N_9025);
nand UO_1057 (O_1057,N_8346,N_9087);
or UO_1058 (O_1058,N_8282,N_9356);
and UO_1059 (O_1059,N_8500,N_9455);
nand UO_1060 (O_1060,N_9075,N_8926);
or UO_1061 (O_1061,N_8503,N_8291);
and UO_1062 (O_1062,N_8920,N_9734);
nand UO_1063 (O_1063,N_8625,N_9206);
and UO_1064 (O_1064,N_8148,N_8556);
nand UO_1065 (O_1065,N_9737,N_9648);
or UO_1066 (O_1066,N_9503,N_9487);
nand UO_1067 (O_1067,N_9050,N_8650);
nand UO_1068 (O_1068,N_8156,N_9988);
nand UO_1069 (O_1069,N_8207,N_8172);
or UO_1070 (O_1070,N_9642,N_9286);
or UO_1071 (O_1071,N_9123,N_8045);
xor UO_1072 (O_1072,N_8421,N_8539);
or UO_1073 (O_1073,N_9445,N_8026);
nand UO_1074 (O_1074,N_9757,N_9825);
nand UO_1075 (O_1075,N_9008,N_8470);
nor UO_1076 (O_1076,N_8696,N_9902);
or UO_1077 (O_1077,N_9677,N_9670);
or UO_1078 (O_1078,N_9309,N_8330);
and UO_1079 (O_1079,N_8101,N_9593);
and UO_1080 (O_1080,N_8646,N_8642);
or UO_1081 (O_1081,N_8875,N_9295);
and UO_1082 (O_1082,N_9855,N_8647);
nor UO_1083 (O_1083,N_8244,N_8851);
or UO_1084 (O_1084,N_8257,N_9906);
or UO_1085 (O_1085,N_8417,N_8834);
nand UO_1086 (O_1086,N_9313,N_8554);
nand UO_1087 (O_1087,N_9360,N_9452);
and UO_1088 (O_1088,N_8417,N_9936);
or UO_1089 (O_1089,N_9875,N_9475);
and UO_1090 (O_1090,N_8950,N_8710);
nor UO_1091 (O_1091,N_9497,N_9188);
nand UO_1092 (O_1092,N_9881,N_9664);
nor UO_1093 (O_1093,N_9628,N_8596);
and UO_1094 (O_1094,N_8043,N_9768);
nor UO_1095 (O_1095,N_8713,N_9667);
or UO_1096 (O_1096,N_9204,N_8847);
and UO_1097 (O_1097,N_8242,N_9036);
nand UO_1098 (O_1098,N_8808,N_9133);
nor UO_1099 (O_1099,N_9861,N_9777);
or UO_1100 (O_1100,N_9534,N_8355);
nand UO_1101 (O_1101,N_8969,N_9572);
nor UO_1102 (O_1102,N_8946,N_8208);
nand UO_1103 (O_1103,N_8415,N_9287);
nor UO_1104 (O_1104,N_9229,N_9404);
nor UO_1105 (O_1105,N_9439,N_8797);
nand UO_1106 (O_1106,N_8682,N_8051);
nor UO_1107 (O_1107,N_9027,N_9603);
or UO_1108 (O_1108,N_9938,N_8932);
or UO_1109 (O_1109,N_8407,N_8975);
nand UO_1110 (O_1110,N_8091,N_9307);
nand UO_1111 (O_1111,N_8646,N_8484);
nor UO_1112 (O_1112,N_8258,N_9795);
nor UO_1113 (O_1113,N_9459,N_9972);
nor UO_1114 (O_1114,N_8576,N_8048);
and UO_1115 (O_1115,N_9251,N_9620);
nor UO_1116 (O_1116,N_9143,N_8987);
nor UO_1117 (O_1117,N_8104,N_9566);
nor UO_1118 (O_1118,N_8822,N_9900);
or UO_1119 (O_1119,N_9542,N_8783);
or UO_1120 (O_1120,N_8905,N_9481);
nor UO_1121 (O_1121,N_8303,N_9660);
or UO_1122 (O_1122,N_9581,N_8477);
and UO_1123 (O_1123,N_8595,N_9075);
nor UO_1124 (O_1124,N_9592,N_8251);
xnor UO_1125 (O_1125,N_9394,N_9170);
nor UO_1126 (O_1126,N_9546,N_8480);
and UO_1127 (O_1127,N_9666,N_8335);
or UO_1128 (O_1128,N_9546,N_9964);
or UO_1129 (O_1129,N_9221,N_9200);
nor UO_1130 (O_1130,N_8511,N_9824);
nor UO_1131 (O_1131,N_9836,N_9566);
nor UO_1132 (O_1132,N_9197,N_9122);
nand UO_1133 (O_1133,N_8640,N_8450);
or UO_1134 (O_1134,N_9146,N_9967);
and UO_1135 (O_1135,N_9103,N_8832);
or UO_1136 (O_1136,N_8206,N_9710);
nand UO_1137 (O_1137,N_9817,N_9986);
nand UO_1138 (O_1138,N_8515,N_9903);
nor UO_1139 (O_1139,N_9311,N_9537);
nor UO_1140 (O_1140,N_9317,N_9424);
or UO_1141 (O_1141,N_8429,N_9027);
nand UO_1142 (O_1142,N_8162,N_8368);
and UO_1143 (O_1143,N_9114,N_9106);
nor UO_1144 (O_1144,N_8446,N_8740);
and UO_1145 (O_1145,N_8269,N_9124);
nand UO_1146 (O_1146,N_8593,N_8439);
nor UO_1147 (O_1147,N_9419,N_8205);
and UO_1148 (O_1148,N_9159,N_8418);
or UO_1149 (O_1149,N_8362,N_9572);
nor UO_1150 (O_1150,N_9888,N_9741);
and UO_1151 (O_1151,N_9246,N_8294);
and UO_1152 (O_1152,N_8912,N_8105);
and UO_1153 (O_1153,N_8451,N_9095);
and UO_1154 (O_1154,N_8055,N_8223);
and UO_1155 (O_1155,N_8550,N_9575);
nand UO_1156 (O_1156,N_9920,N_9309);
nor UO_1157 (O_1157,N_9135,N_9217);
nand UO_1158 (O_1158,N_8740,N_8368);
nand UO_1159 (O_1159,N_8848,N_9358);
nand UO_1160 (O_1160,N_9297,N_9061);
and UO_1161 (O_1161,N_8914,N_9461);
nand UO_1162 (O_1162,N_9593,N_9561);
and UO_1163 (O_1163,N_8452,N_9672);
nand UO_1164 (O_1164,N_8053,N_8206);
and UO_1165 (O_1165,N_9450,N_9199);
and UO_1166 (O_1166,N_8588,N_8435);
nor UO_1167 (O_1167,N_9227,N_9897);
and UO_1168 (O_1168,N_8763,N_8368);
nand UO_1169 (O_1169,N_8971,N_9930);
or UO_1170 (O_1170,N_8669,N_9686);
nor UO_1171 (O_1171,N_8818,N_8767);
nor UO_1172 (O_1172,N_8762,N_9719);
nor UO_1173 (O_1173,N_8760,N_8051);
nand UO_1174 (O_1174,N_8388,N_9194);
or UO_1175 (O_1175,N_8983,N_9594);
and UO_1176 (O_1176,N_9736,N_9636);
nor UO_1177 (O_1177,N_8850,N_8706);
and UO_1178 (O_1178,N_8224,N_8308);
nor UO_1179 (O_1179,N_8735,N_9675);
or UO_1180 (O_1180,N_8783,N_8961);
or UO_1181 (O_1181,N_9000,N_9583);
or UO_1182 (O_1182,N_8825,N_8066);
nand UO_1183 (O_1183,N_9951,N_8579);
or UO_1184 (O_1184,N_9668,N_9860);
nand UO_1185 (O_1185,N_8704,N_9497);
and UO_1186 (O_1186,N_8299,N_9914);
or UO_1187 (O_1187,N_8898,N_9111);
and UO_1188 (O_1188,N_9101,N_9881);
nor UO_1189 (O_1189,N_9499,N_8704);
nand UO_1190 (O_1190,N_9783,N_8736);
nor UO_1191 (O_1191,N_8850,N_8199);
nor UO_1192 (O_1192,N_9775,N_8246);
nor UO_1193 (O_1193,N_9316,N_9870);
nor UO_1194 (O_1194,N_8018,N_9456);
nand UO_1195 (O_1195,N_8274,N_8685);
or UO_1196 (O_1196,N_9783,N_8858);
or UO_1197 (O_1197,N_8180,N_9182);
nor UO_1198 (O_1198,N_9534,N_8367);
nand UO_1199 (O_1199,N_9859,N_9809);
or UO_1200 (O_1200,N_9873,N_8538);
nor UO_1201 (O_1201,N_9189,N_8868);
nand UO_1202 (O_1202,N_9269,N_8165);
nand UO_1203 (O_1203,N_9045,N_9979);
nor UO_1204 (O_1204,N_9651,N_9349);
nor UO_1205 (O_1205,N_8786,N_8612);
nor UO_1206 (O_1206,N_8449,N_8851);
and UO_1207 (O_1207,N_8388,N_9209);
nor UO_1208 (O_1208,N_8063,N_9828);
nand UO_1209 (O_1209,N_9021,N_9002);
and UO_1210 (O_1210,N_9624,N_8502);
or UO_1211 (O_1211,N_9722,N_8632);
nand UO_1212 (O_1212,N_9608,N_8377);
xor UO_1213 (O_1213,N_9506,N_9459);
nand UO_1214 (O_1214,N_8010,N_9110);
and UO_1215 (O_1215,N_9913,N_8283);
or UO_1216 (O_1216,N_8403,N_9625);
and UO_1217 (O_1217,N_9305,N_9242);
nand UO_1218 (O_1218,N_8729,N_8270);
nor UO_1219 (O_1219,N_8123,N_8958);
or UO_1220 (O_1220,N_8216,N_9152);
nor UO_1221 (O_1221,N_8179,N_9118);
or UO_1222 (O_1222,N_9447,N_9098);
nand UO_1223 (O_1223,N_9806,N_9932);
nor UO_1224 (O_1224,N_8983,N_9282);
nor UO_1225 (O_1225,N_9096,N_8214);
nand UO_1226 (O_1226,N_8559,N_9297);
and UO_1227 (O_1227,N_8353,N_8591);
and UO_1228 (O_1228,N_8114,N_8380);
nand UO_1229 (O_1229,N_8780,N_8428);
nor UO_1230 (O_1230,N_8036,N_8620);
or UO_1231 (O_1231,N_9547,N_9051);
or UO_1232 (O_1232,N_9241,N_9660);
or UO_1233 (O_1233,N_8717,N_9105);
nand UO_1234 (O_1234,N_9887,N_9279);
and UO_1235 (O_1235,N_9050,N_9399);
nor UO_1236 (O_1236,N_8843,N_9401);
and UO_1237 (O_1237,N_8843,N_9146);
and UO_1238 (O_1238,N_9707,N_8517);
nor UO_1239 (O_1239,N_8535,N_9836);
nand UO_1240 (O_1240,N_8035,N_8628);
nand UO_1241 (O_1241,N_9463,N_8804);
or UO_1242 (O_1242,N_9289,N_8557);
nand UO_1243 (O_1243,N_9678,N_9864);
nand UO_1244 (O_1244,N_9533,N_8328);
and UO_1245 (O_1245,N_8571,N_9407);
and UO_1246 (O_1246,N_8431,N_8444);
nor UO_1247 (O_1247,N_9381,N_9484);
nor UO_1248 (O_1248,N_8609,N_9712);
nand UO_1249 (O_1249,N_9041,N_8907);
nor UO_1250 (O_1250,N_9536,N_9952);
xnor UO_1251 (O_1251,N_9817,N_8150);
or UO_1252 (O_1252,N_8313,N_9374);
nand UO_1253 (O_1253,N_9054,N_8820);
nand UO_1254 (O_1254,N_8934,N_8713);
or UO_1255 (O_1255,N_8303,N_8445);
nor UO_1256 (O_1256,N_9366,N_9299);
and UO_1257 (O_1257,N_9956,N_9536);
and UO_1258 (O_1258,N_9094,N_9261);
or UO_1259 (O_1259,N_9949,N_9010);
and UO_1260 (O_1260,N_9152,N_8635);
nand UO_1261 (O_1261,N_9671,N_8496);
or UO_1262 (O_1262,N_8958,N_9954);
or UO_1263 (O_1263,N_9790,N_8567);
nor UO_1264 (O_1264,N_9347,N_8721);
nor UO_1265 (O_1265,N_9858,N_9448);
or UO_1266 (O_1266,N_9768,N_8450);
and UO_1267 (O_1267,N_9479,N_9040);
or UO_1268 (O_1268,N_9501,N_8593);
or UO_1269 (O_1269,N_9504,N_9758);
and UO_1270 (O_1270,N_8995,N_9292);
and UO_1271 (O_1271,N_9589,N_8987);
nand UO_1272 (O_1272,N_9360,N_8055);
or UO_1273 (O_1273,N_9564,N_9997);
nand UO_1274 (O_1274,N_9251,N_9401);
nor UO_1275 (O_1275,N_9245,N_9935);
or UO_1276 (O_1276,N_8119,N_9290);
and UO_1277 (O_1277,N_9242,N_8712);
or UO_1278 (O_1278,N_9914,N_8652);
or UO_1279 (O_1279,N_9645,N_9724);
nor UO_1280 (O_1280,N_9369,N_8123);
nand UO_1281 (O_1281,N_9628,N_9061);
or UO_1282 (O_1282,N_9037,N_8491);
nand UO_1283 (O_1283,N_8689,N_8239);
nor UO_1284 (O_1284,N_8755,N_8939);
or UO_1285 (O_1285,N_9506,N_9895);
nand UO_1286 (O_1286,N_9613,N_8613);
or UO_1287 (O_1287,N_9898,N_8271);
nor UO_1288 (O_1288,N_8061,N_9603);
nand UO_1289 (O_1289,N_8904,N_9578);
nand UO_1290 (O_1290,N_9205,N_9658);
and UO_1291 (O_1291,N_9977,N_9249);
nand UO_1292 (O_1292,N_9633,N_9751);
nand UO_1293 (O_1293,N_9437,N_8035);
nand UO_1294 (O_1294,N_8407,N_8661);
and UO_1295 (O_1295,N_8252,N_9384);
or UO_1296 (O_1296,N_8725,N_8939);
nor UO_1297 (O_1297,N_8382,N_9525);
or UO_1298 (O_1298,N_9417,N_8321);
and UO_1299 (O_1299,N_8153,N_9366);
nand UO_1300 (O_1300,N_9830,N_9255);
or UO_1301 (O_1301,N_8600,N_9002);
and UO_1302 (O_1302,N_9001,N_8689);
nand UO_1303 (O_1303,N_9489,N_8380);
and UO_1304 (O_1304,N_8852,N_8718);
or UO_1305 (O_1305,N_8108,N_8133);
or UO_1306 (O_1306,N_9811,N_8982);
and UO_1307 (O_1307,N_8182,N_8737);
and UO_1308 (O_1308,N_9229,N_9271);
and UO_1309 (O_1309,N_8830,N_9393);
nand UO_1310 (O_1310,N_8668,N_9506);
nand UO_1311 (O_1311,N_8125,N_8712);
nand UO_1312 (O_1312,N_9426,N_9354);
or UO_1313 (O_1313,N_9117,N_9498);
and UO_1314 (O_1314,N_9715,N_8670);
nor UO_1315 (O_1315,N_8041,N_9789);
or UO_1316 (O_1316,N_8364,N_8776);
or UO_1317 (O_1317,N_8694,N_9083);
or UO_1318 (O_1318,N_9216,N_9318);
or UO_1319 (O_1319,N_8659,N_9572);
nor UO_1320 (O_1320,N_8765,N_8910);
nand UO_1321 (O_1321,N_9159,N_8367);
or UO_1322 (O_1322,N_8347,N_8764);
or UO_1323 (O_1323,N_8696,N_9758);
or UO_1324 (O_1324,N_9268,N_8441);
nand UO_1325 (O_1325,N_9494,N_9222);
and UO_1326 (O_1326,N_8068,N_9801);
nor UO_1327 (O_1327,N_9428,N_9219);
or UO_1328 (O_1328,N_9694,N_8202);
or UO_1329 (O_1329,N_8862,N_9736);
nor UO_1330 (O_1330,N_8235,N_8451);
nand UO_1331 (O_1331,N_8973,N_8674);
nor UO_1332 (O_1332,N_8965,N_9769);
nand UO_1333 (O_1333,N_8603,N_9613);
or UO_1334 (O_1334,N_9981,N_8203);
nor UO_1335 (O_1335,N_9348,N_9881);
nand UO_1336 (O_1336,N_8249,N_8520);
and UO_1337 (O_1337,N_8120,N_9553);
or UO_1338 (O_1338,N_9851,N_8667);
or UO_1339 (O_1339,N_9528,N_8141);
nor UO_1340 (O_1340,N_9603,N_8541);
and UO_1341 (O_1341,N_8911,N_8197);
and UO_1342 (O_1342,N_9403,N_9755);
or UO_1343 (O_1343,N_8094,N_8320);
nor UO_1344 (O_1344,N_8962,N_8583);
and UO_1345 (O_1345,N_9238,N_8137);
nor UO_1346 (O_1346,N_8976,N_9338);
nor UO_1347 (O_1347,N_9604,N_8582);
and UO_1348 (O_1348,N_8540,N_8494);
nor UO_1349 (O_1349,N_9800,N_9454);
nor UO_1350 (O_1350,N_8248,N_8052);
nand UO_1351 (O_1351,N_9465,N_9617);
or UO_1352 (O_1352,N_8034,N_9979);
and UO_1353 (O_1353,N_8387,N_9836);
or UO_1354 (O_1354,N_8038,N_8868);
nand UO_1355 (O_1355,N_8124,N_9421);
nand UO_1356 (O_1356,N_8802,N_9823);
and UO_1357 (O_1357,N_8432,N_8315);
or UO_1358 (O_1358,N_9549,N_8436);
or UO_1359 (O_1359,N_9757,N_8785);
nand UO_1360 (O_1360,N_8446,N_8686);
and UO_1361 (O_1361,N_8759,N_9575);
or UO_1362 (O_1362,N_8655,N_9775);
or UO_1363 (O_1363,N_8720,N_9279);
nor UO_1364 (O_1364,N_8488,N_9485);
nand UO_1365 (O_1365,N_8115,N_9172);
and UO_1366 (O_1366,N_8974,N_9424);
nand UO_1367 (O_1367,N_8742,N_9506);
nand UO_1368 (O_1368,N_8191,N_9417);
nor UO_1369 (O_1369,N_8516,N_9385);
and UO_1370 (O_1370,N_9386,N_8693);
nor UO_1371 (O_1371,N_8490,N_8564);
and UO_1372 (O_1372,N_9581,N_8495);
nor UO_1373 (O_1373,N_8000,N_9188);
or UO_1374 (O_1374,N_9020,N_8690);
nand UO_1375 (O_1375,N_9570,N_8513);
or UO_1376 (O_1376,N_9515,N_9473);
nor UO_1377 (O_1377,N_8349,N_9313);
or UO_1378 (O_1378,N_9581,N_9990);
nand UO_1379 (O_1379,N_9264,N_9810);
or UO_1380 (O_1380,N_8883,N_9012);
or UO_1381 (O_1381,N_8417,N_8720);
or UO_1382 (O_1382,N_8627,N_9626);
nand UO_1383 (O_1383,N_9616,N_8370);
nand UO_1384 (O_1384,N_9676,N_9281);
and UO_1385 (O_1385,N_9282,N_9543);
or UO_1386 (O_1386,N_8923,N_9947);
or UO_1387 (O_1387,N_9959,N_9187);
nand UO_1388 (O_1388,N_9338,N_8470);
and UO_1389 (O_1389,N_8328,N_9231);
nor UO_1390 (O_1390,N_8368,N_9070);
and UO_1391 (O_1391,N_9403,N_9140);
or UO_1392 (O_1392,N_8847,N_8850);
or UO_1393 (O_1393,N_9786,N_9575);
and UO_1394 (O_1394,N_8218,N_8095);
and UO_1395 (O_1395,N_8960,N_8193);
or UO_1396 (O_1396,N_8189,N_8289);
or UO_1397 (O_1397,N_8742,N_8849);
or UO_1398 (O_1398,N_8155,N_8151);
nor UO_1399 (O_1399,N_8701,N_9468);
and UO_1400 (O_1400,N_9293,N_8167);
and UO_1401 (O_1401,N_8442,N_9285);
xor UO_1402 (O_1402,N_8679,N_9375);
and UO_1403 (O_1403,N_8200,N_8928);
and UO_1404 (O_1404,N_8646,N_8462);
nand UO_1405 (O_1405,N_8821,N_8750);
nor UO_1406 (O_1406,N_8843,N_8748);
or UO_1407 (O_1407,N_9855,N_8095);
or UO_1408 (O_1408,N_9493,N_8783);
nor UO_1409 (O_1409,N_8628,N_9181);
nand UO_1410 (O_1410,N_8174,N_8253);
nor UO_1411 (O_1411,N_8793,N_8136);
nor UO_1412 (O_1412,N_9545,N_9106);
or UO_1413 (O_1413,N_9280,N_8391);
nand UO_1414 (O_1414,N_9060,N_8426);
nor UO_1415 (O_1415,N_9744,N_9786);
nor UO_1416 (O_1416,N_8019,N_9433);
nand UO_1417 (O_1417,N_8561,N_8374);
and UO_1418 (O_1418,N_9137,N_9460);
nand UO_1419 (O_1419,N_9568,N_9997);
or UO_1420 (O_1420,N_8553,N_8230);
nor UO_1421 (O_1421,N_8654,N_8317);
nand UO_1422 (O_1422,N_8610,N_9835);
nand UO_1423 (O_1423,N_9765,N_8717);
xor UO_1424 (O_1424,N_8788,N_9295);
nand UO_1425 (O_1425,N_8035,N_9787);
and UO_1426 (O_1426,N_9132,N_9341);
nand UO_1427 (O_1427,N_9265,N_8405);
nand UO_1428 (O_1428,N_8900,N_9102);
nand UO_1429 (O_1429,N_9980,N_9662);
and UO_1430 (O_1430,N_8923,N_8677);
and UO_1431 (O_1431,N_8357,N_8091);
xor UO_1432 (O_1432,N_8065,N_9423);
or UO_1433 (O_1433,N_9375,N_9558);
nand UO_1434 (O_1434,N_8136,N_9214);
or UO_1435 (O_1435,N_9239,N_9023);
nor UO_1436 (O_1436,N_8458,N_8840);
nor UO_1437 (O_1437,N_9666,N_8905);
nor UO_1438 (O_1438,N_8609,N_9858);
and UO_1439 (O_1439,N_8371,N_9218);
and UO_1440 (O_1440,N_8162,N_9930);
and UO_1441 (O_1441,N_8395,N_9722);
or UO_1442 (O_1442,N_8271,N_9490);
nor UO_1443 (O_1443,N_8209,N_8426);
or UO_1444 (O_1444,N_8551,N_9203);
nor UO_1445 (O_1445,N_9094,N_8505);
or UO_1446 (O_1446,N_9895,N_9466);
or UO_1447 (O_1447,N_9694,N_9804);
nor UO_1448 (O_1448,N_8017,N_9955);
nor UO_1449 (O_1449,N_8255,N_9786);
or UO_1450 (O_1450,N_9832,N_9267);
nand UO_1451 (O_1451,N_8798,N_8612);
nand UO_1452 (O_1452,N_8391,N_8213);
and UO_1453 (O_1453,N_8632,N_8909);
or UO_1454 (O_1454,N_8756,N_8923);
and UO_1455 (O_1455,N_8611,N_8901);
nor UO_1456 (O_1456,N_9194,N_9265);
and UO_1457 (O_1457,N_9346,N_8349);
and UO_1458 (O_1458,N_8326,N_9352);
xnor UO_1459 (O_1459,N_9792,N_8503);
nor UO_1460 (O_1460,N_9827,N_9246);
or UO_1461 (O_1461,N_8787,N_9276);
nor UO_1462 (O_1462,N_8777,N_9203);
nor UO_1463 (O_1463,N_9148,N_9079);
or UO_1464 (O_1464,N_8621,N_8610);
nand UO_1465 (O_1465,N_8859,N_8388);
or UO_1466 (O_1466,N_8974,N_8744);
and UO_1467 (O_1467,N_8870,N_8223);
nand UO_1468 (O_1468,N_8535,N_9106);
nor UO_1469 (O_1469,N_8323,N_8448);
nor UO_1470 (O_1470,N_9377,N_9375);
or UO_1471 (O_1471,N_8331,N_9971);
or UO_1472 (O_1472,N_9130,N_8856);
and UO_1473 (O_1473,N_9405,N_9720);
nor UO_1474 (O_1474,N_8416,N_8433);
nor UO_1475 (O_1475,N_8158,N_8540);
nand UO_1476 (O_1476,N_9406,N_8424);
or UO_1477 (O_1477,N_9755,N_8431);
or UO_1478 (O_1478,N_8859,N_8041);
and UO_1479 (O_1479,N_9041,N_9518);
nand UO_1480 (O_1480,N_8496,N_9599);
nor UO_1481 (O_1481,N_8988,N_9067);
nor UO_1482 (O_1482,N_8713,N_8656);
or UO_1483 (O_1483,N_9013,N_9382);
nand UO_1484 (O_1484,N_8186,N_9166);
or UO_1485 (O_1485,N_8411,N_9341);
and UO_1486 (O_1486,N_9813,N_8702);
and UO_1487 (O_1487,N_8928,N_9260);
and UO_1488 (O_1488,N_8834,N_9160);
or UO_1489 (O_1489,N_8895,N_9861);
nand UO_1490 (O_1490,N_9020,N_8230);
or UO_1491 (O_1491,N_9223,N_9227);
nand UO_1492 (O_1492,N_9328,N_8899);
and UO_1493 (O_1493,N_8435,N_8587);
or UO_1494 (O_1494,N_9319,N_8613);
nand UO_1495 (O_1495,N_9251,N_8969);
nor UO_1496 (O_1496,N_9223,N_8990);
and UO_1497 (O_1497,N_8949,N_8992);
or UO_1498 (O_1498,N_9344,N_8275);
nor UO_1499 (O_1499,N_9457,N_9367);
endmodule